module basic_2500_25000_3000_4_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18935,N_18936,N_18937,N_18938,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19024,N_19025,N_19026,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19076,N_19077,N_19078,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19412,N_19413,N_19414,N_19415,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19600,N_19602,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19623,N_19624,N_19625,N_19626,N_19628,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19787,N_19788,N_19789,N_19790,N_19791,N_19793,N_19794,N_19795,N_19796,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19907,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20168,N_20169,N_20170,N_20171,N_20172,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20210,N_20211,N_20212,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20865,N_20867,N_20868,N_20870,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21060,N_21061,N_21062,N_21063,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21127,N_21128,N_21129,N_21130,N_21131,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21205,N_21206,N_21207,N_21208,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21364,N_21365,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21735,N_21736,N_21737,N_21738,N_21739,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21748,N_21749,N_21750,N_21751,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21798,N_21799,N_21800,N_21801,N_21802,N_21804,N_21805,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21962,N_21963,N_21964,N_21965,N_21967,N_21968,N_21969,N_21970,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22170,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22267,N_22268,N_22269,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22405,N_22406,N_22407,N_22408,N_22410,N_22411,N_22412,N_22414,N_22415,N_22416,N_22417,N_22418,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22447,N_22448,N_22449,N_22450,N_22451,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22498,N_22499,N_22500,N_22501,N_22502,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22681,N_22682,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22971,N_22972,N_22973,N_22974,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23251,N_23252,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23286,N_23287,N_23288,N_23289,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23326,N_23327,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23431,N_23432,N_23433,N_23434,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23516,N_23517,N_23518,N_23519,N_23521,N_23522,N_23523,N_23524,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24188,N_24189,N_24190,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24223,N_24224,N_24225,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24532,N_24533,N_24534,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24552,N_24553,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24582,N_24583,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24959,N_24960,N_24961,N_24962,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998;
nand U0 (N_0,In_1376,In_267);
nor U1 (N_1,In_610,In_268);
xor U2 (N_2,In_1160,In_1334);
or U3 (N_3,In_272,In_1758);
nor U4 (N_4,In_2109,In_2408);
and U5 (N_5,In_790,In_1071);
and U6 (N_6,In_882,In_943);
or U7 (N_7,In_2240,In_257);
nand U8 (N_8,In_2200,In_2445);
xnor U9 (N_9,In_180,In_1797);
and U10 (N_10,In_710,In_1668);
or U11 (N_11,In_2428,In_477);
nand U12 (N_12,In_2104,In_1685);
or U13 (N_13,In_1875,In_1229);
xnor U14 (N_14,In_1741,In_2176);
or U15 (N_15,In_766,In_2482);
nand U16 (N_16,In_2019,In_1426);
or U17 (N_17,In_701,In_1844);
and U18 (N_18,In_826,In_2301);
nor U19 (N_19,In_1309,In_1399);
nand U20 (N_20,In_2426,In_2323);
xnor U21 (N_21,In_193,In_2497);
xor U22 (N_22,In_577,In_2233);
nand U23 (N_23,In_630,In_437);
nand U24 (N_24,In_1020,In_217);
or U25 (N_25,In_2366,In_2364);
nor U26 (N_26,In_467,In_1582);
xnor U27 (N_27,In_1489,In_445);
or U28 (N_28,In_1450,In_874);
and U29 (N_29,In_612,In_1626);
or U30 (N_30,In_2272,In_672);
or U31 (N_31,In_768,In_1266);
and U32 (N_32,In_1834,In_512);
or U33 (N_33,In_744,In_136);
and U34 (N_34,In_2420,In_1500);
xor U35 (N_35,In_1195,In_2419);
nor U36 (N_36,In_2477,In_165);
or U37 (N_37,In_1038,In_533);
xnor U38 (N_38,In_1134,In_2368);
nand U39 (N_39,In_2441,In_1287);
xnor U40 (N_40,In_2444,In_434);
or U41 (N_41,In_667,In_1454);
nor U42 (N_42,In_1833,In_671);
nor U43 (N_43,In_2250,In_849);
nor U44 (N_44,In_1567,In_461);
nand U45 (N_45,In_572,In_100);
nand U46 (N_46,In_604,In_1885);
or U47 (N_47,In_2427,In_448);
or U48 (N_48,In_2094,In_1724);
or U49 (N_49,In_1164,In_1107);
nand U50 (N_50,In_10,In_704);
or U51 (N_51,In_651,In_236);
or U52 (N_52,In_760,In_1536);
xor U53 (N_53,In_1416,In_812);
and U54 (N_54,In_2350,In_1637);
nor U55 (N_55,In_1288,In_1609);
xnor U56 (N_56,In_989,In_1005);
xnor U57 (N_57,In_739,In_947);
and U58 (N_58,In_1186,In_631);
xor U59 (N_59,In_639,In_1417);
or U60 (N_60,In_775,In_195);
nand U61 (N_61,In_780,In_753);
nand U62 (N_62,In_1520,In_2300);
and U63 (N_63,In_1806,In_147);
and U64 (N_64,In_404,In_2005);
xnor U65 (N_65,In_728,In_2378);
and U66 (N_66,In_1613,In_1838);
nor U67 (N_67,In_107,In_1383);
xnor U68 (N_68,In_2040,In_1384);
and U69 (N_69,In_1608,In_2479);
nor U70 (N_70,In_1854,In_465);
nor U71 (N_71,In_441,In_2412);
xor U72 (N_72,In_1277,In_2084);
xnor U73 (N_73,In_1678,In_1720);
or U74 (N_74,In_1718,In_1088);
and U75 (N_75,In_1174,In_1996);
xnor U76 (N_76,In_61,In_212);
nor U77 (N_77,In_749,In_2192);
xnor U78 (N_78,In_2168,In_1397);
and U79 (N_79,In_1717,In_2133);
and U80 (N_80,In_718,In_1605);
nor U81 (N_81,In_1433,In_488);
or U82 (N_82,In_65,In_2145);
or U83 (N_83,In_1377,In_603);
xnor U84 (N_84,In_9,In_2173);
nor U85 (N_85,In_1056,In_618);
or U86 (N_86,In_620,In_1335);
and U87 (N_87,In_1872,In_93);
and U88 (N_88,In_14,In_647);
nor U89 (N_89,In_1575,In_2373);
xnor U90 (N_90,In_1201,In_1727);
xor U91 (N_91,In_1460,In_1736);
nor U92 (N_92,In_2238,In_2032);
nor U93 (N_93,In_2248,In_1853);
nor U94 (N_94,In_978,In_872);
and U95 (N_95,In_2092,In_1901);
and U96 (N_96,In_1928,In_1580);
and U97 (N_97,In_1480,In_1658);
and U98 (N_98,In_929,In_52);
nand U99 (N_99,In_997,In_1369);
and U100 (N_100,In_820,In_1595);
and U101 (N_101,In_712,In_540);
nor U102 (N_102,In_1802,In_1703);
or U103 (N_103,In_164,In_1324);
xnor U104 (N_104,In_506,In_2020);
nor U105 (N_105,In_11,In_956);
and U106 (N_106,In_931,In_1294);
nor U107 (N_107,In_135,In_1991);
xnor U108 (N_108,In_19,In_88);
or U109 (N_109,In_412,In_421);
or U110 (N_110,In_991,In_178);
xor U111 (N_111,In_1654,In_1221);
or U112 (N_112,In_1856,In_132);
or U113 (N_113,In_1765,In_411);
and U114 (N_114,In_1541,In_1624);
nand U115 (N_115,In_853,In_748);
nor U116 (N_116,In_582,In_414);
nand U117 (N_117,In_764,In_1601);
or U118 (N_118,In_1869,In_288);
or U119 (N_119,In_1400,In_115);
or U120 (N_120,In_1864,In_1877);
xnor U121 (N_121,In_2421,In_2202);
and U122 (N_122,In_525,In_1262);
nor U123 (N_123,In_2338,In_648);
xor U124 (N_124,In_703,In_2181);
and U125 (N_125,In_1213,In_2125);
nor U126 (N_126,In_1126,In_1919);
nor U127 (N_127,In_1968,In_2050);
nor U128 (N_128,In_2,In_811);
nor U129 (N_129,In_677,In_139);
or U130 (N_130,In_1322,In_1403);
xor U131 (N_131,In_20,In_1625);
xnor U132 (N_132,In_1807,In_1546);
nand U133 (N_133,In_1503,In_2186);
nor U134 (N_134,In_1990,In_2322);
xnor U135 (N_135,In_1175,In_646);
nand U136 (N_136,In_1822,In_1731);
xor U137 (N_137,In_863,In_1574);
or U138 (N_138,In_311,In_885);
and U139 (N_139,In_2253,In_1571);
nor U140 (N_140,In_1182,In_1540);
xor U141 (N_141,In_1616,In_487);
or U142 (N_142,In_711,In_659);
or U143 (N_143,In_299,In_291);
and U144 (N_144,In_963,In_2370);
nor U145 (N_145,In_1842,In_522);
xnor U146 (N_146,In_758,In_293);
nor U147 (N_147,In_1845,In_1451);
or U148 (N_148,In_755,In_1131);
nand U149 (N_149,In_1693,In_1803);
nor U150 (N_150,In_2470,In_541);
or U151 (N_151,In_190,In_786);
xnor U152 (N_152,In_1396,In_1315);
and U153 (N_153,In_1169,In_2351);
nor U154 (N_154,In_804,In_120);
nand U155 (N_155,In_296,In_407);
and U156 (N_156,In_355,In_420);
or U157 (N_157,In_568,In_2185);
or U158 (N_158,In_2078,In_2222);
xor U159 (N_159,In_211,In_726);
and U160 (N_160,In_206,In_1022);
or U161 (N_161,In_2073,In_301);
nor U162 (N_162,In_1095,In_317);
nand U163 (N_163,In_2262,In_59);
or U164 (N_164,In_449,In_71);
or U165 (N_165,In_1897,In_1830);
xor U166 (N_166,In_2226,In_1430);
or U167 (N_167,In_1677,In_208);
nand U168 (N_168,In_2483,In_1961);
or U169 (N_169,In_452,In_1326);
nor U170 (N_170,In_957,In_539);
or U171 (N_171,In_782,In_1860);
nor U172 (N_172,In_2435,In_968);
or U173 (N_173,In_2465,In_1255);
nand U174 (N_174,In_1237,In_2190);
or U175 (N_175,In_2027,In_2221);
nand U176 (N_176,In_1495,In_429);
xnor U177 (N_177,In_2362,In_1627);
nor U178 (N_178,In_1774,In_1332);
nor U179 (N_179,In_495,In_1336);
nand U180 (N_180,In_2052,In_1712);
and U181 (N_181,In_2007,In_2093);
nand U182 (N_182,In_737,In_96);
xnor U183 (N_183,In_413,In_2254);
xnor U184 (N_184,In_632,In_1463);
and U185 (N_185,In_1874,In_2402);
nand U186 (N_186,In_91,In_877);
nor U187 (N_187,In_1550,In_555);
nor U188 (N_188,In_1614,In_2360);
or U189 (N_189,In_1775,In_2212);
and U190 (N_190,In_1713,In_846);
or U191 (N_191,In_1032,In_468);
or U192 (N_192,In_891,In_2072);
nand U193 (N_193,In_1259,In_1445);
nand U194 (N_194,In_1374,In_1871);
nor U195 (N_195,In_312,In_593);
and U196 (N_196,In_779,In_1523);
or U197 (N_197,In_546,In_1346);
and U198 (N_198,In_2227,In_2228);
nor U199 (N_199,In_388,In_225);
and U200 (N_200,In_2009,In_1778);
or U201 (N_201,In_1344,In_1392);
or U202 (N_202,In_1225,In_1719);
xor U203 (N_203,In_1317,In_852);
or U204 (N_204,In_2180,In_1749);
and U205 (N_205,In_2275,In_2217);
nand U206 (N_206,In_975,In_218);
and U207 (N_207,In_376,In_490);
xor U208 (N_208,In_538,In_660);
nand U209 (N_209,In_600,In_2344);
xnor U210 (N_210,In_1795,In_273);
and U211 (N_211,In_650,In_1341);
nor U212 (N_212,In_2404,In_909);
xor U213 (N_213,In_365,In_1615);
or U214 (N_214,In_1528,In_1552);
and U215 (N_215,In_1069,In_860);
and U216 (N_216,In_1908,In_1849);
and U217 (N_217,In_2144,In_1880);
and U218 (N_218,In_1359,In_1440);
nand U219 (N_219,In_1436,In_1810);
nor U220 (N_220,In_867,In_1846);
and U221 (N_221,In_2423,In_606);
or U222 (N_222,In_2039,In_1618);
and U223 (N_223,In_2043,In_430);
xor U224 (N_224,In_2438,In_1178);
or U225 (N_225,In_150,In_1085);
nor U226 (N_226,In_1584,In_742);
or U227 (N_227,In_1339,In_1272);
nand U228 (N_228,In_1610,In_489);
nor U229 (N_229,In_1558,In_727);
and U230 (N_230,In_500,In_1380);
or U231 (N_231,In_1502,In_2156);
and U232 (N_232,In_2111,In_901);
and U233 (N_233,In_2236,In_2433);
xor U234 (N_234,In_824,In_591);
or U235 (N_235,In_1044,In_761);
nor U236 (N_236,In_2270,In_1027);
xnor U237 (N_237,In_431,In_274);
and U238 (N_238,In_282,In_2242);
nor U239 (N_239,In_2259,In_1192);
xor U240 (N_240,In_415,In_230);
xor U241 (N_241,In_1021,In_2401);
and U242 (N_242,In_2274,In_287);
and U243 (N_243,In_2127,In_1357);
and U244 (N_244,In_887,In_1282);
or U245 (N_245,In_474,In_941);
nand U246 (N_246,In_2225,In_1508);
nor U247 (N_247,In_1559,In_1010);
nand U248 (N_248,In_239,In_1941);
or U249 (N_249,In_2058,In_1406);
nand U250 (N_250,In_92,In_1239);
xnor U251 (N_251,In_1865,In_916);
xor U252 (N_252,In_1666,In_1870);
and U253 (N_253,In_2021,In_390);
or U254 (N_254,In_2055,In_558);
and U255 (N_255,In_141,In_1829);
and U256 (N_256,In_173,In_2167);
or U257 (N_257,In_1424,In_1475);
or U258 (N_258,In_810,In_2387);
nor U259 (N_259,In_1141,In_1114);
nand U260 (N_260,In_391,In_279);
or U261 (N_261,In_2237,In_1012);
xor U262 (N_262,In_203,In_1757);
xnor U263 (N_263,In_318,In_1222);
or U264 (N_264,In_1868,In_394);
and U265 (N_265,In_479,In_1078);
nor U266 (N_266,In_1443,In_2276);
nand U267 (N_267,In_1814,In_2099);
nand U268 (N_268,In_1112,In_2291);
or U269 (N_269,In_416,In_1123);
or U270 (N_270,In_1902,In_987);
nand U271 (N_271,In_484,In_2385);
nor U272 (N_272,In_2100,In_116);
nand U273 (N_273,In_194,In_1441);
nand U274 (N_274,In_2082,In_2067);
or U275 (N_275,In_2205,In_2008);
or U276 (N_276,In_1016,In_1240);
nor U277 (N_277,In_513,In_2393);
or U278 (N_278,In_866,In_1045);
nand U279 (N_279,In_2106,In_640);
nor U280 (N_280,In_2210,In_1375);
or U281 (N_281,In_1951,In_1136);
or U282 (N_282,In_1993,In_1997);
nand U283 (N_283,In_974,In_72);
and U284 (N_284,In_372,In_16);
or U285 (N_285,In_486,In_1548);
xnor U286 (N_286,In_30,In_470);
xnor U287 (N_287,In_1364,In_652);
nand U288 (N_288,In_1345,In_2048);
nand U289 (N_289,In_175,In_1825);
or U290 (N_290,In_386,In_472);
and U291 (N_291,In_324,In_63);
nor U292 (N_292,In_119,In_126);
xnor U293 (N_293,In_2462,In_1682);
nor U294 (N_294,In_1140,In_1799);
and U295 (N_295,In_39,In_585);
xnor U296 (N_296,In_2353,In_145);
xnor U297 (N_297,In_2391,In_1630);
or U298 (N_298,In_1563,In_532);
and U299 (N_299,In_1572,In_936);
xor U300 (N_300,In_314,In_2495);
nor U301 (N_301,In_396,In_155);
or U302 (N_302,In_1118,In_1210);
and U303 (N_303,In_1035,In_1894);
nor U304 (N_304,In_1385,In_2189);
and U305 (N_305,In_499,In_2498);
nor U306 (N_306,In_1779,In_966);
and U307 (N_307,In_2003,In_1623);
nand U308 (N_308,In_2273,In_436);
nand U309 (N_309,In_1776,In_1804);
nand U310 (N_310,In_1879,In_2339);
nor U311 (N_311,In_1269,In_1578);
and U312 (N_312,In_409,In_1931);
xor U313 (N_313,In_837,In_578);
or U314 (N_314,In_818,In_998);
nand U315 (N_315,In_1363,In_1181);
nor U316 (N_316,In_2386,In_1152);
nand U317 (N_317,In_913,In_142);
and U318 (N_318,In_520,In_1587);
nand U319 (N_319,In_1412,In_265);
or U320 (N_320,In_596,In_1120);
or U321 (N_321,In_156,In_215);
and U322 (N_322,In_2400,In_221);
and U323 (N_323,In_366,In_1543);
nand U324 (N_324,In_1947,In_839);
nor U325 (N_325,In_1596,In_1442);
nand U326 (N_326,In_1413,In_1808);
nor U327 (N_327,In_319,In_625);
and U328 (N_328,In_1236,In_378);
or U329 (N_329,In_1905,In_1862);
xnor U330 (N_330,In_861,In_1819);
and U331 (N_331,In_530,In_1672);
nor U332 (N_332,In_1890,In_833);
and U333 (N_333,In_90,In_2114);
nor U334 (N_334,In_224,In_759);
nand U335 (N_335,In_2436,In_2249);
or U336 (N_336,In_781,In_1809);
and U337 (N_337,In_329,In_334);
nor U338 (N_338,In_393,In_571);
or U339 (N_339,In_534,In_444);
nand U340 (N_340,In_2229,In_463);
nor U341 (N_341,In_1831,In_37);
and U342 (N_342,In_1135,In_1592);
and U343 (N_343,In_1937,In_1281);
xnor U344 (N_344,In_2329,In_1469);
or U345 (N_345,In_457,In_382);
nor U346 (N_346,In_2153,In_564);
or U347 (N_347,In_106,In_1292);
and U348 (N_348,In_1411,In_621);
xnor U349 (N_349,In_216,In_1057);
nor U350 (N_350,In_285,In_1594);
nand U351 (N_351,In_1629,In_447);
nand U352 (N_352,In_1318,In_800);
nand U353 (N_353,In_5,In_910);
nand U354 (N_354,In_1086,In_982);
or U355 (N_355,In_1093,In_1542);
or U356 (N_356,In_649,In_1952);
and U357 (N_357,In_1177,In_1545);
xnor U358 (N_358,In_517,In_439);
nor U359 (N_359,In_1137,In_1517);
nor U360 (N_360,In_1008,In_2247);
nor U361 (N_361,In_54,In_563);
nor U362 (N_362,In_1483,In_716);
and U363 (N_363,In_2284,In_1246);
and U364 (N_364,In_18,In_2407);
nor U365 (N_365,In_1052,In_2065);
nor U366 (N_366,In_2297,In_1063);
xnor U367 (N_367,In_140,In_1024);
or U368 (N_368,In_960,In_556);
or U369 (N_369,In_1402,In_1659);
nor U370 (N_370,In_1015,In_2054);
nand U371 (N_371,In_1832,In_2450);
xor U372 (N_372,In_1194,In_1168);
or U373 (N_373,In_774,In_478);
nor U374 (N_374,In_1461,In_617);
or U375 (N_375,In_398,In_1235);
nor U376 (N_376,In_2178,In_772);
nor U377 (N_377,In_2231,In_197);
nor U378 (N_378,In_904,In_49);
and U379 (N_379,In_1945,In_395);
xor U380 (N_380,In_903,In_2251);
and U381 (N_381,In_2484,In_246);
and U382 (N_382,In_1191,In_406);
nand U383 (N_383,In_2403,In_1171);
nor U384 (N_384,In_1496,In_1906);
or U385 (N_385,In_1922,In_1689);
nor U386 (N_386,In_2471,In_1547);
xor U387 (N_387,In_2266,In_961);
xor U388 (N_388,In_1766,In_501);
nor U389 (N_389,In_362,In_2416);
nand U390 (N_390,In_2463,In_1189);
or U391 (N_391,In_2460,In_1805);
nand U392 (N_392,In_1939,In_1458);
and U393 (N_393,In_167,In_1938);
nor U394 (N_394,In_953,In_454);
nor U395 (N_395,In_1007,In_2046);
nor U396 (N_396,In_1139,In_569);
and U397 (N_397,In_1102,In_33);
and U398 (N_398,In_553,In_2327);
nand U399 (N_399,In_109,In_1300);
nand U400 (N_400,In_907,In_1531);
or U401 (N_401,In_1072,In_276);
and U402 (N_402,In_973,In_1153);
or U403 (N_403,In_1661,In_746);
nor U404 (N_404,In_954,In_1600);
or U405 (N_405,In_1656,In_886);
nand U406 (N_406,In_580,In_0);
and U407 (N_407,In_2146,In_1509);
and U408 (N_408,In_504,In_2488);
and U409 (N_409,In_2234,In_1151);
or U410 (N_410,In_151,In_952);
and U411 (N_411,In_1641,In_423);
nand U412 (N_412,In_769,In_1167);
and U413 (N_413,In_2135,In_686);
xor U414 (N_414,In_432,In_1207);
xnor U415 (N_415,In_427,In_995);
or U416 (N_416,In_2278,In_2434);
nor U417 (N_417,In_349,In_552);
nor U418 (N_418,In_1821,In_127);
xor U419 (N_419,In_1964,In_1342);
nand U420 (N_420,In_834,In_1081);
nand U421 (N_421,In_1075,In_1042);
or U422 (N_422,In_1639,In_1188);
nor U423 (N_423,In_47,In_1067);
and U424 (N_424,In_1034,In_1728);
xnor U425 (N_425,In_1493,In_2295);
xnor U426 (N_426,In_2105,In_1549);
xor U427 (N_427,In_41,In_1234);
nor U428 (N_428,In_1681,In_1405);
or U429 (N_429,In_1455,In_12);
nor U430 (N_430,In_567,In_1539);
xor U431 (N_431,In_868,In_841);
xor U432 (N_432,In_2023,In_335);
and U433 (N_433,In_1013,In_1270);
nand U434 (N_434,In_1511,In_1092);
nor U435 (N_435,In_408,In_505);
xor U436 (N_436,In_1459,In_2367);
xor U437 (N_437,In_205,In_583);
nand U438 (N_438,In_1696,In_152);
nand U439 (N_439,In_923,In_2244);
and U440 (N_440,In_1187,In_401);
or U441 (N_441,In_374,In_777);
or U442 (N_442,In_2151,In_1017);
xnor U443 (N_443,In_1217,In_653);
nand U444 (N_444,In_1843,In_1476);
xnor U445 (N_445,In_1635,In_1570);
or U446 (N_446,In_1209,In_964);
xnor U447 (N_447,In_51,In_252);
xor U448 (N_448,In_1138,In_1491);
nor U449 (N_449,In_549,In_2321);
nand U450 (N_450,In_146,In_730);
and U451 (N_451,In_2045,In_524);
nor U452 (N_452,In_1710,In_985);
nand U453 (N_453,In_828,In_2493);
nor U454 (N_454,In_232,In_697);
nor U455 (N_455,In_1555,In_2036);
nor U456 (N_456,In_690,In_2429);
xor U457 (N_457,In_1740,In_1621);
and U458 (N_458,In_2203,In_1884);
and U459 (N_459,In_825,In_1488);
and U460 (N_460,In_247,In_707);
and U461 (N_461,In_566,In_1895);
and U462 (N_462,In_1647,In_25);
nand U463 (N_463,In_1915,In_1573);
nor U464 (N_464,In_2044,In_666);
nand U465 (N_465,In_1047,In_1735);
or U466 (N_466,In_482,In_1011);
nor U467 (N_467,In_1338,In_199);
nor U468 (N_468,In_2410,In_1473);
xor U469 (N_469,In_2143,In_1836);
and U470 (N_470,In_1053,In_2121);
nor U471 (N_471,In_1589,In_1598);
or U472 (N_472,In_68,In_1888);
or U473 (N_473,In_1204,In_2258);
or U474 (N_474,In_1242,In_2209);
nand U475 (N_475,In_1394,In_1859);
nor U476 (N_476,In_1887,In_658);
nand U477 (N_477,In_2457,In_1756);
and U478 (N_478,In_1663,In_871);
or U479 (N_479,In_1801,In_1307);
nand U480 (N_480,In_1506,In_1535);
nor U481 (N_481,In_363,In_1927);
or U482 (N_482,In_204,In_138);
or U483 (N_483,In_17,In_638);
nor U484 (N_484,In_519,In_2454);
or U485 (N_485,In_1470,In_696);
nand U486 (N_486,In_2208,In_1226);
nand U487 (N_487,In_958,In_1759);
or U488 (N_488,In_1839,In_361);
nor U489 (N_489,In_2383,In_969);
and U490 (N_490,In_2490,In_1427);
or U491 (N_491,In_2346,In_1366);
nand U492 (N_492,In_1699,In_627);
or U493 (N_493,In_1694,In_1704);
xnor U494 (N_494,In_392,In_1108);
xor U495 (N_495,In_2037,In_1328);
or U496 (N_496,In_2392,In_1590);
nand U497 (N_497,In_1068,In_1622);
nor U498 (N_498,In_1737,In_1122);
or U499 (N_499,In_2195,In_60);
xor U500 (N_500,In_2010,In_1505);
nor U501 (N_501,In_590,In_521);
xnor U502 (N_502,In_1127,In_1244);
nand U503 (N_503,In_300,In_1583);
xnor U504 (N_504,In_2431,In_817);
nand U505 (N_505,In_1428,In_1302);
xnor U506 (N_506,In_2069,In_2118);
nand U507 (N_507,In_1308,In_2224);
xor U508 (N_508,In_2316,In_1972);
or U509 (N_509,In_160,In_1079);
and U510 (N_510,In_543,In_2031);
or U511 (N_511,In_1636,In_1841);
nand U512 (N_512,In_1278,In_424);
nand U513 (N_513,In_2356,In_237);
and U514 (N_514,In_1373,In_1665);
and U515 (N_515,In_1899,In_636);
nand U516 (N_516,In_26,In_15);
and U517 (N_517,In_713,In_1049);
nand U518 (N_518,In_1331,In_2306);
nor U519 (N_519,In_641,In_7);
nor U520 (N_520,In_1132,In_1730);
nand U521 (N_521,In_1227,In_1003);
xnor U522 (N_522,In_1299,In_1247);
or U523 (N_523,In_428,In_937);
or U524 (N_524,In_2458,In_2241);
nand U525 (N_525,In_557,In_2096);
or U526 (N_526,In_453,In_575);
nor U527 (N_527,In_1564,In_767);
or U528 (N_528,In_614,In_1232);
and U529 (N_529,In_1419,In_1638);
or U530 (N_530,In_1984,In_1203);
and U531 (N_531,In_75,In_1914);
and U532 (N_532,In_2230,In_895);
nor U533 (N_533,In_1723,In_2365);
nand U534 (N_534,In_360,In_793);
xnor U535 (N_535,In_370,In_2310);
xnor U536 (N_536,In_1408,In_1918);
or U537 (N_537,In_341,In_900);
xor U538 (N_538,In_1319,In_400);
nand U539 (N_539,In_1023,In_367);
nand U540 (N_540,In_1347,In_229);
and U541 (N_541,In_1512,In_1599);
nor U542 (N_542,In_2331,In_21);
xnor U543 (N_543,In_383,In_1943);
and U544 (N_544,In_545,In_1125);
or U545 (N_545,In_305,In_1597);
or U546 (N_546,In_2349,In_1738);
and U547 (N_547,In_1208,In_2164);
nand U548 (N_548,In_1368,In_2219);
nand U549 (N_549,In_705,In_1286);
or U550 (N_550,In_698,In_128);
nand U551 (N_551,In_83,In_2455);
or U552 (N_552,In_1471,In_1429);
and U553 (N_553,In_1979,In_464);
and U554 (N_554,In_1848,In_2131);
nand U555 (N_555,In_785,In_2459);
xor U556 (N_556,In_562,In_1077);
xnor U557 (N_557,In_113,In_1401);
or U558 (N_558,In_309,In_1165);
xor U559 (N_559,In_1504,In_2424);
nand U560 (N_560,In_1688,In_896);
nor U561 (N_561,In_210,In_2080);
or U562 (N_562,In_356,In_570);
nand U563 (N_563,In_605,In_914);
xnor U564 (N_564,In_890,In_249);
and U565 (N_565,In_222,In_2481);
and U566 (N_566,In_1513,In_1031);
or U567 (N_567,In_121,In_1333);
and U568 (N_568,In_1781,In_1327);
xnor U569 (N_569,In_2000,In_70);
and U570 (N_570,In_359,In_2475);
xor U571 (N_571,In_337,In_1904);
nor U572 (N_572,In_1974,In_440);
xor U573 (N_573,In_48,In_323);
and U574 (N_574,In_1533,In_1812);
or U575 (N_575,In_1753,In_50);
nand U576 (N_576,In_674,In_2303);
and U577 (N_577,In_2439,In_1323);
or U578 (N_578,In_2359,In_2313);
nand U579 (N_579,In_635,In_2442);
and U580 (N_580,In_1019,In_1002);
nor U581 (N_581,In_1129,In_2187);
xnor U582 (N_582,In_2053,In_795);
nor U583 (N_583,In_1721,In_2290);
xor U584 (N_584,In_1372,In_1486);
nand U585 (N_585,In_770,In_202);
xor U586 (N_586,In_1387,In_2088);
or U587 (N_587,In_1645,In_2281);
nor U588 (N_588,In_657,In_2485);
nand U589 (N_589,In_548,In_2380);
and U590 (N_590,In_1527,In_1743);
or U591 (N_591,In_1569,In_27);
or U592 (N_592,In_2004,In_878);
nand U593 (N_593,In_816,In_784);
nand U594 (N_594,In_949,In_435);
nor U595 (N_595,In_1850,In_1263);
or U596 (N_596,In_1530,In_1407);
nand U597 (N_597,In_1867,In_1734);
and U598 (N_598,In_2026,In_628);
and U599 (N_599,In_1485,In_1708);
and U600 (N_600,In_1257,In_848);
nor U601 (N_601,In_2223,In_125);
xnor U602 (N_602,In_357,In_932);
xnor U603 (N_603,In_1726,In_446);
nor U604 (N_604,In_351,In_1390);
xnor U605 (N_605,In_1432,In_879);
nor U606 (N_606,In_1883,In_1041);
xor U607 (N_607,In_2279,In_1437);
nor U608 (N_608,In_1296,In_1274);
nor U609 (N_609,In_715,In_842);
nand U610 (N_610,In_771,In_220);
and U611 (N_611,In_656,In_2411);
xnor U612 (N_612,In_238,In_559);
or U613 (N_613,In_888,In_1691);
nor U614 (N_614,In_2396,In_1362);
and U615 (N_615,In_1790,In_214);
xnor U616 (N_616,In_251,In_494);
or U617 (N_617,In_1568,In_661);
nor U618 (N_618,In_322,In_1946);
nor U619 (N_619,In_2038,In_1130);
nor U620 (N_620,In_2204,In_241);
nand U621 (N_621,In_972,In_1218);
xor U622 (N_622,In_2174,In_2449);
xor U623 (N_623,In_1183,In_719);
nand U624 (N_624,In_1418,In_2070);
xnor U625 (N_625,In_801,In_283);
nor U626 (N_626,In_123,In_368);
and U627 (N_627,In_1611,In_69);
xnor U628 (N_628,In_192,In_1316);
or U629 (N_629,In_2018,In_1709);
and U630 (N_630,In_1456,In_1082);
nor U631 (N_631,In_231,In_1393);
and U632 (N_632,In_2478,In_516);
and U633 (N_633,In_1982,In_1907);
and U634 (N_634,In_1361,In_1930);
xnor U635 (N_635,In_223,In_1414);
nand U636 (N_636,In_1702,In_892);
or U637 (N_637,In_1644,In_2372);
nand U638 (N_638,In_1145,In_1791);
xnor U639 (N_639,In_384,In_1815);
and U640 (N_640,In_1190,In_971);
or U641 (N_641,In_1117,In_144);
xor U642 (N_642,In_2116,In_1422);
or U643 (N_643,In_794,In_1561);
nand U644 (N_644,In_1477,In_1722);
xnor U645 (N_645,In_765,In_1746);
nor U646 (N_646,In_2137,In_1421);
nor U647 (N_647,In_1748,In_78);
and U648 (N_648,In_1576,In_62);
xor U649 (N_649,In_668,In_942);
nand U650 (N_650,In_1811,In_1352);
nor U651 (N_651,In_2304,In_1415);
or U652 (N_652,In_2352,In_2013);
xor U653 (N_653,In_1275,In_364);
nor U654 (N_654,In_1097,In_1649);
and U655 (N_655,In_1462,In_2496);
and U656 (N_656,In_1510,In_1714);
xnor U657 (N_657,In_1763,In_2452);
xor U658 (N_658,In_1650,In_859);
xnor U659 (N_659,In_1917,In_1813);
xnor U660 (N_660,In_2057,In_1707);
nor U661 (N_661,In_2083,In_2134);
or U662 (N_662,In_622,In_97);
or U663 (N_663,In_920,In_1745);
and U664 (N_664,In_258,In_616);
and U665 (N_665,In_28,In_1881);
or U666 (N_666,In_1863,In_1004);
nand U667 (N_667,In_2399,In_831);
or U668 (N_668,In_1617,In_1925);
nor U669 (N_669,In_1976,In_425);
xnor U670 (N_670,In_921,In_1655);
nand U671 (N_671,In_22,In_598);
xor U672 (N_672,In_280,In_684);
nand U673 (N_673,In_528,In_762);
xnor U674 (N_674,In_665,In_2155);
and U675 (N_675,In_108,In_2294);
or U676 (N_676,In_845,In_2160);
nand U677 (N_677,In_321,In_1764);
or U678 (N_678,In_74,In_870);
or U679 (N_679,In_81,In_1690);
nand U680 (N_680,In_417,In_2172);
xnor U681 (N_681,In_1657,In_2271);
nand U682 (N_682,In_43,In_976);
nand U683 (N_683,In_53,In_1607);
nand U684 (N_684,In_1050,In_254);
nand U685 (N_685,In_1784,In_1264);
nor U686 (N_686,In_2169,In_980);
or U687 (N_687,In_798,In_1716);
and U688 (N_688,In_700,In_756);
or U689 (N_689,In_2206,In_333);
xnor U690 (N_690,In_1760,In_2193);
nand U691 (N_691,In_161,In_1310);
nor U692 (N_692,In_1942,In_1478);
and U693 (N_693,In_862,In_2309);
nand U694 (N_694,In_118,In_1431);
xor U695 (N_695,In_24,In_2071);
xor U696 (N_696,In_579,In_344);
and U697 (N_697,In_295,In_1566);
or U698 (N_698,In_788,In_2025);
nor U699 (N_699,In_58,In_2148);
and U700 (N_700,In_1783,In_912);
nor U701 (N_701,In_2371,In_476);
xor U702 (N_702,In_67,In_1184);
xnor U703 (N_703,In_181,In_945);
nand U704 (N_704,In_338,In_1230);
nand U705 (N_705,In_189,In_1211);
nand U706 (N_706,In_171,In_2467);
nand U707 (N_707,In_930,In_905);
nor U708 (N_708,In_1754,In_286);
nor U709 (N_709,In_259,In_1148);
nor U710 (N_710,In_992,In_399);
or U711 (N_711,In_881,In_455);
nand U712 (N_712,In_745,In_1116);
nor U713 (N_713,In_693,In_602);
xnor U714 (N_714,In_1579,In_1163);
xor U715 (N_715,In_763,In_469);
xnor U716 (N_716,In_1553,In_1816);
nor U717 (N_717,In_154,In_918);
nand U718 (N_718,In_1398,In_1284);
and U719 (N_719,In_645,In_1978);
nor U720 (N_720,In_1484,In_170);
nor U721 (N_721,In_1971,In_1761);
nand U722 (N_722,In_1143,In_460);
xnor U723 (N_723,In_1667,In_1981);
and U724 (N_724,In_2334,In_561);
xnor U725 (N_725,In_2162,In_948);
or U726 (N_726,In_1149,In_422);
nor U727 (N_727,In_2090,In_2140);
xor U728 (N_728,In_2122,In_122);
nand U729 (N_729,In_473,In_2474);
xor U730 (N_730,In_102,In_1642);
nand U731 (N_731,In_1103,In_483);
nand U732 (N_732,In_1534,In_840);
nor U733 (N_733,In_419,In_1909);
nand U734 (N_734,In_253,In_2354);
xnor U735 (N_735,In_796,In_1354);
or U736 (N_736,In_1891,In_847);
and U737 (N_737,In_2029,In_134);
or U738 (N_738,In_681,In_1243);
nor U739 (N_739,In_1061,In_176);
and U740 (N_740,In_228,In_1365);
xnor U741 (N_741,In_1351,In_1283);
or U742 (N_742,In_902,In_213);
xor U743 (N_743,In_38,In_1936);
or U744 (N_744,In_2138,In_2074);
nand U745 (N_745,In_2199,In_1565);
and U746 (N_746,In_1468,In_1772);
nor U747 (N_747,In_1646,In_544);
nand U748 (N_748,In_339,In_1381);
or U749 (N_749,In_1046,In_724);
and U750 (N_750,In_1593,In_1196);
nor U751 (N_751,In_1673,In_1725);
or U752 (N_752,In_369,In_1054);
or U753 (N_753,In_1501,In_1554);
or U754 (N_754,In_1119,In_2123);
or U755 (N_755,In_6,In_2126);
nor U756 (N_756,In_1507,In_1293);
nand U757 (N_757,In_456,In_36);
nor U758 (N_758,In_2317,In_2188);
or U759 (N_759,In_2293,In_1643);
nor U760 (N_760,In_2447,In_1121);
and U761 (N_761,In_537,In_1532);
xor U762 (N_762,In_1018,In_13);
nor U763 (N_763,In_1986,In_29);
and U764 (N_764,In_1700,In_1560);
or U765 (N_765,In_1098,In_535);
xor U766 (N_766,In_679,In_644);
nor U767 (N_767,In_1739,In_209);
nand U768 (N_768,In_2063,In_1064);
xnor U769 (N_769,In_375,In_669);
nand U770 (N_770,In_2285,In_2480);
or U771 (N_771,In_1929,In_1219);
nand U772 (N_772,In_114,In_2343);
and U773 (N_773,In_2299,In_1285);
xor U774 (N_774,In_875,In_137);
xor U775 (N_775,In_536,In_819);
nand U776 (N_776,In_723,In_970);
and U777 (N_777,In_1193,In_2024);
nand U778 (N_778,In_2184,In_56);
or U779 (N_779,In_2430,In_73);
xor U780 (N_780,In_962,In_2499);
nand U781 (N_781,In_2214,In_2473);
or U782 (N_782,In_2283,In_776);
or U783 (N_783,In_1751,In_1873);
and U784 (N_784,In_2318,In_523);
and U785 (N_785,In_347,In_2002);
xor U786 (N_786,In_2425,In_865);
and U787 (N_787,In_1014,In_1304);
nand U788 (N_788,In_2066,In_1048);
or U789 (N_789,In_2014,In_1957);
nand U790 (N_790,In_402,In_1826);
xnor U791 (N_791,In_725,In_2269);
and U792 (N_792,In_201,In_433);
nor U793 (N_793,In_385,In_1084);
or U794 (N_794,In_2159,In_1518);
nor U795 (N_795,In_1172,In_2119);
nand U796 (N_796,In_471,In_695);
and U797 (N_797,In_1228,In_2157);
nor U798 (N_798,In_481,In_492);
nand U799 (N_799,In_791,In_2077);
or U800 (N_800,In_2260,In_2357);
and U801 (N_801,In_242,In_2194);
nand U802 (N_802,In_2158,In_1755);
nand U803 (N_803,In_554,In_2256);
and U804 (N_804,In_34,In_1037);
and U805 (N_805,In_491,In_2312);
nor U806 (N_806,In_675,In_1367);
or U807 (N_807,In_177,In_2413);
and U808 (N_808,In_1612,In_757);
and U809 (N_809,In_1106,In_2136);
and U810 (N_810,In_1000,In_1271);
and U811 (N_811,In_1290,In_1231);
nand U812 (N_812,In_1386,In_1241);
or U813 (N_813,In_1298,In_1798);
nor U814 (N_814,In_884,In_735);
xnor U815 (N_815,In_2142,In_1773);
nor U816 (N_816,In_1249,In_168);
or U817 (N_817,In_1620,In_4);
and U818 (N_818,In_542,In_1752);
nand U819 (N_819,In_935,In_2163);
nor U820 (N_820,In_2108,In_1892);
nor U821 (N_821,In_1628,In_1967);
and U822 (N_822,In_2220,In_1988);
or U823 (N_823,In_270,In_1524);
or U824 (N_824,In_1706,In_908);
or U825 (N_825,In_1147,In_162);
nor U826 (N_826,In_1684,In_2418);
nor U827 (N_827,In_306,In_988);
and U828 (N_828,In_166,In_1581);
and U829 (N_829,In_172,In_1128);
xnor U830 (N_830,In_670,In_103);
or U831 (N_831,In_2453,In_1337);
or U832 (N_832,In_99,In_2064);
and U833 (N_833,In_85,In_2179);
xor U834 (N_834,In_1670,In_2451);
xnor U835 (N_835,In_592,In_637);
nor U836 (N_836,In_906,In_1840);
nor U837 (N_837,In_1994,In_2056);
nand U838 (N_838,In_1954,In_2437);
nor U839 (N_839,In_917,In_2374);
nor U840 (N_840,In_1250,In_1519);
xor U841 (N_841,In_619,In_1932);
nor U842 (N_842,In_1349,In_1715);
nand U843 (N_843,In_1467,In_94);
xnor U844 (N_844,In_2390,In_2120);
xor U845 (N_845,In_1640,In_2129);
or U846 (N_846,In_1744,In_2311);
or U847 (N_847,In_1115,In_1675);
xor U848 (N_848,In_2280,In_714);
nand U849 (N_849,In_1197,In_1662);
nand U850 (N_850,In_1060,In_1479);
xnor U851 (N_851,In_2326,In_938);
or U852 (N_852,In_315,In_560);
nand U853 (N_853,In_1124,In_983);
xnor U854 (N_854,In_2051,In_1083);
xnor U855 (N_855,In_856,In_2182);
nand U856 (N_856,In_1348,In_2468);
nand U857 (N_857,In_379,In_959);
xnor U858 (N_858,In_946,In_2132);
nor U859 (N_859,In_750,In_40);
xnor U860 (N_860,In_2409,In_244);
or U861 (N_861,In_1977,In_741);
nor U862 (N_862,In_371,In_1787);
and U863 (N_863,In_1162,In_1664);
nand U864 (N_864,In_387,In_1793);
xor U865 (N_865,In_792,In_1792);
nor U866 (N_866,In_1215,In_699);
nor U867 (N_867,In_1769,In_326);
and U868 (N_868,In_328,In_1855);
or U869 (N_869,In_1556,In_2110);
xnor U870 (N_870,In_747,In_1161);
nor U871 (N_871,In_733,In_450);
xor U872 (N_872,In_925,In_2487);
nor U873 (N_873,In_944,In_1370);
and U874 (N_874,In_153,In_2389);
xnor U875 (N_875,In_1750,In_149);
xnor U876 (N_876,In_680,In_965);
nand U877 (N_877,In_397,In_1173);
nor U878 (N_878,In_1490,In_502);
and U879 (N_879,In_1652,In_263);
nand U880 (N_880,In_2308,In_1698);
nand U881 (N_881,In_2089,In_1898);
xnor U882 (N_882,In_1603,In_897);
or U883 (N_883,In_1216,In_823);
xor U884 (N_884,In_2012,In_1733);
or U885 (N_885,In_1926,In_990);
and U886 (N_886,In_802,In_996);
nand U887 (N_887,In_1295,In_740);
nand U888 (N_888,In_787,In_1066);
nor U889 (N_889,In_1537,In_316);
nand U890 (N_890,In_607,In_1371);
nor U891 (N_891,In_143,In_2147);
and U892 (N_892,In_1975,In_1314);
nor U893 (N_893,In_940,In_188);
or U894 (N_894,In_981,In_292);
or U895 (N_895,In_185,In_1785);
or U896 (N_896,In_2028,In_587);
xor U897 (N_897,In_284,In_207);
nand U898 (N_898,In_1770,In_1481);
nor U899 (N_899,In_803,In_2211);
and U900 (N_900,In_1320,In_1492);
or U901 (N_901,In_308,In_1212);
nor U902 (N_902,In_511,In_2022);
or U903 (N_903,In_692,In_2232);
nand U904 (N_904,In_2149,In_2097);
nor U905 (N_905,In_84,In_389);
nand U906 (N_906,In_994,In_2325);
or U907 (N_907,In_507,In_979);
xor U908 (N_908,In_2115,In_325);
nor U909 (N_909,In_2098,In_1494);
and U910 (N_910,In_1953,In_307);
nor U911 (N_911,In_2047,In_1109);
xnor U912 (N_912,In_2033,In_2264);
nand U913 (N_913,In_80,In_1747);
xor U914 (N_914,In_1439,In_233);
xor U915 (N_915,In_1962,In_130);
nand U916 (N_916,In_1142,In_2015);
nand U917 (N_917,In_1692,In_1999);
or U918 (N_918,In_898,In_547);
or U919 (N_919,In_1094,In_44);
nand U920 (N_920,In_2388,In_117);
or U921 (N_921,In_805,In_1073);
xor U922 (N_922,In_1395,In_678);
nand U923 (N_923,In_163,In_595);
nand U924 (N_924,In_508,In_2161);
nor U925 (N_925,In_459,In_250);
or U926 (N_926,In_934,In_169);
xor U927 (N_927,In_815,In_1096);
or U928 (N_928,In_1516,In_32);
or U929 (N_929,In_133,In_2361);
nor U930 (N_930,In_2282,In_1653);
or U931 (N_931,In_2006,In_2476);
and U932 (N_932,In_2177,In_2286);
nand U933 (N_933,In_183,In_275);
nor U934 (N_934,In_509,In_2001);
nor U935 (N_935,In_57,In_1206);
xnor U936 (N_936,In_79,In_588);
nand U937 (N_937,In_939,In_1233);
nand U938 (N_938,In_1444,In_227);
and U939 (N_939,In_993,In_191);
or U940 (N_940,In_1026,In_2075);
or U941 (N_941,In_2382,In_1200);
and U942 (N_942,In_821,In_1425);
and U943 (N_943,In_124,In_1100);
and U944 (N_944,In_1289,In_924);
and U945 (N_945,In_1697,In_928);
and U946 (N_946,In_1028,In_1449);
xnor U947 (N_947,In_1036,In_1070);
or U948 (N_948,In_95,In_1062);
xnor U949 (N_949,In_864,In_2255);
and U950 (N_950,In_2375,In_1280);
or U951 (N_951,In_687,In_807);
and U952 (N_952,In_876,In_332);
nand U953 (N_953,In_1861,In_2086);
nor U954 (N_954,In_350,In_673);
and U955 (N_955,In_663,In_1438);
nor U956 (N_956,In_2492,In_1985);
or U957 (N_957,In_1378,In_354);
nand U958 (N_958,In_1823,In_1391);
nand U959 (N_959,In_1410,In_1987);
xnor U960 (N_960,In_1144,In_1434);
xnor U961 (N_961,In_1998,In_915);
nor U962 (N_962,In_1525,In_129);
nand U963 (N_963,In_1159,In_184);
xnor U964 (N_964,In_813,In_2102);
nand U965 (N_965,In_1633,In_89);
xor U966 (N_966,In_2085,In_1522);
nand U967 (N_967,In_2261,In_466);
nor U968 (N_968,In_854,In_1514);
xnor U969 (N_969,In_2113,In_256);
nor U970 (N_970,In_294,In_1866);
nor U971 (N_971,In_2287,In_262);
xor U972 (N_972,In_2213,In_1956);
nor U973 (N_973,In_754,In_226);
nand U974 (N_974,In_196,In_1916);
xor U975 (N_975,In_1648,In_1340);
or U976 (N_976,In_1835,In_1457);
nand U977 (N_977,In_2333,In_1355);
or U978 (N_978,In_1279,In_799);
nand U979 (N_979,In_573,In_551);
and U980 (N_980,In_240,In_2059);
nor U981 (N_981,In_1260,In_1992);
or U982 (N_982,In_1055,In_1273);
nor U983 (N_983,In_926,In_1448);
nand U984 (N_984,In_751,In_1220);
xor U985 (N_985,In_855,In_1452);
or U986 (N_986,In_1935,In_2197);
or U987 (N_987,In_2252,In_1912);
nor U988 (N_988,In_1472,In_1179);
nor U989 (N_989,In_721,In_1150);
or U990 (N_990,In_2397,In_731);
and U991 (N_991,In_527,In_403);
xor U992 (N_992,In_1482,In_873);
xnor U993 (N_993,In_2041,In_2332);
xor U994 (N_994,In_1251,In_31);
nand U995 (N_995,In_2154,In_443);
nor U996 (N_996,In_664,In_1155);
xor U997 (N_997,In_1950,In_1960);
xor U998 (N_998,In_844,In_633);
and U999 (N_999,In_586,In_1631);
nand U1000 (N_1000,In_574,In_1133);
xnor U1001 (N_1001,In_581,In_1995);
nand U1002 (N_1002,In_1767,In_2472);
nor U1003 (N_1003,In_1329,In_1464);
and U1004 (N_1004,In_531,In_1586);
nor U1005 (N_1005,In_1205,In_76);
or U1006 (N_1006,In_778,In_613);
xnor U1007 (N_1007,In_1498,In_654);
nor U1008 (N_1008,In_101,In_2358);
and U1009 (N_1009,In_2128,In_688);
nor U1010 (N_1010,In_1313,In_1214);
nand U1011 (N_1011,In_832,In_2298);
xnor U1012 (N_1012,In_2414,In_1);
and U1013 (N_1013,In_880,In_426);
and U1014 (N_1014,In_245,In_1969);
xnor U1015 (N_1015,In_1059,In_597);
nor U1016 (N_1016,In_1350,In_510);
nor U1017 (N_1017,In_2117,In_858);
nor U1018 (N_1018,In_1920,In_1786);
nor U1019 (N_1019,In_2081,In_1256);
nor U1020 (N_1020,In_1267,In_2296);
xor U1021 (N_1021,In_683,In_2381);
or U1022 (N_1022,In_1983,In_1409);
and U1023 (N_1023,In_503,In_1944);
nand U1024 (N_1024,In_986,In_2062);
nand U1025 (N_1025,In_1252,In_599);
or U1026 (N_1026,In_2235,In_264);
xnor U1027 (N_1027,In_662,In_2494);
xor U1028 (N_1028,In_2183,In_2324);
or U1029 (N_1029,In_951,In_148);
and U1030 (N_1030,In_565,In_1858);
or U1031 (N_1031,In_290,In_2405);
or U1032 (N_1032,In_836,In_23);
nor U1033 (N_1033,In_105,In_2017);
and U1034 (N_1034,In_1889,In_1199);
xor U1035 (N_1035,In_1305,In_2035);
or U1036 (N_1036,In_977,In_405);
nand U1037 (N_1037,In_514,In_2363);
or U1038 (N_1038,In_2216,In_1933);
nor U1039 (N_1039,In_1113,In_104);
xnor U1040 (N_1040,In_410,In_1632);
or U1041 (N_1041,In_234,In_303);
xnor U1042 (N_1042,In_2491,In_2469);
xor U1043 (N_1043,In_485,In_1301);
and U1044 (N_1044,In_1817,In_1404);
or U1045 (N_1045,In_1446,In_655);
xnor U1046 (N_1046,In_87,In_1687);
xor U1047 (N_1047,In_624,In_243);
xnor U1048 (N_1048,In_894,In_623);
or U1049 (N_1049,In_626,In_1911);
and U1050 (N_1050,In_2215,In_1557);
nand U1051 (N_1051,In_174,In_1297);
nand U1052 (N_1052,In_1306,In_2302);
xnor U1053 (N_1053,In_277,In_111);
and U1054 (N_1054,In_2076,In_752);
xnor U1055 (N_1055,In_806,In_1253);
or U1056 (N_1056,In_1966,In_2170);
xor U1057 (N_1057,In_1660,In_1923);
xnor U1058 (N_1058,In_380,In_1076);
nor U1059 (N_1059,In_2446,In_289);
nand U1060 (N_1060,In_2340,In_1245);
xnor U1061 (N_1061,In_2239,In_2384);
and U1062 (N_1062,In_2201,In_1980);
or U1063 (N_1063,In_850,In_1265);
nor U1064 (N_1064,In_526,In_2489);
and U1065 (N_1065,In_1970,In_1033);
nand U1066 (N_1066,In_729,In_1099);
nor U1067 (N_1067,In_1358,In_2448);
nor U1068 (N_1068,In_1157,In_2198);
nand U1069 (N_1069,In_1955,In_830);
nand U1070 (N_1070,In_2345,In_1827);
xnor U1071 (N_1071,In_1356,In_2049);
xor U1072 (N_1072,In_1105,In_438);
nand U1073 (N_1073,In_1521,In_1453);
and U1074 (N_1074,In_1820,In_498);
or U1075 (N_1075,In_1158,In_927);
or U1076 (N_1076,In_736,In_1258);
nor U1077 (N_1077,In_615,In_2335);
xor U1078 (N_1078,In_2464,In_1674);
or U1079 (N_1079,In_1585,In_2440);
nor U1080 (N_1080,In_1303,In_1497);
nor U1081 (N_1081,In_584,In_709);
or U1082 (N_1082,In_1818,In_893);
nand U1083 (N_1083,In_1591,In_550);
xnor U1084 (N_1084,In_1176,In_2277);
nand U1085 (N_1085,In_45,In_1789);
nor U1086 (N_1086,In_2139,In_1009);
nand U1087 (N_1087,In_2443,In_86);
and U1088 (N_1088,In_2265,In_2263);
or U1089 (N_1089,In_2395,In_358);
xnor U1090 (N_1090,In_1958,In_642);
and U1091 (N_1091,In_2289,In_2030);
or U1092 (N_1092,In_1388,In_1882);
and U1093 (N_1093,In_1679,In_1794);
nor U1094 (N_1094,In_373,In_342);
xor U1095 (N_1095,In_331,In_1465);
nor U1096 (N_1096,In_1254,In_260);
nand U1097 (N_1097,In_3,In_496);
or U1098 (N_1098,In_42,In_2348);
xnor U1099 (N_1099,In_717,In_2042);
and U1100 (N_1100,In_2466,In_1705);
or U1101 (N_1101,In_1065,In_689);
nor U1102 (N_1102,In_1768,In_266);
nor U1103 (N_1103,In_198,In_827);
xnor U1104 (N_1104,In_2101,In_200);
nand U1105 (N_1105,In_1154,In_1837);
nor U1106 (N_1106,In_1973,In_722);
and U1107 (N_1107,In_789,In_1852);
and U1108 (N_1108,In_1291,In_2307);
nand U1109 (N_1109,In_2034,In_304);
or U1110 (N_1110,In_98,In_899);
xor U1111 (N_1111,In_999,In_1669);
nor U1112 (N_1112,In_2292,In_2369);
xnor U1113 (N_1113,In_1900,In_2245);
and U1114 (N_1114,In_1551,In_2011);
nor U1115 (N_1115,In_2061,In_1876);
nor U1116 (N_1116,In_2377,In_157);
and U1117 (N_1117,In_1261,In_1886);
nor U1118 (N_1118,In_2243,In_377);
nand U1119 (N_1119,In_1824,In_2456);
nor U1120 (N_1120,In_1924,In_1110);
xor U1121 (N_1121,In_159,In_1777);
or U1122 (N_1122,In_589,In_829);
nand U1123 (N_1123,In_1683,In_35);
and U1124 (N_1124,In_643,In_2103);
xnor U1125 (N_1125,In_2347,In_2175);
and U1126 (N_1126,In_1965,In_1544);
nand U1127 (N_1127,In_271,In_2112);
and U1128 (N_1128,In_2130,In_1379);
nand U1129 (N_1129,In_732,In_1857);
nor U1130 (N_1130,In_1090,In_694);
nand U1131 (N_1131,In_66,In_2246);
and U1132 (N_1132,In_1711,In_2016);
nor U1133 (N_1133,In_857,In_1111);
xor U1134 (N_1134,In_835,In_2422);
nand U1135 (N_1135,In_2107,In_851);
nand U1136 (N_1136,In_77,In_1588);
and U1137 (N_1137,In_2319,In_1940);
nor U1138 (N_1138,In_685,In_1104);
or U1139 (N_1139,In_327,In_353);
and U1140 (N_1140,In_110,In_352);
or U1141 (N_1141,In_2355,In_1878);
nor U1142 (N_1142,In_346,In_1529);
nand U1143 (N_1143,In_1276,In_348);
nand U1144 (N_1144,In_1732,In_1382);
nor U1145 (N_1145,In_340,In_1602);
nor U1146 (N_1146,In_1043,In_1782);
nor U1147 (N_1147,In_278,In_1146);
nand U1148 (N_1148,In_720,In_1680);
nand U1149 (N_1149,In_1312,In_702);
nor U1150 (N_1150,In_1166,In_343);
nand U1151 (N_1151,In_2415,In_691);
and U1152 (N_1152,In_1701,In_883);
nand U1153 (N_1153,In_1224,In_112);
xor U1154 (N_1154,In_493,In_1089);
nor U1155 (N_1155,In_475,In_2336);
and U1156 (N_1156,In_809,In_773);
nor U1157 (N_1157,In_2342,In_2257);
and U1158 (N_1158,In_2207,In_8);
xor U1159 (N_1159,In_1989,In_950);
or U1160 (N_1160,In_330,In_734);
nand U1161 (N_1161,In_2095,In_46);
or U1162 (N_1162,In_1959,In_594);
nor U1163 (N_1163,In_1619,In_1025);
and U1164 (N_1164,In_442,In_158);
or U1165 (N_1165,In_1729,In_480);
nor U1166 (N_1166,In_186,In_2305);
or U1167 (N_1167,In_911,In_922);
or U1168 (N_1168,In_1058,In_984);
nand U1169 (N_1169,In_313,In_1001);
xor U1170 (N_1170,In_1771,In_2141);
nor U1171 (N_1171,In_235,In_1435);
nand U1172 (N_1172,In_1051,In_1671);
xor U1173 (N_1173,In_1847,In_219);
or U1174 (N_1174,In_611,In_1788);
xnor U1175 (N_1175,In_1087,In_814);
nand U1176 (N_1176,In_1562,In_1180);
xor U1177 (N_1177,In_82,In_497);
xnor U1178 (N_1178,In_1466,In_797);
xnor U1179 (N_1179,In_381,In_336);
xnor U1180 (N_1180,In_822,In_2486);
nor U1181 (N_1181,In_320,In_1198);
xnor U1182 (N_1182,In_1343,In_1360);
or U1183 (N_1183,In_2152,In_2417);
xor U1184 (N_1184,In_515,In_1423);
or U1185 (N_1185,In_1040,In_1101);
and U1186 (N_1186,In_1896,In_1796);
or U1187 (N_1187,In_187,In_462);
nand U1188 (N_1188,In_706,In_869);
and U1189 (N_1189,In_2150,In_1762);
xnor U1190 (N_1190,In_1893,In_955);
or U1191 (N_1191,In_1851,In_1676);
xor U1192 (N_1192,In_743,In_576);
and U1193 (N_1193,In_1039,In_2060);
nor U1194 (N_1194,In_1634,In_1515);
nand U1195 (N_1195,In_601,In_2087);
and U1196 (N_1196,In_1185,In_297);
nand U1197 (N_1197,In_738,In_2376);
or U1198 (N_1198,In_2341,In_1742);
and U1199 (N_1199,In_255,In_2328);
and U1200 (N_1200,In_1091,In_518);
nor U1201 (N_1201,In_131,In_1499);
and U1202 (N_1202,In_310,In_2124);
nand U1203 (N_1203,In_1170,In_281);
nor U1204 (N_1204,In_919,In_2196);
xnor U1205 (N_1205,In_1695,In_783);
nor U1206 (N_1206,In_451,In_1910);
and U1207 (N_1207,In_1800,In_2337);
nand U1208 (N_1208,In_2191,In_1311);
or U1209 (N_1209,In_1325,In_2379);
xor U1210 (N_1210,In_261,In_302);
or U1211 (N_1211,In_2314,In_843);
nand U1212 (N_1212,In_1330,In_1903);
and U1213 (N_1213,In_2288,In_2171);
or U1214 (N_1214,In_2166,In_2461);
xnor U1215 (N_1215,In_1248,In_1526);
nand U1216 (N_1216,In_2320,In_1538);
nand U1217 (N_1217,In_1963,In_269);
nor U1218 (N_1218,In_1238,In_609);
or U1219 (N_1219,In_418,In_1913);
xnor U1220 (N_1220,In_1321,In_676);
nand U1221 (N_1221,In_2079,In_1651);
nand U1222 (N_1222,In_248,In_1202);
nor U1223 (N_1223,In_298,In_608);
or U1224 (N_1224,In_808,In_1029);
xor U1225 (N_1225,In_345,In_2398);
xor U1226 (N_1226,In_1030,In_1686);
xor U1227 (N_1227,In_2091,In_1420);
xor U1228 (N_1228,In_1577,In_1080);
nor U1229 (N_1229,In_933,In_1780);
nand U1230 (N_1230,In_1948,In_1074);
or U1231 (N_1231,In_2267,In_634);
and U1232 (N_1232,In_1156,In_55);
xnor U1233 (N_1233,In_1474,In_1828);
nand U1234 (N_1234,In_2330,In_1389);
nand U1235 (N_1235,In_182,In_1223);
nand U1236 (N_1236,In_629,In_889);
xor U1237 (N_1237,In_1949,In_529);
nand U1238 (N_1238,In_2432,In_1006);
and U1239 (N_1239,In_2068,In_2315);
nor U1240 (N_1240,In_2394,In_1934);
and U1241 (N_1241,In_2165,In_1353);
xor U1242 (N_1242,In_1268,In_682);
nand U1243 (N_1243,In_708,In_1604);
xor U1244 (N_1244,In_179,In_2406);
and U1245 (N_1245,In_1447,In_1921);
nor U1246 (N_1246,In_1487,In_458);
and U1247 (N_1247,In_2268,In_2218);
nand U1248 (N_1248,In_967,In_64);
or U1249 (N_1249,In_1606,In_838);
nand U1250 (N_1250,In_302,In_1984);
or U1251 (N_1251,In_2009,In_2000);
xor U1252 (N_1252,In_772,In_257);
or U1253 (N_1253,In_2492,In_1157);
xor U1254 (N_1254,In_1781,In_2260);
and U1255 (N_1255,In_2045,In_1943);
or U1256 (N_1256,In_1279,In_945);
or U1257 (N_1257,In_1096,In_1028);
nor U1258 (N_1258,In_1925,In_1398);
xnor U1259 (N_1259,In_1943,In_2489);
nand U1260 (N_1260,In_70,In_1077);
nor U1261 (N_1261,In_851,In_742);
and U1262 (N_1262,In_1959,In_2491);
nor U1263 (N_1263,In_1653,In_1004);
or U1264 (N_1264,In_831,In_2174);
xnor U1265 (N_1265,In_1217,In_318);
or U1266 (N_1266,In_1122,In_71);
and U1267 (N_1267,In_1741,In_1244);
or U1268 (N_1268,In_1516,In_883);
nand U1269 (N_1269,In_329,In_449);
xnor U1270 (N_1270,In_376,In_139);
or U1271 (N_1271,In_520,In_2132);
or U1272 (N_1272,In_1361,In_1677);
and U1273 (N_1273,In_116,In_413);
xor U1274 (N_1274,In_1102,In_2247);
and U1275 (N_1275,In_1734,In_1877);
xnor U1276 (N_1276,In_2351,In_408);
nand U1277 (N_1277,In_1351,In_547);
xnor U1278 (N_1278,In_701,In_1733);
xor U1279 (N_1279,In_2460,In_692);
or U1280 (N_1280,In_1831,In_1208);
xor U1281 (N_1281,In_989,In_680);
and U1282 (N_1282,In_51,In_2340);
or U1283 (N_1283,In_902,In_835);
xor U1284 (N_1284,In_130,In_2117);
nand U1285 (N_1285,In_1976,In_731);
nand U1286 (N_1286,In_463,In_813);
nor U1287 (N_1287,In_1266,In_1424);
nor U1288 (N_1288,In_990,In_1776);
and U1289 (N_1289,In_482,In_2391);
nand U1290 (N_1290,In_196,In_663);
nand U1291 (N_1291,In_849,In_1567);
nand U1292 (N_1292,In_394,In_400);
nor U1293 (N_1293,In_837,In_1909);
nand U1294 (N_1294,In_414,In_1193);
xnor U1295 (N_1295,In_1740,In_2291);
nor U1296 (N_1296,In_2260,In_1795);
nand U1297 (N_1297,In_1199,In_2073);
nor U1298 (N_1298,In_1485,In_784);
xnor U1299 (N_1299,In_2266,In_1975);
nor U1300 (N_1300,In_1811,In_293);
and U1301 (N_1301,In_1676,In_1719);
or U1302 (N_1302,In_16,In_74);
or U1303 (N_1303,In_2095,In_54);
or U1304 (N_1304,In_939,In_109);
or U1305 (N_1305,In_319,In_1539);
nor U1306 (N_1306,In_1973,In_703);
nor U1307 (N_1307,In_439,In_1430);
and U1308 (N_1308,In_1018,In_1283);
or U1309 (N_1309,In_1453,In_1405);
nand U1310 (N_1310,In_2187,In_2059);
xor U1311 (N_1311,In_1087,In_1777);
and U1312 (N_1312,In_1187,In_831);
xor U1313 (N_1313,In_1805,In_621);
nor U1314 (N_1314,In_509,In_510);
and U1315 (N_1315,In_307,In_1523);
xnor U1316 (N_1316,In_1609,In_2427);
or U1317 (N_1317,In_1828,In_375);
and U1318 (N_1318,In_868,In_382);
nor U1319 (N_1319,In_1721,In_326);
nor U1320 (N_1320,In_1916,In_971);
and U1321 (N_1321,In_2193,In_855);
xor U1322 (N_1322,In_1125,In_728);
and U1323 (N_1323,In_2061,In_313);
nand U1324 (N_1324,In_582,In_140);
nor U1325 (N_1325,In_755,In_1215);
nor U1326 (N_1326,In_551,In_404);
nor U1327 (N_1327,In_1848,In_825);
nor U1328 (N_1328,In_1162,In_1737);
and U1329 (N_1329,In_1761,In_2223);
and U1330 (N_1330,In_1205,In_1974);
or U1331 (N_1331,In_976,In_38);
and U1332 (N_1332,In_1773,In_1506);
or U1333 (N_1333,In_2167,In_1482);
and U1334 (N_1334,In_127,In_1573);
xor U1335 (N_1335,In_783,In_353);
and U1336 (N_1336,In_1411,In_32);
and U1337 (N_1337,In_1699,In_654);
and U1338 (N_1338,In_1551,In_1360);
nor U1339 (N_1339,In_414,In_2345);
or U1340 (N_1340,In_1390,In_1286);
and U1341 (N_1341,In_2034,In_436);
nand U1342 (N_1342,In_784,In_789);
or U1343 (N_1343,In_1342,In_1006);
xor U1344 (N_1344,In_480,In_58);
or U1345 (N_1345,In_2187,In_1535);
and U1346 (N_1346,In_2422,In_1387);
and U1347 (N_1347,In_226,In_1327);
or U1348 (N_1348,In_677,In_999);
and U1349 (N_1349,In_1670,In_451);
or U1350 (N_1350,In_70,In_356);
or U1351 (N_1351,In_950,In_1596);
xor U1352 (N_1352,In_241,In_2373);
and U1353 (N_1353,In_2244,In_1398);
xor U1354 (N_1354,In_1977,In_511);
and U1355 (N_1355,In_1149,In_1171);
nor U1356 (N_1356,In_2005,In_353);
nor U1357 (N_1357,In_1854,In_1154);
and U1358 (N_1358,In_1429,In_820);
nand U1359 (N_1359,In_168,In_1762);
xnor U1360 (N_1360,In_422,In_2230);
xor U1361 (N_1361,In_1375,In_1191);
xor U1362 (N_1362,In_167,In_1524);
nand U1363 (N_1363,In_32,In_2196);
or U1364 (N_1364,In_1930,In_1773);
and U1365 (N_1365,In_1391,In_2017);
nor U1366 (N_1366,In_55,In_2208);
nor U1367 (N_1367,In_2071,In_899);
and U1368 (N_1368,In_1260,In_162);
nand U1369 (N_1369,In_1486,In_587);
nand U1370 (N_1370,In_2172,In_2270);
or U1371 (N_1371,In_1307,In_1257);
or U1372 (N_1372,In_1785,In_2362);
and U1373 (N_1373,In_1129,In_444);
and U1374 (N_1374,In_599,In_2226);
and U1375 (N_1375,In_702,In_2320);
or U1376 (N_1376,In_355,In_2046);
xor U1377 (N_1377,In_421,In_1314);
or U1378 (N_1378,In_906,In_2455);
and U1379 (N_1379,In_771,In_2392);
nor U1380 (N_1380,In_1456,In_545);
or U1381 (N_1381,In_571,In_1800);
nand U1382 (N_1382,In_1721,In_775);
or U1383 (N_1383,In_425,In_485);
and U1384 (N_1384,In_262,In_2232);
or U1385 (N_1385,In_2205,In_198);
nor U1386 (N_1386,In_1005,In_37);
or U1387 (N_1387,In_54,In_342);
or U1388 (N_1388,In_1118,In_83);
nand U1389 (N_1389,In_2486,In_1359);
xnor U1390 (N_1390,In_1493,In_2414);
and U1391 (N_1391,In_2167,In_2061);
and U1392 (N_1392,In_2047,In_900);
xnor U1393 (N_1393,In_1003,In_654);
nand U1394 (N_1394,In_731,In_227);
nor U1395 (N_1395,In_940,In_1853);
or U1396 (N_1396,In_2124,In_1225);
nand U1397 (N_1397,In_764,In_354);
nand U1398 (N_1398,In_1326,In_181);
nor U1399 (N_1399,In_924,In_217);
or U1400 (N_1400,In_1571,In_1914);
or U1401 (N_1401,In_701,In_1686);
or U1402 (N_1402,In_1738,In_848);
xor U1403 (N_1403,In_1588,In_1324);
and U1404 (N_1404,In_2361,In_933);
or U1405 (N_1405,In_1480,In_690);
xor U1406 (N_1406,In_2063,In_1229);
or U1407 (N_1407,In_1540,In_1121);
nand U1408 (N_1408,In_1683,In_1493);
and U1409 (N_1409,In_1335,In_255);
nor U1410 (N_1410,In_695,In_325);
or U1411 (N_1411,In_67,In_266);
nand U1412 (N_1412,In_342,In_1621);
or U1413 (N_1413,In_712,In_650);
and U1414 (N_1414,In_2110,In_636);
nand U1415 (N_1415,In_2385,In_777);
and U1416 (N_1416,In_2157,In_1984);
xor U1417 (N_1417,In_2334,In_1204);
xnor U1418 (N_1418,In_1884,In_2191);
and U1419 (N_1419,In_379,In_243);
nor U1420 (N_1420,In_2376,In_2381);
xnor U1421 (N_1421,In_71,In_1178);
nor U1422 (N_1422,In_1330,In_1782);
nor U1423 (N_1423,In_198,In_1152);
nor U1424 (N_1424,In_596,In_2212);
nor U1425 (N_1425,In_133,In_2188);
xnor U1426 (N_1426,In_1416,In_953);
or U1427 (N_1427,In_1476,In_2174);
or U1428 (N_1428,In_342,In_1958);
xnor U1429 (N_1429,In_2212,In_405);
nor U1430 (N_1430,In_46,In_959);
and U1431 (N_1431,In_2094,In_1254);
nor U1432 (N_1432,In_333,In_870);
xor U1433 (N_1433,In_2428,In_1073);
and U1434 (N_1434,In_2318,In_1502);
xor U1435 (N_1435,In_58,In_1187);
or U1436 (N_1436,In_362,In_63);
xor U1437 (N_1437,In_490,In_1083);
and U1438 (N_1438,In_141,In_1833);
or U1439 (N_1439,In_696,In_1750);
nor U1440 (N_1440,In_1124,In_2004);
or U1441 (N_1441,In_535,In_820);
nor U1442 (N_1442,In_483,In_948);
nor U1443 (N_1443,In_1887,In_2096);
xor U1444 (N_1444,In_2414,In_1115);
nor U1445 (N_1445,In_1808,In_1502);
or U1446 (N_1446,In_128,In_571);
and U1447 (N_1447,In_580,In_2277);
or U1448 (N_1448,In_2365,In_1521);
and U1449 (N_1449,In_216,In_2475);
nor U1450 (N_1450,In_1168,In_557);
nand U1451 (N_1451,In_1626,In_1101);
or U1452 (N_1452,In_2465,In_1020);
or U1453 (N_1453,In_465,In_396);
or U1454 (N_1454,In_1291,In_1030);
nand U1455 (N_1455,In_1399,In_1517);
nor U1456 (N_1456,In_1061,In_1916);
nor U1457 (N_1457,In_1609,In_1598);
nand U1458 (N_1458,In_101,In_19);
nand U1459 (N_1459,In_2124,In_2472);
and U1460 (N_1460,In_1773,In_26);
and U1461 (N_1461,In_2489,In_1208);
and U1462 (N_1462,In_1197,In_1736);
or U1463 (N_1463,In_1396,In_843);
nand U1464 (N_1464,In_1371,In_407);
nor U1465 (N_1465,In_1230,In_2165);
and U1466 (N_1466,In_243,In_629);
nand U1467 (N_1467,In_2030,In_1900);
xnor U1468 (N_1468,In_1750,In_844);
or U1469 (N_1469,In_1223,In_868);
and U1470 (N_1470,In_223,In_315);
or U1471 (N_1471,In_40,In_373);
or U1472 (N_1472,In_370,In_1321);
or U1473 (N_1473,In_1184,In_1013);
or U1474 (N_1474,In_1366,In_2375);
and U1475 (N_1475,In_1170,In_765);
or U1476 (N_1476,In_2150,In_455);
and U1477 (N_1477,In_1757,In_1030);
xnor U1478 (N_1478,In_187,In_1369);
nand U1479 (N_1479,In_2131,In_1913);
and U1480 (N_1480,In_768,In_2257);
and U1481 (N_1481,In_1074,In_1523);
nor U1482 (N_1482,In_904,In_590);
xor U1483 (N_1483,In_2225,In_427);
or U1484 (N_1484,In_565,In_1928);
xnor U1485 (N_1485,In_674,In_10);
nand U1486 (N_1486,In_1413,In_1799);
xor U1487 (N_1487,In_1901,In_833);
and U1488 (N_1488,In_1935,In_957);
nor U1489 (N_1489,In_292,In_488);
or U1490 (N_1490,In_1440,In_786);
and U1491 (N_1491,In_283,In_2076);
and U1492 (N_1492,In_2294,In_1859);
or U1493 (N_1493,In_1339,In_1508);
or U1494 (N_1494,In_478,In_770);
nor U1495 (N_1495,In_438,In_77);
nand U1496 (N_1496,In_688,In_1738);
nand U1497 (N_1497,In_529,In_1955);
and U1498 (N_1498,In_1193,In_652);
xor U1499 (N_1499,In_1753,In_1438);
xor U1500 (N_1500,In_970,In_234);
or U1501 (N_1501,In_2302,In_265);
or U1502 (N_1502,In_2172,In_123);
xor U1503 (N_1503,In_832,In_1503);
or U1504 (N_1504,In_522,In_778);
nor U1505 (N_1505,In_905,In_331);
or U1506 (N_1506,In_1381,In_2381);
and U1507 (N_1507,In_1444,In_177);
or U1508 (N_1508,In_854,In_2219);
or U1509 (N_1509,In_1114,In_1942);
nor U1510 (N_1510,In_971,In_2056);
xor U1511 (N_1511,In_1885,In_1401);
nor U1512 (N_1512,In_2321,In_2101);
nand U1513 (N_1513,In_1970,In_1941);
nor U1514 (N_1514,In_538,In_1904);
or U1515 (N_1515,In_1457,In_2242);
or U1516 (N_1516,In_2190,In_976);
nand U1517 (N_1517,In_2306,In_1102);
and U1518 (N_1518,In_1612,In_1236);
or U1519 (N_1519,In_1771,In_107);
nor U1520 (N_1520,In_295,In_285);
and U1521 (N_1521,In_31,In_311);
xor U1522 (N_1522,In_2262,In_1244);
xnor U1523 (N_1523,In_1017,In_750);
and U1524 (N_1524,In_1798,In_943);
and U1525 (N_1525,In_2257,In_581);
nand U1526 (N_1526,In_637,In_331);
or U1527 (N_1527,In_1644,In_1918);
nand U1528 (N_1528,In_1791,In_2225);
and U1529 (N_1529,In_1437,In_1007);
and U1530 (N_1530,In_646,In_2327);
nor U1531 (N_1531,In_1052,In_1865);
nand U1532 (N_1532,In_1979,In_2090);
xnor U1533 (N_1533,In_1893,In_59);
or U1534 (N_1534,In_2294,In_2307);
nand U1535 (N_1535,In_479,In_947);
and U1536 (N_1536,In_918,In_1507);
or U1537 (N_1537,In_2146,In_1729);
and U1538 (N_1538,In_220,In_163);
xor U1539 (N_1539,In_1370,In_1246);
nor U1540 (N_1540,In_2417,In_1191);
or U1541 (N_1541,In_630,In_2226);
or U1542 (N_1542,In_2082,In_280);
or U1543 (N_1543,In_625,In_1384);
nand U1544 (N_1544,In_1551,In_119);
nand U1545 (N_1545,In_144,In_1206);
xnor U1546 (N_1546,In_2086,In_986);
nor U1547 (N_1547,In_1800,In_2006);
xnor U1548 (N_1548,In_2168,In_1181);
nor U1549 (N_1549,In_1318,In_1259);
nor U1550 (N_1550,In_368,In_396);
xnor U1551 (N_1551,In_877,In_1780);
and U1552 (N_1552,In_1796,In_1515);
xnor U1553 (N_1553,In_2098,In_1759);
or U1554 (N_1554,In_960,In_2333);
xnor U1555 (N_1555,In_2226,In_259);
xnor U1556 (N_1556,In_2034,In_2031);
or U1557 (N_1557,In_908,In_909);
nand U1558 (N_1558,In_1662,In_681);
xor U1559 (N_1559,In_626,In_1176);
nor U1560 (N_1560,In_338,In_216);
nor U1561 (N_1561,In_527,In_901);
nand U1562 (N_1562,In_1492,In_878);
nand U1563 (N_1563,In_1725,In_1541);
nand U1564 (N_1564,In_1466,In_328);
and U1565 (N_1565,In_235,In_1568);
or U1566 (N_1566,In_304,In_1154);
nor U1567 (N_1567,In_1470,In_1181);
or U1568 (N_1568,In_2352,In_2412);
nor U1569 (N_1569,In_1516,In_1072);
nand U1570 (N_1570,In_1808,In_1921);
nand U1571 (N_1571,In_157,In_1098);
nand U1572 (N_1572,In_410,In_1320);
and U1573 (N_1573,In_1425,In_1011);
and U1574 (N_1574,In_1089,In_355);
and U1575 (N_1575,In_2126,In_1404);
xor U1576 (N_1576,In_1134,In_1622);
nor U1577 (N_1577,In_546,In_339);
and U1578 (N_1578,In_809,In_132);
or U1579 (N_1579,In_958,In_436);
or U1580 (N_1580,In_663,In_359);
nand U1581 (N_1581,In_125,In_2151);
xor U1582 (N_1582,In_1363,In_1530);
nand U1583 (N_1583,In_1677,In_2035);
nand U1584 (N_1584,In_922,In_1005);
nand U1585 (N_1585,In_1819,In_1288);
and U1586 (N_1586,In_1561,In_1159);
nand U1587 (N_1587,In_703,In_915);
xor U1588 (N_1588,In_635,In_1012);
or U1589 (N_1589,In_23,In_1949);
xnor U1590 (N_1590,In_804,In_1968);
nand U1591 (N_1591,In_2010,In_1108);
and U1592 (N_1592,In_1129,In_1560);
and U1593 (N_1593,In_213,In_2061);
or U1594 (N_1594,In_213,In_2337);
or U1595 (N_1595,In_1551,In_549);
xnor U1596 (N_1596,In_1821,In_215);
xnor U1597 (N_1597,In_2108,In_1539);
and U1598 (N_1598,In_1162,In_2310);
or U1599 (N_1599,In_842,In_699);
and U1600 (N_1600,In_1292,In_2103);
xnor U1601 (N_1601,In_900,In_2119);
nand U1602 (N_1602,In_1730,In_2483);
nand U1603 (N_1603,In_493,In_1184);
nor U1604 (N_1604,In_1903,In_1438);
nor U1605 (N_1605,In_1989,In_818);
and U1606 (N_1606,In_264,In_1452);
and U1607 (N_1607,In_1371,In_479);
or U1608 (N_1608,In_755,In_245);
and U1609 (N_1609,In_1188,In_621);
nand U1610 (N_1610,In_668,In_1544);
or U1611 (N_1611,In_1719,In_1867);
or U1612 (N_1612,In_667,In_884);
nand U1613 (N_1613,In_2238,In_1947);
nor U1614 (N_1614,In_2461,In_62);
nor U1615 (N_1615,In_1135,In_704);
nand U1616 (N_1616,In_1372,In_2175);
nand U1617 (N_1617,In_1779,In_2410);
xor U1618 (N_1618,In_1833,In_1696);
and U1619 (N_1619,In_208,In_955);
xor U1620 (N_1620,In_798,In_2211);
or U1621 (N_1621,In_1337,In_1173);
or U1622 (N_1622,In_2323,In_333);
and U1623 (N_1623,In_395,In_674);
and U1624 (N_1624,In_762,In_552);
nor U1625 (N_1625,In_207,In_185);
nor U1626 (N_1626,In_1045,In_103);
or U1627 (N_1627,In_2441,In_1352);
nor U1628 (N_1628,In_2372,In_1290);
or U1629 (N_1629,In_1360,In_966);
and U1630 (N_1630,In_443,In_350);
xnor U1631 (N_1631,In_1401,In_2399);
or U1632 (N_1632,In_260,In_1032);
and U1633 (N_1633,In_888,In_889);
or U1634 (N_1634,In_1524,In_1190);
xor U1635 (N_1635,In_1849,In_1025);
nor U1636 (N_1636,In_2255,In_900);
xnor U1637 (N_1637,In_1619,In_1886);
nand U1638 (N_1638,In_2257,In_1047);
nor U1639 (N_1639,In_1977,In_1410);
nand U1640 (N_1640,In_969,In_1812);
or U1641 (N_1641,In_44,In_1469);
and U1642 (N_1642,In_2470,In_1322);
or U1643 (N_1643,In_687,In_1301);
nor U1644 (N_1644,In_794,In_929);
nor U1645 (N_1645,In_497,In_238);
and U1646 (N_1646,In_783,In_2358);
xnor U1647 (N_1647,In_517,In_1547);
and U1648 (N_1648,In_536,In_488);
nand U1649 (N_1649,In_2217,In_1025);
nand U1650 (N_1650,In_1409,In_1283);
xor U1651 (N_1651,In_2400,In_196);
nand U1652 (N_1652,In_1992,In_1245);
nand U1653 (N_1653,In_983,In_1037);
or U1654 (N_1654,In_816,In_860);
nand U1655 (N_1655,In_1054,In_2121);
nand U1656 (N_1656,In_19,In_1029);
and U1657 (N_1657,In_2399,In_944);
xnor U1658 (N_1658,In_515,In_700);
or U1659 (N_1659,In_1873,In_718);
or U1660 (N_1660,In_763,In_2049);
xnor U1661 (N_1661,In_2351,In_1805);
or U1662 (N_1662,In_1628,In_1434);
and U1663 (N_1663,In_1671,In_1622);
nor U1664 (N_1664,In_214,In_506);
nor U1665 (N_1665,In_2382,In_873);
or U1666 (N_1666,In_494,In_1663);
or U1667 (N_1667,In_2401,In_677);
nor U1668 (N_1668,In_2427,In_274);
nor U1669 (N_1669,In_323,In_696);
or U1670 (N_1670,In_177,In_1486);
or U1671 (N_1671,In_2065,In_805);
xnor U1672 (N_1672,In_1269,In_1994);
xor U1673 (N_1673,In_348,In_426);
and U1674 (N_1674,In_157,In_608);
or U1675 (N_1675,In_2435,In_1530);
or U1676 (N_1676,In_1349,In_1643);
and U1677 (N_1677,In_815,In_148);
and U1678 (N_1678,In_58,In_145);
or U1679 (N_1679,In_653,In_367);
or U1680 (N_1680,In_64,In_2379);
nand U1681 (N_1681,In_1470,In_539);
or U1682 (N_1682,In_1404,In_1626);
nor U1683 (N_1683,In_1108,In_519);
nor U1684 (N_1684,In_1317,In_1307);
nor U1685 (N_1685,In_2441,In_1931);
xnor U1686 (N_1686,In_1339,In_56);
and U1687 (N_1687,In_815,In_1890);
nor U1688 (N_1688,In_378,In_979);
nand U1689 (N_1689,In_3,In_1968);
nand U1690 (N_1690,In_2338,In_996);
and U1691 (N_1691,In_397,In_2323);
or U1692 (N_1692,In_3,In_1373);
nand U1693 (N_1693,In_2068,In_569);
xor U1694 (N_1694,In_447,In_652);
xnor U1695 (N_1695,In_1061,In_1142);
nand U1696 (N_1696,In_55,In_1878);
nand U1697 (N_1697,In_1227,In_1735);
or U1698 (N_1698,In_318,In_1654);
xor U1699 (N_1699,In_358,In_1565);
and U1700 (N_1700,In_218,In_988);
or U1701 (N_1701,In_953,In_1775);
nor U1702 (N_1702,In_555,In_377);
and U1703 (N_1703,In_606,In_1784);
or U1704 (N_1704,In_539,In_583);
xor U1705 (N_1705,In_2107,In_52);
or U1706 (N_1706,In_608,In_481);
and U1707 (N_1707,In_1531,In_2215);
and U1708 (N_1708,In_919,In_2139);
nand U1709 (N_1709,In_2377,In_1578);
and U1710 (N_1710,In_1577,In_1275);
nor U1711 (N_1711,In_1578,In_611);
nand U1712 (N_1712,In_114,In_1333);
nand U1713 (N_1713,In_636,In_1221);
and U1714 (N_1714,In_1593,In_1368);
and U1715 (N_1715,In_1536,In_2188);
xor U1716 (N_1716,In_2068,In_456);
or U1717 (N_1717,In_2420,In_549);
nor U1718 (N_1718,In_886,In_10);
nand U1719 (N_1719,In_1922,In_316);
and U1720 (N_1720,In_260,In_381);
and U1721 (N_1721,In_1396,In_987);
nor U1722 (N_1722,In_1366,In_1139);
or U1723 (N_1723,In_593,In_1051);
or U1724 (N_1724,In_325,In_2418);
xnor U1725 (N_1725,In_991,In_395);
nor U1726 (N_1726,In_928,In_1282);
nand U1727 (N_1727,In_1410,In_590);
xnor U1728 (N_1728,In_1108,In_2280);
xnor U1729 (N_1729,In_1374,In_496);
and U1730 (N_1730,In_193,In_1817);
nor U1731 (N_1731,In_843,In_1050);
and U1732 (N_1732,In_2133,In_2066);
or U1733 (N_1733,In_857,In_716);
nor U1734 (N_1734,In_1133,In_1401);
xnor U1735 (N_1735,In_1434,In_537);
or U1736 (N_1736,In_60,In_147);
xnor U1737 (N_1737,In_1424,In_302);
and U1738 (N_1738,In_1814,In_2245);
nor U1739 (N_1739,In_1953,In_2263);
xnor U1740 (N_1740,In_1004,In_1576);
and U1741 (N_1741,In_2497,In_592);
nand U1742 (N_1742,In_1591,In_2149);
and U1743 (N_1743,In_2193,In_333);
or U1744 (N_1744,In_267,In_488);
nand U1745 (N_1745,In_505,In_621);
nand U1746 (N_1746,In_824,In_1046);
nand U1747 (N_1747,In_895,In_1005);
nand U1748 (N_1748,In_1257,In_867);
xor U1749 (N_1749,In_1829,In_1438);
nand U1750 (N_1750,In_729,In_1635);
or U1751 (N_1751,In_1433,In_947);
xor U1752 (N_1752,In_2308,In_780);
nand U1753 (N_1753,In_1761,In_776);
or U1754 (N_1754,In_1530,In_475);
nor U1755 (N_1755,In_979,In_1636);
xnor U1756 (N_1756,In_133,In_555);
or U1757 (N_1757,In_2192,In_1476);
xor U1758 (N_1758,In_770,In_1293);
nand U1759 (N_1759,In_719,In_1619);
or U1760 (N_1760,In_2082,In_1817);
nand U1761 (N_1761,In_1443,In_653);
nand U1762 (N_1762,In_335,In_2141);
and U1763 (N_1763,In_1145,In_161);
nor U1764 (N_1764,In_1327,In_2134);
and U1765 (N_1765,In_2150,In_109);
nor U1766 (N_1766,In_833,In_1);
nor U1767 (N_1767,In_93,In_1528);
or U1768 (N_1768,In_1673,In_1128);
nor U1769 (N_1769,In_694,In_19);
and U1770 (N_1770,In_1456,In_1756);
nand U1771 (N_1771,In_2278,In_7);
nor U1772 (N_1772,In_323,In_377);
nand U1773 (N_1773,In_365,In_2177);
and U1774 (N_1774,In_377,In_370);
and U1775 (N_1775,In_2119,In_315);
or U1776 (N_1776,In_1528,In_705);
nand U1777 (N_1777,In_2490,In_1608);
nand U1778 (N_1778,In_1332,In_1963);
xor U1779 (N_1779,In_280,In_2136);
xor U1780 (N_1780,In_2385,In_1738);
and U1781 (N_1781,In_195,In_726);
nand U1782 (N_1782,In_2395,In_972);
nor U1783 (N_1783,In_304,In_887);
nor U1784 (N_1784,In_2073,In_2499);
xnor U1785 (N_1785,In_654,In_1231);
or U1786 (N_1786,In_582,In_1457);
nand U1787 (N_1787,In_1572,In_1575);
and U1788 (N_1788,In_1765,In_83);
xnor U1789 (N_1789,In_1978,In_1083);
nor U1790 (N_1790,In_2097,In_1060);
nor U1791 (N_1791,In_1602,In_1713);
nand U1792 (N_1792,In_1846,In_1292);
xnor U1793 (N_1793,In_709,In_433);
nor U1794 (N_1794,In_597,In_1068);
or U1795 (N_1795,In_1158,In_573);
nor U1796 (N_1796,In_99,In_819);
or U1797 (N_1797,In_1712,In_349);
nor U1798 (N_1798,In_1520,In_370);
nor U1799 (N_1799,In_577,In_376);
nand U1800 (N_1800,In_1386,In_2200);
xnor U1801 (N_1801,In_1929,In_462);
xnor U1802 (N_1802,In_896,In_1205);
nand U1803 (N_1803,In_2151,In_1839);
and U1804 (N_1804,In_1170,In_1032);
nand U1805 (N_1805,In_2046,In_878);
or U1806 (N_1806,In_2446,In_2296);
nand U1807 (N_1807,In_1210,In_2220);
or U1808 (N_1808,In_1709,In_843);
or U1809 (N_1809,In_20,In_416);
xor U1810 (N_1810,In_2171,In_1240);
nand U1811 (N_1811,In_1595,In_1548);
or U1812 (N_1812,In_924,In_277);
xnor U1813 (N_1813,In_1633,In_2494);
or U1814 (N_1814,In_1544,In_319);
and U1815 (N_1815,In_2482,In_908);
and U1816 (N_1816,In_1781,In_405);
or U1817 (N_1817,In_1028,In_1447);
xnor U1818 (N_1818,In_2105,In_1148);
xnor U1819 (N_1819,In_87,In_2060);
and U1820 (N_1820,In_469,In_1122);
xnor U1821 (N_1821,In_1815,In_1548);
xor U1822 (N_1822,In_91,In_1299);
xor U1823 (N_1823,In_2108,In_1757);
nor U1824 (N_1824,In_1003,In_610);
nand U1825 (N_1825,In_602,In_1679);
nor U1826 (N_1826,In_725,In_2355);
xor U1827 (N_1827,In_1967,In_2325);
xor U1828 (N_1828,In_1818,In_1953);
xor U1829 (N_1829,In_1348,In_2150);
and U1830 (N_1830,In_983,In_2360);
xnor U1831 (N_1831,In_1093,In_725);
and U1832 (N_1832,In_1642,In_1695);
nor U1833 (N_1833,In_1209,In_1981);
nand U1834 (N_1834,In_1297,In_1323);
xor U1835 (N_1835,In_1317,In_616);
nor U1836 (N_1836,In_2105,In_882);
nor U1837 (N_1837,In_892,In_823);
xnor U1838 (N_1838,In_513,In_423);
or U1839 (N_1839,In_619,In_2313);
and U1840 (N_1840,In_2390,In_1153);
nand U1841 (N_1841,In_2348,In_1776);
nand U1842 (N_1842,In_2055,In_1744);
nor U1843 (N_1843,In_1940,In_627);
nor U1844 (N_1844,In_1102,In_1316);
nor U1845 (N_1845,In_2455,In_896);
and U1846 (N_1846,In_1703,In_1396);
xnor U1847 (N_1847,In_664,In_413);
xnor U1848 (N_1848,In_2331,In_1280);
or U1849 (N_1849,In_985,In_1159);
xor U1850 (N_1850,In_957,In_276);
and U1851 (N_1851,In_360,In_1859);
nor U1852 (N_1852,In_2332,In_57);
or U1853 (N_1853,In_549,In_1433);
or U1854 (N_1854,In_1913,In_2177);
and U1855 (N_1855,In_1478,In_505);
xnor U1856 (N_1856,In_2315,In_1427);
nand U1857 (N_1857,In_808,In_1900);
nor U1858 (N_1858,In_2163,In_1416);
xnor U1859 (N_1859,In_693,In_700);
nor U1860 (N_1860,In_1555,In_77);
xnor U1861 (N_1861,In_1043,In_686);
xor U1862 (N_1862,In_1650,In_1284);
or U1863 (N_1863,In_1902,In_215);
nor U1864 (N_1864,In_1785,In_1314);
or U1865 (N_1865,In_2306,In_295);
or U1866 (N_1866,In_541,In_1430);
nor U1867 (N_1867,In_709,In_1672);
nand U1868 (N_1868,In_1622,In_2109);
and U1869 (N_1869,In_194,In_461);
nor U1870 (N_1870,In_1567,In_2160);
and U1871 (N_1871,In_2320,In_421);
nor U1872 (N_1872,In_574,In_1745);
xor U1873 (N_1873,In_447,In_857);
xnor U1874 (N_1874,In_1545,In_1833);
and U1875 (N_1875,In_1452,In_1235);
xor U1876 (N_1876,In_1137,In_315);
xnor U1877 (N_1877,In_850,In_891);
nand U1878 (N_1878,In_153,In_300);
xnor U1879 (N_1879,In_2400,In_1847);
xor U1880 (N_1880,In_1690,In_1092);
or U1881 (N_1881,In_740,In_247);
xor U1882 (N_1882,In_1627,In_391);
xnor U1883 (N_1883,In_1778,In_2027);
nor U1884 (N_1884,In_2059,In_283);
nor U1885 (N_1885,In_813,In_1789);
nand U1886 (N_1886,In_2198,In_2190);
xnor U1887 (N_1887,In_388,In_1712);
nand U1888 (N_1888,In_1413,In_1038);
nand U1889 (N_1889,In_2073,In_2242);
or U1890 (N_1890,In_99,In_2080);
or U1891 (N_1891,In_7,In_2251);
nor U1892 (N_1892,In_2417,In_588);
and U1893 (N_1893,In_2186,In_1472);
or U1894 (N_1894,In_2006,In_2232);
nand U1895 (N_1895,In_2433,In_2320);
and U1896 (N_1896,In_19,In_835);
or U1897 (N_1897,In_2265,In_2063);
or U1898 (N_1898,In_508,In_75);
or U1899 (N_1899,In_1158,In_1754);
or U1900 (N_1900,In_377,In_2221);
nand U1901 (N_1901,In_1819,In_2005);
nand U1902 (N_1902,In_306,In_1622);
or U1903 (N_1903,In_943,In_1910);
xor U1904 (N_1904,In_1209,In_2067);
or U1905 (N_1905,In_175,In_726);
nor U1906 (N_1906,In_2250,In_1385);
nand U1907 (N_1907,In_1490,In_2006);
or U1908 (N_1908,In_1278,In_2481);
nor U1909 (N_1909,In_1760,In_1877);
or U1910 (N_1910,In_507,In_343);
xnor U1911 (N_1911,In_1577,In_1030);
or U1912 (N_1912,In_2356,In_508);
and U1913 (N_1913,In_292,In_160);
or U1914 (N_1914,In_1406,In_425);
nand U1915 (N_1915,In_701,In_588);
or U1916 (N_1916,In_2158,In_1301);
and U1917 (N_1917,In_351,In_742);
nor U1918 (N_1918,In_940,In_325);
nor U1919 (N_1919,In_425,In_1813);
and U1920 (N_1920,In_960,In_1415);
or U1921 (N_1921,In_573,In_1436);
nor U1922 (N_1922,In_1152,In_1189);
nor U1923 (N_1923,In_131,In_332);
and U1924 (N_1924,In_2181,In_1655);
xor U1925 (N_1925,In_2409,In_130);
and U1926 (N_1926,In_720,In_593);
xor U1927 (N_1927,In_1392,In_564);
xnor U1928 (N_1928,In_2012,In_75);
or U1929 (N_1929,In_1215,In_124);
or U1930 (N_1930,In_1959,In_528);
and U1931 (N_1931,In_1553,In_1926);
nor U1932 (N_1932,In_1785,In_180);
nand U1933 (N_1933,In_605,In_2343);
or U1934 (N_1934,In_2249,In_959);
nand U1935 (N_1935,In_1133,In_142);
and U1936 (N_1936,In_1438,In_173);
xnor U1937 (N_1937,In_886,In_1964);
and U1938 (N_1938,In_1934,In_2196);
nand U1939 (N_1939,In_1324,In_1288);
nor U1940 (N_1940,In_1889,In_1654);
and U1941 (N_1941,In_1128,In_397);
and U1942 (N_1942,In_1356,In_582);
nand U1943 (N_1943,In_1709,In_2197);
or U1944 (N_1944,In_2378,In_1680);
or U1945 (N_1945,In_2366,In_2105);
or U1946 (N_1946,In_1158,In_2048);
nand U1947 (N_1947,In_89,In_2138);
or U1948 (N_1948,In_2431,In_517);
or U1949 (N_1949,In_1882,In_28);
nor U1950 (N_1950,In_405,In_1550);
xor U1951 (N_1951,In_2360,In_133);
xnor U1952 (N_1952,In_2079,In_691);
nor U1953 (N_1953,In_757,In_1706);
xnor U1954 (N_1954,In_2351,In_972);
nand U1955 (N_1955,In_461,In_2242);
and U1956 (N_1956,In_1628,In_2290);
or U1957 (N_1957,In_1920,In_2362);
xnor U1958 (N_1958,In_2251,In_1624);
nor U1959 (N_1959,In_1398,In_1239);
nor U1960 (N_1960,In_663,In_1770);
nand U1961 (N_1961,In_14,In_239);
xor U1962 (N_1962,In_1625,In_921);
xnor U1963 (N_1963,In_93,In_1193);
nor U1964 (N_1964,In_2374,In_434);
xor U1965 (N_1965,In_938,In_1235);
nor U1966 (N_1966,In_694,In_2483);
or U1967 (N_1967,In_115,In_2337);
xnor U1968 (N_1968,In_1549,In_1663);
and U1969 (N_1969,In_2107,In_454);
nand U1970 (N_1970,In_411,In_394);
nand U1971 (N_1971,In_1541,In_2295);
and U1972 (N_1972,In_122,In_2128);
xnor U1973 (N_1973,In_1513,In_731);
xor U1974 (N_1974,In_56,In_333);
xnor U1975 (N_1975,In_1571,In_1618);
or U1976 (N_1976,In_2224,In_2330);
nor U1977 (N_1977,In_1760,In_1765);
or U1978 (N_1978,In_848,In_1507);
or U1979 (N_1979,In_522,In_1045);
nor U1980 (N_1980,In_1023,In_787);
and U1981 (N_1981,In_528,In_1413);
nand U1982 (N_1982,In_289,In_1361);
xor U1983 (N_1983,In_1497,In_897);
nand U1984 (N_1984,In_1175,In_2372);
nand U1985 (N_1985,In_1037,In_1436);
nand U1986 (N_1986,In_1540,In_427);
or U1987 (N_1987,In_949,In_492);
xnor U1988 (N_1988,In_562,In_103);
nor U1989 (N_1989,In_281,In_347);
or U1990 (N_1990,In_1965,In_54);
xor U1991 (N_1991,In_1265,In_595);
and U1992 (N_1992,In_1109,In_2459);
xnor U1993 (N_1993,In_136,In_2475);
nand U1994 (N_1994,In_2389,In_317);
nand U1995 (N_1995,In_877,In_305);
nand U1996 (N_1996,In_1897,In_1378);
nor U1997 (N_1997,In_627,In_750);
and U1998 (N_1998,In_953,In_2069);
or U1999 (N_1999,In_966,In_1940);
nand U2000 (N_2000,In_2277,In_2210);
and U2001 (N_2001,In_1472,In_1048);
nand U2002 (N_2002,In_674,In_696);
or U2003 (N_2003,In_1362,In_543);
nand U2004 (N_2004,In_180,In_200);
or U2005 (N_2005,In_813,In_1961);
xor U2006 (N_2006,In_1286,In_1652);
nand U2007 (N_2007,In_1499,In_1978);
and U2008 (N_2008,In_805,In_552);
nand U2009 (N_2009,In_386,In_2481);
or U2010 (N_2010,In_1617,In_432);
xor U2011 (N_2011,In_2240,In_1641);
and U2012 (N_2012,In_1644,In_230);
nand U2013 (N_2013,In_803,In_2183);
or U2014 (N_2014,In_1183,In_497);
nand U2015 (N_2015,In_686,In_2331);
and U2016 (N_2016,In_2418,In_731);
xnor U2017 (N_2017,In_0,In_1376);
xor U2018 (N_2018,In_959,In_528);
nor U2019 (N_2019,In_843,In_408);
nand U2020 (N_2020,In_715,In_2496);
and U2021 (N_2021,In_424,In_1172);
and U2022 (N_2022,In_148,In_1204);
nor U2023 (N_2023,In_1191,In_1014);
xor U2024 (N_2024,In_418,In_2188);
nor U2025 (N_2025,In_2383,In_1455);
or U2026 (N_2026,In_237,In_1127);
nand U2027 (N_2027,In_845,In_258);
xor U2028 (N_2028,In_1827,In_2184);
and U2029 (N_2029,In_1577,In_1880);
nand U2030 (N_2030,In_937,In_1259);
and U2031 (N_2031,In_1935,In_1621);
and U2032 (N_2032,In_2221,In_430);
and U2033 (N_2033,In_2189,In_2086);
nor U2034 (N_2034,In_1069,In_661);
xnor U2035 (N_2035,In_192,In_1226);
and U2036 (N_2036,In_1873,In_963);
nor U2037 (N_2037,In_1977,In_876);
nand U2038 (N_2038,In_1315,In_542);
nand U2039 (N_2039,In_155,In_1011);
xnor U2040 (N_2040,In_2424,In_1193);
or U2041 (N_2041,In_482,In_942);
nand U2042 (N_2042,In_1646,In_1321);
nand U2043 (N_2043,In_2310,In_40);
nor U2044 (N_2044,In_131,In_482);
nor U2045 (N_2045,In_365,In_1769);
and U2046 (N_2046,In_1112,In_1520);
and U2047 (N_2047,In_1347,In_1957);
nand U2048 (N_2048,In_1589,In_64);
or U2049 (N_2049,In_626,In_1975);
or U2050 (N_2050,In_2320,In_2397);
nand U2051 (N_2051,In_772,In_1787);
and U2052 (N_2052,In_720,In_32);
and U2053 (N_2053,In_1094,In_1836);
nand U2054 (N_2054,In_393,In_2343);
and U2055 (N_2055,In_848,In_240);
nor U2056 (N_2056,In_1702,In_2351);
and U2057 (N_2057,In_2018,In_630);
nor U2058 (N_2058,In_1952,In_1530);
and U2059 (N_2059,In_1471,In_2314);
or U2060 (N_2060,In_1712,In_2128);
and U2061 (N_2061,In_1113,In_252);
nor U2062 (N_2062,In_1657,In_1459);
nor U2063 (N_2063,In_860,In_337);
nand U2064 (N_2064,In_401,In_911);
nor U2065 (N_2065,In_379,In_2326);
and U2066 (N_2066,In_1077,In_1018);
nor U2067 (N_2067,In_10,In_788);
xor U2068 (N_2068,In_1134,In_434);
nor U2069 (N_2069,In_398,In_1833);
nand U2070 (N_2070,In_1581,In_1804);
nor U2071 (N_2071,In_2443,In_1833);
or U2072 (N_2072,In_929,In_1989);
or U2073 (N_2073,In_949,In_654);
nand U2074 (N_2074,In_119,In_2135);
or U2075 (N_2075,In_1768,In_657);
and U2076 (N_2076,In_307,In_819);
nand U2077 (N_2077,In_1490,In_1937);
nor U2078 (N_2078,In_1653,In_1155);
or U2079 (N_2079,In_1046,In_1218);
or U2080 (N_2080,In_665,In_411);
nor U2081 (N_2081,In_913,In_1333);
or U2082 (N_2082,In_1767,In_1165);
xnor U2083 (N_2083,In_46,In_1608);
nand U2084 (N_2084,In_2032,In_2178);
xnor U2085 (N_2085,In_472,In_1115);
nor U2086 (N_2086,In_1583,In_579);
or U2087 (N_2087,In_2002,In_2241);
or U2088 (N_2088,In_87,In_1602);
and U2089 (N_2089,In_2170,In_1036);
or U2090 (N_2090,In_767,In_779);
xor U2091 (N_2091,In_1260,In_1318);
nor U2092 (N_2092,In_895,In_1141);
nor U2093 (N_2093,In_1971,In_685);
or U2094 (N_2094,In_301,In_1558);
nor U2095 (N_2095,In_1006,In_1044);
and U2096 (N_2096,In_1414,In_1155);
and U2097 (N_2097,In_732,In_1529);
and U2098 (N_2098,In_214,In_1878);
or U2099 (N_2099,In_2386,In_2300);
xor U2100 (N_2100,In_288,In_1658);
or U2101 (N_2101,In_638,In_703);
nand U2102 (N_2102,In_423,In_1297);
and U2103 (N_2103,In_1617,In_2321);
or U2104 (N_2104,In_2,In_1034);
xor U2105 (N_2105,In_1945,In_2293);
xor U2106 (N_2106,In_837,In_913);
nor U2107 (N_2107,In_476,In_1856);
xor U2108 (N_2108,In_1181,In_259);
xnor U2109 (N_2109,In_666,In_564);
xor U2110 (N_2110,In_2297,In_1625);
xor U2111 (N_2111,In_530,In_1281);
and U2112 (N_2112,In_106,In_2166);
xnor U2113 (N_2113,In_2345,In_474);
and U2114 (N_2114,In_389,In_1572);
and U2115 (N_2115,In_2145,In_625);
or U2116 (N_2116,In_759,In_438);
and U2117 (N_2117,In_873,In_2352);
nand U2118 (N_2118,In_2275,In_1288);
nor U2119 (N_2119,In_100,In_930);
or U2120 (N_2120,In_1285,In_1038);
or U2121 (N_2121,In_113,In_1550);
nor U2122 (N_2122,In_2243,In_641);
xnor U2123 (N_2123,In_191,In_1396);
nor U2124 (N_2124,In_24,In_2393);
and U2125 (N_2125,In_1314,In_1044);
xnor U2126 (N_2126,In_1555,In_2471);
nor U2127 (N_2127,In_1874,In_794);
or U2128 (N_2128,In_2172,In_1353);
nor U2129 (N_2129,In_2336,In_835);
nor U2130 (N_2130,In_1054,In_1392);
and U2131 (N_2131,In_590,In_1797);
nand U2132 (N_2132,In_0,In_787);
or U2133 (N_2133,In_1208,In_691);
and U2134 (N_2134,In_1448,In_1090);
nand U2135 (N_2135,In_477,In_659);
xor U2136 (N_2136,In_2379,In_786);
and U2137 (N_2137,In_696,In_336);
nor U2138 (N_2138,In_23,In_1341);
xor U2139 (N_2139,In_1382,In_2177);
xnor U2140 (N_2140,In_1687,In_1590);
and U2141 (N_2141,In_1361,In_1296);
nor U2142 (N_2142,In_1202,In_665);
or U2143 (N_2143,In_1328,In_2250);
nor U2144 (N_2144,In_742,In_2201);
nor U2145 (N_2145,In_1785,In_803);
nor U2146 (N_2146,In_280,In_2469);
and U2147 (N_2147,In_940,In_762);
xnor U2148 (N_2148,In_2083,In_1781);
nand U2149 (N_2149,In_1993,In_1465);
nand U2150 (N_2150,In_2164,In_2469);
nor U2151 (N_2151,In_187,In_258);
and U2152 (N_2152,In_1156,In_2060);
nand U2153 (N_2153,In_1658,In_380);
nand U2154 (N_2154,In_169,In_2402);
xor U2155 (N_2155,In_698,In_2067);
and U2156 (N_2156,In_529,In_2254);
xnor U2157 (N_2157,In_537,In_2289);
or U2158 (N_2158,In_475,In_1110);
or U2159 (N_2159,In_715,In_264);
nor U2160 (N_2160,In_1562,In_2425);
xor U2161 (N_2161,In_1045,In_95);
nor U2162 (N_2162,In_450,In_1845);
nor U2163 (N_2163,In_2415,In_1665);
nand U2164 (N_2164,In_2396,In_603);
xor U2165 (N_2165,In_1141,In_2035);
nor U2166 (N_2166,In_1740,In_1377);
nor U2167 (N_2167,In_517,In_972);
xnor U2168 (N_2168,In_1676,In_703);
nor U2169 (N_2169,In_745,In_2020);
or U2170 (N_2170,In_1748,In_880);
nand U2171 (N_2171,In_403,In_172);
xor U2172 (N_2172,In_872,In_531);
and U2173 (N_2173,In_862,In_2057);
nand U2174 (N_2174,In_2446,In_1121);
nor U2175 (N_2175,In_997,In_1570);
nand U2176 (N_2176,In_2431,In_2063);
nand U2177 (N_2177,In_1396,In_2177);
nor U2178 (N_2178,In_1513,In_2070);
or U2179 (N_2179,In_2076,In_2401);
and U2180 (N_2180,In_1386,In_258);
nor U2181 (N_2181,In_682,In_2031);
and U2182 (N_2182,In_587,In_745);
xnor U2183 (N_2183,In_1347,In_267);
or U2184 (N_2184,In_138,In_1362);
or U2185 (N_2185,In_1711,In_1807);
nor U2186 (N_2186,In_1812,In_420);
nor U2187 (N_2187,In_259,In_898);
or U2188 (N_2188,In_1196,In_1875);
xor U2189 (N_2189,In_1533,In_362);
xor U2190 (N_2190,In_642,In_1504);
nand U2191 (N_2191,In_181,In_164);
nor U2192 (N_2192,In_232,In_184);
or U2193 (N_2193,In_749,In_596);
and U2194 (N_2194,In_1736,In_1474);
nor U2195 (N_2195,In_481,In_1607);
nor U2196 (N_2196,In_1532,In_2486);
xor U2197 (N_2197,In_498,In_2240);
nor U2198 (N_2198,In_1036,In_489);
and U2199 (N_2199,In_493,In_2129);
and U2200 (N_2200,In_1445,In_1961);
nand U2201 (N_2201,In_2014,In_237);
nor U2202 (N_2202,In_1643,In_508);
and U2203 (N_2203,In_340,In_402);
nor U2204 (N_2204,In_1509,In_83);
and U2205 (N_2205,In_2103,In_1288);
nand U2206 (N_2206,In_246,In_1963);
and U2207 (N_2207,In_173,In_1809);
nor U2208 (N_2208,In_794,In_2472);
xor U2209 (N_2209,In_839,In_585);
xor U2210 (N_2210,In_1335,In_1957);
nand U2211 (N_2211,In_2166,In_1201);
or U2212 (N_2212,In_1549,In_273);
or U2213 (N_2213,In_926,In_816);
nand U2214 (N_2214,In_2241,In_2356);
and U2215 (N_2215,In_2178,In_1298);
xnor U2216 (N_2216,In_494,In_1465);
xnor U2217 (N_2217,In_1263,In_2067);
and U2218 (N_2218,In_687,In_1542);
and U2219 (N_2219,In_2362,In_1666);
or U2220 (N_2220,In_2161,In_1037);
and U2221 (N_2221,In_2114,In_308);
or U2222 (N_2222,In_1918,In_1378);
or U2223 (N_2223,In_470,In_837);
and U2224 (N_2224,In_1712,In_973);
xor U2225 (N_2225,In_930,In_1809);
nand U2226 (N_2226,In_1361,In_633);
nor U2227 (N_2227,In_542,In_1702);
nand U2228 (N_2228,In_1870,In_1410);
nor U2229 (N_2229,In_154,In_934);
or U2230 (N_2230,In_1676,In_1214);
nand U2231 (N_2231,In_827,In_684);
and U2232 (N_2232,In_700,In_558);
or U2233 (N_2233,In_74,In_543);
xor U2234 (N_2234,In_808,In_787);
and U2235 (N_2235,In_831,In_1893);
nand U2236 (N_2236,In_1830,In_1695);
nand U2237 (N_2237,In_825,In_1988);
xor U2238 (N_2238,In_1552,In_1990);
nor U2239 (N_2239,In_945,In_2399);
nor U2240 (N_2240,In_417,In_167);
or U2241 (N_2241,In_55,In_794);
nand U2242 (N_2242,In_440,In_1608);
xnor U2243 (N_2243,In_381,In_483);
and U2244 (N_2244,In_530,In_1980);
and U2245 (N_2245,In_993,In_927);
nand U2246 (N_2246,In_2434,In_1100);
and U2247 (N_2247,In_1346,In_2200);
nand U2248 (N_2248,In_205,In_1766);
nor U2249 (N_2249,In_1973,In_1513);
and U2250 (N_2250,In_89,In_888);
or U2251 (N_2251,In_1639,In_1414);
nand U2252 (N_2252,In_1959,In_2171);
nor U2253 (N_2253,In_578,In_1155);
nor U2254 (N_2254,In_2450,In_446);
nand U2255 (N_2255,In_1441,In_1759);
and U2256 (N_2256,In_1305,In_150);
xnor U2257 (N_2257,In_1378,In_819);
and U2258 (N_2258,In_656,In_1830);
nand U2259 (N_2259,In_902,In_86);
and U2260 (N_2260,In_611,In_362);
xor U2261 (N_2261,In_2237,In_1554);
xor U2262 (N_2262,In_838,In_1040);
xor U2263 (N_2263,In_484,In_2246);
xor U2264 (N_2264,In_1016,In_1299);
and U2265 (N_2265,In_2274,In_851);
or U2266 (N_2266,In_27,In_1660);
and U2267 (N_2267,In_1376,In_2365);
nor U2268 (N_2268,In_148,In_102);
nor U2269 (N_2269,In_1739,In_150);
or U2270 (N_2270,In_2245,In_470);
nand U2271 (N_2271,In_1080,In_1926);
and U2272 (N_2272,In_105,In_1265);
and U2273 (N_2273,In_14,In_2417);
or U2274 (N_2274,In_1269,In_1211);
nor U2275 (N_2275,In_1582,In_557);
and U2276 (N_2276,In_854,In_310);
xnor U2277 (N_2277,In_1063,In_1694);
and U2278 (N_2278,In_1791,In_1504);
xnor U2279 (N_2279,In_1198,In_1895);
or U2280 (N_2280,In_1996,In_320);
and U2281 (N_2281,In_232,In_405);
nor U2282 (N_2282,In_773,In_531);
and U2283 (N_2283,In_811,In_195);
nor U2284 (N_2284,In_802,In_1208);
xnor U2285 (N_2285,In_710,In_1415);
and U2286 (N_2286,In_1850,In_908);
nor U2287 (N_2287,In_982,In_760);
or U2288 (N_2288,In_1122,In_201);
and U2289 (N_2289,In_1989,In_323);
nand U2290 (N_2290,In_264,In_779);
and U2291 (N_2291,In_466,In_1924);
nand U2292 (N_2292,In_1335,In_710);
nand U2293 (N_2293,In_1373,In_1427);
nand U2294 (N_2294,In_1027,In_2340);
xor U2295 (N_2295,In_494,In_865);
or U2296 (N_2296,In_2436,In_1694);
nand U2297 (N_2297,In_846,In_267);
nand U2298 (N_2298,In_2152,In_704);
nand U2299 (N_2299,In_1032,In_2311);
xor U2300 (N_2300,In_8,In_811);
or U2301 (N_2301,In_1885,In_2444);
xnor U2302 (N_2302,In_1291,In_1806);
nand U2303 (N_2303,In_1984,In_1358);
nor U2304 (N_2304,In_2489,In_569);
or U2305 (N_2305,In_1794,In_1926);
nor U2306 (N_2306,In_870,In_1796);
xor U2307 (N_2307,In_2146,In_402);
or U2308 (N_2308,In_980,In_1085);
and U2309 (N_2309,In_913,In_2);
xor U2310 (N_2310,In_2155,In_822);
nand U2311 (N_2311,In_2069,In_1394);
and U2312 (N_2312,In_685,In_2328);
xnor U2313 (N_2313,In_340,In_2055);
xnor U2314 (N_2314,In_2483,In_1780);
nand U2315 (N_2315,In_1742,In_1734);
nand U2316 (N_2316,In_797,In_1664);
and U2317 (N_2317,In_2364,In_83);
and U2318 (N_2318,In_1582,In_795);
or U2319 (N_2319,In_1956,In_929);
nand U2320 (N_2320,In_1613,In_83);
xor U2321 (N_2321,In_299,In_137);
or U2322 (N_2322,In_1141,In_1656);
and U2323 (N_2323,In_2131,In_2386);
xor U2324 (N_2324,In_466,In_1974);
or U2325 (N_2325,In_786,In_767);
nand U2326 (N_2326,In_337,In_1023);
nand U2327 (N_2327,In_813,In_960);
xnor U2328 (N_2328,In_728,In_1913);
or U2329 (N_2329,In_1178,In_813);
xor U2330 (N_2330,In_1195,In_1048);
or U2331 (N_2331,In_87,In_296);
nand U2332 (N_2332,In_702,In_619);
and U2333 (N_2333,In_1334,In_1265);
nor U2334 (N_2334,In_2078,In_33);
and U2335 (N_2335,In_1667,In_2071);
nor U2336 (N_2336,In_1538,In_256);
nor U2337 (N_2337,In_958,In_256);
nor U2338 (N_2338,In_813,In_1816);
nor U2339 (N_2339,In_450,In_1359);
nand U2340 (N_2340,In_1519,In_1041);
and U2341 (N_2341,In_2385,In_655);
nand U2342 (N_2342,In_192,In_1699);
nand U2343 (N_2343,In_175,In_2002);
nor U2344 (N_2344,In_2449,In_1945);
nand U2345 (N_2345,In_1537,In_623);
nor U2346 (N_2346,In_2092,In_992);
nor U2347 (N_2347,In_2292,In_1453);
or U2348 (N_2348,In_1421,In_259);
and U2349 (N_2349,In_905,In_530);
xor U2350 (N_2350,In_1083,In_2424);
nand U2351 (N_2351,In_1759,In_702);
and U2352 (N_2352,In_330,In_322);
and U2353 (N_2353,In_1702,In_2458);
nand U2354 (N_2354,In_186,In_943);
nor U2355 (N_2355,In_69,In_529);
nand U2356 (N_2356,In_2434,In_2481);
nand U2357 (N_2357,In_314,In_1142);
nor U2358 (N_2358,In_1842,In_1366);
xor U2359 (N_2359,In_1930,In_1248);
or U2360 (N_2360,In_1428,In_2255);
nand U2361 (N_2361,In_583,In_2238);
nand U2362 (N_2362,In_79,In_996);
or U2363 (N_2363,In_1574,In_1299);
nor U2364 (N_2364,In_2251,In_1590);
xnor U2365 (N_2365,In_976,In_1736);
nor U2366 (N_2366,In_1030,In_878);
xor U2367 (N_2367,In_811,In_2032);
and U2368 (N_2368,In_1726,In_4);
nand U2369 (N_2369,In_947,In_1458);
or U2370 (N_2370,In_1891,In_1416);
nand U2371 (N_2371,In_1681,In_363);
or U2372 (N_2372,In_2215,In_566);
or U2373 (N_2373,In_1400,In_1175);
xnor U2374 (N_2374,In_210,In_1708);
and U2375 (N_2375,In_1010,In_2267);
nor U2376 (N_2376,In_868,In_608);
xnor U2377 (N_2377,In_1275,In_307);
and U2378 (N_2378,In_270,In_2);
and U2379 (N_2379,In_286,In_1462);
xor U2380 (N_2380,In_39,In_1414);
and U2381 (N_2381,In_838,In_2019);
nand U2382 (N_2382,In_2368,In_122);
xnor U2383 (N_2383,In_1931,In_1696);
nor U2384 (N_2384,In_183,In_685);
or U2385 (N_2385,In_1535,In_1278);
nand U2386 (N_2386,In_1565,In_470);
nor U2387 (N_2387,In_2211,In_272);
or U2388 (N_2388,In_690,In_1476);
nor U2389 (N_2389,In_436,In_2372);
nand U2390 (N_2390,In_2357,In_475);
or U2391 (N_2391,In_662,In_173);
nor U2392 (N_2392,In_1657,In_1226);
xor U2393 (N_2393,In_688,In_392);
nor U2394 (N_2394,In_1126,In_2203);
nand U2395 (N_2395,In_437,In_2416);
and U2396 (N_2396,In_2491,In_1085);
and U2397 (N_2397,In_1717,In_2161);
xnor U2398 (N_2398,In_678,In_1464);
xnor U2399 (N_2399,In_1765,In_2327);
nand U2400 (N_2400,In_2218,In_2091);
nor U2401 (N_2401,In_2141,In_74);
nor U2402 (N_2402,In_2031,In_228);
nor U2403 (N_2403,In_1503,In_986);
nand U2404 (N_2404,In_840,In_1783);
and U2405 (N_2405,In_705,In_787);
and U2406 (N_2406,In_2397,In_434);
xor U2407 (N_2407,In_30,In_110);
xor U2408 (N_2408,In_1905,In_355);
xnor U2409 (N_2409,In_949,In_1993);
nand U2410 (N_2410,In_2050,In_1862);
or U2411 (N_2411,In_2119,In_2166);
xnor U2412 (N_2412,In_294,In_310);
nor U2413 (N_2413,In_80,In_343);
or U2414 (N_2414,In_2013,In_1188);
nand U2415 (N_2415,In_576,In_1038);
nand U2416 (N_2416,In_339,In_205);
nand U2417 (N_2417,In_528,In_2324);
and U2418 (N_2418,In_376,In_26);
or U2419 (N_2419,In_1792,In_1681);
nand U2420 (N_2420,In_960,In_173);
or U2421 (N_2421,In_2099,In_2458);
or U2422 (N_2422,In_1420,In_1049);
nand U2423 (N_2423,In_2465,In_2141);
xnor U2424 (N_2424,In_666,In_1202);
nand U2425 (N_2425,In_1255,In_423);
nor U2426 (N_2426,In_1514,In_1173);
and U2427 (N_2427,In_1894,In_774);
nand U2428 (N_2428,In_1218,In_664);
nor U2429 (N_2429,In_312,In_944);
nand U2430 (N_2430,In_670,In_1221);
and U2431 (N_2431,In_1689,In_1455);
nor U2432 (N_2432,In_1103,In_2394);
xor U2433 (N_2433,In_1966,In_1025);
or U2434 (N_2434,In_1004,In_1280);
nor U2435 (N_2435,In_1936,In_2396);
nor U2436 (N_2436,In_572,In_810);
or U2437 (N_2437,In_561,In_1303);
nand U2438 (N_2438,In_1594,In_631);
nor U2439 (N_2439,In_1013,In_2467);
nand U2440 (N_2440,In_1057,In_1372);
xnor U2441 (N_2441,In_1010,In_2004);
and U2442 (N_2442,In_1752,In_1440);
nor U2443 (N_2443,In_432,In_2337);
xor U2444 (N_2444,In_831,In_1720);
xnor U2445 (N_2445,In_1289,In_2378);
nor U2446 (N_2446,In_1630,In_709);
and U2447 (N_2447,In_2143,In_2007);
nor U2448 (N_2448,In_909,In_1895);
nand U2449 (N_2449,In_96,In_441);
or U2450 (N_2450,In_673,In_1081);
or U2451 (N_2451,In_2256,In_1378);
or U2452 (N_2452,In_515,In_1553);
nor U2453 (N_2453,In_1543,In_154);
nand U2454 (N_2454,In_2229,In_1618);
xnor U2455 (N_2455,In_938,In_2185);
and U2456 (N_2456,In_1954,In_440);
or U2457 (N_2457,In_1168,In_622);
nor U2458 (N_2458,In_2483,In_152);
nor U2459 (N_2459,In_2140,In_907);
nor U2460 (N_2460,In_2430,In_1397);
and U2461 (N_2461,In_2016,In_794);
nand U2462 (N_2462,In_1991,In_2493);
and U2463 (N_2463,In_977,In_1878);
or U2464 (N_2464,In_2010,In_2345);
nand U2465 (N_2465,In_1246,In_2428);
or U2466 (N_2466,In_1018,In_1429);
nor U2467 (N_2467,In_2471,In_2283);
nand U2468 (N_2468,In_1537,In_584);
and U2469 (N_2469,In_2199,In_1729);
and U2470 (N_2470,In_973,In_1498);
and U2471 (N_2471,In_860,In_1592);
nor U2472 (N_2472,In_403,In_1530);
and U2473 (N_2473,In_18,In_2409);
xor U2474 (N_2474,In_1336,In_1519);
nor U2475 (N_2475,In_2151,In_850);
or U2476 (N_2476,In_1017,In_852);
xor U2477 (N_2477,In_1842,In_295);
nor U2478 (N_2478,In_624,In_1399);
xor U2479 (N_2479,In_1987,In_2102);
nand U2480 (N_2480,In_447,In_2409);
nor U2481 (N_2481,In_1026,In_1140);
nand U2482 (N_2482,In_2483,In_233);
xor U2483 (N_2483,In_229,In_222);
nand U2484 (N_2484,In_2092,In_2097);
nand U2485 (N_2485,In_995,In_100);
and U2486 (N_2486,In_1248,In_2267);
xnor U2487 (N_2487,In_1941,In_1127);
nand U2488 (N_2488,In_1385,In_2350);
nand U2489 (N_2489,In_1547,In_429);
nor U2490 (N_2490,In_1901,In_1868);
nor U2491 (N_2491,In_52,In_2023);
xnor U2492 (N_2492,In_1748,In_1498);
and U2493 (N_2493,In_1881,In_2470);
or U2494 (N_2494,In_2314,In_1136);
and U2495 (N_2495,In_1756,In_2377);
nand U2496 (N_2496,In_2441,In_182);
and U2497 (N_2497,In_634,In_1047);
nor U2498 (N_2498,In_2013,In_1852);
nor U2499 (N_2499,In_1997,In_2065);
xnor U2500 (N_2500,In_371,In_303);
nand U2501 (N_2501,In_2224,In_2041);
nor U2502 (N_2502,In_317,In_1444);
nand U2503 (N_2503,In_1558,In_561);
or U2504 (N_2504,In_315,In_1011);
nor U2505 (N_2505,In_1046,In_413);
xor U2506 (N_2506,In_1828,In_2348);
xor U2507 (N_2507,In_1351,In_886);
or U2508 (N_2508,In_714,In_916);
nand U2509 (N_2509,In_1589,In_2124);
nor U2510 (N_2510,In_1451,In_529);
or U2511 (N_2511,In_2486,In_2204);
or U2512 (N_2512,In_1856,In_383);
nand U2513 (N_2513,In_706,In_1);
nor U2514 (N_2514,In_1756,In_186);
nor U2515 (N_2515,In_2084,In_1605);
nand U2516 (N_2516,In_1167,In_1984);
and U2517 (N_2517,In_2177,In_92);
nor U2518 (N_2518,In_1188,In_269);
and U2519 (N_2519,In_2208,In_270);
nor U2520 (N_2520,In_2279,In_1664);
and U2521 (N_2521,In_1428,In_704);
nand U2522 (N_2522,In_1271,In_1172);
and U2523 (N_2523,In_2359,In_512);
nor U2524 (N_2524,In_1020,In_1365);
nor U2525 (N_2525,In_1162,In_813);
or U2526 (N_2526,In_2464,In_2409);
nand U2527 (N_2527,In_1782,In_131);
nand U2528 (N_2528,In_2442,In_2048);
or U2529 (N_2529,In_2072,In_40);
nor U2530 (N_2530,In_1745,In_297);
and U2531 (N_2531,In_805,In_1798);
nor U2532 (N_2532,In_630,In_1822);
and U2533 (N_2533,In_89,In_76);
nor U2534 (N_2534,In_1726,In_1993);
or U2535 (N_2535,In_762,In_1978);
nand U2536 (N_2536,In_274,In_931);
nor U2537 (N_2537,In_844,In_237);
and U2538 (N_2538,In_369,In_1016);
nor U2539 (N_2539,In_1035,In_1574);
or U2540 (N_2540,In_2196,In_979);
nor U2541 (N_2541,In_2499,In_2096);
nor U2542 (N_2542,In_2466,In_1389);
nor U2543 (N_2543,In_757,In_1175);
xor U2544 (N_2544,In_2094,In_784);
nor U2545 (N_2545,In_983,In_38);
nor U2546 (N_2546,In_851,In_382);
and U2547 (N_2547,In_2260,In_1462);
xor U2548 (N_2548,In_993,In_467);
or U2549 (N_2549,In_395,In_558);
or U2550 (N_2550,In_1203,In_1503);
nand U2551 (N_2551,In_1541,In_125);
nor U2552 (N_2552,In_1196,In_1736);
or U2553 (N_2553,In_2383,In_372);
or U2554 (N_2554,In_443,In_1195);
xnor U2555 (N_2555,In_874,In_1489);
and U2556 (N_2556,In_2140,In_2311);
nand U2557 (N_2557,In_2092,In_631);
xnor U2558 (N_2558,In_959,In_2193);
nor U2559 (N_2559,In_1867,In_2250);
nor U2560 (N_2560,In_822,In_550);
nand U2561 (N_2561,In_2095,In_1639);
or U2562 (N_2562,In_2414,In_2475);
nor U2563 (N_2563,In_634,In_490);
xor U2564 (N_2564,In_1686,In_1218);
xor U2565 (N_2565,In_1028,In_2430);
nand U2566 (N_2566,In_953,In_2481);
nor U2567 (N_2567,In_2257,In_651);
or U2568 (N_2568,In_2033,In_1933);
or U2569 (N_2569,In_1602,In_169);
nor U2570 (N_2570,In_1756,In_785);
and U2571 (N_2571,In_2131,In_1354);
nand U2572 (N_2572,In_1943,In_528);
and U2573 (N_2573,In_873,In_1389);
and U2574 (N_2574,In_2079,In_1103);
xor U2575 (N_2575,In_1440,In_918);
and U2576 (N_2576,In_2315,In_1267);
nor U2577 (N_2577,In_1284,In_2384);
and U2578 (N_2578,In_1619,In_741);
xor U2579 (N_2579,In_574,In_45);
nor U2580 (N_2580,In_226,In_2299);
nand U2581 (N_2581,In_1199,In_1818);
xnor U2582 (N_2582,In_158,In_2070);
nor U2583 (N_2583,In_2225,In_896);
xor U2584 (N_2584,In_128,In_537);
nand U2585 (N_2585,In_805,In_2085);
nand U2586 (N_2586,In_2182,In_1762);
or U2587 (N_2587,In_2199,In_1327);
nand U2588 (N_2588,In_68,In_2190);
nor U2589 (N_2589,In_1436,In_62);
nand U2590 (N_2590,In_1577,In_721);
xor U2591 (N_2591,In_962,In_2131);
nand U2592 (N_2592,In_1755,In_1646);
or U2593 (N_2593,In_1666,In_758);
or U2594 (N_2594,In_1657,In_2323);
and U2595 (N_2595,In_1448,In_2032);
nor U2596 (N_2596,In_1291,In_121);
nand U2597 (N_2597,In_1476,In_1839);
or U2598 (N_2598,In_987,In_43);
nand U2599 (N_2599,In_1078,In_1226);
nand U2600 (N_2600,In_83,In_922);
or U2601 (N_2601,In_1177,In_1034);
or U2602 (N_2602,In_372,In_1624);
or U2603 (N_2603,In_402,In_1852);
nor U2604 (N_2604,In_1405,In_774);
and U2605 (N_2605,In_1820,In_464);
nand U2606 (N_2606,In_1208,In_1005);
xor U2607 (N_2607,In_68,In_2093);
nand U2608 (N_2608,In_405,In_2430);
or U2609 (N_2609,In_1720,In_1187);
and U2610 (N_2610,In_1959,In_968);
nor U2611 (N_2611,In_385,In_1006);
nor U2612 (N_2612,In_1658,In_2029);
xor U2613 (N_2613,In_1284,In_1926);
nor U2614 (N_2614,In_537,In_1080);
nor U2615 (N_2615,In_1362,In_1895);
xor U2616 (N_2616,In_1577,In_110);
or U2617 (N_2617,In_1739,In_937);
or U2618 (N_2618,In_1702,In_578);
nor U2619 (N_2619,In_1640,In_459);
nor U2620 (N_2620,In_2083,In_215);
and U2621 (N_2621,In_1684,In_2292);
xnor U2622 (N_2622,In_654,In_2278);
nand U2623 (N_2623,In_1466,In_2088);
xnor U2624 (N_2624,In_249,In_1641);
xor U2625 (N_2625,In_1454,In_2322);
nand U2626 (N_2626,In_1967,In_1435);
nand U2627 (N_2627,In_1206,In_923);
and U2628 (N_2628,In_1871,In_24);
or U2629 (N_2629,In_2041,In_2067);
and U2630 (N_2630,In_292,In_2284);
nand U2631 (N_2631,In_1263,In_738);
or U2632 (N_2632,In_1643,In_1087);
xnor U2633 (N_2633,In_643,In_2281);
xor U2634 (N_2634,In_2091,In_1500);
nand U2635 (N_2635,In_344,In_535);
nor U2636 (N_2636,In_1104,In_2158);
nand U2637 (N_2637,In_205,In_2076);
or U2638 (N_2638,In_1672,In_1038);
and U2639 (N_2639,In_530,In_324);
xnor U2640 (N_2640,In_1183,In_1847);
nor U2641 (N_2641,In_1242,In_19);
nor U2642 (N_2642,In_475,In_1565);
and U2643 (N_2643,In_582,In_210);
or U2644 (N_2644,In_649,In_236);
nor U2645 (N_2645,In_2380,In_745);
and U2646 (N_2646,In_1765,In_2097);
and U2647 (N_2647,In_2247,In_1996);
or U2648 (N_2648,In_1032,In_1984);
nand U2649 (N_2649,In_1371,In_1410);
and U2650 (N_2650,In_76,In_1375);
or U2651 (N_2651,In_535,In_257);
nand U2652 (N_2652,In_20,In_2152);
or U2653 (N_2653,In_44,In_1475);
nor U2654 (N_2654,In_1081,In_2412);
and U2655 (N_2655,In_1020,In_633);
xnor U2656 (N_2656,In_2293,In_907);
and U2657 (N_2657,In_2081,In_1350);
nor U2658 (N_2658,In_1338,In_1614);
xnor U2659 (N_2659,In_1036,In_2137);
nand U2660 (N_2660,In_1899,In_34);
nor U2661 (N_2661,In_536,In_1959);
nor U2662 (N_2662,In_1585,In_180);
nand U2663 (N_2663,In_1893,In_82);
xor U2664 (N_2664,In_746,In_1128);
xor U2665 (N_2665,In_2322,In_1334);
nand U2666 (N_2666,In_478,In_1373);
nor U2667 (N_2667,In_984,In_2050);
or U2668 (N_2668,In_1358,In_1970);
nand U2669 (N_2669,In_2252,In_720);
and U2670 (N_2670,In_1497,In_1735);
nand U2671 (N_2671,In_1038,In_481);
or U2672 (N_2672,In_2114,In_1998);
or U2673 (N_2673,In_1935,In_217);
xnor U2674 (N_2674,In_1689,In_2328);
or U2675 (N_2675,In_1414,In_2469);
nand U2676 (N_2676,In_778,In_377);
nand U2677 (N_2677,In_831,In_1915);
and U2678 (N_2678,In_2272,In_557);
and U2679 (N_2679,In_1334,In_1491);
and U2680 (N_2680,In_1940,In_761);
nor U2681 (N_2681,In_628,In_1505);
nand U2682 (N_2682,In_215,In_934);
xnor U2683 (N_2683,In_950,In_79);
or U2684 (N_2684,In_1847,In_262);
nor U2685 (N_2685,In_1634,In_204);
nand U2686 (N_2686,In_1460,In_1163);
and U2687 (N_2687,In_1134,In_1456);
or U2688 (N_2688,In_1570,In_2005);
or U2689 (N_2689,In_860,In_1636);
or U2690 (N_2690,In_1365,In_1843);
and U2691 (N_2691,In_1498,In_1681);
nor U2692 (N_2692,In_1054,In_2198);
or U2693 (N_2693,In_1741,In_1264);
nor U2694 (N_2694,In_282,In_577);
nor U2695 (N_2695,In_560,In_1506);
nand U2696 (N_2696,In_943,In_38);
and U2697 (N_2697,In_74,In_2241);
and U2698 (N_2698,In_300,In_2382);
xnor U2699 (N_2699,In_1587,In_1049);
nand U2700 (N_2700,In_2175,In_1460);
nand U2701 (N_2701,In_839,In_20);
and U2702 (N_2702,In_813,In_405);
and U2703 (N_2703,In_995,In_258);
nand U2704 (N_2704,In_2002,In_1649);
and U2705 (N_2705,In_1060,In_681);
nor U2706 (N_2706,In_1734,In_1689);
and U2707 (N_2707,In_2344,In_2196);
and U2708 (N_2708,In_454,In_208);
or U2709 (N_2709,In_944,In_372);
nor U2710 (N_2710,In_1941,In_1024);
nor U2711 (N_2711,In_1931,In_191);
nor U2712 (N_2712,In_811,In_1359);
nor U2713 (N_2713,In_129,In_232);
or U2714 (N_2714,In_1936,In_2231);
xnor U2715 (N_2715,In_1198,In_716);
or U2716 (N_2716,In_611,In_1509);
or U2717 (N_2717,In_820,In_1293);
or U2718 (N_2718,In_1166,In_1101);
and U2719 (N_2719,In_721,In_68);
and U2720 (N_2720,In_1469,In_2028);
and U2721 (N_2721,In_1318,In_2367);
xnor U2722 (N_2722,In_2184,In_927);
nand U2723 (N_2723,In_2206,In_183);
or U2724 (N_2724,In_2038,In_125);
or U2725 (N_2725,In_2381,In_761);
and U2726 (N_2726,In_141,In_2334);
nor U2727 (N_2727,In_14,In_2331);
xor U2728 (N_2728,In_195,In_1243);
and U2729 (N_2729,In_1521,In_2227);
nand U2730 (N_2730,In_1675,In_536);
or U2731 (N_2731,In_809,In_347);
xor U2732 (N_2732,In_1373,In_2346);
and U2733 (N_2733,In_277,In_314);
and U2734 (N_2734,In_1870,In_1011);
xor U2735 (N_2735,In_1988,In_2289);
xnor U2736 (N_2736,In_2407,In_896);
xor U2737 (N_2737,In_1384,In_1548);
nand U2738 (N_2738,In_1167,In_1455);
and U2739 (N_2739,In_580,In_2164);
or U2740 (N_2740,In_1818,In_1730);
xnor U2741 (N_2741,In_366,In_1709);
nor U2742 (N_2742,In_1529,In_2104);
and U2743 (N_2743,In_869,In_2002);
nor U2744 (N_2744,In_1635,In_634);
or U2745 (N_2745,In_1646,In_1856);
and U2746 (N_2746,In_1989,In_361);
nor U2747 (N_2747,In_450,In_1276);
xnor U2748 (N_2748,In_1589,In_268);
xor U2749 (N_2749,In_994,In_1039);
nor U2750 (N_2750,In_1798,In_342);
nor U2751 (N_2751,In_1836,In_150);
or U2752 (N_2752,In_1257,In_1553);
xor U2753 (N_2753,In_1323,In_932);
xor U2754 (N_2754,In_1183,In_1818);
nor U2755 (N_2755,In_1086,In_1178);
xnor U2756 (N_2756,In_517,In_1327);
nand U2757 (N_2757,In_1911,In_520);
nand U2758 (N_2758,In_850,In_2298);
and U2759 (N_2759,In_556,In_1607);
and U2760 (N_2760,In_771,In_2430);
nor U2761 (N_2761,In_1155,In_2234);
or U2762 (N_2762,In_792,In_2214);
nand U2763 (N_2763,In_744,In_71);
nor U2764 (N_2764,In_976,In_2019);
nand U2765 (N_2765,In_89,In_1972);
and U2766 (N_2766,In_1978,In_2078);
and U2767 (N_2767,In_2087,In_763);
nor U2768 (N_2768,In_1556,In_777);
and U2769 (N_2769,In_1273,In_285);
or U2770 (N_2770,In_2166,In_468);
nand U2771 (N_2771,In_452,In_769);
xnor U2772 (N_2772,In_449,In_1313);
xnor U2773 (N_2773,In_1033,In_1854);
or U2774 (N_2774,In_2465,In_1262);
nor U2775 (N_2775,In_1002,In_2224);
nand U2776 (N_2776,In_171,In_116);
and U2777 (N_2777,In_8,In_2388);
nor U2778 (N_2778,In_1122,In_337);
or U2779 (N_2779,In_1992,In_677);
nor U2780 (N_2780,In_1107,In_2142);
xor U2781 (N_2781,In_20,In_2334);
xor U2782 (N_2782,In_685,In_1437);
and U2783 (N_2783,In_249,In_2414);
and U2784 (N_2784,In_1841,In_1625);
nand U2785 (N_2785,In_751,In_1193);
or U2786 (N_2786,In_1600,In_1996);
and U2787 (N_2787,In_1898,In_1540);
nor U2788 (N_2788,In_899,In_162);
and U2789 (N_2789,In_2417,In_1661);
nand U2790 (N_2790,In_487,In_1069);
xnor U2791 (N_2791,In_487,In_530);
or U2792 (N_2792,In_1242,In_448);
or U2793 (N_2793,In_695,In_357);
nor U2794 (N_2794,In_1848,In_258);
xnor U2795 (N_2795,In_1209,In_233);
or U2796 (N_2796,In_608,In_2313);
and U2797 (N_2797,In_1527,In_2232);
and U2798 (N_2798,In_1318,In_1468);
xor U2799 (N_2799,In_2,In_317);
nand U2800 (N_2800,In_1734,In_2200);
nand U2801 (N_2801,In_2335,In_1);
nor U2802 (N_2802,In_1447,In_1117);
nand U2803 (N_2803,In_189,In_2228);
xor U2804 (N_2804,In_1826,In_1106);
and U2805 (N_2805,In_451,In_2187);
or U2806 (N_2806,In_2185,In_122);
and U2807 (N_2807,In_1400,In_486);
xor U2808 (N_2808,In_1422,In_837);
and U2809 (N_2809,In_1844,In_2388);
nand U2810 (N_2810,In_1676,In_835);
nand U2811 (N_2811,In_2357,In_1371);
and U2812 (N_2812,In_2011,In_2203);
nand U2813 (N_2813,In_2446,In_970);
nor U2814 (N_2814,In_2443,In_197);
or U2815 (N_2815,In_2326,In_2415);
nand U2816 (N_2816,In_1253,In_1084);
xor U2817 (N_2817,In_1588,In_145);
nand U2818 (N_2818,In_389,In_1272);
xnor U2819 (N_2819,In_728,In_489);
xor U2820 (N_2820,In_506,In_1307);
and U2821 (N_2821,In_957,In_1733);
or U2822 (N_2822,In_295,In_196);
or U2823 (N_2823,In_153,In_1638);
nor U2824 (N_2824,In_2464,In_1762);
or U2825 (N_2825,In_1597,In_942);
nor U2826 (N_2826,In_1957,In_1893);
xnor U2827 (N_2827,In_487,In_1281);
nand U2828 (N_2828,In_2274,In_593);
and U2829 (N_2829,In_1351,In_2404);
and U2830 (N_2830,In_1258,In_1818);
xnor U2831 (N_2831,In_1531,In_1351);
or U2832 (N_2832,In_383,In_2239);
xor U2833 (N_2833,In_273,In_272);
or U2834 (N_2834,In_116,In_2103);
and U2835 (N_2835,In_1349,In_35);
or U2836 (N_2836,In_1183,In_917);
and U2837 (N_2837,In_395,In_1630);
nor U2838 (N_2838,In_2421,In_1267);
nand U2839 (N_2839,In_1758,In_421);
xor U2840 (N_2840,In_553,In_445);
and U2841 (N_2841,In_494,In_261);
or U2842 (N_2842,In_1385,In_2337);
nor U2843 (N_2843,In_1669,In_2173);
nand U2844 (N_2844,In_319,In_862);
or U2845 (N_2845,In_628,In_2344);
nor U2846 (N_2846,In_127,In_938);
and U2847 (N_2847,In_838,In_936);
and U2848 (N_2848,In_1473,In_2290);
or U2849 (N_2849,In_523,In_1643);
and U2850 (N_2850,In_2439,In_1385);
nand U2851 (N_2851,In_688,In_421);
nor U2852 (N_2852,In_2053,In_1440);
and U2853 (N_2853,In_2259,In_1339);
nand U2854 (N_2854,In_1373,In_2369);
nor U2855 (N_2855,In_2232,In_2210);
nor U2856 (N_2856,In_1306,In_1281);
xor U2857 (N_2857,In_2352,In_957);
nand U2858 (N_2858,In_1506,In_741);
or U2859 (N_2859,In_1903,In_926);
and U2860 (N_2860,In_616,In_548);
and U2861 (N_2861,In_1237,In_879);
nor U2862 (N_2862,In_638,In_924);
xnor U2863 (N_2863,In_2121,In_2095);
xor U2864 (N_2864,In_851,In_1442);
nand U2865 (N_2865,In_1140,In_137);
or U2866 (N_2866,In_380,In_106);
nor U2867 (N_2867,In_1371,In_1879);
xnor U2868 (N_2868,In_1027,In_1771);
nand U2869 (N_2869,In_1229,In_1974);
and U2870 (N_2870,In_717,In_558);
and U2871 (N_2871,In_724,In_1274);
and U2872 (N_2872,In_471,In_2437);
nand U2873 (N_2873,In_705,In_2413);
nor U2874 (N_2874,In_649,In_2391);
or U2875 (N_2875,In_1291,In_22);
nor U2876 (N_2876,In_2359,In_1322);
and U2877 (N_2877,In_2154,In_893);
nand U2878 (N_2878,In_1487,In_1180);
and U2879 (N_2879,In_257,In_1769);
nor U2880 (N_2880,In_2094,In_921);
xor U2881 (N_2881,In_429,In_535);
nor U2882 (N_2882,In_2402,In_629);
xnor U2883 (N_2883,In_1810,In_1716);
nor U2884 (N_2884,In_345,In_938);
nor U2885 (N_2885,In_1780,In_56);
xor U2886 (N_2886,In_1717,In_2297);
nor U2887 (N_2887,In_854,In_2149);
xnor U2888 (N_2888,In_1548,In_1070);
nand U2889 (N_2889,In_1326,In_524);
and U2890 (N_2890,In_1659,In_1572);
nand U2891 (N_2891,In_193,In_2342);
xnor U2892 (N_2892,In_2274,In_353);
and U2893 (N_2893,In_994,In_1995);
xor U2894 (N_2894,In_2254,In_929);
nor U2895 (N_2895,In_575,In_454);
xor U2896 (N_2896,In_2071,In_1107);
xor U2897 (N_2897,In_100,In_2108);
xor U2898 (N_2898,In_1035,In_678);
nand U2899 (N_2899,In_947,In_283);
xor U2900 (N_2900,In_2355,In_40);
or U2901 (N_2901,In_1123,In_811);
xor U2902 (N_2902,In_597,In_215);
and U2903 (N_2903,In_716,In_824);
xor U2904 (N_2904,In_373,In_1536);
or U2905 (N_2905,In_114,In_2333);
nor U2906 (N_2906,In_1863,In_863);
and U2907 (N_2907,In_1879,In_1865);
xnor U2908 (N_2908,In_466,In_553);
nand U2909 (N_2909,In_1533,In_1080);
or U2910 (N_2910,In_596,In_2130);
xor U2911 (N_2911,In_1563,In_362);
or U2912 (N_2912,In_92,In_379);
xor U2913 (N_2913,In_1892,In_178);
nand U2914 (N_2914,In_1843,In_2162);
nand U2915 (N_2915,In_915,In_224);
nor U2916 (N_2916,In_2487,In_137);
and U2917 (N_2917,In_1428,In_635);
or U2918 (N_2918,In_153,In_554);
and U2919 (N_2919,In_1568,In_1080);
and U2920 (N_2920,In_1813,In_733);
xnor U2921 (N_2921,In_1049,In_181);
xor U2922 (N_2922,In_513,In_2480);
nor U2923 (N_2923,In_550,In_1306);
xnor U2924 (N_2924,In_164,In_1054);
nor U2925 (N_2925,In_62,In_1241);
and U2926 (N_2926,In_978,In_1266);
and U2927 (N_2927,In_880,In_2168);
or U2928 (N_2928,In_635,In_1838);
or U2929 (N_2929,In_232,In_1592);
nand U2930 (N_2930,In_265,In_1337);
xnor U2931 (N_2931,In_2428,In_244);
xor U2932 (N_2932,In_1436,In_790);
nor U2933 (N_2933,In_925,In_1082);
nand U2934 (N_2934,In_142,In_1505);
nor U2935 (N_2935,In_1262,In_1880);
nor U2936 (N_2936,In_887,In_631);
nor U2937 (N_2937,In_1714,In_346);
xor U2938 (N_2938,In_1085,In_288);
nand U2939 (N_2939,In_2344,In_369);
nand U2940 (N_2940,In_1197,In_226);
nor U2941 (N_2941,In_597,In_65);
xor U2942 (N_2942,In_1444,In_1485);
or U2943 (N_2943,In_2007,In_1730);
nor U2944 (N_2944,In_2436,In_129);
or U2945 (N_2945,In_1148,In_1081);
nand U2946 (N_2946,In_665,In_771);
or U2947 (N_2947,In_645,In_1659);
nand U2948 (N_2948,In_1138,In_1970);
or U2949 (N_2949,In_958,In_322);
xor U2950 (N_2950,In_1923,In_2458);
and U2951 (N_2951,In_1319,In_1213);
nand U2952 (N_2952,In_528,In_1016);
nand U2953 (N_2953,In_786,In_959);
xor U2954 (N_2954,In_1052,In_1478);
xor U2955 (N_2955,In_382,In_757);
xor U2956 (N_2956,In_809,In_926);
nor U2957 (N_2957,In_68,In_44);
xor U2958 (N_2958,In_1551,In_2277);
nor U2959 (N_2959,In_109,In_737);
nand U2960 (N_2960,In_1784,In_2474);
nor U2961 (N_2961,In_390,In_2494);
xor U2962 (N_2962,In_574,In_705);
and U2963 (N_2963,In_514,In_2103);
or U2964 (N_2964,In_1033,In_252);
nor U2965 (N_2965,In_2386,In_1229);
xor U2966 (N_2966,In_1744,In_2306);
nor U2967 (N_2967,In_573,In_96);
and U2968 (N_2968,In_666,In_2420);
xor U2969 (N_2969,In_1805,In_154);
and U2970 (N_2970,In_2064,In_1103);
nor U2971 (N_2971,In_1018,In_2163);
and U2972 (N_2972,In_689,In_1571);
xor U2973 (N_2973,In_431,In_2183);
nand U2974 (N_2974,In_557,In_1214);
xnor U2975 (N_2975,In_2142,In_414);
xnor U2976 (N_2976,In_1260,In_2029);
or U2977 (N_2977,In_2419,In_2193);
and U2978 (N_2978,In_2478,In_1831);
xnor U2979 (N_2979,In_1353,In_1724);
nor U2980 (N_2980,In_966,In_1155);
nand U2981 (N_2981,In_511,In_400);
nor U2982 (N_2982,In_2252,In_1870);
and U2983 (N_2983,In_1651,In_346);
xor U2984 (N_2984,In_281,In_1565);
xnor U2985 (N_2985,In_1788,In_124);
or U2986 (N_2986,In_1654,In_321);
nand U2987 (N_2987,In_723,In_1728);
or U2988 (N_2988,In_1563,In_337);
nor U2989 (N_2989,In_2324,In_2085);
and U2990 (N_2990,In_1317,In_594);
or U2991 (N_2991,In_972,In_1858);
nand U2992 (N_2992,In_1262,In_1588);
xnor U2993 (N_2993,In_1705,In_82);
or U2994 (N_2994,In_978,In_2180);
nor U2995 (N_2995,In_2383,In_2073);
nor U2996 (N_2996,In_1821,In_1467);
nand U2997 (N_2997,In_2185,In_2319);
nand U2998 (N_2998,In_2046,In_1204);
xnor U2999 (N_2999,In_349,In_1532);
and U3000 (N_3000,In_429,In_309);
nor U3001 (N_3001,In_1866,In_1994);
nand U3002 (N_3002,In_1488,In_2282);
nor U3003 (N_3003,In_836,In_2204);
or U3004 (N_3004,In_1733,In_881);
nand U3005 (N_3005,In_1690,In_2312);
or U3006 (N_3006,In_196,In_1054);
xnor U3007 (N_3007,In_103,In_765);
xor U3008 (N_3008,In_709,In_430);
and U3009 (N_3009,In_2020,In_1100);
and U3010 (N_3010,In_1161,In_1629);
and U3011 (N_3011,In_25,In_462);
and U3012 (N_3012,In_1965,In_2106);
and U3013 (N_3013,In_1631,In_637);
nor U3014 (N_3014,In_1070,In_1754);
or U3015 (N_3015,In_905,In_1120);
nor U3016 (N_3016,In_1136,In_2154);
nor U3017 (N_3017,In_2495,In_650);
and U3018 (N_3018,In_236,In_1394);
and U3019 (N_3019,In_1953,In_1122);
and U3020 (N_3020,In_622,In_2418);
xnor U3021 (N_3021,In_433,In_1600);
or U3022 (N_3022,In_976,In_2088);
and U3023 (N_3023,In_631,In_2414);
xor U3024 (N_3024,In_2173,In_1899);
nand U3025 (N_3025,In_93,In_1137);
nor U3026 (N_3026,In_2077,In_2319);
nand U3027 (N_3027,In_121,In_426);
xor U3028 (N_3028,In_2331,In_416);
or U3029 (N_3029,In_1202,In_817);
nand U3030 (N_3030,In_1749,In_1814);
nor U3031 (N_3031,In_657,In_522);
nand U3032 (N_3032,In_1599,In_2373);
and U3033 (N_3033,In_436,In_1353);
or U3034 (N_3034,In_15,In_2181);
or U3035 (N_3035,In_301,In_68);
nor U3036 (N_3036,In_2040,In_901);
and U3037 (N_3037,In_461,In_363);
and U3038 (N_3038,In_41,In_157);
xor U3039 (N_3039,In_164,In_643);
and U3040 (N_3040,In_1886,In_1128);
xor U3041 (N_3041,In_1936,In_1898);
nand U3042 (N_3042,In_481,In_2075);
nand U3043 (N_3043,In_2024,In_934);
and U3044 (N_3044,In_1071,In_700);
and U3045 (N_3045,In_1428,In_140);
xor U3046 (N_3046,In_1269,In_687);
and U3047 (N_3047,In_2327,In_703);
and U3048 (N_3048,In_895,In_1875);
nand U3049 (N_3049,In_1270,In_662);
nand U3050 (N_3050,In_1916,In_930);
or U3051 (N_3051,In_988,In_1548);
and U3052 (N_3052,In_922,In_2458);
or U3053 (N_3053,In_2139,In_2150);
nor U3054 (N_3054,In_1165,In_86);
nor U3055 (N_3055,In_1891,In_109);
nand U3056 (N_3056,In_2356,In_2425);
nand U3057 (N_3057,In_2405,In_607);
or U3058 (N_3058,In_536,In_415);
nor U3059 (N_3059,In_1642,In_702);
or U3060 (N_3060,In_2134,In_1469);
nand U3061 (N_3061,In_2251,In_1262);
nor U3062 (N_3062,In_1363,In_766);
nand U3063 (N_3063,In_626,In_1249);
nand U3064 (N_3064,In_306,In_1084);
nor U3065 (N_3065,In_603,In_1329);
xnor U3066 (N_3066,In_1708,In_1955);
and U3067 (N_3067,In_132,In_578);
xnor U3068 (N_3068,In_1254,In_2130);
and U3069 (N_3069,In_2475,In_1305);
nor U3070 (N_3070,In_1776,In_1560);
xnor U3071 (N_3071,In_151,In_411);
xor U3072 (N_3072,In_1407,In_1597);
nand U3073 (N_3073,In_726,In_40);
and U3074 (N_3074,In_1151,In_1908);
nand U3075 (N_3075,In_631,In_798);
nand U3076 (N_3076,In_713,In_210);
xnor U3077 (N_3077,In_1915,In_957);
nand U3078 (N_3078,In_1472,In_1207);
nor U3079 (N_3079,In_728,In_380);
xor U3080 (N_3080,In_1076,In_1177);
nor U3081 (N_3081,In_1244,In_2163);
nand U3082 (N_3082,In_90,In_1723);
nand U3083 (N_3083,In_424,In_1757);
xor U3084 (N_3084,In_218,In_13);
or U3085 (N_3085,In_1191,In_1746);
or U3086 (N_3086,In_1149,In_2040);
xor U3087 (N_3087,In_66,In_1018);
and U3088 (N_3088,In_744,In_2178);
or U3089 (N_3089,In_2,In_3);
or U3090 (N_3090,In_2232,In_1497);
or U3091 (N_3091,In_1304,In_581);
and U3092 (N_3092,In_2455,In_1064);
and U3093 (N_3093,In_34,In_2420);
or U3094 (N_3094,In_2484,In_641);
xor U3095 (N_3095,In_1228,In_1383);
xnor U3096 (N_3096,In_347,In_2465);
nor U3097 (N_3097,In_1360,In_2003);
xnor U3098 (N_3098,In_644,In_1653);
or U3099 (N_3099,In_1402,In_1325);
xnor U3100 (N_3100,In_2426,In_1768);
nor U3101 (N_3101,In_2189,In_559);
xor U3102 (N_3102,In_989,In_1905);
nor U3103 (N_3103,In_456,In_2384);
or U3104 (N_3104,In_556,In_455);
nand U3105 (N_3105,In_864,In_326);
nor U3106 (N_3106,In_1674,In_263);
nand U3107 (N_3107,In_2056,In_2080);
nand U3108 (N_3108,In_1369,In_1077);
nand U3109 (N_3109,In_2227,In_1836);
xnor U3110 (N_3110,In_850,In_1605);
and U3111 (N_3111,In_296,In_1760);
nor U3112 (N_3112,In_1597,In_2104);
or U3113 (N_3113,In_351,In_1592);
nand U3114 (N_3114,In_137,In_1527);
nor U3115 (N_3115,In_2162,In_1339);
xor U3116 (N_3116,In_157,In_2198);
xnor U3117 (N_3117,In_1138,In_1208);
and U3118 (N_3118,In_2459,In_2217);
xor U3119 (N_3119,In_283,In_1272);
nor U3120 (N_3120,In_1897,In_2342);
nand U3121 (N_3121,In_262,In_1868);
nand U3122 (N_3122,In_1022,In_483);
nor U3123 (N_3123,In_194,In_1226);
or U3124 (N_3124,In_1194,In_686);
nand U3125 (N_3125,In_214,In_330);
nand U3126 (N_3126,In_1953,In_361);
nor U3127 (N_3127,In_1144,In_1452);
and U3128 (N_3128,In_720,In_1782);
nand U3129 (N_3129,In_1997,In_340);
nand U3130 (N_3130,In_443,In_538);
or U3131 (N_3131,In_2248,In_2032);
and U3132 (N_3132,In_344,In_1065);
or U3133 (N_3133,In_941,In_1130);
or U3134 (N_3134,In_486,In_1231);
xor U3135 (N_3135,In_790,In_2044);
xor U3136 (N_3136,In_943,In_2307);
nor U3137 (N_3137,In_2474,In_2486);
nor U3138 (N_3138,In_2003,In_628);
and U3139 (N_3139,In_382,In_2164);
or U3140 (N_3140,In_276,In_1331);
and U3141 (N_3141,In_71,In_229);
and U3142 (N_3142,In_113,In_1102);
or U3143 (N_3143,In_1871,In_688);
nor U3144 (N_3144,In_712,In_428);
nand U3145 (N_3145,In_846,In_302);
nand U3146 (N_3146,In_1045,In_1683);
nor U3147 (N_3147,In_2297,In_64);
nor U3148 (N_3148,In_1322,In_1789);
xor U3149 (N_3149,In_14,In_937);
nor U3150 (N_3150,In_1142,In_1406);
or U3151 (N_3151,In_1425,In_991);
xnor U3152 (N_3152,In_2057,In_262);
or U3153 (N_3153,In_1076,In_680);
xor U3154 (N_3154,In_953,In_1489);
or U3155 (N_3155,In_436,In_1797);
nand U3156 (N_3156,In_1264,In_507);
xnor U3157 (N_3157,In_2407,In_40);
nor U3158 (N_3158,In_612,In_1370);
nand U3159 (N_3159,In_1711,In_2386);
or U3160 (N_3160,In_833,In_1839);
nand U3161 (N_3161,In_1168,In_1498);
nand U3162 (N_3162,In_2098,In_219);
or U3163 (N_3163,In_1713,In_1583);
nor U3164 (N_3164,In_715,In_1698);
or U3165 (N_3165,In_2096,In_2155);
and U3166 (N_3166,In_2422,In_1599);
and U3167 (N_3167,In_2198,In_191);
or U3168 (N_3168,In_1787,In_1496);
nor U3169 (N_3169,In_2308,In_2493);
xor U3170 (N_3170,In_1806,In_1323);
or U3171 (N_3171,In_185,In_117);
and U3172 (N_3172,In_2374,In_736);
and U3173 (N_3173,In_1146,In_1377);
or U3174 (N_3174,In_594,In_1545);
nand U3175 (N_3175,In_87,In_867);
or U3176 (N_3176,In_2335,In_1703);
xor U3177 (N_3177,In_1966,In_1343);
nand U3178 (N_3178,In_751,In_1796);
or U3179 (N_3179,In_1586,In_2340);
xor U3180 (N_3180,In_1181,In_2435);
xor U3181 (N_3181,In_1998,In_835);
xor U3182 (N_3182,In_1416,In_1720);
nand U3183 (N_3183,In_2256,In_2037);
nor U3184 (N_3184,In_2049,In_680);
or U3185 (N_3185,In_2396,In_1209);
nor U3186 (N_3186,In_517,In_1246);
or U3187 (N_3187,In_1261,In_1973);
nand U3188 (N_3188,In_2470,In_341);
and U3189 (N_3189,In_1991,In_894);
and U3190 (N_3190,In_149,In_1961);
xor U3191 (N_3191,In_1136,In_1170);
nand U3192 (N_3192,In_1640,In_940);
xnor U3193 (N_3193,In_1561,In_1127);
xnor U3194 (N_3194,In_698,In_2353);
xor U3195 (N_3195,In_978,In_1949);
and U3196 (N_3196,In_1692,In_1295);
or U3197 (N_3197,In_1951,In_587);
xor U3198 (N_3198,In_171,In_2345);
or U3199 (N_3199,In_1729,In_2324);
and U3200 (N_3200,In_1944,In_1719);
nand U3201 (N_3201,In_1963,In_1629);
and U3202 (N_3202,In_1640,In_1047);
and U3203 (N_3203,In_1492,In_2061);
xnor U3204 (N_3204,In_1665,In_1026);
nor U3205 (N_3205,In_87,In_1501);
nor U3206 (N_3206,In_1266,In_941);
nor U3207 (N_3207,In_2292,In_1754);
xnor U3208 (N_3208,In_1291,In_784);
or U3209 (N_3209,In_1176,In_2036);
nand U3210 (N_3210,In_111,In_1948);
xnor U3211 (N_3211,In_1080,In_971);
nand U3212 (N_3212,In_1301,In_1510);
xnor U3213 (N_3213,In_938,In_2404);
nor U3214 (N_3214,In_2380,In_1740);
nand U3215 (N_3215,In_818,In_803);
nand U3216 (N_3216,In_1294,In_1453);
xnor U3217 (N_3217,In_2405,In_84);
or U3218 (N_3218,In_114,In_1155);
nor U3219 (N_3219,In_800,In_1601);
nor U3220 (N_3220,In_1907,In_495);
and U3221 (N_3221,In_2198,In_31);
or U3222 (N_3222,In_2179,In_959);
nand U3223 (N_3223,In_1107,In_763);
xnor U3224 (N_3224,In_1953,In_418);
xor U3225 (N_3225,In_2196,In_1176);
nor U3226 (N_3226,In_1225,In_609);
xor U3227 (N_3227,In_1561,In_935);
and U3228 (N_3228,In_2277,In_381);
nor U3229 (N_3229,In_1942,In_74);
xor U3230 (N_3230,In_459,In_318);
nand U3231 (N_3231,In_1885,In_132);
nor U3232 (N_3232,In_463,In_336);
xor U3233 (N_3233,In_2212,In_0);
or U3234 (N_3234,In_1393,In_1752);
or U3235 (N_3235,In_2460,In_1098);
xnor U3236 (N_3236,In_1175,In_2430);
nor U3237 (N_3237,In_1524,In_702);
nor U3238 (N_3238,In_1746,In_1058);
xor U3239 (N_3239,In_1771,In_863);
xnor U3240 (N_3240,In_613,In_2295);
or U3241 (N_3241,In_1405,In_498);
nand U3242 (N_3242,In_180,In_1879);
xor U3243 (N_3243,In_205,In_1166);
nor U3244 (N_3244,In_2440,In_2313);
and U3245 (N_3245,In_1353,In_1496);
or U3246 (N_3246,In_627,In_133);
or U3247 (N_3247,In_1307,In_627);
xnor U3248 (N_3248,In_224,In_225);
xor U3249 (N_3249,In_1500,In_1905);
or U3250 (N_3250,In_2264,In_2222);
nor U3251 (N_3251,In_552,In_2154);
and U3252 (N_3252,In_1758,In_228);
nand U3253 (N_3253,In_224,In_272);
xor U3254 (N_3254,In_1379,In_79);
nor U3255 (N_3255,In_2216,In_83);
and U3256 (N_3256,In_338,In_896);
or U3257 (N_3257,In_2364,In_336);
xor U3258 (N_3258,In_2413,In_1731);
or U3259 (N_3259,In_1541,In_2328);
and U3260 (N_3260,In_2122,In_8);
nand U3261 (N_3261,In_1372,In_2320);
and U3262 (N_3262,In_1827,In_1076);
or U3263 (N_3263,In_1372,In_1381);
and U3264 (N_3264,In_2006,In_2099);
nand U3265 (N_3265,In_2342,In_597);
nand U3266 (N_3266,In_1492,In_506);
and U3267 (N_3267,In_1648,In_1764);
xnor U3268 (N_3268,In_1341,In_2262);
or U3269 (N_3269,In_208,In_1771);
nand U3270 (N_3270,In_1447,In_2192);
or U3271 (N_3271,In_1225,In_1118);
nor U3272 (N_3272,In_443,In_1535);
xor U3273 (N_3273,In_2170,In_1619);
nand U3274 (N_3274,In_2482,In_17);
nor U3275 (N_3275,In_616,In_480);
nor U3276 (N_3276,In_512,In_2271);
or U3277 (N_3277,In_830,In_1510);
or U3278 (N_3278,In_108,In_587);
or U3279 (N_3279,In_490,In_1221);
or U3280 (N_3280,In_1628,In_1023);
and U3281 (N_3281,In_1684,In_1381);
nor U3282 (N_3282,In_812,In_32);
nand U3283 (N_3283,In_1377,In_663);
and U3284 (N_3284,In_1497,In_1831);
nand U3285 (N_3285,In_1357,In_2200);
xor U3286 (N_3286,In_366,In_723);
nand U3287 (N_3287,In_1991,In_900);
and U3288 (N_3288,In_2381,In_2294);
nand U3289 (N_3289,In_2018,In_483);
or U3290 (N_3290,In_2432,In_1555);
xnor U3291 (N_3291,In_1191,In_2234);
and U3292 (N_3292,In_1673,In_1672);
or U3293 (N_3293,In_631,In_2351);
nor U3294 (N_3294,In_2194,In_465);
nor U3295 (N_3295,In_1902,In_1478);
and U3296 (N_3296,In_1755,In_331);
xnor U3297 (N_3297,In_1777,In_182);
and U3298 (N_3298,In_1960,In_2440);
nor U3299 (N_3299,In_1732,In_934);
xor U3300 (N_3300,In_1288,In_1350);
nor U3301 (N_3301,In_662,In_1232);
xor U3302 (N_3302,In_2016,In_1735);
xor U3303 (N_3303,In_284,In_142);
xor U3304 (N_3304,In_462,In_1131);
or U3305 (N_3305,In_16,In_1704);
nand U3306 (N_3306,In_2120,In_1873);
and U3307 (N_3307,In_204,In_42);
nor U3308 (N_3308,In_1938,In_215);
nand U3309 (N_3309,In_59,In_1946);
or U3310 (N_3310,In_814,In_2202);
nor U3311 (N_3311,In_2212,In_2059);
and U3312 (N_3312,In_64,In_197);
nand U3313 (N_3313,In_1654,In_1504);
and U3314 (N_3314,In_830,In_1322);
nand U3315 (N_3315,In_1912,In_2009);
and U3316 (N_3316,In_810,In_1757);
xor U3317 (N_3317,In_2160,In_1611);
nor U3318 (N_3318,In_308,In_1569);
nor U3319 (N_3319,In_1448,In_1287);
or U3320 (N_3320,In_280,In_1901);
nor U3321 (N_3321,In_1760,In_2297);
and U3322 (N_3322,In_556,In_1599);
or U3323 (N_3323,In_1602,In_1755);
xnor U3324 (N_3324,In_793,In_1183);
nand U3325 (N_3325,In_2340,In_183);
and U3326 (N_3326,In_49,In_1169);
or U3327 (N_3327,In_611,In_751);
xnor U3328 (N_3328,In_1249,In_971);
or U3329 (N_3329,In_229,In_184);
nor U3330 (N_3330,In_259,In_1173);
xnor U3331 (N_3331,In_1815,In_1297);
nand U3332 (N_3332,In_298,In_1308);
nor U3333 (N_3333,In_74,In_2338);
and U3334 (N_3334,In_622,In_2202);
and U3335 (N_3335,In_711,In_2084);
nor U3336 (N_3336,In_2444,In_2210);
and U3337 (N_3337,In_1345,In_1274);
xor U3338 (N_3338,In_2160,In_1415);
and U3339 (N_3339,In_2338,In_2187);
xnor U3340 (N_3340,In_1578,In_1205);
nand U3341 (N_3341,In_1786,In_906);
and U3342 (N_3342,In_2442,In_674);
and U3343 (N_3343,In_2424,In_1052);
nor U3344 (N_3344,In_698,In_469);
nor U3345 (N_3345,In_2486,In_1535);
nor U3346 (N_3346,In_1543,In_307);
nand U3347 (N_3347,In_980,In_2143);
nor U3348 (N_3348,In_8,In_67);
nor U3349 (N_3349,In_59,In_458);
nand U3350 (N_3350,In_2043,In_1145);
xnor U3351 (N_3351,In_290,In_574);
or U3352 (N_3352,In_1963,In_994);
and U3353 (N_3353,In_25,In_1153);
and U3354 (N_3354,In_2441,In_1776);
nand U3355 (N_3355,In_544,In_1075);
nand U3356 (N_3356,In_306,In_1039);
nor U3357 (N_3357,In_258,In_2398);
nor U3358 (N_3358,In_1424,In_1508);
or U3359 (N_3359,In_123,In_1973);
xor U3360 (N_3360,In_777,In_1037);
xnor U3361 (N_3361,In_1525,In_913);
nor U3362 (N_3362,In_1751,In_2380);
and U3363 (N_3363,In_1424,In_551);
nor U3364 (N_3364,In_228,In_2280);
xnor U3365 (N_3365,In_1697,In_2042);
xnor U3366 (N_3366,In_331,In_1651);
and U3367 (N_3367,In_43,In_823);
and U3368 (N_3368,In_797,In_2102);
nand U3369 (N_3369,In_413,In_717);
and U3370 (N_3370,In_2423,In_2106);
nand U3371 (N_3371,In_171,In_1468);
and U3372 (N_3372,In_1453,In_1039);
xnor U3373 (N_3373,In_456,In_139);
or U3374 (N_3374,In_1816,In_1561);
nand U3375 (N_3375,In_2079,In_2151);
or U3376 (N_3376,In_2053,In_197);
nor U3377 (N_3377,In_763,In_2317);
nor U3378 (N_3378,In_2457,In_1618);
and U3379 (N_3379,In_1090,In_1493);
or U3380 (N_3380,In_2474,In_785);
nand U3381 (N_3381,In_517,In_2373);
and U3382 (N_3382,In_1581,In_435);
nor U3383 (N_3383,In_2186,In_934);
or U3384 (N_3384,In_1490,In_1277);
or U3385 (N_3385,In_820,In_1291);
and U3386 (N_3386,In_966,In_1836);
nand U3387 (N_3387,In_895,In_1144);
or U3388 (N_3388,In_812,In_1705);
nand U3389 (N_3389,In_28,In_2243);
xnor U3390 (N_3390,In_1051,In_311);
nand U3391 (N_3391,In_1946,In_1705);
nand U3392 (N_3392,In_1690,In_1038);
or U3393 (N_3393,In_2452,In_1140);
nor U3394 (N_3394,In_2093,In_989);
xor U3395 (N_3395,In_131,In_47);
xor U3396 (N_3396,In_2065,In_2181);
nor U3397 (N_3397,In_899,In_2267);
nor U3398 (N_3398,In_1629,In_2211);
and U3399 (N_3399,In_200,In_2217);
nor U3400 (N_3400,In_2315,In_1911);
nor U3401 (N_3401,In_2332,In_1139);
nor U3402 (N_3402,In_1746,In_1640);
xnor U3403 (N_3403,In_1159,In_769);
xnor U3404 (N_3404,In_2327,In_569);
nor U3405 (N_3405,In_1394,In_1853);
nand U3406 (N_3406,In_1398,In_1525);
nor U3407 (N_3407,In_1331,In_2251);
and U3408 (N_3408,In_1085,In_1547);
xnor U3409 (N_3409,In_40,In_309);
nand U3410 (N_3410,In_813,In_21);
nand U3411 (N_3411,In_2022,In_1219);
nor U3412 (N_3412,In_1686,In_341);
or U3413 (N_3413,In_258,In_218);
nand U3414 (N_3414,In_1355,In_1116);
nand U3415 (N_3415,In_1038,In_1056);
or U3416 (N_3416,In_1541,In_2061);
or U3417 (N_3417,In_494,In_1951);
nor U3418 (N_3418,In_1874,In_1639);
nor U3419 (N_3419,In_2190,In_2123);
nor U3420 (N_3420,In_1188,In_2310);
or U3421 (N_3421,In_200,In_2238);
nand U3422 (N_3422,In_93,In_1979);
nor U3423 (N_3423,In_844,In_787);
or U3424 (N_3424,In_2171,In_12);
nand U3425 (N_3425,In_329,In_1330);
and U3426 (N_3426,In_54,In_2307);
nand U3427 (N_3427,In_739,In_282);
nand U3428 (N_3428,In_1941,In_214);
nand U3429 (N_3429,In_2055,In_1731);
or U3430 (N_3430,In_878,In_1562);
nor U3431 (N_3431,In_1754,In_154);
nor U3432 (N_3432,In_326,In_1390);
and U3433 (N_3433,In_2087,In_872);
or U3434 (N_3434,In_116,In_527);
or U3435 (N_3435,In_1330,In_1229);
xor U3436 (N_3436,In_1276,In_2354);
or U3437 (N_3437,In_589,In_2458);
xor U3438 (N_3438,In_1707,In_646);
xnor U3439 (N_3439,In_1996,In_202);
and U3440 (N_3440,In_1318,In_405);
or U3441 (N_3441,In_2349,In_2430);
or U3442 (N_3442,In_1354,In_1954);
xor U3443 (N_3443,In_787,In_432);
and U3444 (N_3444,In_1488,In_432);
or U3445 (N_3445,In_492,In_2015);
or U3446 (N_3446,In_488,In_2303);
nand U3447 (N_3447,In_49,In_2225);
and U3448 (N_3448,In_1252,In_725);
and U3449 (N_3449,In_1380,In_411);
xor U3450 (N_3450,In_985,In_596);
nor U3451 (N_3451,In_92,In_1681);
or U3452 (N_3452,In_762,In_2403);
and U3453 (N_3453,In_1506,In_195);
xor U3454 (N_3454,In_2269,In_990);
nand U3455 (N_3455,In_618,In_745);
and U3456 (N_3456,In_2441,In_1418);
and U3457 (N_3457,In_1423,In_748);
nor U3458 (N_3458,In_2231,In_2084);
and U3459 (N_3459,In_2331,In_1606);
nand U3460 (N_3460,In_31,In_39);
nand U3461 (N_3461,In_75,In_2002);
or U3462 (N_3462,In_2356,In_326);
nor U3463 (N_3463,In_375,In_1090);
or U3464 (N_3464,In_2108,In_599);
and U3465 (N_3465,In_440,In_1425);
or U3466 (N_3466,In_1686,In_2402);
nor U3467 (N_3467,In_1182,In_102);
nand U3468 (N_3468,In_2170,In_1218);
and U3469 (N_3469,In_1854,In_839);
xor U3470 (N_3470,In_221,In_420);
and U3471 (N_3471,In_2108,In_593);
nor U3472 (N_3472,In_1640,In_2040);
nand U3473 (N_3473,In_1503,In_923);
and U3474 (N_3474,In_1078,In_2025);
nor U3475 (N_3475,In_1522,In_183);
xnor U3476 (N_3476,In_1789,In_546);
or U3477 (N_3477,In_1572,In_774);
nand U3478 (N_3478,In_1277,In_1609);
nor U3479 (N_3479,In_592,In_1933);
nand U3480 (N_3480,In_399,In_471);
nor U3481 (N_3481,In_1362,In_278);
or U3482 (N_3482,In_309,In_1414);
nand U3483 (N_3483,In_1160,In_143);
or U3484 (N_3484,In_1193,In_2455);
and U3485 (N_3485,In_2331,In_1831);
and U3486 (N_3486,In_1352,In_1064);
xnor U3487 (N_3487,In_621,In_1015);
nor U3488 (N_3488,In_1665,In_7);
or U3489 (N_3489,In_1018,In_241);
xor U3490 (N_3490,In_1017,In_2070);
or U3491 (N_3491,In_561,In_553);
nor U3492 (N_3492,In_1866,In_1305);
nand U3493 (N_3493,In_2224,In_1012);
and U3494 (N_3494,In_1799,In_2272);
nor U3495 (N_3495,In_1132,In_1363);
nand U3496 (N_3496,In_581,In_747);
nand U3497 (N_3497,In_628,In_203);
nand U3498 (N_3498,In_1408,In_2468);
nand U3499 (N_3499,In_1006,In_1582);
or U3500 (N_3500,In_1979,In_202);
or U3501 (N_3501,In_2060,In_518);
or U3502 (N_3502,In_483,In_705);
nor U3503 (N_3503,In_769,In_320);
nand U3504 (N_3504,In_732,In_216);
xor U3505 (N_3505,In_627,In_62);
or U3506 (N_3506,In_802,In_1326);
and U3507 (N_3507,In_1852,In_2301);
nand U3508 (N_3508,In_1162,In_2056);
and U3509 (N_3509,In_2142,In_2362);
and U3510 (N_3510,In_2036,In_1073);
nand U3511 (N_3511,In_42,In_936);
nor U3512 (N_3512,In_544,In_2195);
or U3513 (N_3513,In_2021,In_2227);
or U3514 (N_3514,In_1307,In_136);
xor U3515 (N_3515,In_1213,In_1792);
xnor U3516 (N_3516,In_2030,In_1858);
xnor U3517 (N_3517,In_1848,In_105);
nor U3518 (N_3518,In_1021,In_198);
or U3519 (N_3519,In_1039,In_1949);
and U3520 (N_3520,In_1751,In_1543);
or U3521 (N_3521,In_1209,In_370);
nor U3522 (N_3522,In_574,In_986);
or U3523 (N_3523,In_2395,In_1520);
nor U3524 (N_3524,In_85,In_1747);
nor U3525 (N_3525,In_1664,In_1485);
nor U3526 (N_3526,In_1707,In_1241);
nor U3527 (N_3527,In_710,In_1747);
xnor U3528 (N_3528,In_637,In_1799);
and U3529 (N_3529,In_1453,In_1956);
nand U3530 (N_3530,In_2297,In_2098);
xnor U3531 (N_3531,In_1993,In_2182);
nor U3532 (N_3532,In_2047,In_2101);
and U3533 (N_3533,In_1255,In_1100);
nor U3534 (N_3534,In_502,In_791);
and U3535 (N_3535,In_1096,In_567);
nand U3536 (N_3536,In_2482,In_2334);
xnor U3537 (N_3537,In_1843,In_1481);
nand U3538 (N_3538,In_1157,In_568);
nor U3539 (N_3539,In_1159,In_1351);
nand U3540 (N_3540,In_1894,In_517);
nor U3541 (N_3541,In_2326,In_24);
xor U3542 (N_3542,In_2045,In_1177);
and U3543 (N_3543,In_203,In_2440);
xnor U3544 (N_3544,In_2090,In_1892);
xnor U3545 (N_3545,In_271,In_2079);
and U3546 (N_3546,In_1810,In_1294);
nor U3547 (N_3547,In_1586,In_157);
and U3548 (N_3548,In_1093,In_316);
or U3549 (N_3549,In_560,In_278);
xnor U3550 (N_3550,In_207,In_1158);
nor U3551 (N_3551,In_1373,In_1881);
nor U3552 (N_3552,In_92,In_2271);
or U3553 (N_3553,In_1967,In_470);
or U3554 (N_3554,In_1189,In_1885);
xor U3555 (N_3555,In_257,In_2196);
xnor U3556 (N_3556,In_574,In_1456);
nand U3557 (N_3557,In_1515,In_2118);
nand U3558 (N_3558,In_1013,In_707);
and U3559 (N_3559,In_1552,In_24);
nand U3560 (N_3560,In_610,In_864);
or U3561 (N_3561,In_2401,In_1491);
nand U3562 (N_3562,In_93,In_978);
nand U3563 (N_3563,In_2470,In_286);
and U3564 (N_3564,In_1247,In_1566);
xor U3565 (N_3565,In_1833,In_226);
xnor U3566 (N_3566,In_1789,In_1674);
and U3567 (N_3567,In_578,In_1243);
nand U3568 (N_3568,In_724,In_939);
or U3569 (N_3569,In_1231,In_386);
nor U3570 (N_3570,In_666,In_1658);
nand U3571 (N_3571,In_172,In_1657);
or U3572 (N_3572,In_34,In_2233);
and U3573 (N_3573,In_2005,In_136);
nand U3574 (N_3574,In_221,In_1940);
and U3575 (N_3575,In_261,In_1662);
and U3576 (N_3576,In_1759,In_689);
and U3577 (N_3577,In_2038,In_855);
nor U3578 (N_3578,In_2042,In_1149);
or U3579 (N_3579,In_1214,In_267);
nor U3580 (N_3580,In_1999,In_950);
nand U3581 (N_3581,In_1564,In_746);
or U3582 (N_3582,In_2035,In_2103);
nand U3583 (N_3583,In_746,In_2149);
or U3584 (N_3584,In_1236,In_1610);
xor U3585 (N_3585,In_255,In_1258);
nor U3586 (N_3586,In_1607,In_2367);
or U3587 (N_3587,In_1722,In_843);
nor U3588 (N_3588,In_1225,In_2133);
nor U3589 (N_3589,In_2262,In_1839);
and U3590 (N_3590,In_2413,In_1015);
nand U3591 (N_3591,In_2358,In_1068);
or U3592 (N_3592,In_1540,In_604);
and U3593 (N_3593,In_518,In_866);
xnor U3594 (N_3594,In_1738,In_2318);
or U3595 (N_3595,In_1487,In_1681);
and U3596 (N_3596,In_1561,In_831);
nor U3597 (N_3597,In_312,In_2277);
nor U3598 (N_3598,In_2408,In_1304);
and U3599 (N_3599,In_1258,In_1359);
xnor U3600 (N_3600,In_1437,In_622);
nor U3601 (N_3601,In_167,In_2013);
nand U3602 (N_3602,In_983,In_1650);
and U3603 (N_3603,In_2075,In_1617);
xor U3604 (N_3604,In_1072,In_1140);
or U3605 (N_3605,In_1151,In_946);
nand U3606 (N_3606,In_1725,In_1895);
nand U3607 (N_3607,In_2136,In_23);
nor U3608 (N_3608,In_2029,In_895);
or U3609 (N_3609,In_338,In_1143);
xor U3610 (N_3610,In_916,In_1062);
or U3611 (N_3611,In_1714,In_39);
nand U3612 (N_3612,In_1304,In_971);
and U3613 (N_3613,In_1423,In_1997);
nand U3614 (N_3614,In_776,In_766);
nand U3615 (N_3615,In_447,In_254);
nor U3616 (N_3616,In_1445,In_2333);
nor U3617 (N_3617,In_707,In_1908);
xnor U3618 (N_3618,In_806,In_496);
or U3619 (N_3619,In_482,In_885);
nand U3620 (N_3620,In_1050,In_831);
or U3621 (N_3621,In_1055,In_340);
nand U3622 (N_3622,In_2054,In_1571);
or U3623 (N_3623,In_2232,In_1745);
nor U3624 (N_3624,In_460,In_979);
or U3625 (N_3625,In_2049,In_1338);
nor U3626 (N_3626,In_1065,In_690);
xor U3627 (N_3627,In_1060,In_1985);
and U3628 (N_3628,In_1814,In_166);
or U3629 (N_3629,In_1245,In_1645);
xor U3630 (N_3630,In_2396,In_1328);
nor U3631 (N_3631,In_417,In_2293);
or U3632 (N_3632,In_1552,In_249);
nand U3633 (N_3633,In_498,In_1112);
nand U3634 (N_3634,In_2478,In_199);
xnor U3635 (N_3635,In_2040,In_685);
nand U3636 (N_3636,In_1037,In_2407);
nand U3637 (N_3637,In_1203,In_1385);
and U3638 (N_3638,In_58,In_983);
xnor U3639 (N_3639,In_606,In_739);
nand U3640 (N_3640,In_2469,In_960);
xor U3641 (N_3641,In_2110,In_1538);
and U3642 (N_3642,In_1971,In_251);
xor U3643 (N_3643,In_1122,In_388);
or U3644 (N_3644,In_246,In_1429);
or U3645 (N_3645,In_1818,In_297);
and U3646 (N_3646,In_1369,In_2402);
xnor U3647 (N_3647,In_1256,In_132);
nor U3648 (N_3648,In_338,In_2240);
xnor U3649 (N_3649,In_1194,In_565);
nand U3650 (N_3650,In_1945,In_579);
or U3651 (N_3651,In_247,In_1650);
or U3652 (N_3652,In_1436,In_1595);
or U3653 (N_3653,In_1084,In_806);
or U3654 (N_3654,In_1230,In_1804);
nor U3655 (N_3655,In_2367,In_1031);
nand U3656 (N_3656,In_2065,In_900);
and U3657 (N_3657,In_2115,In_1114);
or U3658 (N_3658,In_1249,In_1349);
and U3659 (N_3659,In_2256,In_394);
nor U3660 (N_3660,In_1755,In_1077);
or U3661 (N_3661,In_2484,In_334);
xnor U3662 (N_3662,In_388,In_320);
xnor U3663 (N_3663,In_1072,In_1689);
or U3664 (N_3664,In_174,In_2462);
nand U3665 (N_3665,In_305,In_2230);
or U3666 (N_3666,In_315,In_1432);
nor U3667 (N_3667,In_343,In_1176);
xnor U3668 (N_3668,In_1098,In_1040);
xnor U3669 (N_3669,In_79,In_606);
nor U3670 (N_3670,In_1158,In_698);
xnor U3671 (N_3671,In_173,In_1777);
nor U3672 (N_3672,In_551,In_932);
nor U3673 (N_3673,In_865,In_868);
nor U3674 (N_3674,In_111,In_1567);
xor U3675 (N_3675,In_1944,In_195);
or U3676 (N_3676,In_623,In_2227);
nor U3677 (N_3677,In_1029,In_1435);
and U3678 (N_3678,In_2205,In_2433);
nor U3679 (N_3679,In_157,In_1442);
or U3680 (N_3680,In_886,In_954);
nand U3681 (N_3681,In_211,In_635);
and U3682 (N_3682,In_221,In_817);
xor U3683 (N_3683,In_48,In_1835);
nor U3684 (N_3684,In_389,In_1623);
xor U3685 (N_3685,In_1939,In_828);
and U3686 (N_3686,In_2214,In_1166);
xor U3687 (N_3687,In_58,In_550);
nor U3688 (N_3688,In_2416,In_197);
or U3689 (N_3689,In_1168,In_600);
nand U3690 (N_3690,In_974,In_189);
nor U3691 (N_3691,In_107,In_2118);
nand U3692 (N_3692,In_371,In_1923);
nand U3693 (N_3693,In_1161,In_2050);
and U3694 (N_3694,In_1046,In_1650);
nor U3695 (N_3695,In_1012,In_2096);
nand U3696 (N_3696,In_148,In_1613);
and U3697 (N_3697,In_2396,In_2324);
xor U3698 (N_3698,In_2055,In_1646);
xor U3699 (N_3699,In_593,In_1370);
nor U3700 (N_3700,In_1690,In_2350);
or U3701 (N_3701,In_321,In_1758);
nor U3702 (N_3702,In_2465,In_528);
nand U3703 (N_3703,In_1097,In_72);
or U3704 (N_3704,In_882,In_2142);
nand U3705 (N_3705,In_578,In_1146);
and U3706 (N_3706,In_318,In_2006);
nand U3707 (N_3707,In_966,In_1200);
or U3708 (N_3708,In_1207,In_296);
xor U3709 (N_3709,In_1047,In_1986);
xnor U3710 (N_3710,In_1827,In_1268);
nor U3711 (N_3711,In_613,In_204);
and U3712 (N_3712,In_2423,In_1173);
and U3713 (N_3713,In_88,In_1890);
and U3714 (N_3714,In_1020,In_1051);
nand U3715 (N_3715,In_2241,In_2351);
xor U3716 (N_3716,In_1479,In_1016);
nor U3717 (N_3717,In_2119,In_223);
or U3718 (N_3718,In_2479,In_186);
nor U3719 (N_3719,In_2154,In_387);
nor U3720 (N_3720,In_842,In_980);
xnor U3721 (N_3721,In_2466,In_829);
nand U3722 (N_3722,In_1380,In_1861);
or U3723 (N_3723,In_1183,In_1560);
nand U3724 (N_3724,In_261,In_1697);
or U3725 (N_3725,In_1670,In_596);
nand U3726 (N_3726,In_288,In_1157);
nor U3727 (N_3727,In_1457,In_801);
or U3728 (N_3728,In_22,In_2287);
nand U3729 (N_3729,In_2474,In_2273);
nor U3730 (N_3730,In_1433,In_206);
xor U3731 (N_3731,In_2242,In_1578);
xnor U3732 (N_3732,In_1098,In_1607);
or U3733 (N_3733,In_1436,In_2480);
nand U3734 (N_3734,In_428,In_805);
and U3735 (N_3735,In_1529,In_459);
and U3736 (N_3736,In_1582,In_1467);
nor U3737 (N_3737,In_723,In_1537);
nand U3738 (N_3738,In_1853,In_1867);
nand U3739 (N_3739,In_35,In_1337);
and U3740 (N_3740,In_2438,In_2188);
and U3741 (N_3741,In_1347,In_1410);
and U3742 (N_3742,In_1543,In_1777);
nand U3743 (N_3743,In_264,In_1329);
and U3744 (N_3744,In_1039,In_739);
xor U3745 (N_3745,In_2199,In_1189);
nor U3746 (N_3746,In_1192,In_11);
nor U3747 (N_3747,In_1094,In_2251);
nand U3748 (N_3748,In_958,In_610);
and U3749 (N_3749,In_1873,In_1690);
and U3750 (N_3750,In_2242,In_2128);
or U3751 (N_3751,In_1711,In_1198);
and U3752 (N_3752,In_2284,In_1154);
or U3753 (N_3753,In_550,In_2174);
and U3754 (N_3754,In_163,In_361);
nor U3755 (N_3755,In_2211,In_108);
xnor U3756 (N_3756,In_691,In_398);
nor U3757 (N_3757,In_911,In_2254);
and U3758 (N_3758,In_2418,In_20);
or U3759 (N_3759,In_2136,In_2075);
nand U3760 (N_3760,In_2243,In_1960);
and U3761 (N_3761,In_1083,In_2386);
xnor U3762 (N_3762,In_1861,In_1770);
xnor U3763 (N_3763,In_332,In_697);
nand U3764 (N_3764,In_818,In_1513);
or U3765 (N_3765,In_1306,In_2254);
and U3766 (N_3766,In_519,In_1653);
and U3767 (N_3767,In_685,In_2284);
xnor U3768 (N_3768,In_2464,In_2240);
or U3769 (N_3769,In_1858,In_2165);
xor U3770 (N_3770,In_1596,In_1361);
xor U3771 (N_3771,In_1643,In_1806);
nor U3772 (N_3772,In_1511,In_2258);
or U3773 (N_3773,In_473,In_1471);
nand U3774 (N_3774,In_2180,In_1572);
nor U3775 (N_3775,In_194,In_2095);
or U3776 (N_3776,In_1203,In_78);
and U3777 (N_3777,In_513,In_2076);
nand U3778 (N_3778,In_1939,In_667);
nor U3779 (N_3779,In_1824,In_1745);
or U3780 (N_3780,In_1495,In_872);
nand U3781 (N_3781,In_2278,In_1637);
nor U3782 (N_3782,In_1503,In_1785);
xor U3783 (N_3783,In_2160,In_567);
nand U3784 (N_3784,In_2453,In_1169);
nor U3785 (N_3785,In_263,In_1129);
nor U3786 (N_3786,In_887,In_2102);
nor U3787 (N_3787,In_415,In_2314);
xnor U3788 (N_3788,In_2305,In_55);
nand U3789 (N_3789,In_2475,In_1702);
nor U3790 (N_3790,In_1246,In_1597);
xnor U3791 (N_3791,In_2277,In_1188);
and U3792 (N_3792,In_1773,In_1742);
or U3793 (N_3793,In_2144,In_2227);
nand U3794 (N_3794,In_1298,In_325);
nor U3795 (N_3795,In_722,In_2405);
xnor U3796 (N_3796,In_2300,In_1703);
and U3797 (N_3797,In_1747,In_1862);
nor U3798 (N_3798,In_1335,In_64);
or U3799 (N_3799,In_1723,In_258);
xor U3800 (N_3800,In_865,In_2375);
xor U3801 (N_3801,In_610,In_1606);
xor U3802 (N_3802,In_766,In_1212);
xor U3803 (N_3803,In_197,In_723);
and U3804 (N_3804,In_1713,In_1697);
and U3805 (N_3805,In_1405,In_2376);
nor U3806 (N_3806,In_391,In_837);
nor U3807 (N_3807,In_1557,In_48);
nand U3808 (N_3808,In_1901,In_2328);
and U3809 (N_3809,In_904,In_1340);
nand U3810 (N_3810,In_317,In_970);
xnor U3811 (N_3811,In_2249,In_264);
nand U3812 (N_3812,In_937,In_1865);
xnor U3813 (N_3813,In_2388,In_1151);
nor U3814 (N_3814,In_2399,In_1811);
nand U3815 (N_3815,In_1808,In_578);
nor U3816 (N_3816,In_480,In_1039);
nor U3817 (N_3817,In_1347,In_1808);
nor U3818 (N_3818,In_717,In_724);
xnor U3819 (N_3819,In_423,In_311);
nand U3820 (N_3820,In_960,In_390);
nor U3821 (N_3821,In_2334,In_508);
nand U3822 (N_3822,In_86,In_2346);
nor U3823 (N_3823,In_848,In_970);
xnor U3824 (N_3824,In_726,In_1672);
xor U3825 (N_3825,In_1664,In_305);
and U3826 (N_3826,In_714,In_334);
nor U3827 (N_3827,In_736,In_725);
nor U3828 (N_3828,In_1426,In_1457);
xnor U3829 (N_3829,In_1586,In_547);
nand U3830 (N_3830,In_2275,In_367);
nor U3831 (N_3831,In_111,In_658);
xor U3832 (N_3832,In_885,In_1767);
xnor U3833 (N_3833,In_461,In_2463);
and U3834 (N_3834,In_350,In_1162);
nor U3835 (N_3835,In_1015,In_650);
or U3836 (N_3836,In_1679,In_1212);
nor U3837 (N_3837,In_1594,In_1112);
and U3838 (N_3838,In_2290,In_2005);
xor U3839 (N_3839,In_1915,In_860);
nand U3840 (N_3840,In_1503,In_850);
nor U3841 (N_3841,In_862,In_39);
or U3842 (N_3842,In_2222,In_1401);
or U3843 (N_3843,In_365,In_1520);
xnor U3844 (N_3844,In_1590,In_2169);
xor U3845 (N_3845,In_1168,In_1174);
and U3846 (N_3846,In_1478,In_2161);
or U3847 (N_3847,In_1884,In_434);
nand U3848 (N_3848,In_868,In_234);
and U3849 (N_3849,In_720,In_2116);
xnor U3850 (N_3850,In_1756,In_2237);
or U3851 (N_3851,In_967,In_639);
xnor U3852 (N_3852,In_1281,In_194);
nand U3853 (N_3853,In_302,In_348);
and U3854 (N_3854,In_2229,In_2134);
xnor U3855 (N_3855,In_543,In_1434);
and U3856 (N_3856,In_2069,In_1878);
nand U3857 (N_3857,In_2232,In_802);
nor U3858 (N_3858,In_1657,In_1817);
and U3859 (N_3859,In_2226,In_1981);
xor U3860 (N_3860,In_825,In_985);
nand U3861 (N_3861,In_1761,In_1488);
nor U3862 (N_3862,In_2241,In_1232);
nor U3863 (N_3863,In_1239,In_1275);
or U3864 (N_3864,In_821,In_709);
nand U3865 (N_3865,In_509,In_1925);
or U3866 (N_3866,In_828,In_17);
and U3867 (N_3867,In_2369,In_1548);
xor U3868 (N_3868,In_1344,In_2425);
or U3869 (N_3869,In_1393,In_1758);
xor U3870 (N_3870,In_840,In_995);
or U3871 (N_3871,In_2040,In_1951);
or U3872 (N_3872,In_1726,In_39);
xor U3873 (N_3873,In_1326,In_317);
nor U3874 (N_3874,In_2028,In_2457);
and U3875 (N_3875,In_1585,In_1960);
and U3876 (N_3876,In_1286,In_1276);
and U3877 (N_3877,In_2199,In_1902);
xor U3878 (N_3878,In_107,In_1136);
nor U3879 (N_3879,In_932,In_425);
xor U3880 (N_3880,In_71,In_1090);
nand U3881 (N_3881,In_631,In_1646);
and U3882 (N_3882,In_2034,In_1673);
xor U3883 (N_3883,In_1182,In_446);
and U3884 (N_3884,In_1629,In_1550);
and U3885 (N_3885,In_2143,In_2075);
xor U3886 (N_3886,In_2223,In_2069);
and U3887 (N_3887,In_1889,In_1933);
xor U3888 (N_3888,In_2257,In_930);
and U3889 (N_3889,In_472,In_707);
and U3890 (N_3890,In_2459,In_1435);
nor U3891 (N_3891,In_1782,In_1622);
nor U3892 (N_3892,In_2278,In_1482);
nand U3893 (N_3893,In_1142,In_1003);
or U3894 (N_3894,In_473,In_205);
or U3895 (N_3895,In_445,In_1219);
or U3896 (N_3896,In_1338,In_658);
nor U3897 (N_3897,In_512,In_1066);
nor U3898 (N_3898,In_471,In_1284);
and U3899 (N_3899,In_1386,In_1919);
xnor U3900 (N_3900,In_976,In_1266);
nor U3901 (N_3901,In_1179,In_2407);
xor U3902 (N_3902,In_1561,In_2158);
nand U3903 (N_3903,In_1026,In_635);
xnor U3904 (N_3904,In_2111,In_1619);
xor U3905 (N_3905,In_1294,In_356);
nand U3906 (N_3906,In_1551,In_1426);
nor U3907 (N_3907,In_918,In_48);
nand U3908 (N_3908,In_2148,In_649);
nor U3909 (N_3909,In_1078,In_1873);
nand U3910 (N_3910,In_2138,In_1760);
and U3911 (N_3911,In_1165,In_642);
nor U3912 (N_3912,In_1341,In_421);
and U3913 (N_3913,In_452,In_2118);
or U3914 (N_3914,In_912,In_547);
xnor U3915 (N_3915,In_1700,In_2135);
xor U3916 (N_3916,In_1878,In_443);
nor U3917 (N_3917,In_1937,In_2278);
and U3918 (N_3918,In_302,In_77);
xor U3919 (N_3919,In_1077,In_1790);
xnor U3920 (N_3920,In_271,In_2474);
nand U3921 (N_3921,In_1101,In_1106);
nand U3922 (N_3922,In_312,In_1667);
nand U3923 (N_3923,In_1886,In_1021);
nand U3924 (N_3924,In_930,In_2204);
or U3925 (N_3925,In_2273,In_2352);
nand U3926 (N_3926,In_1072,In_1569);
xnor U3927 (N_3927,In_982,In_414);
or U3928 (N_3928,In_2135,In_1979);
nor U3929 (N_3929,In_1456,In_942);
xor U3930 (N_3930,In_1305,In_1678);
and U3931 (N_3931,In_1565,In_1430);
nor U3932 (N_3932,In_1100,In_2330);
nand U3933 (N_3933,In_1328,In_2294);
nor U3934 (N_3934,In_2346,In_927);
nor U3935 (N_3935,In_1068,In_1522);
nand U3936 (N_3936,In_2376,In_2093);
and U3937 (N_3937,In_578,In_2403);
xnor U3938 (N_3938,In_2135,In_2030);
xnor U3939 (N_3939,In_1492,In_1834);
or U3940 (N_3940,In_789,In_1896);
nor U3941 (N_3941,In_1623,In_742);
and U3942 (N_3942,In_29,In_2297);
xor U3943 (N_3943,In_1269,In_2149);
or U3944 (N_3944,In_912,In_1264);
or U3945 (N_3945,In_1233,In_2340);
nor U3946 (N_3946,In_288,In_2365);
nor U3947 (N_3947,In_1518,In_1844);
xor U3948 (N_3948,In_594,In_957);
xor U3949 (N_3949,In_557,In_1575);
nor U3950 (N_3950,In_2054,In_1907);
nor U3951 (N_3951,In_610,In_2213);
xnor U3952 (N_3952,In_1250,In_410);
nor U3953 (N_3953,In_187,In_1365);
and U3954 (N_3954,In_2217,In_679);
xnor U3955 (N_3955,In_904,In_2429);
or U3956 (N_3956,In_2092,In_2232);
or U3957 (N_3957,In_2308,In_1323);
nor U3958 (N_3958,In_325,In_1636);
nor U3959 (N_3959,In_1496,In_816);
xnor U3960 (N_3960,In_528,In_2143);
xor U3961 (N_3961,In_2397,In_102);
or U3962 (N_3962,In_1623,In_291);
and U3963 (N_3963,In_1632,In_820);
nor U3964 (N_3964,In_879,In_1412);
xnor U3965 (N_3965,In_3,In_377);
and U3966 (N_3966,In_864,In_842);
xnor U3967 (N_3967,In_1555,In_1681);
and U3968 (N_3968,In_827,In_722);
or U3969 (N_3969,In_310,In_1842);
nor U3970 (N_3970,In_151,In_879);
nand U3971 (N_3971,In_284,In_644);
nor U3972 (N_3972,In_282,In_1585);
nand U3973 (N_3973,In_1567,In_225);
nand U3974 (N_3974,In_2387,In_1160);
and U3975 (N_3975,In_2430,In_1347);
xor U3976 (N_3976,In_2446,In_1170);
xnor U3977 (N_3977,In_2452,In_331);
nor U3978 (N_3978,In_2388,In_1393);
and U3979 (N_3979,In_1430,In_1119);
or U3980 (N_3980,In_711,In_1826);
and U3981 (N_3981,In_945,In_2098);
or U3982 (N_3982,In_1190,In_939);
nor U3983 (N_3983,In_529,In_45);
or U3984 (N_3984,In_1180,In_1208);
nor U3985 (N_3985,In_903,In_523);
and U3986 (N_3986,In_37,In_2453);
nand U3987 (N_3987,In_2208,In_1232);
xor U3988 (N_3988,In_2441,In_1773);
nand U3989 (N_3989,In_497,In_2249);
nor U3990 (N_3990,In_1668,In_1291);
nand U3991 (N_3991,In_2081,In_1913);
nand U3992 (N_3992,In_883,In_266);
and U3993 (N_3993,In_2368,In_113);
xor U3994 (N_3994,In_498,In_2467);
and U3995 (N_3995,In_251,In_1587);
and U3996 (N_3996,In_949,In_898);
nand U3997 (N_3997,In_1792,In_1557);
nand U3998 (N_3998,In_318,In_693);
nor U3999 (N_3999,In_1930,In_1660);
or U4000 (N_4000,In_1289,In_1313);
nand U4001 (N_4001,In_777,In_1378);
nor U4002 (N_4002,In_1604,In_111);
nand U4003 (N_4003,In_1300,In_434);
xnor U4004 (N_4004,In_1158,In_960);
and U4005 (N_4005,In_796,In_1652);
nand U4006 (N_4006,In_444,In_830);
nand U4007 (N_4007,In_1319,In_1474);
nand U4008 (N_4008,In_1245,In_88);
xnor U4009 (N_4009,In_1200,In_517);
or U4010 (N_4010,In_1964,In_1582);
or U4011 (N_4011,In_923,In_860);
nand U4012 (N_4012,In_825,In_1531);
xnor U4013 (N_4013,In_1575,In_1490);
nor U4014 (N_4014,In_668,In_912);
and U4015 (N_4015,In_1962,In_1915);
nand U4016 (N_4016,In_258,In_1748);
or U4017 (N_4017,In_228,In_211);
xor U4018 (N_4018,In_2333,In_1650);
and U4019 (N_4019,In_2299,In_2162);
xnor U4020 (N_4020,In_395,In_2072);
nand U4021 (N_4021,In_1879,In_755);
and U4022 (N_4022,In_1022,In_1692);
nand U4023 (N_4023,In_1946,In_474);
and U4024 (N_4024,In_2367,In_2116);
nor U4025 (N_4025,In_1336,In_1792);
nor U4026 (N_4026,In_896,In_1515);
xnor U4027 (N_4027,In_1856,In_1657);
nor U4028 (N_4028,In_194,In_1099);
nor U4029 (N_4029,In_2096,In_548);
or U4030 (N_4030,In_222,In_2345);
or U4031 (N_4031,In_2422,In_213);
or U4032 (N_4032,In_261,In_2186);
or U4033 (N_4033,In_1314,In_103);
xor U4034 (N_4034,In_1385,In_1499);
or U4035 (N_4035,In_1528,In_1892);
xor U4036 (N_4036,In_360,In_905);
xor U4037 (N_4037,In_2169,In_1488);
xor U4038 (N_4038,In_2131,In_1445);
and U4039 (N_4039,In_1679,In_1519);
or U4040 (N_4040,In_2236,In_1331);
or U4041 (N_4041,In_557,In_2176);
nand U4042 (N_4042,In_1503,In_640);
and U4043 (N_4043,In_2010,In_1860);
nor U4044 (N_4044,In_637,In_519);
or U4045 (N_4045,In_895,In_105);
nand U4046 (N_4046,In_1714,In_1533);
and U4047 (N_4047,In_813,In_2148);
nand U4048 (N_4048,In_1814,In_838);
or U4049 (N_4049,In_65,In_925);
nand U4050 (N_4050,In_1469,In_1219);
and U4051 (N_4051,In_958,In_768);
and U4052 (N_4052,In_1819,In_1567);
nand U4053 (N_4053,In_2074,In_2170);
and U4054 (N_4054,In_1753,In_451);
xor U4055 (N_4055,In_811,In_1110);
xor U4056 (N_4056,In_1291,In_965);
xor U4057 (N_4057,In_1786,In_378);
nand U4058 (N_4058,In_1561,In_292);
nand U4059 (N_4059,In_883,In_634);
and U4060 (N_4060,In_618,In_1576);
xor U4061 (N_4061,In_735,In_865);
or U4062 (N_4062,In_1762,In_1109);
nor U4063 (N_4063,In_664,In_1415);
nor U4064 (N_4064,In_1560,In_1971);
xnor U4065 (N_4065,In_289,In_542);
and U4066 (N_4066,In_1934,In_2174);
xor U4067 (N_4067,In_1690,In_1970);
and U4068 (N_4068,In_454,In_2446);
or U4069 (N_4069,In_1163,In_1879);
nor U4070 (N_4070,In_1771,In_1800);
and U4071 (N_4071,In_365,In_553);
xor U4072 (N_4072,In_535,In_1936);
xnor U4073 (N_4073,In_1015,In_1318);
nand U4074 (N_4074,In_612,In_51);
or U4075 (N_4075,In_1735,In_364);
xnor U4076 (N_4076,In_250,In_1915);
nand U4077 (N_4077,In_2226,In_237);
xnor U4078 (N_4078,In_77,In_945);
and U4079 (N_4079,In_1750,In_1277);
nor U4080 (N_4080,In_2081,In_1432);
and U4081 (N_4081,In_580,In_2156);
xor U4082 (N_4082,In_1221,In_579);
and U4083 (N_4083,In_2200,In_873);
xor U4084 (N_4084,In_1132,In_884);
and U4085 (N_4085,In_2338,In_1351);
and U4086 (N_4086,In_1022,In_275);
xnor U4087 (N_4087,In_408,In_1133);
and U4088 (N_4088,In_2219,In_2194);
xor U4089 (N_4089,In_178,In_2259);
and U4090 (N_4090,In_2005,In_261);
xor U4091 (N_4091,In_2222,In_1269);
or U4092 (N_4092,In_373,In_1197);
and U4093 (N_4093,In_1941,In_2478);
nor U4094 (N_4094,In_1820,In_276);
or U4095 (N_4095,In_1318,In_974);
nand U4096 (N_4096,In_508,In_1183);
or U4097 (N_4097,In_29,In_1569);
nor U4098 (N_4098,In_2297,In_1295);
xnor U4099 (N_4099,In_2022,In_599);
and U4100 (N_4100,In_2220,In_1523);
or U4101 (N_4101,In_817,In_48);
nand U4102 (N_4102,In_1044,In_291);
xnor U4103 (N_4103,In_1379,In_1327);
nand U4104 (N_4104,In_1765,In_232);
xnor U4105 (N_4105,In_1221,In_1809);
and U4106 (N_4106,In_1118,In_1642);
xnor U4107 (N_4107,In_2214,In_954);
xnor U4108 (N_4108,In_1709,In_1537);
or U4109 (N_4109,In_1549,In_753);
nand U4110 (N_4110,In_335,In_2342);
nor U4111 (N_4111,In_1790,In_2018);
nand U4112 (N_4112,In_1663,In_2305);
nor U4113 (N_4113,In_1054,In_1891);
and U4114 (N_4114,In_363,In_918);
nor U4115 (N_4115,In_1352,In_2008);
and U4116 (N_4116,In_2488,In_1791);
xor U4117 (N_4117,In_967,In_858);
or U4118 (N_4118,In_133,In_770);
or U4119 (N_4119,In_190,In_804);
and U4120 (N_4120,In_2157,In_2191);
xnor U4121 (N_4121,In_24,In_320);
nand U4122 (N_4122,In_639,In_2343);
and U4123 (N_4123,In_183,In_1959);
xnor U4124 (N_4124,In_2178,In_1327);
and U4125 (N_4125,In_603,In_639);
or U4126 (N_4126,In_277,In_1974);
and U4127 (N_4127,In_1156,In_356);
nor U4128 (N_4128,In_2336,In_592);
or U4129 (N_4129,In_332,In_1585);
nand U4130 (N_4130,In_2082,In_335);
nand U4131 (N_4131,In_1645,In_1335);
and U4132 (N_4132,In_1882,In_1272);
xor U4133 (N_4133,In_2313,In_2166);
or U4134 (N_4134,In_939,In_1559);
nand U4135 (N_4135,In_88,In_2138);
or U4136 (N_4136,In_532,In_740);
or U4137 (N_4137,In_2320,In_2437);
nor U4138 (N_4138,In_784,In_1723);
or U4139 (N_4139,In_2252,In_848);
xnor U4140 (N_4140,In_2238,In_2022);
and U4141 (N_4141,In_947,In_1869);
and U4142 (N_4142,In_1892,In_264);
or U4143 (N_4143,In_1608,In_1687);
nand U4144 (N_4144,In_583,In_2302);
xnor U4145 (N_4145,In_2029,In_219);
nor U4146 (N_4146,In_908,In_5);
nand U4147 (N_4147,In_384,In_838);
nor U4148 (N_4148,In_1085,In_745);
nor U4149 (N_4149,In_773,In_1737);
or U4150 (N_4150,In_111,In_2330);
and U4151 (N_4151,In_554,In_1607);
and U4152 (N_4152,In_1373,In_664);
nand U4153 (N_4153,In_201,In_1111);
nor U4154 (N_4154,In_2007,In_1524);
and U4155 (N_4155,In_1651,In_1447);
nor U4156 (N_4156,In_915,In_1988);
xnor U4157 (N_4157,In_1885,In_1073);
xnor U4158 (N_4158,In_1002,In_880);
nor U4159 (N_4159,In_738,In_2120);
nand U4160 (N_4160,In_17,In_2331);
nor U4161 (N_4161,In_2322,In_1683);
nor U4162 (N_4162,In_2000,In_1122);
and U4163 (N_4163,In_2051,In_1822);
or U4164 (N_4164,In_1418,In_1241);
nand U4165 (N_4165,In_1517,In_645);
or U4166 (N_4166,In_702,In_155);
xor U4167 (N_4167,In_814,In_57);
nand U4168 (N_4168,In_1112,In_985);
nor U4169 (N_4169,In_496,In_2174);
nand U4170 (N_4170,In_153,In_2320);
xnor U4171 (N_4171,In_1293,In_644);
xnor U4172 (N_4172,In_2403,In_428);
and U4173 (N_4173,In_1101,In_2090);
nor U4174 (N_4174,In_2318,In_1621);
and U4175 (N_4175,In_1419,In_1629);
xnor U4176 (N_4176,In_87,In_1924);
nor U4177 (N_4177,In_898,In_341);
xnor U4178 (N_4178,In_1786,In_2272);
nor U4179 (N_4179,In_2365,In_2420);
xnor U4180 (N_4180,In_193,In_1844);
nand U4181 (N_4181,In_580,In_1933);
nor U4182 (N_4182,In_1532,In_1511);
and U4183 (N_4183,In_564,In_2120);
nand U4184 (N_4184,In_312,In_2178);
xor U4185 (N_4185,In_434,In_1190);
nand U4186 (N_4186,In_1679,In_1836);
or U4187 (N_4187,In_478,In_1652);
and U4188 (N_4188,In_1029,In_769);
nand U4189 (N_4189,In_1787,In_2420);
nand U4190 (N_4190,In_1745,In_794);
xnor U4191 (N_4191,In_1675,In_531);
and U4192 (N_4192,In_1907,In_799);
xor U4193 (N_4193,In_834,In_2401);
nor U4194 (N_4194,In_2317,In_856);
nor U4195 (N_4195,In_694,In_2457);
or U4196 (N_4196,In_790,In_647);
or U4197 (N_4197,In_1320,In_1981);
and U4198 (N_4198,In_1682,In_1805);
nor U4199 (N_4199,In_1721,In_2435);
or U4200 (N_4200,In_1443,In_963);
nand U4201 (N_4201,In_2264,In_6);
nor U4202 (N_4202,In_1909,In_2298);
xnor U4203 (N_4203,In_1839,In_2037);
and U4204 (N_4204,In_2202,In_39);
nor U4205 (N_4205,In_2152,In_1677);
and U4206 (N_4206,In_157,In_1091);
xor U4207 (N_4207,In_1987,In_63);
or U4208 (N_4208,In_657,In_982);
nand U4209 (N_4209,In_2493,In_497);
nor U4210 (N_4210,In_817,In_1520);
xnor U4211 (N_4211,In_346,In_457);
or U4212 (N_4212,In_1510,In_2393);
and U4213 (N_4213,In_2237,In_520);
nand U4214 (N_4214,In_1975,In_1103);
nand U4215 (N_4215,In_1376,In_2477);
and U4216 (N_4216,In_1280,In_321);
nand U4217 (N_4217,In_1478,In_964);
and U4218 (N_4218,In_17,In_1225);
nand U4219 (N_4219,In_1396,In_2364);
nand U4220 (N_4220,In_555,In_1365);
or U4221 (N_4221,In_16,In_2157);
or U4222 (N_4222,In_839,In_595);
nor U4223 (N_4223,In_1716,In_131);
or U4224 (N_4224,In_149,In_2171);
xor U4225 (N_4225,In_1034,In_1543);
and U4226 (N_4226,In_95,In_1693);
xor U4227 (N_4227,In_443,In_726);
or U4228 (N_4228,In_1028,In_668);
and U4229 (N_4229,In_607,In_216);
xnor U4230 (N_4230,In_1224,In_2437);
nor U4231 (N_4231,In_1398,In_1309);
and U4232 (N_4232,In_2307,In_2417);
and U4233 (N_4233,In_685,In_813);
xnor U4234 (N_4234,In_2120,In_2311);
or U4235 (N_4235,In_718,In_1877);
nand U4236 (N_4236,In_62,In_255);
nand U4237 (N_4237,In_2208,In_1815);
and U4238 (N_4238,In_729,In_1123);
nor U4239 (N_4239,In_1831,In_1609);
nor U4240 (N_4240,In_1539,In_970);
and U4241 (N_4241,In_940,In_1428);
and U4242 (N_4242,In_335,In_1955);
nor U4243 (N_4243,In_533,In_1304);
nor U4244 (N_4244,In_1922,In_812);
or U4245 (N_4245,In_332,In_898);
nand U4246 (N_4246,In_1839,In_2332);
nand U4247 (N_4247,In_2409,In_1542);
or U4248 (N_4248,In_308,In_2190);
nor U4249 (N_4249,In_574,In_2060);
or U4250 (N_4250,In_1421,In_1505);
xor U4251 (N_4251,In_1530,In_1305);
or U4252 (N_4252,In_256,In_111);
nand U4253 (N_4253,In_1012,In_2170);
nor U4254 (N_4254,In_1720,In_2041);
nand U4255 (N_4255,In_464,In_978);
or U4256 (N_4256,In_1402,In_367);
xor U4257 (N_4257,In_975,In_428);
or U4258 (N_4258,In_2238,In_2287);
nor U4259 (N_4259,In_1230,In_2100);
nor U4260 (N_4260,In_1002,In_135);
nor U4261 (N_4261,In_514,In_1541);
or U4262 (N_4262,In_1342,In_394);
and U4263 (N_4263,In_76,In_1976);
nand U4264 (N_4264,In_1731,In_904);
nor U4265 (N_4265,In_1753,In_1986);
or U4266 (N_4266,In_665,In_2477);
nand U4267 (N_4267,In_1232,In_440);
and U4268 (N_4268,In_249,In_1021);
and U4269 (N_4269,In_1220,In_567);
and U4270 (N_4270,In_2490,In_2483);
and U4271 (N_4271,In_1796,In_237);
xor U4272 (N_4272,In_416,In_548);
nand U4273 (N_4273,In_2359,In_1868);
xor U4274 (N_4274,In_400,In_920);
nor U4275 (N_4275,In_504,In_368);
nor U4276 (N_4276,In_692,In_1642);
xor U4277 (N_4277,In_128,In_1591);
or U4278 (N_4278,In_2334,In_2188);
xnor U4279 (N_4279,In_323,In_1799);
or U4280 (N_4280,In_2325,In_2045);
or U4281 (N_4281,In_1545,In_2054);
or U4282 (N_4282,In_1432,In_1016);
xor U4283 (N_4283,In_1956,In_2203);
nor U4284 (N_4284,In_1765,In_1677);
or U4285 (N_4285,In_58,In_258);
xor U4286 (N_4286,In_1608,In_1773);
nand U4287 (N_4287,In_895,In_614);
nor U4288 (N_4288,In_868,In_1366);
nand U4289 (N_4289,In_115,In_514);
nand U4290 (N_4290,In_2331,In_2005);
xnor U4291 (N_4291,In_1238,In_887);
or U4292 (N_4292,In_475,In_1820);
or U4293 (N_4293,In_2094,In_381);
nand U4294 (N_4294,In_667,In_2453);
and U4295 (N_4295,In_881,In_74);
nand U4296 (N_4296,In_2237,In_1022);
or U4297 (N_4297,In_695,In_1276);
or U4298 (N_4298,In_859,In_2489);
nor U4299 (N_4299,In_1102,In_1030);
nand U4300 (N_4300,In_920,In_103);
nor U4301 (N_4301,In_2055,In_1901);
and U4302 (N_4302,In_200,In_1375);
xor U4303 (N_4303,In_762,In_1168);
nor U4304 (N_4304,In_420,In_683);
xnor U4305 (N_4305,In_447,In_1068);
and U4306 (N_4306,In_1994,In_1242);
xor U4307 (N_4307,In_559,In_627);
or U4308 (N_4308,In_1883,In_211);
xor U4309 (N_4309,In_2468,In_693);
and U4310 (N_4310,In_1465,In_2453);
and U4311 (N_4311,In_2478,In_1398);
nand U4312 (N_4312,In_2217,In_189);
nand U4313 (N_4313,In_128,In_2306);
nand U4314 (N_4314,In_1740,In_327);
nand U4315 (N_4315,In_2230,In_1960);
and U4316 (N_4316,In_1580,In_1968);
or U4317 (N_4317,In_853,In_2010);
or U4318 (N_4318,In_1291,In_941);
xor U4319 (N_4319,In_1901,In_136);
and U4320 (N_4320,In_1304,In_2168);
or U4321 (N_4321,In_2322,In_1141);
or U4322 (N_4322,In_1973,In_159);
nor U4323 (N_4323,In_2447,In_1468);
and U4324 (N_4324,In_1157,In_2036);
nor U4325 (N_4325,In_362,In_1440);
and U4326 (N_4326,In_730,In_1500);
or U4327 (N_4327,In_1751,In_2095);
nor U4328 (N_4328,In_366,In_2488);
nand U4329 (N_4329,In_1624,In_265);
and U4330 (N_4330,In_1472,In_940);
and U4331 (N_4331,In_705,In_1030);
or U4332 (N_4332,In_420,In_1241);
xnor U4333 (N_4333,In_2120,In_779);
xor U4334 (N_4334,In_1821,In_2091);
xnor U4335 (N_4335,In_972,In_1066);
xor U4336 (N_4336,In_521,In_1207);
and U4337 (N_4337,In_294,In_764);
or U4338 (N_4338,In_53,In_800);
and U4339 (N_4339,In_1369,In_886);
or U4340 (N_4340,In_2308,In_1005);
nor U4341 (N_4341,In_1792,In_1641);
nor U4342 (N_4342,In_992,In_2154);
or U4343 (N_4343,In_557,In_2465);
xor U4344 (N_4344,In_329,In_196);
nor U4345 (N_4345,In_2468,In_1610);
nand U4346 (N_4346,In_77,In_2089);
nor U4347 (N_4347,In_1256,In_2328);
or U4348 (N_4348,In_843,In_1795);
and U4349 (N_4349,In_2463,In_2052);
xnor U4350 (N_4350,In_760,In_70);
or U4351 (N_4351,In_659,In_2246);
xnor U4352 (N_4352,In_97,In_2181);
or U4353 (N_4353,In_469,In_2361);
nor U4354 (N_4354,In_2493,In_1555);
or U4355 (N_4355,In_535,In_2087);
and U4356 (N_4356,In_46,In_880);
and U4357 (N_4357,In_467,In_1640);
xor U4358 (N_4358,In_144,In_846);
nand U4359 (N_4359,In_1403,In_1424);
nor U4360 (N_4360,In_2417,In_2097);
or U4361 (N_4361,In_1473,In_196);
nor U4362 (N_4362,In_1102,In_936);
or U4363 (N_4363,In_1859,In_2365);
and U4364 (N_4364,In_787,In_327);
nand U4365 (N_4365,In_2164,In_1608);
or U4366 (N_4366,In_1776,In_1231);
and U4367 (N_4367,In_1654,In_1542);
and U4368 (N_4368,In_219,In_294);
nor U4369 (N_4369,In_1623,In_1636);
xnor U4370 (N_4370,In_1930,In_983);
and U4371 (N_4371,In_2293,In_1910);
or U4372 (N_4372,In_370,In_1339);
xor U4373 (N_4373,In_1711,In_2390);
or U4374 (N_4374,In_2496,In_970);
and U4375 (N_4375,In_1304,In_1349);
or U4376 (N_4376,In_2436,In_415);
xnor U4377 (N_4377,In_736,In_199);
nor U4378 (N_4378,In_887,In_2372);
and U4379 (N_4379,In_1663,In_93);
or U4380 (N_4380,In_1363,In_674);
and U4381 (N_4381,In_2139,In_1540);
xnor U4382 (N_4382,In_281,In_964);
or U4383 (N_4383,In_435,In_624);
and U4384 (N_4384,In_435,In_337);
xor U4385 (N_4385,In_1950,In_663);
and U4386 (N_4386,In_1251,In_2120);
xor U4387 (N_4387,In_1016,In_676);
and U4388 (N_4388,In_1724,In_351);
or U4389 (N_4389,In_2077,In_2413);
and U4390 (N_4390,In_774,In_1488);
nor U4391 (N_4391,In_2429,In_1829);
or U4392 (N_4392,In_1805,In_2199);
or U4393 (N_4393,In_236,In_1608);
nor U4394 (N_4394,In_627,In_82);
or U4395 (N_4395,In_1044,In_1239);
nor U4396 (N_4396,In_1431,In_1991);
nor U4397 (N_4397,In_2387,In_1105);
nor U4398 (N_4398,In_979,In_1615);
nand U4399 (N_4399,In_1150,In_491);
or U4400 (N_4400,In_1487,In_637);
nand U4401 (N_4401,In_81,In_1744);
nand U4402 (N_4402,In_1329,In_257);
or U4403 (N_4403,In_1407,In_229);
and U4404 (N_4404,In_325,In_1802);
and U4405 (N_4405,In_401,In_2014);
nand U4406 (N_4406,In_1535,In_2364);
or U4407 (N_4407,In_1851,In_2056);
and U4408 (N_4408,In_2145,In_1996);
or U4409 (N_4409,In_410,In_1786);
xor U4410 (N_4410,In_1571,In_1427);
xnor U4411 (N_4411,In_1612,In_1193);
nor U4412 (N_4412,In_1968,In_1900);
xnor U4413 (N_4413,In_1449,In_1094);
xor U4414 (N_4414,In_1672,In_1946);
nand U4415 (N_4415,In_1285,In_701);
nand U4416 (N_4416,In_1639,In_1830);
nand U4417 (N_4417,In_1618,In_1710);
xor U4418 (N_4418,In_1661,In_445);
and U4419 (N_4419,In_1359,In_1272);
xnor U4420 (N_4420,In_601,In_1029);
or U4421 (N_4421,In_1213,In_2392);
nand U4422 (N_4422,In_247,In_1827);
or U4423 (N_4423,In_212,In_342);
and U4424 (N_4424,In_1459,In_891);
or U4425 (N_4425,In_664,In_113);
nand U4426 (N_4426,In_2384,In_2359);
xor U4427 (N_4427,In_476,In_209);
nand U4428 (N_4428,In_466,In_140);
nand U4429 (N_4429,In_1982,In_881);
nor U4430 (N_4430,In_310,In_2461);
nand U4431 (N_4431,In_852,In_1759);
xor U4432 (N_4432,In_1511,In_2184);
xor U4433 (N_4433,In_2073,In_2392);
xor U4434 (N_4434,In_928,In_179);
or U4435 (N_4435,In_813,In_1282);
nor U4436 (N_4436,In_2140,In_1967);
xor U4437 (N_4437,In_2180,In_2143);
nand U4438 (N_4438,In_49,In_174);
and U4439 (N_4439,In_302,In_1936);
or U4440 (N_4440,In_251,In_952);
nor U4441 (N_4441,In_309,In_894);
nor U4442 (N_4442,In_2470,In_2462);
nand U4443 (N_4443,In_1879,In_210);
nor U4444 (N_4444,In_301,In_2126);
or U4445 (N_4445,In_1572,In_703);
or U4446 (N_4446,In_486,In_748);
or U4447 (N_4447,In_1111,In_2211);
xor U4448 (N_4448,In_1033,In_1264);
or U4449 (N_4449,In_2327,In_1609);
and U4450 (N_4450,In_1024,In_2231);
and U4451 (N_4451,In_937,In_1474);
or U4452 (N_4452,In_301,In_2438);
and U4453 (N_4453,In_343,In_986);
nand U4454 (N_4454,In_652,In_2152);
and U4455 (N_4455,In_199,In_1012);
or U4456 (N_4456,In_837,In_248);
or U4457 (N_4457,In_1930,In_1784);
or U4458 (N_4458,In_845,In_50);
nor U4459 (N_4459,In_2166,In_326);
xnor U4460 (N_4460,In_664,In_1819);
and U4461 (N_4461,In_1503,In_11);
or U4462 (N_4462,In_2457,In_861);
and U4463 (N_4463,In_256,In_2360);
and U4464 (N_4464,In_1204,In_1492);
nor U4465 (N_4465,In_2262,In_462);
or U4466 (N_4466,In_1832,In_1590);
xnor U4467 (N_4467,In_1267,In_279);
and U4468 (N_4468,In_1597,In_473);
or U4469 (N_4469,In_2211,In_1860);
xor U4470 (N_4470,In_1796,In_1196);
nand U4471 (N_4471,In_393,In_1320);
nor U4472 (N_4472,In_1514,In_1085);
and U4473 (N_4473,In_351,In_510);
and U4474 (N_4474,In_2437,In_1179);
nor U4475 (N_4475,In_1766,In_709);
nor U4476 (N_4476,In_1409,In_980);
xnor U4477 (N_4477,In_720,In_1209);
nor U4478 (N_4478,In_2232,In_2273);
or U4479 (N_4479,In_1741,In_2073);
nor U4480 (N_4480,In_1109,In_1755);
or U4481 (N_4481,In_2357,In_334);
and U4482 (N_4482,In_1550,In_2121);
xor U4483 (N_4483,In_1085,In_592);
xor U4484 (N_4484,In_1097,In_1969);
and U4485 (N_4485,In_177,In_51);
nor U4486 (N_4486,In_501,In_993);
or U4487 (N_4487,In_1656,In_124);
xnor U4488 (N_4488,In_2311,In_697);
nand U4489 (N_4489,In_1993,In_617);
or U4490 (N_4490,In_1443,In_1520);
or U4491 (N_4491,In_972,In_942);
or U4492 (N_4492,In_87,In_1674);
nor U4493 (N_4493,In_1705,In_863);
or U4494 (N_4494,In_859,In_758);
xnor U4495 (N_4495,In_62,In_34);
nand U4496 (N_4496,In_2246,In_1815);
xnor U4497 (N_4497,In_94,In_1282);
or U4498 (N_4498,In_2216,In_2420);
xnor U4499 (N_4499,In_2293,In_2246);
nor U4500 (N_4500,In_1020,In_1745);
or U4501 (N_4501,In_2342,In_2324);
and U4502 (N_4502,In_529,In_1711);
nor U4503 (N_4503,In_107,In_1982);
xor U4504 (N_4504,In_70,In_1145);
xor U4505 (N_4505,In_415,In_2188);
and U4506 (N_4506,In_1502,In_2194);
xor U4507 (N_4507,In_1849,In_445);
nand U4508 (N_4508,In_2454,In_1566);
and U4509 (N_4509,In_760,In_1135);
nand U4510 (N_4510,In_1182,In_2209);
xnor U4511 (N_4511,In_391,In_1413);
nand U4512 (N_4512,In_2166,In_1980);
nor U4513 (N_4513,In_2060,In_1541);
and U4514 (N_4514,In_460,In_2349);
nor U4515 (N_4515,In_318,In_2102);
and U4516 (N_4516,In_2119,In_1903);
nand U4517 (N_4517,In_1088,In_820);
or U4518 (N_4518,In_1760,In_8);
xnor U4519 (N_4519,In_1760,In_545);
and U4520 (N_4520,In_0,In_201);
or U4521 (N_4521,In_1322,In_1757);
or U4522 (N_4522,In_1742,In_1055);
or U4523 (N_4523,In_979,In_1392);
nand U4524 (N_4524,In_1074,In_1053);
and U4525 (N_4525,In_850,In_323);
xnor U4526 (N_4526,In_2299,In_1384);
and U4527 (N_4527,In_2105,In_1412);
nor U4528 (N_4528,In_684,In_252);
or U4529 (N_4529,In_1670,In_1479);
or U4530 (N_4530,In_1121,In_1160);
and U4531 (N_4531,In_1764,In_2392);
or U4532 (N_4532,In_1879,In_2317);
and U4533 (N_4533,In_2357,In_2485);
or U4534 (N_4534,In_482,In_2317);
xor U4535 (N_4535,In_2430,In_2419);
xnor U4536 (N_4536,In_1858,In_2158);
nor U4537 (N_4537,In_2299,In_1142);
xor U4538 (N_4538,In_103,In_358);
nand U4539 (N_4539,In_1616,In_2415);
nand U4540 (N_4540,In_1467,In_1364);
nor U4541 (N_4541,In_902,In_1046);
xnor U4542 (N_4542,In_1386,In_2058);
nand U4543 (N_4543,In_1817,In_993);
nor U4544 (N_4544,In_1553,In_2350);
nand U4545 (N_4545,In_1228,In_720);
nand U4546 (N_4546,In_237,In_2000);
nor U4547 (N_4547,In_1628,In_2437);
nand U4548 (N_4548,In_1303,In_1910);
nand U4549 (N_4549,In_1915,In_385);
or U4550 (N_4550,In_1203,In_60);
or U4551 (N_4551,In_795,In_1315);
and U4552 (N_4552,In_724,In_520);
or U4553 (N_4553,In_2456,In_523);
xnor U4554 (N_4554,In_1140,In_2081);
or U4555 (N_4555,In_114,In_1540);
and U4556 (N_4556,In_1822,In_2124);
xor U4557 (N_4557,In_173,In_1072);
nand U4558 (N_4558,In_1332,In_1317);
xor U4559 (N_4559,In_1731,In_1899);
xor U4560 (N_4560,In_1586,In_2082);
and U4561 (N_4561,In_1646,In_1496);
and U4562 (N_4562,In_2321,In_888);
xnor U4563 (N_4563,In_1317,In_1230);
nand U4564 (N_4564,In_2366,In_449);
and U4565 (N_4565,In_1391,In_829);
or U4566 (N_4566,In_834,In_1724);
and U4567 (N_4567,In_1700,In_1556);
nand U4568 (N_4568,In_1026,In_1756);
nand U4569 (N_4569,In_683,In_838);
nor U4570 (N_4570,In_635,In_1983);
or U4571 (N_4571,In_1515,In_1151);
and U4572 (N_4572,In_273,In_28);
or U4573 (N_4573,In_1146,In_347);
and U4574 (N_4574,In_295,In_1643);
nor U4575 (N_4575,In_277,In_1543);
and U4576 (N_4576,In_1258,In_1445);
nor U4577 (N_4577,In_2062,In_800);
nor U4578 (N_4578,In_826,In_654);
nand U4579 (N_4579,In_2404,In_561);
nand U4580 (N_4580,In_1531,In_554);
xor U4581 (N_4581,In_1640,In_632);
nand U4582 (N_4582,In_1616,In_1557);
nor U4583 (N_4583,In_1931,In_2177);
nor U4584 (N_4584,In_1716,In_2491);
nor U4585 (N_4585,In_755,In_2);
nand U4586 (N_4586,In_82,In_2176);
or U4587 (N_4587,In_875,In_1137);
nand U4588 (N_4588,In_1055,In_624);
xor U4589 (N_4589,In_24,In_662);
nand U4590 (N_4590,In_887,In_1005);
xor U4591 (N_4591,In_1299,In_1395);
or U4592 (N_4592,In_1875,In_200);
xor U4593 (N_4593,In_2077,In_2445);
nand U4594 (N_4594,In_1039,In_195);
xor U4595 (N_4595,In_954,In_971);
xor U4596 (N_4596,In_2130,In_2045);
nand U4597 (N_4597,In_2142,In_488);
and U4598 (N_4598,In_1049,In_2065);
and U4599 (N_4599,In_454,In_2234);
xor U4600 (N_4600,In_1039,In_1014);
or U4601 (N_4601,In_1041,In_35);
xor U4602 (N_4602,In_1832,In_1728);
and U4603 (N_4603,In_214,In_658);
nand U4604 (N_4604,In_1935,In_1871);
xor U4605 (N_4605,In_2148,In_1928);
nor U4606 (N_4606,In_1502,In_959);
nand U4607 (N_4607,In_1335,In_2356);
or U4608 (N_4608,In_829,In_1428);
xnor U4609 (N_4609,In_232,In_1454);
nor U4610 (N_4610,In_116,In_563);
nor U4611 (N_4611,In_434,In_1112);
and U4612 (N_4612,In_1746,In_1086);
nor U4613 (N_4613,In_2011,In_1093);
or U4614 (N_4614,In_1696,In_251);
nand U4615 (N_4615,In_2364,In_989);
nand U4616 (N_4616,In_1487,In_1920);
nand U4617 (N_4617,In_369,In_2481);
nand U4618 (N_4618,In_1492,In_2168);
nand U4619 (N_4619,In_1423,In_1668);
xor U4620 (N_4620,In_1089,In_1482);
xor U4621 (N_4621,In_1329,In_2375);
xnor U4622 (N_4622,In_1570,In_1781);
and U4623 (N_4623,In_1019,In_379);
nor U4624 (N_4624,In_2044,In_308);
nor U4625 (N_4625,In_1510,In_2168);
nor U4626 (N_4626,In_1616,In_1684);
xnor U4627 (N_4627,In_663,In_690);
nor U4628 (N_4628,In_1565,In_1591);
and U4629 (N_4629,In_1022,In_1671);
and U4630 (N_4630,In_363,In_893);
xnor U4631 (N_4631,In_217,In_1945);
or U4632 (N_4632,In_456,In_2066);
xnor U4633 (N_4633,In_1668,In_1950);
xnor U4634 (N_4634,In_842,In_1663);
or U4635 (N_4635,In_662,In_1763);
nor U4636 (N_4636,In_1957,In_40);
xor U4637 (N_4637,In_2127,In_959);
nand U4638 (N_4638,In_1066,In_1005);
nor U4639 (N_4639,In_1546,In_25);
or U4640 (N_4640,In_231,In_1924);
and U4641 (N_4641,In_129,In_48);
and U4642 (N_4642,In_2161,In_274);
nor U4643 (N_4643,In_721,In_1288);
xnor U4644 (N_4644,In_648,In_875);
xnor U4645 (N_4645,In_2470,In_1827);
nor U4646 (N_4646,In_2229,In_1135);
nor U4647 (N_4647,In_1602,In_1946);
nand U4648 (N_4648,In_1271,In_2164);
nor U4649 (N_4649,In_773,In_33);
nand U4650 (N_4650,In_790,In_1735);
or U4651 (N_4651,In_113,In_1088);
nand U4652 (N_4652,In_2323,In_1480);
and U4653 (N_4653,In_1182,In_29);
xnor U4654 (N_4654,In_996,In_360);
and U4655 (N_4655,In_1851,In_2365);
nand U4656 (N_4656,In_1157,In_2076);
nand U4657 (N_4657,In_2464,In_1269);
xnor U4658 (N_4658,In_1836,In_2226);
nand U4659 (N_4659,In_1083,In_624);
or U4660 (N_4660,In_1956,In_1709);
xor U4661 (N_4661,In_429,In_61);
nand U4662 (N_4662,In_2088,In_1655);
nand U4663 (N_4663,In_1590,In_1849);
and U4664 (N_4664,In_1403,In_1778);
nand U4665 (N_4665,In_1133,In_2233);
or U4666 (N_4666,In_377,In_256);
and U4667 (N_4667,In_2023,In_1384);
and U4668 (N_4668,In_1067,In_1808);
or U4669 (N_4669,In_2143,In_678);
and U4670 (N_4670,In_416,In_157);
or U4671 (N_4671,In_927,In_2396);
xnor U4672 (N_4672,In_833,In_523);
xnor U4673 (N_4673,In_676,In_2010);
and U4674 (N_4674,In_622,In_186);
nand U4675 (N_4675,In_1828,In_291);
nand U4676 (N_4676,In_2233,In_1887);
or U4677 (N_4677,In_1392,In_986);
xnor U4678 (N_4678,In_1876,In_2234);
nand U4679 (N_4679,In_1909,In_838);
nand U4680 (N_4680,In_1066,In_1087);
nor U4681 (N_4681,In_2249,In_162);
or U4682 (N_4682,In_861,In_967);
or U4683 (N_4683,In_756,In_723);
nand U4684 (N_4684,In_1778,In_1907);
or U4685 (N_4685,In_2181,In_1039);
xor U4686 (N_4686,In_1571,In_654);
and U4687 (N_4687,In_2126,In_57);
or U4688 (N_4688,In_2300,In_331);
or U4689 (N_4689,In_2282,In_565);
or U4690 (N_4690,In_1206,In_2061);
nand U4691 (N_4691,In_258,In_753);
nand U4692 (N_4692,In_2325,In_38);
xor U4693 (N_4693,In_1650,In_675);
nor U4694 (N_4694,In_97,In_600);
or U4695 (N_4695,In_2234,In_2323);
nor U4696 (N_4696,In_212,In_1034);
and U4697 (N_4697,In_1286,In_2124);
nor U4698 (N_4698,In_1880,In_1718);
nand U4699 (N_4699,In_2359,In_510);
xor U4700 (N_4700,In_99,In_1244);
or U4701 (N_4701,In_394,In_2024);
xor U4702 (N_4702,In_1658,In_652);
nand U4703 (N_4703,In_1782,In_2368);
nor U4704 (N_4704,In_792,In_1362);
or U4705 (N_4705,In_1135,In_90);
or U4706 (N_4706,In_1709,In_354);
xnor U4707 (N_4707,In_997,In_1385);
nor U4708 (N_4708,In_2062,In_330);
nand U4709 (N_4709,In_84,In_611);
nand U4710 (N_4710,In_1610,In_2497);
nor U4711 (N_4711,In_1171,In_611);
xor U4712 (N_4712,In_2190,In_805);
xor U4713 (N_4713,In_1109,In_481);
nor U4714 (N_4714,In_2352,In_610);
xor U4715 (N_4715,In_1065,In_1716);
xor U4716 (N_4716,In_684,In_2353);
or U4717 (N_4717,In_1091,In_228);
and U4718 (N_4718,In_1459,In_1128);
xnor U4719 (N_4719,In_1642,In_1493);
xor U4720 (N_4720,In_704,In_1709);
and U4721 (N_4721,In_1935,In_586);
xor U4722 (N_4722,In_2113,In_1105);
nor U4723 (N_4723,In_1917,In_107);
and U4724 (N_4724,In_1054,In_1285);
or U4725 (N_4725,In_15,In_2065);
nand U4726 (N_4726,In_1005,In_2368);
nand U4727 (N_4727,In_1619,In_1733);
xor U4728 (N_4728,In_2233,In_1799);
or U4729 (N_4729,In_917,In_2104);
nand U4730 (N_4730,In_2220,In_262);
nand U4731 (N_4731,In_2321,In_182);
nor U4732 (N_4732,In_1898,In_2193);
xor U4733 (N_4733,In_943,In_2044);
and U4734 (N_4734,In_2472,In_2228);
nor U4735 (N_4735,In_1275,In_502);
xnor U4736 (N_4736,In_1945,In_304);
nand U4737 (N_4737,In_1580,In_194);
and U4738 (N_4738,In_398,In_1088);
nor U4739 (N_4739,In_734,In_1341);
nand U4740 (N_4740,In_460,In_239);
and U4741 (N_4741,In_1459,In_2390);
and U4742 (N_4742,In_430,In_2468);
nor U4743 (N_4743,In_956,In_174);
xor U4744 (N_4744,In_1177,In_1673);
nor U4745 (N_4745,In_1561,In_2133);
nor U4746 (N_4746,In_1561,In_2239);
nand U4747 (N_4747,In_829,In_1417);
and U4748 (N_4748,In_1778,In_687);
and U4749 (N_4749,In_1122,In_1178);
nor U4750 (N_4750,In_1268,In_691);
nor U4751 (N_4751,In_1672,In_1284);
or U4752 (N_4752,In_138,In_900);
nor U4753 (N_4753,In_722,In_1001);
xor U4754 (N_4754,In_1408,In_287);
nor U4755 (N_4755,In_928,In_1383);
xnor U4756 (N_4756,In_1890,In_2115);
nand U4757 (N_4757,In_39,In_654);
nand U4758 (N_4758,In_2230,In_2197);
xnor U4759 (N_4759,In_2261,In_1611);
or U4760 (N_4760,In_2304,In_353);
nand U4761 (N_4761,In_1292,In_8);
and U4762 (N_4762,In_2278,In_2008);
or U4763 (N_4763,In_266,In_2166);
and U4764 (N_4764,In_1927,In_7);
and U4765 (N_4765,In_1846,In_1343);
xnor U4766 (N_4766,In_2391,In_2337);
xor U4767 (N_4767,In_1568,In_1173);
and U4768 (N_4768,In_186,In_760);
nand U4769 (N_4769,In_1888,In_882);
or U4770 (N_4770,In_185,In_2417);
nand U4771 (N_4771,In_1268,In_167);
xor U4772 (N_4772,In_1465,In_1300);
or U4773 (N_4773,In_297,In_1989);
and U4774 (N_4774,In_691,In_1683);
nor U4775 (N_4775,In_459,In_346);
xor U4776 (N_4776,In_1836,In_1705);
or U4777 (N_4777,In_275,In_396);
nor U4778 (N_4778,In_1989,In_1547);
xor U4779 (N_4779,In_525,In_2327);
and U4780 (N_4780,In_993,In_1782);
and U4781 (N_4781,In_2249,In_892);
and U4782 (N_4782,In_1793,In_2339);
nand U4783 (N_4783,In_248,In_1843);
xor U4784 (N_4784,In_1976,In_2433);
nor U4785 (N_4785,In_1739,In_345);
nand U4786 (N_4786,In_2266,In_1054);
nand U4787 (N_4787,In_680,In_1779);
nand U4788 (N_4788,In_1259,In_1487);
and U4789 (N_4789,In_1470,In_98);
nor U4790 (N_4790,In_399,In_1258);
or U4791 (N_4791,In_1309,In_1723);
and U4792 (N_4792,In_2410,In_1961);
or U4793 (N_4793,In_705,In_794);
xnor U4794 (N_4794,In_2271,In_1245);
or U4795 (N_4795,In_1144,In_1616);
xor U4796 (N_4796,In_615,In_2088);
or U4797 (N_4797,In_1519,In_293);
nor U4798 (N_4798,In_2095,In_90);
or U4799 (N_4799,In_1860,In_1949);
nor U4800 (N_4800,In_893,In_1103);
and U4801 (N_4801,In_2392,In_577);
and U4802 (N_4802,In_1620,In_648);
nor U4803 (N_4803,In_1671,In_700);
nand U4804 (N_4804,In_1470,In_2212);
nor U4805 (N_4805,In_1895,In_750);
and U4806 (N_4806,In_1165,In_1435);
and U4807 (N_4807,In_746,In_2006);
or U4808 (N_4808,In_1166,In_2393);
and U4809 (N_4809,In_2443,In_1848);
and U4810 (N_4810,In_1012,In_1664);
or U4811 (N_4811,In_276,In_1898);
and U4812 (N_4812,In_353,In_1612);
and U4813 (N_4813,In_951,In_1946);
xor U4814 (N_4814,In_1445,In_1419);
xor U4815 (N_4815,In_2187,In_2134);
or U4816 (N_4816,In_2366,In_386);
nor U4817 (N_4817,In_727,In_1435);
xor U4818 (N_4818,In_734,In_2333);
and U4819 (N_4819,In_270,In_1510);
xor U4820 (N_4820,In_1874,In_568);
xnor U4821 (N_4821,In_1456,In_313);
nand U4822 (N_4822,In_428,In_421);
or U4823 (N_4823,In_1470,In_282);
nor U4824 (N_4824,In_1940,In_996);
xor U4825 (N_4825,In_1742,In_1595);
or U4826 (N_4826,In_1549,In_1650);
xor U4827 (N_4827,In_1067,In_952);
or U4828 (N_4828,In_462,In_1406);
xnor U4829 (N_4829,In_1745,In_439);
nor U4830 (N_4830,In_1803,In_1666);
nor U4831 (N_4831,In_73,In_2128);
or U4832 (N_4832,In_1435,In_264);
nor U4833 (N_4833,In_2270,In_2454);
nand U4834 (N_4834,In_1659,In_1824);
and U4835 (N_4835,In_1992,In_1592);
xor U4836 (N_4836,In_980,In_1293);
nand U4837 (N_4837,In_1956,In_2210);
xnor U4838 (N_4838,In_2156,In_1755);
nand U4839 (N_4839,In_2419,In_2489);
xnor U4840 (N_4840,In_2184,In_101);
nor U4841 (N_4841,In_1597,In_2475);
and U4842 (N_4842,In_947,In_1789);
xnor U4843 (N_4843,In_1440,In_170);
nand U4844 (N_4844,In_2364,In_191);
nor U4845 (N_4845,In_1878,In_1653);
xor U4846 (N_4846,In_1304,In_1923);
nand U4847 (N_4847,In_805,In_686);
nand U4848 (N_4848,In_1648,In_1923);
nand U4849 (N_4849,In_1207,In_1520);
nor U4850 (N_4850,In_2436,In_2256);
nor U4851 (N_4851,In_735,In_1186);
or U4852 (N_4852,In_2084,In_1751);
and U4853 (N_4853,In_820,In_314);
nand U4854 (N_4854,In_1349,In_349);
xor U4855 (N_4855,In_1116,In_2388);
nor U4856 (N_4856,In_1729,In_44);
xnor U4857 (N_4857,In_656,In_1560);
and U4858 (N_4858,In_1717,In_748);
nand U4859 (N_4859,In_1233,In_104);
nor U4860 (N_4860,In_1706,In_1623);
nand U4861 (N_4861,In_2243,In_2258);
nand U4862 (N_4862,In_661,In_2004);
xor U4863 (N_4863,In_2342,In_1433);
nand U4864 (N_4864,In_2250,In_2138);
nor U4865 (N_4865,In_839,In_2203);
nand U4866 (N_4866,In_1346,In_662);
or U4867 (N_4867,In_2254,In_1054);
xor U4868 (N_4868,In_578,In_2413);
and U4869 (N_4869,In_1654,In_1693);
nand U4870 (N_4870,In_184,In_1110);
or U4871 (N_4871,In_1168,In_1478);
and U4872 (N_4872,In_1882,In_391);
and U4873 (N_4873,In_859,In_911);
and U4874 (N_4874,In_1900,In_2182);
and U4875 (N_4875,In_1466,In_943);
xor U4876 (N_4876,In_1938,In_141);
and U4877 (N_4877,In_1254,In_2172);
and U4878 (N_4878,In_1625,In_899);
nor U4879 (N_4879,In_674,In_1859);
nand U4880 (N_4880,In_1681,In_538);
nor U4881 (N_4881,In_1675,In_59);
xnor U4882 (N_4882,In_1984,In_378);
nand U4883 (N_4883,In_1400,In_2315);
nor U4884 (N_4884,In_2199,In_464);
nor U4885 (N_4885,In_1535,In_1251);
or U4886 (N_4886,In_2083,In_859);
nand U4887 (N_4887,In_1970,In_1079);
nand U4888 (N_4888,In_1972,In_1247);
nor U4889 (N_4889,In_2313,In_2278);
and U4890 (N_4890,In_404,In_1958);
nor U4891 (N_4891,In_315,In_2035);
nand U4892 (N_4892,In_117,In_878);
nor U4893 (N_4893,In_1806,In_1819);
and U4894 (N_4894,In_1265,In_1675);
xor U4895 (N_4895,In_472,In_1258);
nor U4896 (N_4896,In_1114,In_587);
and U4897 (N_4897,In_87,In_994);
and U4898 (N_4898,In_988,In_2284);
or U4899 (N_4899,In_1548,In_1939);
or U4900 (N_4900,In_1456,In_1569);
and U4901 (N_4901,In_819,In_1619);
or U4902 (N_4902,In_1785,In_570);
or U4903 (N_4903,In_2180,In_1779);
xor U4904 (N_4904,In_1274,In_2406);
or U4905 (N_4905,In_1323,In_764);
or U4906 (N_4906,In_427,In_1849);
xor U4907 (N_4907,In_478,In_2171);
nor U4908 (N_4908,In_204,In_1618);
nor U4909 (N_4909,In_767,In_2036);
xor U4910 (N_4910,In_1443,In_439);
and U4911 (N_4911,In_851,In_333);
nand U4912 (N_4912,In_1799,In_67);
and U4913 (N_4913,In_1146,In_1736);
xnor U4914 (N_4914,In_219,In_2309);
xnor U4915 (N_4915,In_611,In_1433);
nor U4916 (N_4916,In_1540,In_40);
xor U4917 (N_4917,In_669,In_2239);
nand U4918 (N_4918,In_1773,In_443);
or U4919 (N_4919,In_1853,In_2290);
and U4920 (N_4920,In_2314,In_479);
or U4921 (N_4921,In_4,In_1137);
xor U4922 (N_4922,In_2040,In_297);
or U4923 (N_4923,In_1353,In_277);
nor U4924 (N_4924,In_1253,In_449);
and U4925 (N_4925,In_1330,In_461);
xnor U4926 (N_4926,In_2139,In_895);
xor U4927 (N_4927,In_1185,In_1653);
xor U4928 (N_4928,In_237,In_978);
and U4929 (N_4929,In_1207,In_1597);
nor U4930 (N_4930,In_2057,In_2123);
nand U4931 (N_4931,In_592,In_2153);
or U4932 (N_4932,In_2171,In_641);
xor U4933 (N_4933,In_517,In_851);
nand U4934 (N_4934,In_2477,In_624);
and U4935 (N_4935,In_424,In_1977);
or U4936 (N_4936,In_2317,In_493);
or U4937 (N_4937,In_493,In_380);
and U4938 (N_4938,In_2121,In_1540);
and U4939 (N_4939,In_2053,In_1565);
nand U4940 (N_4940,In_512,In_977);
and U4941 (N_4941,In_323,In_263);
nand U4942 (N_4942,In_429,In_1697);
nand U4943 (N_4943,In_1522,In_523);
nor U4944 (N_4944,In_1806,In_1843);
nor U4945 (N_4945,In_826,In_605);
or U4946 (N_4946,In_1119,In_469);
and U4947 (N_4947,In_654,In_556);
xnor U4948 (N_4948,In_501,In_533);
or U4949 (N_4949,In_1507,In_2435);
nand U4950 (N_4950,In_191,In_779);
nand U4951 (N_4951,In_753,In_1279);
xor U4952 (N_4952,In_852,In_759);
nand U4953 (N_4953,In_1890,In_1526);
and U4954 (N_4954,In_755,In_1730);
or U4955 (N_4955,In_2395,In_182);
nor U4956 (N_4956,In_496,In_2163);
nand U4957 (N_4957,In_2457,In_1302);
xor U4958 (N_4958,In_550,In_233);
nor U4959 (N_4959,In_1586,In_559);
nor U4960 (N_4960,In_1052,In_802);
nand U4961 (N_4961,In_605,In_348);
xnor U4962 (N_4962,In_1695,In_1192);
or U4963 (N_4963,In_1299,In_449);
xor U4964 (N_4964,In_223,In_2311);
or U4965 (N_4965,In_856,In_2075);
or U4966 (N_4966,In_1277,In_1338);
nand U4967 (N_4967,In_1706,In_2311);
nand U4968 (N_4968,In_1792,In_773);
nand U4969 (N_4969,In_2293,In_302);
xor U4970 (N_4970,In_110,In_820);
xnor U4971 (N_4971,In_1728,In_889);
and U4972 (N_4972,In_448,In_511);
or U4973 (N_4973,In_1833,In_150);
nor U4974 (N_4974,In_2116,In_1416);
xnor U4975 (N_4975,In_848,In_2324);
nand U4976 (N_4976,In_1826,In_2471);
nor U4977 (N_4977,In_927,In_1377);
and U4978 (N_4978,In_446,In_988);
and U4979 (N_4979,In_1833,In_2234);
nor U4980 (N_4980,In_2320,In_1548);
nand U4981 (N_4981,In_818,In_2236);
and U4982 (N_4982,In_2319,In_2325);
nand U4983 (N_4983,In_2477,In_174);
and U4984 (N_4984,In_2258,In_1887);
or U4985 (N_4985,In_949,In_2060);
nand U4986 (N_4986,In_2042,In_2228);
xnor U4987 (N_4987,In_2066,In_1103);
nor U4988 (N_4988,In_1352,In_2264);
nor U4989 (N_4989,In_2082,In_2331);
xnor U4990 (N_4990,In_2106,In_1273);
nand U4991 (N_4991,In_1544,In_1178);
nor U4992 (N_4992,In_1326,In_1115);
nor U4993 (N_4993,In_1406,In_321);
nor U4994 (N_4994,In_1776,In_813);
and U4995 (N_4995,In_286,In_196);
xnor U4996 (N_4996,In_347,In_253);
nor U4997 (N_4997,In_897,In_614);
xnor U4998 (N_4998,In_1938,In_1676);
or U4999 (N_4999,In_1680,In_1085);
or U5000 (N_5000,In_2424,In_1890);
nand U5001 (N_5001,In_2005,In_1763);
nor U5002 (N_5002,In_1814,In_1986);
nor U5003 (N_5003,In_526,In_2279);
nor U5004 (N_5004,In_509,In_1362);
nand U5005 (N_5005,In_956,In_1829);
or U5006 (N_5006,In_437,In_2027);
nor U5007 (N_5007,In_1147,In_1562);
xor U5008 (N_5008,In_1104,In_2310);
and U5009 (N_5009,In_1279,In_317);
nor U5010 (N_5010,In_887,In_74);
xor U5011 (N_5011,In_1861,In_479);
xnor U5012 (N_5012,In_755,In_2176);
nand U5013 (N_5013,In_2382,In_338);
or U5014 (N_5014,In_679,In_438);
and U5015 (N_5015,In_1989,In_2383);
nand U5016 (N_5016,In_556,In_323);
nand U5017 (N_5017,In_2067,In_1318);
nand U5018 (N_5018,In_55,In_1112);
nor U5019 (N_5019,In_436,In_1396);
nor U5020 (N_5020,In_1754,In_1627);
xnor U5021 (N_5021,In_2241,In_1656);
nor U5022 (N_5022,In_1662,In_1812);
xnor U5023 (N_5023,In_903,In_613);
xor U5024 (N_5024,In_1719,In_2448);
nand U5025 (N_5025,In_2446,In_1494);
xor U5026 (N_5026,In_39,In_200);
nand U5027 (N_5027,In_909,In_2120);
or U5028 (N_5028,In_2319,In_1495);
and U5029 (N_5029,In_1283,In_1338);
or U5030 (N_5030,In_229,In_93);
xor U5031 (N_5031,In_1142,In_1445);
and U5032 (N_5032,In_1631,In_2417);
or U5033 (N_5033,In_1148,In_1075);
xnor U5034 (N_5034,In_1038,In_888);
nand U5035 (N_5035,In_96,In_2138);
nand U5036 (N_5036,In_126,In_1495);
nand U5037 (N_5037,In_280,In_403);
nor U5038 (N_5038,In_498,In_1693);
or U5039 (N_5039,In_2296,In_1881);
nand U5040 (N_5040,In_83,In_1551);
or U5041 (N_5041,In_2353,In_12);
nor U5042 (N_5042,In_1858,In_887);
and U5043 (N_5043,In_1467,In_71);
and U5044 (N_5044,In_329,In_1913);
xnor U5045 (N_5045,In_482,In_237);
nor U5046 (N_5046,In_630,In_2293);
nor U5047 (N_5047,In_158,In_1233);
or U5048 (N_5048,In_1661,In_145);
nor U5049 (N_5049,In_2061,In_1130);
nor U5050 (N_5050,In_1706,In_2374);
xnor U5051 (N_5051,In_946,In_460);
nor U5052 (N_5052,In_1824,In_1849);
nand U5053 (N_5053,In_1643,In_1450);
nor U5054 (N_5054,In_1288,In_1883);
nor U5055 (N_5055,In_1080,In_726);
nand U5056 (N_5056,In_1072,In_1938);
and U5057 (N_5057,In_2451,In_1508);
nand U5058 (N_5058,In_2060,In_2233);
nand U5059 (N_5059,In_761,In_618);
or U5060 (N_5060,In_395,In_1224);
nand U5061 (N_5061,In_1468,In_1146);
nand U5062 (N_5062,In_384,In_1200);
and U5063 (N_5063,In_1963,In_1543);
and U5064 (N_5064,In_1785,In_438);
nand U5065 (N_5065,In_1744,In_2270);
nand U5066 (N_5066,In_2170,In_2470);
and U5067 (N_5067,In_1723,In_1965);
nand U5068 (N_5068,In_717,In_1305);
xor U5069 (N_5069,In_803,In_2187);
nand U5070 (N_5070,In_2418,In_275);
nor U5071 (N_5071,In_2429,In_1267);
xor U5072 (N_5072,In_882,In_2015);
xor U5073 (N_5073,In_2027,In_1766);
xor U5074 (N_5074,In_619,In_1312);
and U5075 (N_5075,In_772,In_1613);
nand U5076 (N_5076,In_980,In_1899);
xor U5077 (N_5077,In_171,In_1230);
or U5078 (N_5078,In_437,In_1518);
nor U5079 (N_5079,In_1318,In_1435);
nand U5080 (N_5080,In_2051,In_1503);
xor U5081 (N_5081,In_73,In_2357);
nand U5082 (N_5082,In_1838,In_2155);
and U5083 (N_5083,In_339,In_955);
or U5084 (N_5084,In_756,In_621);
nand U5085 (N_5085,In_2391,In_781);
xnor U5086 (N_5086,In_515,In_759);
and U5087 (N_5087,In_1049,In_2010);
or U5088 (N_5088,In_2078,In_1301);
xor U5089 (N_5089,In_120,In_1779);
or U5090 (N_5090,In_1197,In_1187);
nand U5091 (N_5091,In_1312,In_922);
and U5092 (N_5092,In_2268,In_1838);
or U5093 (N_5093,In_549,In_984);
nor U5094 (N_5094,In_362,In_1278);
nor U5095 (N_5095,In_1401,In_2317);
or U5096 (N_5096,In_319,In_1131);
xnor U5097 (N_5097,In_903,In_1660);
xnor U5098 (N_5098,In_1105,In_664);
nor U5099 (N_5099,In_2419,In_949);
xor U5100 (N_5100,In_684,In_254);
and U5101 (N_5101,In_1015,In_1530);
nand U5102 (N_5102,In_248,In_1477);
and U5103 (N_5103,In_456,In_42);
xnor U5104 (N_5104,In_2342,In_1474);
nor U5105 (N_5105,In_1883,In_1657);
xnor U5106 (N_5106,In_27,In_1097);
xnor U5107 (N_5107,In_1420,In_395);
or U5108 (N_5108,In_2297,In_188);
nand U5109 (N_5109,In_2216,In_976);
and U5110 (N_5110,In_2215,In_1297);
or U5111 (N_5111,In_751,In_465);
nor U5112 (N_5112,In_2400,In_1468);
nand U5113 (N_5113,In_2311,In_125);
nand U5114 (N_5114,In_2208,In_286);
xor U5115 (N_5115,In_1932,In_2449);
nor U5116 (N_5116,In_54,In_2121);
or U5117 (N_5117,In_433,In_1700);
xor U5118 (N_5118,In_1229,In_96);
and U5119 (N_5119,In_2139,In_2172);
nand U5120 (N_5120,In_780,In_1210);
nand U5121 (N_5121,In_384,In_2039);
nand U5122 (N_5122,In_1465,In_1101);
nor U5123 (N_5123,In_1510,In_1936);
and U5124 (N_5124,In_600,In_1234);
nand U5125 (N_5125,In_1626,In_1949);
nand U5126 (N_5126,In_1171,In_659);
or U5127 (N_5127,In_820,In_1035);
and U5128 (N_5128,In_2118,In_93);
xnor U5129 (N_5129,In_1585,In_2088);
and U5130 (N_5130,In_832,In_723);
nor U5131 (N_5131,In_1583,In_1144);
nor U5132 (N_5132,In_2281,In_2144);
nor U5133 (N_5133,In_374,In_2443);
nand U5134 (N_5134,In_2244,In_356);
xnor U5135 (N_5135,In_819,In_501);
and U5136 (N_5136,In_1761,In_2184);
or U5137 (N_5137,In_116,In_2368);
nand U5138 (N_5138,In_2435,In_2175);
xor U5139 (N_5139,In_1984,In_1342);
nor U5140 (N_5140,In_452,In_2106);
nor U5141 (N_5141,In_1006,In_2437);
or U5142 (N_5142,In_1347,In_1430);
or U5143 (N_5143,In_2127,In_1248);
and U5144 (N_5144,In_1395,In_2311);
nor U5145 (N_5145,In_1447,In_1831);
or U5146 (N_5146,In_687,In_1099);
nand U5147 (N_5147,In_2061,In_1535);
and U5148 (N_5148,In_248,In_1403);
nor U5149 (N_5149,In_2368,In_2208);
or U5150 (N_5150,In_383,In_524);
and U5151 (N_5151,In_932,In_240);
xnor U5152 (N_5152,In_1696,In_1244);
or U5153 (N_5153,In_2469,In_1545);
or U5154 (N_5154,In_485,In_791);
and U5155 (N_5155,In_717,In_389);
or U5156 (N_5156,In_1939,In_1531);
nand U5157 (N_5157,In_2372,In_438);
xnor U5158 (N_5158,In_1184,In_1275);
xor U5159 (N_5159,In_2162,In_643);
xnor U5160 (N_5160,In_214,In_2197);
or U5161 (N_5161,In_1998,In_878);
and U5162 (N_5162,In_1880,In_1466);
or U5163 (N_5163,In_1741,In_1194);
nand U5164 (N_5164,In_2094,In_2409);
and U5165 (N_5165,In_990,In_1005);
xor U5166 (N_5166,In_2093,In_794);
nor U5167 (N_5167,In_1801,In_2412);
nand U5168 (N_5168,In_571,In_1836);
nand U5169 (N_5169,In_1029,In_817);
nand U5170 (N_5170,In_1406,In_69);
or U5171 (N_5171,In_1515,In_318);
nor U5172 (N_5172,In_1040,In_1451);
nor U5173 (N_5173,In_914,In_137);
and U5174 (N_5174,In_1752,In_682);
or U5175 (N_5175,In_1152,In_1139);
nor U5176 (N_5176,In_2319,In_806);
and U5177 (N_5177,In_318,In_748);
nor U5178 (N_5178,In_1587,In_1805);
nor U5179 (N_5179,In_382,In_2144);
and U5180 (N_5180,In_1267,In_778);
nand U5181 (N_5181,In_1496,In_1037);
xnor U5182 (N_5182,In_2151,In_1631);
nor U5183 (N_5183,In_1589,In_359);
and U5184 (N_5184,In_2497,In_55);
and U5185 (N_5185,In_255,In_2152);
xnor U5186 (N_5186,In_683,In_6);
nand U5187 (N_5187,In_1623,In_545);
xor U5188 (N_5188,In_891,In_1399);
nor U5189 (N_5189,In_912,In_64);
and U5190 (N_5190,In_1335,In_2190);
and U5191 (N_5191,In_1370,In_45);
xor U5192 (N_5192,In_1251,In_2248);
xnor U5193 (N_5193,In_615,In_482);
nor U5194 (N_5194,In_376,In_2043);
or U5195 (N_5195,In_290,In_1491);
xor U5196 (N_5196,In_2095,In_2379);
xnor U5197 (N_5197,In_1790,In_470);
nor U5198 (N_5198,In_2220,In_403);
or U5199 (N_5199,In_499,In_1344);
nand U5200 (N_5200,In_1784,In_912);
nor U5201 (N_5201,In_2379,In_2173);
nand U5202 (N_5202,In_2459,In_1064);
and U5203 (N_5203,In_386,In_1973);
nor U5204 (N_5204,In_2249,In_961);
nand U5205 (N_5205,In_2126,In_489);
xor U5206 (N_5206,In_1036,In_2334);
and U5207 (N_5207,In_2483,In_581);
or U5208 (N_5208,In_1548,In_1579);
nor U5209 (N_5209,In_794,In_2484);
or U5210 (N_5210,In_613,In_564);
and U5211 (N_5211,In_1048,In_1356);
and U5212 (N_5212,In_1803,In_2170);
nor U5213 (N_5213,In_2130,In_709);
and U5214 (N_5214,In_125,In_832);
and U5215 (N_5215,In_1438,In_1410);
xor U5216 (N_5216,In_49,In_1817);
nand U5217 (N_5217,In_2431,In_433);
or U5218 (N_5218,In_163,In_1208);
xnor U5219 (N_5219,In_2303,In_825);
or U5220 (N_5220,In_1105,In_1041);
or U5221 (N_5221,In_1527,In_633);
nand U5222 (N_5222,In_484,In_138);
nand U5223 (N_5223,In_914,In_717);
nor U5224 (N_5224,In_1649,In_1660);
xor U5225 (N_5225,In_248,In_1019);
xnor U5226 (N_5226,In_864,In_226);
and U5227 (N_5227,In_1038,In_1911);
nor U5228 (N_5228,In_1750,In_207);
and U5229 (N_5229,In_1505,In_2362);
or U5230 (N_5230,In_17,In_908);
nand U5231 (N_5231,In_250,In_1597);
or U5232 (N_5232,In_827,In_365);
nand U5233 (N_5233,In_15,In_1635);
and U5234 (N_5234,In_2362,In_1770);
and U5235 (N_5235,In_1627,In_668);
nor U5236 (N_5236,In_2205,In_2352);
nand U5237 (N_5237,In_633,In_1557);
nor U5238 (N_5238,In_1674,In_2434);
and U5239 (N_5239,In_2323,In_2272);
nand U5240 (N_5240,In_1229,In_25);
nand U5241 (N_5241,In_46,In_677);
or U5242 (N_5242,In_2161,In_1014);
and U5243 (N_5243,In_1708,In_1334);
nand U5244 (N_5244,In_695,In_1569);
xor U5245 (N_5245,In_1129,In_878);
nor U5246 (N_5246,In_116,In_822);
xnor U5247 (N_5247,In_1988,In_1406);
nand U5248 (N_5248,In_1210,In_492);
or U5249 (N_5249,In_689,In_779);
or U5250 (N_5250,In_2327,In_2167);
xor U5251 (N_5251,In_363,In_1968);
xor U5252 (N_5252,In_1408,In_197);
and U5253 (N_5253,In_2320,In_238);
and U5254 (N_5254,In_501,In_39);
and U5255 (N_5255,In_2148,In_1171);
xnor U5256 (N_5256,In_2436,In_2111);
or U5257 (N_5257,In_352,In_1971);
nand U5258 (N_5258,In_2018,In_2022);
nor U5259 (N_5259,In_1009,In_1231);
nor U5260 (N_5260,In_2288,In_1796);
or U5261 (N_5261,In_741,In_811);
nor U5262 (N_5262,In_1731,In_1318);
or U5263 (N_5263,In_1883,In_127);
or U5264 (N_5264,In_125,In_1207);
or U5265 (N_5265,In_1427,In_528);
nor U5266 (N_5266,In_1964,In_320);
nor U5267 (N_5267,In_1034,In_1665);
or U5268 (N_5268,In_1135,In_159);
or U5269 (N_5269,In_321,In_580);
or U5270 (N_5270,In_2458,In_585);
and U5271 (N_5271,In_2354,In_2296);
nor U5272 (N_5272,In_81,In_990);
or U5273 (N_5273,In_1272,In_210);
xnor U5274 (N_5274,In_363,In_460);
and U5275 (N_5275,In_68,In_1659);
nand U5276 (N_5276,In_2280,In_1055);
or U5277 (N_5277,In_2358,In_461);
or U5278 (N_5278,In_1890,In_218);
nand U5279 (N_5279,In_2375,In_2460);
or U5280 (N_5280,In_1317,In_64);
and U5281 (N_5281,In_1127,In_2475);
xor U5282 (N_5282,In_927,In_879);
and U5283 (N_5283,In_1732,In_1332);
and U5284 (N_5284,In_315,In_1377);
and U5285 (N_5285,In_1826,In_1194);
nand U5286 (N_5286,In_1322,In_832);
nand U5287 (N_5287,In_745,In_1688);
nand U5288 (N_5288,In_2483,In_2134);
nand U5289 (N_5289,In_706,In_2386);
or U5290 (N_5290,In_1707,In_1746);
nor U5291 (N_5291,In_635,In_1747);
and U5292 (N_5292,In_1666,In_1362);
nor U5293 (N_5293,In_1938,In_251);
xor U5294 (N_5294,In_1668,In_1843);
and U5295 (N_5295,In_558,In_743);
and U5296 (N_5296,In_250,In_1790);
nor U5297 (N_5297,In_2352,In_1407);
or U5298 (N_5298,In_2253,In_1733);
and U5299 (N_5299,In_277,In_1990);
or U5300 (N_5300,In_1601,In_2436);
nand U5301 (N_5301,In_1205,In_706);
nand U5302 (N_5302,In_2243,In_200);
nor U5303 (N_5303,In_1642,In_300);
xor U5304 (N_5304,In_1899,In_1413);
xor U5305 (N_5305,In_494,In_294);
nand U5306 (N_5306,In_1995,In_1236);
nor U5307 (N_5307,In_1250,In_678);
nand U5308 (N_5308,In_581,In_2482);
and U5309 (N_5309,In_2109,In_2206);
xor U5310 (N_5310,In_2214,In_1801);
and U5311 (N_5311,In_1144,In_1973);
xnor U5312 (N_5312,In_935,In_2389);
xor U5313 (N_5313,In_1411,In_1500);
or U5314 (N_5314,In_2125,In_82);
xor U5315 (N_5315,In_330,In_1745);
nor U5316 (N_5316,In_657,In_1939);
or U5317 (N_5317,In_1995,In_1093);
and U5318 (N_5318,In_1558,In_1443);
nor U5319 (N_5319,In_622,In_1268);
nor U5320 (N_5320,In_1363,In_1481);
and U5321 (N_5321,In_884,In_1544);
xor U5322 (N_5322,In_1825,In_157);
nor U5323 (N_5323,In_1046,In_1595);
nor U5324 (N_5324,In_533,In_2231);
or U5325 (N_5325,In_347,In_1471);
nor U5326 (N_5326,In_692,In_499);
nor U5327 (N_5327,In_2206,In_2094);
xor U5328 (N_5328,In_749,In_41);
nand U5329 (N_5329,In_337,In_2217);
nor U5330 (N_5330,In_704,In_1548);
nor U5331 (N_5331,In_2419,In_1982);
xnor U5332 (N_5332,In_1775,In_481);
xor U5333 (N_5333,In_1915,In_1955);
xnor U5334 (N_5334,In_92,In_1929);
and U5335 (N_5335,In_2168,In_296);
xor U5336 (N_5336,In_1882,In_2458);
and U5337 (N_5337,In_2439,In_1340);
nand U5338 (N_5338,In_1995,In_370);
xor U5339 (N_5339,In_520,In_896);
nand U5340 (N_5340,In_1100,In_92);
and U5341 (N_5341,In_545,In_617);
or U5342 (N_5342,In_1114,In_269);
nand U5343 (N_5343,In_533,In_1080);
or U5344 (N_5344,In_185,In_983);
and U5345 (N_5345,In_1207,In_1052);
or U5346 (N_5346,In_243,In_828);
and U5347 (N_5347,In_65,In_2083);
xor U5348 (N_5348,In_161,In_847);
and U5349 (N_5349,In_891,In_1995);
xor U5350 (N_5350,In_1887,In_776);
nand U5351 (N_5351,In_21,In_1447);
nand U5352 (N_5352,In_659,In_1444);
nor U5353 (N_5353,In_858,In_2011);
nor U5354 (N_5354,In_838,In_222);
xnor U5355 (N_5355,In_620,In_1922);
and U5356 (N_5356,In_781,In_810);
nand U5357 (N_5357,In_2286,In_2370);
nand U5358 (N_5358,In_461,In_325);
nor U5359 (N_5359,In_1791,In_1779);
or U5360 (N_5360,In_1127,In_2443);
and U5361 (N_5361,In_2340,In_237);
nand U5362 (N_5362,In_651,In_2330);
nand U5363 (N_5363,In_462,In_802);
and U5364 (N_5364,In_2421,In_1179);
nor U5365 (N_5365,In_225,In_852);
xnor U5366 (N_5366,In_829,In_1367);
and U5367 (N_5367,In_2351,In_1338);
nor U5368 (N_5368,In_847,In_1201);
and U5369 (N_5369,In_1748,In_2212);
nor U5370 (N_5370,In_1061,In_1070);
xnor U5371 (N_5371,In_2446,In_2318);
nand U5372 (N_5372,In_2148,In_580);
nor U5373 (N_5373,In_1684,In_1561);
or U5374 (N_5374,In_326,In_628);
nor U5375 (N_5375,In_1777,In_2334);
xnor U5376 (N_5376,In_1057,In_1412);
and U5377 (N_5377,In_819,In_411);
nand U5378 (N_5378,In_2261,In_86);
nand U5379 (N_5379,In_753,In_191);
nand U5380 (N_5380,In_1789,In_1524);
and U5381 (N_5381,In_1546,In_564);
and U5382 (N_5382,In_1223,In_1069);
nor U5383 (N_5383,In_1312,In_224);
and U5384 (N_5384,In_1984,In_1749);
xor U5385 (N_5385,In_1235,In_889);
nor U5386 (N_5386,In_1905,In_2494);
nor U5387 (N_5387,In_1401,In_1286);
and U5388 (N_5388,In_184,In_2131);
xnor U5389 (N_5389,In_35,In_167);
and U5390 (N_5390,In_1555,In_1112);
or U5391 (N_5391,In_1449,In_248);
nand U5392 (N_5392,In_453,In_2090);
nor U5393 (N_5393,In_120,In_343);
xor U5394 (N_5394,In_1008,In_30);
and U5395 (N_5395,In_1905,In_1601);
xnor U5396 (N_5396,In_439,In_2105);
xor U5397 (N_5397,In_2477,In_2162);
nor U5398 (N_5398,In_1670,In_1449);
nand U5399 (N_5399,In_808,In_1379);
xnor U5400 (N_5400,In_1967,In_1608);
xor U5401 (N_5401,In_1339,In_484);
or U5402 (N_5402,In_880,In_1835);
and U5403 (N_5403,In_692,In_1787);
nand U5404 (N_5404,In_1860,In_2166);
or U5405 (N_5405,In_1366,In_1331);
xor U5406 (N_5406,In_548,In_1945);
and U5407 (N_5407,In_1932,In_2314);
xor U5408 (N_5408,In_1581,In_782);
xor U5409 (N_5409,In_1128,In_1469);
nor U5410 (N_5410,In_1737,In_186);
nand U5411 (N_5411,In_131,In_2196);
or U5412 (N_5412,In_1848,In_380);
and U5413 (N_5413,In_1988,In_127);
xnor U5414 (N_5414,In_1169,In_1487);
or U5415 (N_5415,In_873,In_772);
nand U5416 (N_5416,In_1609,In_248);
and U5417 (N_5417,In_2369,In_31);
nand U5418 (N_5418,In_859,In_37);
or U5419 (N_5419,In_2215,In_189);
nor U5420 (N_5420,In_425,In_286);
xnor U5421 (N_5421,In_162,In_2089);
nand U5422 (N_5422,In_1594,In_2298);
nand U5423 (N_5423,In_1166,In_1137);
and U5424 (N_5424,In_2422,In_1962);
nand U5425 (N_5425,In_348,In_2117);
xor U5426 (N_5426,In_1269,In_1620);
xnor U5427 (N_5427,In_1500,In_851);
nand U5428 (N_5428,In_2333,In_2050);
nand U5429 (N_5429,In_297,In_778);
and U5430 (N_5430,In_922,In_1020);
nor U5431 (N_5431,In_2239,In_2328);
nand U5432 (N_5432,In_817,In_306);
nor U5433 (N_5433,In_2168,In_1086);
nand U5434 (N_5434,In_229,In_2334);
and U5435 (N_5435,In_1205,In_1303);
nor U5436 (N_5436,In_2408,In_1061);
and U5437 (N_5437,In_1868,In_738);
nor U5438 (N_5438,In_1282,In_1331);
nand U5439 (N_5439,In_501,In_19);
nand U5440 (N_5440,In_856,In_706);
or U5441 (N_5441,In_314,In_323);
xnor U5442 (N_5442,In_2052,In_763);
nor U5443 (N_5443,In_976,In_1748);
nor U5444 (N_5444,In_176,In_2165);
nand U5445 (N_5445,In_900,In_160);
and U5446 (N_5446,In_1573,In_2266);
nand U5447 (N_5447,In_1304,In_909);
nand U5448 (N_5448,In_1965,In_682);
or U5449 (N_5449,In_842,In_219);
nand U5450 (N_5450,In_797,In_423);
or U5451 (N_5451,In_2293,In_1007);
nand U5452 (N_5452,In_2495,In_1134);
xor U5453 (N_5453,In_949,In_1371);
nor U5454 (N_5454,In_1195,In_1017);
or U5455 (N_5455,In_1165,In_772);
xor U5456 (N_5456,In_2115,In_1923);
nor U5457 (N_5457,In_2069,In_2158);
nor U5458 (N_5458,In_1527,In_1878);
nor U5459 (N_5459,In_1151,In_453);
nand U5460 (N_5460,In_421,In_1595);
or U5461 (N_5461,In_1440,In_1790);
or U5462 (N_5462,In_1165,In_490);
nor U5463 (N_5463,In_1298,In_1736);
or U5464 (N_5464,In_607,In_486);
nor U5465 (N_5465,In_2057,In_1962);
xor U5466 (N_5466,In_2101,In_2050);
nand U5467 (N_5467,In_1114,In_1488);
and U5468 (N_5468,In_514,In_1283);
xnor U5469 (N_5469,In_262,In_475);
nand U5470 (N_5470,In_1889,In_2477);
or U5471 (N_5471,In_172,In_1816);
xnor U5472 (N_5472,In_942,In_241);
or U5473 (N_5473,In_1358,In_1531);
and U5474 (N_5474,In_1272,In_1572);
nor U5475 (N_5475,In_332,In_191);
and U5476 (N_5476,In_2098,In_1824);
xor U5477 (N_5477,In_204,In_2217);
or U5478 (N_5478,In_677,In_60);
or U5479 (N_5479,In_1439,In_1545);
nor U5480 (N_5480,In_629,In_109);
xor U5481 (N_5481,In_920,In_1622);
or U5482 (N_5482,In_509,In_300);
nor U5483 (N_5483,In_487,In_1004);
or U5484 (N_5484,In_176,In_142);
nand U5485 (N_5485,In_681,In_2256);
or U5486 (N_5486,In_328,In_1810);
xor U5487 (N_5487,In_1992,In_409);
xnor U5488 (N_5488,In_836,In_506);
and U5489 (N_5489,In_1061,In_866);
nand U5490 (N_5490,In_1403,In_1937);
nor U5491 (N_5491,In_2135,In_75);
or U5492 (N_5492,In_1853,In_2250);
nor U5493 (N_5493,In_1672,In_1034);
and U5494 (N_5494,In_2013,In_222);
xor U5495 (N_5495,In_1141,In_1897);
or U5496 (N_5496,In_512,In_1226);
xnor U5497 (N_5497,In_2279,In_448);
nor U5498 (N_5498,In_361,In_2461);
nand U5499 (N_5499,In_2253,In_1031);
nor U5500 (N_5500,In_680,In_2169);
xor U5501 (N_5501,In_2282,In_1784);
xnor U5502 (N_5502,In_1879,In_1594);
xor U5503 (N_5503,In_1626,In_2121);
nor U5504 (N_5504,In_64,In_1612);
nand U5505 (N_5505,In_618,In_1088);
xor U5506 (N_5506,In_1255,In_1770);
nor U5507 (N_5507,In_1935,In_168);
xor U5508 (N_5508,In_1919,In_684);
or U5509 (N_5509,In_1418,In_908);
xor U5510 (N_5510,In_29,In_1823);
or U5511 (N_5511,In_524,In_1495);
or U5512 (N_5512,In_858,In_393);
or U5513 (N_5513,In_2111,In_141);
or U5514 (N_5514,In_1274,In_2);
or U5515 (N_5515,In_632,In_1341);
nand U5516 (N_5516,In_1218,In_340);
xor U5517 (N_5517,In_330,In_261);
nand U5518 (N_5518,In_1509,In_2469);
nor U5519 (N_5519,In_969,In_2178);
or U5520 (N_5520,In_971,In_964);
and U5521 (N_5521,In_2443,In_1280);
nand U5522 (N_5522,In_2196,In_1674);
nand U5523 (N_5523,In_2380,In_1630);
or U5524 (N_5524,In_1374,In_1770);
and U5525 (N_5525,In_154,In_2173);
nand U5526 (N_5526,In_45,In_209);
xnor U5527 (N_5527,In_716,In_1272);
xor U5528 (N_5528,In_1092,In_499);
nand U5529 (N_5529,In_1270,In_749);
nand U5530 (N_5530,In_558,In_465);
nand U5531 (N_5531,In_2154,In_1893);
nand U5532 (N_5532,In_309,In_2419);
nand U5533 (N_5533,In_1126,In_1385);
nand U5534 (N_5534,In_1872,In_1755);
and U5535 (N_5535,In_566,In_340);
or U5536 (N_5536,In_2043,In_1741);
xnor U5537 (N_5537,In_1876,In_1751);
and U5538 (N_5538,In_1785,In_1344);
or U5539 (N_5539,In_2388,In_1696);
nand U5540 (N_5540,In_1232,In_246);
xnor U5541 (N_5541,In_1331,In_333);
and U5542 (N_5542,In_1399,In_1353);
xnor U5543 (N_5543,In_108,In_1001);
and U5544 (N_5544,In_1997,In_622);
and U5545 (N_5545,In_6,In_1374);
xnor U5546 (N_5546,In_1612,In_1843);
or U5547 (N_5547,In_1323,In_252);
nor U5548 (N_5548,In_419,In_261);
xnor U5549 (N_5549,In_1845,In_2343);
and U5550 (N_5550,In_1819,In_52);
xnor U5551 (N_5551,In_1785,In_322);
and U5552 (N_5552,In_296,In_46);
nor U5553 (N_5553,In_2148,In_2135);
xnor U5554 (N_5554,In_1466,In_166);
nand U5555 (N_5555,In_37,In_1178);
and U5556 (N_5556,In_193,In_2219);
and U5557 (N_5557,In_2301,In_1591);
nor U5558 (N_5558,In_2347,In_2062);
nand U5559 (N_5559,In_1441,In_330);
and U5560 (N_5560,In_174,In_2076);
or U5561 (N_5561,In_1258,In_1944);
nor U5562 (N_5562,In_2245,In_1101);
or U5563 (N_5563,In_1230,In_2394);
nand U5564 (N_5564,In_1185,In_995);
nand U5565 (N_5565,In_711,In_1166);
or U5566 (N_5566,In_159,In_1199);
and U5567 (N_5567,In_1849,In_1180);
nor U5568 (N_5568,In_2178,In_846);
nand U5569 (N_5569,In_671,In_512);
xnor U5570 (N_5570,In_1738,In_330);
nand U5571 (N_5571,In_479,In_2220);
or U5572 (N_5572,In_1979,In_792);
or U5573 (N_5573,In_1114,In_2277);
nand U5574 (N_5574,In_751,In_1070);
nor U5575 (N_5575,In_2185,In_315);
nor U5576 (N_5576,In_0,In_1743);
and U5577 (N_5577,In_947,In_1545);
nor U5578 (N_5578,In_841,In_2117);
xor U5579 (N_5579,In_1843,In_1799);
and U5580 (N_5580,In_903,In_343);
xnor U5581 (N_5581,In_301,In_2338);
nor U5582 (N_5582,In_191,In_2052);
or U5583 (N_5583,In_1470,In_1503);
nand U5584 (N_5584,In_323,In_573);
or U5585 (N_5585,In_1166,In_334);
or U5586 (N_5586,In_1575,In_1270);
or U5587 (N_5587,In_2061,In_540);
or U5588 (N_5588,In_822,In_2399);
nor U5589 (N_5589,In_831,In_1218);
nand U5590 (N_5590,In_692,In_2417);
or U5591 (N_5591,In_2089,In_1852);
and U5592 (N_5592,In_832,In_457);
nor U5593 (N_5593,In_2285,In_531);
and U5594 (N_5594,In_1376,In_1132);
and U5595 (N_5595,In_1807,In_185);
or U5596 (N_5596,In_2185,In_1994);
or U5597 (N_5597,In_2013,In_1825);
xnor U5598 (N_5598,In_1,In_158);
xor U5599 (N_5599,In_639,In_2090);
xor U5600 (N_5600,In_2169,In_821);
nor U5601 (N_5601,In_2262,In_605);
and U5602 (N_5602,In_1524,In_1340);
and U5603 (N_5603,In_2467,In_2258);
xnor U5604 (N_5604,In_889,In_2086);
or U5605 (N_5605,In_2215,In_313);
or U5606 (N_5606,In_1282,In_2281);
and U5607 (N_5607,In_2204,In_816);
nand U5608 (N_5608,In_2408,In_2157);
nor U5609 (N_5609,In_1363,In_601);
xor U5610 (N_5610,In_1271,In_710);
xnor U5611 (N_5611,In_1016,In_129);
nor U5612 (N_5612,In_737,In_29);
xor U5613 (N_5613,In_1357,In_371);
nand U5614 (N_5614,In_2143,In_1068);
and U5615 (N_5615,In_2093,In_1743);
nand U5616 (N_5616,In_387,In_1144);
or U5617 (N_5617,In_660,In_769);
nor U5618 (N_5618,In_1412,In_792);
or U5619 (N_5619,In_1944,In_1928);
and U5620 (N_5620,In_949,In_178);
and U5621 (N_5621,In_1183,In_450);
xor U5622 (N_5622,In_1043,In_357);
xor U5623 (N_5623,In_829,In_456);
nor U5624 (N_5624,In_1501,In_1331);
and U5625 (N_5625,In_572,In_695);
xnor U5626 (N_5626,In_2232,In_1308);
nand U5627 (N_5627,In_1368,In_2408);
xor U5628 (N_5628,In_870,In_2228);
and U5629 (N_5629,In_1648,In_2019);
xor U5630 (N_5630,In_1146,In_1111);
xnor U5631 (N_5631,In_2040,In_1332);
nor U5632 (N_5632,In_2164,In_1386);
nor U5633 (N_5633,In_1239,In_2104);
nor U5634 (N_5634,In_896,In_2341);
nand U5635 (N_5635,In_507,In_2346);
or U5636 (N_5636,In_434,In_32);
xnor U5637 (N_5637,In_557,In_386);
and U5638 (N_5638,In_1712,In_1068);
and U5639 (N_5639,In_2297,In_2131);
or U5640 (N_5640,In_306,In_123);
xnor U5641 (N_5641,In_2033,In_494);
nand U5642 (N_5642,In_2184,In_2260);
or U5643 (N_5643,In_1194,In_2153);
nand U5644 (N_5644,In_1822,In_782);
and U5645 (N_5645,In_829,In_175);
xnor U5646 (N_5646,In_572,In_468);
nand U5647 (N_5647,In_2072,In_2017);
nor U5648 (N_5648,In_1737,In_561);
nor U5649 (N_5649,In_2230,In_1071);
nand U5650 (N_5650,In_1050,In_2494);
nor U5651 (N_5651,In_2366,In_496);
nand U5652 (N_5652,In_2319,In_984);
xnor U5653 (N_5653,In_1121,In_2212);
nand U5654 (N_5654,In_267,In_941);
xnor U5655 (N_5655,In_1766,In_42);
or U5656 (N_5656,In_2434,In_1975);
nand U5657 (N_5657,In_2086,In_87);
xor U5658 (N_5658,In_1224,In_1519);
xnor U5659 (N_5659,In_2451,In_2481);
or U5660 (N_5660,In_2047,In_836);
nand U5661 (N_5661,In_1643,In_1038);
nand U5662 (N_5662,In_861,In_435);
nand U5663 (N_5663,In_2349,In_607);
and U5664 (N_5664,In_1656,In_2104);
nand U5665 (N_5665,In_1464,In_883);
nor U5666 (N_5666,In_868,In_968);
nor U5667 (N_5667,In_2286,In_1190);
xnor U5668 (N_5668,In_2187,In_667);
and U5669 (N_5669,In_1559,In_2056);
xnor U5670 (N_5670,In_2428,In_955);
nand U5671 (N_5671,In_1359,In_2106);
nand U5672 (N_5672,In_16,In_1571);
nor U5673 (N_5673,In_572,In_1928);
and U5674 (N_5674,In_819,In_1355);
nand U5675 (N_5675,In_871,In_373);
nand U5676 (N_5676,In_1521,In_1619);
xor U5677 (N_5677,In_2240,In_613);
xnor U5678 (N_5678,In_1329,In_977);
nor U5679 (N_5679,In_985,In_1709);
or U5680 (N_5680,In_507,In_1355);
nand U5681 (N_5681,In_1385,In_610);
nand U5682 (N_5682,In_386,In_267);
nand U5683 (N_5683,In_1676,In_1477);
or U5684 (N_5684,In_623,In_2085);
nand U5685 (N_5685,In_509,In_1058);
or U5686 (N_5686,In_2314,In_2311);
xor U5687 (N_5687,In_755,In_39);
and U5688 (N_5688,In_666,In_393);
and U5689 (N_5689,In_355,In_1207);
or U5690 (N_5690,In_1377,In_1684);
or U5691 (N_5691,In_821,In_392);
or U5692 (N_5692,In_81,In_1801);
xor U5693 (N_5693,In_1254,In_1884);
nor U5694 (N_5694,In_1510,In_1442);
nand U5695 (N_5695,In_101,In_609);
xor U5696 (N_5696,In_1768,In_1472);
xor U5697 (N_5697,In_21,In_412);
or U5698 (N_5698,In_851,In_601);
or U5699 (N_5699,In_1419,In_23);
and U5700 (N_5700,In_2163,In_1868);
nand U5701 (N_5701,In_2146,In_1493);
xor U5702 (N_5702,In_519,In_1746);
and U5703 (N_5703,In_1323,In_1686);
nor U5704 (N_5704,In_1913,In_914);
nor U5705 (N_5705,In_2032,In_10);
and U5706 (N_5706,In_738,In_1315);
xor U5707 (N_5707,In_72,In_789);
xor U5708 (N_5708,In_350,In_800);
nor U5709 (N_5709,In_1399,In_118);
xnor U5710 (N_5710,In_370,In_0);
or U5711 (N_5711,In_2371,In_2225);
xnor U5712 (N_5712,In_2329,In_850);
nor U5713 (N_5713,In_1325,In_46);
xnor U5714 (N_5714,In_966,In_1648);
and U5715 (N_5715,In_1802,In_1923);
nand U5716 (N_5716,In_1555,In_1207);
nor U5717 (N_5717,In_934,In_2184);
or U5718 (N_5718,In_1460,In_1431);
nand U5719 (N_5719,In_1118,In_2319);
or U5720 (N_5720,In_1391,In_1888);
and U5721 (N_5721,In_2436,In_1393);
nand U5722 (N_5722,In_161,In_453);
nand U5723 (N_5723,In_1599,In_1647);
and U5724 (N_5724,In_145,In_1341);
or U5725 (N_5725,In_1703,In_904);
or U5726 (N_5726,In_22,In_1423);
nor U5727 (N_5727,In_322,In_1892);
nand U5728 (N_5728,In_1412,In_2281);
or U5729 (N_5729,In_2375,In_1911);
nand U5730 (N_5730,In_1454,In_1005);
and U5731 (N_5731,In_1749,In_702);
nor U5732 (N_5732,In_606,In_1950);
xor U5733 (N_5733,In_2454,In_1071);
nand U5734 (N_5734,In_610,In_768);
nor U5735 (N_5735,In_1672,In_13);
xor U5736 (N_5736,In_1416,In_1244);
nand U5737 (N_5737,In_2490,In_840);
xnor U5738 (N_5738,In_2219,In_786);
xnor U5739 (N_5739,In_1286,In_695);
or U5740 (N_5740,In_615,In_242);
xnor U5741 (N_5741,In_1657,In_104);
nand U5742 (N_5742,In_439,In_1139);
and U5743 (N_5743,In_829,In_1496);
or U5744 (N_5744,In_133,In_1378);
or U5745 (N_5745,In_2,In_2128);
and U5746 (N_5746,In_1363,In_594);
or U5747 (N_5747,In_577,In_2161);
or U5748 (N_5748,In_631,In_1665);
nand U5749 (N_5749,In_2300,In_842);
nand U5750 (N_5750,In_1741,In_1135);
nor U5751 (N_5751,In_703,In_2216);
nand U5752 (N_5752,In_1669,In_665);
or U5753 (N_5753,In_1716,In_38);
nand U5754 (N_5754,In_460,In_2055);
nor U5755 (N_5755,In_2188,In_2264);
or U5756 (N_5756,In_534,In_2297);
or U5757 (N_5757,In_2221,In_761);
and U5758 (N_5758,In_1868,In_2091);
xor U5759 (N_5759,In_49,In_1891);
nand U5760 (N_5760,In_2370,In_802);
xnor U5761 (N_5761,In_2189,In_1056);
nor U5762 (N_5762,In_352,In_19);
and U5763 (N_5763,In_1990,In_161);
nand U5764 (N_5764,In_2310,In_2174);
or U5765 (N_5765,In_1692,In_856);
xor U5766 (N_5766,In_1790,In_49);
nand U5767 (N_5767,In_1592,In_1153);
nand U5768 (N_5768,In_1762,In_2155);
nor U5769 (N_5769,In_1376,In_2363);
and U5770 (N_5770,In_288,In_627);
and U5771 (N_5771,In_2309,In_129);
nor U5772 (N_5772,In_2439,In_1517);
nor U5773 (N_5773,In_1069,In_2030);
nor U5774 (N_5774,In_2182,In_693);
or U5775 (N_5775,In_1579,In_1088);
nor U5776 (N_5776,In_1545,In_959);
or U5777 (N_5777,In_1744,In_654);
nand U5778 (N_5778,In_2017,In_84);
xor U5779 (N_5779,In_421,In_2309);
and U5780 (N_5780,In_134,In_569);
nand U5781 (N_5781,In_660,In_132);
nand U5782 (N_5782,In_2468,In_1252);
or U5783 (N_5783,In_815,In_50);
and U5784 (N_5784,In_686,In_291);
nor U5785 (N_5785,In_66,In_1411);
and U5786 (N_5786,In_1114,In_874);
xnor U5787 (N_5787,In_782,In_1227);
nor U5788 (N_5788,In_2421,In_2391);
nand U5789 (N_5789,In_1612,In_794);
or U5790 (N_5790,In_1189,In_305);
xor U5791 (N_5791,In_1977,In_2067);
nand U5792 (N_5792,In_212,In_2496);
nand U5793 (N_5793,In_861,In_926);
and U5794 (N_5794,In_1344,In_2184);
or U5795 (N_5795,In_1485,In_701);
nand U5796 (N_5796,In_2052,In_1084);
or U5797 (N_5797,In_993,In_1278);
nand U5798 (N_5798,In_214,In_1973);
nor U5799 (N_5799,In_735,In_2080);
nand U5800 (N_5800,In_405,In_503);
nand U5801 (N_5801,In_437,In_320);
or U5802 (N_5802,In_192,In_1175);
and U5803 (N_5803,In_438,In_638);
or U5804 (N_5804,In_1144,In_130);
and U5805 (N_5805,In_1326,In_2340);
xor U5806 (N_5806,In_1844,In_1019);
nand U5807 (N_5807,In_133,In_394);
xnor U5808 (N_5808,In_919,In_952);
or U5809 (N_5809,In_2394,In_1511);
xor U5810 (N_5810,In_1463,In_944);
xnor U5811 (N_5811,In_2246,In_825);
xnor U5812 (N_5812,In_1842,In_2493);
nor U5813 (N_5813,In_177,In_547);
and U5814 (N_5814,In_2109,In_1603);
and U5815 (N_5815,In_872,In_7);
xnor U5816 (N_5816,In_364,In_2359);
nand U5817 (N_5817,In_188,In_1724);
and U5818 (N_5818,In_914,In_1812);
nor U5819 (N_5819,In_882,In_184);
xnor U5820 (N_5820,In_1325,In_1627);
nand U5821 (N_5821,In_497,In_1635);
nor U5822 (N_5822,In_908,In_1387);
xor U5823 (N_5823,In_1113,In_2195);
nand U5824 (N_5824,In_427,In_679);
xnor U5825 (N_5825,In_2484,In_2011);
nor U5826 (N_5826,In_2282,In_1446);
nand U5827 (N_5827,In_1403,In_1964);
or U5828 (N_5828,In_1914,In_1540);
nor U5829 (N_5829,In_1185,In_820);
or U5830 (N_5830,In_1425,In_232);
or U5831 (N_5831,In_1049,In_1972);
or U5832 (N_5832,In_467,In_2456);
nand U5833 (N_5833,In_135,In_2044);
or U5834 (N_5834,In_718,In_1696);
nor U5835 (N_5835,In_1970,In_183);
or U5836 (N_5836,In_785,In_362);
or U5837 (N_5837,In_521,In_1787);
xnor U5838 (N_5838,In_1233,In_1252);
nor U5839 (N_5839,In_2373,In_2407);
xor U5840 (N_5840,In_998,In_47);
nor U5841 (N_5841,In_2160,In_2080);
or U5842 (N_5842,In_2315,In_2392);
nor U5843 (N_5843,In_447,In_1644);
nand U5844 (N_5844,In_1945,In_160);
nor U5845 (N_5845,In_2492,In_1750);
xor U5846 (N_5846,In_2486,In_147);
and U5847 (N_5847,In_1754,In_355);
and U5848 (N_5848,In_1132,In_1012);
nand U5849 (N_5849,In_2110,In_1998);
or U5850 (N_5850,In_2024,In_1751);
and U5851 (N_5851,In_2371,In_514);
and U5852 (N_5852,In_728,In_1460);
xnor U5853 (N_5853,In_870,In_1649);
and U5854 (N_5854,In_261,In_700);
or U5855 (N_5855,In_2157,In_1043);
and U5856 (N_5856,In_1689,In_2021);
nor U5857 (N_5857,In_2081,In_1383);
nand U5858 (N_5858,In_1746,In_904);
or U5859 (N_5859,In_2216,In_1849);
xnor U5860 (N_5860,In_679,In_842);
xnor U5861 (N_5861,In_878,In_397);
or U5862 (N_5862,In_324,In_1146);
nand U5863 (N_5863,In_1751,In_200);
nor U5864 (N_5864,In_659,In_2096);
nor U5865 (N_5865,In_708,In_1758);
xnor U5866 (N_5866,In_1018,In_1501);
and U5867 (N_5867,In_802,In_826);
nor U5868 (N_5868,In_1342,In_1300);
nor U5869 (N_5869,In_438,In_1568);
nand U5870 (N_5870,In_663,In_1943);
and U5871 (N_5871,In_356,In_1948);
xor U5872 (N_5872,In_2491,In_1457);
or U5873 (N_5873,In_1050,In_471);
nor U5874 (N_5874,In_1106,In_1361);
and U5875 (N_5875,In_1771,In_1734);
nor U5876 (N_5876,In_2074,In_2274);
or U5877 (N_5877,In_768,In_290);
xnor U5878 (N_5878,In_2471,In_2461);
nand U5879 (N_5879,In_1021,In_2422);
and U5880 (N_5880,In_1751,In_624);
nor U5881 (N_5881,In_81,In_1771);
nand U5882 (N_5882,In_1277,In_1875);
xor U5883 (N_5883,In_1297,In_2059);
or U5884 (N_5884,In_294,In_1582);
or U5885 (N_5885,In_304,In_1042);
nand U5886 (N_5886,In_161,In_174);
nand U5887 (N_5887,In_653,In_2378);
or U5888 (N_5888,In_958,In_1023);
nor U5889 (N_5889,In_668,In_1050);
or U5890 (N_5890,In_1538,In_535);
nor U5891 (N_5891,In_2400,In_1575);
and U5892 (N_5892,In_858,In_1732);
and U5893 (N_5893,In_875,In_250);
and U5894 (N_5894,In_672,In_194);
xnor U5895 (N_5895,In_2197,In_1972);
and U5896 (N_5896,In_916,In_1025);
nor U5897 (N_5897,In_1504,In_232);
or U5898 (N_5898,In_1455,In_560);
xor U5899 (N_5899,In_1763,In_859);
nand U5900 (N_5900,In_497,In_327);
and U5901 (N_5901,In_257,In_2433);
and U5902 (N_5902,In_75,In_2352);
nand U5903 (N_5903,In_2311,In_520);
xnor U5904 (N_5904,In_740,In_1178);
and U5905 (N_5905,In_1489,In_89);
or U5906 (N_5906,In_900,In_1617);
nand U5907 (N_5907,In_280,In_1231);
or U5908 (N_5908,In_1261,In_17);
and U5909 (N_5909,In_1194,In_576);
nand U5910 (N_5910,In_413,In_938);
or U5911 (N_5911,In_1051,In_2168);
or U5912 (N_5912,In_1875,In_2025);
and U5913 (N_5913,In_503,In_1464);
or U5914 (N_5914,In_94,In_1627);
and U5915 (N_5915,In_999,In_159);
nand U5916 (N_5916,In_1933,In_2012);
xnor U5917 (N_5917,In_1774,In_633);
and U5918 (N_5918,In_1481,In_1772);
xor U5919 (N_5919,In_133,In_719);
xor U5920 (N_5920,In_1181,In_1112);
nand U5921 (N_5921,In_58,In_887);
nand U5922 (N_5922,In_1485,In_1028);
nor U5923 (N_5923,In_1141,In_214);
nand U5924 (N_5924,In_1209,In_2160);
and U5925 (N_5925,In_1059,In_1625);
nand U5926 (N_5926,In_815,In_1951);
and U5927 (N_5927,In_492,In_875);
nor U5928 (N_5928,In_1633,In_2410);
nand U5929 (N_5929,In_103,In_1842);
nand U5930 (N_5930,In_332,In_1178);
xnor U5931 (N_5931,In_1386,In_2211);
nor U5932 (N_5932,In_1729,In_138);
xnor U5933 (N_5933,In_2491,In_522);
nand U5934 (N_5934,In_2156,In_1495);
nand U5935 (N_5935,In_1064,In_151);
xnor U5936 (N_5936,In_525,In_672);
xor U5937 (N_5937,In_200,In_96);
nand U5938 (N_5938,In_172,In_2049);
nand U5939 (N_5939,In_2189,In_635);
nor U5940 (N_5940,In_1084,In_2118);
nand U5941 (N_5941,In_1366,In_2464);
or U5942 (N_5942,In_564,In_2046);
and U5943 (N_5943,In_587,In_1530);
nand U5944 (N_5944,In_24,In_745);
or U5945 (N_5945,In_285,In_2376);
and U5946 (N_5946,In_734,In_1552);
xnor U5947 (N_5947,In_2484,In_727);
and U5948 (N_5948,In_811,In_250);
nor U5949 (N_5949,In_315,In_1018);
nor U5950 (N_5950,In_1095,In_2119);
or U5951 (N_5951,In_2470,In_451);
xor U5952 (N_5952,In_2152,In_2450);
or U5953 (N_5953,In_2264,In_71);
or U5954 (N_5954,In_1339,In_659);
and U5955 (N_5955,In_1955,In_775);
and U5956 (N_5956,In_1254,In_1351);
nand U5957 (N_5957,In_892,In_2392);
nor U5958 (N_5958,In_773,In_2077);
nand U5959 (N_5959,In_915,In_340);
nand U5960 (N_5960,In_2078,In_901);
xnor U5961 (N_5961,In_39,In_1442);
nand U5962 (N_5962,In_1780,In_770);
and U5963 (N_5963,In_248,In_2434);
nand U5964 (N_5964,In_2368,In_1640);
and U5965 (N_5965,In_800,In_1325);
and U5966 (N_5966,In_177,In_2493);
nand U5967 (N_5967,In_1110,In_377);
and U5968 (N_5968,In_1935,In_1364);
nand U5969 (N_5969,In_1393,In_1006);
and U5970 (N_5970,In_853,In_1138);
nand U5971 (N_5971,In_562,In_2321);
xor U5972 (N_5972,In_423,In_202);
nor U5973 (N_5973,In_1398,In_542);
and U5974 (N_5974,In_1279,In_1378);
nand U5975 (N_5975,In_2071,In_1742);
xnor U5976 (N_5976,In_593,In_2383);
and U5977 (N_5977,In_1785,In_639);
or U5978 (N_5978,In_1748,In_2368);
or U5979 (N_5979,In_819,In_76);
xnor U5980 (N_5980,In_1512,In_1486);
and U5981 (N_5981,In_743,In_1538);
nand U5982 (N_5982,In_419,In_2198);
nand U5983 (N_5983,In_2349,In_346);
and U5984 (N_5984,In_2163,In_1966);
and U5985 (N_5985,In_1807,In_1201);
xnor U5986 (N_5986,In_1861,In_497);
xnor U5987 (N_5987,In_382,In_231);
and U5988 (N_5988,In_75,In_1655);
nor U5989 (N_5989,In_1906,In_1091);
nand U5990 (N_5990,In_2258,In_728);
and U5991 (N_5991,In_498,In_1985);
and U5992 (N_5992,In_2214,In_87);
nor U5993 (N_5993,In_857,In_1883);
or U5994 (N_5994,In_1464,In_2366);
nand U5995 (N_5995,In_2101,In_1053);
and U5996 (N_5996,In_805,In_294);
and U5997 (N_5997,In_2411,In_503);
xnor U5998 (N_5998,In_838,In_1741);
nor U5999 (N_5999,In_1440,In_168);
xor U6000 (N_6000,In_2218,In_929);
nand U6001 (N_6001,In_1923,In_2050);
or U6002 (N_6002,In_551,In_1690);
and U6003 (N_6003,In_623,In_1483);
nand U6004 (N_6004,In_349,In_1266);
nand U6005 (N_6005,In_669,In_1881);
nand U6006 (N_6006,In_163,In_2471);
nor U6007 (N_6007,In_983,In_2027);
xor U6008 (N_6008,In_728,In_1633);
nand U6009 (N_6009,In_81,In_468);
xnor U6010 (N_6010,In_1866,In_2005);
or U6011 (N_6011,In_867,In_2165);
or U6012 (N_6012,In_2279,In_1421);
or U6013 (N_6013,In_79,In_2482);
and U6014 (N_6014,In_364,In_152);
nand U6015 (N_6015,In_424,In_392);
and U6016 (N_6016,In_1231,In_1766);
xor U6017 (N_6017,In_2415,In_2295);
xor U6018 (N_6018,In_424,In_1032);
and U6019 (N_6019,In_797,In_2043);
nor U6020 (N_6020,In_2390,In_1104);
nor U6021 (N_6021,In_1828,In_438);
nand U6022 (N_6022,In_1527,In_1854);
nand U6023 (N_6023,In_2449,In_625);
nor U6024 (N_6024,In_1174,In_1339);
and U6025 (N_6025,In_1647,In_1504);
and U6026 (N_6026,In_269,In_355);
nor U6027 (N_6027,In_524,In_456);
nand U6028 (N_6028,In_786,In_511);
nor U6029 (N_6029,In_966,In_2013);
xor U6030 (N_6030,In_1553,In_2144);
and U6031 (N_6031,In_754,In_173);
or U6032 (N_6032,In_2242,In_315);
or U6033 (N_6033,In_2146,In_849);
xnor U6034 (N_6034,In_212,In_1813);
and U6035 (N_6035,In_1555,In_2346);
or U6036 (N_6036,In_1750,In_1688);
or U6037 (N_6037,In_2445,In_2400);
or U6038 (N_6038,In_1845,In_618);
or U6039 (N_6039,In_2388,In_2024);
or U6040 (N_6040,In_1467,In_1743);
xor U6041 (N_6041,In_544,In_1873);
xnor U6042 (N_6042,In_1043,In_1929);
nand U6043 (N_6043,In_981,In_680);
nor U6044 (N_6044,In_2497,In_807);
or U6045 (N_6045,In_600,In_1839);
nand U6046 (N_6046,In_1751,In_563);
nor U6047 (N_6047,In_251,In_122);
nor U6048 (N_6048,In_1008,In_699);
or U6049 (N_6049,In_1995,In_524);
nand U6050 (N_6050,In_1159,In_965);
nor U6051 (N_6051,In_1806,In_18);
and U6052 (N_6052,In_661,In_2448);
and U6053 (N_6053,In_1918,In_499);
or U6054 (N_6054,In_1842,In_219);
nor U6055 (N_6055,In_264,In_1048);
nor U6056 (N_6056,In_2038,In_2050);
or U6057 (N_6057,In_1839,In_1080);
and U6058 (N_6058,In_963,In_1950);
or U6059 (N_6059,In_1915,In_2173);
nand U6060 (N_6060,In_692,In_1360);
nand U6061 (N_6061,In_665,In_1476);
or U6062 (N_6062,In_1225,In_722);
xor U6063 (N_6063,In_1990,In_1882);
nand U6064 (N_6064,In_1953,In_961);
and U6065 (N_6065,In_1595,In_2063);
nor U6066 (N_6066,In_2334,In_524);
nor U6067 (N_6067,In_997,In_503);
nor U6068 (N_6068,In_243,In_30);
xor U6069 (N_6069,In_970,In_1767);
nand U6070 (N_6070,In_553,In_629);
nand U6071 (N_6071,In_166,In_406);
nor U6072 (N_6072,In_1902,In_2022);
nor U6073 (N_6073,In_413,In_2493);
xor U6074 (N_6074,In_2486,In_905);
nor U6075 (N_6075,In_651,In_1426);
nand U6076 (N_6076,In_423,In_1882);
nor U6077 (N_6077,In_2142,In_1847);
nand U6078 (N_6078,In_2258,In_752);
nand U6079 (N_6079,In_1562,In_1781);
or U6080 (N_6080,In_1301,In_1008);
and U6081 (N_6081,In_2150,In_387);
or U6082 (N_6082,In_2169,In_2096);
and U6083 (N_6083,In_781,In_484);
nor U6084 (N_6084,In_2100,In_1738);
or U6085 (N_6085,In_1921,In_1383);
or U6086 (N_6086,In_1491,In_1279);
nor U6087 (N_6087,In_2184,In_1314);
and U6088 (N_6088,In_209,In_818);
nor U6089 (N_6089,In_491,In_1617);
nand U6090 (N_6090,In_2326,In_345);
or U6091 (N_6091,In_1206,In_1279);
xor U6092 (N_6092,In_724,In_2319);
xor U6093 (N_6093,In_1681,In_995);
nor U6094 (N_6094,In_341,In_588);
and U6095 (N_6095,In_1699,In_801);
nand U6096 (N_6096,In_1551,In_1760);
or U6097 (N_6097,In_226,In_2125);
nand U6098 (N_6098,In_2260,In_1112);
nor U6099 (N_6099,In_1034,In_506);
or U6100 (N_6100,In_1920,In_2442);
and U6101 (N_6101,In_143,In_1922);
nand U6102 (N_6102,In_436,In_1295);
nor U6103 (N_6103,In_2093,In_1744);
nand U6104 (N_6104,In_918,In_1260);
nand U6105 (N_6105,In_804,In_1376);
nand U6106 (N_6106,In_947,In_1535);
and U6107 (N_6107,In_176,In_260);
xor U6108 (N_6108,In_2319,In_703);
xor U6109 (N_6109,In_2383,In_2108);
or U6110 (N_6110,In_1272,In_2381);
nor U6111 (N_6111,In_38,In_1460);
nand U6112 (N_6112,In_734,In_1321);
nand U6113 (N_6113,In_2403,In_569);
and U6114 (N_6114,In_1928,In_2022);
or U6115 (N_6115,In_552,In_976);
nor U6116 (N_6116,In_1766,In_1747);
and U6117 (N_6117,In_1531,In_1133);
xnor U6118 (N_6118,In_1455,In_1938);
or U6119 (N_6119,In_453,In_1016);
nand U6120 (N_6120,In_1609,In_920);
xor U6121 (N_6121,In_497,In_477);
or U6122 (N_6122,In_604,In_2274);
xnor U6123 (N_6123,In_968,In_1484);
or U6124 (N_6124,In_820,In_992);
and U6125 (N_6125,In_24,In_1232);
nor U6126 (N_6126,In_328,In_742);
xnor U6127 (N_6127,In_89,In_879);
and U6128 (N_6128,In_1585,In_612);
xor U6129 (N_6129,In_1524,In_1059);
nand U6130 (N_6130,In_359,In_1014);
nor U6131 (N_6131,In_830,In_2372);
and U6132 (N_6132,In_494,In_728);
or U6133 (N_6133,In_1641,In_1386);
xor U6134 (N_6134,In_17,In_173);
or U6135 (N_6135,In_776,In_1908);
and U6136 (N_6136,In_1178,In_421);
and U6137 (N_6137,In_2255,In_361);
and U6138 (N_6138,In_1711,In_1345);
xnor U6139 (N_6139,In_2429,In_1531);
and U6140 (N_6140,In_1410,In_2279);
xnor U6141 (N_6141,In_2318,In_140);
xnor U6142 (N_6142,In_1930,In_1666);
xor U6143 (N_6143,In_36,In_1940);
nand U6144 (N_6144,In_572,In_1852);
xor U6145 (N_6145,In_2300,In_1073);
xnor U6146 (N_6146,In_1659,In_822);
or U6147 (N_6147,In_901,In_1268);
and U6148 (N_6148,In_2042,In_460);
nand U6149 (N_6149,In_1194,In_2211);
nand U6150 (N_6150,In_908,In_894);
and U6151 (N_6151,In_1970,In_1077);
nand U6152 (N_6152,In_2183,In_2215);
nor U6153 (N_6153,In_2002,In_2082);
xnor U6154 (N_6154,In_2428,In_1123);
or U6155 (N_6155,In_1003,In_115);
nand U6156 (N_6156,In_477,In_1449);
nand U6157 (N_6157,In_2002,In_1293);
xor U6158 (N_6158,In_1841,In_209);
xor U6159 (N_6159,In_1297,In_1537);
or U6160 (N_6160,In_2251,In_310);
and U6161 (N_6161,In_2086,In_551);
and U6162 (N_6162,In_1404,In_884);
or U6163 (N_6163,In_1443,In_1947);
and U6164 (N_6164,In_71,In_2408);
or U6165 (N_6165,In_1264,In_749);
and U6166 (N_6166,In_1789,In_361);
xor U6167 (N_6167,In_869,In_596);
xor U6168 (N_6168,In_725,In_2371);
and U6169 (N_6169,In_1782,In_2205);
nor U6170 (N_6170,In_2249,In_1865);
nor U6171 (N_6171,In_2003,In_2399);
nand U6172 (N_6172,In_1414,In_1645);
nand U6173 (N_6173,In_283,In_124);
nor U6174 (N_6174,In_897,In_1909);
nor U6175 (N_6175,In_2462,In_968);
nand U6176 (N_6176,In_265,In_98);
and U6177 (N_6177,In_246,In_2481);
xnor U6178 (N_6178,In_1171,In_2445);
nand U6179 (N_6179,In_1222,In_2427);
nor U6180 (N_6180,In_283,In_2106);
and U6181 (N_6181,In_1873,In_2127);
nor U6182 (N_6182,In_1532,In_2279);
xnor U6183 (N_6183,In_2430,In_2147);
nand U6184 (N_6184,In_1409,In_2103);
nor U6185 (N_6185,In_252,In_267);
or U6186 (N_6186,In_1288,In_2352);
or U6187 (N_6187,In_212,In_2084);
nor U6188 (N_6188,In_865,In_2119);
nand U6189 (N_6189,In_499,In_1150);
nand U6190 (N_6190,In_1226,In_1448);
xor U6191 (N_6191,In_472,In_1355);
nand U6192 (N_6192,In_1170,In_1925);
or U6193 (N_6193,In_531,In_1602);
nand U6194 (N_6194,In_2291,In_820);
nor U6195 (N_6195,In_390,In_1378);
and U6196 (N_6196,In_1126,In_476);
nor U6197 (N_6197,In_96,In_2111);
xor U6198 (N_6198,In_210,In_1748);
or U6199 (N_6199,In_972,In_1492);
nor U6200 (N_6200,In_2454,In_2342);
nor U6201 (N_6201,In_55,In_1181);
or U6202 (N_6202,In_2411,In_838);
nor U6203 (N_6203,In_1099,In_1484);
or U6204 (N_6204,In_966,In_766);
nor U6205 (N_6205,In_2361,In_745);
xor U6206 (N_6206,In_108,In_1314);
nor U6207 (N_6207,In_2290,In_119);
nor U6208 (N_6208,In_2154,In_335);
or U6209 (N_6209,In_2204,In_1371);
nor U6210 (N_6210,In_1777,In_761);
and U6211 (N_6211,In_1592,In_785);
nor U6212 (N_6212,In_541,In_1547);
and U6213 (N_6213,In_990,In_571);
nand U6214 (N_6214,In_833,In_2345);
and U6215 (N_6215,In_2228,In_1898);
and U6216 (N_6216,In_1059,In_2268);
nor U6217 (N_6217,In_1755,In_2107);
and U6218 (N_6218,In_597,In_77);
and U6219 (N_6219,In_1590,In_866);
nor U6220 (N_6220,In_286,In_102);
or U6221 (N_6221,In_1875,In_1341);
nor U6222 (N_6222,In_898,In_1033);
xnor U6223 (N_6223,In_1566,In_16);
nand U6224 (N_6224,In_1501,In_2171);
or U6225 (N_6225,In_719,In_2340);
and U6226 (N_6226,In_2078,In_699);
nor U6227 (N_6227,In_452,In_518);
and U6228 (N_6228,In_270,In_21);
xor U6229 (N_6229,In_775,In_2246);
or U6230 (N_6230,In_500,In_383);
nand U6231 (N_6231,In_1074,In_1463);
xor U6232 (N_6232,In_1997,In_2340);
nand U6233 (N_6233,In_285,In_77);
nand U6234 (N_6234,In_16,In_422);
or U6235 (N_6235,In_2113,In_1286);
or U6236 (N_6236,In_1985,In_1424);
and U6237 (N_6237,In_1708,In_2137);
and U6238 (N_6238,In_1647,In_812);
or U6239 (N_6239,In_299,In_1903);
nor U6240 (N_6240,In_1266,In_1049);
xnor U6241 (N_6241,In_932,In_1923);
nand U6242 (N_6242,In_1468,In_7);
nand U6243 (N_6243,In_1072,In_496);
and U6244 (N_6244,In_1336,In_2372);
xnor U6245 (N_6245,In_2016,In_66);
and U6246 (N_6246,In_895,In_2108);
or U6247 (N_6247,In_1873,In_1091);
xnor U6248 (N_6248,In_1883,In_806);
xor U6249 (N_6249,In_2439,In_1383);
nand U6250 (N_6250,N_2419,N_957);
or U6251 (N_6251,N_2850,N_4936);
or U6252 (N_6252,N_4448,N_5244);
or U6253 (N_6253,N_735,N_2004);
and U6254 (N_6254,N_5723,N_881);
xor U6255 (N_6255,N_5786,N_2692);
xor U6256 (N_6256,N_1282,N_1538);
nor U6257 (N_6257,N_5222,N_534);
and U6258 (N_6258,N_1874,N_1217);
xnor U6259 (N_6259,N_4264,N_619);
or U6260 (N_6260,N_3363,N_4668);
nand U6261 (N_6261,N_5151,N_3462);
and U6262 (N_6262,N_759,N_213);
xor U6263 (N_6263,N_4380,N_3421);
nor U6264 (N_6264,N_4968,N_1916);
and U6265 (N_6265,N_1494,N_3960);
or U6266 (N_6266,N_5612,N_2813);
xor U6267 (N_6267,N_1179,N_1246);
and U6268 (N_6268,N_2729,N_771);
or U6269 (N_6269,N_2477,N_5897);
xnor U6270 (N_6270,N_2639,N_5141);
and U6271 (N_6271,N_318,N_1511);
xor U6272 (N_6272,N_562,N_991);
xor U6273 (N_6273,N_2833,N_3236);
or U6274 (N_6274,N_1257,N_5026);
or U6275 (N_6275,N_5339,N_6037);
xnor U6276 (N_6276,N_5662,N_4760);
or U6277 (N_6277,N_5163,N_414);
nor U6278 (N_6278,N_6129,N_1161);
and U6279 (N_6279,N_1480,N_3802);
nand U6280 (N_6280,N_196,N_937);
or U6281 (N_6281,N_4869,N_3476);
xnor U6282 (N_6282,N_2698,N_5099);
or U6283 (N_6283,N_5461,N_5988);
and U6284 (N_6284,N_5443,N_6202);
nand U6285 (N_6285,N_4884,N_3153);
xnor U6286 (N_6286,N_4171,N_2634);
nor U6287 (N_6287,N_2664,N_4710);
xnor U6288 (N_6288,N_2459,N_512);
and U6289 (N_6289,N_3357,N_1514);
nor U6290 (N_6290,N_751,N_5186);
xor U6291 (N_6291,N_337,N_4081);
nor U6292 (N_6292,N_5715,N_3339);
or U6293 (N_6293,N_4323,N_3602);
and U6294 (N_6294,N_967,N_1771);
xor U6295 (N_6295,N_5757,N_1615);
and U6296 (N_6296,N_5279,N_5420);
nor U6297 (N_6297,N_2542,N_4395);
or U6298 (N_6298,N_2082,N_3195);
nand U6299 (N_6299,N_2605,N_6091);
or U6300 (N_6300,N_2307,N_546);
or U6301 (N_6301,N_4570,N_335);
nor U6302 (N_6302,N_1095,N_6025);
or U6303 (N_6303,N_5345,N_1327);
nor U6304 (N_6304,N_1387,N_3453);
and U6305 (N_6305,N_1752,N_2925);
xor U6306 (N_6306,N_378,N_2481);
or U6307 (N_6307,N_2952,N_648);
and U6308 (N_6308,N_2855,N_3582);
xor U6309 (N_6309,N_679,N_3310);
nand U6310 (N_6310,N_1507,N_3758);
xor U6311 (N_6311,N_3924,N_3514);
or U6312 (N_6312,N_1144,N_3850);
nor U6313 (N_6313,N_3832,N_5908);
or U6314 (N_6314,N_4466,N_68);
and U6315 (N_6315,N_3835,N_2876);
nor U6316 (N_6316,N_906,N_2453);
xnor U6317 (N_6317,N_30,N_4990);
xnor U6318 (N_6318,N_3724,N_3364);
nor U6319 (N_6319,N_670,N_260);
nand U6320 (N_6320,N_899,N_83);
or U6321 (N_6321,N_4140,N_4182);
nor U6322 (N_6322,N_4533,N_998);
or U6323 (N_6323,N_1982,N_4090);
and U6324 (N_6324,N_1026,N_1961);
and U6325 (N_6325,N_6046,N_1096);
or U6326 (N_6326,N_531,N_3399);
nand U6327 (N_6327,N_5840,N_1590);
or U6328 (N_6328,N_2073,N_980);
and U6329 (N_6329,N_3171,N_3134);
or U6330 (N_6330,N_2878,N_601);
or U6331 (N_6331,N_1394,N_2918);
nor U6332 (N_6332,N_2875,N_935);
and U6333 (N_6333,N_2900,N_3435);
nor U6334 (N_6334,N_2144,N_5935);
and U6335 (N_6335,N_5713,N_1067);
or U6336 (N_6336,N_270,N_4126);
xnor U6337 (N_6337,N_3212,N_4260);
or U6338 (N_6338,N_6128,N_3854);
xor U6339 (N_6339,N_6130,N_4746);
xnor U6340 (N_6340,N_2044,N_1234);
xnor U6341 (N_6341,N_1287,N_3772);
xor U6342 (N_6342,N_5714,N_3270);
xnor U6343 (N_6343,N_4941,N_3899);
or U6344 (N_6344,N_1662,N_1586);
xnor U6345 (N_6345,N_234,N_5783);
nand U6346 (N_6346,N_2815,N_246);
and U6347 (N_6347,N_2390,N_668);
nand U6348 (N_6348,N_5301,N_3788);
or U6349 (N_6349,N_1636,N_1297);
and U6350 (N_6350,N_6189,N_1952);
or U6351 (N_6351,N_683,N_2566);
and U6352 (N_6352,N_3222,N_482);
xor U6353 (N_6353,N_3331,N_770);
xnor U6354 (N_6354,N_3573,N_2725);
nor U6355 (N_6355,N_133,N_359);
nand U6356 (N_6356,N_457,N_3035);
xnor U6357 (N_6357,N_5242,N_4994);
nor U6358 (N_6358,N_1675,N_2688);
xor U6359 (N_6359,N_2425,N_1539);
nand U6360 (N_6360,N_2197,N_1105);
nand U6361 (N_6361,N_3709,N_760);
nor U6362 (N_6362,N_1948,N_1187);
and U6363 (N_6363,N_2146,N_1435);
nand U6364 (N_6364,N_6170,N_1657);
nand U6365 (N_6365,N_2801,N_5766);
and U6366 (N_6366,N_5216,N_3137);
nand U6367 (N_6367,N_2030,N_3030);
nand U6368 (N_6368,N_5109,N_186);
nor U6369 (N_6369,N_388,N_5860);
nor U6370 (N_6370,N_1763,N_3671);
nand U6371 (N_6371,N_694,N_3235);
nor U6372 (N_6372,N_4714,N_3563);
xnor U6373 (N_6373,N_4978,N_5655);
xor U6374 (N_6374,N_4161,N_2136);
and U6375 (N_6375,N_3086,N_2402);
nor U6376 (N_6376,N_91,N_2284);
or U6377 (N_6377,N_983,N_3087);
xnor U6378 (N_6378,N_324,N_1998);
and U6379 (N_6379,N_680,N_5588);
or U6380 (N_6380,N_5843,N_4834);
or U6381 (N_6381,N_5466,N_4654);
nand U6382 (N_6382,N_1608,N_1888);
nor U6383 (N_6383,N_6214,N_664);
nor U6384 (N_6384,N_2189,N_530);
and U6385 (N_6385,N_6087,N_1019);
and U6386 (N_6386,N_2223,N_916);
and U6387 (N_6387,N_1614,N_5075);
xnor U6388 (N_6388,N_1623,N_154);
or U6389 (N_6389,N_2192,N_2145);
nor U6390 (N_6390,N_4987,N_69);
and U6391 (N_6391,N_2661,N_2973);
or U6392 (N_6392,N_3711,N_6161);
nor U6393 (N_6393,N_3938,N_2831);
and U6394 (N_6394,N_2045,N_5862);
nand U6395 (N_6395,N_4179,N_349);
xor U6396 (N_6396,N_2507,N_112);
or U6397 (N_6397,N_4275,N_1534);
xor U6398 (N_6398,N_3538,N_5215);
nand U6399 (N_6399,N_3750,N_1001);
xor U6400 (N_6400,N_277,N_1053);
and U6401 (N_6401,N_5039,N_1783);
and U6402 (N_6402,N_4369,N_3604);
or U6403 (N_6403,N_1780,N_3038);
xnor U6404 (N_6404,N_4979,N_4751);
xnor U6405 (N_6405,N_3775,N_4461);
or U6406 (N_6406,N_387,N_254);
nor U6407 (N_6407,N_3676,N_779);
or U6408 (N_6408,N_5219,N_1685);
nor U6409 (N_6409,N_5097,N_4669);
nand U6410 (N_6410,N_3877,N_3239);
or U6411 (N_6411,N_459,N_3044);
xor U6412 (N_6412,N_5023,N_2247);
nor U6413 (N_6413,N_4356,N_6104);
xnor U6414 (N_6414,N_2093,N_3168);
or U6415 (N_6415,N_3401,N_3492);
nor U6416 (N_6416,N_2074,N_4449);
or U6417 (N_6417,N_127,N_4358);
or U6418 (N_6418,N_4084,N_369);
or U6419 (N_6419,N_1581,N_5237);
and U6420 (N_6420,N_56,N_4089);
xor U6421 (N_6421,N_2000,N_4837);
xor U6422 (N_6422,N_4201,N_361);
or U6423 (N_6423,N_1092,N_5596);
and U6424 (N_6424,N_2777,N_2956);
xor U6425 (N_6425,N_1183,N_542);
xor U6426 (N_6426,N_1410,N_2274);
nor U6427 (N_6427,N_5487,N_4057);
xnor U6428 (N_6428,N_1812,N_2894);
and U6429 (N_6429,N_3360,N_4619);
and U6430 (N_6430,N_2779,N_2613);
nand U6431 (N_6431,N_4243,N_4687);
and U6432 (N_6432,N_1547,N_237);
xor U6433 (N_6433,N_1602,N_5368);
nor U6434 (N_6434,N_3585,N_6102);
xnor U6435 (N_6435,N_4145,N_5498);
nand U6436 (N_6436,N_3342,N_2685);
and U6437 (N_6437,N_1071,N_3062);
nor U6438 (N_6438,N_3697,N_4276);
xnor U6439 (N_6439,N_4332,N_2844);
xor U6440 (N_6440,N_820,N_3741);
nand U6441 (N_6441,N_926,N_5058);
nor U6442 (N_6442,N_2965,N_1831);
xnor U6443 (N_6443,N_1641,N_2842);
nor U6444 (N_6444,N_556,N_5479);
xnor U6445 (N_6445,N_5797,N_4068);
or U6446 (N_6446,N_189,N_1673);
and U6447 (N_6447,N_5974,N_2428);
or U6448 (N_6448,N_2335,N_1157);
and U6449 (N_6449,N_3547,N_4956);
nand U6450 (N_6450,N_195,N_1809);
nand U6451 (N_6451,N_5520,N_1726);
xnor U6452 (N_6452,N_936,N_6139);
or U6453 (N_6453,N_624,N_5040);
nor U6454 (N_6454,N_5327,N_351);
or U6455 (N_6455,N_1400,N_2187);
and U6456 (N_6456,N_1192,N_2058);
xnor U6457 (N_6457,N_2746,N_1527);
or U6458 (N_6458,N_1566,N_3747);
and U6459 (N_6459,N_2487,N_190);
nand U6460 (N_6460,N_4388,N_1296);
nor U6461 (N_6461,N_1665,N_1989);
nor U6462 (N_6462,N_5235,N_4190);
and U6463 (N_6463,N_1865,N_2737);
or U6464 (N_6464,N_2961,N_3792);
nor U6465 (N_6465,N_5440,N_1362);
and U6466 (N_6466,N_423,N_5674);
nand U6467 (N_6467,N_2429,N_5232);
xor U6468 (N_6468,N_232,N_1174);
nor U6469 (N_6469,N_1194,N_5730);
nor U6470 (N_6470,N_4665,N_5119);
xnor U6471 (N_6471,N_4697,N_1344);
or U6472 (N_6472,N_824,N_2728);
nor U6473 (N_6473,N_2277,N_1462);
and U6474 (N_6474,N_876,N_3945);
nand U6475 (N_6475,N_2349,N_3033);
xnor U6476 (N_6476,N_1986,N_4125);
nand U6477 (N_6477,N_3932,N_1895);
nor U6478 (N_6478,N_3480,N_1628);
xnor U6479 (N_6479,N_2934,N_1571);
and U6480 (N_6480,N_5115,N_5229);
or U6481 (N_6481,N_5250,N_2577);
nor U6482 (N_6482,N_2440,N_2549);
nand U6483 (N_6483,N_170,N_5568);
nand U6484 (N_6484,N_2430,N_3147);
or U6485 (N_6485,N_5424,N_4390);
or U6486 (N_6486,N_104,N_1508);
nand U6487 (N_6487,N_910,N_4952);
xnor U6488 (N_6488,N_4902,N_3415);
nor U6489 (N_6489,N_5589,N_3594);
nand U6490 (N_6490,N_1184,N_5855);
or U6491 (N_6491,N_501,N_4009);
or U6492 (N_6492,N_2214,N_442);
nor U6493 (N_6493,N_6133,N_333);
and U6494 (N_6494,N_1559,N_4501);
xnor U6495 (N_6495,N_3943,N_2932);
nor U6496 (N_6496,N_6076,N_5310);
or U6497 (N_6497,N_2867,N_2422);
or U6498 (N_6498,N_275,N_5519);
nand U6499 (N_6499,N_1149,N_1464);
nand U6500 (N_6500,N_3979,N_5885);
nand U6501 (N_6501,N_2881,N_3181);
nor U6502 (N_6502,N_2583,N_5972);
xor U6503 (N_6503,N_3733,N_5298);
and U6504 (N_6504,N_4823,N_959);
xnor U6505 (N_6505,N_390,N_1080);
nand U6506 (N_6506,N_3634,N_4895);
xor U6507 (N_6507,N_3882,N_2745);
or U6508 (N_6508,N_5156,N_4546);
nor U6509 (N_6509,N_1625,N_430);
and U6510 (N_6510,N_3528,N_2805);
xnor U6511 (N_6511,N_996,N_5257);
and U6512 (N_6512,N_5426,N_3474);
nor U6513 (N_6513,N_979,N_2470);
or U6514 (N_6514,N_5936,N_6230);
xor U6515 (N_6515,N_4860,N_4228);
and U6516 (N_6516,N_1438,N_2946);
and U6517 (N_6517,N_3897,N_5140);
nand U6518 (N_6518,N_426,N_904);
nor U6519 (N_6519,N_75,N_4176);
and U6520 (N_6520,N_1553,N_4139);
nor U6521 (N_6521,N_3626,N_4119);
xor U6522 (N_6522,N_5388,N_1849);
and U6523 (N_6523,N_746,N_1315);
and U6524 (N_6524,N_4883,N_1512);
and U6525 (N_6525,N_1687,N_2165);
nand U6526 (N_6526,N_3083,N_2753);
nor U6527 (N_6527,N_1843,N_2076);
nand U6528 (N_6528,N_1899,N_4970);
nand U6529 (N_6529,N_1801,N_1690);
nor U6530 (N_6530,N_4118,N_3145);
and U6531 (N_6531,N_1802,N_174);
and U6532 (N_6532,N_3196,N_1521);
nor U6533 (N_6533,N_1627,N_4564);
nor U6534 (N_6534,N_702,N_2739);
or U6535 (N_6535,N_51,N_5954);
nand U6536 (N_6536,N_3131,N_852);
xor U6537 (N_6537,N_2062,N_2523);
nor U6538 (N_6538,N_2863,N_3478);
nand U6539 (N_6539,N_2399,N_4728);
xnor U6540 (N_6540,N_6233,N_1087);
nand U6541 (N_6541,N_3632,N_224);
nor U6542 (N_6542,N_1269,N_607);
or U6543 (N_6543,N_5819,N_265);
or U6544 (N_6544,N_3531,N_3746);
and U6545 (N_6545,N_3079,N_4498);
xnor U6546 (N_6546,N_3851,N_4023);
nor U6547 (N_6547,N_544,N_5325);
nor U6548 (N_6548,N_3276,N_3163);
and U6549 (N_6549,N_1249,N_3948);
or U6550 (N_6550,N_5861,N_3905);
xnor U6551 (N_6551,N_3922,N_2304);
nand U6552 (N_6552,N_541,N_5690);
or U6553 (N_6553,N_2511,N_5491);
or U6554 (N_6554,N_1607,N_4378);
and U6555 (N_6555,N_1500,N_373);
nor U6556 (N_6556,N_866,N_1205);
xor U6557 (N_6557,N_6231,N_5642);
nor U6558 (N_6558,N_4286,N_6034);
and U6559 (N_6559,N_784,N_2173);
and U6560 (N_6560,N_5403,N_5961);
and U6561 (N_6561,N_5335,N_6144);
nand U6562 (N_6562,N_6010,N_2079);
nand U6563 (N_6563,N_1000,N_159);
and U6564 (N_6564,N_3779,N_4166);
nand U6565 (N_6565,N_5656,N_3810);
nor U6566 (N_6566,N_4097,N_235);
and U6567 (N_6567,N_804,N_131);
nand U6568 (N_6568,N_5727,N_3328);
xnor U6569 (N_6569,N_5210,N_5285);
nor U6570 (N_6570,N_4039,N_1537);
nor U6571 (N_6571,N_215,N_4284);
xnor U6572 (N_6572,N_5636,N_4165);
nor U6573 (N_6573,N_3853,N_1397);
or U6574 (N_6574,N_4329,N_4297);
and U6575 (N_6575,N_2704,N_2107);
and U6576 (N_6576,N_5469,N_1902);
nand U6577 (N_6577,N_3368,N_4984);
xor U6578 (N_6578,N_1453,N_5680);
and U6579 (N_6579,N_1746,N_5181);
xor U6580 (N_6580,N_2614,N_1474);
or U6581 (N_6581,N_4447,N_3645);
xnor U6582 (N_6582,N_4861,N_6106);
nor U6583 (N_6583,N_840,N_3156);
or U6584 (N_6584,N_2023,N_5201);
xor U6585 (N_6585,N_2412,N_2182);
or U6586 (N_6586,N_4818,N_473);
xnor U6587 (N_6587,N_288,N_720);
nor U6588 (N_6588,N_212,N_2160);
or U6589 (N_6589,N_615,N_3094);
or U6590 (N_6590,N_3097,N_4105);
or U6591 (N_6591,N_3283,N_1492);
nand U6592 (N_6592,N_4515,N_545);
or U6593 (N_6593,N_4168,N_300);
nor U6594 (N_6594,N_2503,N_660);
and U6595 (N_6595,N_4472,N_6248);
xnor U6596 (N_6596,N_3801,N_3683);
nand U6597 (N_6597,N_3844,N_6093);
or U6598 (N_6598,N_3429,N_5079);
or U6599 (N_6599,N_1093,N_995);
and U6600 (N_6600,N_1245,N_2967);
or U6601 (N_6601,N_5386,N_4602);
and U6602 (N_6602,N_2858,N_5299);
nor U6603 (N_6603,N_3170,N_2959);
and U6604 (N_6604,N_126,N_2366);
and U6605 (N_6605,N_4905,N_5598);
and U6606 (N_6606,N_4368,N_3680);
and U6607 (N_6607,N_1178,N_2015);
xnor U6608 (N_6608,N_6049,N_4942);
or U6609 (N_6609,N_209,N_3228);
or U6610 (N_6610,N_393,N_5551);
nor U6611 (N_6611,N_1248,N_102);
and U6612 (N_6612,N_1484,N_1025);
nor U6613 (N_6613,N_4010,N_78);
and U6614 (N_6614,N_2830,N_4565);
or U6615 (N_6615,N_1782,N_3976);
and U6616 (N_6616,N_5130,N_2052);
nor U6617 (N_6617,N_2536,N_5146);
or U6618 (N_6618,N_263,N_1635);
and U6619 (N_6619,N_3858,N_732);
xor U6620 (N_6620,N_5619,N_2373);
and U6621 (N_6621,N_1437,N_3815);
xor U6622 (N_6622,N_1414,N_486);
nand U6623 (N_6623,N_3544,N_441);
xnor U6624 (N_6624,N_1605,N_5166);
xor U6625 (N_6625,N_4212,N_2191);
or U6626 (N_6626,N_5184,N_5107);
and U6627 (N_6627,N_1263,N_3609);
nor U6628 (N_6628,N_5004,N_5595);
xor U6629 (N_6629,N_4328,N_5007);
or U6630 (N_6630,N_5068,N_5764);
and U6631 (N_6631,N_3172,N_383);
or U6632 (N_6632,N_281,N_2267);
xnor U6633 (N_6633,N_2190,N_4012);
nand U6634 (N_6634,N_5530,N_6113);
xor U6635 (N_6635,N_157,N_1969);
and U6636 (N_6636,N_1363,N_192);
xor U6637 (N_6637,N_3365,N_1044);
nor U6638 (N_6638,N_3424,N_5615);
or U6639 (N_6639,N_5353,N_2841);
nand U6640 (N_6640,N_5472,N_201);
nand U6641 (N_6641,N_1243,N_3417);
nor U6642 (N_6642,N_6220,N_460);
and U6643 (N_6643,N_1117,N_5775);
xnor U6644 (N_6644,N_4918,N_5822);
xnor U6645 (N_6645,N_6016,N_3606);
and U6646 (N_6646,N_4406,N_219);
and U6647 (N_6647,N_3329,N_5883);
xnor U6648 (N_6648,N_4024,N_3866);
or U6649 (N_6649,N_4028,N_2572);
or U6650 (N_6650,N_4571,N_462);
or U6651 (N_6651,N_2749,N_5895);
nor U6652 (N_6652,N_183,N_834);
and U6653 (N_6653,N_1284,N_5916);
and U6654 (N_6654,N_4926,N_844);
and U6655 (N_6655,N_164,N_2468);
and U6656 (N_6656,N_2683,N_3341);
and U6657 (N_6657,N_1398,N_4739);
xor U6658 (N_6658,N_1086,N_2380);
xnor U6659 (N_6659,N_1038,N_2393);
nand U6660 (N_6660,N_1762,N_4185);
nor U6661 (N_6661,N_2620,N_5580);
or U6662 (N_6662,N_5042,N_4399);
or U6663 (N_6663,N_5652,N_2090);
nand U6664 (N_6664,N_3440,N_1409);
nand U6665 (N_6665,N_2703,N_2126);
xnor U6666 (N_6666,N_6239,N_650);
or U6667 (N_6667,N_1382,N_53);
nor U6668 (N_6668,N_5422,N_1108);
nand U6669 (N_6669,N_3317,N_2993);
or U6670 (N_6670,N_4698,N_1046);
nor U6671 (N_6671,N_3846,N_1562);
xnor U6672 (N_6672,N_4340,N_2303);
or U6673 (N_6673,N_4433,N_4988);
nor U6674 (N_6674,N_3005,N_5060);
xnor U6675 (N_6675,N_941,N_3787);
or U6676 (N_6676,N_4704,N_5625);
nor U6677 (N_6677,N_1525,N_2239);
and U6678 (N_6678,N_242,N_2242);
xor U6679 (N_6679,N_4281,N_3358);
and U6680 (N_6680,N_3126,N_4662);
nor U6681 (N_6681,N_3238,N_3583);
and U6682 (N_6682,N_3860,N_6115);
xor U6683 (N_6683,N_790,N_4705);
nand U6684 (N_6684,N_3845,N_141);
and U6685 (N_6685,N_2883,N_5952);
nor U6686 (N_6686,N_3588,N_758);
nand U6687 (N_6687,N_3613,N_4341);
and U6688 (N_6688,N_107,N_1923);
and U6689 (N_6689,N_569,N_1360);
nor U6690 (N_6690,N_5356,N_649);
nor U6691 (N_6691,N_1262,N_4349);
nand U6692 (N_6692,N_1754,N_437);
nor U6693 (N_6693,N_166,N_843);
xor U6694 (N_6694,N_4436,N_6185);
nor U6695 (N_6695,N_778,N_1709);
nand U6696 (N_6696,N_4977,N_2760);
and U6697 (N_6697,N_940,N_4856);
nor U6698 (N_6698,N_3425,N_5884);
and U6699 (N_6699,N_1227,N_792);
and U6700 (N_6700,N_5372,N_3121);
nor U6701 (N_6701,N_2035,N_3678);
and U6702 (N_6702,N_5923,N_1036);
xor U6703 (N_6703,N_4736,N_3279);
nand U6704 (N_6704,N_1370,N_450);
nor U6705 (N_6705,N_5521,N_6172);
xor U6706 (N_6706,N_492,N_6216);
nor U6707 (N_6707,N_1676,N_5581);
nand U6708 (N_6708,N_2155,N_1721);
nand U6709 (N_6709,N_791,N_6029);
and U6710 (N_6710,N_2263,N_5332);
xnor U6711 (N_6711,N_2465,N_5560);
or U6712 (N_6712,N_749,N_833);
nand U6713 (N_6713,N_4469,N_3157);
nor U6714 (N_6714,N_2457,N_1153);
or U6715 (N_6715,N_6234,N_3495);
and U6716 (N_6716,N_2313,N_3702);
or U6717 (N_6717,N_2852,N_1633);
nand U6718 (N_6718,N_1114,N_5864);
xor U6719 (N_6719,N_3112,N_5261);
nand U6720 (N_6720,N_4732,N_1666);
xor U6721 (N_6721,N_2942,N_475);
or U6722 (N_6722,N_3370,N_1548);
or U6723 (N_6723,N_6116,N_3513);
or U6724 (N_6724,N_2874,N_608);
or U6725 (N_6725,N_2928,N_5437);
or U6726 (N_6726,N_1416,N_823);
and U6727 (N_6727,N_1867,N_3655);
nand U6728 (N_6728,N_2645,N_1293);
xor U6729 (N_6729,N_2843,N_2835);
and U6730 (N_6730,N_1079,N_5901);
or U6731 (N_6731,N_4370,N_575);
or U6732 (N_6732,N_1037,N_1112);
and U6733 (N_6733,N_5430,N_2362);
nor U6734 (N_6734,N_4239,N_6074);
nand U6735 (N_6735,N_3596,N_5925);
nor U6736 (N_6736,N_576,N_4867);
or U6737 (N_6737,N_3891,N_4077);
nor U6738 (N_6738,N_933,N_695);
xnor U6739 (N_6739,N_3493,N_231);
and U6740 (N_6740,N_2348,N_2570);
nor U6741 (N_6741,N_5116,N_2418);
xnor U6742 (N_6742,N_4876,N_200);
nor U6743 (N_6743,N_603,N_5792);
and U6744 (N_6744,N_2127,N_5648);
nor U6745 (N_6745,N_3612,N_1835);
or U6746 (N_6746,N_3773,N_273);
xor U6747 (N_6747,N_3307,N_2772);
and U6748 (N_6748,N_3359,N_2195);
and U6749 (N_6749,N_4808,N_5022);
nand U6750 (N_6750,N_954,N_2217);
and U6751 (N_6751,N_1172,N_5164);
xor U6752 (N_6752,N_1714,N_2715);
xor U6753 (N_6753,N_832,N_1704);
nand U6754 (N_6754,N_3862,N_1354);
and U6755 (N_6755,N_4361,N_5756);
and U6756 (N_6756,N_3334,N_2383);
and U6757 (N_6757,N_4133,N_1945);
and U6758 (N_6758,N_3377,N_2101);
nor U6759 (N_6759,N_3049,N_1335);
and U6760 (N_6760,N_4699,N_2764);
nand U6761 (N_6761,N_2085,N_2886);
or U6762 (N_6762,N_2110,N_5523);
and U6763 (N_6763,N_3286,N_2269);
and U6764 (N_6764,N_3,N_5276);
or U6765 (N_6765,N_3490,N_2621);
or U6766 (N_6766,N_5451,N_2616);
and U6767 (N_6767,N_5738,N_5937);
xnor U6768 (N_6768,N_2199,N_4385);
and U6769 (N_6769,N_24,N_2610);
or U6770 (N_6770,N_4874,N_2655);
nand U6771 (N_6771,N_3111,N_911);
and U6772 (N_6772,N_4333,N_1824);
or U6773 (N_6773,N_298,N_1732);
nand U6774 (N_6774,N_3176,N_561);
or U6775 (N_6775,N_1604,N_2276);
or U6776 (N_6776,N_41,N_4167);
nor U6777 (N_6777,N_3575,N_3139);
nor U6778 (N_6778,N_5962,N_1064);
and U6779 (N_6779,N_5611,N_3109);
nand U6780 (N_6780,N_1121,N_171);
xor U6781 (N_6781,N_5758,N_2172);
nor U6782 (N_6782,N_5616,N_5429);
nor U6783 (N_6783,N_3125,N_3208);
nor U6784 (N_6784,N_1300,N_4871);
xor U6785 (N_6785,N_4849,N_1374);
xnor U6786 (N_6786,N_3175,N_5460);
and U6787 (N_6787,N_3644,N_5989);
nand U6788 (N_6788,N_3791,N_4989);
or U6789 (N_6789,N_2262,N_377);
nand U6790 (N_6790,N_4787,N_4692);
xnor U6791 (N_6791,N_5270,N_1057);
nor U6792 (N_6792,N_4144,N_2921);
xnor U6793 (N_6793,N_5526,N_767);
nor U6794 (N_6794,N_4650,N_2294);
or U6795 (N_6795,N_4016,N_1680);
and U6796 (N_6796,N_4935,N_3501);
xnor U6797 (N_6797,N_5438,N_4269);
nor U6798 (N_6798,N_1584,N_3592);
or U6799 (N_6799,N_4881,N_2648);
nand U6800 (N_6800,N_4074,N_3523);
nand U6801 (N_6801,N_4523,N_2953);
nand U6802 (N_6802,N_2857,N_3375);
and U6803 (N_6803,N_6164,N_1218);
xnor U6804 (N_6804,N_1613,N_5112);
or U6805 (N_6805,N_2067,N_286);
nor U6806 (N_6806,N_5868,N_3918);
xnor U6807 (N_6807,N_4790,N_5145);
nand U6808 (N_6808,N_5142,N_392);
and U6809 (N_6809,N_2471,N_106);
nor U6810 (N_6810,N_3879,N_5516);
nor U6811 (N_6811,N_4587,N_3980);
or U6812 (N_6812,N_5506,N_3962);
xnor U6813 (N_6813,N_598,N_2241);
xnor U6814 (N_6814,N_4236,N_3275);
and U6815 (N_6815,N_6053,N_4589);
nor U6816 (N_6816,N_197,N_1392);
xor U6817 (N_6817,N_956,N_2945);
nand U6818 (N_6818,N_3008,N_2326);
or U6819 (N_6819,N_1533,N_1499);
or U6820 (N_6820,N_2594,N_1442);
xor U6821 (N_6821,N_5557,N_4581);
xnor U6822 (N_6822,N_4457,N_4347);
or U6823 (N_6823,N_1799,N_497);
nor U6824 (N_6824,N_1180,N_5820);
or U6825 (N_6825,N_4715,N_3202);
nand U6826 (N_6826,N_3473,N_4481);
nor U6827 (N_6827,N_3201,N_5473);
xnor U6828 (N_6828,N_4671,N_6014);
nand U6829 (N_6829,N_2754,N_1850);
nand U6830 (N_6830,N_5105,N_5635);
and U6831 (N_6831,N_5384,N_1707);
or U6832 (N_6832,N_326,N_2096);
or U6833 (N_6833,N_978,N_3818);
xnor U6834 (N_6834,N_5048,N_4439);
nor U6835 (N_6835,N_6048,N_3244);
and U6836 (N_6836,N_2297,N_2124);
or U6837 (N_6837,N_1399,N_3713);
xor U6838 (N_6838,N_2563,N_3039);
xnor U6839 (N_6839,N_5791,N_5544);
and U6840 (N_6840,N_1871,N_2152);
or U6841 (N_6841,N_3714,N_348);
xnor U6842 (N_6842,N_3593,N_4301);
xor U6843 (N_6843,N_5501,N_4204);
xnor U6844 (N_6844,N_1672,N_4688);
nor U6845 (N_6845,N_5025,N_2154);
and U6846 (N_6846,N_3068,N_1439);
or U6847 (N_6847,N_5179,N_5759);
or U6848 (N_6848,N_4793,N_5476);
nor U6849 (N_6849,N_2135,N_368);
xor U6850 (N_6850,N_4259,N_1786);
or U6851 (N_6851,N_3718,N_1330);
or U6852 (N_6852,N_4888,N_942);
or U6853 (N_6853,N_1186,N_4401);
xor U6854 (N_6854,N_6150,N_2464);
nor U6855 (N_6855,N_6162,N_1198);
nand U6856 (N_6856,N_2824,N_747);
nand U6857 (N_6857,N_1190,N_4096);
or U6858 (N_6858,N_1358,N_6182);
nor U6859 (N_6859,N_4740,N_3053);
or U6860 (N_6860,N_2580,N_1466);
xnor U6861 (N_6861,N_6138,N_1649);
xnor U6862 (N_6862,N_3469,N_3665);
and U6863 (N_6863,N_5303,N_3635);
xnor U6864 (N_6864,N_5034,N_5765);
xor U6865 (N_6865,N_1570,N_740);
xnor U6866 (N_6866,N_2376,N_6072);
nand U6867 (N_6867,N_425,N_4304);
and U6868 (N_6868,N_2714,N_3366);
xnor U6869 (N_6869,N_2736,N_1827);
and U6870 (N_6870,N_1642,N_4073);
xor U6871 (N_6871,N_907,N_3150);
xor U6872 (N_6872,N_4135,N_1066);
xor U6873 (N_6873,N_3653,N_5856);
and U6874 (N_6874,N_4858,N_1430);
xor U6875 (N_6875,N_5609,N_5188);
nor U6876 (N_6876,N_846,N_2530);
nor U6877 (N_6877,N_1241,N_3650);
and U6878 (N_6878,N_5087,N_1289);
nand U6879 (N_6879,N_5505,N_3597);
nor U6880 (N_6880,N_3871,N_2557);
nor U6881 (N_6881,N_593,N_4949);
nor U6882 (N_6882,N_522,N_3901);
nor U6883 (N_6883,N_1599,N_3082);
nor U6884 (N_6884,N_3254,N_3507);
and U6885 (N_6885,N_5576,N_4120);
xor U6886 (N_6886,N_3013,N_1195);
and U6887 (N_6887,N_2889,N_4257);
and U6888 (N_6888,N_4218,N_2581);
xnor U6889 (N_6889,N_2435,N_6188);
and U6890 (N_6890,N_510,N_2500);
nor U6891 (N_6891,N_2028,N_5468);
nor U6892 (N_6892,N_5789,N_5315);
nor U6893 (N_6893,N_2892,N_2514);
nand U6894 (N_6894,N_2183,N_884);
and U6895 (N_6895,N_592,N_636);
xor U6896 (N_6896,N_5209,N_198);
and U6897 (N_6897,N_4263,N_5369);
or U6898 (N_6898,N_2646,N_3231);
nor U6899 (N_6899,N_3065,N_5871);
nand U6900 (N_6900,N_1776,N_3926);
and U6901 (N_6901,N_3011,N_1529);
nand U6902 (N_6902,N_3725,N_137);
or U6903 (N_6903,N_511,N_5444);
xor U6904 (N_6904,N_2521,N_3610);
and U6905 (N_6905,N_4649,N_815);
xnor U6906 (N_6906,N_4202,N_2273);
nand U6907 (N_6907,N_80,N_4075);
and U6908 (N_6908,N_2005,N_4048);
and U6909 (N_6909,N_5161,N_2582);
or U6910 (N_6910,N_4015,N_5133);
nand U6911 (N_6911,N_3372,N_4062);
nor U6912 (N_6912,N_550,N_4534);
nor U6913 (N_6913,N_5610,N_5517);
nor U6914 (N_6914,N_1415,N_2251);
or U6915 (N_6915,N_5147,N_950);
and U6916 (N_6916,N_6103,N_4458);
and U6917 (N_6917,N_697,N_3771);
xor U6918 (N_6918,N_5349,N_2598);
xnor U6919 (N_6919,N_2927,N_1637);
nand U6920 (N_6920,N_2227,N_558);
or U6921 (N_6921,N_2210,N_2653);
and U6922 (N_6922,N_2163,N_711);
or U6923 (N_6923,N_178,N_2708);
or U6924 (N_6924,N_4441,N_3284);
nand U6925 (N_6925,N_1449,N_1182);
and U6926 (N_6926,N_5340,N_3198);
nor U6927 (N_6927,N_4093,N_3981);
nand U6928 (N_6928,N_4644,N_4529);
and U6929 (N_6929,N_5717,N_5608);
or U6930 (N_6930,N_2472,N_1683);
nand U6931 (N_6931,N_4786,N_574);
nand U6932 (N_6932,N_429,N_338);
nand U6933 (N_6933,N_2543,N_2094);
nor U6934 (N_6934,N_5903,N_4708);
xor U6935 (N_6935,N_4810,N_1332);
or U6936 (N_6936,N_657,N_5352);
nand U6937 (N_6937,N_4959,N_5344);
nor U6938 (N_6938,N_1928,N_651);
or U6939 (N_6939,N_2391,N_2185);
and U6940 (N_6940,N_1705,N_5628);
nand U6941 (N_6941,N_6082,N_4756);
or U6942 (N_6942,N_1115,N_4833);
or U6943 (N_6943,N_864,N_1237);
and U6944 (N_6944,N_4478,N_2914);
xnor U6945 (N_6945,N_2149,N_5940);
or U6946 (N_6946,N_739,N_2596);
nor U6947 (N_6947,N_3302,N_2558);
nand U6948 (N_6948,N_1991,N_1225);
xor U6949 (N_6949,N_2575,N_1727);
or U6950 (N_6950,N_4554,N_1554);
nand U6951 (N_6951,N_2010,N_1440);
nand U6952 (N_6952,N_3048,N_4953);
nand U6953 (N_6953,N_1338,N_4758);
or U6954 (N_6954,N_2834,N_1101);
or U6955 (N_6955,N_3463,N_4321);
or U6956 (N_6956,N_1953,N_3784);
nor U6957 (N_6957,N_5876,N_1622);
nand U6958 (N_6958,N_1598,N_4307);
nor U6959 (N_6959,N_2782,N_3522);
or U6960 (N_6960,N_100,N_90);
xnor U6961 (N_6961,N_5328,N_860);
and U6962 (N_6962,N_4651,N_5996);
nor U6963 (N_6963,N_5915,N_5886);
or U6964 (N_6964,N_3600,N_2997);
nor U6965 (N_6965,N_6121,N_974);
nor U6966 (N_6966,N_4049,N_4006);
or U6967 (N_6967,N_4213,N_5997);
nand U6968 (N_6968,N_3663,N_4707);
and U6969 (N_6969,N_4637,N_203);
nor U6970 (N_6970,N_323,N_1306);
nand U6971 (N_6971,N_4224,N_4785);
or U6972 (N_6972,N_3595,N_1450);
or U6973 (N_6973,N_4421,N_1476);
nand U6974 (N_6974,N_5666,N_156);
xnor U6975 (N_6975,N_4625,N_5118);
or U6976 (N_6976,N_5192,N_4552);
xnor U6977 (N_6977,N_4415,N_1388);
nand U6978 (N_6978,N_3542,N_3019);
xnor U6979 (N_6979,N_3022,N_4509);
and U6980 (N_6980,N_3023,N_5376);
nor U6981 (N_6981,N_3915,N_1658);
nand U6982 (N_6982,N_1168,N_1291);
and U6983 (N_6983,N_3271,N_5818);
nor U6984 (N_6984,N_5016,N_3701);
or U6985 (N_6985,N_4045,N_6141);
or U6986 (N_6986,N_2527,N_3861);
or U6987 (N_6987,N_3859,N_4617);
or U6988 (N_6988,N_3735,N_924);
or U6989 (N_6989,N_4851,N_5572);
and U6990 (N_6990,N_1972,N_755);
nor U6991 (N_6991,N_3719,N_2219);
and U6992 (N_6992,N_750,N_3889);
nand U6993 (N_6993,N_1869,N_2268);
nand U6994 (N_6994,N_3620,N_5917);
or U6995 (N_6995,N_2098,N_6078);
nand U6996 (N_6996,N_5504,N_1294);
nor U6997 (N_6997,N_5162,N_3917);
nor U6998 (N_6998,N_525,N_708);
nand U6999 (N_6999,N_5343,N_3624);
nand U7000 (N_7000,N_2649,N_1017);
or U7001 (N_7001,N_1318,N_2460);
and U7002 (N_7002,N_1693,N_6131);
nand U7003 (N_7003,N_2666,N_3770);
nor U7004 (N_7004,N_4836,N_5136);
nand U7005 (N_7005,N_421,N_2803);
nand U7006 (N_7006,N_330,N_1934);
nand U7007 (N_7007,N_1942,N_5383);
and U7008 (N_7008,N_2323,N_3726);
or U7009 (N_7009,N_1757,N_1795);
and U7010 (N_7010,N_4271,N_5603);
and U7011 (N_7011,N_2164,N_193);
nand U7012 (N_7012,N_2659,N_4893);
xor U7013 (N_7013,N_217,N_3902);
nor U7014 (N_7014,N_5907,N_1818);
or U7015 (N_7015,N_3654,N_6064);
xor U7016 (N_7016,N_2908,N_1131);
nor U7017 (N_7017,N_230,N_989);
or U7018 (N_7018,N_15,N_4930);
nand U7019 (N_7019,N_3812,N_2775);
xor U7020 (N_7020,N_3436,N_5143);
xnor U7021 (N_7021,N_5051,N_4676);
xor U7022 (N_7022,N_3706,N_3525);
xnor U7023 (N_7023,N_3057,N_5676);
nor U7024 (N_7024,N_2463,N_2896);
and U7025 (N_7025,N_1573,N_3857);
nand U7026 (N_7026,N_3727,N_2133);
or U7027 (N_7027,N_713,N_4319);
or U7028 (N_7028,N_977,N_2924);
and U7029 (N_7029,N_5367,N_160);
nand U7030 (N_7030,N_5309,N_2034);
and U7031 (N_7031,N_2591,N_822);
and U7032 (N_7032,N_4208,N_4947);
nand U7033 (N_7033,N_3229,N_5433);
and U7034 (N_7034,N_3067,N_4684);
nor U7035 (N_7035,N_5238,N_3076);
and U7036 (N_7036,N_2498,N_3353);
nand U7037 (N_7037,N_2589,N_727);
and U7038 (N_7038,N_2235,N_1612);
nor U7039 (N_7039,N_1356,N_3682);
nor U7040 (N_7040,N_4295,N_2092);
xor U7041 (N_7041,N_2909,N_412);
or U7042 (N_7042,N_976,N_2439);
xor U7043 (N_7043,N_3004,N_1830);
nand U7044 (N_7044,N_2826,N_2111);
and U7045 (N_7045,N_134,N_4663);
and U7046 (N_7046,N_1591,N_4070);
nand U7047 (N_7047,N_4528,N_3452);
nand U7048 (N_7048,N_3280,N_3349);
xnor U7049 (N_7049,N_606,N_8);
or U7050 (N_7050,N_3330,N_2663);
xor U7051 (N_7051,N_2193,N_4857);
or U7052 (N_7052,N_1197,N_1487);
nor U7053 (N_7053,N_5522,N_3472);
or U7054 (N_7054,N_3158,N_3562);
nor U7055 (N_7055,N_5207,N_2140);
xnor U7056 (N_7056,N_2941,N_6187);
xnor U7057 (N_7057,N_5928,N_4765);
and U7058 (N_7058,N_2237,N_1550);
xnor U7059 (N_7059,N_6083,N_5102);
nor U7060 (N_7060,N_4468,N_4664);
or U7061 (N_7061,N_1145,N_1299);
and U7062 (N_7062,N_264,N_684);
nor U7063 (N_7063,N_5629,N_3132);
nor U7064 (N_7064,N_2702,N_1567);
xnor U7065 (N_7065,N_413,N_4598);
or U7066 (N_7066,N_2780,N_2705);
nand U7067 (N_7067,N_3273,N_2341);
nand U7068 (N_7068,N_3977,N_4624);
xnor U7069 (N_7069,N_4872,N_3817);
and U7070 (N_7070,N_3386,N_2416);
nand U7071 (N_7071,N_4686,N_2446);
xnor U7072 (N_7072,N_3517,N_394);
and U7073 (N_7073,N_2990,N_4334);
nand U7074 (N_7074,N_3355,N_4277);
nor U7075 (N_7075,N_2986,N_763);
nand U7076 (N_7076,N_1715,N_4721);
and U7077 (N_7077,N_6105,N_1024);
or U7078 (N_7078,N_5793,N_2740);
nand U7079 (N_7079,N_2748,N_3564);
nand U7080 (N_7080,N_4398,N_5632);
or U7081 (N_7081,N_3045,N_4037);
xnor U7082 (N_7082,N_3904,N_3740);
nand U7083 (N_7083,N_5671,N_1971);
and U7084 (N_7084,N_1582,N_6092);
and U7085 (N_7085,N_5231,N_1563);
nand U7086 (N_7086,N_2475,N_1983);
xnor U7087 (N_7087,N_428,N_4675);
nand U7088 (N_7088,N_293,N_638);
nor U7089 (N_7089,N_2677,N_1954);
nand U7090 (N_7090,N_5803,N_3849);
nor U7091 (N_7091,N_5844,N_5638);
xor U7092 (N_7092,N_4287,N_6244);
or U7093 (N_7093,N_2727,N_1708);
nor U7094 (N_7094,N_4229,N_2494);
xnor U7095 (N_7095,N_540,N_4210);
nand U7096 (N_7096,N_2171,N_3214);
nor U7097 (N_7097,N_1674,N_5267);
xnor U7098 (N_7098,N_3789,N_6003);
xnor U7099 (N_7099,N_2524,N_4240);
or U7100 (N_7100,N_5200,N_4711);
nor U7101 (N_7101,N_3242,N_243);
nor U7102 (N_7102,N_3821,N_4738);
xor U7103 (N_7103,N_295,N_4771);
or U7104 (N_7104,N_4379,N_5427);
xor U7105 (N_7105,N_5599,N_3409);
nor U7106 (N_7106,N_3230,N_5260);
and U7107 (N_7107,N_1697,N_5155);
nor U7108 (N_7108,N_5556,N_6237);
xnor U7109 (N_7109,N_4789,N_5975);
nor U7110 (N_7110,N_3282,N_5302);
or U7111 (N_7111,N_4517,N_571);
or U7112 (N_7112,N_5072,N_5736);
xor U7113 (N_7113,N_2515,N_1012);
nand U7114 (N_7114,N_447,N_4909);
or U7115 (N_7115,N_1617,N_285);
nor U7116 (N_7116,N_3919,N_3520);
and U7117 (N_7117,N_919,N_5695);
and U7118 (N_7118,N_3983,N_1651);
xor U7119 (N_7119,N_449,N_455);
xor U7120 (N_7120,N_1307,N_3872);
xnor U7121 (N_7121,N_176,N_494);
or U7122 (N_7122,N_2037,N_4843);
nor U7123 (N_7123,N_2337,N_3998);
nand U7124 (N_7124,N_5098,N_1775);
nand U7125 (N_7125,N_3055,N_2324);
or U7126 (N_7126,N_2054,N_1610);
xnor U7127 (N_7127,N_2793,N_1428);
and U7128 (N_7128,N_5721,N_161);
nor U7129 (N_7129,N_1130,N_1258);
xnor U7130 (N_7130,N_2233,N_119);
xnor U7131 (N_7131,N_287,N_4585);
and U7132 (N_7132,N_3975,N_6004);
nor U7133 (N_7133,N_4932,N_6160);
nand U7134 (N_7134,N_2050,N_2121);
xnor U7135 (N_7135,N_4772,N_3081);
nor U7136 (N_7136,N_4646,N_4335);
and U7137 (N_7137,N_2778,N_1208);
and U7138 (N_7138,N_752,N_1040);
or U7139 (N_7139,N_89,N_2053);
nand U7140 (N_7140,N_6000,N_5241);
nand U7141 (N_7141,N_1417,N_3699);
xnor U7142 (N_7142,N_2599,N_2290);
nand U7143 (N_7143,N_5976,N_3296);
xor U7144 (N_7144,N_1910,N_1433);
and U7145 (N_7145,N_4805,N_1256);
or U7146 (N_7146,N_1055,N_5248);
nand U7147 (N_7147,N_4716,N_4017);
nand U7148 (N_7148,N_2496,N_88);
and U7149 (N_7149,N_4803,N_2560);
or U7150 (N_7150,N_3692,N_2593);
or U7151 (N_7151,N_4656,N_4414);
xor U7152 (N_7152,N_5600,N_5507);
nor U7153 (N_7153,N_3888,N_3077);
and U7154 (N_7154,N_3058,N_1845);
nor U7155 (N_7155,N_2933,N_2456);
nand U7156 (N_7156,N_2696,N_2266);
xnor U7157 (N_7157,N_1764,N_4485);
nor U7158 (N_7158,N_2679,N_4261);
nor U7159 (N_7159,N_1993,N_2768);
and U7160 (N_7160,N_2635,N_3974);
and U7161 (N_7161,N_1810,N_3894);
nor U7162 (N_7162,N_3169,N_3205);
xor U7163 (N_7163,N_4615,N_1456);
xor U7164 (N_7164,N_4886,N_1594);
nand U7165 (N_7165,N_4974,N_1968);
and U7166 (N_7166,N_2903,N_3864);
xor U7167 (N_7167,N_4755,N_1203);
nand U7168 (N_7168,N_3289,N_3732);
nor U7169 (N_7169,N_5641,N_1842);
nor U7170 (N_7170,N_6026,N_2710);
nor U7171 (N_7171,N_6148,N_2438);
or U7172 (N_7172,N_1551,N_1070);
xor U7173 (N_7173,N_4377,N_2811);
or U7174 (N_7174,N_1848,N_5284);
nor U7175 (N_7175,N_4995,N_4034);
nand U7176 (N_7176,N_1309,N_1290);
nor U7177 (N_7177,N_1473,N_3190);
or U7178 (N_7178,N_1897,N_4887);
and U7179 (N_7179,N_4597,N_1232);
xnor U7180 (N_7180,N_590,N_4497);
or U7181 (N_7181,N_4059,N_3426);
and U7182 (N_7182,N_4940,N_2493);
xnor U7183 (N_7183,N_6027,N_367);
nor U7184 (N_7184,N_2226,N_94);
or U7185 (N_7185,N_5452,N_3220);
nor U7186 (N_7186,N_4289,N_2166);
and U7187 (N_7187,N_889,N_3098);
xor U7188 (N_7188,N_155,N_4992);
nor U7189 (N_7189,N_4998,N_432);
xnor U7190 (N_7190,N_3599,N_6174);
nor U7191 (N_7191,N_1520,N_4150);
nand U7192 (N_7192,N_1231,N_4853);
and U7193 (N_7193,N_1261,N_431);
or U7194 (N_7194,N_1997,N_5390);
xnor U7195 (N_7195,N_1833,N_2433);
or U7196 (N_7196,N_6001,N_5618);
or U7197 (N_7197,N_5964,N_40);
nor U7198 (N_7198,N_4759,N_1013);
xor U7199 (N_7199,N_774,N_2300);
xor U7200 (N_7200,N_5348,N_4524);
or U7201 (N_7201,N_4894,N_1750);
xnor U7202 (N_7202,N_5467,N_1844);
and U7203 (N_7203,N_2660,N_43);
nor U7204 (N_7204,N_583,N_1924);
nand U7205 (N_7205,N_4163,N_1408);
nand U7206 (N_7206,N_4969,N_2822);
xnor U7207 (N_7207,N_4722,N_2490);
or U7208 (N_7208,N_1002,N_2495);
or U7209 (N_7209,N_5991,N_3154);
xor U7210 (N_7210,N_4351,N_3548);
or U7211 (N_7211,N_5245,N_3410);
nor U7212 (N_7212,N_4922,N_2364);
and U7213 (N_7213,N_4639,N_5306);
and U7214 (N_7214,N_908,N_95);
and U7215 (N_7215,N_61,N_3785);
or U7216 (N_7216,N_2678,N_3167);
nand U7217 (N_7217,N_1285,N_3475);
xnor U7218 (N_7218,N_2355,N_6222);
xor U7219 (N_7219,N_5586,N_1058);
or U7220 (N_7220,N_2077,N_585);
or U7221 (N_7221,N_1821,N_2427);
nand U7222 (N_7222,N_2257,N_4242);
nor U7223 (N_7223,N_5347,N_2861);
nor U7224 (N_7224,N_5739,N_2551);
nor U7225 (N_7225,N_775,N_2120);
xnor U7226 (N_7226,N_4413,N_3040);
xor U7227 (N_7227,N_812,N_5399);
or U7228 (N_7228,N_4661,N_2032);
and U7229 (N_7229,N_4801,N_4632);
nor U7230 (N_7230,N_5767,N_1758);
nor U7231 (N_7231,N_2352,N_1069);
xnor U7232 (N_7232,N_5681,N_4519);
or U7233 (N_7233,N_5410,N_211);
xnor U7234 (N_7234,N_4143,N_5341);
nor U7235 (N_7235,N_4769,N_764);
and U7236 (N_7236,N_2206,N_1741);
or U7237 (N_7237,N_5373,N_5673);
xor U7238 (N_7238,N_1371,N_2319);
xor U7239 (N_7239,N_5134,N_2372);
xor U7240 (N_7240,N_4683,N_3551);
nor U7241 (N_7241,N_5813,N_120);
and U7242 (N_7242,N_5891,N_2985);
xor U7243 (N_7243,N_396,N_2443);
xor U7244 (N_7244,N_2363,N_987);
and U7245 (N_7245,N_3848,N_2756);
and U7246 (N_7246,N_4822,N_2499);
nor U7247 (N_7247,N_1710,N_2264);
or U7248 (N_7248,N_4806,N_5396);
and U7249 (N_7249,N_1756,N_1921);
and U7250 (N_7250,N_921,N_3451);
or U7251 (N_7251,N_4076,N_5640);
or U7252 (N_7252,N_5731,N_1907);
and U7253 (N_7253,N_855,N_4791);
or U7254 (N_7254,N_3947,N_1886);
nor U7255 (N_7255,N_1985,N_2134);
nand U7256 (N_7256,N_5003,N_336);
nand U7257 (N_7257,N_766,N_2712);
and U7258 (N_7258,N_3344,N_402);
xor U7259 (N_7259,N_1646,N_2535);
nand U7260 (N_7260,N_5689,N_3972);
or U7261 (N_7261,N_5949,N_4363);
and U7262 (N_7262,N_3601,N_2123);
or U7263 (N_7263,N_586,N_5251);
and U7264 (N_7264,N_6009,N_4745);
nand U7265 (N_7265,N_1063,N_4718);
and U7266 (N_7266,N_5571,N_958);
or U7267 (N_7267,N_537,N_930);
or U7268 (N_7268,N_4612,N_3191);
nor U7269 (N_7269,N_3411,N_165);
nand U7270 (N_7270,N_549,N_2293);
nand U7271 (N_7271,N_1722,N_5761);
nor U7272 (N_7272,N_294,N_5024);
nand U7273 (N_7273,N_3050,N_1155);
xor U7274 (N_7274,N_4044,N_2167);
or U7275 (N_7275,N_1944,N_3518);
nor U7276 (N_7276,N_672,N_4047);
or U7277 (N_7277,N_3863,N_1789);
nor U7278 (N_7278,N_2381,N_4904);
xor U7279 (N_7279,N_2969,N_5358);
nand U7280 (N_7280,N_5033,N_3325);
xor U7281 (N_7281,N_5150,N_3103);
nand U7282 (N_7282,N_4957,N_796);
and U7283 (N_7283,N_4903,N_4305);
nor U7284 (N_7284,N_5545,N_6194);
xor U7285 (N_7285,N_2272,N_464);
and U7286 (N_7286,N_5114,N_4249);
or U7287 (N_7287,N_4149,N_808);
nand U7288 (N_7288,N_1339,N_5707);
xnor U7289 (N_7289,N_3651,N_810);
and U7290 (N_7290,N_5898,N_5780);
nand U7291 (N_7291,N_1540,N_3839);
xor U7292 (N_7292,N_2970,N_948);
xor U7293 (N_7293,N_4170,N_1126);
nor U7294 (N_7294,N_3394,N_5018);
and U7295 (N_7295,N_5199,N_3657);
xnor U7296 (N_7296,N_4146,N_415);
nor U7297 (N_7297,N_3967,N_305);
nand U7298 (N_7298,N_5675,N_3796);
or U7299 (N_7299,N_2420,N_1419);
nand U7300 (N_7300,N_1288,N_737);
xnor U7301 (N_7301,N_6070,N_5918);
nand U7302 (N_7302,N_3584,N_1878);
nor U7303 (N_7303,N_2643,N_4101);
or U7304 (N_7304,N_2147,N_2365);
nor U7305 (N_7305,N_4035,N_1882);
nand U7306 (N_7306,N_1049,N_4440);
nand U7307 (N_7307,N_4636,N_1832);
nand U7308 (N_7308,N_1738,N_613);
xor U7309 (N_7309,N_2488,N_1380);
xor U7310 (N_7310,N_1367,N_2912);
nor U7311 (N_7311,N_3498,N_152);
or U7312 (N_7312,N_972,N_2713);
nand U7313 (N_7313,N_4870,N_3722);
or U7314 (N_7314,N_1901,N_4303);
and U7315 (N_7315,N_3433,N_187);
nor U7316 (N_7316,N_5657,N_4628);
xnor U7317 (N_7317,N_1863,N_39);
xor U7318 (N_7318,N_5566,N_1378);
or U7319 (N_7319,N_2812,N_505);
nor U7320 (N_7320,N_4187,N_2553);
nand U7321 (N_7321,N_3799,N_5541);
xor U7322 (N_7322,N_3586,N_890);
nor U7323 (N_7323,N_594,N_5875);
xor U7324 (N_7324,N_665,N_3142);
nand U7325 (N_7325,N_2170,N_2466);
nand U7326 (N_7326,N_5499,N_1937);
and U7327 (N_7327,N_2392,N_4512);
xor U7328 (N_7328,N_2602,N_4200);
nand U7329 (N_7329,N_975,N_587);
nor U7330 (N_7330,N_786,N_4109);
nor U7331 (N_7331,N_1751,N_738);
nand U7332 (N_7332,N_1120,N_4371);
xor U7333 (N_7333,N_5627,N_973);
or U7334 (N_7334,N_247,N_1276);
or U7335 (N_7335,N_1894,N_6175);
and U7336 (N_7336,N_1468,N_2086);
nor U7337 (N_7337,N_3970,N_3226);
xnor U7338 (N_7338,N_5318,N_2522);
or U7339 (N_7339,N_1723,N_3376);
xor U7340 (N_7340,N_1914,N_3287);
and U7341 (N_7341,N_2358,N_4846);
or U7342 (N_7342,N_1039,N_646);
and U7343 (N_7343,N_4244,N_1015);
xor U7344 (N_7344,N_6008,N_986);
or U7345 (N_7345,N_754,N_1814);
or U7346 (N_7346,N_5858,N_118);
nor U7347 (N_7347,N_3332,N_2027);
nor U7348 (N_7348,N_5160,N_762);
nand U7349 (N_7349,N_5266,N_2485);
nand U7350 (N_7350,N_4325,N_1618);
or U7351 (N_7351,N_221,N_4164);
nand U7352 (N_7352,N_5183,N_2821);
xnor U7353 (N_7353,N_682,N_4719);
nor U7354 (N_7354,N_5196,N_6245);
nor U7355 (N_7355,N_3569,N_4584);
xor U7356 (N_7356,N_5233,N_4196);
xnor U7357 (N_7357,N_4106,N_4174);
nand U7358 (N_7358,N_2827,N_1890);
nand U7359 (N_7359,N_4720,N_3161);
nor U7360 (N_7360,N_5665,N_2650);
xor U7361 (N_7361,N_2568,N_2747);
and U7362 (N_7362,N_1811,N_5649);
or U7363 (N_7363,N_2117,N_2359);
xnor U7364 (N_7364,N_4815,N_5203);
nand U7365 (N_7365,N_944,N_6213);
nand U7366 (N_7366,N_3929,N_1766);
nor U7367 (N_7367,N_2295,N_616);
and U7368 (N_7368,N_6192,N_4116);
or U7369 (N_7369,N_4831,N_4254);
xnor U7370 (N_7370,N_3233,N_714);
nand U7371 (N_7371,N_3465,N_2444);
xor U7372 (N_7372,N_5733,N_625);
nand U7373 (N_7373,N_5661,N_3255);
or U7374 (N_7374,N_2087,N_2078);
nor U7375 (N_7375,N_1696,N_2630);
nand U7376 (N_7376,N_3428,N_5920);
xor U7377 (N_7377,N_2325,N_3712);
nand U7378 (N_7378,N_82,N_353);
xnor U7379 (N_7379,N_3819,N_3389);
nor U7380 (N_7380,N_4911,N_4616);
or U7381 (N_7381,N_2516,N_5838);
or U7382 (N_7382,N_5494,N_2051);
or U7383 (N_7383,N_4850,N_3780);
xor U7384 (N_7384,N_2992,N_3499);
nand U7385 (N_7385,N_5182,N_4400);
nor U7386 (N_7386,N_811,N_923);
xnor U7387 (N_7387,N_487,N_2652);
nand U7388 (N_7388,N_4948,N_4580);
xor U7389 (N_7389,N_1060,N_1561);
nor U7390 (N_7390,N_1328,N_1434);
or U7391 (N_7391,N_6153,N_3350);
nand U7392 (N_7392,N_1150,N_640);
or U7393 (N_7393,N_6117,N_4794);
and U7394 (N_7394,N_3274,N_3427);
xor U7395 (N_7395,N_2243,N_1072);
or U7396 (N_7396,N_6055,N_4192);
and U7397 (N_7397,N_465,N_620);
or U7398 (N_7398,N_1728,N_2988);
nor U7399 (N_7399,N_3505,N_249);
and U7400 (N_7400,N_4812,N_1405);
and U7401 (N_7401,N_4586,N_1045);
nor U7402 (N_7402,N_2492,N_146);
or U7403 (N_7403,N_5088,N_2021);
xor U7404 (N_7404,N_5511,N_4582);
or U7405 (N_7405,N_2351,N_4925);
nor U7406 (N_7406,N_491,N_5418);
nand U7407 (N_7407,N_4638,N_4717);
nand U7408 (N_7408,N_3118,N_6235);
xor U7409 (N_7409,N_3378,N_6040);
and U7410 (N_7410,N_5056,N_3304);
nor U7411 (N_7411,N_4897,N_2478);
nand U7412 (N_7412,N_6193,N_3723);
nor U7413 (N_7413,N_1855,N_5311);
nor U7414 (N_7414,N_3800,N_3767);
and U7415 (N_7415,N_4194,N_4470);
or U7416 (N_7416,N_6181,N_3354);
xnor U7417 (N_7417,N_5967,N_3669);
nor U7418 (N_7418,N_4342,N_4521);
xor U7419 (N_7419,N_5821,N_1459);
and U7420 (N_7420,N_5036,N_1477);
xnor U7421 (N_7421,N_1535,N_2387);
xor U7422 (N_7422,N_4535,N_1124);
nor U7423 (N_7423,N_3855,N_3380);
or U7424 (N_7424,N_5924,N_5324);
and U7425 (N_7425,N_3072,N_1059);
xor U7426 (N_7426,N_5194,N_5702);
or U7427 (N_7427,N_4423,N_599);
or U7428 (N_7428,N_4350,N_272);
xor U7429 (N_7429,N_5679,N_5559);
xnor U7430 (N_7430,N_4014,N_6065);
or U7431 (N_7431,N_5490,N_3406);
or U7432 (N_7432,N_518,N_787);
xnor U7433 (N_7433,N_4784,N_301);
nor U7434 (N_7434,N_3696,N_4982);
nand U7435 (N_7435,N_3768,N_6126);
or U7436 (N_7436,N_1215,N_2287);
nand U7437 (N_7437,N_2317,N_6191);
xnor U7438 (N_7438,N_2541,N_113);
or U7439 (N_7439,N_637,N_2567);
xnor U7440 (N_7440,N_4838,N_5113);
nand U7441 (N_7441,N_1984,N_6045);
nor U7442 (N_7442,N_5239,N_5771);
or U7443 (N_7443,N_4429,N_1699);
nor U7444 (N_7444,N_1495,N_185);
nor U7445 (N_7445,N_3288,N_2971);
nand U7446 (N_7446,N_878,N_478);
or U7447 (N_7447,N_536,N_3322);
or U7448 (N_7448,N_4030,N_1966);
nand U7449 (N_7449,N_2800,N_1426);
nand U7450 (N_7450,N_4777,N_52);
or U7451 (N_7451,N_4306,N_5032);
and U7452 (N_7452,N_5806,N_4060);
or U7453 (N_7453,N_5346,N_4382);
nand U7454 (N_7454,N_1840,N_5696);
nand U7455 (N_7455,N_3534,N_4504);
and U7456 (N_7456,N_3266,N_2244);
xnor U7457 (N_7457,N_1054,N_3034);
nor U7458 (N_7458,N_800,N_4693);
and U7459 (N_7459,N_2699,N_1220);
and U7460 (N_7460,N_2207,N_4256);
nand U7461 (N_7461,N_2936,N_4343);
nor U7462 (N_7462,N_6217,N_5685);
xnor U7463 (N_7463,N_5380,N_4555);
nand U7464 (N_7464,N_3687,N_420);
xnor U7465 (N_7465,N_1127,N_3952);
and U7466 (N_7466,N_5381,N_181);
nor U7467 (N_7467,N_3241,N_3843);
nand U7468 (N_7468,N_3369,N_4302);
xnor U7469 (N_7469,N_573,N_5084);
nand U7470 (N_7470,N_5043,N_4908);
or U7471 (N_7471,N_5191,N_3443);
nand U7472 (N_7472,N_2270,N_2717);
nand U7473 (N_7473,N_5259,N_5449);
xnor U7474 (N_7474,N_5799,N_3146);
or U7475 (N_7475,N_5703,N_1645);
and U7476 (N_7476,N_3958,N_1703);
or U7477 (N_7477,N_2431,N_117);
nand U7478 (N_7478,N_3704,N_5172);
and U7479 (N_7479,N_3323,N_3338);
nor U7480 (N_7480,N_5121,N_4768);
or U7481 (N_7481,N_4199,N_372);
or U7482 (N_7482,N_716,N_2213);
nand U7483 (N_7483,N_2963,N_5177);
nor U7484 (N_7484,N_4128,N_5061);
or U7485 (N_7485,N_3277,N_115);
or U7486 (N_7486,N_3984,N_3661);
or U7487 (N_7487,N_1572,N_2411);
or U7488 (N_7488,N_4551,N_4420);
xor U7489 (N_7489,N_4250,N_1498);
or U7490 (N_7490,N_1029,N_3910);
or U7491 (N_7491,N_701,N_2633);
or U7492 (N_7492,N_686,N_297);
or U7493 (N_7493,N_2203,N_6120);
xor U7494 (N_7494,N_5197,N_17);
nand U7495 (N_7495,N_3509,N_951);
or U7496 (N_7496,N_3400,N_780);
nor U7497 (N_7497,N_3056,N_1216);
nor U7498 (N_7498,N_5307,N_4309);
nor U7499 (N_7499,N_2406,N_5850);
and U7500 (N_7500,N_6219,N_458);
nor U7501 (N_7501,N_5879,N_5078);
xor U7502 (N_7502,N_2068,N_5104);
xnor U7503 (N_7503,N_5847,N_2681);
and U7504 (N_7504,N_1292,N_220);
nor U7505 (N_7505,N_3590,N_5319);
nand U7506 (N_7506,N_938,N_2513);
nand U7507 (N_7507,N_4462,N_6018);
xor U7508 (N_7508,N_578,N_3611);
nor U7509 (N_7509,N_5909,N_5286);
nor U7510 (N_7510,N_3259,N_3824);
nand U7511 (N_7511,N_2565,N_73);
xnor U7512 (N_7512,N_4840,N_3892);
and U7513 (N_7513,N_2520,N_5206);
nand U7514 (N_7514,N_1541,N_1252);
and U7515 (N_7515,N_4703,N_3623);
nand U7516 (N_7516,N_404,N_5314);
xor U7517 (N_7517,N_5020,N_854);
nand U7518 (N_7518,N_4367,N_554);
and U7519 (N_7519,N_2629,N_5458);
and U7520 (N_7520,N_6052,N_5525);
or U7521 (N_7521,N_2157,N_191);
xor U7522 (N_7522,N_5035,N_2070);
and U7523 (N_7523,N_3006,N_2707);
and U7524 (N_7524,N_5371,N_2766);
or U7525 (N_7525,N_835,N_5798);
xor U7526 (N_7526,N_2923,N_5021);
nor U7527 (N_7527,N_4104,N_3786);
nor U7528 (N_7528,N_631,N_3337);
and U7529 (N_7529,N_2236,N_5462);
nand U7530 (N_7530,N_4184,N_568);
xor U7531 (N_7531,N_27,N_4802);
or U7532 (N_7532,N_2836,N_5019);
or U7533 (N_7533,N_1624,N_5497);
xnor U7534 (N_7534,N_4241,N_1911);
nor U7535 (N_7535,N_3989,N_2389);
xor U7536 (N_7536,N_3615,N_1929);
nor U7537 (N_7537,N_2758,N_4003);
nand U7538 (N_7538,N_4518,N_4387);
and U7539 (N_7539,N_3825,N_1211);
and U7540 (N_7540,N_4091,N_4300);
or U7541 (N_7541,N_282,N_1253);
nand U7542 (N_7542,N_4937,N_2250);
nand U7543 (N_7543,N_3579,N_3061);
nor U7544 (N_7544,N_5981,N_3324);
or U7545 (N_7545,N_6006,N_3434);
xor U7546 (N_7546,N_4419,N_4227);
and U7547 (N_7547,N_20,N_1643);
or U7548 (N_7548,N_3301,N_2198);
nor U7549 (N_7549,N_2920,N_4058);
xor U7550 (N_7550,N_5230,N_5361);
nand U7551 (N_7551,N_4431,N_5175);
and U7552 (N_7552,N_2105,N_98);
xnor U7553 (N_7553,N_519,N_4331);
nand U7554 (N_7554,N_6143,N_3466);
xnor U7555 (N_7555,N_5622,N_6023);
nor U7556 (N_7556,N_4183,N_817);
xnor U7557 (N_7557,N_6154,N_642);
nand U7558 (N_7558,N_6124,N_3384);
and U7559 (N_7559,N_2890,N_1436);
nor U7560 (N_7560,N_177,N_5453);
and U7561 (N_7561,N_4267,N_1207);
nand U7562 (N_7562,N_5828,N_311);
nand U7563 (N_7563,N_4337,N_3160);
xor U7564 (N_7564,N_3488,N_173);
nor U7565 (N_7565,N_5538,N_595);
xnor U7566 (N_7566,N_3261,N_3636);
xnor U7567 (N_7567,N_2026,N_2018);
nor U7568 (N_7568,N_999,N_2469);
and U7569 (N_7569,N_514,N_861);
nand U7570 (N_7570,N_5379,N_2724);
xnor U7571 (N_7571,N_5484,N_2128);
nand U7572 (N_7572,N_70,N_1011);
or U7573 (N_7573,N_597,N_4082);
or U7574 (N_7574,N_5167,N_205);
nand U7575 (N_7575,N_2828,N_1107);
and U7576 (N_7576,N_2309,N_2571);
nand U7577 (N_7577,N_3291,N_3633);
xnor U7578 (N_7578,N_179,N_5054);
nor U7579 (N_7579,N_2075,N_4544);
nand U7580 (N_7580,N_2489,N_5726);
xor U7581 (N_7581,N_5455,N_858);
and U7582 (N_7582,N_5005,N_5591);
nor U7583 (N_7583,N_2281,N_532);
and U7584 (N_7584,N_507,N_278);
nor U7585 (N_7585,N_1669,N_1509);
nand U7586 (N_7586,N_6022,N_4873);
nand U7587 (N_7587,N_4878,N_1796);
or U7588 (N_7588,N_1176,N_4134);
or U7589 (N_7589,N_4537,N_3165);
nor U7590 (N_7590,N_2388,N_4748);
xor U7591 (N_7591,N_3245,N_4473);
and U7592 (N_7592,N_4880,N_5770);
nand U7593 (N_7593,N_6069,N_2298);
and U7594 (N_7594,N_250,N_632);
and U7595 (N_7595,N_1056,N_2680);
xnor U7596 (N_7596,N_1469,N_2333);
and U7597 (N_7597,N_5569,N_2);
or U7598 (N_7598,N_204,N_5254);
or U7599 (N_7599,N_6132,N_1236);
nand U7600 (N_7600,N_2730,N_4923);
nand U7601 (N_7601,N_6084,N_1712);
or U7602 (N_7602,N_3105,N_2043);
nor U7603 (N_7603,N_5735,N_5890);
nor U7604 (N_7604,N_1444,N_6032);
nor U7605 (N_7605,N_5710,N_5228);
or U7606 (N_7606,N_5777,N_1418);
nand U7607 (N_7607,N_1140,N_4631);
xor U7608 (N_7608,N_1725,N_3021);
or U7609 (N_7609,N_1395,N_2512);
xnor U7610 (N_7610,N_1630,N_4063);
xor U7611 (N_7611,N_1099,N_3320);
nand U7612 (N_7612,N_3379,N_6173);
or U7613 (N_7613,N_2002,N_993);
nand U7614 (N_7614,N_6206,N_4079);
nand U7615 (N_7615,N_1103,N_4951);
nand U7616 (N_7616,N_327,N_2011);
nand U7617 (N_7617,N_4590,N_214);
and U7618 (N_7618,N_3898,N_48);
and U7619 (N_7619,N_551,N_4859);
xnor U7620 (N_7620,N_4326,N_947);
nand U7621 (N_7621,N_3903,N_757);
nor U7622 (N_7622,N_3893,N_6068);
and U7623 (N_7623,N_2249,N_5979);
nor U7624 (N_7624,N_6013,N_946);
xor U7625 (N_7625,N_3764,N_4914);
nor U7626 (N_7626,N_5333,N_22);
nor U7627 (N_7627,N_969,N_1488);
nor U7628 (N_7628,N_785,N_3700);
or U7629 (N_7629,N_2574,N_4416);
xor U7630 (N_7630,N_4556,N_1407);
or U7631 (N_7631,N_5337,N_2301);
xnor U7632 (N_7632,N_2024,N_3047);
or U7633 (N_7633,N_5263,N_6215);
nand U7634 (N_7634,N_3923,N_1313);
or U7635 (N_7635,N_3571,N_6236);
and U7636 (N_7636,N_3281,N_4442);
xnor U7637 (N_7637,N_1677,N_3123);
nand U7638 (N_7638,N_79,N_150);
xor U7639 (N_7639,N_1239,N_3135);
nand U7640 (N_7640,N_4002,N_1887);
or U7641 (N_7641,N_6089,N_2072);
xnor U7642 (N_7642,N_2253,N_456);
nand U7643 (N_7643,N_4659,N_1560);
nand U7644 (N_7644,N_5577,N_1129);
or U7645 (N_7645,N_3553,N_5866);
and U7646 (N_7646,N_1479,N_370);
xnor U7647 (N_7647,N_1639,N_5931);
nor U7648 (N_7648,N_1519,N_4816);
and U7649 (N_7649,N_3144,N_3080);
nand U7650 (N_7650,N_5584,N_3710);
nor U7651 (N_7651,N_3769,N_1386);
and U7652 (N_7652,N_5763,N_2585);
nor U7653 (N_7653,N_3151,N_503);
nor U7654 (N_7654,N_3729,N_3197);
or U7655 (N_7655,N_2131,N_6180);
nand U7656 (N_7656,N_2099,N_1082);
nand U7657 (N_7657,N_2866,N_1041);
nor U7658 (N_7658,N_11,N_5408);
or U7659 (N_7659,N_2279,N_768);
or U7660 (N_7660,N_206,N_5126);
nand U7661 (N_7661,N_1377,N_5436);
or U7662 (N_7662,N_513,N_3182);
nor U7663 (N_7663,N_1368,N_882);
xnor U7664 (N_7664,N_2231,N_2588);
nand U7665 (N_7665,N_3141,N_661);
or U7666 (N_7666,N_5063,N_516);
xnor U7667 (N_7667,N_1956,N_3388);
and U7668 (N_7668,N_3674,N_4879);
xnor U7669 (N_7669,N_962,N_1737);
and U7670 (N_7670,N_310,N_5459);
xor U7671 (N_7671,N_3477,N_2672);
xnor U7672 (N_7672,N_5047,N_2221);
nor U7673 (N_7673,N_4538,N_4946);
nor U7674 (N_7674,N_3577,N_1047);
nand U7675 (N_7675,N_5509,N_87);
or U7676 (N_7676,N_2721,N_3026);
nor U7677 (N_7677,N_4110,N_5428);
xnor U7678 (N_7678,N_44,N_1557);
xnor U7679 (N_7679,N_5253,N_2825);
nor U7680 (N_7680,N_1793,N_2377);
xnor U7681 (N_7681,N_3757,N_162);
nand U7682 (N_7682,N_612,N_2950);
and U7683 (N_7683,N_3420,N_4629);
and U7684 (N_7684,N_2919,N_1891);
xor U7685 (N_7685,N_1277,N_4298);
and U7686 (N_7686,N_1122,N_4087);
xnor U7687 (N_7687,N_520,N_5788);
or U7688 (N_7688,N_4247,N_5995);
nand U7689 (N_7689,N_3968,N_1884);
or U7690 (N_7690,N_3237,N_3091);
xnor U7691 (N_7691,N_1491,N_703);
nor U7692 (N_7692,N_5496,N_1100);
nor U7693 (N_7693,N_6123,N_2547);
or U7694 (N_7694,N_5090,N_1652);
and U7695 (N_7695,N_322,N_4724);
nor U7696 (N_7696,N_1686,N_1189);
xor U7697 (N_7697,N_3503,N_2119);
xnor U7698 (N_7698,N_158,N_6203);
nand U7699 (N_7699,N_4296,N_2106);
or U7700 (N_7700,N_182,N_1128);
nor U7701 (N_7701,N_1791,N_4730);
nand U7702 (N_7702,N_5193,N_2265);
and U7703 (N_7703,N_1564,N_3148);
or U7704 (N_7704,N_4643,N_1081);
and U7705 (N_7705,N_1679,N_60);
nand U7706 (N_7706,N_1424,N_5249);
nand U7707 (N_7707,N_5658,N_535);
nor U7708 (N_7708,N_1626,N_1873);
nand U7709 (N_7709,N_5587,N_2423);
or U7710 (N_7710,N_3536,N_3951);
nor U7711 (N_7711,N_809,N_5744);
and U7712 (N_7712,N_611,N_3015);
xnor U7713 (N_7713,N_4548,N_1585);
or U7714 (N_7714,N_2139,N_4417);
nand U7715 (N_7715,N_2371,N_4839);
nor U7716 (N_7716,N_3054,N_5317);
nand U7717 (N_7717,N_5776,N_5796);
nor U7718 (N_7718,N_5906,N_5668);
xor U7719 (N_7719,N_1503,N_6047);
or U7720 (N_7720,N_2720,N_3174);
nand U7721 (N_7721,N_2305,N_4945);
xnor U7722 (N_7722,N_4410,N_3550);
and U7723 (N_7723,N_848,N_2846);
and U7724 (N_7724,N_403,N_1960);
and U7725 (N_7725,N_3119,N_523);
nor U7726 (N_7726,N_6136,N_5712);
or U7727 (N_7727,N_3820,N_5138);
xor U7728 (N_7728,N_756,N_1778);
and U7729 (N_7729,N_5863,N_1536);
nor U7730 (N_7730,N_581,N_37);
xor U7731 (N_7731,N_5,N_466);
or U7732 (N_7732,N_3189,N_4225);
or U7733 (N_7733,N_1493,N_3689);
nor U7734 (N_7734,N_4050,N_782);
and U7735 (N_7735,N_872,N_5705);
xor U7736 (N_7736,N_4274,N_2104);
or U7737 (N_7737,N_2538,N_533);
nor U7738 (N_7738,N_3804,N_2658);
and U7739 (N_7739,N_5070,N_3025);
or U7740 (N_7740,N_5540,N_5910);
or U7741 (N_7741,N_1772,N_1346);
nor U7742 (N_7742,N_2991,N_5174);
xor U7743 (N_7743,N_3956,N_3540);
nor U7744 (N_7744,N_4215,N_4652);
and U7745 (N_7745,N_1281,N_887);
nand U7746 (N_7746,N_690,N_5617);
nand U7747 (N_7747,N_5291,N_4177);
nand U7748 (N_7748,N_2204,N_5647);
nand U7749 (N_7749,N_4130,N_4040);
xor U7750 (N_7750,N_2719,N_614);
xnor U7751 (N_7751,N_2864,N_5585);
nand U7752 (N_7752,N_2690,N_1247);
nor U7753 (N_7753,N_4188,N_6240);
and U7754 (N_7754,N_2968,N_3185);
nor U7755 (N_7755,N_3219,N_382);
and U7756 (N_7756,N_839,N_3308);
xnor U7757 (N_7757,N_5510,N_5123);
and U7758 (N_7758,N_1876,N_1266);
nor U7759 (N_7759,N_5305,N_2949);
and U7760 (N_7760,N_1250,N_4020);
nor U7761 (N_7761,N_5272,N_3944);
nor U7762 (N_7762,N_728,N_3414);
nand U7763 (N_7763,N_3691,N_841);
nor U7764 (N_7764,N_4310,N_5189);
and U7765 (N_7765,N_5450,N_267);
nor U7766 (N_7766,N_172,N_5406);
and U7767 (N_7767,N_5983,N_4435);
and U7768 (N_7768,N_1199,N_4696);
nand U7769 (N_7769,N_3002,N_66);
xor U7770 (N_7770,N_2102,N_4999);
xnor U7771 (N_7771,N_1326,N_863);
or U7772 (N_7772,N_3159,N_2254);
nor U7773 (N_7773,N_5304,N_5289);
nor U7774 (N_7774,N_4854,N_2532);
xnor U7775 (N_7775,N_3253,N_4702);
nand U7776 (N_7776,N_2142,N_480);
xor U7777 (N_7777,N_1141,N_3649);
nand U7778 (N_7778,N_2394,N_2771);
nand U7779 (N_7779,N_2141,N_3445);
nor U7780 (N_7780,N_3878,N_2008);
nor U7781 (N_7781,N_5360,N_4527);
nor U7782 (N_7782,N_5513,N_5008);
or U7783 (N_7783,N_5811,N_2794);
nand U7784 (N_7784,N_964,N_2865);
xnor U7785 (N_7785,N_4678,N_3753);
nor U7786 (N_7786,N_4614,N_1736);
or U7787 (N_7787,N_4315,N_3629);
and U7788 (N_7788,N_857,N_725);
xnor U7789 (N_7789,N_6081,N_5256);
and U7790 (N_7790,N_3639,N_1621);
nor U7791 (N_7791,N_3693,N_99);
nand U7792 (N_7792,N_802,N_6086);
or U7793 (N_7793,N_1321,N_1596);
xor U7794 (N_7794,N_2676,N_399);
xnor U7795 (N_7795,N_3217,N_4931);
and U7796 (N_7796,N_4670,N_81);
nor U7797 (N_7797,N_5605,N_1829);
or U7798 (N_7798,N_3656,N_918);
and U7799 (N_7799,N_3961,N_2201);
or U7800 (N_7800,N_1768,N_3315);
nor U7801 (N_7801,N_2671,N_3688);
or U7802 (N_7802,N_1868,N_2767);
xnor U7803 (N_7803,N_5366,N_3432);
xor U7804 (N_7804,N_2285,N_5000);
or U7805 (N_7805,N_6096,N_3865);
and U7806 (N_7806,N_2966,N_332);
nor U7807 (N_7807,N_2508,N_5800);
nand U7808 (N_7808,N_92,N_4682);
or U7809 (N_7809,N_453,N_1089);
nand U7810 (N_7810,N_1753,N_5128);
xnor U7811 (N_7811,N_2806,N_5583);
nor U7812 (N_7812,N_2597,N_3367);
or U7813 (N_7813,N_5902,N_5782);
xor U7814 (N_7814,N_4543,N_2336);
nor U7815 (N_7815,N_320,N_1376);
or U7816 (N_7816,N_5578,N_1214);
xor U7817 (N_7817,N_2175,N_704);
and U7818 (N_7818,N_521,N_4882);
nand U7819 (N_7819,N_5899,N_3412);
or U7820 (N_7820,N_5554,N_3748);
nor U7821 (N_7821,N_508,N_6031);
nor U7822 (N_7822,N_1912,N_5139);
nor U7823 (N_7823,N_3444,N_3578);
xor U7824 (N_7824,N_2505,N_1233);
nor U7825 (N_7825,N_1749,N_605);
or U7826 (N_7826,N_245,N_5006);
or U7827 (N_7827,N_4151,N_709);
and U7828 (N_7828,N_4727,N_1030);
xor U7829 (N_7829,N_5409,N_2980);
nand U7830 (N_7830,N_1773,N_4511);
nor U7831 (N_7831,N_5830,N_5077);
nand U7832 (N_7832,N_1532,N_2669);
xnor U7833 (N_7833,N_506,N_5528);
and U7834 (N_7834,N_4288,N_62);
xor U7835 (N_7835,N_386,N_4131);
nor U7836 (N_7836,N_4603,N_2368);
xor U7837 (N_7837,N_2603,N_1936);
and U7838 (N_7838,N_5129,N_5454);
or U7839 (N_7839,N_5246,N_898);
or U7840 (N_7840,N_4072,N_826);
nor U7841 (N_7841,N_6019,N_4056);
or U7842 (N_7842,N_3965,N_6036);
and U7843 (N_7843,N_5966,N_1678);
or U7844 (N_7844,N_3075,N_4437);
or U7845 (N_7845,N_4115,N_602);
and U7846 (N_7846,N_862,N_4835);
and U7847 (N_7847,N_4993,N_2773);
xor U7848 (N_7848,N_2788,N_5031);
and U7849 (N_7849,N_3316,N_25);
or U7850 (N_7850,N_2911,N_207);
and U7851 (N_7851,N_939,N_539);
nor U7852 (N_7852,N_563,N_2095);
or U7853 (N_7853,N_5567,N_1974);
nor U7854 (N_7854,N_2944,N_3736);
xor U7855 (N_7855,N_5385,N_4348);
nor U7856 (N_7856,N_3290,N_3964);
or U7857 (N_7857,N_2901,N_3647);
and U7858 (N_7858,N_427,N_742);
xnor U7859 (N_7859,N_6238,N_6077);
nor U7860 (N_7860,N_1689,N_1385);
nor U7861 (N_7861,N_5417,N_2384);
xor U7862 (N_7862,N_3920,N_5948);
xnor U7863 (N_7863,N_49,N_1851);
and U7864 (N_7864,N_524,N_5607);
and U7865 (N_7865,N_3224,N_3457);
and U7866 (N_7866,N_3293,N_699);
nand U7867 (N_7867,N_5377,N_3751);
nor U7868 (N_7868,N_4653,N_4322);
xor U7869 (N_7869,N_547,N_1661);
nand U7870 (N_7870,N_4299,N_1893);
nor U7871 (N_7871,N_4513,N_417);
and U7872 (N_7872,N_108,N_4889);
nand U7873 (N_7873,N_2763,N_1154);
and U7874 (N_7874,N_5968,N_6108);
and U7875 (N_7875,N_1526,N_3052);
or U7876 (N_7876,N_6101,N_865);
xnor U7877 (N_7877,N_2994,N_2962);
or U7878 (N_7878,N_266,N_3831);
and U7879 (N_7879,N_2506,N_1373);
nor U7880 (N_7880,N_5651,N_2784);
nor U7881 (N_7881,N_3921,N_144);
nor U7882 (N_7882,N_3166,N_4607);
nand U7883 (N_7883,N_5117,N_3742);
and U7884 (N_7884,N_2636,N_5880);
nor U7885 (N_7885,N_6088,N_3382);
and U7886 (N_7886,N_4103,N_229);
or U7887 (N_7887,N_5204,N_4430);
nand U7888 (N_7888,N_3717,N_873);
nor U7889 (N_7889,N_5755,N_1946);
xnor U7890 (N_7890,N_1021,N_3392);
xnor U7891 (N_7891,N_4981,N_623);
xor U7892 (N_7892,N_2220,N_5414);
nor U7893 (N_7893,N_1431,N_5853);
or U7894 (N_7894,N_3558,N_5514);
or U7895 (N_7895,N_621,N_5293);
nand U7896 (N_7896,N_306,N_2622);
xnor U7897 (N_7897,N_3568,N_6062);
xnor U7898 (N_7898,N_2718,N_1007);
nor U7899 (N_7899,N_5872,N_1322);
and U7900 (N_7900,N_454,N_3591);
nand U7901 (N_7901,N_3455,N_3456);
or U7902 (N_7902,N_4499,N_6020);
and U7903 (N_7903,N_5748,N_45);
and U7904 (N_7904,N_2329,N_4443);
and U7905 (N_7905,N_6050,N_4339);
nand U7906 (N_7906,N_5963,N_5725);
or U7907 (N_7907,N_1042,N_2482);
nand U7908 (N_7908,N_943,N_3515);
nand U7909 (N_7909,N_6205,N_4912);
xnor U7910 (N_7910,N_1967,N_5802);
or U7911 (N_7911,N_1465,N_1302);
xor U7912 (N_7912,N_1005,N_1695);
nor U7913 (N_7913,N_4827,N_1146);
nor U7914 (N_7914,N_1404,N_5687);
nand U7915 (N_7915,N_4588,N_1552);
xnor U7916 (N_7916,N_2529,N_4069);
nand U7917 (N_7917,N_6232,N_1977);
xor U7918 (N_7918,N_1317,N_3218);
nor U7919 (N_7919,N_5784,N_932);
xnor U7920 (N_7920,N_2751,N_2049);
and U7921 (N_7921,N_5180,N_2256);
nor U7922 (N_7922,N_3931,N_4910);
or U7923 (N_7923,N_5805,N_5153);
xor U7924 (N_7924,N_1808,N_6225);
and U7925 (N_7925,N_2548,N_1244);
xnor U7926 (N_7926,N_3668,N_2619);
and U7927 (N_7927,N_5407,N_1955);
and U7928 (N_7928,N_46,N_2510);
nand U7929 (N_7929,N_4633,N_1134);
nor U7930 (N_7930,N_6060,N_2022);
nor U7931 (N_7931,N_2148,N_3069);
and U7932 (N_7932,N_1730,N_3418);
or U7933 (N_7933,N_1461,N_2330);
nor U7934 (N_7934,N_3298,N_1104);
and U7935 (N_7935,N_4029,N_2315);
nor U7936 (N_7936,N_4487,N_1530);
nand U7937 (N_7937,N_344,N_3694);
or U7938 (N_7938,N_3811,N_3827);
nor U7939 (N_7939,N_2851,N_4531);
nor U7940 (N_7940,N_2999,N_2103);
nor U7941 (N_7941,N_1990,N_2039);
xor U7942 (N_7942,N_2958,N_2525);
xnor U7943 (N_7943,N_1455,N_3285);
or U7944 (N_7944,N_5412,N_5958);
xor U7945 (N_7945,N_4622,N_3303);
nor U7946 (N_7946,N_927,N_3177);
nand U7947 (N_7947,N_4962,N_5338);
nor U7948 (N_7948,N_153,N_3576);
and U7949 (N_7949,N_1838,N_4173);
nand U7950 (N_7950,N_1137,N_5842);
or U7951 (N_7951,N_358,N_5463);
and U7952 (N_7952,N_2960,N_1892);
and U7953 (N_7953,N_2899,N_2211);
nand U7954 (N_7954,N_5882,N_3737);
and U7955 (N_7955,N_5320,N_3130);
nor U7956 (N_7956,N_2654,N_6169);
xor U7957 (N_7957,N_3439,N_5478);
nand U7958 (N_7958,N_407,N_2013);
nor U7959 (N_7959,N_6051,N_1308);
or U7960 (N_7960,N_3180,N_5398);
nor U7961 (N_7961,N_1739,N_1853);
nand U7962 (N_7962,N_5394,N_5745);
nor U7963 (N_7963,N_4735,N_4763);
nor U7964 (N_7964,N_5779,N_1212);
nor U7965 (N_7965,N_4885,N_825);
and U7966 (N_7966,N_3059,N_1485);
or U7967 (N_7967,N_3085,N_451);
or U7968 (N_7968,N_1803,N_2564);
and U7969 (N_7969,N_5683,N_4660);
and U7970 (N_7970,N_2951,N_4061);
nand U7971 (N_7971,N_1729,N_3876);
xor U7972 (N_7972,N_3880,N_629);
nor U7973 (N_7973,N_1787,N_3625);
and U7974 (N_7974,N_2759,N_2356);
or U7975 (N_7975,N_3908,N_3708);
and U7976 (N_7976,N_3933,N_3211);
nand U7977 (N_7977,N_5841,N_6163);
nor U7978 (N_7978,N_3188,N_3982);
nor U7979 (N_7979,N_345,N_1483);
and U7980 (N_7980,N_4685,N_4292);
nand U7981 (N_7981,N_3063,N_2795);
xnor U7982 (N_7982,N_357,N_2504);
and U7983 (N_7983,N_2407,N_19);
and U7984 (N_7984,N_2556,N_5846);
nand U7985 (N_7985,N_3805,N_3607);
nand U7986 (N_7986,N_5218,N_1116);
nor U7987 (N_7987,N_5283,N_5225);
and U7988 (N_7988,N_2445,N_4530);
and U7989 (N_7989,N_1094,N_2686);
and U7990 (N_7990,N_2202,N_5258);
and U7991 (N_7991,N_5375,N_1767);
and U7992 (N_7992,N_1769,N_2109);
nor U7993 (N_7993,N_1048,N_3695);
and U7994 (N_7994,N_3306,N_2340);
nand U7995 (N_7995,N_4976,N_3830);
or U7996 (N_7996,N_4809,N_1333);
nand U7997 (N_7997,N_3108,N_4214);
or U7998 (N_7998,N_1909,N_3017);
nor U7999 (N_7999,N_990,N_2291);
and U8000 (N_8000,N_1740,N_1716);
and U8001 (N_8001,N_4041,N_5405);
nor U8002 (N_8002,N_5643,N_3232);
or U8003 (N_8003,N_3099,N_1340);
and U8004 (N_8004,N_5960,N_33);
nor U8005 (N_8005,N_5382,N_142);
nand U8006 (N_8006,N_5835,N_3685);
or U8007 (N_8007,N_5125,N_4964);
or U8008 (N_8008,N_2016,N_816);
nor U8009 (N_8009,N_5865,N_1004);
nor U8010 (N_8010,N_2059,N_4559);
nor U8011 (N_8011,N_4444,N_3036);
xnor U8012 (N_8012,N_4270,N_2700);
xor U8013 (N_8013,N_6179,N_1403);
or U8014 (N_8014,N_1609,N_5495);
or U8015 (N_8015,N_5718,N_5080);
nand U8016 (N_8016,N_696,N_4967);
and U8017 (N_8017,N_1717,N_4921);
or U8018 (N_8018,N_1359,N_4391);
nand U8019 (N_8019,N_3874,N_3760);
nand U8020 (N_8020,N_5456,N_140);
and U8021 (N_8021,N_2064,N_1181);
xor U8022 (N_8022,N_2151,N_1034);
nor U8023 (N_8023,N_5911,N_2722);
and U8024 (N_8024,N_5085,N_1524);
and U8025 (N_8025,N_1323,N_4396);
nand U8026 (N_8026,N_4038,N_1350);
nand U8027 (N_8027,N_4207,N_1265);
or U8028 (N_8028,N_1429,N_1201);
or U8029 (N_8029,N_5737,N_4232);
nand U8030 (N_8030,N_3385,N_1052);
or U8031 (N_8031,N_2343,N_1546);
xnor U8032 (N_8032,N_3541,N_579);
xnor U8033 (N_8033,N_3936,N_2344);
or U8034 (N_8034,N_6085,N_4273);
and U8035 (N_8035,N_3340,N_3703);
nand U8036 (N_8036,N_2060,N_4807);
xnor U8037 (N_8037,N_2450,N_4355);
or U8038 (N_8038,N_5488,N_2451);
or U8039 (N_8039,N_5448,N_875);
xnor U8040 (N_8040,N_5236,N_5481);
xnor U8041 (N_8041,N_4085,N_4514);
nand U8042 (N_8042,N_6211,N_3533);
or U8043 (N_8043,N_4409,N_1068);
nand U8044 (N_8044,N_1904,N_2012);
and U8045 (N_8045,N_868,N_5404);
xnor U8046 (N_8046,N_4475,N_2578);
nand U8047 (N_8047,N_1118,N_5442);
xor U8048 (N_8048,N_1268,N_5190);
or U8049 (N_8049,N_1731,N_269);
xnor U8050 (N_8050,N_5678,N_4674);
nand U8051 (N_8051,N_1545,N_4268);
and U8052 (N_8052,N_2224,N_5471);
nor U8053 (N_8053,N_1913,N_3618);
nor U8054 (N_8054,N_5992,N_96);
nor U8055 (N_8055,N_5743,N_2893);
nor U8056 (N_8056,N_47,N_5321);
or U8057 (N_8057,N_3110,N_3104);
or U8058 (N_8058,N_3822,N_1760);
nor U8059 (N_8059,N_2215,N_5893);
xor U8060 (N_8060,N_2476,N_3630);
or U8061 (N_8061,N_4752,N_3016);
and U8062 (N_8062,N_4797,N_4095);
xnor U8063 (N_8063,N_3555,N_3603);
nor U8064 (N_8064,N_4099,N_5573);
nand U8065 (N_8065,N_101,N_893);
nor U8066 (N_8066,N_1502,N_34);
nand U8067 (N_8067,N_2546,N_2888);
and U8068 (N_8068,N_4027,N_3847);
xor U8069 (N_8069,N_4474,N_124);
and U8070 (N_8070,N_1640,N_5827);
and U8071 (N_8071,N_903,N_5998);
nand U8072 (N_8072,N_5867,N_5808);
nor U8073 (N_8073,N_3124,N_2930);
nand U8074 (N_8074,N_4064,N_1980);
and U8075 (N_8075,N_3416,N_3252);
nor U8076 (N_8076,N_1959,N_4924);
and U8077 (N_8077,N_291,N_5439);
nor U8078 (N_8078,N_4754,N_3554);
nor U8079 (N_8079,N_4618,N_1062);
and U8080 (N_8080,N_2706,N_4454);
and U8081 (N_8081,N_6146,N_5905);
nand U8082 (N_8082,N_1489,N_3362);
xnor U8083 (N_8083,N_813,N_4036);
or U8084 (N_8084,N_4451,N_1917);
or U8085 (N_8085,N_3178,N_2606);
or U8086 (N_8086,N_5854,N_5594);
xnor U8087 (N_8087,N_5527,N_498);
nor U8088 (N_8088,N_2562,N_5205);
nand U8089 (N_8089,N_2177,N_5754);
and U8090 (N_8090,N_557,N_3046);
nor U8091 (N_8091,N_4804,N_5824);
nand U8092 (N_8092,N_365,N_2063);
or U8093 (N_8093,N_2873,N_5053);
or U8094 (N_8094,N_1166,N_3543);
and U8095 (N_8095,N_1076,N_2877);
xnor U8096 (N_8096,N_4896,N_5814);
xnor U8097 (N_8097,N_1965,N_1033);
xnor U8098 (N_8098,N_4279,N_1660);
xor U8099 (N_8099,N_4681,N_248);
nand U8100 (N_8100,N_4353,N_5815);
nor U8101 (N_8101,N_5280,N_3450);
nor U8102 (N_8102,N_2716,N_745);
nor U8103 (N_8103,N_827,N_5202);
xor U8104 (N_8104,N_2168,N_2761);
nor U8105 (N_8105,N_85,N_2410);
or U8106 (N_8106,N_4197,N_3890);
nand U8107 (N_8107,N_334,N_1303);
nor U8108 (N_8108,N_3464,N_1132);
and U8109 (N_8109,N_1384,N_559);
or U8110 (N_8110,N_4492,N_3200);
nand U8111 (N_8111,N_1077,N_2286);
and U8112 (N_8112,N_2238,N_4635);
nor U8113 (N_8113,N_1542,N_103);
nand U8114 (N_8114,N_5027,N_4733);
xnor U8115 (N_8115,N_440,N_552);
nand U8116 (N_8116,N_3486,N_1016);
and U8117 (N_8117,N_2038,N_3950);
or U8118 (N_8118,N_5252,N_715);
and U8119 (N_8119,N_2937,N_3114);
nor U8120 (N_8120,N_4216,N_1003);
nand U8121 (N_8121,N_630,N_3422);
nor U8122 (N_8122,N_617,N_645);
nor U8123 (N_8123,N_2682,N_5392);
xnor U8124 (N_8124,N_2228,N_3345);
nor U8125 (N_8125,N_2158,N_5878);
and U8126 (N_8126,N_28,N_1347);
nor U8127 (N_8127,N_830,N_1125);
nor U8128 (N_8128,N_4737,N_1908);
xor U8129 (N_8129,N_4054,N_1938);
nand U8130 (N_8130,N_0,N_596);
nand U8131 (N_8131,N_67,N_4359);
and U8132 (N_8132,N_685,N_3715);
or U8133 (N_8133,N_2982,N_3681);
or U8134 (N_8134,N_1097,N_2357);
xor U8135 (N_8135,N_2640,N_2838);
xnor U8136 (N_8136,N_2150,N_3249);
nor U8137 (N_8137,N_1601,N_1595);
and U8138 (N_8138,N_1226,N_1941);
nand U8139 (N_8139,N_356,N_5441);
nand U8140 (N_8140,N_4152,N_4980);
and U8141 (N_8141,N_2975,N_1486);
and U8142 (N_8142,N_2137,N_1825);
nor U8143 (N_8143,N_5606,N_2816);
and U8144 (N_8144,N_2755,N_2776);
and U8145 (N_8145,N_4767,N_5601);
and U8146 (N_8146,N_2687,N_317);
or U8147 (N_8147,N_2314,N_32);
and U8148 (N_8148,N_6044,N_3679);
xor U8149 (N_8149,N_3614,N_829);
or U8150 (N_8150,N_1319,N_3884);
and U8151 (N_8151,N_121,N_3129);
nor U8152 (N_8152,N_408,N_3209);
nand U8153 (N_8153,N_1310,N_707);
nor U8154 (N_8154,N_2823,N_945);
and U8155 (N_8155,N_5312,N_4460);
and U8156 (N_8156,N_1574,N_3793);
nor U8157 (N_8157,N_2732,N_6043);
and U8158 (N_8158,N_2260,N_2693);
nor U8159 (N_8159,N_5214,N_2948);
nand U8160 (N_8160,N_3617,N_5851);
nor U8161 (N_8161,N_4961,N_3260);
and U8162 (N_8162,N_2007,N_1949);
nor U8163 (N_8163,N_3896,N_2607);
nor U8164 (N_8164,N_3117,N_5550);
and U8165 (N_8165,N_5930,N_3734);
and U8166 (N_8166,N_6007,N_5211);
and U8167 (N_8167,N_3074,N_331);
and U8168 (N_8168,N_5274,N_257);
and U8169 (N_8169,N_2787,N_5700);
nand U8170 (N_8170,N_896,N_2984);
xor U8171 (N_8171,N_678,N_111);
nor U8172 (N_8172,N_5009,N_1522);
nand U8173 (N_8173,N_1196,N_6228);
nand U8174 (N_8174,N_529,N_5873);
nand U8175 (N_8175,N_2205,N_4505);
or U8176 (N_8176,N_1841,N_3037);
nor U8177 (N_8177,N_783,N_3347);
nand U8178 (N_8178,N_5029,N_5401);
nand U8179 (N_8179,N_4169,N_5010);
nand U8180 (N_8180,N_5492,N_2130);
and U8181 (N_8181,N_4493,N_6147);
nor U8182 (N_8182,N_5095,N_346);
xor U8183 (N_8183,N_321,N_891);
nand U8184 (N_8184,N_4820,N_307);
or U8185 (N_8185,N_5127,N_3264);
or U8186 (N_8186,N_818,N_4386);
and U8187 (N_8187,N_2845,N_1006);
or U8188 (N_8188,N_566,N_5938);
and U8189 (N_8189,N_1135,N_5413);
and U8190 (N_8190,N_6114,N_6042);
nor U8191 (N_8191,N_1401,N_842);
nor U8192 (N_8192,N_655,N_1926);
nand U8193 (N_8193,N_5590,N_5664);
nand U8194 (N_8194,N_3459,N_4129);
or U8195 (N_8195,N_3461,N_4594);
or U8196 (N_8196,N_1457,N_4362);
and U8197 (N_8197,N_2590,N_6002);
nor U8198 (N_8198,N_3716,N_2531);
and U8199 (N_8199,N_4158,N_643);
xnor U8200 (N_8200,N_1663,N_653);
nand U8201 (N_8201,N_4219,N_1334);
xnor U8202 (N_8202,N_2662,N_1366);
xnor U8203 (N_8203,N_5859,N_2856);
nand U8204 (N_8204,N_4154,N_1513);
nor U8205 (N_8205,N_3744,N_3999);
and U8206 (N_8206,N_4826,N_4053);
nor U8207 (N_8207,N_4778,N_5751);
nor U8208 (N_8208,N_6176,N_2118);
nor U8209 (N_8209,N_3662,N_1578);
xor U8210 (N_8210,N_4055,N_3024);
nand U8211 (N_8211,N_4226,N_1238);
nor U8212 (N_8212,N_1847,N_3743);
or U8213 (N_8213,N_2208,N_3895);
and U8214 (N_8214,N_400,N_4569);
nor U8215 (N_8215,N_3374,N_3511);
and U8216 (N_8216,N_65,N_6149);
or U8217 (N_8217,N_5212,N_381);
or U8218 (N_8218,N_2647,N_2957);
xor U8219 (N_8219,N_717,N_4621);
xnor U8220 (N_8220,N_5065,N_1828);
or U8221 (N_8221,N_1579,N_5724);
nand U8222 (N_8222,N_1009,N_1518);
xnor U8223 (N_8223,N_2651,N_1251);
xnor U8224 (N_8224,N_1365,N_3834);
or U8225 (N_8225,N_3403,N_2674);
xnor U8226 (N_8226,N_5132,N_5178);
and U8227 (N_8227,N_4747,N_584);
or U8228 (N_8228,N_3441,N_1682);
and U8229 (N_8229,N_6155,N_3502);
xor U8230 (N_8230,N_3949,N_4795);
or U8231 (N_8231,N_626,N_2031);
xnor U8232 (N_8232,N_1681,N_5168);
xor U8233 (N_8233,N_128,N_3913);
or U8234 (N_8234,N_3806,N_6166);
nor U8235 (N_8235,N_4832,N_710);
nand U8236 (N_8236,N_2926,N_663);
and U8237 (N_8237,N_5999,N_5547);
nand U8238 (N_8238,N_3140,N_422);
and U8239 (N_8239,N_225,N_5941);
xnor U8240 (N_8240,N_1906,N_4189);
and U8241 (N_8241,N_6186,N_3248);
and U8242 (N_8242,N_2454,N_1784);
and U8243 (N_8243,N_5355,N_1823);
or U8244 (N_8244,N_238,N_2480);
or U8245 (N_8245,N_2491,N_1691);
xnor U8246 (N_8246,N_666,N_1898);
xnor U8247 (N_8247,N_1506,N_4463);
nand U8248 (N_8248,N_1947,N_4262);
or U8249 (N_8249,N_3387,N_1856);
nor U8250 (N_8250,N_3487,N_4235);
xor U8251 (N_8251,N_3155,N_1406);
or U8252 (N_8252,N_3297,N_5135);
xnor U8253 (N_8253,N_3572,N_5106);
nor U8254 (N_8254,N_1454,N_5268);
nor U8255 (N_8255,N_23,N_2370);
and U8256 (N_8256,N_1228,N_5533);
xnor U8257 (N_8257,N_920,N_1061);
xnor U8258 (N_8258,N_1915,N_4971);
nand U8259 (N_8259,N_5329,N_718);
and U8260 (N_8260,N_2334,N_5817);
nand U8261 (N_8261,N_2289,N_4788);
nor U8262 (N_8262,N_5623,N_3991);
nand U8263 (N_8263,N_4963,N_2066);
nand U8264 (N_8264,N_1857,N_5630);
or U8265 (N_8265,N_283,N_5322);
nor U8266 (N_8266,N_1975,N_4111);
nor U8267 (N_8267,N_6209,N_2484);
xor U8268 (N_8268,N_5049,N_4251);
xnor U8269 (N_8269,N_3752,N_885);
or U8270 (N_8270,N_1994,N_722);
nand U8271 (N_8271,N_691,N_2895);
nor U8272 (N_8272,N_3537,N_5787);
or U8273 (N_8273,N_313,N_5316);
xnor U8274 (N_8274,N_3447,N_3527);
or U8275 (N_8275,N_2887,N_3470);
or U8276 (N_8276,N_4958,N_4113);
xnor U8277 (N_8277,N_3766,N_4366);
or U8278 (N_8278,N_216,N_1805);
nor U8279 (N_8279,N_3090,N_3431);
nor U8280 (N_8280,N_5447,N_3164);
and U8281 (N_8281,N_4490,N_485);
or U8282 (N_8282,N_2837,N_5953);
xor U8283 (N_8283,N_5887,N_1345);
and U8284 (N_8284,N_125,N_3985);
nand U8285 (N_8285,N_543,N_3953);
nor U8286 (N_8286,N_3643,N_4596);
and U8287 (N_8287,N_1866,N_5892);
nand U8288 (N_8288,N_1467,N_168);
and U8289 (N_8289,N_5111,N_5066);
and U8290 (N_8290,N_5959,N_2258);
or U8291 (N_8291,N_1701,N_985);
nor U8292 (N_8292,N_5508,N_5069);
or U8293 (N_8293,N_1962,N_1349);
xnor U8294 (N_8294,N_600,N_5631);
nand U8295 (N_8295,N_5536,N_5602);
and U8296 (N_8296,N_6226,N_3881);
xor U8297 (N_8297,N_3526,N_5970);
nand U8298 (N_8298,N_2047,N_639);
nor U8299 (N_8299,N_59,N_1698);
or U8300 (N_8300,N_5720,N_4453);
nand U8301 (N_8301,N_222,N_2282);
or U8302 (N_8302,N_419,N_2232);
nor U8303 (N_8303,N_3084,N_3508);
nand U8304 (N_8304,N_1978,N_4324);
xnor U8305 (N_8305,N_4175,N_5524);
nor U8306 (N_8306,N_244,N_1619);
and U8307 (N_8307,N_362,N_3621);
xor U8308 (N_8308,N_4764,N_21);
xnor U8309 (N_8309,N_5187,N_1213);
and U8310 (N_8310,N_2808,N_609);
and U8311 (N_8311,N_4920,N_634);
xnor U8312 (N_8312,N_3808,N_4694);
or U8313 (N_8313,N_1448,N_2587);
and U8314 (N_8314,N_6024,N_1744);
xor U8315 (N_8315,N_5402,N_3395);
and U8316 (N_8316,N_3828,N_3029);
or U8317 (N_8317,N_3988,N_3622);
nor U8318 (N_8318,N_1528,N_1343);
and U8319 (N_8319,N_1859,N_2804);
or U8320 (N_8320,N_2347,N_5483);
nor U8321 (N_8321,N_226,N_1589);
nor U8322 (N_8322,N_385,N_3018);
and U8323 (N_8323,N_3934,N_6199);
nor U8324 (N_8324,N_4679,N_1999);
xor U8325 (N_8325,N_2972,N_4071);
nor U8326 (N_8326,N_3423,N_2245);
or U8327 (N_8327,N_3954,N_1372);
nand U8328 (N_8328,N_5874,N_3381);
xor U8329 (N_8329,N_731,N_5985);
nand U8330 (N_8330,N_188,N_4000);
nor U8331 (N_8331,N_2796,N_5845);
xnor U8332 (N_8332,N_4540,N_953);
xor U8333 (N_8333,N_1920,N_4673);
or U8334 (N_8334,N_2448,N_341);
nor U8335 (N_8335,N_1804,N_3348);
xnor U8336 (N_8336,N_5028,N_2526);
nand U8337 (N_8337,N_2798,N_6183);
nand U8338 (N_8338,N_4013,N_5969);
xor U8339 (N_8339,N_479,N_4108);
xnor U8340 (N_8340,N_1880,N_4847);
nand U8341 (N_8341,N_2528,N_2741);
nand U8342 (N_8342,N_5549,N_3187);
and U8343 (N_8343,N_1951,N_1110);
nor U8344 (N_8344,N_743,N_4180);
nor U8345 (N_8345,N_2417,N_6190);
nand U8346 (N_8346,N_4502,N_1162);
nand U8347 (N_8347,N_4729,N_1413);
xor U8348 (N_8348,N_5363,N_5912);
or U8349 (N_8349,N_4445,N_2910);
nor U8350 (N_8350,N_1050,N_439);
nand U8351 (N_8351,N_853,N_4938);
nor U8352 (N_8352,N_3100,N_3535);
and U8353 (N_8353,N_3497,N_1078);
and U8354 (N_8354,N_3326,N_2361);
and U8355 (N_8355,N_4234,N_309);
and U8356 (N_8356,N_5255,N_6059);
xor U8357 (N_8357,N_5485,N_1193);
or U8358 (N_8358,N_1576,N_374);
nand U8359 (N_8359,N_2642,N_5742);
xnor U8360 (N_8360,N_1632,N_676);
nor U8361 (N_8361,N_3001,N_97);
xor U8362 (N_8362,N_527,N_4983);
nor U8363 (N_8363,N_3567,N_2312);
xor U8364 (N_8364,N_3642,N_5082);
nor U8365 (N_8365,N_2200,N_5971);
nor U8366 (N_8366,N_2112,N_2360);
nor U8367 (N_8367,N_4845,N_1644);
and U8368 (N_8368,N_2550,N_2432);
xor U8369 (N_8369,N_64,N_4828);
nand U8370 (N_8370,N_4848,N_2332);
or U8371 (N_8371,N_3371,N_4480);
and U8372 (N_8372,N_384,N_3809);
and U8373 (N_8373,N_2632,N_3781);
nor U8374 (N_8374,N_799,N_366);
or U8375 (N_8375,N_2001,N_3813);
xnor U8376 (N_8376,N_4901,N_1451);
xnor U8377 (N_8377,N_3987,N_4577);
and U8378 (N_8378,N_1235,N_3143);
nand U8379 (N_8379,N_2559,N_3120);
and U8380 (N_8380,N_4147,N_4381);
or U8381 (N_8381,N_2020,N_5747);
and U8382 (N_8382,N_6033,N_5790);
nand U8383 (N_8383,N_1221,N_4365);
and U8384 (N_8384,N_3268,N_4640);
nor U8385 (N_8385,N_411,N_1136);
and U8386 (N_8386,N_729,N_1724);
nor U8387 (N_8387,N_2255,N_984);
or U8388 (N_8388,N_2497,N_1151);
nor U8389 (N_8389,N_4316,N_18);
xnor U8390 (N_8390,N_2981,N_262);
and U8391 (N_8391,N_3027,N_5185);
nand U8392 (N_8392,N_5176,N_3608);
and U8393 (N_8393,N_1272,N_2913);
xnor U8394 (N_8394,N_3546,N_4450);
nor U8395 (N_8395,N_5290,N_1837);
nor U8396 (N_8396,N_194,N_3852);
xor U8397 (N_8397,N_2989,N_1656);
or U8398 (N_8398,N_6201,N_3935);
or U8399 (N_8399,N_3794,N_4623);
nor U8400 (N_8400,N_3581,N_5432);
and U8401 (N_8401,N_4522,N_279);
or U8402 (N_8402,N_5342,N_2057);
nor U8403 (N_8403,N_2089,N_4627);
or U8404 (N_8404,N_1458,N_1797);
xor U8405 (N_8405,N_1481,N_3996);
xnor U8406 (N_8406,N_2283,N_4294);
xor U8407 (N_8407,N_3419,N_1446);
and U8408 (N_8408,N_4726,N_4562);
or U8409 (N_8409,N_2539,N_3257);
nor U8410 (N_8410,N_2955,N_3869);
nor U8411 (N_8411,N_3512,N_3942);
nand U8412 (N_8412,N_3529,N_4766);
nor U8413 (N_8413,N_4186,N_4647);
or U8414 (N_8414,N_4438,N_5223);
or U8415 (N_8415,N_1885,N_256);
nand U8416 (N_8416,N_4915,N_1620);
nor U8417 (N_8417,N_1790,N_2017);
nor U8418 (N_8418,N_795,N_5749);
and U8419 (N_8419,N_4051,N_5644);
xnor U8420 (N_8420,N_555,N_4278);
xnor U8421 (N_8421,N_1,N_4172);
and U8422 (N_8422,N_4741,N_57);
nand U8423 (N_8423,N_1133,N_3373);
nand U8424 (N_8424,N_5278,N_3405);
or U8425 (N_8425,N_280,N_5620);
nand U8426 (N_8426,N_5387,N_5762);
nand U8427 (N_8427,N_3705,N_5781);
xnor U8428 (N_8428,N_1770,N_1445);
or U8429 (N_8429,N_5746,N_3867);
nand U8430 (N_8430,N_2791,N_13);
xor U8431 (N_8431,N_3556,N_3838);
nand U8432 (N_8432,N_2230,N_1964);
xor U8433 (N_8433,N_3032,N_1813);
or U8434 (N_8434,N_1357,N_4563);
nand U8435 (N_8435,N_677,N_4193);
xor U8436 (N_8436,N_5654,N_3745);
xnor U8437 (N_8437,N_147,N_4255);
nand U8438 (N_8438,N_5728,N_761);
nand U8439 (N_8439,N_641,N_1119);
and U8440 (N_8440,N_2061,N_1452);
nand U8441 (N_8441,N_35,N_719);
nor U8442 (N_8442,N_1301,N_2194);
nor U8443 (N_8443,N_1351,N_1858);
nand U8444 (N_8444,N_3269,N_667);
xnor U8445 (N_8445,N_4479,N_4312);
nand U8446 (N_8446,N_3318,N_435);
nand U8447 (N_8447,N_289,N_3641);
and U8448 (N_8448,N_5684,N_1970);
or U8449 (N_8449,N_1713,N_2935);
nor U8450 (N_8450,N_2734,N_3116);
xor U8451 (N_8451,N_5563,N_2978);
and U8452 (N_8452,N_5101,N_16);
nand U8453 (N_8453,N_410,N_2641);
xor U8454 (N_8454,N_1447,N_3684);
and U8455 (N_8455,N_5423,N_3313);
nand U8456 (N_8456,N_2405,N_2625);
xor U8457 (N_8457,N_2216,N_2338);
nor U8458 (N_8458,N_5778,N_2473);
or U8459 (N_8459,N_5092,N_4620);
and U8460 (N_8460,N_5772,N_2153);
and U8461 (N_8461,N_4568,N_3295);
nand U8462 (N_8462,N_223,N_4088);
nand U8463 (N_8463,N_1383,N_922);
and U8464 (N_8464,N_4412,N_688);
xnor U8465 (N_8465,N_2519,N_3969);
or U8466 (N_8466,N_3471,N_4780);
nand U8467 (N_8467,N_433,N_2770);
or U8468 (N_8468,N_1482,N_5067);
or U8469 (N_8469,N_4567,N_5165);
nand U8470 (N_8470,N_1188,N_5704);
and U8471 (N_8471,N_3516,N_5045);
xnor U8472 (N_8472,N_2656,N_401);
nand U8473 (N_8473,N_914,N_6107);
xnor U8474 (N_8474,N_4865,N_5558);
nand U8475 (N_8475,N_1336,N_1032);
nand U8476 (N_8476,N_6135,N_4507);
nor U8477 (N_8477,N_1020,N_6061);
nor U8478 (N_8478,N_1390,N_4898);
or U8479 (N_8479,N_3873,N_3738);
and U8480 (N_8480,N_1298,N_438);
nand U8481 (N_8481,N_4222,N_2280);
nand U8482 (N_8482,N_1720,N_2872);
xor U8483 (N_8483,N_3251,N_2308);
or U8484 (N_8484,N_3173,N_6200);
xnor U8485 (N_8485,N_3138,N_6165);
and U8486 (N_8486,N_2534,N_604);
xnor U8487 (N_8487,N_2592,N_934);
xor U8488 (N_8488,N_5832,N_2084);
and U8489 (N_8489,N_2302,N_2346);
nand U8490 (N_8490,N_949,N_5943);
and U8491 (N_8491,N_445,N_5900);
nor U8492 (N_8492,N_1209,N_6241);
nand U8493 (N_8493,N_3664,N_5978);
xor U8494 (N_8494,N_4018,N_354);
and U8495 (N_8495,N_4892,N_6119);
nand U8496 (N_8496,N_2848,N_1896);
nand U8497 (N_8497,N_1580,N_1544);
nor U8498 (N_8498,N_548,N_1774);
nor U8499 (N_8499,N_1175,N_409);
or U8500 (N_8500,N_2917,N_471);
or U8501 (N_8501,N_1996,N_849);
xnor U8502 (N_8502,N_4404,N_1684);
nand U8503 (N_8503,N_5836,N_4258);
and U8504 (N_8504,N_493,N_1501);
and U8505 (N_8505,N_3605,N_5670);
xnor U8506 (N_8506,N_314,N_5173);
and U8507 (N_8507,N_4583,N_4744);
nor U8508 (N_8508,N_6167,N_2108);
xor U8509 (N_8509,N_4238,N_3995);
and U8510 (N_8510,N_2752,N_4648);
or U8511 (N_8511,N_2915,N_218);
xor U8512 (N_8512,N_55,N_5287);
xor U8513 (N_8513,N_328,N_5269);
or U8514 (N_8514,N_4428,N_5158);
and U8515 (N_8515,N_1381,N_5927);
xor U8516 (N_8516,N_6140,N_4609);
nand U8517 (N_8517,N_4604,N_180);
or U8518 (N_8518,N_3149,N_1364);
xnor U8519 (N_8519,N_3911,N_582);
or U8520 (N_8520,N_3955,N_2400);
or U8521 (N_8521,N_1995,N_1305);
nor U8522 (N_8522,N_452,N_3043);
and U8523 (N_8523,N_4749,N_1931);
xor U8524 (N_8524,N_3096,N_389);
nand U8525 (N_8525,N_316,N_5297);
or U8526 (N_8526,N_3698,N_355);
or U8527 (N_8527,N_5553,N_1073);
or U8528 (N_8528,N_4542,N_960);
or U8529 (N_8529,N_1014,N_4906);
or U8530 (N_8530,N_74,N_871);
xnor U8531 (N_8531,N_2631,N_4237);
and U8532 (N_8532,N_3003,N_4798);
and U8533 (N_8533,N_1688,N_2797);
nand U8534 (N_8534,N_6218,N_4844);
and U8535 (N_8535,N_5706,N_1113);
and U8536 (N_8536,N_5708,N_2742);
or U8537 (N_8537,N_4083,N_398);
and U8538 (N_8538,N_3448,N_4231);
nor U8539 (N_8539,N_5055,N_5041);
or U8540 (N_8540,N_4731,N_1102);
nand U8541 (N_8541,N_4761,N_4605);
nand U8542 (N_8542,N_4346,N_5013);
xnor U8543 (N_8543,N_528,N_4575);
xnor U8544 (N_8544,N_5653,N_4464);
or U8545 (N_8545,N_2132,N_5682);
xnor U8546 (N_8546,N_3300,N_652);
xnor U8547 (N_8547,N_981,N_3336);
nor U8548 (N_8548,N_5534,N_5932);
nand U8549 (N_8549,N_2350,N_4770);
nand U8550 (N_8550,N_1389,N_5955);
or U8551 (N_8551,N_5834,N_424);
xnor U8552 (N_8552,N_1271,N_894);
and U8553 (N_8553,N_2600,N_3028);
nand U8554 (N_8554,N_3925,N_736);
or U8555 (N_8555,N_3073,N_4389);
nand U8556 (N_8556,N_4917,N_3807);
xor U8557 (N_8557,N_3460,N_3759);
and U8558 (N_8558,N_5334,N_2275);
and U8559 (N_8559,N_5308,N_2996);
nand U8560 (N_8560,N_77,N_3203);
xnor U8561 (N_8561,N_5425,N_3754);
xor U8562 (N_8562,N_2733,N_3299);
nor U8563 (N_8563,N_1743,N_2943);
or U8564 (N_8564,N_470,N_5365);
or U8565 (N_8565,N_4043,N_2386);
or U8566 (N_8566,N_6243,N_167);
nand U8567 (N_8567,N_5752,N_1883);
nor U8568 (N_8568,N_982,N_2618);
or U8569 (N_8569,N_1755,N_2169);
xor U8570 (N_8570,N_12,N_3914);
xnor U8571 (N_8571,N_5548,N_765);
or U8572 (N_8572,N_10,N_1939);
nand U8573 (N_8573,N_1023,N_3309);
or U8574 (N_8574,N_4320,N_3530);
xor U8575 (N_8575,N_5131,N_472);
and U8576 (N_8576,N_5816,N_5939);
nor U8577 (N_8577,N_1324,N_3184);
nor U8578 (N_8578,N_2518,N_4508);
or U8579 (N_8579,N_5947,N_5753);
xnor U8580 (N_8580,N_4471,N_3707);
nand U8581 (N_8581,N_5677,N_4890);
nand U8582 (N_8582,N_4489,N_36);
or U8583 (N_8583,N_3658,N_2907);
and U8584 (N_8584,N_5389,N_3078);
and U8585 (N_8585,N_2397,N_5400);
or U8586 (N_8586,N_712,N_3646);
nor U8587 (N_8587,N_2817,N_4392);
nand U8588 (N_8588,N_2181,N_4318);
nand U8589 (N_8589,N_5120,N_4313);
nand U8590 (N_8590,N_4875,N_2612);
nand U8591 (N_8591,N_3826,N_4965);
or U8592 (N_8592,N_5195,N_6137);
and U8593 (N_8593,N_3803,N_4246);
or U8594 (N_8594,N_5881,N_5982);
or U8595 (N_8595,N_3009,N_4817);
xnor U8596 (N_8596,N_2544,N_2902);
and U8597 (N_8597,N_406,N_6090);
nand U8598 (N_8598,N_339,N_5956);
nand U8599 (N_8599,N_6122,N_6197);
xor U8600 (N_8600,N_5391,N_4159);
or U8601 (N_8601,N_6157,N_4067);
and U8602 (N_8602,N_1515,N_271);
nor U8603 (N_8603,N_915,N_5493);
or U8604 (N_8604,N_892,N_1393);
and U8605 (N_8605,N_1935,N_284);
xnor U8606 (N_8606,N_538,N_3265);
and U8607 (N_8607,N_2483,N_4712);
or U8608 (N_8608,N_5351,N_4972);
or U8609 (N_8609,N_2743,N_42);
and U8610 (N_8610,N_5565,N_4434);
or U8611 (N_8611,N_93,N_5052);
nand U8612 (N_8612,N_2159,N_5542);
nand U8613 (N_8613,N_644,N_1852);
xnor U8614 (N_8614,N_1142,N_4352);
xnor U8615 (N_8615,N_700,N_6171);
xor U8616 (N_8616,N_5904,N_3107);
nand U8617 (N_8617,N_1304,N_2299);
xnor U8618 (N_8618,N_5633,N_1631);
and U8619 (N_8619,N_136,N_5660);
xor U8620 (N_8620,N_2617,N_1820);
nand U8621 (N_8621,N_5059,N_4008);
nor U8622 (N_8622,N_570,N_902);
xnor U8623 (N_8623,N_4360,N_123);
xnor U8624 (N_8624,N_3966,N_3589);
xor U8625 (N_8625,N_4645,N_312);
nand U8626 (N_8626,N_2916,N_3937);
nand U8627 (N_8627,N_1311,N_3071);
nand U8628 (N_8628,N_5224,N_1734);
and U8629 (N_8629,N_4553,N_3404);
xor U8630 (N_8630,N_6056,N_3587);
nor U8631 (N_8631,N_1008,N_4539);
or U8632 (N_8632,N_2019,N_1230);
nand U8633 (N_8633,N_5639,N_5370);
and U8634 (N_8634,N_2447,N_5914);
and U8635 (N_8635,N_4824,N_4545);
xor U8636 (N_8636,N_888,N_276);
nand U8637 (N_8637,N_2415,N_1106);
and U8638 (N_8638,N_3193,N_1123);
nand U8639 (N_8639,N_1671,N_3670);
xnor U8640 (N_8640,N_1084,N_748);
or U8641 (N_8641,N_4452,N_4734);
and U8642 (N_8642,N_199,N_1718);
xnor U8643 (N_8643,N_1264,N_6038);
nand U8644 (N_8644,N_474,N_2849);
or U8645 (N_8645,N_674,N_662);
nor U8646 (N_8646,N_1259,N_2818);
nor U8647 (N_8647,N_5411,N_4799);
and U8648 (N_8648,N_4944,N_2318);
or U8649 (N_8649,N_814,N_772);
xnor U8650 (N_8650,N_3356,N_1839);
nand U8651 (N_8651,N_2367,N_4007);
or U8652 (N_8652,N_6112,N_1925);
or U8653 (N_8653,N_1283,N_3101);
and U8654 (N_8654,N_228,N_4672);
nand U8655 (N_8655,N_693,N_909);
and U8656 (N_8656,N_463,N_5445);
and U8657 (N_8657,N_502,N_4022);
nor U8658 (N_8658,N_3906,N_5446);
xor U8659 (N_8659,N_706,N_1510);
or U8660 (N_8660,N_3127,N_1160);
nand U8661 (N_8661,N_138,N_2378);
nor U8662 (N_8662,N_3246,N_5221);
and U8663 (N_8663,N_867,N_4573);
or U8664 (N_8664,N_2088,N_1879);
and U8665 (N_8665,N_6210,N_4308);
and U8666 (N_8666,N_2040,N_965);
nand U8667 (N_8667,N_4411,N_1427);
and U8668 (N_8668,N_2862,N_1788);
and U8669 (N_8669,N_1355,N_4344);
xnor U8670 (N_8670,N_4252,N_1497);
and U8671 (N_8671,N_4456,N_3437);
nor U8672 (N_8672,N_1577,N_3064);
nor U8673 (N_8673,N_1600,N_6110);
xor U8674 (N_8674,N_1314,N_1028);
and U8675 (N_8675,N_1278,N_1224);
xor U8676 (N_8676,N_5711,N_1933);
or U8677 (N_8677,N_4566,N_4496);
nand U8678 (N_8678,N_2810,N_4557);
xnor U8679 (N_8679,N_1864,N_5692);
nor U8680 (N_8680,N_994,N_1138);
xnor U8681 (N_8681,N_3199,N_1275);
and U8682 (N_8682,N_1504,N_4138);
or U8683 (N_8683,N_3095,N_2860);
nand U8684 (N_8684,N_2184,N_1861);
xor U8685 (N_8685,N_6158,N_2854);
and U8686 (N_8686,N_509,N_2331);
nor U8687 (N_8687,N_3321,N_1807);
nor U8688 (N_8688,N_3262,N_5110);
nand U8689 (N_8689,N_798,N_2879);
nand U8690 (N_8690,N_6247,N_9);
nand U8691 (N_8691,N_3408,N_1463);
and U8692 (N_8692,N_1159,N_325);
xnor U8693 (N_8693,N_5993,N_5535);
and U8694 (N_8694,N_776,N_5672);
nand U8695 (N_8695,N_5288,N_1402);
or U8696 (N_8696,N_6095,N_4001);
xor U8697 (N_8697,N_1834,N_1988);
nand U8698 (N_8698,N_3532,N_5688);
xnor U8699 (N_8699,N_3816,N_1846);
and U8700 (N_8700,N_4122,N_6118);
and U8701 (N_8701,N_1587,N_970);
nand U8702 (N_8702,N_443,N_6054);
nand U8703 (N_8703,N_2502,N_3194);
and U8704 (N_8704,N_1420,N_5539);
nor U8705 (N_8705,N_831,N_6134);
or U8706 (N_8706,N_3481,N_4592);
nor U8707 (N_8707,N_5994,N_1152);
nor U8708 (N_8708,N_2786,N_2977);
nand U8709 (N_8709,N_1817,N_3559);
nand U8710 (N_8710,N_14,N_395);
or U8711 (N_8711,N_1664,N_5489);
and U8712 (N_8712,N_721,N_1286);
xnor U8713 (N_8713,N_4899,N_5243);
nor U8714 (N_8714,N_5050,N_1973);
and U8715 (N_8715,N_4338,N_4383);
nor U8716 (N_8716,N_4330,N_5323);
nand U8717 (N_8717,N_5208,N_3616);
nor U8718 (N_8718,N_3042,N_1273);
and U8719 (N_8719,N_2212,N_5475);
xnor U8720 (N_8720,N_5934,N_929);
and U8721 (N_8721,N_2025,N_724);
or U8722 (N_8722,N_3731,N_851);
or U8723 (N_8723,N_610,N_622);
and U8724 (N_8724,N_5592,N_467);
nand U8725 (N_8725,N_5393,N_1950);
nor U8726 (N_8726,N_838,N_2691);
nor U8727 (N_8727,N_1411,N_4955);
or U8728 (N_8728,N_3012,N_5922);
xor U8729 (N_8729,N_3978,N_5839);
and U8730 (N_8730,N_1862,N_3335);
and U8731 (N_8731,N_5296,N_5604);
or U8732 (N_8732,N_3088,N_2404);
xor U8733 (N_8733,N_1147,N_654);
xnor U8734 (N_8734,N_3504,N_416);
xnor U8735 (N_8735,N_2379,N_253);
or U8736 (N_8736,N_2408,N_5062);
or U8737 (N_8737,N_4424,N_1331);
nand U8738 (N_8738,N_3234,N_1655);
xnor U8739 (N_8739,N_793,N_801);
xnor U8740 (N_8740,N_2871,N_2322);
or U8741 (N_8741,N_4700,N_4495);
xnor U8742 (N_8742,N_2847,N_3352);
nand U8743 (N_8743,N_5144,N_3762);
nor U8744 (N_8744,N_6224,N_4265);
xnor U8745 (N_8745,N_2441,N_1027);
nand U8746 (N_8746,N_2840,N_4290);
nor U8747 (N_8747,N_2769,N_4021);
nand U8748 (N_8748,N_5532,N_2069);
or U8749 (N_8749,N_4004,N_4427);
or U8750 (N_8750,N_3267,N_4230);
or U8751 (N_8751,N_3842,N_3247);
nor U8752 (N_8752,N_4520,N_1341);
and U8753 (N_8753,N_6030,N_2987);
or U8754 (N_8754,N_340,N_3797);
nor U8755 (N_8755,N_4503,N_2998);
and U8756 (N_8756,N_2462,N_2940);
and U8757 (N_8757,N_202,N_5124);
xor U8758 (N_8758,N_4484,N_6125);
nor U8759 (N_8759,N_2382,N_5415);
or U8760 (N_8760,N_477,N_1085);
or U8761 (N_8761,N_274,N_4483);
xnor U8762 (N_8762,N_5465,N_3204);
or U8763 (N_8763,N_4792,N_692);
nand U8764 (N_8764,N_6178,N_5096);
nor U8765 (N_8765,N_819,N_3941);
and U8766 (N_8766,N_4031,N_239);
nand U8767 (N_8767,N_2750,N_3215);
nor U8768 (N_8768,N_4779,N_5152);
nor U8769 (N_8769,N_488,N_1375);
nor U8770 (N_8770,N_5226,N_3292);
and U8771 (N_8771,N_564,N_1352);
and U8772 (N_8772,N_4314,N_850);
or U8773 (N_8773,N_5977,N_5621);
and U8774 (N_8774,N_3959,N_2774);
nand U8775 (N_8775,N_2080,N_3560);
or U8776 (N_8776,N_1735,N_2697);
nor U8777 (N_8777,N_3739,N_1881);
or U8778 (N_8778,N_4929,N_4868);
or U8779 (N_8779,N_3319,N_4819);
or U8780 (N_8780,N_2353,N_5650);
or U8781 (N_8781,N_5014,N_836);
nor U8782 (N_8782,N_3089,N_1010);
and U8783 (N_8783,N_1759,N_671);
xnor U8784 (N_8784,N_5582,N_1761);
xnor U8785 (N_8785,N_1979,N_4900);
and U8786 (N_8786,N_3628,N_869);
and U8787 (N_8787,N_1742,N_4613);
xnor U8788 (N_8788,N_3223,N_5869);
nor U8789 (N_8789,N_1441,N_109);
nand U8790 (N_8790,N_148,N_3992);
xnor U8791 (N_8791,N_1391,N_3361);
xnor U8792 (N_8792,N_2114,N_63);
nor U8793 (N_8793,N_2885,N_2041);
nor U8794 (N_8794,N_5740,N_1583);
or U8795 (N_8795,N_4774,N_5667);
nor U8796 (N_8796,N_656,N_5281);
xnor U8797 (N_8797,N_560,N_5614);
nand U8798 (N_8798,N_5825,N_304);
and U8799 (N_8799,N_2113,N_130);
or U8800 (N_8800,N_2176,N_261);
xnor U8801 (N_8801,N_5331,N_469);
xor U8802 (N_8802,N_5613,N_3798);
nor U8803 (N_8803,N_3122,N_490);
and U8804 (N_8804,N_797,N_4121);
nor U8805 (N_8805,N_5693,N_4691);
nand U8806 (N_8806,N_2442,N_5076);
nand U8807 (N_8807,N_2891,N_3886);
nor U8808 (N_8808,N_255,N_6208);
xor U8809 (N_8809,N_803,N_2807);
and U8810 (N_8810,N_744,N_2785);
or U8811 (N_8811,N_659,N_31);
and U8812 (N_8812,N_4525,N_4641);
or U8813 (N_8813,N_905,N_1634);
nand U8814 (N_8814,N_4601,N_149);
nor U8815 (N_8815,N_4107,N_669);
nor U8816 (N_8816,N_476,N_4725);
and U8817 (N_8817,N_5794,N_5100);
and U8818 (N_8818,N_726,N_4100);
nor U8819 (N_8819,N_329,N_5240);
xor U8820 (N_8820,N_3549,N_4695);
xnor U8821 (N_8821,N_1164,N_2311);
and U8822 (N_8822,N_1765,N_1667);
and U8823 (N_8823,N_4510,N_3210);
xnor U8824 (N_8824,N_3631,N_4599);
nor U8825 (N_8825,N_4842,N_837);
nor U8826 (N_8826,N_4123,N_6159);
nor U8827 (N_8827,N_5234,N_2586);
or U8828 (N_8828,N_5474,N_3256);
nor U8829 (N_8829,N_2218,N_2540);
and U8830 (N_8830,N_3776,N_132);
nor U8831 (N_8831,N_4217,N_2627);
or U8832 (N_8832,N_3449,N_4211);
and U8833 (N_8833,N_3783,N_1379);
xor U8834 (N_8834,N_319,N_6142);
xnor U8835 (N_8835,N_1822,N_1202);
nand U8836 (N_8836,N_2694,N_6198);
xor U8837 (N_8837,N_698,N_4114);
or U8838 (N_8838,N_3659,N_5154);
or U8839 (N_8839,N_3482,N_3391);
nand U8840 (N_8840,N_58,N_1517);
xnor U8841 (N_8841,N_2437,N_2474);
or U8842 (N_8842,N_2517,N_5555);
xnor U8843 (N_8843,N_4248,N_2820);
xor U8844 (N_8844,N_1930,N_504);
or U8845 (N_8845,N_1185,N_1280);
and U8846 (N_8846,N_3986,N_2180);
and U8847 (N_8847,N_5694,N_2657);
nor U8848 (N_8848,N_5951,N_3728);
or U8849 (N_8849,N_2426,N_4127);
or U8850 (N_8850,N_5336,N_5768);
nor U8851 (N_8851,N_375,N_4376);
or U8852 (N_8852,N_4354,N_5374);
nor U8853 (N_8853,N_3856,N_4397);
nor U8854 (N_8854,N_828,N_4094);
or U8855 (N_8855,N_2675,N_963);
nand U8856 (N_8856,N_4446,N_1222);
nand U8857 (N_8857,N_4630,N_2604);
nor U8858 (N_8858,N_992,N_2455);
and U8859 (N_8859,N_3402,N_2979);
and U8860 (N_8860,N_901,N_4374);
xor U8861 (N_8861,N_2976,N_4536);
nand U8862 (N_8862,N_3413,N_5722);
and U8863 (N_8863,N_3997,N_2832);
nor U8864 (N_8864,N_116,N_1325);
and U8865 (N_8865,N_2974,N_3500);
xnor U8866 (N_8866,N_2509,N_3721);
and U8867 (N_8867,N_3552,N_3483);
or U8868 (N_8868,N_3557,N_5264);
xnor U8869 (N_8869,N_635,N_2595);
nor U8870 (N_8870,N_1206,N_2762);
nand U8871 (N_8871,N_4723,N_821);
xor U8872 (N_8872,N_3311,N_1171);
nand U8873 (N_8873,N_5823,N_3314);
xor U8874 (N_8874,N_5457,N_6079);
nand U8875 (N_8875,N_3020,N_210);
nand U8876 (N_8876,N_553,N_4282);
nand U8877 (N_8877,N_5561,N_3390);
or U8878 (N_8878,N_4667,N_4713);
nor U8879 (N_8879,N_1565,N_2609);
nand U8880 (N_8880,N_4829,N_769);
or U8881 (N_8881,N_3939,N_3225);
xnor U8882 (N_8882,N_4494,N_3051);
xor U8883 (N_8883,N_4706,N_4950);
or U8884 (N_8884,N_2744,N_5015);
nor U8885 (N_8885,N_2882,N_3829);
nand U8886 (N_8886,N_931,N_3666);
nor U8887 (N_8887,N_1745,N_3900);
nor U8888 (N_8888,N_1659,N_5570);
and U8889 (N_8889,N_2802,N_805);
xnor U8890 (N_8890,N_3814,N_5543);
nor U8891 (N_8891,N_4052,N_859);
or U8892 (N_8892,N_2424,N_1875);
and U8893 (N_8893,N_928,N_5064);
nor U8894 (N_8894,N_5933,N_3885);
nor U8895 (N_8895,N_2819,N_4285);
nand U8896 (N_8896,N_380,N_3383);
nand U8897 (N_8897,N_1139,N_5275);
and U8898 (N_8898,N_5942,N_4541);
and U8899 (N_8899,N_3206,N_3930);
or U8900 (N_8900,N_3667,N_2906);
or U8901 (N_8901,N_3672,N_436);
nor U8902 (N_8902,N_2234,N_5419);
xor U8903 (N_8903,N_1569,N_4205);
nor U8904 (N_8904,N_5073,N_1035);
xnor U8905 (N_8905,N_143,N_3565);
xor U8906 (N_8906,N_4657,N_633);
nor U8907 (N_8907,N_5038,N_405);
or U8908 (N_8908,N_446,N_1919);
or U8909 (N_8909,N_1575,N_4336);
nand U8910 (N_8910,N_2161,N_1022);
and U8911 (N_8911,N_3000,N_5987);
or U8912 (N_8912,N_3186,N_870);
nand U8913 (N_8913,N_5913,N_4005);
and U8914 (N_8914,N_227,N_1549);
xor U8915 (N_8915,N_5094,N_3946);
nand U8916 (N_8916,N_6021,N_4156);
or U8917 (N_8917,N_303,N_6035);
nor U8918 (N_8918,N_4357,N_2278);
nor U8919 (N_8919,N_6109,N_2637);
or U8920 (N_8920,N_5877,N_5294);
or U8921 (N_8921,N_2042,N_2248);
nor U8922 (N_8922,N_6249,N_4591);
or U8923 (N_8923,N_5929,N_2569);
and U8924 (N_8924,N_2573,N_5926);
xor U8925 (N_8925,N_1854,N_3213);
and U8926 (N_8926,N_2246,N_258);
nand U8927 (N_8927,N_3398,N_5537);
or U8928 (N_8928,N_1396,N_2100);
nand U8929 (N_8929,N_2839,N_2723);
or U8930 (N_8930,N_3675,N_5122);
xnor U8931 (N_8931,N_2374,N_2321);
and U8932 (N_8932,N_968,N_1320);
xnor U8933 (N_8933,N_1943,N_2789);
nand U8934 (N_8934,N_4762,N_3393);
nand U8935 (N_8935,N_4384,N_3278);
or U8936 (N_8936,N_1074,N_1777);
or U8937 (N_8937,N_2869,N_2116);
or U8938 (N_8938,N_2396,N_1976);
nor U8939 (N_8939,N_4291,N_495);
xnor U8940 (N_8940,N_2644,N_1075);
and U8941 (N_8941,N_4579,N_577);
xnor U8942 (N_8942,N_5699,N_1900);
or U8943 (N_8943,N_3093,N_5108);
or U8944 (N_8944,N_4600,N_5919);
or U8945 (N_8945,N_169,N_5350);
and U8946 (N_8946,N_1733,N_5719);
or U8947 (N_8947,N_4209,N_5562);
and U8948 (N_8948,N_895,N_6177);
nor U8949 (N_8949,N_6099,N_5807);
nand U8950 (N_8950,N_4866,N_4928);
or U8951 (N_8951,N_2029,N_925);
or U8952 (N_8952,N_658,N_1472);
nor U8953 (N_8953,N_2670,N_3627);
xnor U8954 (N_8954,N_741,N_2395);
or U8955 (N_8955,N_1158,N_5857);
and U8956 (N_8956,N_3638,N_1329);
nand U8957 (N_8957,N_2905,N_302);
and U8958 (N_8958,N_3496,N_1109);
nand U8959 (N_8959,N_883,N_5833);
nand U8960 (N_8960,N_4608,N_1279);
and U8961 (N_8961,N_4960,N_3484);
xor U8962 (N_8962,N_997,N_2398);
nor U8963 (N_8963,N_2259,N_789);
or U8964 (N_8964,N_966,N_1412);
or U8965 (N_8965,N_4919,N_4);
nor U8966 (N_8966,N_6111,N_2091);
nand U8967 (N_8967,N_1611,N_5944);
xnor U8968 (N_8968,N_5012,N_4709);
nand U8969 (N_8969,N_1792,N_3446);
xor U8970 (N_8970,N_6005,N_733);
or U8971 (N_8971,N_3438,N_5579);
nor U8972 (N_8972,N_3870,N_730);
xnor U8973 (N_8973,N_4293,N_2479);
or U8974 (N_8974,N_5081,N_879);
and U8975 (N_8975,N_7,N_4796);
and U8976 (N_8976,N_1987,N_5512);
nand U8977 (N_8977,N_4939,N_4933);
nor U8978 (N_8978,N_589,N_4782);
nor U8979 (N_8979,N_753,N_5395);
nor U8980 (N_8980,N_2327,N_5750);
nor U8981 (N_8981,N_6242,N_1143);
xor U8982 (N_8982,N_5359,N_5277);
nand U8983 (N_8983,N_5716,N_54);
or U8984 (N_8984,N_4066,N_3912);
nand U8985 (N_8985,N_5773,N_5741);
nand U8986 (N_8986,N_2115,N_1470);
nor U8987 (N_8987,N_4927,N_4393);
nand U8988 (N_8988,N_4578,N_5169);
xor U8989 (N_8989,N_1148,N_4418);
or U8990 (N_8990,N_1165,N_5801);
xnor U8991 (N_8991,N_1668,N_5593);
nand U8992 (N_8992,N_5044,N_5265);
nand U8993 (N_8993,N_3510,N_4642);
nand U8994 (N_8994,N_4019,N_6195);
nor U8995 (N_8995,N_1648,N_2545);
nand U8996 (N_8996,N_4574,N_1836);
nor U8997 (N_8997,N_2288,N_1992);
nor U8998 (N_8998,N_2859,N_1903);
or U8999 (N_8999,N_777,N_2125);
nor U9000 (N_9000,N_1255,N_4477);
nor U9001 (N_9001,N_1423,N_988);
nand U9002 (N_9002,N_3041,N_2868);
or U9003 (N_9003,N_1958,N_1877);
xnor U9004 (N_9004,N_1254,N_4080);
or U9005 (N_9005,N_4634,N_4162);
or U9006 (N_9006,N_38,N_6246);
xor U9007 (N_9007,N_565,N_5464);
nor U9008 (N_9008,N_6097,N_371);
xor U9009 (N_9009,N_6227,N_4046);
nand U9010 (N_9010,N_3263,N_4141);
xnor U9011 (N_9011,N_4221,N_4506);
or U9012 (N_9012,N_3790,N_448);
and U9013 (N_9013,N_2033,N_1088);
or U9014 (N_9014,N_900,N_6223);
nand U9015 (N_9015,N_3580,N_5001);
xnor U9016 (N_9016,N_4155,N_2271);
xor U9017 (N_9017,N_4491,N_1270);
nor U9018 (N_9018,N_397,N_4272);
xnor U9019 (N_9019,N_4181,N_1653);
nand U9020 (N_9020,N_1443,N_4610);
xnor U9021 (N_9021,N_5965,N_1826);
or U9022 (N_9022,N_955,N_1957);
nand U9023 (N_9023,N_5957,N_468);
and U9024 (N_9024,N_2898,N_4943);
or U9025 (N_9025,N_4560,N_3561);
nor U9026 (N_9026,N_4042,N_6011);
and U9027 (N_9027,N_5990,N_6012);
nor U9028 (N_9028,N_886,N_4345);
nand U9029 (N_9029,N_4776,N_4220);
and U9030 (N_9030,N_360,N_3491);
nor U9031 (N_9031,N_3183,N_3868);
nand U9032 (N_9032,N_1348,N_5326);
nand U9033 (N_9033,N_1274,N_5669);
xor U9034 (N_9034,N_2792,N_2385);
and U9035 (N_9035,N_3795,N_3566);
nand U9036 (N_9036,N_2414,N_3458);
and U9037 (N_9037,N_3574,N_5362);
and U9038 (N_9038,N_2083,N_588);
xor U9039 (N_9039,N_2665,N_913);
or U9040 (N_9040,N_352,N_5057);
or U9041 (N_9041,N_4011,N_2964);
xnor U9042 (N_9042,N_2615,N_4078);
nand U9043 (N_9043,N_2601,N_1816);
or U9044 (N_9044,N_4595,N_5645);
or U9045 (N_9045,N_1647,N_5691);
nor U9046 (N_9046,N_2156,N_1592);
nor U9047 (N_9047,N_3207,N_489);
or U9048 (N_9048,N_3907,N_5888);
nand U9049 (N_9049,N_1889,N_2065);
nand U9050 (N_9050,N_4593,N_1860);
and U9051 (N_9051,N_4966,N_6041);
or U9052 (N_9052,N_4891,N_4701);
and U9053 (N_9053,N_2375,N_5159);
and U9054 (N_9054,N_5273,N_2790);
nand U9055 (N_9055,N_2579,N_3327);
nor U9056 (N_9056,N_3506,N_4855);
nor U9057 (N_9057,N_874,N_3066);
or U9058 (N_9058,N_2097,N_5826);
nand U9059 (N_9059,N_4863,N_3749);
xor U9060 (N_9060,N_350,N_2561);
or U9061 (N_9061,N_3765,N_3619);
xor U9062 (N_9062,N_84,N_2229);
nor U9063 (N_9063,N_1819,N_4032);
and U9064 (N_9064,N_5148,N_4124);
nand U9065 (N_9065,N_4690,N_5663);
or U9066 (N_9066,N_2608,N_912);
and U9067 (N_9067,N_5950,N_880);
or U9068 (N_9068,N_794,N_2138);
nand U9069 (N_9069,N_5227,N_4526);
xor U9070 (N_9070,N_76,N_105);
and U9071 (N_9071,N_628,N_4814);
and U9072 (N_9072,N_2081,N_5300);
and U9073 (N_9073,N_342,N_175);
and U9074 (N_9074,N_4086,N_4153);
or U9075 (N_9075,N_5894,N_5531);
xnor U9076 (N_9076,N_952,N_3333);
nand U9077 (N_9077,N_1091,N_3673);
or U9078 (N_9078,N_1432,N_4550);
nand U9079 (N_9079,N_5829,N_2623);
xor U9080 (N_9080,N_6080,N_4025);
or U9081 (N_9081,N_2413,N_1588);
or U9082 (N_9082,N_5089,N_627);
or U9083 (N_9083,N_5482,N_5037);
and U9084 (N_9084,N_2328,N_5729);
and U9085 (N_9085,N_1603,N_3648);
nor U9086 (N_9086,N_2983,N_1700);
and U9087 (N_9087,N_500,N_2354);
and U9088 (N_9088,N_4576,N_1260);
and U9089 (N_9089,N_1927,N_496);
or U9090 (N_9090,N_1872,N_1051);
nand U9091 (N_9091,N_6098,N_6152);
nand U9092 (N_9092,N_2306,N_2342);
xor U9093 (N_9093,N_4916,N_3774);
and U9094 (N_9094,N_2701,N_591);
and U9095 (N_9095,N_5984,N_2668);
nand U9096 (N_9096,N_1191,N_2014);
nor U9097 (N_9097,N_845,N_5149);
nand U9098 (N_9098,N_3113,N_5921);
nand U9099 (N_9099,N_4206,N_1240);
and U9100 (N_9100,N_2209,N_6063);
xor U9101 (N_9101,N_4112,N_308);
nand U9102 (N_9102,N_4626,N_4253);
nor U9103 (N_9103,N_3524,N_5785);
and U9104 (N_9104,N_3777,N_4364);
and U9105 (N_9105,N_723,N_1083);
and U9106 (N_9106,N_971,N_4266);
nor U9107 (N_9107,N_6151,N_4408);
and U9108 (N_9108,N_5271,N_444);
xor U9109 (N_9109,N_6075,N_5986);
or U9110 (N_9110,N_2292,N_687);
or U9111 (N_9111,N_961,N_208);
xor U9112 (N_9112,N_2880,N_5480);
nor U9113 (N_9113,N_1785,N_2225);
and U9114 (N_9114,N_3973,N_3014);
or U9115 (N_9115,N_3570,N_1922);
xor U9116 (N_9116,N_1204,N_4280);
nor U9117 (N_9117,N_4198,N_5837);
nor U9118 (N_9118,N_2162,N_2781);
nor U9119 (N_9119,N_1167,N_6028);
nor U9120 (N_9120,N_1748,N_2006);
or U9121 (N_9121,N_2947,N_3519);
or U9122 (N_9122,N_2048,N_5626);
nand U9123 (N_9123,N_1219,N_461);
nand U9124 (N_9124,N_4813,N_4907);
or U9125 (N_9125,N_1353,N_3963);
xor U9126 (N_9126,N_343,N_4373);
nand U9127 (N_9127,N_3598,N_2884);
nor U9128 (N_9128,N_3652,N_4486);
xor U9129 (N_9129,N_1616,N_2409);
nor U9130 (N_9130,N_1312,N_1606);
or U9131 (N_9131,N_2799,N_6);
and U9132 (N_9132,N_3841,N_5564);
or U9133 (N_9133,N_5624,N_6057);
or U9134 (N_9134,N_1090,N_2122);
nor U9135 (N_9135,N_3778,N_2611);
or U9136 (N_9136,N_5809,N_1638);
xnor U9137 (N_9137,N_1779,N_499);
xor U9138 (N_9138,N_2533,N_1223);
xnor U9139 (N_9139,N_1490,N_3677);
nor U9140 (N_9140,N_4191,N_1650);
xnor U9141 (N_9141,N_580,N_145);
xor U9142 (N_9142,N_4422,N_391);
or U9143 (N_9143,N_3007,N_2814);
xor U9144 (N_9144,N_3192,N_163);
and U9145 (N_9145,N_240,N_572);
nor U9146 (N_9146,N_807,N_5503);
nor U9147 (N_9147,N_233,N_5546);
xnor U9148 (N_9148,N_1556,N_6212);
or U9149 (N_9149,N_5812,N_3396);
nand U9150 (N_9150,N_1478,N_5434);
nand U9151 (N_9151,N_4658,N_4689);
and U9152 (N_9152,N_114,N_6094);
and U9153 (N_9153,N_1706,N_3092);
xor U9154 (N_9154,N_4549,N_618);
xnor U9155 (N_9155,N_5500,N_4742);
nand U9156 (N_9156,N_4033,N_2310);
nand U9157 (N_9157,N_2003,N_5171);
or U9158 (N_9158,N_5357,N_4402);
xnor U9159 (N_9159,N_4677,N_2922);
or U9160 (N_9160,N_3250,N_3221);
nand U9161 (N_9161,N_1670,N_3216);
or U9162 (N_9162,N_5945,N_3010);
or U9163 (N_9163,N_2261,N_2196);
nor U9164 (N_9164,N_72,N_4403);
xor U9165 (N_9165,N_5354,N_1558);
nor U9166 (N_9166,N_4825,N_315);
nand U9167 (N_9167,N_1918,N_4311);
and U9168 (N_9168,N_184,N_5774);
nor U9169 (N_9169,N_5378,N_5364);
nand U9170 (N_9170,N_2461,N_3272);
nor U9171 (N_9171,N_3305,N_6156);
nand U9172 (N_9172,N_5686,N_1692);
and U9173 (N_9173,N_3312,N_2929);
xnor U9174 (N_9174,N_6058,N_5502);
or U9175 (N_9175,N_2576,N_5831);
nor U9176 (N_9176,N_4877,N_71);
nor U9177 (N_9177,N_5011,N_3916);
or U9178 (N_9178,N_5157,N_3840);
xor U9179 (N_9179,N_5732,N_3258);
or U9180 (N_9180,N_5574,N_4178);
or U9181 (N_9181,N_3690,N_4783);
nand U9182 (N_9182,N_5217,N_2369);
xor U9183 (N_9183,N_1369,N_4500);
or U9184 (N_9184,N_481,N_6067);
nand U9185 (N_9185,N_4223,N_1806);
and U9186 (N_9186,N_2421,N_5220);
xnor U9187 (N_9187,N_6015,N_2995);
and U9188 (N_9188,N_363,N_1543);
and U9189 (N_9189,N_3070,N_2434);
or U9190 (N_9190,N_4666,N_4195);
nand U9191 (N_9191,N_1210,N_3227);
nand U9192 (N_9192,N_3640,N_3115);
nand U9193 (N_9193,N_3782,N_4862);
or U9194 (N_9194,N_3294,N_4117);
and U9195 (N_9195,N_6207,N_1593);
nor U9196 (N_9196,N_1981,N_5292);
nand U9197 (N_9197,N_3489,N_3133);
or U9198 (N_9198,N_2056,N_5030);
or U9199 (N_9199,N_2345,N_4372);
and U9200 (N_9200,N_4680,N_1940);
or U9201 (N_9201,N_5247,N_3660);
nor U9202 (N_9202,N_6071,N_5946);
xnor U9203 (N_9203,N_5529,N_4092);
or U9204 (N_9204,N_135,N_4426);
nor U9205 (N_9205,N_3909,N_1629);
or U9206 (N_9206,N_4572,N_1229);
and U9207 (N_9207,N_3539,N_5017);
and U9208 (N_9208,N_5198,N_1337);
nand U9209 (N_9209,N_2296,N_3343);
or U9210 (N_9210,N_2711,N_3823);
nand U9211 (N_9211,N_3994,N_2726);
or U9212 (N_9212,N_734,N_5470);
nand U9213 (N_9213,N_2684,N_1471);
or U9214 (N_9214,N_3102,N_3467);
and U9215 (N_9215,N_4841,N_4954);
nand U9216 (N_9216,N_2452,N_4102);
and U9217 (N_9217,N_2436,N_1719);
and U9218 (N_9218,N_2554,N_5810);
xor U9219 (N_9219,N_379,N_1018);
and U9220 (N_9220,N_5477,N_129);
xnor U9221 (N_9221,N_4973,N_1781);
nor U9222 (N_9222,N_2809,N_1163);
nor U9223 (N_9223,N_6127,N_110);
nor U9224 (N_9224,N_2829,N_897);
or U9225 (N_9225,N_1932,N_2853);
nor U9226 (N_9226,N_1065,N_5435);
and U9227 (N_9227,N_3521,N_6184);
or U9228 (N_9228,N_2628,N_4516);
or U9229 (N_9229,N_2222,N_788);
and U9230 (N_9230,N_4991,N_1531);
xor U9231 (N_9231,N_292,N_3761);
nor U9232 (N_9232,N_1963,N_5709);
nor U9233 (N_9233,N_4547,N_1555);
and U9234 (N_9234,N_3875,N_3957);
or U9235 (N_9235,N_3927,N_6039);
nor U9236 (N_9236,N_3479,N_5973);
xnor U9237 (N_9237,N_4611,N_4407);
and U9238 (N_9238,N_5416,N_4476);
xnor U9239 (N_9239,N_3106,N_3940);
xnor U9240 (N_9240,N_5002,N_4317);
or U9241 (N_9241,N_5486,N_241);
or U9242 (N_9242,N_1798,N_6100);
nand U9243 (N_9243,N_139,N_86);
nor U9244 (N_9244,N_3152,N_5597);
or U9245 (N_9245,N_1747,N_3993);
or U9246 (N_9246,N_3128,N_4157);
or U9247 (N_9247,N_5046,N_2939);
nand U9248 (N_9248,N_567,N_5637);
and U9249 (N_9249,N_3240,N_4132);
and U9250 (N_9250,N_4488,N_5103);
or U9251 (N_9251,N_4753,N_5295);
and U9252 (N_9252,N_5282,N_3755);
nor U9253 (N_9253,N_3971,N_1177);
nor U9254 (N_9254,N_26,N_4655);
xor U9255 (N_9255,N_2129,N_4781);
or U9256 (N_9256,N_2954,N_5896);
nor U9257 (N_9257,N_268,N_5575);
and U9258 (N_9258,N_4996,N_1342);
or U9259 (N_9259,N_376,N_299);
or U9260 (N_9260,N_2904,N_4864);
nor U9261 (N_9261,N_2188,N_5137);
or U9262 (N_9262,N_1361,N_483);
and U9263 (N_9263,N_1316,N_4405);
nor U9264 (N_9264,N_1267,N_4606);
nor U9265 (N_9265,N_2870,N_2555);
and U9266 (N_9266,N_1711,N_4098);
nand U9267 (N_9267,N_5262,N_5870);
nand U9268 (N_9268,N_290,N_4233);
xnor U9269 (N_9269,N_2501,N_2240);
nand U9270 (N_9270,N_50,N_781);
nor U9271 (N_9271,N_6229,N_3430);
and U9272 (N_9272,N_705,N_5698);
nand U9273 (N_9273,N_2046,N_5071);
nor U9274 (N_9274,N_2735,N_2731);
nand U9275 (N_9275,N_4465,N_4425);
or U9276 (N_9276,N_4203,N_1523);
and U9277 (N_9277,N_5421,N_689);
or U9278 (N_9278,N_4142,N_1242);
nor U9279 (N_9279,N_2783,N_296);
and U9280 (N_9280,N_1098,N_151);
nand U9281 (N_9281,N_2449,N_2178);
and U9282 (N_9282,N_4065,N_4830);
and U9283 (N_9283,N_1516,N_4934);
and U9284 (N_9284,N_3031,N_252);
or U9285 (N_9285,N_6073,N_517);
nor U9286 (N_9286,N_4743,N_3468);
xor U9287 (N_9287,N_3637,N_3928);
and U9288 (N_9288,N_773,N_4283);
or U9289 (N_9289,N_1422,N_681);
xnor U9290 (N_9290,N_5848,N_4160);
nor U9291 (N_9291,N_3162,N_3485);
nor U9292 (N_9292,N_1295,N_434);
and U9293 (N_9293,N_5330,N_675);
nand U9294 (N_9294,N_364,N_1815);
nor U9295 (N_9295,N_3833,N_5697);
or U9296 (N_9296,N_2320,N_5515);
or U9297 (N_9297,N_6168,N_5091);
nand U9298 (N_9298,N_5646,N_1043);
nor U9299 (N_9299,N_3837,N_2486);
or U9300 (N_9300,N_2401,N_2938);
and U9301 (N_9301,N_3686,N_4137);
nand U9302 (N_9302,N_4026,N_847);
and U9303 (N_9303,N_2624,N_3346);
nand U9304 (N_9304,N_3730,N_2055);
nand U9305 (N_9305,N_3351,N_3179);
and U9306 (N_9306,N_2667,N_4459);
nor U9307 (N_9307,N_3407,N_3883);
nand U9308 (N_9308,N_1425,N_3756);
nand U9309 (N_9309,N_1156,N_1702);
nand U9310 (N_9310,N_5734,N_4913);
nor U9311 (N_9311,N_259,N_5701);
nand U9312 (N_9312,N_5849,N_2252);
and U9313 (N_9313,N_4773,N_4757);
xnor U9314 (N_9314,N_1654,N_6017);
nand U9315 (N_9315,N_5397,N_1870);
and U9316 (N_9316,N_5659,N_29);
or U9317 (N_9317,N_4852,N_5170);
and U9318 (N_9318,N_1460,N_4455);
xor U9319 (N_9319,N_3397,N_6145);
xor U9320 (N_9320,N_4148,N_6196);
nand U9321 (N_9321,N_5086,N_4245);
nor U9322 (N_9322,N_1475,N_4811);
nor U9323 (N_9323,N_1031,N_3442);
nand U9324 (N_9324,N_3545,N_6204);
nand U9325 (N_9325,N_4327,N_2709);
and U9326 (N_9326,N_3887,N_1505);
and U9327 (N_9327,N_3454,N_6066);
or U9328 (N_9328,N_1421,N_4394);
or U9329 (N_9329,N_4800,N_5769);
xnor U9330 (N_9330,N_2931,N_3990);
nor U9331 (N_9331,N_6221,N_877);
and U9332 (N_9332,N_5313,N_2467);
and U9333 (N_9333,N_5804,N_5852);
xor U9334 (N_9334,N_4136,N_3136);
nor U9335 (N_9335,N_1597,N_526);
xor U9336 (N_9336,N_2316,N_2584);
and U9337 (N_9337,N_2071,N_5083);
or U9338 (N_9338,N_5634,N_4997);
or U9339 (N_9339,N_2339,N_515);
nor U9340 (N_9340,N_2673,N_4975);
and U9341 (N_9341,N_2626,N_4558);
or U9342 (N_9342,N_2403,N_2897);
and U9343 (N_9343,N_1568,N_2036);
xor U9344 (N_9344,N_418,N_2552);
nand U9345 (N_9345,N_1111,N_3763);
and U9346 (N_9346,N_4775,N_2695);
nor U9347 (N_9347,N_4986,N_2174);
nand U9348 (N_9348,N_2738,N_1200);
nand U9349 (N_9349,N_4482,N_2638);
and U9350 (N_9350,N_1173,N_4821);
or U9351 (N_9351,N_5980,N_2689);
or U9352 (N_9352,N_856,N_2009);
and U9353 (N_9353,N_647,N_673);
or U9354 (N_9354,N_5552,N_4561);
nor U9355 (N_9355,N_1496,N_3060);
nor U9356 (N_9356,N_917,N_5889);
and U9357 (N_9357,N_5093,N_5074);
and U9358 (N_9358,N_2765,N_1170);
nor U9359 (N_9359,N_5760,N_5795);
nor U9360 (N_9360,N_3720,N_1694);
or U9361 (N_9361,N_484,N_2143);
xor U9362 (N_9362,N_1169,N_3836);
and U9363 (N_9363,N_2458,N_122);
or U9364 (N_9364,N_2537,N_806);
nor U9365 (N_9365,N_5431,N_3494);
and U9366 (N_9366,N_236,N_4985);
nand U9367 (N_9367,N_4375,N_1905);
nand U9368 (N_9368,N_2757,N_4467);
nor U9369 (N_9369,N_1794,N_4532);
nor U9370 (N_9370,N_3243,N_5518);
nor U9371 (N_9371,N_4432,N_1800);
nor U9372 (N_9372,N_4750,N_251);
and U9373 (N_9373,N_2186,N_347);
and U9374 (N_9374,N_5213,N_2179);
xnor U9375 (N_9375,N_5151,N_3844);
nor U9376 (N_9376,N_867,N_5223);
nand U9377 (N_9377,N_1657,N_1032);
or U9378 (N_9378,N_4097,N_6235);
nor U9379 (N_9379,N_1485,N_5498);
and U9380 (N_9380,N_1716,N_1764);
xor U9381 (N_9381,N_5590,N_6007);
or U9382 (N_9382,N_5138,N_951);
or U9383 (N_9383,N_2553,N_5636);
and U9384 (N_9384,N_5632,N_4226);
xnor U9385 (N_9385,N_2314,N_4712);
or U9386 (N_9386,N_1513,N_3799);
or U9387 (N_9387,N_2220,N_4485);
nor U9388 (N_9388,N_5400,N_358);
xnor U9389 (N_9389,N_1225,N_865);
nor U9390 (N_9390,N_1221,N_4904);
nor U9391 (N_9391,N_2182,N_2459);
nand U9392 (N_9392,N_4683,N_4774);
nand U9393 (N_9393,N_2112,N_1857);
nor U9394 (N_9394,N_1921,N_5062);
and U9395 (N_9395,N_4039,N_1158);
nand U9396 (N_9396,N_4866,N_4370);
or U9397 (N_9397,N_1407,N_4238);
xnor U9398 (N_9398,N_967,N_3758);
nand U9399 (N_9399,N_5738,N_1216);
or U9400 (N_9400,N_1990,N_339);
nand U9401 (N_9401,N_5454,N_2619);
xor U9402 (N_9402,N_4407,N_4603);
and U9403 (N_9403,N_3286,N_5966);
nand U9404 (N_9404,N_5830,N_2342);
or U9405 (N_9405,N_2294,N_4234);
or U9406 (N_9406,N_573,N_5614);
and U9407 (N_9407,N_2071,N_3129);
nand U9408 (N_9408,N_2513,N_5625);
nor U9409 (N_9409,N_3450,N_57);
nor U9410 (N_9410,N_5030,N_3606);
and U9411 (N_9411,N_75,N_5510);
or U9412 (N_9412,N_2642,N_2798);
xor U9413 (N_9413,N_5811,N_2671);
xor U9414 (N_9414,N_2370,N_634);
nor U9415 (N_9415,N_2781,N_3473);
xor U9416 (N_9416,N_2372,N_5569);
nand U9417 (N_9417,N_1170,N_4690);
xnor U9418 (N_9418,N_2820,N_5118);
xor U9419 (N_9419,N_1829,N_1003);
or U9420 (N_9420,N_4462,N_4483);
and U9421 (N_9421,N_2450,N_5731);
nor U9422 (N_9422,N_5218,N_3544);
nor U9423 (N_9423,N_2095,N_3493);
nand U9424 (N_9424,N_2574,N_5945);
nor U9425 (N_9425,N_5323,N_4247);
or U9426 (N_9426,N_3942,N_2949);
xor U9427 (N_9427,N_1688,N_3158);
nor U9428 (N_9428,N_2824,N_1387);
and U9429 (N_9429,N_1798,N_3910);
or U9430 (N_9430,N_4004,N_6233);
and U9431 (N_9431,N_1499,N_1203);
or U9432 (N_9432,N_1207,N_2464);
and U9433 (N_9433,N_1820,N_4353);
or U9434 (N_9434,N_2570,N_1852);
nand U9435 (N_9435,N_4153,N_2866);
or U9436 (N_9436,N_261,N_4667);
and U9437 (N_9437,N_539,N_133);
and U9438 (N_9438,N_4276,N_5682);
xnor U9439 (N_9439,N_779,N_429);
or U9440 (N_9440,N_2408,N_1551);
nand U9441 (N_9441,N_1696,N_4302);
and U9442 (N_9442,N_1921,N_1096);
nand U9443 (N_9443,N_5153,N_2684);
or U9444 (N_9444,N_3496,N_1694);
or U9445 (N_9445,N_4565,N_524);
nand U9446 (N_9446,N_5735,N_3524);
nand U9447 (N_9447,N_3749,N_1061);
xor U9448 (N_9448,N_4223,N_4877);
xnor U9449 (N_9449,N_4434,N_3743);
and U9450 (N_9450,N_4691,N_120);
nand U9451 (N_9451,N_1784,N_905);
xor U9452 (N_9452,N_2323,N_406);
and U9453 (N_9453,N_5923,N_141);
nor U9454 (N_9454,N_3742,N_2413);
xor U9455 (N_9455,N_2961,N_1829);
or U9456 (N_9456,N_401,N_80);
xnor U9457 (N_9457,N_435,N_425);
or U9458 (N_9458,N_1569,N_5976);
nor U9459 (N_9459,N_5301,N_6050);
xnor U9460 (N_9460,N_4346,N_2418);
xnor U9461 (N_9461,N_3695,N_2426);
nand U9462 (N_9462,N_4088,N_5903);
nor U9463 (N_9463,N_4471,N_1978);
xnor U9464 (N_9464,N_2116,N_1887);
xor U9465 (N_9465,N_5939,N_4392);
or U9466 (N_9466,N_5365,N_3223);
or U9467 (N_9467,N_1771,N_2118);
nand U9468 (N_9468,N_612,N_2259);
nand U9469 (N_9469,N_4062,N_2994);
nand U9470 (N_9470,N_3125,N_606);
and U9471 (N_9471,N_5155,N_5124);
or U9472 (N_9472,N_998,N_3441);
and U9473 (N_9473,N_6037,N_3669);
nand U9474 (N_9474,N_1043,N_2363);
or U9475 (N_9475,N_6076,N_1367);
nor U9476 (N_9476,N_1974,N_3245);
nand U9477 (N_9477,N_4527,N_3299);
or U9478 (N_9478,N_1699,N_5977);
and U9479 (N_9479,N_1237,N_564);
nor U9480 (N_9480,N_5107,N_2490);
nor U9481 (N_9481,N_4841,N_4966);
xnor U9482 (N_9482,N_5803,N_5962);
or U9483 (N_9483,N_2123,N_5687);
xnor U9484 (N_9484,N_2220,N_3095);
nand U9485 (N_9485,N_4099,N_1652);
nand U9486 (N_9486,N_4275,N_1585);
xnor U9487 (N_9487,N_1602,N_456);
and U9488 (N_9488,N_5630,N_5404);
and U9489 (N_9489,N_2709,N_4630);
nor U9490 (N_9490,N_4721,N_4413);
or U9491 (N_9491,N_4154,N_5261);
or U9492 (N_9492,N_2277,N_2324);
nor U9493 (N_9493,N_3014,N_3375);
or U9494 (N_9494,N_1912,N_4288);
xor U9495 (N_9495,N_1130,N_1474);
and U9496 (N_9496,N_673,N_181);
xor U9497 (N_9497,N_63,N_4950);
and U9498 (N_9498,N_4419,N_1642);
nor U9499 (N_9499,N_2679,N_100);
nor U9500 (N_9500,N_3245,N_3643);
nor U9501 (N_9501,N_6007,N_4789);
nand U9502 (N_9502,N_3112,N_5000);
or U9503 (N_9503,N_2275,N_4750);
and U9504 (N_9504,N_4661,N_4003);
or U9505 (N_9505,N_3714,N_1424);
and U9506 (N_9506,N_401,N_892);
and U9507 (N_9507,N_1225,N_318);
xnor U9508 (N_9508,N_434,N_2752);
and U9509 (N_9509,N_1842,N_6019);
and U9510 (N_9510,N_2909,N_256);
xor U9511 (N_9511,N_4171,N_4264);
and U9512 (N_9512,N_3378,N_3476);
or U9513 (N_9513,N_6141,N_5878);
nand U9514 (N_9514,N_1892,N_6029);
nand U9515 (N_9515,N_1222,N_5280);
or U9516 (N_9516,N_1004,N_2837);
or U9517 (N_9517,N_3142,N_1817);
and U9518 (N_9518,N_2461,N_5773);
nor U9519 (N_9519,N_6099,N_5947);
nor U9520 (N_9520,N_3929,N_1004);
nor U9521 (N_9521,N_2340,N_3480);
nand U9522 (N_9522,N_5391,N_2763);
nand U9523 (N_9523,N_2514,N_2714);
nor U9524 (N_9524,N_5570,N_2023);
nor U9525 (N_9525,N_3031,N_3958);
and U9526 (N_9526,N_2954,N_966);
nand U9527 (N_9527,N_4154,N_152);
nor U9528 (N_9528,N_3963,N_2157);
nand U9529 (N_9529,N_309,N_869);
xor U9530 (N_9530,N_3304,N_4575);
xor U9531 (N_9531,N_1865,N_5732);
or U9532 (N_9532,N_5728,N_3971);
nor U9533 (N_9533,N_4513,N_2112);
nand U9534 (N_9534,N_984,N_2511);
or U9535 (N_9535,N_2328,N_2295);
nand U9536 (N_9536,N_2988,N_5696);
and U9537 (N_9537,N_3445,N_4335);
xnor U9538 (N_9538,N_3065,N_5104);
or U9539 (N_9539,N_6094,N_4425);
nand U9540 (N_9540,N_1856,N_720);
xnor U9541 (N_9541,N_1423,N_488);
or U9542 (N_9542,N_5052,N_914);
and U9543 (N_9543,N_3787,N_4495);
nor U9544 (N_9544,N_831,N_1976);
nor U9545 (N_9545,N_547,N_982);
xnor U9546 (N_9546,N_4209,N_250);
nand U9547 (N_9547,N_2720,N_1697);
or U9548 (N_9548,N_2029,N_4074);
nor U9549 (N_9549,N_4574,N_337);
xnor U9550 (N_9550,N_4727,N_232);
nand U9551 (N_9551,N_5373,N_385);
and U9552 (N_9552,N_6137,N_552);
xor U9553 (N_9553,N_3747,N_3375);
xor U9554 (N_9554,N_3361,N_1632);
xnor U9555 (N_9555,N_4066,N_6195);
or U9556 (N_9556,N_5230,N_4787);
or U9557 (N_9557,N_1245,N_4225);
nand U9558 (N_9558,N_3128,N_1834);
and U9559 (N_9559,N_3847,N_4713);
and U9560 (N_9560,N_5375,N_1909);
nor U9561 (N_9561,N_4477,N_822);
and U9562 (N_9562,N_5982,N_1356);
nor U9563 (N_9563,N_290,N_5427);
nand U9564 (N_9564,N_3564,N_1676);
nor U9565 (N_9565,N_395,N_4321);
nor U9566 (N_9566,N_1041,N_5488);
and U9567 (N_9567,N_1666,N_1325);
or U9568 (N_9568,N_2135,N_2407);
or U9569 (N_9569,N_3065,N_2755);
or U9570 (N_9570,N_5237,N_357);
xnor U9571 (N_9571,N_5146,N_1534);
xnor U9572 (N_9572,N_1430,N_2313);
xor U9573 (N_9573,N_4852,N_5914);
nand U9574 (N_9574,N_2259,N_1623);
nor U9575 (N_9575,N_5396,N_1934);
xor U9576 (N_9576,N_2683,N_4113);
nand U9577 (N_9577,N_4559,N_6144);
xnor U9578 (N_9578,N_6180,N_5489);
and U9579 (N_9579,N_2882,N_5504);
or U9580 (N_9580,N_3550,N_6038);
xor U9581 (N_9581,N_2688,N_5776);
nor U9582 (N_9582,N_1565,N_5581);
or U9583 (N_9583,N_1493,N_4679);
nor U9584 (N_9584,N_5200,N_122);
and U9585 (N_9585,N_5755,N_2832);
nor U9586 (N_9586,N_3673,N_2425);
and U9587 (N_9587,N_2759,N_418);
nor U9588 (N_9588,N_4037,N_1663);
nor U9589 (N_9589,N_3591,N_3343);
xnor U9590 (N_9590,N_3142,N_1482);
or U9591 (N_9591,N_216,N_5733);
xor U9592 (N_9592,N_6018,N_5309);
nor U9593 (N_9593,N_1549,N_6117);
nand U9594 (N_9594,N_4385,N_4906);
xor U9595 (N_9595,N_4762,N_3670);
nand U9596 (N_9596,N_4353,N_2100);
nand U9597 (N_9597,N_3325,N_2801);
and U9598 (N_9598,N_5580,N_27);
and U9599 (N_9599,N_5211,N_1256);
nand U9600 (N_9600,N_5294,N_5435);
or U9601 (N_9601,N_433,N_4460);
nor U9602 (N_9602,N_6056,N_2038);
and U9603 (N_9603,N_1197,N_1958);
nand U9604 (N_9604,N_4502,N_3301);
nand U9605 (N_9605,N_4904,N_781);
or U9606 (N_9606,N_1489,N_5659);
or U9607 (N_9607,N_3177,N_3525);
xor U9608 (N_9608,N_671,N_3375);
and U9609 (N_9609,N_2469,N_3748);
or U9610 (N_9610,N_2887,N_2265);
xnor U9611 (N_9611,N_1141,N_4282);
and U9612 (N_9612,N_1239,N_3653);
xor U9613 (N_9613,N_1548,N_38);
and U9614 (N_9614,N_954,N_2651);
and U9615 (N_9615,N_2878,N_3487);
and U9616 (N_9616,N_1954,N_2145);
and U9617 (N_9617,N_2548,N_1380);
nor U9618 (N_9618,N_4711,N_1062);
xor U9619 (N_9619,N_3784,N_1637);
and U9620 (N_9620,N_947,N_4154);
nand U9621 (N_9621,N_5304,N_4645);
xor U9622 (N_9622,N_3810,N_2784);
nand U9623 (N_9623,N_870,N_3546);
or U9624 (N_9624,N_4032,N_1444);
xor U9625 (N_9625,N_583,N_2306);
xor U9626 (N_9626,N_165,N_1011);
nor U9627 (N_9627,N_928,N_3060);
nor U9628 (N_9628,N_4899,N_3782);
or U9629 (N_9629,N_3784,N_2938);
or U9630 (N_9630,N_4463,N_581);
xor U9631 (N_9631,N_964,N_4782);
nor U9632 (N_9632,N_784,N_5397);
or U9633 (N_9633,N_1596,N_4464);
xor U9634 (N_9634,N_2363,N_2648);
xor U9635 (N_9635,N_3632,N_2608);
xnor U9636 (N_9636,N_3150,N_5190);
xor U9637 (N_9637,N_2915,N_3189);
nand U9638 (N_9638,N_139,N_6232);
or U9639 (N_9639,N_4566,N_5236);
nand U9640 (N_9640,N_1605,N_106);
nor U9641 (N_9641,N_1461,N_2511);
nand U9642 (N_9642,N_3476,N_3978);
nor U9643 (N_9643,N_3405,N_3600);
and U9644 (N_9644,N_5211,N_135);
nand U9645 (N_9645,N_2766,N_1421);
and U9646 (N_9646,N_5046,N_3003);
nand U9647 (N_9647,N_4320,N_2965);
nor U9648 (N_9648,N_1360,N_448);
nand U9649 (N_9649,N_880,N_5143);
nand U9650 (N_9650,N_2371,N_4478);
xnor U9651 (N_9651,N_1054,N_1327);
nor U9652 (N_9652,N_3182,N_5694);
nor U9653 (N_9653,N_5009,N_1620);
xnor U9654 (N_9654,N_3883,N_3855);
nand U9655 (N_9655,N_5465,N_5585);
and U9656 (N_9656,N_3301,N_2976);
xnor U9657 (N_9657,N_2457,N_686);
nand U9658 (N_9658,N_1702,N_3025);
xor U9659 (N_9659,N_4998,N_1362);
nand U9660 (N_9660,N_2786,N_2359);
nand U9661 (N_9661,N_1985,N_5140);
nor U9662 (N_9662,N_5303,N_5133);
nand U9663 (N_9663,N_5175,N_299);
nand U9664 (N_9664,N_6142,N_2405);
and U9665 (N_9665,N_5000,N_4313);
or U9666 (N_9666,N_770,N_3406);
and U9667 (N_9667,N_2091,N_5980);
and U9668 (N_9668,N_3274,N_3763);
and U9669 (N_9669,N_5362,N_1520);
nor U9670 (N_9670,N_1578,N_2558);
xor U9671 (N_9671,N_5452,N_1905);
xnor U9672 (N_9672,N_2775,N_947);
or U9673 (N_9673,N_6140,N_6150);
or U9674 (N_9674,N_4320,N_1706);
xor U9675 (N_9675,N_2159,N_236);
xnor U9676 (N_9676,N_2806,N_2119);
nor U9677 (N_9677,N_2798,N_453);
or U9678 (N_9678,N_3492,N_5790);
or U9679 (N_9679,N_2633,N_5746);
or U9680 (N_9680,N_6124,N_4952);
xor U9681 (N_9681,N_1104,N_418);
xnor U9682 (N_9682,N_2748,N_2211);
nand U9683 (N_9683,N_5198,N_5515);
xnor U9684 (N_9684,N_1282,N_5309);
nand U9685 (N_9685,N_2346,N_3813);
and U9686 (N_9686,N_2268,N_5557);
or U9687 (N_9687,N_3851,N_4293);
nand U9688 (N_9688,N_4445,N_6156);
nand U9689 (N_9689,N_1795,N_2454);
or U9690 (N_9690,N_2161,N_2139);
xnor U9691 (N_9691,N_2810,N_3748);
nand U9692 (N_9692,N_5227,N_2912);
or U9693 (N_9693,N_2832,N_3344);
nor U9694 (N_9694,N_41,N_2218);
or U9695 (N_9695,N_4499,N_4603);
nor U9696 (N_9696,N_3291,N_3120);
and U9697 (N_9697,N_1954,N_32);
xor U9698 (N_9698,N_3090,N_1848);
xnor U9699 (N_9699,N_6135,N_1281);
nor U9700 (N_9700,N_977,N_1017);
and U9701 (N_9701,N_4701,N_5683);
or U9702 (N_9702,N_2449,N_4992);
nor U9703 (N_9703,N_2077,N_6081);
nor U9704 (N_9704,N_1785,N_937);
nor U9705 (N_9705,N_3071,N_5887);
or U9706 (N_9706,N_728,N_1359);
and U9707 (N_9707,N_5442,N_828);
nor U9708 (N_9708,N_2114,N_5732);
nand U9709 (N_9709,N_3219,N_1450);
or U9710 (N_9710,N_2780,N_5820);
or U9711 (N_9711,N_34,N_5066);
and U9712 (N_9712,N_5397,N_5399);
xor U9713 (N_9713,N_1199,N_1714);
and U9714 (N_9714,N_2510,N_4665);
nand U9715 (N_9715,N_3528,N_196);
nand U9716 (N_9716,N_1561,N_1919);
nand U9717 (N_9717,N_2014,N_2431);
or U9718 (N_9718,N_2269,N_5057);
xnor U9719 (N_9719,N_2393,N_1119);
nor U9720 (N_9720,N_3262,N_2826);
xor U9721 (N_9721,N_2481,N_6190);
nor U9722 (N_9722,N_101,N_2684);
nand U9723 (N_9723,N_2424,N_2970);
xor U9724 (N_9724,N_3226,N_2380);
and U9725 (N_9725,N_4422,N_3179);
nand U9726 (N_9726,N_422,N_4373);
nor U9727 (N_9727,N_5549,N_1980);
xnor U9728 (N_9728,N_5460,N_582);
xor U9729 (N_9729,N_1884,N_4631);
xor U9730 (N_9730,N_4077,N_878);
or U9731 (N_9731,N_6046,N_3662);
nor U9732 (N_9732,N_446,N_3620);
nand U9733 (N_9733,N_205,N_5263);
and U9734 (N_9734,N_4101,N_5463);
and U9735 (N_9735,N_523,N_3323);
xnor U9736 (N_9736,N_5122,N_4315);
or U9737 (N_9737,N_4676,N_4953);
nand U9738 (N_9738,N_4861,N_215);
nor U9739 (N_9739,N_2297,N_191);
nor U9740 (N_9740,N_4598,N_2491);
or U9741 (N_9741,N_933,N_4205);
nor U9742 (N_9742,N_3918,N_4715);
xnor U9743 (N_9743,N_6195,N_2318);
nand U9744 (N_9744,N_348,N_1314);
nand U9745 (N_9745,N_2120,N_5830);
nand U9746 (N_9746,N_2133,N_5356);
or U9747 (N_9747,N_5584,N_2779);
nor U9748 (N_9748,N_1238,N_979);
and U9749 (N_9749,N_996,N_1967);
or U9750 (N_9750,N_492,N_1494);
xnor U9751 (N_9751,N_5558,N_6015);
and U9752 (N_9752,N_975,N_1825);
and U9753 (N_9753,N_74,N_4243);
or U9754 (N_9754,N_513,N_1985);
xnor U9755 (N_9755,N_1268,N_1935);
xnor U9756 (N_9756,N_4735,N_4944);
or U9757 (N_9757,N_1047,N_4229);
xor U9758 (N_9758,N_1372,N_6175);
nor U9759 (N_9759,N_4288,N_4326);
and U9760 (N_9760,N_3760,N_3844);
and U9761 (N_9761,N_4688,N_5156);
and U9762 (N_9762,N_4924,N_4550);
nand U9763 (N_9763,N_2180,N_400);
or U9764 (N_9764,N_3829,N_1500);
or U9765 (N_9765,N_1013,N_4624);
xor U9766 (N_9766,N_4150,N_1120);
and U9767 (N_9767,N_6187,N_5899);
and U9768 (N_9768,N_1276,N_2089);
xor U9769 (N_9769,N_1031,N_5123);
nand U9770 (N_9770,N_4471,N_531);
xor U9771 (N_9771,N_2686,N_3172);
nand U9772 (N_9772,N_5167,N_4259);
xor U9773 (N_9773,N_5363,N_3913);
and U9774 (N_9774,N_4762,N_251);
nand U9775 (N_9775,N_206,N_984);
or U9776 (N_9776,N_156,N_2847);
nor U9777 (N_9777,N_4201,N_3801);
or U9778 (N_9778,N_5072,N_3611);
or U9779 (N_9779,N_2585,N_894);
xnor U9780 (N_9780,N_3385,N_909);
nand U9781 (N_9781,N_2057,N_5093);
or U9782 (N_9782,N_5934,N_942);
and U9783 (N_9783,N_810,N_4908);
and U9784 (N_9784,N_5611,N_117);
or U9785 (N_9785,N_1423,N_5753);
and U9786 (N_9786,N_173,N_4052);
nand U9787 (N_9787,N_5735,N_1139);
and U9788 (N_9788,N_5618,N_2456);
nor U9789 (N_9789,N_4187,N_6186);
xor U9790 (N_9790,N_5533,N_3919);
nand U9791 (N_9791,N_4940,N_4374);
nor U9792 (N_9792,N_2915,N_4219);
nor U9793 (N_9793,N_2372,N_5442);
or U9794 (N_9794,N_5868,N_4109);
nand U9795 (N_9795,N_6243,N_3315);
and U9796 (N_9796,N_4275,N_4969);
or U9797 (N_9797,N_4903,N_703);
xor U9798 (N_9798,N_1693,N_5850);
xnor U9799 (N_9799,N_4909,N_5503);
nor U9800 (N_9800,N_4527,N_4779);
and U9801 (N_9801,N_5835,N_4421);
nand U9802 (N_9802,N_4955,N_1685);
xor U9803 (N_9803,N_2583,N_1311);
nor U9804 (N_9804,N_3135,N_3649);
or U9805 (N_9805,N_1798,N_3759);
or U9806 (N_9806,N_2483,N_5482);
or U9807 (N_9807,N_6073,N_58);
and U9808 (N_9808,N_3057,N_945);
and U9809 (N_9809,N_3385,N_5076);
and U9810 (N_9810,N_4429,N_1059);
xor U9811 (N_9811,N_1180,N_5049);
nor U9812 (N_9812,N_5434,N_2212);
nand U9813 (N_9813,N_1093,N_1981);
nand U9814 (N_9814,N_204,N_75);
and U9815 (N_9815,N_4221,N_3064);
or U9816 (N_9816,N_4871,N_3326);
nor U9817 (N_9817,N_3430,N_1537);
or U9818 (N_9818,N_3342,N_2946);
nand U9819 (N_9819,N_4121,N_2162);
or U9820 (N_9820,N_2829,N_6140);
nand U9821 (N_9821,N_4236,N_1606);
and U9822 (N_9822,N_286,N_2468);
nand U9823 (N_9823,N_3278,N_4540);
nor U9824 (N_9824,N_207,N_5354);
and U9825 (N_9825,N_5182,N_353);
nor U9826 (N_9826,N_2820,N_3673);
xor U9827 (N_9827,N_2010,N_4845);
xor U9828 (N_9828,N_3532,N_5514);
nand U9829 (N_9829,N_14,N_5399);
xor U9830 (N_9830,N_1999,N_133);
or U9831 (N_9831,N_897,N_2849);
xor U9832 (N_9832,N_3329,N_1015);
nor U9833 (N_9833,N_4574,N_4787);
nor U9834 (N_9834,N_2876,N_1315);
or U9835 (N_9835,N_4386,N_2994);
and U9836 (N_9836,N_903,N_2015);
xnor U9837 (N_9837,N_2824,N_5036);
or U9838 (N_9838,N_3069,N_5135);
or U9839 (N_9839,N_1803,N_3357);
or U9840 (N_9840,N_6209,N_2952);
nor U9841 (N_9841,N_1877,N_1189);
nand U9842 (N_9842,N_953,N_1239);
and U9843 (N_9843,N_3197,N_6082);
xor U9844 (N_9844,N_4376,N_3735);
nor U9845 (N_9845,N_1739,N_3757);
nand U9846 (N_9846,N_4194,N_2428);
nor U9847 (N_9847,N_533,N_2835);
nand U9848 (N_9848,N_959,N_3685);
xnor U9849 (N_9849,N_5792,N_3675);
xnor U9850 (N_9850,N_1187,N_891);
and U9851 (N_9851,N_1475,N_3592);
or U9852 (N_9852,N_2724,N_5398);
nand U9853 (N_9853,N_4818,N_3093);
nand U9854 (N_9854,N_1223,N_681);
or U9855 (N_9855,N_4843,N_4378);
xnor U9856 (N_9856,N_5699,N_2942);
nand U9857 (N_9857,N_1098,N_2522);
and U9858 (N_9858,N_4693,N_2873);
nor U9859 (N_9859,N_5916,N_1442);
xnor U9860 (N_9860,N_5115,N_3093);
xnor U9861 (N_9861,N_2606,N_3539);
nor U9862 (N_9862,N_5960,N_3299);
nor U9863 (N_9863,N_4111,N_4707);
nand U9864 (N_9864,N_3623,N_1525);
nand U9865 (N_9865,N_1046,N_1660);
nor U9866 (N_9866,N_205,N_923);
nor U9867 (N_9867,N_5549,N_4300);
and U9868 (N_9868,N_4187,N_1885);
xor U9869 (N_9869,N_4554,N_2013);
nand U9870 (N_9870,N_3772,N_3206);
nor U9871 (N_9871,N_4564,N_5570);
or U9872 (N_9872,N_4931,N_3093);
nor U9873 (N_9873,N_2444,N_2711);
nor U9874 (N_9874,N_2508,N_3801);
or U9875 (N_9875,N_5457,N_3750);
nor U9876 (N_9876,N_4672,N_311);
nor U9877 (N_9877,N_4363,N_3750);
nand U9878 (N_9878,N_5891,N_608);
xor U9879 (N_9879,N_4656,N_1338);
or U9880 (N_9880,N_938,N_1851);
nor U9881 (N_9881,N_4600,N_701);
and U9882 (N_9882,N_3597,N_2051);
xor U9883 (N_9883,N_2353,N_3157);
xnor U9884 (N_9884,N_1427,N_642);
nor U9885 (N_9885,N_6059,N_2924);
and U9886 (N_9886,N_5773,N_553);
nor U9887 (N_9887,N_1990,N_3955);
and U9888 (N_9888,N_1377,N_321);
nor U9889 (N_9889,N_3145,N_5867);
xnor U9890 (N_9890,N_3110,N_4845);
nor U9891 (N_9891,N_3065,N_1759);
nand U9892 (N_9892,N_81,N_5824);
and U9893 (N_9893,N_3711,N_2895);
nor U9894 (N_9894,N_3749,N_5260);
or U9895 (N_9895,N_1284,N_5169);
xnor U9896 (N_9896,N_2067,N_1098);
xor U9897 (N_9897,N_3580,N_75);
xnor U9898 (N_9898,N_5700,N_46);
nor U9899 (N_9899,N_6033,N_5296);
and U9900 (N_9900,N_4533,N_2483);
nand U9901 (N_9901,N_1005,N_5067);
nand U9902 (N_9902,N_4033,N_693);
nor U9903 (N_9903,N_1624,N_1829);
and U9904 (N_9904,N_2813,N_1851);
xor U9905 (N_9905,N_3350,N_1176);
nand U9906 (N_9906,N_3590,N_1233);
nor U9907 (N_9907,N_4144,N_3979);
nand U9908 (N_9908,N_4850,N_4502);
nand U9909 (N_9909,N_5317,N_1561);
nor U9910 (N_9910,N_2161,N_2746);
and U9911 (N_9911,N_2559,N_4186);
nand U9912 (N_9912,N_2665,N_3940);
nor U9913 (N_9913,N_4341,N_4905);
nor U9914 (N_9914,N_5860,N_2753);
nand U9915 (N_9915,N_5595,N_3572);
nor U9916 (N_9916,N_2941,N_6060);
nor U9917 (N_9917,N_2063,N_2428);
or U9918 (N_9918,N_505,N_1177);
nor U9919 (N_9919,N_3351,N_5104);
nand U9920 (N_9920,N_2963,N_1790);
nand U9921 (N_9921,N_2586,N_4052);
nor U9922 (N_9922,N_5432,N_5312);
nor U9923 (N_9923,N_2459,N_171);
nor U9924 (N_9924,N_639,N_1612);
and U9925 (N_9925,N_1106,N_4104);
nor U9926 (N_9926,N_3285,N_4841);
xor U9927 (N_9927,N_2880,N_370);
or U9928 (N_9928,N_3307,N_228);
or U9929 (N_9929,N_2731,N_4649);
or U9930 (N_9930,N_5468,N_1898);
nor U9931 (N_9931,N_3680,N_1910);
nor U9932 (N_9932,N_1897,N_3488);
and U9933 (N_9933,N_1475,N_2150);
nor U9934 (N_9934,N_5231,N_5979);
nor U9935 (N_9935,N_4810,N_4996);
nand U9936 (N_9936,N_4534,N_3835);
xor U9937 (N_9937,N_3402,N_3116);
nor U9938 (N_9938,N_4256,N_1341);
or U9939 (N_9939,N_195,N_3788);
nor U9940 (N_9940,N_3909,N_5466);
xor U9941 (N_9941,N_3131,N_165);
nor U9942 (N_9942,N_3075,N_3889);
xnor U9943 (N_9943,N_6038,N_6214);
xnor U9944 (N_9944,N_2182,N_734);
nor U9945 (N_9945,N_120,N_3455);
nand U9946 (N_9946,N_1431,N_4186);
or U9947 (N_9947,N_4719,N_1170);
nand U9948 (N_9948,N_2010,N_610);
nand U9949 (N_9949,N_5784,N_1675);
nand U9950 (N_9950,N_4858,N_5486);
nor U9951 (N_9951,N_1988,N_4583);
nor U9952 (N_9952,N_330,N_2334);
and U9953 (N_9953,N_3235,N_1927);
nor U9954 (N_9954,N_5588,N_508);
nor U9955 (N_9955,N_927,N_2137);
and U9956 (N_9956,N_4871,N_3838);
xnor U9957 (N_9957,N_3540,N_1730);
or U9958 (N_9958,N_4095,N_2609);
and U9959 (N_9959,N_2699,N_4391);
or U9960 (N_9960,N_3504,N_2650);
and U9961 (N_9961,N_2915,N_1505);
xor U9962 (N_9962,N_5259,N_4405);
and U9963 (N_9963,N_1567,N_2743);
and U9964 (N_9964,N_2346,N_1872);
nor U9965 (N_9965,N_5548,N_1005);
and U9966 (N_9966,N_5445,N_5199);
nand U9967 (N_9967,N_2873,N_4917);
xor U9968 (N_9968,N_3916,N_248);
or U9969 (N_9969,N_1904,N_5643);
nand U9970 (N_9970,N_4280,N_1579);
and U9971 (N_9971,N_2957,N_1484);
or U9972 (N_9972,N_1607,N_1287);
xor U9973 (N_9973,N_5419,N_2575);
and U9974 (N_9974,N_1639,N_3773);
or U9975 (N_9975,N_5153,N_4705);
and U9976 (N_9976,N_2458,N_4824);
xnor U9977 (N_9977,N_2036,N_328);
or U9978 (N_9978,N_2069,N_1353);
xnor U9979 (N_9979,N_1249,N_2739);
xnor U9980 (N_9980,N_3361,N_5648);
or U9981 (N_9981,N_1237,N_5556);
and U9982 (N_9982,N_2474,N_4816);
and U9983 (N_9983,N_533,N_6090);
and U9984 (N_9984,N_5711,N_2410);
xnor U9985 (N_9985,N_1944,N_3003);
nand U9986 (N_9986,N_4897,N_758);
and U9987 (N_9987,N_4761,N_2610);
or U9988 (N_9988,N_994,N_5109);
and U9989 (N_9989,N_458,N_411);
nand U9990 (N_9990,N_4709,N_3099);
xor U9991 (N_9991,N_2614,N_4822);
nor U9992 (N_9992,N_3736,N_572);
xor U9993 (N_9993,N_1788,N_1308);
nand U9994 (N_9994,N_5542,N_1696);
or U9995 (N_9995,N_4163,N_4745);
xnor U9996 (N_9996,N_657,N_945);
and U9997 (N_9997,N_3597,N_2424);
nor U9998 (N_9998,N_2133,N_2560);
xnor U9999 (N_9999,N_1422,N_3122);
nor U10000 (N_10000,N_5382,N_3140);
nand U10001 (N_10001,N_27,N_4920);
and U10002 (N_10002,N_5980,N_5520);
xnor U10003 (N_10003,N_2729,N_5759);
nand U10004 (N_10004,N_1263,N_3580);
nor U10005 (N_10005,N_5875,N_2691);
and U10006 (N_10006,N_1485,N_4610);
or U10007 (N_10007,N_3161,N_1599);
and U10008 (N_10008,N_4138,N_5553);
or U10009 (N_10009,N_4987,N_1058);
nor U10010 (N_10010,N_4669,N_4502);
xor U10011 (N_10011,N_2084,N_2740);
xnor U10012 (N_10012,N_4950,N_1398);
nand U10013 (N_10013,N_5254,N_2421);
or U10014 (N_10014,N_1301,N_616);
or U10015 (N_10015,N_2501,N_5602);
or U10016 (N_10016,N_2530,N_181);
nor U10017 (N_10017,N_594,N_5683);
nor U10018 (N_10018,N_3658,N_1020);
and U10019 (N_10019,N_1494,N_6248);
or U10020 (N_10020,N_431,N_405);
or U10021 (N_10021,N_4005,N_3317);
and U10022 (N_10022,N_1512,N_4031);
nand U10023 (N_10023,N_4352,N_6071);
and U10024 (N_10024,N_833,N_795);
nor U10025 (N_10025,N_3376,N_1249);
nand U10026 (N_10026,N_1813,N_5489);
xnor U10027 (N_10027,N_1631,N_3354);
and U10028 (N_10028,N_1316,N_1858);
and U10029 (N_10029,N_4259,N_5893);
xnor U10030 (N_10030,N_1578,N_5344);
nand U10031 (N_10031,N_1092,N_2533);
xnor U10032 (N_10032,N_4862,N_3595);
nand U10033 (N_10033,N_5715,N_2588);
and U10034 (N_10034,N_1819,N_2102);
nand U10035 (N_10035,N_1575,N_5607);
xor U10036 (N_10036,N_5842,N_5856);
nor U10037 (N_10037,N_2638,N_1005);
nand U10038 (N_10038,N_3427,N_4200);
nor U10039 (N_10039,N_3642,N_790);
xnor U10040 (N_10040,N_2336,N_765);
nand U10041 (N_10041,N_1703,N_1688);
nand U10042 (N_10042,N_6109,N_2431);
nor U10043 (N_10043,N_2768,N_5533);
nor U10044 (N_10044,N_1779,N_1933);
or U10045 (N_10045,N_1385,N_3523);
xor U10046 (N_10046,N_1200,N_2325);
nor U10047 (N_10047,N_4697,N_1709);
or U10048 (N_10048,N_1005,N_93);
xor U10049 (N_10049,N_1354,N_1522);
or U10050 (N_10050,N_5100,N_49);
nor U10051 (N_10051,N_6054,N_4830);
xnor U10052 (N_10052,N_3156,N_4913);
nand U10053 (N_10053,N_96,N_2439);
and U10054 (N_10054,N_1459,N_1257);
xnor U10055 (N_10055,N_4447,N_250);
nand U10056 (N_10056,N_4045,N_3886);
and U10057 (N_10057,N_4722,N_202);
xnor U10058 (N_10058,N_2768,N_2835);
or U10059 (N_10059,N_3998,N_741);
or U10060 (N_10060,N_2084,N_5904);
nand U10061 (N_10061,N_6156,N_5529);
or U10062 (N_10062,N_5268,N_1260);
nor U10063 (N_10063,N_4396,N_6088);
or U10064 (N_10064,N_4159,N_1696);
xor U10065 (N_10065,N_521,N_4855);
and U10066 (N_10066,N_2451,N_5664);
nor U10067 (N_10067,N_2020,N_1143);
and U10068 (N_10068,N_3454,N_5453);
xnor U10069 (N_10069,N_1332,N_4003);
and U10070 (N_10070,N_505,N_2748);
or U10071 (N_10071,N_4322,N_5558);
and U10072 (N_10072,N_2385,N_3535);
nor U10073 (N_10073,N_1402,N_5541);
and U10074 (N_10074,N_5104,N_4333);
xnor U10075 (N_10075,N_2053,N_1756);
nand U10076 (N_10076,N_4625,N_1310);
or U10077 (N_10077,N_5978,N_777);
xnor U10078 (N_10078,N_3304,N_5020);
and U10079 (N_10079,N_1286,N_2733);
nand U10080 (N_10080,N_4860,N_796);
and U10081 (N_10081,N_348,N_3575);
and U10082 (N_10082,N_2062,N_3355);
nor U10083 (N_10083,N_2066,N_4571);
nor U10084 (N_10084,N_6016,N_1656);
or U10085 (N_10085,N_3326,N_3538);
and U10086 (N_10086,N_2446,N_1133);
xor U10087 (N_10087,N_960,N_2768);
and U10088 (N_10088,N_6003,N_1550);
nand U10089 (N_10089,N_2236,N_2268);
nor U10090 (N_10090,N_5023,N_2539);
xnor U10091 (N_10091,N_3833,N_3927);
or U10092 (N_10092,N_1286,N_2858);
nor U10093 (N_10093,N_1668,N_1181);
or U10094 (N_10094,N_4552,N_3626);
or U10095 (N_10095,N_4072,N_3462);
nand U10096 (N_10096,N_935,N_366);
nor U10097 (N_10097,N_2352,N_1734);
xor U10098 (N_10098,N_4749,N_4964);
nand U10099 (N_10099,N_126,N_145);
nor U10100 (N_10100,N_79,N_163);
xor U10101 (N_10101,N_5663,N_893);
or U10102 (N_10102,N_3772,N_891);
xnor U10103 (N_10103,N_4558,N_1425);
xnor U10104 (N_10104,N_4673,N_4763);
nor U10105 (N_10105,N_4028,N_3162);
xor U10106 (N_10106,N_5499,N_5468);
and U10107 (N_10107,N_1053,N_5125);
nand U10108 (N_10108,N_2492,N_5183);
nor U10109 (N_10109,N_2709,N_4001);
nand U10110 (N_10110,N_922,N_5218);
nand U10111 (N_10111,N_2585,N_2794);
or U10112 (N_10112,N_2870,N_219);
or U10113 (N_10113,N_1187,N_1830);
xnor U10114 (N_10114,N_782,N_5836);
or U10115 (N_10115,N_5004,N_4660);
xnor U10116 (N_10116,N_4392,N_100);
and U10117 (N_10117,N_1141,N_5662);
or U10118 (N_10118,N_5051,N_5592);
xnor U10119 (N_10119,N_2934,N_2418);
or U10120 (N_10120,N_420,N_2405);
or U10121 (N_10121,N_2878,N_887);
and U10122 (N_10122,N_2920,N_4235);
nand U10123 (N_10123,N_1106,N_5991);
or U10124 (N_10124,N_1207,N_444);
nand U10125 (N_10125,N_3445,N_5331);
nand U10126 (N_10126,N_706,N_4352);
nor U10127 (N_10127,N_1469,N_1856);
and U10128 (N_10128,N_5673,N_210);
xnor U10129 (N_10129,N_2574,N_1285);
and U10130 (N_10130,N_4795,N_3056);
xor U10131 (N_10131,N_2159,N_1313);
nand U10132 (N_10132,N_5861,N_4615);
or U10133 (N_10133,N_5397,N_4008);
nor U10134 (N_10134,N_537,N_51);
nor U10135 (N_10135,N_4515,N_1570);
and U10136 (N_10136,N_4803,N_3531);
or U10137 (N_10137,N_1614,N_5099);
nor U10138 (N_10138,N_2622,N_1522);
xor U10139 (N_10139,N_5858,N_5044);
and U10140 (N_10140,N_3890,N_1513);
or U10141 (N_10141,N_3113,N_6105);
and U10142 (N_10142,N_1539,N_4593);
nand U10143 (N_10143,N_1338,N_258);
and U10144 (N_10144,N_6117,N_5362);
and U10145 (N_10145,N_5612,N_6007);
nor U10146 (N_10146,N_963,N_2891);
nor U10147 (N_10147,N_1873,N_1353);
xor U10148 (N_10148,N_372,N_6202);
nand U10149 (N_10149,N_3866,N_3590);
nor U10150 (N_10150,N_1245,N_558);
and U10151 (N_10151,N_635,N_4140);
and U10152 (N_10152,N_5469,N_5282);
nand U10153 (N_10153,N_5382,N_1822);
xor U10154 (N_10154,N_5847,N_6072);
nor U10155 (N_10155,N_1404,N_3862);
and U10156 (N_10156,N_1687,N_1799);
nand U10157 (N_10157,N_4474,N_1155);
nand U10158 (N_10158,N_311,N_1106);
and U10159 (N_10159,N_5652,N_3282);
nand U10160 (N_10160,N_251,N_3042);
xor U10161 (N_10161,N_5201,N_2530);
or U10162 (N_10162,N_4670,N_2018);
and U10163 (N_10163,N_1193,N_5774);
nor U10164 (N_10164,N_894,N_2386);
nor U10165 (N_10165,N_386,N_5904);
nor U10166 (N_10166,N_4951,N_6008);
or U10167 (N_10167,N_4596,N_3838);
or U10168 (N_10168,N_5627,N_4310);
nand U10169 (N_10169,N_1292,N_5408);
nand U10170 (N_10170,N_4125,N_2471);
nand U10171 (N_10171,N_2847,N_2550);
and U10172 (N_10172,N_3492,N_4981);
or U10173 (N_10173,N_1752,N_4481);
and U10174 (N_10174,N_3554,N_868);
nor U10175 (N_10175,N_5517,N_1315);
xor U10176 (N_10176,N_447,N_2659);
or U10177 (N_10177,N_384,N_2216);
nand U10178 (N_10178,N_753,N_1325);
nand U10179 (N_10179,N_5148,N_3573);
xor U10180 (N_10180,N_1142,N_2501);
or U10181 (N_10181,N_4631,N_6177);
nor U10182 (N_10182,N_682,N_4945);
nand U10183 (N_10183,N_5475,N_3116);
nand U10184 (N_10184,N_1815,N_1953);
or U10185 (N_10185,N_3517,N_1058);
or U10186 (N_10186,N_1572,N_4891);
nand U10187 (N_10187,N_4651,N_3506);
xnor U10188 (N_10188,N_3919,N_5469);
and U10189 (N_10189,N_4798,N_4091);
nor U10190 (N_10190,N_1215,N_422);
nor U10191 (N_10191,N_2653,N_5006);
xnor U10192 (N_10192,N_5568,N_5928);
nor U10193 (N_10193,N_1752,N_3213);
xor U10194 (N_10194,N_184,N_2977);
or U10195 (N_10195,N_346,N_4053);
and U10196 (N_10196,N_667,N_717);
xnor U10197 (N_10197,N_1719,N_4654);
or U10198 (N_10198,N_4808,N_5641);
xnor U10199 (N_10199,N_1054,N_3835);
or U10200 (N_10200,N_2275,N_3259);
nor U10201 (N_10201,N_6189,N_4684);
xor U10202 (N_10202,N_3125,N_83);
nand U10203 (N_10203,N_1738,N_4669);
xor U10204 (N_10204,N_1283,N_5414);
and U10205 (N_10205,N_5894,N_314);
or U10206 (N_10206,N_2874,N_2344);
and U10207 (N_10207,N_2226,N_3871);
nor U10208 (N_10208,N_2628,N_1287);
or U10209 (N_10209,N_984,N_3609);
or U10210 (N_10210,N_613,N_55);
nand U10211 (N_10211,N_5546,N_1541);
or U10212 (N_10212,N_6124,N_2773);
xnor U10213 (N_10213,N_363,N_4934);
and U10214 (N_10214,N_2928,N_2262);
nor U10215 (N_10215,N_328,N_6210);
xnor U10216 (N_10216,N_1402,N_1414);
and U10217 (N_10217,N_2130,N_3990);
and U10218 (N_10218,N_4912,N_3932);
and U10219 (N_10219,N_3591,N_2435);
xnor U10220 (N_10220,N_5749,N_4523);
nand U10221 (N_10221,N_4309,N_5873);
nand U10222 (N_10222,N_5576,N_1429);
xor U10223 (N_10223,N_2725,N_3228);
xnor U10224 (N_10224,N_1513,N_137);
xor U10225 (N_10225,N_1961,N_559);
and U10226 (N_10226,N_1926,N_1050);
nand U10227 (N_10227,N_1315,N_154);
or U10228 (N_10228,N_5169,N_5143);
or U10229 (N_10229,N_3979,N_5082);
nand U10230 (N_10230,N_4697,N_2776);
nand U10231 (N_10231,N_5746,N_1818);
xor U10232 (N_10232,N_2572,N_4106);
and U10233 (N_10233,N_6105,N_3394);
and U10234 (N_10234,N_4072,N_4890);
nand U10235 (N_10235,N_2464,N_5003);
or U10236 (N_10236,N_3109,N_5245);
or U10237 (N_10237,N_3139,N_3021);
nor U10238 (N_10238,N_1920,N_5711);
or U10239 (N_10239,N_1263,N_5075);
xnor U10240 (N_10240,N_546,N_4431);
xnor U10241 (N_10241,N_4041,N_3300);
nand U10242 (N_10242,N_3126,N_1227);
nand U10243 (N_10243,N_2503,N_4650);
nand U10244 (N_10244,N_2895,N_5775);
and U10245 (N_10245,N_3012,N_4938);
or U10246 (N_10246,N_4880,N_2269);
nand U10247 (N_10247,N_1501,N_5165);
or U10248 (N_10248,N_4575,N_3601);
nor U10249 (N_10249,N_3914,N_6042);
and U10250 (N_10250,N_2040,N_5892);
xor U10251 (N_10251,N_1010,N_3038);
or U10252 (N_10252,N_1393,N_480);
or U10253 (N_10253,N_1314,N_3342);
and U10254 (N_10254,N_4827,N_495);
nand U10255 (N_10255,N_5362,N_4102);
nand U10256 (N_10256,N_4433,N_1961);
and U10257 (N_10257,N_4068,N_1425);
or U10258 (N_10258,N_4319,N_3462);
nor U10259 (N_10259,N_3962,N_4575);
and U10260 (N_10260,N_2951,N_3526);
or U10261 (N_10261,N_5761,N_4729);
xor U10262 (N_10262,N_2087,N_1014);
nand U10263 (N_10263,N_4396,N_3656);
nand U10264 (N_10264,N_1814,N_4977);
xor U10265 (N_10265,N_2699,N_303);
nor U10266 (N_10266,N_6121,N_1201);
and U10267 (N_10267,N_2705,N_5331);
nand U10268 (N_10268,N_3132,N_4824);
xnor U10269 (N_10269,N_2287,N_4931);
xor U10270 (N_10270,N_2661,N_3339);
nand U10271 (N_10271,N_176,N_4902);
and U10272 (N_10272,N_5260,N_5110);
nand U10273 (N_10273,N_1660,N_184);
or U10274 (N_10274,N_4034,N_4552);
nand U10275 (N_10275,N_103,N_1736);
or U10276 (N_10276,N_5237,N_4288);
or U10277 (N_10277,N_341,N_1292);
nor U10278 (N_10278,N_5479,N_213);
xor U10279 (N_10279,N_2170,N_3191);
or U10280 (N_10280,N_3470,N_124);
xor U10281 (N_10281,N_4273,N_573);
and U10282 (N_10282,N_4184,N_577);
and U10283 (N_10283,N_5443,N_1036);
or U10284 (N_10284,N_4071,N_1615);
nor U10285 (N_10285,N_2908,N_1310);
nand U10286 (N_10286,N_1072,N_4620);
or U10287 (N_10287,N_3832,N_652);
nor U10288 (N_10288,N_6139,N_2726);
xnor U10289 (N_10289,N_3896,N_6014);
nor U10290 (N_10290,N_3564,N_162);
nor U10291 (N_10291,N_6115,N_1466);
and U10292 (N_10292,N_5285,N_342);
xor U10293 (N_10293,N_424,N_2851);
xor U10294 (N_10294,N_3154,N_4477);
nand U10295 (N_10295,N_3505,N_6073);
nor U10296 (N_10296,N_3370,N_2897);
nor U10297 (N_10297,N_3344,N_3756);
nand U10298 (N_10298,N_3429,N_3889);
nor U10299 (N_10299,N_5909,N_1591);
xor U10300 (N_10300,N_2014,N_6038);
nor U10301 (N_10301,N_4709,N_4379);
or U10302 (N_10302,N_1189,N_1530);
nand U10303 (N_10303,N_4249,N_2053);
nor U10304 (N_10304,N_3795,N_3022);
or U10305 (N_10305,N_3892,N_4652);
xor U10306 (N_10306,N_2362,N_6189);
and U10307 (N_10307,N_145,N_225);
and U10308 (N_10308,N_3903,N_4817);
nand U10309 (N_10309,N_2249,N_1199);
and U10310 (N_10310,N_1300,N_2915);
nor U10311 (N_10311,N_1962,N_3486);
nand U10312 (N_10312,N_2395,N_5993);
and U10313 (N_10313,N_3028,N_3954);
or U10314 (N_10314,N_442,N_2653);
and U10315 (N_10315,N_4037,N_5471);
or U10316 (N_10316,N_3038,N_5370);
nand U10317 (N_10317,N_4785,N_3312);
nand U10318 (N_10318,N_3263,N_3695);
and U10319 (N_10319,N_1295,N_2269);
xor U10320 (N_10320,N_1795,N_5697);
nand U10321 (N_10321,N_2603,N_2260);
and U10322 (N_10322,N_4613,N_93);
or U10323 (N_10323,N_2730,N_5902);
or U10324 (N_10324,N_1658,N_3955);
xnor U10325 (N_10325,N_1845,N_5130);
xor U10326 (N_10326,N_596,N_1336);
nor U10327 (N_10327,N_2722,N_1746);
xor U10328 (N_10328,N_921,N_2679);
or U10329 (N_10329,N_3206,N_1223);
xor U10330 (N_10330,N_5648,N_3823);
and U10331 (N_10331,N_4628,N_3004);
nor U10332 (N_10332,N_6162,N_5645);
nand U10333 (N_10333,N_5672,N_5351);
xor U10334 (N_10334,N_2355,N_4458);
nor U10335 (N_10335,N_934,N_451);
xor U10336 (N_10336,N_5056,N_2277);
nor U10337 (N_10337,N_6206,N_4552);
xor U10338 (N_10338,N_1991,N_5611);
nor U10339 (N_10339,N_717,N_4383);
or U10340 (N_10340,N_3645,N_3917);
nand U10341 (N_10341,N_5691,N_3209);
xnor U10342 (N_10342,N_2577,N_6070);
nand U10343 (N_10343,N_2129,N_2245);
nand U10344 (N_10344,N_2517,N_689);
or U10345 (N_10345,N_3739,N_2534);
nand U10346 (N_10346,N_5646,N_1670);
xor U10347 (N_10347,N_937,N_1753);
nand U10348 (N_10348,N_5084,N_3585);
nor U10349 (N_10349,N_1823,N_3275);
xnor U10350 (N_10350,N_725,N_2253);
xor U10351 (N_10351,N_1291,N_4663);
and U10352 (N_10352,N_2270,N_3752);
xor U10353 (N_10353,N_3775,N_2340);
xnor U10354 (N_10354,N_5447,N_1133);
or U10355 (N_10355,N_5202,N_6237);
xor U10356 (N_10356,N_5754,N_2581);
or U10357 (N_10357,N_3326,N_2400);
xor U10358 (N_10358,N_5184,N_6056);
xor U10359 (N_10359,N_3404,N_569);
or U10360 (N_10360,N_4629,N_5469);
nor U10361 (N_10361,N_2882,N_2809);
nand U10362 (N_10362,N_794,N_5430);
nor U10363 (N_10363,N_4060,N_3513);
nand U10364 (N_10364,N_4830,N_4559);
xor U10365 (N_10365,N_572,N_893);
and U10366 (N_10366,N_1698,N_2632);
and U10367 (N_10367,N_1000,N_5833);
or U10368 (N_10368,N_3362,N_4895);
nor U10369 (N_10369,N_3065,N_4807);
or U10370 (N_10370,N_4198,N_8);
or U10371 (N_10371,N_1200,N_1426);
xnor U10372 (N_10372,N_3806,N_3661);
or U10373 (N_10373,N_3843,N_1764);
nand U10374 (N_10374,N_3343,N_2668);
nand U10375 (N_10375,N_3305,N_2);
nor U10376 (N_10376,N_983,N_1687);
xnor U10377 (N_10377,N_5084,N_5357);
and U10378 (N_10378,N_2482,N_3825);
nor U10379 (N_10379,N_2475,N_6184);
xor U10380 (N_10380,N_838,N_5939);
or U10381 (N_10381,N_1137,N_3847);
nand U10382 (N_10382,N_3750,N_3578);
and U10383 (N_10383,N_5829,N_2712);
xnor U10384 (N_10384,N_5359,N_1712);
nand U10385 (N_10385,N_319,N_4220);
or U10386 (N_10386,N_4176,N_1566);
nand U10387 (N_10387,N_832,N_5798);
nand U10388 (N_10388,N_3942,N_5149);
and U10389 (N_10389,N_4045,N_1627);
xor U10390 (N_10390,N_4735,N_4744);
and U10391 (N_10391,N_2326,N_3282);
nor U10392 (N_10392,N_5788,N_3396);
or U10393 (N_10393,N_5799,N_259);
xor U10394 (N_10394,N_4986,N_3384);
nand U10395 (N_10395,N_1896,N_1934);
nand U10396 (N_10396,N_4831,N_4939);
or U10397 (N_10397,N_4293,N_1336);
nor U10398 (N_10398,N_2409,N_2518);
and U10399 (N_10399,N_1753,N_6093);
and U10400 (N_10400,N_3085,N_1771);
nand U10401 (N_10401,N_5763,N_931);
or U10402 (N_10402,N_5218,N_4174);
xnor U10403 (N_10403,N_2300,N_2209);
and U10404 (N_10404,N_3921,N_4283);
or U10405 (N_10405,N_1040,N_1855);
and U10406 (N_10406,N_3822,N_1671);
nand U10407 (N_10407,N_2021,N_3590);
xor U10408 (N_10408,N_80,N_2722);
nor U10409 (N_10409,N_2206,N_3482);
nand U10410 (N_10410,N_4752,N_1364);
nand U10411 (N_10411,N_2239,N_5869);
xnor U10412 (N_10412,N_4670,N_5077);
nor U10413 (N_10413,N_2272,N_701);
nand U10414 (N_10414,N_4340,N_5073);
nand U10415 (N_10415,N_2828,N_4106);
xor U10416 (N_10416,N_5044,N_6151);
and U10417 (N_10417,N_5792,N_1035);
or U10418 (N_10418,N_4502,N_3534);
or U10419 (N_10419,N_1072,N_2292);
or U10420 (N_10420,N_6143,N_1996);
or U10421 (N_10421,N_263,N_5678);
nor U10422 (N_10422,N_3061,N_4422);
xnor U10423 (N_10423,N_11,N_5708);
or U10424 (N_10424,N_6059,N_5717);
or U10425 (N_10425,N_2375,N_1215);
nand U10426 (N_10426,N_2997,N_1701);
or U10427 (N_10427,N_4373,N_2966);
or U10428 (N_10428,N_5398,N_1704);
nand U10429 (N_10429,N_950,N_949);
nand U10430 (N_10430,N_4690,N_1120);
xnor U10431 (N_10431,N_5219,N_1025);
or U10432 (N_10432,N_4167,N_4631);
xnor U10433 (N_10433,N_3261,N_2482);
or U10434 (N_10434,N_4415,N_3471);
nand U10435 (N_10435,N_1871,N_2425);
and U10436 (N_10436,N_4949,N_4718);
or U10437 (N_10437,N_2924,N_3485);
xnor U10438 (N_10438,N_3333,N_4635);
nand U10439 (N_10439,N_288,N_3117);
or U10440 (N_10440,N_6141,N_5164);
xnor U10441 (N_10441,N_3536,N_4063);
nor U10442 (N_10442,N_1012,N_2719);
or U10443 (N_10443,N_778,N_3970);
or U10444 (N_10444,N_6124,N_4174);
and U10445 (N_10445,N_4449,N_3796);
nor U10446 (N_10446,N_3100,N_2535);
or U10447 (N_10447,N_3035,N_1046);
nor U10448 (N_10448,N_6192,N_1085);
xor U10449 (N_10449,N_250,N_5277);
or U10450 (N_10450,N_637,N_65);
xnor U10451 (N_10451,N_4128,N_2468);
nor U10452 (N_10452,N_1531,N_3751);
xnor U10453 (N_10453,N_2104,N_1054);
or U10454 (N_10454,N_2214,N_2280);
xnor U10455 (N_10455,N_1502,N_204);
and U10456 (N_10456,N_1905,N_5828);
nor U10457 (N_10457,N_545,N_3538);
nand U10458 (N_10458,N_1505,N_1723);
and U10459 (N_10459,N_3118,N_5606);
xnor U10460 (N_10460,N_5787,N_6099);
or U10461 (N_10461,N_2132,N_2380);
nand U10462 (N_10462,N_3081,N_4748);
nor U10463 (N_10463,N_30,N_414);
and U10464 (N_10464,N_4384,N_183);
or U10465 (N_10465,N_5304,N_4751);
and U10466 (N_10466,N_4115,N_1394);
or U10467 (N_10467,N_3068,N_2418);
and U10468 (N_10468,N_5033,N_2534);
and U10469 (N_10469,N_2623,N_3496);
nand U10470 (N_10470,N_2082,N_3397);
xor U10471 (N_10471,N_3616,N_108);
nand U10472 (N_10472,N_2942,N_4202);
and U10473 (N_10473,N_5185,N_1365);
nor U10474 (N_10474,N_3426,N_1710);
xor U10475 (N_10475,N_1424,N_4821);
nand U10476 (N_10476,N_4351,N_1332);
xor U10477 (N_10477,N_3118,N_3664);
xor U10478 (N_10478,N_3417,N_3693);
or U10479 (N_10479,N_4136,N_4985);
nor U10480 (N_10480,N_3388,N_5015);
or U10481 (N_10481,N_4785,N_1311);
and U10482 (N_10482,N_2527,N_4037);
nand U10483 (N_10483,N_5968,N_377);
xor U10484 (N_10484,N_5242,N_4394);
or U10485 (N_10485,N_6176,N_1717);
nand U10486 (N_10486,N_5918,N_545);
nand U10487 (N_10487,N_5918,N_3241);
nor U10488 (N_10488,N_4347,N_6018);
or U10489 (N_10489,N_5953,N_4793);
and U10490 (N_10490,N_2384,N_2156);
xnor U10491 (N_10491,N_5111,N_5547);
and U10492 (N_10492,N_3665,N_5153);
or U10493 (N_10493,N_1476,N_5744);
or U10494 (N_10494,N_4555,N_2901);
xor U10495 (N_10495,N_2395,N_710);
and U10496 (N_10496,N_616,N_2807);
or U10497 (N_10497,N_2895,N_724);
or U10498 (N_10498,N_4364,N_5392);
xnor U10499 (N_10499,N_4479,N_4111);
nand U10500 (N_10500,N_663,N_29);
nor U10501 (N_10501,N_2796,N_4133);
xor U10502 (N_10502,N_273,N_3516);
nor U10503 (N_10503,N_5392,N_1040);
nand U10504 (N_10504,N_4825,N_1662);
nor U10505 (N_10505,N_3461,N_5143);
and U10506 (N_10506,N_2875,N_4993);
and U10507 (N_10507,N_2796,N_4239);
nor U10508 (N_10508,N_4308,N_987);
xnor U10509 (N_10509,N_5883,N_1749);
nand U10510 (N_10510,N_3929,N_4338);
and U10511 (N_10511,N_4357,N_2634);
xnor U10512 (N_10512,N_4244,N_265);
xor U10513 (N_10513,N_2307,N_1686);
nor U10514 (N_10514,N_4293,N_4266);
or U10515 (N_10515,N_1166,N_4095);
or U10516 (N_10516,N_2536,N_4396);
xnor U10517 (N_10517,N_5478,N_793);
nor U10518 (N_10518,N_5907,N_4663);
and U10519 (N_10519,N_1916,N_3149);
and U10520 (N_10520,N_6021,N_2070);
xnor U10521 (N_10521,N_3317,N_4998);
nor U10522 (N_10522,N_819,N_5655);
or U10523 (N_10523,N_5668,N_1046);
nand U10524 (N_10524,N_4913,N_4700);
nor U10525 (N_10525,N_5118,N_437);
or U10526 (N_10526,N_476,N_2018);
xnor U10527 (N_10527,N_3839,N_451);
or U10528 (N_10528,N_1485,N_1317);
and U10529 (N_10529,N_1309,N_5572);
nand U10530 (N_10530,N_1483,N_2915);
nor U10531 (N_10531,N_2491,N_2011);
and U10532 (N_10532,N_3133,N_4904);
nand U10533 (N_10533,N_2946,N_2717);
nor U10534 (N_10534,N_5335,N_1009);
xnor U10535 (N_10535,N_1904,N_1703);
nand U10536 (N_10536,N_5819,N_5184);
and U10537 (N_10537,N_3557,N_616);
or U10538 (N_10538,N_3023,N_5403);
nand U10539 (N_10539,N_882,N_5417);
or U10540 (N_10540,N_2926,N_1585);
nand U10541 (N_10541,N_1013,N_5001);
and U10542 (N_10542,N_5996,N_4114);
nor U10543 (N_10543,N_6243,N_5173);
or U10544 (N_10544,N_2888,N_3661);
or U10545 (N_10545,N_386,N_3673);
xor U10546 (N_10546,N_5545,N_1073);
and U10547 (N_10547,N_1482,N_2278);
xnor U10548 (N_10548,N_1249,N_2354);
nor U10549 (N_10549,N_2051,N_5090);
nor U10550 (N_10550,N_1114,N_3477);
nor U10551 (N_10551,N_2388,N_3560);
nor U10552 (N_10552,N_5866,N_6175);
nand U10553 (N_10553,N_4232,N_1197);
xor U10554 (N_10554,N_5586,N_1921);
nor U10555 (N_10555,N_3450,N_1401);
and U10556 (N_10556,N_5888,N_1295);
nand U10557 (N_10557,N_5788,N_1763);
and U10558 (N_10558,N_2377,N_4688);
or U10559 (N_10559,N_739,N_4642);
xnor U10560 (N_10560,N_229,N_2380);
xnor U10561 (N_10561,N_2782,N_5273);
nand U10562 (N_10562,N_2134,N_3487);
or U10563 (N_10563,N_5073,N_1770);
xor U10564 (N_10564,N_811,N_5880);
and U10565 (N_10565,N_505,N_4525);
nand U10566 (N_10566,N_6143,N_2234);
xor U10567 (N_10567,N_3692,N_151);
or U10568 (N_10568,N_6180,N_1993);
and U10569 (N_10569,N_1291,N_5985);
nand U10570 (N_10570,N_3692,N_4031);
or U10571 (N_10571,N_3748,N_3826);
and U10572 (N_10572,N_5689,N_1202);
or U10573 (N_10573,N_4241,N_3720);
and U10574 (N_10574,N_5090,N_2220);
nand U10575 (N_10575,N_2231,N_128);
xor U10576 (N_10576,N_1339,N_1116);
nor U10577 (N_10577,N_327,N_4391);
nor U10578 (N_10578,N_4723,N_3744);
or U10579 (N_10579,N_4833,N_2088);
xor U10580 (N_10580,N_1479,N_1121);
and U10581 (N_10581,N_5870,N_6096);
and U10582 (N_10582,N_253,N_5742);
and U10583 (N_10583,N_356,N_3105);
nor U10584 (N_10584,N_883,N_2999);
or U10585 (N_10585,N_4394,N_4404);
nor U10586 (N_10586,N_3699,N_1391);
xnor U10587 (N_10587,N_2123,N_4653);
or U10588 (N_10588,N_5740,N_3859);
or U10589 (N_10589,N_62,N_855);
xor U10590 (N_10590,N_5826,N_2606);
or U10591 (N_10591,N_672,N_3731);
nor U10592 (N_10592,N_2641,N_2451);
nor U10593 (N_10593,N_5552,N_5077);
nor U10594 (N_10594,N_1752,N_3404);
nand U10595 (N_10595,N_2562,N_2421);
or U10596 (N_10596,N_2114,N_3196);
nand U10597 (N_10597,N_3230,N_5542);
nand U10598 (N_10598,N_1534,N_5706);
xnor U10599 (N_10599,N_2182,N_1298);
nand U10600 (N_10600,N_4046,N_5029);
nand U10601 (N_10601,N_3372,N_5472);
and U10602 (N_10602,N_4214,N_169);
and U10603 (N_10603,N_4733,N_3377);
nor U10604 (N_10604,N_858,N_5789);
xnor U10605 (N_10605,N_4928,N_2410);
nor U10606 (N_10606,N_1064,N_543);
nor U10607 (N_10607,N_3642,N_3427);
nand U10608 (N_10608,N_3026,N_789);
nor U10609 (N_10609,N_2917,N_875);
and U10610 (N_10610,N_6217,N_3749);
xor U10611 (N_10611,N_5417,N_2727);
xnor U10612 (N_10612,N_5920,N_1871);
nand U10613 (N_10613,N_2934,N_4877);
xor U10614 (N_10614,N_1113,N_6135);
nand U10615 (N_10615,N_5554,N_4875);
nor U10616 (N_10616,N_4626,N_1780);
xnor U10617 (N_10617,N_4388,N_343);
nor U10618 (N_10618,N_165,N_6180);
nand U10619 (N_10619,N_3125,N_5225);
nand U10620 (N_10620,N_5752,N_6027);
nor U10621 (N_10621,N_1355,N_3407);
or U10622 (N_10622,N_3969,N_2070);
xnor U10623 (N_10623,N_5906,N_4362);
xor U10624 (N_10624,N_2544,N_4029);
nand U10625 (N_10625,N_3331,N_56);
nand U10626 (N_10626,N_5045,N_5902);
or U10627 (N_10627,N_2731,N_1374);
or U10628 (N_10628,N_4334,N_1074);
or U10629 (N_10629,N_3873,N_86);
nor U10630 (N_10630,N_5135,N_6186);
xor U10631 (N_10631,N_1091,N_5638);
and U10632 (N_10632,N_5618,N_4033);
nand U10633 (N_10633,N_1025,N_2913);
and U10634 (N_10634,N_2280,N_1862);
xnor U10635 (N_10635,N_820,N_3504);
or U10636 (N_10636,N_5955,N_2264);
nand U10637 (N_10637,N_4314,N_3541);
nand U10638 (N_10638,N_3458,N_1899);
nor U10639 (N_10639,N_1857,N_4221);
xnor U10640 (N_10640,N_4000,N_284);
xor U10641 (N_10641,N_5987,N_459);
nand U10642 (N_10642,N_5042,N_3719);
or U10643 (N_10643,N_2556,N_3457);
nand U10644 (N_10644,N_871,N_6014);
nor U10645 (N_10645,N_6179,N_1091);
and U10646 (N_10646,N_3367,N_1910);
and U10647 (N_10647,N_4109,N_4760);
nand U10648 (N_10648,N_1815,N_1180);
nand U10649 (N_10649,N_2307,N_4725);
or U10650 (N_10650,N_781,N_2424);
nor U10651 (N_10651,N_2914,N_2333);
nor U10652 (N_10652,N_5725,N_4864);
nand U10653 (N_10653,N_4033,N_4040);
nand U10654 (N_10654,N_5792,N_1138);
xor U10655 (N_10655,N_3730,N_672);
xor U10656 (N_10656,N_4429,N_3686);
nand U10657 (N_10657,N_4673,N_5571);
nand U10658 (N_10658,N_91,N_3881);
nor U10659 (N_10659,N_4689,N_4365);
nand U10660 (N_10660,N_784,N_616);
or U10661 (N_10661,N_4877,N_89);
nor U10662 (N_10662,N_2492,N_1753);
nand U10663 (N_10663,N_435,N_2416);
xor U10664 (N_10664,N_2095,N_3281);
and U10665 (N_10665,N_2008,N_6239);
nand U10666 (N_10666,N_5418,N_2562);
and U10667 (N_10667,N_2401,N_2012);
or U10668 (N_10668,N_2557,N_6046);
xnor U10669 (N_10669,N_1065,N_6114);
nor U10670 (N_10670,N_1022,N_2834);
and U10671 (N_10671,N_3512,N_2491);
nand U10672 (N_10672,N_4373,N_1135);
nand U10673 (N_10673,N_3773,N_824);
nand U10674 (N_10674,N_2929,N_4320);
xnor U10675 (N_10675,N_2240,N_5662);
or U10676 (N_10676,N_3802,N_4522);
or U10677 (N_10677,N_2475,N_1170);
nor U10678 (N_10678,N_208,N_3385);
or U10679 (N_10679,N_1861,N_4674);
or U10680 (N_10680,N_3242,N_2427);
or U10681 (N_10681,N_4228,N_4160);
nor U10682 (N_10682,N_2969,N_4499);
or U10683 (N_10683,N_1411,N_847);
nand U10684 (N_10684,N_5754,N_4270);
nand U10685 (N_10685,N_2063,N_5243);
nor U10686 (N_10686,N_496,N_1842);
nor U10687 (N_10687,N_5953,N_5069);
xnor U10688 (N_10688,N_2905,N_5168);
nor U10689 (N_10689,N_1933,N_25);
and U10690 (N_10690,N_695,N_116);
or U10691 (N_10691,N_6091,N_2451);
and U10692 (N_10692,N_1231,N_5218);
or U10693 (N_10693,N_5989,N_2599);
xnor U10694 (N_10694,N_5193,N_4440);
xnor U10695 (N_10695,N_5131,N_2781);
and U10696 (N_10696,N_5362,N_4171);
nand U10697 (N_10697,N_1282,N_5788);
and U10698 (N_10698,N_1228,N_1305);
xor U10699 (N_10699,N_2921,N_5212);
xor U10700 (N_10700,N_1731,N_4364);
and U10701 (N_10701,N_3178,N_3774);
xor U10702 (N_10702,N_2547,N_5155);
or U10703 (N_10703,N_3607,N_4265);
xor U10704 (N_10704,N_1602,N_3623);
nand U10705 (N_10705,N_5291,N_5303);
nand U10706 (N_10706,N_5400,N_1513);
nand U10707 (N_10707,N_1661,N_4217);
nand U10708 (N_10708,N_132,N_466);
xor U10709 (N_10709,N_1135,N_1229);
xnor U10710 (N_10710,N_1748,N_5528);
nor U10711 (N_10711,N_4642,N_3633);
xor U10712 (N_10712,N_3290,N_1230);
nor U10713 (N_10713,N_3888,N_832);
xor U10714 (N_10714,N_3872,N_308);
xor U10715 (N_10715,N_5856,N_336);
or U10716 (N_10716,N_4855,N_1876);
nand U10717 (N_10717,N_247,N_5032);
and U10718 (N_10718,N_1901,N_1821);
xnor U10719 (N_10719,N_2745,N_618);
or U10720 (N_10720,N_2753,N_326);
or U10721 (N_10721,N_5588,N_5434);
nor U10722 (N_10722,N_5330,N_1998);
xor U10723 (N_10723,N_452,N_5132);
or U10724 (N_10724,N_5852,N_32);
xnor U10725 (N_10725,N_2403,N_5111);
xor U10726 (N_10726,N_4190,N_2703);
xnor U10727 (N_10727,N_4007,N_1402);
xnor U10728 (N_10728,N_4572,N_415);
xnor U10729 (N_10729,N_1788,N_5944);
or U10730 (N_10730,N_5719,N_4063);
and U10731 (N_10731,N_220,N_5291);
and U10732 (N_10732,N_880,N_3995);
xor U10733 (N_10733,N_4517,N_1550);
nor U10734 (N_10734,N_3101,N_500);
nor U10735 (N_10735,N_4165,N_6016);
nand U10736 (N_10736,N_3551,N_164);
nand U10737 (N_10737,N_434,N_5602);
nand U10738 (N_10738,N_2904,N_611);
or U10739 (N_10739,N_1227,N_1560);
nand U10740 (N_10740,N_6092,N_3390);
and U10741 (N_10741,N_3217,N_2564);
or U10742 (N_10742,N_4947,N_1104);
nand U10743 (N_10743,N_3743,N_2826);
nand U10744 (N_10744,N_239,N_3219);
xnor U10745 (N_10745,N_1455,N_2932);
or U10746 (N_10746,N_5133,N_5092);
and U10747 (N_10747,N_6140,N_189);
or U10748 (N_10748,N_2797,N_5886);
xnor U10749 (N_10749,N_986,N_1838);
and U10750 (N_10750,N_5497,N_2814);
or U10751 (N_10751,N_857,N_1533);
and U10752 (N_10752,N_5343,N_289);
nand U10753 (N_10753,N_891,N_6046);
or U10754 (N_10754,N_2258,N_5573);
and U10755 (N_10755,N_4150,N_4441);
and U10756 (N_10756,N_5546,N_4468);
nand U10757 (N_10757,N_1473,N_1475);
or U10758 (N_10758,N_3001,N_3642);
nand U10759 (N_10759,N_3121,N_692);
or U10760 (N_10760,N_2092,N_4266);
or U10761 (N_10761,N_382,N_4879);
and U10762 (N_10762,N_1744,N_4744);
xnor U10763 (N_10763,N_471,N_445);
nor U10764 (N_10764,N_1643,N_1875);
xnor U10765 (N_10765,N_3888,N_1227);
xor U10766 (N_10766,N_3022,N_3899);
and U10767 (N_10767,N_1076,N_3047);
and U10768 (N_10768,N_2471,N_1833);
nor U10769 (N_10769,N_3756,N_4872);
nor U10770 (N_10770,N_4466,N_1949);
and U10771 (N_10771,N_2309,N_2210);
and U10772 (N_10772,N_2413,N_3630);
or U10773 (N_10773,N_6206,N_3865);
and U10774 (N_10774,N_1234,N_924);
nand U10775 (N_10775,N_4377,N_2937);
nor U10776 (N_10776,N_1034,N_3384);
nor U10777 (N_10777,N_6010,N_1796);
xnor U10778 (N_10778,N_3818,N_999);
nand U10779 (N_10779,N_3252,N_2826);
xnor U10780 (N_10780,N_2817,N_5368);
nand U10781 (N_10781,N_3126,N_2103);
nor U10782 (N_10782,N_1837,N_3569);
nor U10783 (N_10783,N_5277,N_1161);
or U10784 (N_10784,N_1854,N_4651);
or U10785 (N_10785,N_3959,N_2234);
nor U10786 (N_10786,N_1584,N_1327);
nor U10787 (N_10787,N_703,N_4970);
xnor U10788 (N_10788,N_5195,N_130);
or U10789 (N_10789,N_4252,N_4778);
xor U10790 (N_10790,N_5026,N_4179);
or U10791 (N_10791,N_206,N_2192);
and U10792 (N_10792,N_576,N_2899);
or U10793 (N_10793,N_5959,N_5640);
or U10794 (N_10794,N_2009,N_3783);
or U10795 (N_10795,N_2653,N_5330);
nand U10796 (N_10796,N_2962,N_4792);
or U10797 (N_10797,N_4117,N_1816);
or U10798 (N_10798,N_3914,N_290);
nor U10799 (N_10799,N_4333,N_3244);
nand U10800 (N_10800,N_4087,N_3839);
or U10801 (N_10801,N_3806,N_1903);
nor U10802 (N_10802,N_14,N_316);
nand U10803 (N_10803,N_4510,N_1203);
xnor U10804 (N_10804,N_948,N_3835);
nand U10805 (N_10805,N_4372,N_1757);
nand U10806 (N_10806,N_6000,N_4692);
or U10807 (N_10807,N_6026,N_4167);
xor U10808 (N_10808,N_3807,N_4245);
nand U10809 (N_10809,N_1273,N_3060);
xor U10810 (N_10810,N_1773,N_1528);
xor U10811 (N_10811,N_6069,N_2099);
nand U10812 (N_10812,N_5852,N_4122);
and U10813 (N_10813,N_5672,N_3350);
and U10814 (N_10814,N_4012,N_610);
nor U10815 (N_10815,N_4428,N_610);
and U10816 (N_10816,N_5746,N_3501);
xor U10817 (N_10817,N_4816,N_4479);
or U10818 (N_10818,N_3864,N_5922);
or U10819 (N_10819,N_238,N_2185);
nand U10820 (N_10820,N_6200,N_3721);
nand U10821 (N_10821,N_3863,N_1299);
xor U10822 (N_10822,N_1649,N_2156);
nand U10823 (N_10823,N_2498,N_4188);
or U10824 (N_10824,N_578,N_419);
and U10825 (N_10825,N_5189,N_3329);
or U10826 (N_10826,N_2107,N_4489);
xnor U10827 (N_10827,N_2685,N_1852);
or U10828 (N_10828,N_3463,N_3993);
nand U10829 (N_10829,N_3918,N_2817);
nand U10830 (N_10830,N_1359,N_5155);
xor U10831 (N_10831,N_240,N_5341);
xor U10832 (N_10832,N_4816,N_3059);
or U10833 (N_10833,N_3283,N_5460);
nand U10834 (N_10834,N_2363,N_3983);
nor U10835 (N_10835,N_1009,N_3737);
or U10836 (N_10836,N_2324,N_1252);
or U10837 (N_10837,N_5874,N_2300);
or U10838 (N_10838,N_3024,N_4192);
nand U10839 (N_10839,N_5244,N_3271);
nand U10840 (N_10840,N_1832,N_5819);
or U10841 (N_10841,N_1533,N_6240);
nor U10842 (N_10842,N_5930,N_202);
nand U10843 (N_10843,N_1476,N_4383);
nand U10844 (N_10844,N_3838,N_3782);
and U10845 (N_10845,N_6089,N_5085);
and U10846 (N_10846,N_1578,N_5249);
and U10847 (N_10847,N_2235,N_5302);
nand U10848 (N_10848,N_2497,N_4920);
nor U10849 (N_10849,N_4329,N_1364);
or U10850 (N_10850,N_1735,N_5827);
and U10851 (N_10851,N_3449,N_6031);
xnor U10852 (N_10852,N_789,N_2141);
nand U10853 (N_10853,N_3628,N_2029);
nor U10854 (N_10854,N_1746,N_2686);
xor U10855 (N_10855,N_2332,N_6153);
and U10856 (N_10856,N_4840,N_4660);
or U10857 (N_10857,N_2206,N_2612);
or U10858 (N_10858,N_2219,N_261);
or U10859 (N_10859,N_2136,N_2496);
and U10860 (N_10860,N_5967,N_2618);
nand U10861 (N_10861,N_3666,N_1915);
nor U10862 (N_10862,N_5122,N_3226);
xnor U10863 (N_10863,N_5935,N_1284);
nor U10864 (N_10864,N_3422,N_991);
nand U10865 (N_10865,N_1754,N_4244);
xnor U10866 (N_10866,N_5439,N_384);
xor U10867 (N_10867,N_3672,N_1317);
or U10868 (N_10868,N_1473,N_2981);
nor U10869 (N_10869,N_4798,N_3835);
nor U10870 (N_10870,N_4889,N_92);
nor U10871 (N_10871,N_537,N_5427);
xnor U10872 (N_10872,N_3280,N_5825);
xnor U10873 (N_10873,N_3789,N_5650);
or U10874 (N_10874,N_809,N_2087);
nor U10875 (N_10875,N_1932,N_454);
and U10876 (N_10876,N_857,N_1837);
or U10877 (N_10877,N_5329,N_3990);
nand U10878 (N_10878,N_2210,N_1252);
xor U10879 (N_10879,N_4336,N_5016);
nand U10880 (N_10880,N_2289,N_71);
nand U10881 (N_10881,N_5302,N_810);
nor U10882 (N_10882,N_2703,N_2071);
nor U10883 (N_10883,N_5390,N_2594);
and U10884 (N_10884,N_6074,N_6124);
nor U10885 (N_10885,N_1144,N_995);
xor U10886 (N_10886,N_3412,N_2061);
nand U10887 (N_10887,N_3028,N_4334);
nor U10888 (N_10888,N_2135,N_4481);
and U10889 (N_10889,N_2125,N_1780);
and U10890 (N_10890,N_5026,N_6033);
nand U10891 (N_10891,N_1539,N_4265);
nor U10892 (N_10892,N_4009,N_3715);
nor U10893 (N_10893,N_4517,N_2514);
nand U10894 (N_10894,N_2560,N_2361);
nand U10895 (N_10895,N_6141,N_1046);
nor U10896 (N_10896,N_1553,N_2255);
and U10897 (N_10897,N_4589,N_4712);
nor U10898 (N_10898,N_3259,N_1090);
or U10899 (N_10899,N_1591,N_2470);
nand U10900 (N_10900,N_832,N_5424);
nand U10901 (N_10901,N_4061,N_669);
xor U10902 (N_10902,N_3263,N_4990);
and U10903 (N_10903,N_64,N_4730);
and U10904 (N_10904,N_2623,N_2220);
nor U10905 (N_10905,N_1261,N_5147);
xnor U10906 (N_10906,N_514,N_2412);
xor U10907 (N_10907,N_571,N_3444);
xnor U10908 (N_10908,N_4236,N_5974);
and U10909 (N_10909,N_5305,N_6084);
nor U10910 (N_10910,N_104,N_5450);
nor U10911 (N_10911,N_1583,N_3372);
nand U10912 (N_10912,N_381,N_1282);
or U10913 (N_10913,N_5791,N_3614);
nand U10914 (N_10914,N_2575,N_2900);
xnor U10915 (N_10915,N_632,N_611);
or U10916 (N_10916,N_2522,N_625);
or U10917 (N_10917,N_1171,N_481);
and U10918 (N_10918,N_5590,N_3635);
nand U10919 (N_10919,N_2856,N_481);
nor U10920 (N_10920,N_5342,N_1864);
nand U10921 (N_10921,N_5945,N_3367);
nor U10922 (N_10922,N_5551,N_1756);
xor U10923 (N_10923,N_4992,N_5634);
nand U10924 (N_10924,N_2854,N_1708);
and U10925 (N_10925,N_3790,N_5870);
nand U10926 (N_10926,N_5690,N_5042);
nand U10927 (N_10927,N_2469,N_1012);
or U10928 (N_10928,N_3072,N_5391);
nand U10929 (N_10929,N_3791,N_5622);
or U10930 (N_10930,N_477,N_5368);
xor U10931 (N_10931,N_4853,N_3792);
or U10932 (N_10932,N_5486,N_4902);
and U10933 (N_10933,N_5735,N_524);
nand U10934 (N_10934,N_2808,N_1716);
nand U10935 (N_10935,N_3931,N_6187);
xor U10936 (N_10936,N_879,N_5027);
and U10937 (N_10937,N_1910,N_3593);
and U10938 (N_10938,N_4396,N_5935);
nor U10939 (N_10939,N_2890,N_6011);
nor U10940 (N_10940,N_1977,N_762);
nand U10941 (N_10941,N_5037,N_4708);
nand U10942 (N_10942,N_2244,N_1528);
and U10943 (N_10943,N_1356,N_481);
nand U10944 (N_10944,N_1754,N_888);
nor U10945 (N_10945,N_4397,N_2128);
xnor U10946 (N_10946,N_1075,N_5921);
xnor U10947 (N_10947,N_3497,N_1873);
or U10948 (N_10948,N_666,N_4423);
nor U10949 (N_10949,N_2915,N_2415);
or U10950 (N_10950,N_132,N_2663);
nor U10951 (N_10951,N_4798,N_5652);
or U10952 (N_10952,N_5177,N_2430);
or U10953 (N_10953,N_706,N_482);
or U10954 (N_10954,N_2418,N_1053);
or U10955 (N_10955,N_2164,N_2646);
and U10956 (N_10956,N_2643,N_5630);
nor U10957 (N_10957,N_691,N_1545);
and U10958 (N_10958,N_5008,N_841);
nand U10959 (N_10959,N_6181,N_4265);
xor U10960 (N_10960,N_3534,N_5872);
nor U10961 (N_10961,N_555,N_287);
or U10962 (N_10962,N_1770,N_1267);
nor U10963 (N_10963,N_2058,N_609);
nand U10964 (N_10964,N_5475,N_2008);
nand U10965 (N_10965,N_4048,N_4520);
and U10966 (N_10966,N_3076,N_2597);
xnor U10967 (N_10967,N_5572,N_2016);
or U10968 (N_10968,N_2063,N_4080);
and U10969 (N_10969,N_2843,N_5216);
or U10970 (N_10970,N_2765,N_2912);
and U10971 (N_10971,N_257,N_23);
nand U10972 (N_10972,N_399,N_5930);
xnor U10973 (N_10973,N_3520,N_5786);
nor U10974 (N_10974,N_681,N_5500);
and U10975 (N_10975,N_1746,N_5387);
and U10976 (N_10976,N_5453,N_5788);
nor U10977 (N_10977,N_1760,N_5266);
xnor U10978 (N_10978,N_942,N_4048);
xnor U10979 (N_10979,N_4610,N_1233);
and U10980 (N_10980,N_2759,N_1171);
or U10981 (N_10981,N_2330,N_3265);
xnor U10982 (N_10982,N_4209,N_4499);
or U10983 (N_10983,N_1449,N_3020);
or U10984 (N_10984,N_2428,N_1055);
xor U10985 (N_10985,N_36,N_1384);
xnor U10986 (N_10986,N_4759,N_3892);
and U10987 (N_10987,N_2717,N_2053);
nand U10988 (N_10988,N_5497,N_2612);
xor U10989 (N_10989,N_688,N_4991);
nor U10990 (N_10990,N_1206,N_2298);
and U10991 (N_10991,N_1844,N_1472);
xor U10992 (N_10992,N_3092,N_360);
xor U10993 (N_10993,N_3732,N_516);
nand U10994 (N_10994,N_644,N_5939);
nand U10995 (N_10995,N_2783,N_5323);
or U10996 (N_10996,N_4998,N_1929);
xor U10997 (N_10997,N_2479,N_1328);
xor U10998 (N_10998,N_2629,N_4834);
xor U10999 (N_10999,N_2291,N_2430);
and U11000 (N_11000,N_6237,N_339);
and U11001 (N_11001,N_4168,N_814);
nor U11002 (N_11002,N_1126,N_522);
and U11003 (N_11003,N_5804,N_4289);
or U11004 (N_11004,N_5477,N_1724);
nor U11005 (N_11005,N_3179,N_5030);
nand U11006 (N_11006,N_854,N_118);
xor U11007 (N_11007,N_5854,N_2417);
and U11008 (N_11008,N_1867,N_6048);
or U11009 (N_11009,N_2259,N_2738);
or U11010 (N_11010,N_5160,N_5379);
or U11011 (N_11011,N_1011,N_3303);
xor U11012 (N_11012,N_672,N_2148);
nand U11013 (N_11013,N_5343,N_5840);
or U11014 (N_11014,N_670,N_317);
or U11015 (N_11015,N_3407,N_2803);
nor U11016 (N_11016,N_4811,N_3296);
nor U11017 (N_11017,N_1566,N_1488);
nand U11018 (N_11018,N_4451,N_4366);
and U11019 (N_11019,N_1279,N_60);
or U11020 (N_11020,N_5647,N_724);
and U11021 (N_11021,N_1535,N_1214);
xor U11022 (N_11022,N_1006,N_4515);
xnor U11023 (N_11023,N_1033,N_3774);
nand U11024 (N_11024,N_2523,N_1641);
or U11025 (N_11025,N_743,N_3980);
or U11026 (N_11026,N_2545,N_1511);
or U11027 (N_11027,N_3168,N_4981);
nand U11028 (N_11028,N_808,N_2707);
nor U11029 (N_11029,N_2570,N_1484);
nor U11030 (N_11030,N_154,N_2523);
nor U11031 (N_11031,N_1459,N_2195);
and U11032 (N_11032,N_1621,N_395);
nor U11033 (N_11033,N_5623,N_2924);
nand U11034 (N_11034,N_6138,N_934);
xor U11035 (N_11035,N_1200,N_112);
nor U11036 (N_11036,N_2891,N_5719);
and U11037 (N_11037,N_4801,N_690);
nor U11038 (N_11038,N_5508,N_4368);
or U11039 (N_11039,N_4734,N_2849);
or U11040 (N_11040,N_3793,N_1945);
nand U11041 (N_11041,N_1565,N_2828);
or U11042 (N_11042,N_5187,N_6032);
nand U11043 (N_11043,N_461,N_5458);
or U11044 (N_11044,N_4431,N_6039);
or U11045 (N_11045,N_232,N_3410);
xor U11046 (N_11046,N_4077,N_2124);
nand U11047 (N_11047,N_3856,N_430);
nor U11048 (N_11048,N_2628,N_5487);
nor U11049 (N_11049,N_4341,N_5644);
or U11050 (N_11050,N_4747,N_309);
nor U11051 (N_11051,N_4929,N_6221);
xnor U11052 (N_11052,N_4066,N_1303);
nor U11053 (N_11053,N_1159,N_4807);
and U11054 (N_11054,N_5210,N_3072);
xnor U11055 (N_11055,N_3913,N_263);
nor U11056 (N_11056,N_1728,N_1639);
xor U11057 (N_11057,N_4856,N_5466);
xor U11058 (N_11058,N_4003,N_4779);
and U11059 (N_11059,N_3037,N_5144);
or U11060 (N_11060,N_1711,N_3204);
xnor U11061 (N_11061,N_5062,N_1183);
xnor U11062 (N_11062,N_2416,N_1716);
and U11063 (N_11063,N_2147,N_3736);
nor U11064 (N_11064,N_353,N_5344);
and U11065 (N_11065,N_3672,N_16);
and U11066 (N_11066,N_2964,N_5283);
nand U11067 (N_11067,N_5483,N_1878);
and U11068 (N_11068,N_5477,N_1596);
or U11069 (N_11069,N_4065,N_4614);
nor U11070 (N_11070,N_1642,N_4473);
or U11071 (N_11071,N_2158,N_4845);
nand U11072 (N_11072,N_3035,N_3893);
or U11073 (N_11073,N_6059,N_56);
nand U11074 (N_11074,N_519,N_4579);
and U11075 (N_11075,N_5357,N_514);
nor U11076 (N_11076,N_4374,N_1006);
nand U11077 (N_11077,N_2358,N_690);
xnor U11078 (N_11078,N_5828,N_1612);
xnor U11079 (N_11079,N_2658,N_5088);
or U11080 (N_11080,N_2523,N_3794);
xor U11081 (N_11081,N_3966,N_4887);
nand U11082 (N_11082,N_6107,N_1535);
nor U11083 (N_11083,N_525,N_5623);
xor U11084 (N_11084,N_4556,N_556);
or U11085 (N_11085,N_2647,N_2944);
or U11086 (N_11086,N_5111,N_3590);
or U11087 (N_11087,N_1649,N_3516);
or U11088 (N_11088,N_3534,N_3754);
or U11089 (N_11089,N_4950,N_5316);
and U11090 (N_11090,N_2034,N_4210);
nor U11091 (N_11091,N_3771,N_4918);
nand U11092 (N_11092,N_1932,N_3807);
and U11093 (N_11093,N_3289,N_2663);
and U11094 (N_11094,N_5227,N_1683);
or U11095 (N_11095,N_2163,N_1472);
nor U11096 (N_11096,N_5052,N_131);
xnor U11097 (N_11097,N_5751,N_1462);
nand U11098 (N_11098,N_3510,N_3729);
nor U11099 (N_11099,N_3622,N_395);
nor U11100 (N_11100,N_495,N_432);
xor U11101 (N_11101,N_1276,N_5929);
nand U11102 (N_11102,N_273,N_3220);
or U11103 (N_11103,N_2647,N_4640);
nand U11104 (N_11104,N_3844,N_2012);
xor U11105 (N_11105,N_5621,N_3954);
and U11106 (N_11106,N_5938,N_3568);
xor U11107 (N_11107,N_3675,N_4456);
and U11108 (N_11108,N_3687,N_6189);
or U11109 (N_11109,N_1398,N_5580);
or U11110 (N_11110,N_5457,N_6202);
nand U11111 (N_11111,N_4865,N_4514);
nor U11112 (N_11112,N_4130,N_752);
xnor U11113 (N_11113,N_4607,N_1764);
or U11114 (N_11114,N_3401,N_5244);
nand U11115 (N_11115,N_3350,N_1875);
nand U11116 (N_11116,N_6236,N_3833);
nor U11117 (N_11117,N_635,N_5797);
or U11118 (N_11118,N_4354,N_2411);
nand U11119 (N_11119,N_836,N_5309);
xnor U11120 (N_11120,N_2199,N_4835);
nor U11121 (N_11121,N_1579,N_5434);
nand U11122 (N_11122,N_4215,N_3818);
nor U11123 (N_11123,N_5822,N_4996);
xnor U11124 (N_11124,N_3957,N_5445);
nand U11125 (N_11125,N_1230,N_2358);
nand U11126 (N_11126,N_4857,N_1955);
nor U11127 (N_11127,N_4960,N_5254);
xor U11128 (N_11128,N_2827,N_4509);
nand U11129 (N_11129,N_5603,N_1564);
xnor U11130 (N_11130,N_1730,N_1815);
or U11131 (N_11131,N_3798,N_4700);
xor U11132 (N_11132,N_311,N_2319);
or U11133 (N_11133,N_1042,N_2095);
and U11134 (N_11134,N_3485,N_3522);
and U11135 (N_11135,N_4198,N_6072);
xor U11136 (N_11136,N_3134,N_3713);
or U11137 (N_11137,N_5603,N_4960);
nor U11138 (N_11138,N_603,N_5877);
nand U11139 (N_11139,N_4512,N_4370);
or U11140 (N_11140,N_4075,N_2364);
nand U11141 (N_11141,N_4840,N_2776);
or U11142 (N_11142,N_4484,N_139);
nand U11143 (N_11143,N_4572,N_1478);
nand U11144 (N_11144,N_3232,N_905);
nor U11145 (N_11145,N_3739,N_4760);
xnor U11146 (N_11146,N_5221,N_230);
or U11147 (N_11147,N_5915,N_1997);
xor U11148 (N_11148,N_4663,N_4516);
or U11149 (N_11149,N_157,N_3454);
or U11150 (N_11150,N_5364,N_2036);
and U11151 (N_11151,N_1831,N_1715);
nor U11152 (N_11152,N_4878,N_3116);
or U11153 (N_11153,N_3235,N_307);
and U11154 (N_11154,N_3175,N_2140);
or U11155 (N_11155,N_3079,N_5750);
or U11156 (N_11156,N_5722,N_6071);
xor U11157 (N_11157,N_4450,N_153);
or U11158 (N_11158,N_3324,N_1211);
and U11159 (N_11159,N_4718,N_3718);
nor U11160 (N_11160,N_2171,N_5953);
or U11161 (N_11161,N_35,N_204);
nand U11162 (N_11162,N_5384,N_6175);
xnor U11163 (N_11163,N_1331,N_1519);
and U11164 (N_11164,N_586,N_6107);
or U11165 (N_11165,N_4349,N_1161);
nand U11166 (N_11166,N_1515,N_3801);
nand U11167 (N_11167,N_3433,N_1398);
and U11168 (N_11168,N_4886,N_276);
nand U11169 (N_11169,N_193,N_3139);
or U11170 (N_11170,N_6181,N_4389);
or U11171 (N_11171,N_372,N_427);
nand U11172 (N_11172,N_1065,N_6153);
xnor U11173 (N_11173,N_1489,N_3649);
nand U11174 (N_11174,N_1140,N_4231);
nor U11175 (N_11175,N_5733,N_3330);
and U11176 (N_11176,N_4816,N_1483);
or U11177 (N_11177,N_2211,N_2455);
nand U11178 (N_11178,N_296,N_5550);
nand U11179 (N_11179,N_1422,N_5412);
nor U11180 (N_11180,N_3601,N_375);
xor U11181 (N_11181,N_4229,N_2700);
nor U11182 (N_11182,N_2956,N_6205);
xnor U11183 (N_11183,N_2527,N_2747);
nor U11184 (N_11184,N_1122,N_801);
xnor U11185 (N_11185,N_5427,N_5338);
nor U11186 (N_11186,N_5979,N_2156);
nand U11187 (N_11187,N_1800,N_5256);
xnor U11188 (N_11188,N_415,N_1360);
or U11189 (N_11189,N_2371,N_1076);
xor U11190 (N_11190,N_6023,N_4056);
or U11191 (N_11191,N_3548,N_2678);
xor U11192 (N_11192,N_3447,N_2541);
xor U11193 (N_11193,N_3935,N_3937);
and U11194 (N_11194,N_2031,N_1923);
xor U11195 (N_11195,N_2236,N_6114);
nor U11196 (N_11196,N_1458,N_1254);
nor U11197 (N_11197,N_3692,N_4083);
nand U11198 (N_11198,N_5437,N_6075);
or U11199 (N_11199,N_855,N_5854);
nor U11200 (N_11200,N_3634,N_3617);
nor U11201 (N_11201,N_2146,N_3066);
nor U11202 (N_11202,N_3496,N_3693);
and U11203 (N_11203,N_5970,N_2511);
or U11204 (N_11204,N_353,N_4181);
and U11205 (N_11205,N_4833,N_2746);
and U11206 (N_11206,N_2902,N_3058);
nand U11207 (N_11207,N_445,N_1241);
and U11208 (N_11208,N_2030,N_1463);
and U11209 (N_11209,N_518,N_4207);
or U11210 (N_11210,N_2689,N_6081);
xor U11211 (N_11211,N_3985,N_2718);
or U11212 (N_11212,N_5747,N_3975);
and U11213 (N_11213,N_195,N_1876);
xnor U11214 (N_11214,N_2095,N_4179);
and U11215 (N_11215,N_2676,N_5478);
nor U11216 (N_11216,N_1458,N_2507);
nand U11217 (N_11217,N_3782,N_3684);
nor U11218 (N_11218,N_2712,N_1495);
nor U11219 (N_11219,N_2179,N_1848);
nand U11220 (N_11220,N_2936,N_5134);
or U11221 (N_11221,N_3918,N_171);
xnor U11222 (N_11222,N_4451,N_605);
or U11223 (N_11223,N_3533,N_3646);
or U11224 (N_11224,N_4617,N_262);
or U11225 (N_11225,N_3010,N_2531);
or U11226 (N_11226,N_3008,N_2384);
nand U11227 (N_11227,N_4857,N_746);
or U11228 (N_11228,N_1437,N_4732);
or U11229 (N_11229,N_2678,N_2358);
and U11230 (N_11230,N_1570,N_1848);
xor U11231 (N_11231,N_2629,N_1618);
or U11232 (N_11232,N_5673,N_1890);
nand U11233 (N_11233,N_1042,N_3581);
nor U11234 (N_11234,N_452,N_3357);
nand U11235 (N_11235,N_5227,N_928);
and U11236 (N_11236,N_2742,N_2311);
nor U11237 (N_11237,N_3907,N_3232);
nor U11238 (N_11238,N_404,N_3034);
or U11239 (N_11239,N_1027,N_1418);
and U11240 (N_11240,N_4408,N_4789);
and U11241 (N_11241,N_5290,N_3503);
nand U11242 (N_11242,N_1779,N_4557);
xor U11243 (N_11243,N_1773,N_1608);
or U11244 (N_11244,N_1736,N_776);
or U11245 (N_11245,N_834,N_4235);
or U11246 (N_11246,N_4498,N_3603);
or U11247 (N_11247,N_550,N_38);
and U11248 (N_11248,N_2983,N_77);
nand U11249 (N_11249,N_2353,N_4058);
xnor U11250 (N_11250,N_4408,N_2720);
xnor U11251 (N_11251,N_5567,N_6096);
and U11252 (N_11252,N_1336,N_5705);
and U11253 (N_11253,N_1119,N_3602);
xnor U11254 (N_11254,N_4170,N_4738);
and U11255 (N_11255,N_4639,N_4572);
nor U11256 (N_11256,N_5778,N_674);
xnor U11257 (N_11257,N_1185,N_5389);
nor U11258 (N_11258,N_2195,N_3718);
xnor U11259 (N_11259,N_685,N_2705);
and U11260 (N_11260,N_4147,N_3455);
xnor U11261 (N_11261,N_5233,N_663);
and U11262 (N_11262,N_5425,N_2468);
nand U11263 (N_11263,N_881,N_3395);
or U11264 (N_11264,N_4857,N_1302);
nand U11265 (N_11265,N_4995,N_451);
or U11266 (N_11266,N_5754,N_4461);
nand U11267 (N_11267,N_792,N_4711);
or U11268 (N_11268,N_4092,N_6126);
nand U11269 (N_11269,N_2133,N_1926);
and U11270 (N_11270,N_3207,N_1711);
xnor U11271 (N_11271,N_4954,N_3240);
or U11272 (N_11272,N_4620,N_4828);
nor U11273 (N_11273,N_5196,N_3899);
nor U11274 (N_11274,N_1221,N_3808);
xor U11275 (N_11275,N_4689,N_1279);
or U11276 (N_11276,N_5441,N_1335);
xnor U11277 (N_11277,N_1914,N_4613);
and U11278 (N_11278,N_511,N_2009);
nand U11279 (N_11279,N_5370,N_5417);
nor U11280 (N_11280,N_3200,N_6246);
xor U11281 (N_11281,N_1,N_4521);
and U11282 (N_11282,N_4089,N_3047);
nor U11283 (N_11283,N_4479,N_1430);
nor U11284 (N_11284,N_2061,N_2451);
xnor U11285 (N_11285,N_5336,N_3539);
and U11286 (N_11286,N_2721,N_1890);
xor U11287 (N_11287,N_2652,N_3537);
nand U11288 (N_11288,N_4715,N_424);
nand U11289 (N_11289,N_5211,N_5236);
xnor U11290 (N_11290,N_2571,N_5778);
and U11291 (N_11291,N_3301,N_5633);
xnor U11292 (N_11292,N_1175,N_2745);
nand U11293 (N_11293,N_2328,N_2013);
or U11294 (N_11294,N_943,N_2221);
and U11295 (N_11295,N_3031,N_99);
nand U11296 (N_11296,N_1868,N_2560);
xor U11297 (N_11297,N_3545,N_2159);
nand U11298 (N_11298,N_1435,N_1605);
nand U11299 (N_11299,N_1548,N_2725);
nand U11300 (N_11300,N_557,N_3937);
xor U11301 (N_11301,N_1467,N_3446);
xor U11302 (N_11302,N_1641,N_4598);
xnor U11303 (N_11303,N_1539,N_3964);
nand U11304 (N_11304,N_6037,N_930);
xor U11305 (N_11305,N_5828,N_3671);
xnor U11306 (N_11306,N_2988,N_5815);
or U11307 (N_11307,N_3620,N_5174);
nor U11308 (N_11308,N_1434,N_172);
nor U11309 (N_11309,N_6186,N_5245);
and U11310 (N_11310,N_4304,N_3906);
and U11311 (N_11311,N_8,N_4526);
xor U11312 (N_11312,N_2015,N_4551);
or U11313 (N_11313,N_92,N_6002);
nor U11314 (N_11314,N_5183,N_4763);
or U11315 (N_11315,N_1216,N_1007);
nand U11316 (N_11316,N_2091,N_5805);
nand U11317 (N_11317,N_1304,N_2935);
xor U11318 (N_11318,N_2998,N_1118);
nand U11319 (N_11319,N_5002,N_5590);
nor U11320 (N_11320,N_2507,N_2274);
nand U11321 (N_11321,N_1815,N_4234);
xor U11322 (N_11322,N_1138,N_4724);
and U11323 (N_11323,N_98,N_1407);
and U11324 (N_11324,N_3041,N_4240);
xor U11325 (N_11325,N_2885,N_207);
and U11326 (N_11326,N_4279,N_2859);
xnor U11327 (N_11327,N_4121,N_5889);
xnor U11328 (N_11328,N_1897,N_2209);
xnor U11329 (N_11329,N_5692,N_1344);
nand U11330 (N_11330,N_1763,N_1410);
nor U11331 (N_11331,N_2244,N_133);
or U11332 (N_11332,N_5244,N_3993);
nor U11333 (N_11333,N_3163,N_3550);
nand U11334 (N_11334,N_1186,N_988);
xor U11335 (N_11335,N_4161,N_2559);
and U11336 (N_11336,N_5494,N_3975);
xnor U11337 (N_11337,N_852,N_6178);
nand U11338 (N_11338,N_5130,N_1179);
xnor U11339 (N_11339,N_1617,N_4414);
xor U11340 (N_11340,N_2379,N_5133);
xnor U11341 (N_11341,N_1362,N_2203);
or U11342 (N_11342,N_1024,N_5102);
nor U11343 (N_11343,N_6220,N_2632);
xor U11344 (N_11344,N_3238,N_1502);
and U11345 (N_11345,N_4618,N_1617);
nor U11346 (N_11346,N_4177,N_2290);
nor U11347 (N_11347,N_1362,N_3176);
and U11348 (N_11348,N_4609,N_626);
nand U11349 (N_11349,N_4582,N_2412);
nor U11350 (N_11350,N_3326,N_3343);
xnor U11351 (N_11351,N_4205,N_5202);
nor U11352 (N_11352,N_173,N_4567);
or U11353 (N_11353,N_4803,N_644);
xnor U11354 (N_11354,N_8,N_3332);
or U11355 (N_11355,N_3461,N_3480);
or U11356 (N_11356,N_3732,N_1764);
and U11357 (N_11357,N_5567,N_5008);
and U11358 (N_11358,N_2095,N_4106);
nor U11359 (N_11359,N_2343,N_880);
nor U11360 (N_11360,N_610,N_4285);
nor U11361 (N_11361,N_1077,N_4622);
or U11362 (N_11362,N_6187,N_1922);
or U11363 (N_11363,N_2166,N_156);
nand U11364 (N_11364,N_1012,N_899);
nor U11365 (N_11365,N_2106,N_3794);
xnor U11366 (N_11366,N_5372,N_572);
xnor U11367 (N_11367,N_4055,N_5437);
nand U11368 (N_11368,N_2754,N_1029);
and U11369 (N_11369,N_4045,N_1785);
or U11370 (N_11370,N_2662,N_1225);
or U11371 (N_11371,N_3932,N_5210);
xor U11372 (N_11372,N_422,N_5522);
and U11373 (N_11373,N_3157,N_5531);
and U11374 (N_11374,N_1553,N_1631);
nor U11375 (N_11375,N_1501,N_3802);
nand U11376 (N_11376,N_5044,N_2868);
nand U11377 (N_11377,N_5197,N_5699);
and U11378 (N_11378,N_1548,N_2316);
and U11379 (N_11379,N_5142,N_5959);
nor U11380 (N_11380,N_4057,N_3308);
and U11381 (N_11381,N_3235,N_4881);
nor U11382 (N_11382,N_4492,N_2344);
xnor U11383 (N_11383,N_1274,N_6119);
xor U11384 (N_11384,N_5007,N_2350);
nor U11385 (N_11385,N_1301,N_2187);
and U11386 (N_11386,N_1935,N_4932);
or U11387 (N_11387,N_4477,N_3544);
nor U11388 (N_11388,N_440,N_2665);
nand U11389 (N_11389,N_4286,N_5564);
and U11390 (N_11390,N_2736,N_4737);
xor U11391 (N_11391,N_1506,N_6095);
or U11392 (N_11392,N_469,N_850);
xnor U11393 (N_11393,N_2007,N_900);
and U11394 (N_11394,N_693,N_5403);
xor U11395 (N_11395,N_1069,N_4742);
and U11396 (N_11396,N_3152,N_4894);
nor U11397 (N_11397,N_2914,N_1504);
xnor U11398 (N_11398,N_1872,N_1411);
or U11399 (N_11399,N_822,N_3641);
or U11400 (N_11400,N_5211,N_1982);
nand U11401 (N_11401,N_4244,N_1645);
xnor U11402 (N_11402,N_4345,N_4777);
nand U11403 (N_11403,N_4418,N_2366);
nand U11404 (N_11404,N_109,N_3870);
xor U11405 (N_11405,N_4920,N_33);
and U11406 (N_11406,N_6214,N_4406);
and U11407 (N_11407,N_5009,N_2718);
or U11408 (N_11408,N_1243,N_4078);
nand U11409 (N_11409,N_4871,N_4727);
xor U11410 (N_11410,N_4619,N_4028);
nand U11411 (N_11411,N_5729,N_4763);
and U11412 (N_11412,N_4327,N_3323);
nand U11413 (N_11413,N_4891,N_6010);
xnor U11414 (N_11414,N_4471,N_4498);
and U11415 (N_11415,N_2121,N_5700);
nor U11416 (N_11416,N_4434,N_418);
xor U11417 (N_11417,N_4881,N_3151);
nand U11418 (N_11418,N_634,N_1058);
nand U11419 (N_11419,N_3203,N_5904);
and U11420 (N_11420,N_3442,N_6235);
xnor U11421 (N_11421,N_6206,N_3621);
or U11422 (N_11422,N_3611,N_585);
xnor U11423 (N_11423,N_5087,N_178);
xnor U11424 (N_11424,N_295,N_516);
nor U11425 (N_11425,N_1425,N_3405);
nor U11426 (N_11426,N_2488,N_477);
nor U11427 (N_11427,N_3727,N_6070);
nor U11428 (N_11428,N_3412,N_933);
or U11429 (N_11429,N_2796,N_1132);
and U11430 (N_11430,N_2165,N_4249);
xor U11431 (N_11431,N_2794,N_1589);
xor U11432 (N_11432,N_5281,N_4254);
nand U11433 (N_11433,N_4344,N_5516);
nand U11434 (N_11434,N_4435,N_4848);
and U11435 (N_11435,N_5594,N_6212);
nand U11436 (N_11436,N_1433,N_3231);
or U11437 (N_11437,N_5395,N_86);
nor U11438 (N_11438,N_5712,N_3797);
and U11439 (N_11439,N_3298,N_3245);
and U11440 (N_11440,N_4862,N_5606);
nor U11441 (N_11441,N_5679,N_5766);
xor U11442 (N_11442,N_4094,N_5236);
nand U11443 (N_11443,N_1108,N_387);
xnor U11444 (N_11444,N_24,N_5319);
xnor U11445 (N_11445,N_1687,N_5563);
and U11446 (N_11446,N_4113,N_3435);
xnor U11447 (N_11447,N_1326,N_2144);
nand U11448 (N_11448,N_4278,N_3376);
and U11449 (N_11449,N_4549,N_4485);
or U11450 (N_11450,N_5234,N_3067);
and U11451 (N_11451,N_1295,N_2071);
nor U11452 (N_11452,N_2506,N_4027);
and U11453 (N_11453,N_5000,N_979);
xor U11454 (N_11454,N_4692,N_4307);
nor U11455 (N_11455,N_4319,N_3934);
nand U11456 (N_11456,N_1288,N_1453);
nor U11457 (N_11457,N_2864,N_5930);
nand U11458 (N_11458,N_5030,N_368);
or U11459 (N_11459,N_2909,N_1428);
xor U11460 (N_11460,N_2733,N_5775);
and U11461 (N_11461,N_4707,N_4284);
nand U11462 (N_11462,N_1773,N_5373);
and U11463 (N_11463,N_5939,N_4696);
xnor U11464 (N_11464,N_4757,N_5423);
or U11465 (N_11465,N_1290,N_1998);
and U11466 (N_11466,N_1821,N_1150);
nand U11467 (N_11467,N_1107,N_1469);
xor U11468 (N_11468,N_2188,N_3266);
nor U11469 (N_11469,N_3467,N_4648);
and U11470 (N_11470,N_6019,N_1759);
nand U11471 (N_11471,N_902,N_6073);
or U11472 (N_11472,N_3575,N_6081);
or U11473 (N_11473,N_6032,N_3831);
nand U11474 (N_11474,N_1479,N_3850);
and U11475 (N_11475,N_3265,N_1242);
xnor U11476 (N_11476,N_4501,N_2385);
xor U11477 (N_11477,N_4130,N_3388);
nor U11478 (N_11478,N_3563,N_4296);
nor U11479 (N_11479,N_2103,N_3449);
and U11480 (N_11480,N_2080,N_753);
or U11481 (N_11481,N_5493,N_3284);
or U11482 (N_11482,N_689,N_2289);
nand U11483 (N_11483,N_5830,N_6054);
xnor U11484 (N_11484,N_373,N_4208);
and U11485 (N_11485,N_2743,N_6045);
or U11486 (N_11486,N_1940,N_2654);
and U11487 (N_11487,N_4478,N_5257);
xnor U11488 (N_11488,N_4489,N_890);
nand U11489 (N_11489,N_2564,N_4911);
nor U11490 (N_11490,N_4531,N_6016);
and U11491 (N_11491,N_522,N_4679);
nor U11492 (N_11492,N_1341,N_5895);
nand U11493 (N_11493,N_6071,N_1237);
or U11494 (N_11494,N_1174,N_1748);
xor U11495 (N_11495,N_1946,N_7);
xnor U11496 (N_11496,N_4148,N_605);
xor U11497 (N_11497,N_4387,N_3439);
and U11498 (N_11498,N_3859,N_3941);
nand U11499 (N_11499,N_112,N_5408);
nor U11500 (N_11500,N_4250,N_535);
nor U11501 (N_11501,N_5139,N_182);
and U11502 (N_11502,N_2207,N_3281);
or U11503 (N_11503,N_6071,N_4405);
nand U11504 (N_11504,N_2176,N_1389);
nor U11505 (N_11505,N_5040,N_4581);
nor U11506 (N_11506,N_3858,N_6054);
nand U11507 (N_11507,N_5653,N_5470);
and U11508 (N_11508,N_5140,N_5636);
or U11509 (N_11509,N_2967,N_4315);
and U11510 (N_11510,N_4427,N_1794);
xnor U11511 (N_11511,N_1636,N_4856);
xor U11512 (N_11512,N_4438,N_5480);
or U11513 (N_11513,N_3532,N_2928);
or U11514 (N_11514,N_1243,N_3092);
nand U11515 (N_11515,N_4581,N_5123);
xnor U11516 (N_11516,N_550,N_5328);
nand U11517 (N_11517,N_1130,N_2075);
and U11518 (N_11518,N_879,N_5362);
nor U11519 (N_11519,N_893,N_1526);
or U11520 (N_11520,N_6146,N_5634);
nor U11521 (N_11521,N_4037,N_3628);
nor U11522 (N_11522,N_5099,N_176);
xnor U11523 (N_11523,N_574,N_2455);
nand U11524 (N_11524,N_2854,N_2820);
nand U11525 (N_11525,N_2583,N_1957);
xor U11526 (N_11526,N_1629,N_315);
xnor U11527 (N_11527,N_3865,N_3578);
nand U11528 (N_11528,N_3122,N_2287);
and U11529 (N_11529,N_5507,N_6168);
nor U11530 (N_11530,N_499,N_6180);
and U11531 (N_11531,N_1093,N_2977);
nor U11532 (N_11532,N_4843,N_264);
nand U11533 (N_11533,N_2939,N_5843);
and U11534 (N_11534,N_1366,N_4924);
nand U11535 (N_11535,N_5826,N_2788);
xnor U11536 (N_11536,N_5648,N_2349);
and U11537 (N_11537,N_1247,N_6225);
nor U11538 (N_11538,N_2819,N_2926);
xor U11539 (N_11539,N_6207,N_1155);
or U11540 (N_11540,N_1716,N_810);
nor U11541 (N_11541,N_5670,N_2555);
nand U11542 (N_11542,N_4499,N_6207);
xor U11543 (N_11543,N_692,N_3242);
xnor U11544 (N_11544,N_4577,N_198);
or U11545 (N_11545,N_895,N_952);
nor U11546 (N_11546,N_4330,N_4916);
and U11547 (N_11547,N_3890,N_4265);
nand U11548 (N_11548,N_2207,N_4178);
nor U11549 (N_11549,N_3081,N_2467);
and U11550 (N_11550,N_1273,N_4173);
nand U11551 (N_11551,N_1898,N_5098);
nor U11552 (N_11552,N_2904,N_1725);
nand U11553 (N_11553,N_6042,N_5085);
nand U11554 (N_11554,N_5653,N_4910);
nand U11555 (N_11555,N_982,N_4492);
nand U11556 (N_11556,N_1338,N_3550);
or U11557 (N_11557,N_2538,N_2503);
or U11558 (N_11558,N_1377,N_3279);
nor U11559 (N_11559,N_6152,N_906);
nand U11560 (N_11560,N_3057,N_4146);
and U11561 (N_11561,N_5482,N_3959);
and U11562 (N_11562,N_6234,N_2299);
nor U11563 (N_11563,N_634,N_1110);
or U11564 (N_11564,N_3496,N_3651);
nor U11565 (N_11565,N_2855,N_1680);
and U11566 (N_11566,N_5541,N_4830);
xnor U11567 (N_11567,N_2282,N_2185);
xnor U11568 (N_11568,N_387,N_5350);
nor U11569 (N_11569,N_5840,N_4032);
xor U11570 (N_11570,N_1583,N_3151);
nor U11571 (N_11571,N_3258,N_1921);
nand U11572 (N_11572,N_3021,N_2840);
nand U11573 (N_11573,N_2774,N_2293);
xor U11574 (N_11574,N_637,N_5207);
or U11575 (N_11575,N_1242,N_3539);
nor U11576 (N_11576,N_4336,N_5708);
nand U11577 (N_11577,N_254,N_4297);
or U11578 (N_11578,N_2217,N_3325);
nor U11579 (N_11579,N_3182,N_217);
and U11580 (N_11580,N_1729,N_413);
or U11581 (N_11581,N_1347,N_4373);
nor U11582 (N_11582,N_2521,N_2179);
nor U11583 (N_11583,N_1892,N_1327);
xor U11584 (N_11584,N_3583,N_272);
xnor U11585 (N_11585,N_2630,N_3230);
nand U11586 (N_11586,N_37,N_1170);
and U11587 (N_11587,N_4901,N_6151);
xnor U11588 (N_11588,N_2824,N_966);
and U11589 (N_11589,N_5153,N_2502);
nor U11590 (N_11590,N_4121,N_3860);
and U11591 (N_11591,N_5208,N_5286);
xor U11592 (N_11592,N_1386,N_2509);
nor U11593 (N_11593,N_4733,N_709);
or U11594 (N_11594,N_3312,N_2778);
nand U11595 (N_11595,N_1649,N_13);
nor U11596 (N_11596,N_3859,N_351);
or U11597 (N_11597,N_2422,N_2309);
xor U11598 (N_11598,N_4315,N_4387);
and U11599 (N_11599,N_3091,N_5628);
nand U11600 (N_11600,N_5322,N_3472);
nand U11601 (N_11601,N_6211,N_5192);
and U11602 (N_11602,N_3168,N_5381);
xnor U11603 (N_11603,N_4158,N_1144);
or U11604 (N_11604,N_780,N_4586);
nand U11605 (N_11605,N_822,N_5097);
nor U11606 (N_11606,N_3990,N_3981);
or U11607 (N_11607,N_4179,N_4704);
and U11608 (N_11608,N_6169,N_2359);
and U11609 (N_11609,N_3890,N_2036);
or U11610 (N_11610,N_5495,N_5697);
nor U11611 (N_11611,N_97,N_6037);
or U11612 (N_11612,N_2971,N_1692);
xor U11613 (N_11613,N_5904,N_3604);
nor U11614 (N_11614,N_3001,N_106);
and U11615 (N_11615,N_2103,N_2802);
nor U11616 (N_11616,N_829,N_2685);
nand U11617 (N_11617,N_1205,N_3481);
xor U11618 (N_11618,N_2069,N_1089);
nor U11619 (N_11619,N_2069,N_3180);
nand U11620 (N_11620,N_1804,N_2186);
and U11621 (N_11621,N_2918,N_3824);
or U11622 (N_11622,N_585,N_3372);
or U11623 (N_11623,N_5504,N_551);
and U11624 (N_11624,N_757,N_4782);
xor U11625 (N_11625,N_3303,N_649);
nor U11626 (N_11626,N_663,N_3526);
nor U11627 (N_11627,N_3435,N_2065);
or U11628 (N_11628,N_4671,N_645);
nor U11629 (N_11629,N_5279,N_6045);
and U11630 (N_11630,N_5730,N_3098);
or U11631 (N_11631,N_402,N_130);
xor U11632 (N_11632,N_2522,N_5208);
nor U11633 (N_11633,N_6176,N_5830);
nand U11634 (N_11634,N_2153,N_1142);
xor U11635 (N_11635,N_3576,N_1718);
nand U11636 (N_11636,N_2154,N_3104);
xor U11637 (N_11637,N_4243,N_4789);
and U11638 (N_11638,N_1780,N_5699);
nor U11639 (N_11639,N_1297,N_4551);
xor U11640 (N_11640,N_4723,N_2246);
and U11641 (N_11641,N_2608,N_3939);
and U11642 (N_11642,N_1994,N_3788);
and U11643 (N_11643,N_1530,N_1798);
nand U11644 (N_11644,N_658,N_3179);
nor U11645 (N_11645,N_5065,N_4502);
and U11646 (N_11646,N_4178,N_4823);
xor U11647 (N_11647,N_5015,N_5345);
nand U11648 (N_11648,N_4460,N_3965);
or U11649 (N_11649,N_206,N_5075);
and U11650 (N_11650,N_667,N_2989);
nor U11651 (N_11651,N_6011,N_672);
nor U11652 (N_11652,N_3870,N_5695);
nor U11653 (N_11653,N_5673,N_5598);
nor U11654 (N_11654,N_4140,N_4307);
nor U11655 (N_11655,N_3045,N_3436);
xnor U11656 (N_11656,N_1322,N_3759);
nand U11657 (N_11657,N_2908,N_828);
nor U11658 (N_11658,N_128,N_1733);
and U11659 (N_11659,N_5406,N_6222);
nor U11660 (N_11660,N_4054,N_4541);
or U11661 (N_11661,N_4839,N_5525);
xor U11662 (N_11662,N_2035,N_3673);
and U11663 (N_11663,N_2405,N_979);
nand U11664 (N_11664,N_4106,N_517);
nor U11665 (N_11665,N_714,N_1008);
and U11666 (N_11666,N_214,N_6191);
xor U11667 (N_11667,N_5264,N_4446);
nand U11668 (N_11668,N_3591,N_1693);
nor U11669 (N_11669,N_5968,N_1151);
nand U11670 (N_11670,N_2185,N_2474);
nand U11671 (N_11671,N_1183,N_3116);
nor U11672 (N_11672,N_3417,N_933);
nor U11673 (N_11673,N_2442,N_6140);
and U11674 (N_11674,N_380,N_934);
or U11675 (N_11675,N_2679,N_543);
nand U11676 (N_11676,N_1264,N_5987);
nand U11677 (N_11677,N_425,N_946);
xor U11678 (N_11678,N_4198,N_4601);
nand U11679 (N_11679,N_5592,N_107);
and U11680 (N_11680,N_5936,N_1491);
nand U11681 (N_11681,N_1305,N_5565);
or U11682 (N_11682,N_2017,N_4455);
or U11683 (N_11683,N_3556,N_5239);
xnor U11684 (N_11684,N_3120,N_2560);
and U11685 (N_11685,N_5611,N_5476);
nand U11686 (N_11686,N_2585,N_2814);
or U11687 (N_11687,N_6179,N_2608);
nand U11688 (N_11688,N_5181,N_3118);
nor U11689 (N_11689,N_1887,N_6030);
and U11690 (N_11690,N_774,N_1786);
xor U11691 (N_11691,N_1741,N_5092);
nor U11692 (N_11692,N_5721,N_1505);
nand U11693 (N_11693,N_2662,N_2626);
nor U11694 (N_11694,N_1767,N_4904);
and U11695 (N_11695,N_267,N_6163);
nor U11696 (N_11696,N_3968,N_3407);
nor U11697 (N_11697,N_2948,N_5003);
nand U11698 (N_11698,N_5744,N_5010);
or U11699 (N_11699,N_2039,N_1978);
nor U11700 (N_11700,N_5167,N_3352);
xnor U11701 (N_11701,N_2204,N_873);
nor U11702 (N_11702,N_6214,N_3011);
nand U11703 (N_11703,N_2977,N_3600);
xor U11704 (N_11704,N_4768,N_4333);
and U11705 (N_11705,N_5016,N_4015);
nor U11706 (N_11706,N_4307,N_5245);
nor U11707 (N_11707,N_925,N_1925);
nand U11708 (N_11708,N_1099,N_4921);
or U11709 (N_11709,N_3048,N_3649);
nor U11710 (N_11710,N_547,N_2282);
nor U11711 (N_11711,N_3352,N_5742);
or U11712 (N_11712,N_2676,N_287);
and U11713 (N_11713,N_3580,N_4966);
nor U11714 (N_11714,N_1977,N_5149);
and U11715 (N_11715,N_2681,N_4244);
nor U11716 (N_11716,N_3028,N_2530);
nand U11717 (N_11717,N_3994,N_5304);
or U11718 (N_11718,N_1032,N_4846);
xnor U11719 (N_11719,N_4858,N_5609);
and U11720 (N_11720,N_3708,N_5868);
nor U11721 (N_11721,N_4212,N_4575);
nand U11722 (N_11722,N_514,N_296);
and U11723 (N_11723,N_2608,N_2830);
or U11724 (N_11724,N_4832,N_623);
nand U11725 (N_11725,N_4698,N_2982);
nand U11726 (N_11726,N_5603,N_2361);
xor U11727 (N_11727,N_3107,N_491);
nand U11728 (N_11728,N_5211,N_3540);
xor U11729 (N_11729,N_37,N_5738);
or U11730 (N_11730,N_4923,N_590);
or U11731 (N_11731,N_4763,N_3562);
xnor U11732 (N_11732,N_214,N_2596);
xnor U11733 (N_11733,N_2310,N_4070);
nor U11734 (N_11734,N_2940,N_6097);
and U11735 (N_11735,N_1970,N_4729);
xor U11736 (N_11736,N_4417,N_3029);
or U11737 (N_11737,N_2561,N_3147);
or U11738 (N_11738,N_4910,N_4476);
and U11739 (N_11739,N_1220,N_11);
or U11740 (N_11740,N_2428,N_469);
and U11741 (N_11741,N_5640,N_637);
or U11742 (N_11742,N_326,N_3204);
xnor U11743 (N_11743,N_1883,N_4083);
xor U11744 (N_11744,N_455,N_4912);
xor U11745 (N_11745,N_4868,N_5557);
nand U11746 (N_11746,N_4209,N_1404);
nor U11747 (N_11747,N_2346,N_4605);
and U11748 (N_11748,N_2470,N_5609);
nand U11749 (N_11749,N_4751,N_2839);
xor U11750 (N_11750,N_4818,N_3987);
nand U11751 (N_11751,N_2289,N_4581);
xnor U11752 (N_11752,N_5917,N_5780);
nand U11753 (N_11753,N_6097,N_3214);
nand U11754 (N_11754,N_1265,N_2729);
xor U11755 (N_11755,N_5187,N_1792);
xnor U11756 (N_11756,N_5747,N_3697);
nor U11757 (N_11757,N_5549,N_6229);
and U11758 (N_11758,N_6219,N_2763);
and U11759 (N_11759,N_696,N_5964);
xor U11760 (N_11760,N_3986,N_940);
nand U11761 (N_11761,N_5399,N_2292);
and U11762 (N_11762,N_1425,N_1844);
or U11763 (N_11763,N_3098,N_4323);
and U11764 (N_11764,N_2439,N_1217);
and U11765 (N_11765,N_4166,N_2692);
and U11766 (N_11766,N_682,N_3772);
xor U11767 (N_11767,N_4646,N_4510);
and U11768 (N_11768,N_1349,N_1265);
nand U11769 (N_11769,N_1158,N_523);
xor U11770 (N_11770,N_5037,N_4306);
or U11771 (N_11771,N_3715,N_247);
xor U11772 (N_11772,N_2361,N_2678);
and U11773 (N_11773,N_2722,N_4869);
nand U11774 (N_11774,N_3491,N_3494);
and U11775 (N_11775,N_1106,N_4544);
xnor U11776 (N_11776,N_2876,N_2059);
or U11777 (N_11777,N_2515,N_1639);
nand U11778 (N_11778,N_210,N_2186);
nand U11779 (N_11779,N_1464,N_3507);
and U11780 (N_11780,N_4955,N_5253);
and U11781 (N_11781,N_3581,N_4038);
or U11782 (N_11782,N_2504,N_1951);
nor U11783 (N_11783,N_1649,N_155);
or U11784 (N_11784,N_4398,N_4776);
or U11785 (N_11785,N_1544,N_4854);
xnor U11786 (N_11786,N_4227,N_4985);
and U11787 (N_11787,N_4522,N_4108);
or U11788 (N_11788,N_3500,N_3987);
or U11789 (N_11789,N_1072,N_203);
nand U11790 (N_11790,N_2354,N_5522);
nor U11791 (N_11791,N_5247,N_4441);
nor U11792 (N_11792,N_3610,N_4173);
nand U11793 (N_11793,N_1425,N_461);
and U11794 (N_11794,N_5699,N_1147);
or U11795 (N_11795,N_2812,N_221);
and U11796 (N_11796,N_5459,N_1610);
or U11797 (N_11797,N_2703,N_5034);
or U11798 (N_11798,N_1406,N_901);
or U11799 (N_11799,N_1141,N_846);
xor U11800 (N_11800,N_3313,N_3757);
and U11801 (N_11801,N_2194,N_3816);
nand U11802 (N_11802,N_969,N_5982);
nand U11803 (N_11803,N_3114,N_6186);
nor U11804 (N_11804,N_1796,N_6033);
and U11805 (N_11805,N_1728,N_896);
or U11806 (N_11806,N_2566,N_3158);
nand U11807 (N_11807,N_4426,N_3617);
nand U11808 (N_11808,N_1111,N_1092);
nand U11809 (N_11809,N_3317,N_5794);
or U11810 (N_11810,N_1856,N_5592);
and U11811 (N_11811,N_3992,N_3768);
xor U11812 (N_11812,N_4259,N_1766);
nor U11813 (N_11813,N_3281,N_1826);
nor U11814 (N_11814,N_4053,N_978);
nor U11815 (N_11815,N_1363,N_2397);
nor U11816 (N_11816,N_2147,N_4324);
or U11817 (N_11817,N_821,N_1202);
xor U11818 (N_11818,N_1746,N_4479);
nand U11819 (N_11819,N_3656,N_180);
nor U11820 (N_11820,N_3093,N_2914);
nand U11821 (N_11821,N_3106,N_174);
nand U11822 (N_11822,N_5622,N_4704);
nand U11823 (N_11823,N_5979,N_4273);
nor U11824 (N_11824,N_3326,N_5431);
nand U11825 (N_11825,N_1099,N_397);
xnor U11826 (N_11826,N_6105,N_3095);
or U11827 (N_11827,N_1976,N_5061);
nand U11828 (N_11828,N_4432,N_3297);
xnor U11829 (N_11829,N_1960,N_4268);
nand U11830 (N_11830,N_5173,N_4801);
or U11831 (N_11831,N_5388,N_2899);
nor U11832 (N_11832,N_3538,N_6202);
nand U11833 (N_11833,N_1781,N_1278);
xnor U11834 (N_11834,N_1779,N_414);
xnor U11835 (N_11835,N_2937,N_4389);
and U11836 (N_11836,N_5702,N_1899);
nand U11837 (N_11837,N_6214,N_840);
or U11838 (N_11838,N_3729,N_605);
nand U11839 (N_11839,N_3089,N_4617);
or U11840 (N_11840,N_1081,N_3524);
nor U11841 (N_11841,N_877,N_1);
nor U11842 (N_11842,N_5035,N_5656);
nor U11843 (N_11843,N_4640,N_4892);
nand U11844 (N_11844,N_5272,N_299);
nand U11845 (N_11845,N_3779,N_2851);
and U11846 (N_11846,N_3011,N_4036);
nand U11847 (N_11847,N_2451,N_217);
nand U11848 (N_11848,N_4554,N_5064);
and U11849 (N_11849,N_215,N_3547);
xnor U11850 (N_11850,N_4100,N_4256);
nand U11851 (N_11851,N_4205,N_5634);
or U11852 (N_11852,N_619,N_173);
xor U11853 (N_11853,N_1716,N_4619);
or U11854 (N_11854,N_4086,N_5461);
nand U11855 (N_11855,N_2741,N_5585);
or U11856 (N_11856,N_5874,N_1076);
xnor U11857 (N_11857,N_2592,N_668);
and U11858 (N_11858,N_2648,N_5152);
xnor U11859 (N_11859,N_1090,N_3215);
or U11860 (N_11860,N_3062,N_3232);
and U11861 (N_11861,N_5936,N_5050);
and U11862 (N_11862,N_3066,N_4476);
xnor U11863 (N_11863,N_1601,N_6197);
nand U11864 (N_11864,N_1106,N_5018);
nor U11865 (N_11865,N_3627,N_4496);
or U11866 (N_11866,N_5535,N_1701);
and U11867 (N_11867,N_2979,N_2109);
or U11868 (N_11868,N_5593,N_619);
nand U11869 (N_11869,N_703,N_5013);
and U11870 (N_11870,N_5651,N_64);
and U11871 (N_11871,N_5846,N_1876);
or U11872 (N_11872,N_1387,N_1531);
and U11873 (N_11873,N_3846,N_4639);
nand U11874 (N_11874,N_5813,N_3658);
nand U11875 (N_11875,N_4071,N_3800);
nor U11876 (N_11876,N_5984,N_3041);
nor U11877 (N_11877,N_2198,N_1180);
xnor U11878 (N_11878,N_5937,N_626);
or U11879 (N_11879,N_1801,N_971);
and U11880 (N_11880,N_5153,N_584);
or U11881 (N_11881,N_6150,N_5837);
or U11882 (N_11882,N_1013,N_4038);
nor U11883 (N_11883,N_4274,N_254);
xnor U11884 (N_11884,N_4034,N_3441);
or U11885 (N_11885,N_5642,N_595);
xor U11886 (N_11886,N_1673,N_5516);
or U11887 (N_11887,N_2803,N_2496);
nand U11888 (N_11888,N_393,N_2696);
nand U11889 (N_11889,N_883,N_1077);
and U11890 (N_11890,N_4166,N_5038);
nand U11891 (N_11891,N_889,N_2900);
or U11892 (N_11892,N_978,N_5716);
nor U11893 (N_11893,N_876,N_2782);
and U11894 (N_11894,N_5503,N_3192);
nor U11895 (N_11895,N_2834,N_5436);
and U11896 (N_11896,N_5696,N_256);
xor U11897 (N_11897,N_1908,N_3035);
and U11898 (N_11898,N_3818,N_1844);
xnor U11899 (N_11899,N_6006,N_6193);
or U11900 (N_11900,N_3265,N_3380);
nand U11901 (N_11901,N_2906,N_2756);
xnor U11902 (N_11902,N_3181,N_3879);
and U11903 (N_11903,N_488,N_2344);
nor U11904 (N_11904,N_894,N_6060);
nand U11905 (N_11905,N_1875,N_4677);
nor U11906 (N_11906,N_2885,N_3186);
xnor U11907 (N_11907,N_867,N_3834);
and U11908 (N_11908,N_2989,N_2485);
xnor U11909 (N_11909,N_3135,N_1371);
xnor U11910 (N_11910,N_2153,N_272);
nand U11911 (N_11911,N_1481,N_1857);
xor U11912 (N_11912,N_4852,N_3565);
xor U11913 (N_11913,N_1721,N_2939);
nand U11914 (N_11914,N_4335,N_724);
or U11915 (N_11915,N_990,N_918);
and U11916 (N_11916,N_6195,N_1785);
and U11917 (N_11917,N_4269,N_4951);
and U11918 (N_11918,N_5471,N_422);
xor U11919 (N_11919,N_4747,N_3789);
or U11920 (N_11920,N_2106,N_2966);
nor U11921 (N_11921,N_5981,N_4888);
nor U11922 (N_11922,N_1605,N_556);
nor U11923 (N_11923,N_5707,N_267);
xor U11924 (N_11924,N_5245,N_5251);
xor U11925 (N_11925,N_1855,N_5817);
nor U11926 (N_11926,N_95,N_5452);
xnor U11927 (N_11927,N_2966,N_4778);
nand U11928 (N_11928,N_2831,N_3322);
or U11929 (N_11929,N_3927,N_3191);
xnor U11930 (N_11930,N_4669,N_3995);
or U11931 (N_11931,N_3053,N_5179);
nand U11932 (N_11932,N_490,N_2022);
xor U11933 (N_11933,N_3164,N_12);
xnor U11934 (N_11934,N_3747,N_1985);
nor U11935 (N_11935,N_528,N_1815);
or U11936 (N_11936,N_3313,N_5234);
or U11937 (N_11937,N_5838,N_903);
and U11938 (N_11938,N_2611,N_4246);
and U11939 (N_11939,N_5146,N_518);
and U11940 (N_11940,N_435,N_4457);
nand U11941 (N_11941,N_5441,N_5701);
and U11942 (N_11942,N_3008,N_6173);
nand U11943 (N_11943,N_4601,N_5174);
nor U11944 (N_11944,N_5782,N_5807);
xor U11945 (N_11945,N_4818,N_811);
and U11946 (N_11946,N_3361,N_181);
nand U11947 (N_11947,N_4266,N_638);
or U11948 (N_11948,N_1325,N_5427);
and U11949 (N_11949,N_2771,N_4804);
xor U11950 (N_11950,N_3565,N_581);
or U11951 (N_11951,N_3388,N_5904);
nand U11952 (N_11952,N_3240,N_6039);
nor U11953 (N_11953,N_858,N_6199);
or U11954 (N_11954,N_3372,N_6069);
nor U11955 (N_11955,N_1801,N_5054);
or U11956 (N_11956,N_948,N_1288);
xnor U11957 (N_11957,N_3398,N_3042);
and U11958 (N_11958,N_3132,N_428);
nand U11959 (N_11959,N_1194,N_3243);
and U11960 (N_11960,N_4189,N_4986);
and U11961 (N_11961,N_3945,N_2791);
nor U11962 (N_11962,N_2517,N_4085);
or U11963 (N_11963,N_1152,N_5226);
or U11964 (N_11964,N_3403,N_991);
xnor U11965 (N_11965,N_1320,N_2549);
nor U11966 (N_11966,N_3533,N_2213);
or U11967 (N_11967,N_2817,N_3082);
nand U11968 (N_11968,N_5751,N_5398);
xnor U11969 (N_11969,N_3550,N_1729);
and U11970 (N_11970,N_4716,N_1644);
nor U11971 (N_11971,N_1165,N_4282);
or U11972 (N_11972,N_1252,N_6041);
nand U11973 (N_11973,N_3847,N_5887);
and U11974 (N_11974,N_1009,N_4611);
nor U11975 (N_11975,N_2607,N_4766);
or U11976 (N_11976,N_4634,N_4120);
and U11977 (N_11977,N_2711,N_3610);
nand U11978 (N_11978,N_2166,N_5662);
xor U11979 (N_11979,N_1895,N_2886);
nand U11980 (N_11980,N_4144,N_470);
nand U11981 (N_11981,N_2216,N_2653);
and U11982 (N_11982,N_5168,N_3142);
nor U11983 (N_11983,N_2473,N_570);
and U11984 (N_11984,N_4849,N_72);
or U11985 (N_11985,N_2498,N_2533);
or U11986 (N_11986,N_3067,N_1854);
nor U11987 (N_11987,N_2189,N_4261);
nor U11988 (N_11988,N_2857,N_5158);
and U11989 (N_11989,N_5247,N_1521);
nor U11990 (N_11990,N_3679,N_2605);
and U11991 (N_11991,N_573,N_4043);
nand U11992 (N_11992,N_3408,N_301);
or U11993 (N_11993,N_2189,N_2086);
nor U11994 (N_11994,N_3582,N_5976);
or U11995 (N_11995,N_2568,N_4133);
nor U11996 (N_11996,N_4778,N_1738);
xor U11997 (N_11997,N_2490,N_5682);
xor U11998 (N_11998,N_4305,N_2616);
or U11999 (N_11999,N_1814,N_1861);
xnor U12000 (N_12000,N_4699,N_6122);
nand U12001 (N_12001,N_5820,N_4455);
nor U12002 (N_12002,N_5811,N_1624);
xnor U12003 (N_12003,N_1371,N_309);
or U12004 (N_12004,N_5971,N_5193);
or U12005 (N_12005,N_1646,N_1678);
nand U12006 (N_12006,N_5104,N_4822);
or U12007 (N_12007,N_4825,N_4144);
xor U12008 (N_12008,N_1783,N_836);
and U12009 (N_12009,N_370,N_3882);
and U12010 (N_12010,N_3630,N_3406);
or U12011 (N_12011,N_3389,N_4603);
xnor U12012 (N_12012,N_3532,N_2516);
xor U12013 (N_12013,N_2960,N_695);
xor U12014 (N_12014,N_557,N_6137);
and U12015 (N_12015,N_120,N_6167);
or U12016 (N_12016,N_2396,N_1566);
nand U12017 (N_12017,N_3941,N_5703);
nand U12018 (N_12018,N_2476,N_2489);
or U12019 (N_12019,N_3138,N_6072);
xnor U12020 (N_12020,N_5449,N_2289);
and U12021 (N_12021,N_3420,N_1793);
xor U12022 (N_12022,N_5689,N_1015);
nand U12023 (N_12023,N_1727,N_5332);
and U12024 (N_12024,N_3348,N_1132);
or U12025 (N_12025,N_2862,N_4903);
xnor U12026 (N_12026,N_3549,N_32);
and U12027 (N_12027,N_1995,N_4527);
and U12028 (N_12028,N_1109,N_5939);
nand U12029 (N_12029,N_5947,N_4244);
or U12030 (N_12030,N_3081,N_2972);
nor U12031 (N_12031,N_4377,N_2776);
xnor U12032 (N_12032,N_3865,N_3486);
or U12033 (N_12033,N_1517,N_1582);
nand U12034 (N_12034,N_2584,N_748);
xor U12035 (N_12035,N_1044,N_570);
nor U12036 (N_12036,N_4013,N_3824);
nor U12037 (N_12037,N_6213,N_925);
nand U12038 (N_12038,N_4641,N_275);
nand U12039 (N_12039,N_5045,N_2801);
and U12040 (N_12040,N_3826,N_1622);
and U12041 (N_12041,N_5035,N_3194);
and U12042 (N_12042,N_3856,N_4288);
or U12043 (N_12043,N_3845,N_969);
xor U12044 (N_12044,N_4730,N_4710);
or U12045 (N_12045,N_3286,N_5331);
or U12046 (N_12046,N_6043,N_1140);
or U12047 (N_12047,N_5770,N_1740);
or U12048 (N_12048,N_2226,N_2459);
nor U12049 (N_12049,N_4828,N_4714);
nand U12050 (N_12050,N_2299,N_1139);
nor U12051 (N_12051,N_230,N_1744);
or U12052 (N_12052,N_3767,N_5808);
nor U12053 (N_12053,N_3333,N_3285);
and U12054 (N_12054,N_1932,N_4777);
nor U12055 (N_12055,N_2100,N_5604);
xnor U12056 (N_12056,N_3983,N_4906);
xnor U12057 (N_12057,N_4322,N_5919);
nor U12058 (N_12058,N_2699,N_3380);
nand U12059 (N_12059,N_2912,N_5699);
nor U12060 (N_12060,N_6247,N_2088);
nand U12061 (N_12061,N_5761,N_4634);
nand U12062 (N_12062,N_717,N_397);
xnor U12063 (N_12063,N_6011,N_2511);
and U12064 (N_12064,N_52,N_580);
and U12065 (N_12065,N_3497,N_5149);
and U12066 (N_12066,N_599,N_5231);
nor U12067 (N_12067,N_6095,N_44);
or U12068 (N_12068,N_2603,N_5893);
and U12069 (N_12069,N_4804,N_604);
or U12070 (N_12070,N_2579,N_3498);
xor U12071 (N_12071,N_5098,N_981);
or U12072 (N_12072,N_5434,N_4871);
xor U12073 (N_12073,N_2241,N_1637);
xor U12074 (N_12074,N_5729,N_5715);
and U12075 (N_12075,N_922,N_1330);
nor U12076 (N_12076,N_86,N_2628);
xnor U12077 (N_12077,N_1921,N_2501);
nand U12078 (N_12078,N_3328,N_1543);
or U12079 (N_12079,N_4093,N_2912);
or U12080 (N_12080,N_4121,N_3764);
nand U12081 (N_12081,N_4282,N_3526);
nand U12082 (N_12082,N_1300,N_4678);
nor U12083 (N_12083,N_1019,N_4805);
nor U12084 (N_12084,N_4757,N_2567);
and U12085 (N_12085,N_2044,N_4181);
xor U12086 (N_12086,N_2298,N_1967);
nor U12087 (N_12087,N_4547,N_435);
xnor U12088 (N_12088,N_3664,N_4537);
or U12089 (N_12089,N_527,N_5770);
or U12090 (N_12090,N_2717,N_2808);
nand U12091 (N_12091,N_2600,N_4833);
or U12092 (N_12092,N_5662,N_5018);
xnor U12093 (N_12093,N_3706,N_3613);
xor U12094 (N_12094,N_25,N_2158);
nand U12095 (N_12095,N_2736,N_4749);
nand U12096 (N_12096,N_3416,N_1815);
nor U12097 (N_12097,N_1898,N_4742);
and U12098 (N_12098,N_4963,N_2330);
or U12099 (N_12099,N_2526,N_188);
xnor U12100 (N_12100,N_3271,N_1325);
xor U12101 (N_12101,N_38,N_2813);
xnor U12102 (N_12102,N_629,N_282);
or U12103 (N_12103,N_3932,N_1516);
xnor U12104 (N_12104,N_4151,N_4524);
or U12105 (N_12105,N_5414,N_2840);
and U12106 (N_12106,N_2954,N_4225);
xnor U12107 (N_12107,N_3097,N_6249);
nand U12108 (N_12108,N_2402,N_2588);
and U12109 (N_12109,N_2264,N_4921);
nor U12110 (N_12110,N_2891,N_764);
and U12111 (N_12111,N_3720,N_1550);
or U12112 (N_12112,N_3105,N_5520);
nand U12113 (N_12113,N_587,N_1110);
xnor U12114 (N_12114,N_4017,N_5494);
nor U12115 (N_12115,N_1098,N_5498);
nor U12116 (N_12116,N_2731,N_623);
xnor U12117 (N_12117,N_1411,N_4893);
nand U12118 (N_12118,N_1044,N_5418);
or U12119 (N_12119,N_1897,N_2842);
and U12120 (N_12120,N_4092,N_3108);
and U12121 (N_12121,N_4559,N_728);
xnor U12122 (N_12122,N_5967,N_3347);
and U12123 (N_12123,N_2376,N_1356);
xnor U12124 (N_12124,N_3575,N_6157);
nand U12125 (N_12125,N_379,N_168);
or U12126 (N_12126,N_690,N_4431);
nand U12127 (N_12127,N_2289,N_3012);
nand U12128 (N_12128,N_6010,N_2314);
xor U12129 (N_12129,N_2644,N_837);
and U12130 (N_12130,N_2365,N_4159);
or U12131 (N_12131,N_5928,N_4916);
and U12132 (N_12132,N_4806,N_1092);
or U12133 (N_12133,N_824,N_154);
and U12134 (N_12134,N_4248,N_5332);
nand U12135 (N_12135,N_862,N_5592);
nor U12136 (N_12136,N_4292,N_1588);
xnor U12137 (N_12137,N_3587,N_2315);
xnor U12138 (N_12138,N_5862,N_156);
xor U12139 (N_12139,N_4325,N_2397);
xnor U12140 (N_12140,N_5280,N_1021);
xor U12141 (N_12141,N_4768,N_203);
and U12142 (N_12142,N_1897,N_4251);
and U12143 (N_12143,N_693,N_2327);
and U12144 (N_12144,N_4295,N_3693);
nor U12145 (N_12145,N_3862,N_3680);
nor U12146 (N_12146,N_5055,N_5791);
and U12147 (N_12147,N_5946,N_2717);
xnor U12148 (N_12148,N_3285,N_2315);
and U12149 (N_12149,N_2301,N_5684);
nor U12150 (N_12150,N_5160,N_1927);
or U12151 (N_12151,N_2357,N_3834);
and U12152 (N_12152,N_3479,N_2221);
nor U12153 (N_12153,N_4003,N_1731);
xnor U12154 (N_12154,N_2808,N_4704);
nor U12155 (N_12155,N_302,N_913);
nor U12156 (N_12156,N_1142,N_5438);
nor U12157 (N_12157,N_5234,N_5996);
nand U12158 (N_12158,N_299,N_6012);
xnor U12159 (N_12159,N_6158,N_3843);
xor U12160 (N_12160,N_1199,N_2315);
and U12161 (N_12161,N_920,N_742);
or U12162 (N_12162,N_2180,N_6228);
and U12163 (N_12163,N_997,N_3710);
and U12164 (N_12164,N_3484,N_2901);
nor U12165 (N_12165,N_867,N_3364);
or U12166 (N_12166,N_1095,N_1999);
or U12167 (N_12167,N_4634,N_4816);
and U12168 (N_12168,N_3337,N_1302);
and U12169 (N_12169,N_153,N_402);
and U12170 (N_12170,N_1172,N_3988);
nand U12171 (N_12171,N_5060,N_483);
xnor U12172 (N_12172,N_1233,N_4906);
nor U12173 (N_12173,N_4891,N_955);
xor U12174 (N_12174,N_4390,N_1937);
nand U12175 (N_12175,N_5762,N_2018);
nand U12176 (N_12176,N_3125,N_592);
nand U12177 (N_12177,N_1428,N_1756);
or U12178 (N_12178,N_2265,N_1555);
nand U12179 (N_12179,N_74,N_3026);
nand U12180 (N_12180,N_5203,N_840);
xnor U12181 (N_12181,N_4148,N_2747);
or U12182 (N_12182,N_3681,N_201);
and U12183 (N_12183,N_1639,N_1322);
xor U12184 (N_12184,N_4341,N_4123);
nand U12185 (N_12185,N_5398,N_5430);
xor U12186 (N_12186,N_4188,N_6033);
or U12187 (N_12187,N_4212,N_2173);
or U12188 (N_12188,N_5650,N_3296);
nor U12189 (N_12189,N_1474,N_5405);
and U12190 (N_12190,N_4820,N_2079);
nor U12191 (N_12191,N_3669,N_5791);
nand U12192 (N_12192,N_13,N_60);
xnor U12193 (N_12193,N_5104,N_357);
nand U12194 (N_12194,N_1788,N_3699);
or U12195 (N_12195,N_4610,N_2332);
nor U12196 (N_12196,N_3667,N_5241);
xnor U12197 (N_12197,N_1499,N_1794);
xnor U12198 (N_12198,N_5124,N_43);
nor U12199 (N_12199,N_978,N_142);
xnor U12200 (N_12200,N_1284,N_4296);
and U12201 (N_12201,N_4709,N_6227);
nand U12202 (N_12202,N_116,N_1689);
nor U12203 (N_12203,N_4082,N_5848);
and U12204 (N_12204,N_3885,N_915);
nand U12205 (N_12205,N_279,N_3331);
and U12206 (N_12206,N_1829,N_3513);
nor U12207 (N_12207,N_2775,N_4775);
or U12208 (N_12208,N_2859,N_1174);
nand U12209 (N_12209,N_4890,N_1979);
nand U12210 (N_12210,N_6246,N_5612);
nor U12211 (N_12211,N_3674,N_3363);
or U12212 (N_12212,N_3946,N_2524);
xor U12213 (N_12213,N_2760,N_122);
and U12214 (N_12214,N_6121,N_1798);
or U12215 (N_12215,N_1273,N_4803);
nor U12216 (N_12216,N_2302,N_5451);
nand U12217 (N_12217,N_3429,N_1152);
or U12218 (N_12218,N_5110,N_3193);
xnor U12219 (N_12219,N_3667,N_4733);
nand U12220 (N_12220,N_3594,N_718);
nand U12221 (N_12221,N_3028,N_4524);
xnor U12222 (N_12222,N_4978,N_4682);
and U12223 (N_12223,N_415,N_3093);
or U12224 (N_12224,N_1269,N_1007);
nand U12225 (N_12225,N_5282,N_3969);
or U12226 (N_12226,N_715,N_4701);
nor U12227 (N_12227,N_392,N_5549);
xnor U12228 (N_12228,N_971,N_1217);
nand U12229 (N_12229,N_2746,N_1064);
nand U12230 (N_12230,N_1075,N_2277);
nor U12231 (N_12231,N_910,N_1963);
or U12232 (N_12232,N_324,N_1958);
nor U12233 (N_12233,N_4601,N_5426);
nor U12234 (N_12234,N_1200,N_419);
nand U12235 (N_12235,N_3662,N_3021);
or U12236 (N_12236,N_4997,N_4399);
xnor U12237 (N_12237,N_75,N_1429);
and U12238 (N_12238,N_6016,N_6224);
xnor U12239 (N_12239,N_255,N_3230);
nor U12240 (N_12240,N_2881,N_5576);
and U12241 (N_12241,N_1758,N_284);
and U12242 (N_12242,N_3570,N_4173);
nor U12243 (N_12243,N_3011,N_275);
and U12244 (N_12244,N_2673,N_2012);
xnor U12245 (N_12245,N_3891,N_5346);
nor U12246 (N_12246,N_2004,N_1033);
nand U12247 (N_12247,N_2284,N_4836);
and U12248 (N_12248,N_6132,N_5661);
nand U12249 (N_12249,N_3832,N_2739);
xor U12250 (N_12250,N_640,N_4095);
and U12251 (N_12251,N_4376,N_4946);
and U12252 (N_12252,N_3825,N_4005);
nand U12253 (N_12253,N_2112,N_4792);
nor U12254 (N_12254,N_5096,N_3956);
xor U12255 (N_12255,N_4270,N_4913);
xor U12256 (N_12256,N_904,N_608);
or U12257 (N_12257,N_3532,N_1802);
or U12258 (N_12258,N_2629,N_1226);
nand U12259 (N_12259,N_4868,N_5279);
and U12260 (N_12260,N_2479,N_3862);
xnor U12261 (N_12261,N_3587,N_3542);
nor U12262 (N_12262,N_3099,N_1341);
xor U12263 (N_12263,N_1345,N_5132);
and U12264 (N_12264,N_5604,N_4396);
and U12265 (N_12265,N_5865,N_4983);
or U12266 (N_12266,N_4495,N_2639);
nand U12267 (N_12267,N_4831,N_127);
nand U12268 (N_12268,N_5170,N_4679);
xnor U12269 (N_12269,N_4285,N_3333);
or U12270 (N_12270,N_5935,N_2016);
or U12271 (N_12271,N_3595,N_3312);
nand U12272 (N_12272,N_2681,N_629);
xor U12273 (N_12273,N_6193,N_1071);
and U12274 (N_12274,N_2609,N_2341);
or U12275 (N_12275,N_1391,N_6075);
and U12276 (N_12276,N_6003,N_2775);
nand U12277 (N_12277,N_5893,N_5314);
or U12278 (N_12278,N_1542,N_1545);
nand U12279 (N_12279,N_1419,N_5963);
xnor U12280 (N_12280,N_812,N_5237);
xor U12281 (N_12281,N_3589,N_4552);
nor U12282 (N_12282,N_4977,N_5955);
nand U12283 (N_12283,N_5939,N_333);
and U12284 (N_12284,N_2636,N_1163);
and U12285 (N_12285,N_276,N_2514);
and U12286 (N_12286,N_1219,N_3222);
nand U12287 (N_12287,N_1978,N_637);
or U12288 (N_12288,N_2173,N_24);
xnor U12289 (N_12289,N_5598,N_2481);
or U12290 (N_12290,N_2869,N_5455);
or U12291 (N_12291,N_2724,N_1039);
or U12292 (N_12292,N_2143,N_4004);
nand U12293 (N_12293,N_5221,N_3531);
and U12294 (N_12294,N_2913,N_3955);
or U12295 (N_12295,N_1228,N_3416);
and U12296 (N_12296,N_3744,N_5488);
nor U12297 (N_12297,N_5864,N_580);
nor U12298 (N_12298,N_2692,N_4246);
xnor U12299 (N_12299,N_2553,N_5322);
nor U12300 (N_12300,N_3143,N_3485);
nand U12301 (N_12301,N_624,N_3775);
or U12302 (N_12302,N_3267,N_960);
nor U12303 (N_12303,N_294,N_5501);
or U12304 (N_12304,N_5634,N_1755);
nor U12305 (N_12305,N_707,N_2430);
nor U12306 (N_12306,N_5472,N_5391);
or U12307 (N_12307,N_3447,N_1149);
nor U12308 (N_12308,N_5404,N_3532);
and U12309 (N_12309,N_3543,N_471);
nand U12310 (N_12310,N_2160,N_5847);
or U12311 (N_12311,N_3984,N_2088);
and U12312 (N_12312,N_6247,N_2939);
nand U12313 (N_12313,N_5203,N_5868);
xnor U12314 (N_12314,N_3475,N_3062);
and U12315 (N_12315,N_4407,N_2761);
nand U12316 (N_12316,N_609,N_4879);
and U12317 (N_12317,N_3125,N_1887);
and U12318 (N_12318,N_3587,N_5490);
nand U12319 (N_12319,N_2908,N_3757);
nor U12320 (N_12320,N_1218,N_3629);
nand U12321 (N_12321,N_3173,N_2692);
nor U12322 (N_12322,N_3993,N_251);
or U12323 (N_12323,N_3093,N_3187);
nor U12324 (N_12324,N_87,N_711);
and U12325 (N_12325,N_1228,N_940);
or U12326 (N_12326,N_4427,N_3438);
or U12327 (N_12327,N_4295,N_5069);
xor U12328 (N_12328,N_2933,N_5870);
nor U12329 (N_12329,N_2606,N_2029);
xnor U12330 (N_12330,N_4112,N_1894);
or U12331 (N_12331,N_385,N_2762);
nor U12332 (N_12332,N_4080,N_257);
or U12333 (N_12333,N_4419,N_6093);
and U12334 (N_12334,N_2796,N_766);
xor U12335 (N_12335,N_1354,N_4067);
and U12336 (N_12336,N_4413,N_1911);
nand U12337 (N_12337,N_3487,N_1174);
or U12338 (N_12338,N_6223,N_2675);
xnor U12339 (N_12339,N_3571,N_1426);
xnor U12340 (N_12340,N_5264,N_2647);
nand U12341 (N_12341,N_316,N_5329);
xnor U12342 (N_12342,N_5888,N_4429);
xor U12343 (N_12343,N_4814,N_2062);
and U12344 (N_12344,N_2213,N_4042);
or U12345 (N_12345,N_1979,N_5536);
and U12346 (N_12346,N_4163,N_1603);
nor U12347 (N_12347,N_4699,N_4335);
and U12348 (N_12348,N_2978,N_1843);
or U12349 (N_12349,N_646,N_4073);
nand U12350 (N_12350,N_1592,N_3285);
xnor U12351 (N_12351,N_2541,N_888);
nor U12352 (N_12352,N_2239,N_4638);
xnor U12353 (N_12353,N_2244,N_4143);
nand U12354 (N_12354,N_2942,N_5104);
or U12355 (N_12355,N_3153,N_116);
nor U12356 (N_12356,N_6243,N_431);
nand U12357 (N_12357,N_3750,N_1129);
or U12358 (N_12358,N_1309,N_1930);
or U12359 (N_12359,N_1857,N_1967);
nor U12360 (N_12360,N_3939,N_5897);
nor U12361 (N_12361,N_4139,N_85);
nor U12362 (N_12362,N_1932,N_3430);
xnor U12363 (N_12363,N_4793,N_6037);
xor U12364 (N_12364,N_3465,N_428);
or U12365 (N_12365,N_1728,N_3357);
nand U12366 (N_12366,N_1301,N_3656);
nand U12367 (N_12367,N_1662,N_5473);
or U12368 (N_12368,N_2666,N_2858);
xor U12369 (N_12369,N_3868,N_2794);
nor U12370 (N_12370,N_1133,N_5994);
or U12371 (N_12371,N_4560,N_3295);
xor U12372 (N_12372,N_5402,N_1153);
xnor U12373 (N_12373,N_3780,N_4595);
xnor U12374 (N_12374,N_5241,N_5037);
or U12375 (N_12375,N_725,N_5764);
nand U12376 (N_12376,N_4650,N_4590);
nand U12377 (N_12377,N_1756,N_1271);
nand U12378 (N_12378,N_2354,N_5423);
and U12379 (N_12379,N_3136,N_4930);
or U12380 (N_12380,N_4218,N_1885);
xnor U12381 (N_12381,N_3628,N_3606);
nand U12382 (N_12382,N_1869,N_5897);
or U12383 (N_12383,N_1147,N_865);
nor U12384 (N_12384,N_5898,N_1142);
nor U12385 (N_12385,N_2199,N_4082);
or U12386 (N_12386,N_5955,N_5171);
nor U12387 (N_12387,N_2451,N_6097);
nand U12388 (N_12388,N_507,N_921);
or U12389 (N_12389,N_488,N_4247);
xor U12390 (N_12390,N_802,N_5205);
xor U12391 (N_12391,N_933,N_3220);
or U12392 (N_12392,N_5547,N_2073);
nand U12393 (N_12393,N_1193,N_1441);
nor U12394 (N_12394,N_5269,N_857);
xor U12395 (N_12395,N_2390,N_131);
xor U12396 (N_12396,N_2293,N_5658);
and U12397 (N_12397,N_615,N_3369);
and U12398 (N_12398,N_2244,N_1311);
or U12399 (N_12399,N_4681,N_3151);
and U12400 (N_12400,N_1894,N_4985);
nor U12401 (N_12401,N_2047,N_782);
and U12402 (N_12402,N_1844,N_2175);
or U12403 (N_12403,N_4730,N_4291);
or U12404 (N_12404,N_615,N_2592);
xor U12405 (N_12405,N_3833,N_4119);
xor U12406 (N_12406,N_3764,N_2377);
or U12407 (N_12407,N_3941,N_1135);
or U12408 (N_12408,N_1393,N_2543);
nor U12409 (N_12409,N_6028,N_4472);
nand U12410 (N_12410,N_5357,N_2802);
and U12411 (N_12411,N_3505,N_902);
and U12412 (N_12412,N_4279,N_4650);
and U12413 (N_12413,N_1710,N_562);
xor U12414 (N_12414,N_2748,N_1750);
nand U12415 (N_12415,N_2693,N_151);
or U12416 (N_12416,N_240,N_1100);
and U12417 (N_12417,N_673,N_533);
nor U12418 (N_12418,N_3491,N_5520);
or U12419 (N_12419,N_2991,N_2227);
nor U12420 (N_12420,N_5236,N_2685);
or U12421 (N_12421,N_1847,N_6182);
xor U12422 (N_12422,N_2216,N_2912);
nand U12423 (N_12423,N_4689,N_1642);
and U12424 (N_12424,N_2839,N_6016);
xnor U12425 (N_12425,N_3876,N_4822);
nor U12426 (N_12426,N_2284,N_2619);
or U12427 (N_12427,N_1875,N_6186);
or U12428 (N_12428,N_6120,N_2843);
or U12429 (N_12429,N_1974,N_4221);
and U12430 (N_12430,N_324,N_2751);
nand U12431 (N_12431,N_4152,N_4533);
xor U12432 (N_12432,N_5935,N_5757);
and U12433 (N_12433,N_715,N_4505);
xor U12434 (N_12434,N_1681,N_2609);
xnor U12435 (N_12435,N_5678,N_4848);
or U12436 (N_12436,N_5764,N_5309);
or U12437 (N_12437,N_3253,N_3123);
or U12438 (N_12438,N_305,N_215);
nand U12439 (N_12439,N_5220,N_4930);
nor U12440 (N_12440,N_2091,N_4632);
and U12441 (N_12441,N_1469,N_108);
nand U12442 (N_12442,N_5397,N_3117);
xor U12443 (N_12443,N_2020,N_3913);
nor U12444 (N_12444,N_2367,N_5552);
nor U12445 (N_12445,N_4456,N_3067);
and U12446 (N_12446,N_4138,N_3382);
or U12447 (N_12447,N_4145,N_3833);
or U12448 (N_12448,N_3140,N_13);
nand U12449 (N_12449,N_5656,N_3860);
and U12450 (N_12450,N_1023,N_4870);
nor U12451 (N_12451,N_5395,N_2667);
xor U12452 (N_12452,N_4711,N_1030);
or U12453 (N_12453,N_4445,N_901);
or U12454 (N_12454,N_1198,N_6042);
xor U12455 (N_12455,N_1502,N_730);
nand U12456 (N_12456,N_5443,N_3544);
xor U12457 (N_12457,N_4701,N_1686);
xnor U12458 (N_12458,N_153,N_6096);
or U12459 (N_12459,N_1114,N_4464);
and U12460 (N_12460,N_4818,N_6073);
or U12461 (N_12461,N_4671,N_2939);
and U12462 (N_12462,N_187,N_826);
xnor U12463 (N_12463,N_1804,N_1748);
nand U12464 (N_12464,N_4454,N_3354);
nand U12465 (N_12465,N_953,N_2773);
and U12466 (N_12466,N_1890,N_3731);
xor U12467 (N_12467,N_4384,N_4395);
xnor U12468 (N_12468,N_6092,N_4512);
or U12469 (N_12469,N_2170,N_4948);
and U12470 (N_12470,N_5565,N_2070);
or U12471 (N_12471,N_4512,N_1174);
xnor U12472 (N_12472,N_1043,N_4768);
or U12473 (N_12473,N_2164,N_5952);
xnor U12474 (N_12474,N_4849,N_4075);
nor U12475 (N_12475,N_4252,N_607);
and U12476 (N_12476,N_3988,N_1094);
or U12477 (N_12477,N_1986,N_1622);
or U12478 (N_12478,N_787,N_5615);
nor U12479 (N_12479,N_5674,N_698);
xnor U12480 (N_12480,N_1544,N_360);
nand U12481 (N_12481,N_4530,N_2092);
or U12482 (N_12482,N_4005,N_4486);
or U12483 (N_12483,N_4635,N_1921);
nand U12484 (N_12484,N_1814,N_26);
and U12485 (N_12485,N_3475,N_1113);
or U12486 (N_12486,N_2865,N_4030);
nor U12487 (N_12487,N_6,N_1421);
nor U12488 (N_12488,N_2981,N_5227);
xor U12489 (N_12489,N_5349,N_5664);
nand U12490 (N_12490,N_4331,N_5411);
nand U12491 (N_12491,N_2269,N_852);
nand U12492 (N_12492,N_621,N_4844);
and U12493 (N_12493,N_880,N_1111);
xor U12494 (N_12494,N_3013,N_3424);
or U12495 (N_12495,N_95,N_1614);
and U12496 (N_12496,N_240,N_3486);
nand U12497 (N_12497,N_4157,N_1752);
nand U12498 (N_12498,N_245,N_1195);
nor U12499 (N_12499,N_875,N_4860);
nor U12500 (N_12500,N_8661,N_12209);
nand U12501 (N_12501,N_10443,N_8069);
xnor U12502 (N_12502,N_10361,N_11008);
xor U12503 (N_12503,N_6827,N_7705);
and U12504 (N_12504,N_12266,N_10395);
nor U12505 (N_12505,N_10649,N_7302);
and U12506 (N_12506,N_11027,N_6838);
or U12507 (N_12507,N_9445,N_8977);
xor U12508 (N_12508,N_10129,N_10294);
nand U12509 (N_12509,N_9033,N_7391);
xor U12510 (N_12510,N_6820,N_11753);
nor U12511 (N_12511,N_10137,N_12379);
or U12512 (N_12512,N_8966,N_8407);
nor U12513 (N_12513,N_8745,N_8924);
and U12514 (N_12514,N_10892,N_9755);
xor U12515 (N_12515,N_11393,N_11732);
or U12516 (N_12516,N_7155,N_6548);
xor U12517 (N_12517,N_7852,N_9200);
xor U12518 (N_12518,N_10621,N_10567);
and U12519 (N_12519,N_7175,N_6359);
and U12520 (N_12520,N_7859,N_12395);
and U12521 (N_12521,N_11706,N_6357);
nor U12522 (N_12522,N_7899,N_10359);
xor U12523 (N_12523,N_7385,N_12310);
and U12524 (N_12524,N_10504,N_6912);
nand U12525 (N_12525,N_9170,N_6604);
nand U12526 (N_12526,N_10038,N_6979);
and U12527 (N_12527,N_9881,N_8568);
and U12528 (N_12528,N_8831,N_9034);
nor U12529 (N_12529,N_6618,N_9447);
xnor U12530 (N_12530,N_7309,N_11149);
nor U12531 (N_12531,N_7148,N_6261);
or U12532 (N_12532,N_11644,N_11233);
nand U12533 (N_12533,N_8135,N_9645);
nand U12534 (N_12534,N_8373,N_6797);
nand U12535 (N_12535,N_9048,N_12105);
nor U12536 (N_12536,N_8840,N_10100);
xor U12537 (N_12537,N_9801,N_11400);
nor U12538 (N_12538,N_8038,N_6710);
nand U12539 (N_12539,N_9082,N_10419);
nor U12540 (N_12540,N_8438,N_7355);
nor U12541 (N_12541,N_9816,N_12282);
nand U12542 (N_12542,N_11947,N_11476);
or U12543 (N_12543,N_10958,N_7650);
or U12544 (N_12544,N_7916,N_11782);
or U12545 (N_12545,N_9129,N_8029);
nand U12546 (N_12546,N_12474,N_11000);
nand U12547 (N_12547,N_12316,N_10063);
or U12548 (N_12548,N_11990,N_12060);
or U12549 (N_12549,N_11922,N_9997);
or U12550 (N_12550,N_8208,N_6991);
or U12551 (N_12551,N_8781,N_7218);
nand U12552 (N_12552,N_10424,N_10840);
xnor U12553 (N_12553,N_11908,N_6412);
or U12554 (N_12554,N_11110,N_6553);
nand U12555 (N_12555,N_12162,N_6607);
nor U12556 (N_12556,N_8638,N_7131);
and U12557 (N_12557,N_6642,N_7003);
nand U12558 (N_12558,N_12342,N_10043);
or U12559 (N_12559,N_10408,N_6785);
nor U12560 (N_12560,N_7213,N_6254);
nand U12561 (N_12561,N_8269,N_9282);
or U12562 (N_12562,N_8959,N_11394);
nand U12563 (N_12563,N_8921,N_6471);
nand U12564 (N_12564,N_6365,N_11895);
nand U12565 (N_12565,N_10612,N_10596);
nand U12566 (N_12566,N_6321,N_6971);
xor U12567 (N_12567,N_7297,N_6816);
nor U12568 (N_12568,N_6479,N_10029);
xnor U12569 (N_12569,N_12252,N_7629);
xnor U12570 (N_12570,N_11702,N_9285);
xor U12571 (N_12571,N_11247,N_8030);
nor U12572 (N_12572,N_6341,N_11337);
nor U12573 (N_12573,N_8507,N_8355);
nand U12574 (N_12574,N_8992,N_10304);
nor U12575 (N_12575,N_7861,N_8902);
nor U12576 (N_12576,N_9687,N_6324);
nand U12577 (N_12577,N_10289,N_11840);
or U12578 (N_12578,N_11720,N_12038);
or U12579 (N_12579,N_8542,N_7128);
and U12580 (N_12580,N_6812,N_7681);
nor U12581 (N_12581,N_10593,N_10016);
nor U12582 (N_12582,N_11765,N_11596);
or U12583 (N_12583,N_9540,N_9690);
xnor U12584 (N_12584,N_7221,N_9172);
and U12585 (N_12585,N_7634,N_11818);
nor U12586 (N_12586,N_8915,N_10797);
and U12587 (N_12587,N_9704,N_11885);
xnor U12588 (N_12588,N_9156,N_7036);
xnor U12589 (N_12589,N_9731,N_8478);
or U12590 (N_12590,N_9481,N_7961);
and U12591 (N_12591,N_8983,N_11586);
nand U12592 (N_12592,N_9737,N_11570);
or U12593 (N_12593,N_6727,N_7038);
and U12594 (N_12594,N_11347,N_6796);
and U12595 (N_12595,N_7833,N_9449);
nand U12596 (N_12596,N_7589,N_8109);
nor U12597 (N_12597,N_8596,N_6945);
and U12598 (N_12598,N_12225,N_9463);
xnor U12599 (N_12599,N_9496,N_7362);
nand U12600 (N_12600,N_10557,N_8418);
nand U12601 (N_12601,N_11561,N_6925);
nor U12602 (N_12602,N_8648,N_8404);
or U12603 (N_12603,N_10825,N_6378);
nor U12604 (N_12604,N_12423,N_9774);
and U12605 (N_12605,N_7761,N_7834);
and U12606 (N_12606,N_8446,N_12134);
or U12607 (N_12607,N_6251,N_6696);
and U12608 (N_12608,N_7766,N_7569);
xor U12609 (N_12609,N_11637,N_8066);
or U12610 (N_12610,N_6481,N_10343);
nor U12611 (N_12611,N_7363,N_9161);
nand U12612 (N_12612,N_9069,N_11966);
xnor U12613 (N_12613,N_12152,N_12250);
nor U12614 (N_12614,N_6986,N_10113);
or U12615 (N_12615,N_7343,N_11666);
nor U12616 (N_12616,N_7194,N_8681);
xor U12617 (N_12617,N_6538,N_9091);
and U12618 (N_12618,N_8882,N_6454);
or U12619 (N_12619,N_6411,N_8743);
and U12620 (N_12620,N_11698,N_9185);
nor U12621 (N_12621,N_11106,N_8378);
xor U12622 (N_12622,N_11042,N_8195);
xor U12623 (N_12623,N_10975,N_7535);
or U12624 (N_12624,N_10118,N_7494);
nand U12625 (N_12625,N_10358,N_12472);
nand U12626 (N_12626,N_12253,N_7246);
nand U12627 (N_12627,N_6853,N_7395);
or U12628 (N_12628,N_11681,N_7996);
xor U12629 (N_12629,N_8383,N_10320);
nor U12630 (N_12630,N_11556,N_9832);
or U12631 (N_12631,N_6605,N_11204);
or U12632 (N_12632,N_7054,N_7689);
nor U12633 (N_12633,N_7640,N_12207);
nand U12634 (N_12634,N_7524,N_9889);
or U12635 (N_12635,N_9604,N_12206);
nor U12636 (N_12636,N_6596,N_6401);
and U12637 (N_12637,N_7390,N_9166);
or U12638 (N_12638,N_8453,N_9843);
or U12639 (N_12639,N_6757,N_7151);
xor U12640 (N_12640,N_6992,N_8271);
nand U12641 (N_12641,N_7878,N_12285);
or U12642 (N_12642,N_11676,N_9281);
nand U12643 (N_12643,N_6749,N_11932);
nand U12644 (N_12644,N_9833,N_9238);
or U12645 (N_12645,N_9101,N_8943);
and U12646 (N_12646,N_11580,N_11855);
nor U12647 (N_12647,N_7988,N_8939);
nand U12648 (N_12648,N_9940,N_11134);
and U12649 (N_12649,N_8799,N_10644);
and U12650 (N_12650,N_11468,N_9441);
nand U12651 (N_12651,N_11530,N_7215);
or U12652 (N_12652,N_8416,N_12375);
and U12653 (N_12653,N_9002,N_8004);
and U12654 (N_12654,N_12183,N_9005);
nor U12655 (N_12655,N_6988,N_10619);
or U12656 (N_12656,N_11551,N_8744);
xnor U12657 (N_12657,N_9066,N_8337);
nor U12658 (N_12658,N_10149,N_8808);
nor U12659 (N_12659,N_11948,N_10366);
xor U12660 (N_12660,N_8177,N_11653);
xor U12661 (N_12661,N_7152,N_6928);
nor U12662 (N_12662,N_10531,N_11114);
or U12663 (N_12663,N_11542,N_10480);
nor U12664 (N_12664,N_9522,N_9868);
nand U12665 (N_12665,N_11945,N_7884);
nor U12666 (N_12666,N_7006,N_7739);
nor U12667 (N_12667,N_9517,N_9126);
xnor U12668 (N_12668,N_9696,N_12036);
nor U12669 (N_12669,N_8206,N_8136);
nor U12670 (N_12670,N_10292,N_6865);
xor U12671 (N_12671,N_6620,N_7093);
nor U12672 (N_12672,N_10127,N_11788);
xnor U12673 (N_12673,N_10576,N_10182);
or U12674 (N_12674,N_11277,N_12018);
xnor U12675 (N_12675,N_8079,N_8050);
or U12676 (N_12676,N_6415,N_9919);
xnor U12677 (N_12677,N_11744,N_10044);
and U12678 (N_12678,N_9851,N_11179);
nor U12679 (N_12679,N_9885,N_9168);
nor U12680 (N_12680,N_7450,N_9136);
and U12681 (N_12681,N_6655,N_8925);
or U12682 (N_12682,N_9684,N_9403);
or U12683 (N_12683,N_10210,N_7048);
nor U12684 (N_12684,N_6554,N_6332);
or U12685 (N_12685,N_11246,N_7596);
and U12686 (N_12686,N_8161,N_11043);
and U12687 (N_12687,N_7580,N_11010);
nand U12688 (N_12688,N_10515,N_11343);
xnor U12689 (N_12689,N_8131,N_11673);
and U12690 (N_12690,N_10259,N_10664);
nand U12691 (N_12691,N_7860,N_10690);
and U12692 (N_12692,N_9410,N_10401);
and U12693 (N_12693,N_11583,N_8505);
nand U12694 (N_12694,N_9227,N_10048);
and U12695 (N_12695,N_12227,N_7877);
nor U12696 (N_12696,N_9028,N_9310);
and U12697 (N_12697,N_7314,N_8310);
xor U12698 (N_12698,N_7950,N_12411);
or U12699 (N_12699,N_7276,N_7790);
nor U12700 (N_12700,N_9391,N_11998);
nor U12701 (N_12701,N_7258,N_6643);
xnor U12702 (N_12702,N_12066,N_9261);
and U12703 (N_12703,N_6892,N_10122);
and U12704 (N_12704,N_7044,N_10225);
nand U12705 (N_12705,N_12315,N_8462);
xor U12706 (N_12706,N_12112,N_10852);
nand U12707 (N_12707,N_12337,N_11231);
nand U12708 (N_12708,N_8729,N_7331);
nand U12709 (N_12709,N_9207,N_8223);
nand U12710 (N_12710,N_6255,N_9848);
xnor U12711 (N_12711,N_8742,N_6857);
nor U12712 (N_12712,N_9556,N_8819);
xor U12713 (N_12713,N_6661,N_10367);
xor U12714 (N_12714,N_9877,N_8806);
xnor U12715 (N_12715,N_12330,N_9505);
nand U12716 (N_12716,N_6510,N_9717);
nand U12717 (N_12717,N_8608,N_9679);
and U12718 (N_12718,N_8081,N_7100);
nand U12719 (N_12719,N_7898,N_6869);
and U12720 (N_12720,N_7267,N_8919);
nand U12721 (N_12721,N_6649,N_8549);
xnor U12722 (N_12722,N_7020,N_9867);
and U12723 (N_12723,N_6474,N_6648);
or U12724 (N_12724,N_11993,N_10589);
and U12725 (N_12725,N_10125,N_10310);
and U12726 (N_12726,N_11572,N_11991);
and U12727 (N_12727,N_8725,N_9667);
nand U12728 (N_12728,N_9963,N_10828);
xnor U12729 (N_12729,N_11791,N_11079);
nand U12730 (N_12730,N_9659,N_11016);
and U12731 (N_12731,N_11680,N_8242);
and U12732 (N_12732,N_7149,N_7301);
xnor U12733 (N_12733,N_8379,N_10929);
or U12734 (N_12734,N_9305,N_11062);
or U12735 (N_12735,N_12210,N_6692);
nor U12736 (N_12736,N_11241,N_11436);
xnor U12737 (N_12737,N_12384,N_8699);
nor U12738 (N_12738,N_6885,N_9528);
nand U12739 (N_12739,N_11979,N_9652);
or U12740 (N_12740,N_10688,N_6469);
nor U12741 (N_12741,N_7407,N_11208);
and U12742 (N_12742,N_8879,N_12298);
and U12743 (N_12743,N_9964,N_6614);
or U12744 (N_12744,N_9422,N_12326);
nor U12745 (N_12745,N_10347,N_10606);
xnor U12746 (N_12746,N_7467,N_9694);
xnor U12747 (N_12747,N_8702,N_10339);
and U12748 (N_12748,N_10431,N_6296);
or U12749 (N_12749,N_8757,N_10700);
or U12750 (N_12750,N_7853,N_7164);
and U12751 (N_12751,N_11870,N_7216);
nor U12752 (N_12752,N_12392,N_9723);
nand U12753 (N_12753,N_11694,N_11404);
nor U12754 (N_12754,N_6387,N_7291);
xor U12755 (N_12755,N_7599,N_11466);
xnor U12756 (N_12756,N_10434,N_6734);
and U12757 (N_12757,N_9961,N_8394);
or U12758 (N_12758,N_6368,N_10586);
and U12759 (N_12759,N_9140,N_10667);
nand U12760 (N_12760,N_7588,N_6834);
and U12761 (N_12761,N_7266,N_9968);
nor U12762 (N_12762,N_8942,N_11635);
or U12763 (N_12763,N_6899,N_9529);
xor U12764 (N_12764,N_10168,N_6916);
and U12765 (N_12765,N_9749,N_8016);
nand U12766 (N_12766,N_12051,N_12367);
and U12767 (N_12767,N_6644,N_9150);
xor U12768 (N_12768,N_9052,N_12409);
nor U12769 (N_12769,N_7253,N_8412);
nand U12770 (N_12770,N_11035,N_9480);
nor U12771 (N_12771,N_9794,N_6266);
or U12772 (N_12772,N_7747,N_10227);
or U12773 (N_12773,N_7089,N_11884);
and U12774 (N_12774,N_7477,N_11573);
nand U12775 (N_12775,N_8265,N_8555);
or U12776 (N_12776,N_9991,N_6360);
or U12777 (N_12777,N_6337,N_11670);
or U12778 (N_12778,N_6402,N_10337);
nand U12779 (N_12779,N_7320,N_8635);
xor U12780 (N_12780,N_10499,N_8585);
nor U12781 (N_12781,N_9831,N_7686);
nor U12782 (N_12782,N_11777,N_10422);
nor U12783 (N_12783,N_7393,N_12129);
xor U12784 (N_12784,N_11736,N_10174);
xnor U12785 (N_12785,N_7359,N_11140);
nor U12786 (N_12786,N_6430,N_7341);
xor U12787 (N_12787,N_6426,N_9460);
nand U12788 (N_12788,N_9853,N_7364);
or U12789 (N_12789,N_11200,N_7349);
or U12790 (N_12790,N_8762,N_10086);
nand U12791 (N_12791,N_11816,N_9280);
and U12792 (N_12792,N_8457,N_9539);
and U12793 (N_12793,N_11825,N_11202);
and U12794 (N_12794,N_6798,N_10374);
nand U12795 (N_12795,N_11876,N_7000);
xnor U12796 (N_12796,N_8445,N_7967);
xnor U12797 (N_12797,N_6863,N_6712);
xor U12798 (N_12798,N_8282,N_12398);
nor U12799 (N_12799,N_7510,N_7479);
xnor U12800 (N_12800,N_7051,N_7537);
or U12801 (N_12801,N_11856,N_9870);
xor U12802 (N_12802,N_12374,N_7755);
and U12803 (N_12803,N_8261,N_10888);
and U12804 (N_12804,N_9515,N_7010);
or U12805 (N_12805,N_7224,N_7262);
nor U12806 (N_12806,N_9586,N_8114);
nand U12807 (N_12807,N_10509,N_11823);
nand U12808 (N_12808,N_11089,N_12132);
or U12809 (N_12809,N_9419,N_6637);
nor U12810 (N_12810,N_11899,N_8484);
and U12811 (N_12811,N_8251,N_10271);
nand U12812 (N_12812,N_7365,N_8717);
and U12813 (N_12813,N_9404,N_11227);
nor U12814 (N_12814,N_11734,N_7879);
xor U12815 (N_12815,N_6467,N_8633);
xnor U12816 (N_12816,N_8094,N_11216);
and U12817 (N_12817,N_10352,N_10495);
nor U12818 (N_12818,N_11903,N_7613);
or U12819 (N_12819,N_6775,N_8067);
xor U12820 (N_12820,N_7244,N_12102);
nor U12821 (N_12821,N_6790,N_10811);
xor U12822 (N_12822,N_6974,N_8642);
nand U12823 (N_12823,N_12247,N_10270);
nand U12824 (N_12824,N_6830,N_6349);
and U12825 (N_12825,N_10845,N_10212);
or U12826 (N_12826,N_11321,N_9960);
xor U12827 (N_12827,N_7026,N_11951);
xor U12828 (N_12828,N_8887,N_12350);
nand U12829 (N_12829,N_9163,N_11238);
and U12830 (N_12830,N_10282,N_6636);
nand U12831 (N_12831,N_12339,N_8632);
or U12832 (N_12832,N_9437,N_8503);
nand U12833 (N_12833,N_8089,N_11450);
nor U12834 (N_12834,N_10856,N_9372);
nor U12835 (N_12835,N_12381,N_6294);
nand U12836 (N_12836,N_11812,N_7418);
or U12837 (N_12837,N_11795,N_6819);
nand U12838 (N_12838,N_11607,N_9488);
nor U12839 (N_12839,N_8130,N_11444);
nand U12840 (N_12840,N_10588,N_6756);
and U12841 (N_12841,N_10765,N_7982);
nand U12842 (N_12842,N_11934,N_10409);
and U12843 (N_12843,N_11429,N_9023);
nand U12844 (N_12844,N_9278,N_6369);
and U12845 (N_12845,N_6304,N_11156);
xor U12846 (N_12846,N_8519,N_10733);
nand U12847 (N_12847,N_10918,N_8805);
nor U12848 (N_12848,N_9988,N_9535);
xnor U12849 (N_12849,N_9951,N_8422);
nor U12850 (N_12850,N_11701,N_11215);
nand U12851 (N_12851,N_9154,N_6398);
xnor U12852 (N_12852,N_10795,N_8930);
nand U12853 (N_12853,N_8612,N_11581);
nor U12854 (N_12854,N_8928,N_8440);
nor U12855 (N_12855,N_8031,N_8247);
and U12856 (N_12856,N_10123,N_6610);
and U12857 (N_12857,N_11662,N_8591);
xnor U12858 (N_12858,N_7017,N_7007);
xor U12859 (N_12859,N_9550,N_8554);
xnor U12860 (N_12860,N_9167,N_11726);
nand U12861 (N_12861,N_8215,N_9918);
nand U12862 (N_12862,N_11783,N_7389);
xor U12863 (N_12863,N_10972,N_10067);
or U12864 (N_12864,N_10539,N_12061);
or U12865 (N_12865,N_8201,N_10444);
or U12866 (N_12866,N_11700,N_7958);
or U12867 (N_12867,N_11859,N_10732);
or U12868 (N_12868,N_10997,N_9985);
nand U12869 (N_12869,N_11597,N_9318);
and U12870 (N_12870,N_6702,N_12107);
or U12871 (N_12871,N_10948,N_8342);
nand U12872 (N_12872,N_9093,N_7519);
and U12873 (N_12873,N_8617,N_6611);
xor U12874 (N_12874,N_7290,N_10411);
and U12875 (N_12875,N_6285,N_11953);
nand U12876 (N_12876,N_6313,N_11535);
nand U12877 (N_12877,N_10506,N_7584);
nor U12878 (N_12878,N_8352,N_8539);
nor U12879 (N_12879,N_8059,N_6344);
and U12880 (N_12880,N_10559,N_9811);
or U12881 (N_12881,N_8405,N_12160);
or U12882 (N_12882,N_6564,N_8832);
or U12883 (N_12883,N_8687,N_11747);
xor U12884 (N_12884,N_7715,N_10062);
xor U12885 (N_12885,N_12419,N_11128);
xnor U12886 (N_12886,N_10562,N_8403);
nand U12887 (N_12887,N_10010,N_9428);
and U12888 (N_12888,N_9152,N_11467);
xnor U12889 (N_12889,N_6780,N_11316);
xnor U12890 (N_12890,N_10570,N_11577);
and U12891 (N_12891,N_11040,N_9417);
and U12892 (N_12892,N_6958,N_9557);
nand U12893 (N_12893,N_12279,N_8634);
nor U12894 (N_12894,N_12033,N_6488);
or U12895 (N_12895,N_8931,N_10702);
and U12896 (N_12896,N_11323,N_7618);
nor U12897 (N_12897,N_12208,N_10804);
or U12898 (N_12898,N_9654,N_12035);
nand U12899 (N_12899,N_9125,N_11964);
nand U12900 (N_12900,N_7965,N_10818);
nand U12901 (N_12901,N_12261,N_6422);
nor U12902 (N_12902,N_7807,N_10105);
nand U12903 (N_12903,N_7098,N_11199);
xor U12904 (N_12904,N_6837,N_8372);
or U12905 (N_12905,N_10283,N_8237);
nand U12906 (N_12906,N_11956,N_11829);
nor U12907 (N_12907,N_9825,N_11959);
or U12908 (N_12908,N_7606,N_9845);
nand U12909 (N_12909,N_12044,N_9804);
or U12910 (N_12910,N_8852,N_7882);
and U12911 (N_12911,N_11933,N_12133);
nor U12912 (N_12912,N_12139,N_8715);
nand U12913 (N_12913,N_11015,N_6482);
or U12914 (N_12914,N_6399,N_9102);
and U12915 (N_12915,N_6382,N_8151);
and U12916 (N_12916,N_9616,N_10050);
xnor U12917 (N_12917,N_11995,N_7095);
or U12918 (N_12918,N_8837,N_8794);
nor U12919 (N_12919,N_9178,N_8472);
and U12920 (N_12920,N_7876,N_8771);
nor U12921 (N_12921,N_11153,N_6758);
or U12922 (N_12922,N_9976,N_11712);
or U12923 (N_12923,N_8970,N_11348);
xnor U12924 (N_12924,N_10274,N_7452);
xnor U12925 (N_12925,N_9672,N_10145);
xor U12926 (N_12926,N_7917,N_12443);
nand U12927 (N_12927,N_11645,N_9987);
nor U12928 (N_12928,N_7310,N_10971);
nor U12929 (N_12929,N_12106,N_12043);
or U12930 (N_12930,N_6770,N_6279);
nor U12931 (N_12931,N_10141,N_11038);
nor U12932 (N_12932,N_7920,N_7333);
xnor U12933 (N_12933,N_9316,N_9840);
or U12934 (N_12934,N_8768,N_9012);
or U12935 (N_12935,N_7957,N_10998);
and U12936 (N_12936,N_10410,N_8708);
nor U12937 (N_12937,N_11382,N_6322);
or U12938 (N_12938,N_9277,N_10109);
and U12939 (N_12939,N_7931,N_11330);
and U12940 (N_12940,N_7597,N_11674);
or U12941 (N_12941,N_8609,N_9617);
or U12942 (N_12942,N_8267,N_7072);
nand U12943 (N_12943,N_10643,N_8613);
nor U12944 (N_12944,N_9374,N_12294);
or U12945 (N_12945,N_12213,N_7404);
or U12946 (N_12946,N_9958,N_9670);
nand U12947 (N_12947,N_6566,N_12177);
nand U12948 (N_12948,N_6393,N_6966);
nor U12949 (N_12949,N_9354,N_12497);
xnor U12950 (N_12950,N_12414,N_12390);
xnor U12951 (N_12951,N_9903,N_8981);
nand U12952 (N_12952,N_11302,N_10610);
and U12953 (N_12953,N_8597,N_10884);
nor U12954 (N_12954,N_6606,N_8772);
or U12955 (N_12955,N_12237,N_6733);
and U12956 (N_12956,N_6485,N_7008);
nand U12957 (N_12957,N_11313,N_7166);
nor U12958 (N_12958,N_11147,N_6303);
xnor U12959 (N_12959,N_10116,N_9132);
nor U12960 (N_12960,N_8898,N_8938);
nor U12961 (N_12961,N_11102,N_8249);
nor U12962 (N_12962,N_10671,N_7992);
or U12963 (N_12963,N_9145,N_12344);
nand U12964 (N_12964,N_11050,N_11066);
xor U12965 (N_12965,N_8494,N_9138);
and U12966 (N_12966,N_10827,N_7154);
and U12967 (N_12967,N_9079,N_6498);
nand U12968 (N_12968,N_9160,N_10886);
and U12969 (N_12969,N_6846,N_9359);
and U12970 (N_12970,N_8469,N_8964);
nand U12971 (N_12971,N_10778,N_7810);
xnor U12972 (N_12972,N_10368,N_10735);
nor U12973 (N_12973,N_7161,N_8423);
nor U12974 (N_12974,N_12030,N_6372);
xor U12975 (N_12975,N_7822,N_11418);
nand U12976 (N_12976,N_8284,N_8752);
nand U12977 (N_12977,N_8060,N_11322);
nor U12978 (N_12978,N_11285,N_8436);
or U12979 (N_12979,N_7784,N_6257);
or U12980 (N_12980,N_6665,N_10089);
and U12981 (N_12981,N_9920,N_10743);
or U12982 (N_12982,N_6932,N_11270);
nand U12983 (N_12983,N_9324,N_9369);
nor U12984 (N_12984,N_10286,N_9175);
or U12985 (N_12985,N_10486,N_9311);
nor U12986 (N_12986,N_8520,N_9336);
nand U12987 (N_12987,N_7004,N_9613);
nor U12988 (N_12988,N_10860,N_8560);
and U12989 (N_12989,N_6659,N_11594);
nand U12990 (N_12990,N_9839,N_10976);
or U12991 (N_12991,N_7841,N_6558);
xor U12992 (N_12992,N_8967,N_10449);
nor U12993 (N_12993,N_7962,N_10202);
nor U12994 (N_12994,N_10802,N_8172);
xnor U12995 (N_12995,N_12169,N_9551);
xor U12996 (N_12996,N_8605,N_7146);
nor U12997 (N_12997,N_10180,N_11715);
nand U12998 (N_12998,N_9878,N_10071);
nor U12999 (N_12999,N_7240,N_11029);
nand U13000 (N_13000,N_6500,N_11487);
nand U13001 (N_13001,N_9262,N_8798);
and U13002 (N_13002,N_9910,N_11972);
and U13003 (N_13003,N_8953,N_8755);
or U13004 (N_13004,N_10636,N_11006);
or U13005 (N_13005,N_10307,N_10662);
or U13006 (N_13006,N_11863,N_10999);
nor U13007 (N_13007,N_8991,N_6433);
or U13008 (N_13008,N_7986,N_10841);
nor U13009 (N_13009,N_12371,N_11425);
nand U13010 (N_13010,N_9561,N_8510);
and U13011 (N_13011,N_8455,N_7210);
nand U13012 (N_13012,N_12185,N_11297);
and U13013 (N_13013,N_9527,N_8073);
xnor U13014 (N_13014,N_9500,N_7185);
xor U13015 (N_13015,N_9494,N_9884);
and U13016 (N_13016,N_6600,N_10169);
xor U13017 (N_13017,N_9837,N_11937);
xnor U13018 (N_13018,N_11340,N_11447);
nor U13019 (N_13019,N_8111,N_12343);
and U13020 (N_13020,N_9284,N_10949);
or U13021 (N_13021,N_6657,N_11786);
nor U13022 (N_13022,N_11718,N_8684);
or U13023 (N_13023,N_11997,N_12488);
nand U13024 (N_13024,N_10625,N_9942);
xor U13025 (N_13025,N_6813,N_10839);
or U13026 (N_13026,N_8225,N_8792);
and U13027 (N_13027,N_9253,N_9695);
or U13028 (N_13028,N_7081,N_11669);
and U13029 (N_13029,N_11668,N_9116);
and U13030 (N_13030,N_8381,N_11186);
nand U13031 (N_13031,N_11207,N_8302);
nand U13032 (N_13032,N_11707,N_8593);
nand U13033 (N_13033,N_9890,N_12231);
nand U13034 (N_13034,N_11071,N_11046);
and U13035 (N_13035,N_12040,N_7520);
or U13036 (N_13036,N_11251,N_7538);
nor U13037 (N_13037,N_9521,N_10199);
or U13038 (N_13038,N_7406,N_6929);
nor U13039 (N_13039,N_8795,N_11819);
or U13040 (N_13040,N_11733,N_8914);
or U13041 (N_13041,N_11873,N_6994);
nand U13042 (N_13042,N_7358,N_11924);
nor U13043 (N_13043,N_7782,N_7127);
xnor U13044 (N_13044,N_9328,N_6389);
nor U13045 (N_13045,N_12017,N_9053);
xor U13046 (N_13046,N_11176,N_7738);
nor U13047 (N_13047,N_9634,N_11549);
xor U13048 (N_13048,N_12069,N_11505);
xor U13049 (N_13049,N_10981,N_8387);
nor U13050 (N_13050,N_7701,N_11472);
and U13051 (N_13051,N_9498,N_9567);
nand U13052 (N_13052,N_7281,N_11699);
nand U13053 (N_13053,N_11282,N_10575);
and U13054 (N_13054,N_11054,N_9649);
or U13055 (N_13055,N_8784,N_11952);
xor U13056 (N_13056,N_7742,N_10219);
xnor U13057 (N_13057,N_9299,N_8506);
and U13058 (N_13058,N_8780,N_8487);
xor U13059 (N_13059,N_9917,N_8384);
or U13060 (N_13060,N_8489,N_7909);
xor U13061 (N_13061,N_9573,N_9224);
and U13062 (N_13062,N_12013,N_9673);
or U13063 (N_13063,N_7083,N_7059);
nand U13064 (N_13064,N_9797,N_11832);
xor U13065 (N_13065,N_6658,N_9425);
or U13066 (N_13066,N_7202,N_8132);
nand U13067 (N_13067,N_8231,N_7942);
xor U13068 (N_13068,N_7769,N_10291);
and U13069 (N_13069,N_11624,N_7717);
or U13070 (N_13070,N_10396,N_7129);
and U13071 (N_13071,N_10853,N_12348);
nand U13072 (N_13072,N_9476,N_11077);
nor U13073 (N_13073,N_7420,N_7470);
or U13074 (N_13074,N_12446,N_7346);
nand U13075 (N_13075,N_8552,N_12100);
or U13076 (N_13076,N_6949,N_11776);
nor U13077 (N_13077,N_10099,N_9977);
nand U13078 (N_13078,N_10541,N_7970);
nand U13079 (N_13079,N_11957,N_10257);
or U13080 (N_13080,N_12483,N_7071);
nand U13081 (N_13081,N_10558,N_6745);
and U13082 (N_13082,N_8408,N_8474);
nor U13083 (N_13083,N_10036,N_8158);
nand U13084 (N_13084,N_7890,N_9806);
nand U13085 (N_13085,N_9271,N_11705);
or U13086 (N_13086,N_12003,N_11521);
or U13087 (N_13087,N_9531,N_8245);
xor U13088 (N_13088,N_7517,N_10990);
nand U13089 (N_13089,N_11529,N_6981);
xor U13090 (N_13090,N_6326,N_9155);
xnor U13091 (N_13091,N_6268,N_8358);
nor U13092 (N_13092,N_7143,N_10058);
or U13093 (N_13093,N_9744,N_10093);
xor U13094 (N_13094,N_7553,N_8420);
nor U13095 (N_13095,N_9474,N_11223);
nor U13096 (N_13096,N_8450,N_7582);
or U13097 (N_13097,N_8263,N_6452);
nand U13098 (N_13098,N_9073,N_9803);
and U13099 (N_13099,N_10450,N_9137);
nand U13100 (N_13100,N_7602,N_7399);
xor U13101 (N_13101,N_7727,N_11014);
nand U13102 (N_13102,N_6741,N_7227);
xnor U13103 (N_13103,N_10583,N_10960);
xnor U13104 (N_13104,N_8645,N_9644);
nand U13105 (N_13105,N_11004,N_10622);
xor U13106 (N_13106,N_6647,N_9244);
or U13107 (N_13107,N_8181,N_6709);
nand U13108 (N_13108,N_10695,N_9021);
nor U13109 (N_13109,N_9092,N_7340);
or U13110 (N_13110,N_8058,N_9880);
xnor U13111 (N_13111,N_6891,N_10862);
xnor U13112 (N_13112,N_7043,N_11272);
nand U13113 (N_13113,N_12050,N_9757);
and U13114 (N_13114,N_6698,N_6436);
and U13115 (N_13115,N_9603,N_9983);
or U13116 (N_13116,N_11403,N_10684);
nor U13117 (N_13117,N_7022,N_11898);
nand U13118 (N_13118,N_7226,N_12272);
nand U13119 (N_13119,N_9165,N_12292);
xor U13120 (N_13120,N_11619,N_12141);
or U13121 (N_13121,N_8958,N_8351);
xnor U13122 (N_13122,N_6927,N_8148);
and U13123 (N_13123,N_7581,N_9298);
or U13124 (N_13124,N_6650,N_6946);
nor U13125 (N_13125,N_7987,N_8734);
nor U13126 (N_13126,N_10474,N_10922);
or U13127 (N_13127,N_8912,N_11663);
and U13128 (N_13128,N_11742,N_11896);
nor U13129 (N_13129,N_11914,N_11779);
nand U13130 (N_13130,N_9356,N_9675);
xnor U13131 (N_13131,N_7133,N_10630);
xor U13132 (N_13132,N_8262,N_9866);
nor U13133 (N_13133,N_8185,N_11253);
nand U13134 (N_13134,N_7529,N_10142);
or U13135 (N_13135,N_6451,N_12318);
and U13136 (N_13136,N_9429,N_8566);
or U13137 (N_13137,N_9346,N_7242);
xor U13138 (N_13138,N_10108,N_9829);
xnor U13139 (N_13139,N_7062,N_9068);
nor U13140 (N_13140,N_7688,N_8399);
nor U13141 (N_13141,N_10341,N_9483);
xnor U13142 (N_13142,N_6714,N_10773);
nor U13143 (N_13143,N_9911,N_10910);
nor U13144 (N_13144,N_11329,N_11890);
nor U13145 (N_13145,N_10512,N_8210);
nand U13146 (N_13146,N_10849,N_8227);
and U13147 (N_13147,N_10308,N_10387);
xnor U13148 (N_13148,N_7162,N_8301);
and U13149 (N_13149,N_6339,N_12385);
xnor U13150 (N_13150,N_9606,N_6298);
nor U13151 (N_13151,N_8194,N_9376);
nand U13152 (N_13152,N_9657,N_9432);
nand U13153 (N_13153,N_6288,N_9257);
nand U13154 (N_13154,N_6516,N_6286);
xnor U13155 (N_13155,N_10085,N_9856);
xnor U13156 (N_13156,N_9248,N_8588);
nand U13157 (N_13157,N_9229,N_10920);
nand U13158 (N_13158,N_11341,N_11868);
or U13159 (N_13159,N_8544,N_9366);
nor U13160 (N_13160,N_8179,N_10457);
xor U13161 (N_13161,N_8847,N_10383);
nor U13162 (N_13162,N_7296,N_10425);
or U13163 (N_13163,N_11243,N_10554);
nor U13164 (N_13164,N_7892,N_9992);
xor U13165 (N_13165,N_6894,N_9725);
or U13166 (N_13166,N_9276,N_11999);
and U13167 (N_13167,N_6318,N_7433);
nor U13168 (N_13168,N_10460,N_11755);
nor U13169 (N_13169,N_9941,N_7801);
nand U13170 (N_13170,N_11911,N_6703);
nand U13171 (N_13171,N_11120,N_7874);
xor U13172 (N_13172,N_10488,N_9728);
nor U13173 (N_13173,N_12244,N_7424);
xor U13174 (N_13174,N_10574,N_11434);
nand U13175 (N_13175,N_11891,N_11386);
or U13176 (N_13176,N_8511,N_7439);
and U13177 (N_13177,N_10598,N_9904);
nor U13178 (N_13178,N_8033,N_6904);
nand U13179 (N_13179,N_12026,N_7635);
or U13180 (N_13180,N_10633,N_8601);
nand U13181 (N_13181,N_6805,N_8824);
nand U13182 (N_13182,N_12161,N_9680);
and U13183 (N_13183,N_9349,N_8649);
nor U13184 (N_13184,N_8843,N_10076);
or U13185 (N_13185,N_7005,N_8890);
nor U13186 (N_13186,N_6507,N_6954);
nor U13187 (N_13187,N_9860,N_6937);
or U13188 (N_13188,N_6308,N_10171);
or U13189 (N_13189,N_8348,N_9274);
nand U13190 (N_13190,N_6478,N_8916);
or U13191 (N_13191,N_11391,N_9456);
xnor U13192 (N_13192,N_9001,N_10511);
or U13193 (N_13193,N_6706,N_7283);
nand U13194 (N_13194,N_8518,N_7063);
and U13195 (N_13195,N_10111,N_10796);
nand U13196 (N_13196,N_7598,N_10191);
and U13197 (N_13197,N_11003,N_6923);
and U13198 (N_13198,N_6466,N_10415);
or U13199 (N_13199,N_10240,N_6549);
or U13200 (N_13200,N_12383,N_8865);
and U13201 (N_13201,N_8490,N_12267);
or U13202 (N_13202,N_10717,N_8655);
or U13203 (N_13203,N_9553,N_11659);
nand U13204 (N_13204,N_10658,N_9407);
xnor U13205 (N_13205,N_9591,N_12425);
and U13206 (N_13206,N_9895,N_10628);
xor U13207 (N_13207,N_7846,N_7661);
nand U13208 (N_13208,N_11390,N_11492);
or U13209 (N_13209,N_11051,N_10248);
nand U13210 (N_13210,N_11703,N_11536);
nor U13211 (N_13211,N_7702,N_10665);
nor U13212 (N_13212,N_10781,N_6909);
xnor U13213 (N_13213,N_8811,N_11754);
or U13214 (N_13214,N_6594,N_8385);
or U13215 (N_13215,N_9929,N_11910);
or U13216 (N_13216,N_7720,N_9503);
nand U13217 (N_13217,N_7241,N_12144);
nor U13218 (N_13218,N_11608,N_8093);
nand U13219 (N_13219,N_7971,N_8761);
nor U13220 (N_13220,N_8698,N_12116);
and U13221 (N_13221,N_6350,N_7765);
xnor U13222 (N_13222,N_6978,N_7201);
and U13223 (N_13223,N_9711,N_11371);
and U13224 (N_13224,N_7697,N_9159);
nor U13225 (N_13225,N_11475,N_10500);
or U13226 (N_13226,N_9206,N_8000);
or U13227 (N_13227,N_6771,N_9891);
nor U13228 (N_13228,N_8631,N_10580);
xor U13229 (N_13229,N_11546,N_9533);
nand U13230 (N_13230,N_6726,N_9808);
and U13231 (N_13231,N_6367,N_10740);
and U13232 (N_13232,N_9943,N_10678);
xnor U13233 (N_13233,N_7646,N_7076);
or U13234 (N_13234,N_10790,N_8775);
nand U13235 (N_13235,N_10228,N_7668);
xor U13236 (N_13236,N_7388,N_8774);
or U13237 (N_13237,N_6437,N_7550);
xor U13238 (N_13238,N_8018,N_11267);
and U13239 (N_13239,N_8291,N_12095);
nand U13240 (N_13240,N_7248,N_9235);
nand U13241 (N_13241,N_9440,N_9632);
xor U13242 (N_13242,N_12465,N_6400);
nand U13243 (N_13243,N_9542,N_11333);
and U13244 (N_13244,N_8553,N_10775);
nor U13245 (N_13245,N_6501,N_8020);
nand U13246 (N_13246,N_10462,N_9029);
and U13247 (N_13247,N_8306,N_11011);
or U13248 (N_13248,N_6333,N_6730);
nor U13249 (N_13249,N_8512,N_6561);
nor U13250 (N_13250,N_6690,N_10595);
and U13251 (N_13251,N_11469,N_10984);
nand U13252 (N_13252,N_10254,N_8639);
xnor U13253 (N_13253,N_9740,N_10154);
nand U13254 (N_13254,N_6764,N_10049);
xor U13255 (N_13255,N_10683,N_7465);
or U13256 (N_13256,N_8380,N_10745);
or U13257 (N_13257,N_12490,N_9482);
or U13258 (N_13258,N_10088,N_11366);
and U13259 (N_13259,N_11633,N_7798);
xor U13260 (N_13260,N_7699,N_6817);
and U13261 (N_13261,N_10530,N_8234);
nand U13262 (N_13262,N_7559,N_9572);
xor U13263 (N_13263,N_7844,N_9450);
or U13264 (N_13264,N_9350,N_6373);
or U13265 (N_13265,N_12496,N_6645);
and U13266 (N_13266,N_8413,N_11560);
and U13267 (N_13267,N_9260,N_9552);
nor U13268 (N_13268,N_9876,N_8080);
xnor U13269 (N_13269,N_6800,N_11099);
nor U13270 (N_13270,N_7787,N_8178);
and U13271 (N_13271,N_11994,N_8486);
and U13272 (N_13272,N_10681,N_7374);
or U13273 (N_13273,N_10782,N_8107);
nand U13274 (N_13274,N_7126,N_8275);
nor U13275 (N_13275,N_10760,N_11482);
xor U13276 (N_13276,N_11969,N_6867);
xor U13277 (N_13277,N_8314,N_7250);
and U13278 (N_13278,N_8374,N_11100);
nand U13279 (N_13279,N_10523,N_7123);
nor U13280 (N_13280,N_6772,N_10394);
nand U13281 (N_13281,N_12479,N_12216);
nand U13282 (N_13282,N_11078,N_8818);
nor U13283 (N_13283,N_8845,N_10373);
nand U13284 (N_13284,N_10463,N_10054);
nor U13285 (N_13285,N_8697,N_11543);
and U13286 (N_13286,N_9266,N_10503);
or U13287 (N_13287,N_7002,N_6864);
and U13288 (N_13288,N_8285,N_6272);
nand U13289 (N_13289,N_8183,N_9339);
and U13290 (N_13290,N_8312,N_11510);
and U13291 (N_13291,N_9631,N_10332);
xnor U13292 (N_13292,N_7530,N_12219);
nor U13293 (N_13293,N_8941,N_12236);
and U13294 (N_13294,N_6441,N_6397);
and U13295 (N_13295,N_11168,N_10102);
and U13296 (N_13296,N_9058,N_10249);
and U13297 (N_13297,N_7736,N_7514);
and U13298 (N_13298,N_10402,N_9916);
and U13299 (N_13299,N_10390,N_8982);
xnor U13300 (N_13300,N_9059,N_9793);
or U13301 (N_13301,N_10068,N_8705);
or U13302 (N_13302,N_9089,N_10516);
xnor U13303 (N_13303,N_8703,N_8203);
nor U13304 (N_13304,N_10040,N_8854);
or U13305 (N_13305,N_10211,N_10519);
xor U13306 (N_13306,N_10439,N_9511);
and U13307 (N_13307,N_10479,N_6848);
xor U13308 (N_13308,N_10866,N_7721);
xor U13309 (N_13309,N_8102,N_9383);
xor U13310 (N_13310,N_7278,N_6705);
or U13311 (N_13311,N_6667,N_11101);
xor U13312 (N_13312,N_8233,N_7326);
and U13313 (N_13313,N_8504,N_6634);
and U13314 (N_13314,N_11857,N_9642);
nor U13315 (N_13315,N_6940,N_11249);
nor U13316 (N_13316,N_10942,N_6735);
nand U13317 (N_13317,N_6264,N_8565);
nor U13318 (N_13318,N_8628,N_7678);
xnor U13319 (N_13319,N_7413,N_9792);
xnor U13320 (N_13320,N_11848,N_6963);
or U13321 (N_13321,N_6858,N_10932);
xor U13322 (N_13322,N_8259,N_10364);
xnor U13323 (N_13323,N_8133,N_9071);
and U13324 (N_13324,N_9664,N_9751);
xor U13325 (N_13325,N_12417,N_10484);
and U13326 (N_13326,N_7182,N_10883);
and U13327 (N_13327,N_7733,N_7895);
or U13328 (N_13328,N_9842,N_10489);
xnor U13329 (N_13329,N_9615,N_10891);
or U13330 (N_13330,N_6998,N_9022);
nand U13331 (N_13331,N_12092,N_9582);
and U13332 (N_13332,N_6305,N_10008);
or U13333 (N_13333,N_6829,N_10138);
and U13334 (N_13334,N_10003,N_10978);
and U13335 (N_13335,N_9131,N_11511);
nand U13336 (N_13336,N_9746,N_9750);
or U13337 (N_13337,N_11122,N_10490);
nand U13338 (N_13338,N_10639,N_6576);
nor U13339 (N_13339,N_6996,N_11018);
nand U13340 (N_13340,N_9040,N_12265);
nor U13341 (N_13341,N_6582,N_11210);
xnor U13342 (N_13342,N_11162,N_9078);
xnor U13343 (N_13343,N_8760,N_7968);
xnor U13344 (N_13344,N_8447,N_10875);
nor U13345 (N_13345,N_11518,N_6911);
nor U13346 (N_13346,N_8624,N_8305);
and U13347 (N_13347,N_8886,N_9246);
nor U13348 (N_13348,N_7256,N_8714);
and U13349 (N_13349,N_10293,N_6767);
and U13350 (N_13350,N_11728,N_6347);
or U13351 (N_13351,N_9656,N_12099);
xor U13352 (N_13352,N_8759,N_10466);
and U13353 (N_13353,N_9931,N_7140);
nor U13354 (N_13354,N_12150,N_7973);
nor U13355 (N_13355,N_6355,N_10793);
nand U13356 (N_13356,N_7976,N_7921);
xor U13357 (N_13357,N_11360,N_8767);
xnor U13358 (N_13358,N_9643,N_10871);
nor U13359 (N_13359,N_11121,N_12180);
nand U13360 (N_13360,N_10565,N_8421);
xor U13361 (N_13361,N_9894,N_8174);
nand U13362 (N_13362,N_9118,N_9008);
and U13363 (N_13363,N_7471,N_8365);
nor U13364 (N_13364,N_9703,N_9579);
or U13365 (N_13365,N_10597,N_6724);
nor U13366 (N_13366,N_11061,N_6390);
nand U13367 (N_13367,N_7741,N_10017);
xor U13368 (N_13368,N_7758,N_11967);
or U13369 (N_13369,N_12394,N_10447);
xnor U13370 (N_13370,N_10037,N_11031);
nor U13371 (N_13371,N_6964,N_10943);
or U13372 (N_13372,N_9936,N_8191);
or U13373 (N_13373,N_11423,N_10299);
and U13374 (N_13374,N_8517,N_6348);
nor U13375 (N_13375,N_11344,N_11295);
nor U13376 (N_13376,N_6729,N_6574);
and U13377 (N_13377,N_12410,N_6639);
nand U13378 (N_13378,N_7435,N_12334);
nand U13379 (N_13379,N_12270,N_9081);
or U13380 (N_13380,N_12495,N_11656);
or U13381 (N_13381,N_11158,N_11401);
or U13382 (N_13382,N_8783,N_9173);
nor U13383 (N_13383,N_8524,N_8712);
xnor U13384 (N_13384,N_7370,N_10594);
nor U13385 (N_13385,N_10986,N_8475);
nand U13386 (N_13386,N_8527,N_9308);
or U13387 (N_13387,N_11372,N_9726);
or U13388 (N_13388,N_11288,N_8741);
nor U13389 (N_13389,N_11501,N_9063);
xnor U13390 (N_13390,N_11274,N_10448);
nand U13391 (N_13391,N_12325,N_8159);
nor U13392 (N_13392,N_9771,N_7850);
or U13393 (N_13393,N_8454,N_10226);
and U13394 (N_13394,N_12204,N_11451);
nand U13395 (N_13395,N_6434,N_6406);
nand U13396 (N_13396,N_8500,N_7532);
nor U13397 (N_13397,N_7683,N_11229);
xor U13398 (N_13398,N_11654,N_12304);
xnor U13399 (N_13399,N_7745,N_7783);
nand U13400 (N_13400,N_9559,N_9592);
nor U13401 (N_13401,N_6505,N_6654);
or U13402 (N_13402,N_10747,N_10666);
and U13403 (N_13403,N_10236,N_8766);
nand U13404 (N_13404,N_8789,N_9122);
nand U13405 (N_13405,N_10335,N_8564);
or U13406 (N_13406,N_7512,N_10965);
nand U13407 (N_13407,N_11532,N_12477);
nand U13408 (N_13408,N_7605,N_7053);
and U13409 (N_13409,N_10964,N_10090);
xor U13410 (N_13410,N_7662,N_6440);
xnor U13411 (N_13411,N_8693,N_11389);
nor U13412 (N_13412,N_7977,N_10117);
and U13413 (N_13413,N_9758,N_6555);
or U13414 (N_13414,N_10130,N_8957);
and U13415 (N_13415,N_11268,N_8888);
xnor U13416 (N_13416,N_7074,N_11124);
or U13417 (N_13417,N_8270,N_6763);
xor U13418 (N_13418,N_10267,N_10938);
nor U13419 (N_13419,N_6737,N_10529);
nand U13420 (N_13420,N_8220,N_7547);
xnor U13421 (N_13421,N_10200,N_11749);
nor U13422 (N_13422,N_7748,N_7719);
nor U13423 (N_13423,N_8685,N_11385);
and U13424 (N_13424,N_10072,N_12084);
nand U13425 (N_13425,N_7107,N_10417);
nand U13426 (N_13426,N_10715,N_10066);
xnor U13427 (N_13427,N_7934,N_10025);
or U13428 (N_13428,N_11860,N_8777);
xor U13429 (N_13429,N_10455,N_10993);
or U13430 (N_13430,N_8536,N_11762);
nand U13431 (N_13431,N_11965,N_6860);
xnor U13432 (N_13432,N_11093,N_8590);
xnor U13433 (N_13433,N_11763,N_6896);
or U13434 (N_13434,N_6824,N_6751);
nand U13435 (N_13435,N_9705,N_7275);
or U13436 (N_13436,N_9288,N_6617);
nand U13437 (N_13437,N_11355,N_6552);
xor U13438 (N_13438,N_6679,N_11622);
nand U13439 (N_13439,N_9113,N_8678);
nand U13440 (N_13440,N_9187,N_8993);
and U13441 (N_13441,N_8770,N_10263);
or U13442 (N_13442,N_12364,N_7443);
nand U13443 (N_13443,N_7103,N_8753);
or U13444 (N_13444,N_8236,N_11893);
or U13445 (N_13445,N_11799,N_8862);
or U13446 (N_13446,N_9773,N_8187);
nand U13447 (N_13447,N_9562,N_8055);
and U13448 (N_13448,N_7312,N_10679);
or U13449 (N_13449,N_9956,N_6331);
and U13450 (N_13450,N_8754,N_12098);
nand U13451 (N_13451,N_6652,N_7680);
xnor U13452 (N_13452,N_6522,N_7750);
or U13453 (N_13453,N_7457,N_11584);
xnor U13454 (N_13454,N_8496,N_7138);
nor U13455 (N_13455,N_7671,N_8406);
nor U13456 (N_13456,N_7272,N_7405);
nor U13457 (N_13457,N_9423,N_11774);
and U13458 (N_13458,N_10272,N_9761);
or U13459 (N_13459,N_9926,N_10707);
nor U13460 (N_13460,N_8700,N_9312);
xor U13461 (N_13461,N_6989,N_10864);
nor U13462 (N_13462,N_11651,N_10380);
or U13463 (N_13463,N_6301,N_7698);
nor U13464 (N_13464,N_9300,N_8084);
and U13465 (N_13465,N_12289,N_10573);
and U13466 (N_13466,N_8973,N_11064);
nor U13467 (N_13467,N_8526,N_10538);
xor U13468 (N_13468,N_12079,N_9736);
and U13469 (N_13469,N_8790,N_9514);
nor U13470 (N_13470,N_11159,N_9946);
or U13471 (N_13471,N_7409,N_11486);
and U13472 (N_13472,N_12113,N_12428);
and U13473 (N_13473,N_10692,N_11287);
and U13474 (N_13474,N_9371,N_7282);
and U13475 (N_13475,N_11407,N_7648);
nor U13476 (N_13476,N_8615,N_7354);
nor U13477 (N_13477,N_7583,N_12025);
or U13478 (N_13478,N_11955,N_7371);
and U13479 (N_13479,N_6513,N_8116);
nor U13480 (N_13480,N_6589,N_8077);
nor U13481 (N_13481,N_6854,N_8990);
xnor U13482 (N_13482,N_7633,N_12198);
nand U13483 (N_13483,N_6330,N_8786);
xnor U13484 (N_13484,N_11262,N_7025);
or U13485 (N_13485,N_8758,N_11851);
and U13486 (N_13486,N_9196,N_9104);
and U13487 (N_13487,N_7791,N_11284);
nand U13488 (N_13488,N_8849,N_12499);
xor U13489 (N_13489,N_10303,N_12256);
nand U13490 (N_13490,N_8252,N_10354);
or U13491 (N_13491,N_11721,N_11030);
or U13492 (N_13492,N_12466,N_9329);
or U13493 (N_13493,N_9241,N_6850);
and U13494 (N_13494,N_9106,N_6539);
nand U13495 (N_13495,N_10729,N_11443);
or U13496 (N_13496,N_7744,N_10941);
or U13497 (N_13497,N_9430,N_9954);
nand U13498 (N_13498,N_9355,N_7636);
or U13499 (N_13499,N_9915,N_11539);
or U13500 (N_13500,N_12015,N_12074);
xor U13501 (N_13501,N_10893,N_10363);
nor U13502 (N_13502,N_7767,N_8646);
and U13503 (N_13503,N_11837,N_7360);
or U13504 (N_13504,N_6609,N_6948);
nor U13505 (N_13505,N_7084,N_8807);
xnor U13506 (N_13506,N_8255,N_7637);
xnor U13507 (N_13507,N_7848,N_9458);
nor U13508 (N_13508,N_7135,N_9208);
xnor U13509 (N_13509,N_8692,N_9520);
and U13510 (N_13510,N_11614,N_10651);
xnor U13511 (N_13511,N_7819,N_11790);
xnor U13512 (N_13512,N_10318,N_8878);
xor U13513 (N_13513,N_6779,N_10534);
and U13514 (N_13514,N_10264,N_9258);
or U13515 (N_13515,N_11944,N_11565);
nor U13516 (N_13516,N_11609,N_10722);
nor U13517 (N_13517,N_11300,N_12232);
nor U13518 (N_13518,N_10405,N_9786);
nand U13519 (N_13519,N_12331,N_9541);
and U13520 (N_13520,N_11713,N_11769);
and U13521 (N_13521,N_9984,N_8961);
nand U13522 (N_13522,N_10629,N_6438);
xnor U13523 (N_13523,N_8076,N_8117);
xor U13524 (N_13524,N_10126,N_8199);
nor U13525 (N_13525,N_11464,N_9210);
nand U13526 (N_13526,N_10659,N_11378);
nand U13527 (N_13527,N_11299,N_9283);
xnor U13528 (N_13528,N_8235,N_8905);
nor U13529 (N_13529,N_11002,N_8343);
nand U13530 (N_13530,N_8803,N_7918);
or U13531 (N_13531,N_12309,N_8859);
or U13532 (N_13532,N_11242,N_9923);
nand U13533 (N_13533,N_11892,N_11320);
nor U13534 (N_13534,N_6786,N_9538);
nor U13535 (N_13535,N_6922,N_7804);
or U13536 (N_13536,N_12122,N_10301);
nand U13537 (N_13537,N_9906,N_7573);
xor U13538 (N_13538,N_11214,N_6497);
and U13539 (N_13539,N_12352,N_7593);
xor U13540 (N_13540,N_8594,N_8721);
nor U13541 (N_13541,N_9560,N_7797);
and U13542 (N_13542,N_12494,N_10889);
and U13543 (N_13543,N_9762,N_11453);
and U13544 (N_13544,N_7869,N_9663);
nand U13545 (N_13545,N_8561,N_7115);
nor U13546 (N_13546,N_10112,N_9275);
nand U13547 (N_13547,N_12212,N_12439);
and U13548 (N_13548,N_10362,N_8395);
nand U13549 (N_13549,N_9768,N_9590);
nor U13550 (N_13550,N_7066,N_10098);
nand U13551 (N_13551,N_9524,N_12217);
or U13552 (N_13552,N_7628,N_12293);
and U13553 (N_13553,N_7601,N_7261);
and U13554 (N_13554,N_11024,N_11735);
or U13555 (N_13555,N_7109,N_7322);
nand U13556 (N_13556,N_7430,N_8429);
nor U13557 (N_13557,N_8053,N_11617);
xor U13558 (N_13558,N_9944,N_9633);
and U13559 (N_13559,N_10213,N_9189);
and U13560 (N_13560,N_10398,N_6740);
nand U13561 (N_13561,N_9263,N_11647);
or U13562 (N_13562,N_11520,N_8153);
nand U13563 (N_13563,N_12424,N_10386);
xnor U13564 (N_13564,N_11009,N_6748);
and U13565 (N_13565,N_9685,N_10896);
nand U13566 (N_13566,N_7963,N_11927);
xnor U13567 (N_13567,N_9948,N_8891);
or U13568 (N_13568,N_7641,N_8419);
nand U13569 (N_13569,N_6778,N_9169);
xnor U13570 (N_13570,N_6985,N_10399);
and U13571 (N_13571,N_11165,N_7949);
nor U13572 (N_13572,N_8701,N_9015);
xor U13573 (N_13573,N_9264,N_6476);
and U13574 (N_13574,N_6808,N_12358);
nand U13575 (N_13575,N_9031,N_11559);
and U13576 (N_13576,N_8999,N_10528);
and U13577 (N_13577,N_6616,N_9309);
nand U13578 (N_13578,N_6622,N_8357);
nand U13579 (N_13579,N_8192,N_6883);
and U13580 (N_13580,N_7113,N_11416);
xor U13581 (N_13581,N_8576,N_6569);
nand U13582 (N_13582,N_9993,N_7047);
nand U13583 (N_13583,N_11942,N_8737);
or U13584 (N_13584,N_11828,N_10159);
xor U13585 (N_13585,N_12221,N_6546);
xor U13586 (N_13586,N_7657,N_11350);
nand U13587 (N_13587,N_10007,N_11415);
nor U13588 (N_13588,N_9236,N_12165);
nor U13589 (N_13589,N_10708,N_8040);
or U13590 (N_13590,N_10288,N_9577);
nor U13591 (N_13591,N_7415,N_9584);
nor U13592 (N_13592,N_9864,N_6271);
and U13593 (N_13593,N_9914,N_6274);
or U13594 (N_13594,N_11978,N_11351);
nor U13595 (N_13595,N_10750,N_11545);
and U13596 (N_13596,N_10323,N_8866);
nor U13597 (N_13597,N_8595,N_6895);
nand U13598 (N_13598,N_11489,N_7031);
nor U13599 (N_13599,N_7295,N_10569);
or U13600 (N_13600,N_10791,N_7572);
or U13601 (N_13601,N_10718,N_9772);
xor U13602 (N_13602,N_6532,N_11883);
or U13603 (N_13603,N_10009,N_11133);
nand U13604 (N_13604,N_12321,N_11052);
nand U13605 (N_13605,N_10974,N_8344);
and U13606 (N_13606,N_9338,N_9927);
nand U13607 (N_13607,N_7034,N_8332);
and U13608 (N_13608,N_11517,N_6889);
and U13609 (N_13609,N_9384,N_7619);
and U13610 (N_13610,N_9098,N_12391);
or U13611 (N_13611,N_8611,N_10655);
and U13612 (N_13612,N_9061,N_8295);
or U13613 (N_13613,N_8997,N_12475);
xor U13614 (N_13614,N_7590,N_12096);
or U13615 (N_13615,N_10296,N_7578);
nand U13616 (N_13616,N_7845,N_11963);
and U13617 (N_13617,N_8051,N_12008);
xor U13618 (N_13618,N_8048,N_10820);
or U13619 (N_13619,N_9351,N_11196);
nor U13620 (N_13620,N_8830,N_8858);
nand U13621 (N_13621,N_12067,N_11180);
and U13622 (N_13622,N_11096,N_9120);
nand U13623 (N_13623,N_8105,N_6524);
nor U13624 (N_13624,N_11442,N_9759);
nor U13625 (N_13625,N_8716,N_8730);
and U13626 (N_13626,N_7478,N_8460);
nor U13627 (N_13627,N_7574,N_7234);
nand U13628 (N_13628,N_12229,N_12181);
nor U13629 (N_13629,N_11750,N_9969);
and U13630 (N_13630,N_10650,N_8809);
xor U13631 (N_13631,N_7696,N_11353);
or U13632 (N_13632,N_8569,N_6791);
or U13633 (N_13633,N_8995,N_7770);
nor U13634 (N_13634,N_11808,N_12311);
and U13635 (N_13635,N_12354,N_7999);
nor U13636 (N_13636,N_11918,N_10482);
and U13637 (N_13637,N_12249,N_12086);
and U13638 (N_13638,N_11304,N_7298);
nand U13639 (N_13639,N_9901,N_11793);
nor U13640 (N_13640,N_12121,N_7176);
nand U13641 (N_13641,N_7888,N_8096);
nand U13642 (N_13642,N_8173,N_9996);
xnor U13643 (N_13643,N_7233,N_9148);
or U13644 (N_13644,N_10885,N_8965);
nand U13645 (N_13645,N_11634,N_6720);
or U13646 (N_13646,N_7425,N_6766);
or U13647 (N_13647,N_6997,N_11687);
nand U13648 (N_13648,N_9042,N_12332);
and U13649 (N_13649,N_9849,N_9314);
and U13650 (N_13650,N_6792,N_12324);
xor U13651 (N_13651,N_12262,N_7369);
and U13652 (N_13652,N_7082,N_6587);
nand U13653 (N_13653,N_7608,N_12159);
nand U13654 (N_13654,N_7463,N_8128);
or U13655 (N_13655,N_7088,N_9327);
or U13656 (N_13656,N_12357,N_6551);
xnor U13657 (N_13657,N_6833,N_10926);
xnor U13658 (N_13658,N_7300,N_7252);
nand U13659 (N_13659,N_11345,N_11796);
nor U13660 (N_13660,N_8012,N_11692);
nor U13661 (N_13661,N_7440,N_7419);
or U13662 (N_13662,N_12029,N_8028);
or U13663 (N_13663,N_6877,N_8435);
xnor U13664 (N_13664,N_8198,N_12489);
nor U13665 (N_13665,N_10897,N_9569);
nand U13666 (N_13666,N_12214,N_10222);
nor U13667 (N_13667,N_8495,N_10193);
nand U13668 (N_13668,N_11976,N_8196);
nor U13669 (N_13669,N_12455,N_11235);
nor U13670 (N_13670,N_7579,N_6844);
nor U13671 (N_13671,N_9228,N_6852);
nor U13672 (N_13672,N_9405,N_11514);
and U13673 (N_13673,N_8926,N_11902);
and U13674 (N_13674,N_6376,N_11301);
xor U13675 (N_13675,N_10391,N_7870);
xnor U13676 (N_13676,N_8672,N_10055);
or U13677 (N_13677,N_11387,N_7183);
nand U13678 (N_13678,N_10526,N_12083);
nand U13679 (N_13679,N_9732,N_8589);
and U13680 (N_13680,N_12349,N_6646);
xnor U13681 (N_13681,N_8550,N_9818);
or U13682 (N_13682,N_7604,N_9909);
and U13683 (N_13683,N_10737,N_11915);
nand U13684 (N_13684,N_9477,N_7188);
nand U13685 (N_13685,N_8340,N_11912);
nand U13686 (N_13686,N_9835,N_6457);
or U13687 (N_13687,N_7778,N_7693);
nand U13688 (N_13688,N_6473,N_6884);
nand U13689 (N_13689,N_9495,N_7667);
and U13690 (N_13690,N_9268,N_9861);
or U13691 (N_13691,N_9686,N_7886);
nand U13692 (N_13692,N_6859,N_12138);
xor U13693 (N_13693,N_11810,N_12173);
or U13694 (N_13694,N_8671,N_8562);
nand U13695 (N_13695,N_9401,N_12062);
and U13696 (N_13696,N_7703,N_7624);
and U13697 (N_13697,N_10471,N_11368);
and U13698 (N_13698,N_7672,N_11611);
nand U13699 (N_13699,N_12047,N_6739);
nor U13700 (N_13700,N_6874,N_7380);
xnor U13701 (N_13701,N_11612,N_9857);
and U13702 (N_13702,N_7414,N_9121);
nor U13703 (N_13703,N_6362,N_10340);
nand U13704 (N_13704,N_11724,N_9380);
nor U13705 (N_13705,N_8354,N_11727);
nand U13706 (N_13706,N_6270,N_8679);
nand U13707 (N_13707,N_10921,N_11456);
or U13708 (N_13708,N_7142,N_11977);
xor U13709 (N_13709,N_12218,N_11454);
and U13710 (N_13710,N_7914,N_8061);
nand U13711 (N_13711,N_11588,N_11354);
nor U13712 (N_13712,N_8557,N_12422);
xor U13713 (N_13713,N_8298,N_8683);
nand U13714 (N_13714,N_10031,N_7935);
nand U13715 (N_13715,N_9427,N_7857);
nand U13716 (N_13716,N_6902,N_9824);
nand U13717 (N_13717,N_8971,N_10376);
nor U13718 (N_13718,N_7793,N_9085);
and U13719 (N_13719,N_6828,N_6625);
nor U13720 (N_13720,N_7459,N_10095);
xor U13721 (N_13721,N_7058,N_6375);
nand U13722 (N_13722,N_9504,N_10652);
and U13723 (N_13723,N_8563,N_9546);
nand U13724 (N_13724,N_8944,N_7610);
xnor U13725 (N_13725,N_10907,N_9734);
xor U13726 (N_13726,N_11576,N_8308);
xor U13727 (N_13727,N_9526,N_10438);
xor U13728 (N_13728,N_6420,N_8664);
and U13729 (N_13729,N_7565,N_11748);
and U13730 (N_13730,N_9830,N_6431);
nor U13731 (N_13731,N_12118,N_12431);
or U13732 (N_13732,N_10550,N_7577);
nor U13733 (N_13733,N_8936,N_10317);
nor U13734 (N_13734,N_9888,N_9345);
xnor U13735 (N_13735,N_12238,N_11904);
nor U13736 (N_13736,N_11982,N_11265);
or U13737 (N_13737,N_11789,N_10768);
and U13738 (N_13738,N_8892,N_9897);
or U13739 (N_13739,N_8022,N_7908);
or U13740 (N_13740,N_10546,N_10520);
nand U13741 (N_13741,N_11600,N_8071);
or U13742 (N_13742,N_12421,N_9074);
and U13743 (N_13743,N_7627,N_7557);
xor U13744 (N_13744,N_10469,N_7196);
nand U13745 (N_13745,N_10925,N_7099);
nor U13746 (N_13746,N_7503,N_11237);
nor U13747 (N_13747,N_9935,N_9139);
and U13748 (N_13748,N_8796,N_10899);
nand U13749 (N_13749,N_6956,N_8145);
nand U13750 (N_13750,N_7776,N_12020);
and U13751 (N_13751,N_9697,N_12104);
nand U13752 (N_13752,N_12070,N_9373);
or U13753 (N_13753,N_11621,N_8253);
nand U13754 (N_13754,N_10545,N_7891);
nor U13755 (N_13755,N_7592,N_7737);
xor U13756 (N_13756,N_10114,N_7652);
or U13757 (N_13757,N_9791,N_9415);
xor U13758 (N_13758,N_11308,N_7487);
and U13759 (N_13759,N_11759,N_6464);
or U13760 (N_13760,N_9265,N_9434);
nor U13761 (N_13761,N_7486,N_11784);
or U13762 (N_13762,N_6718,N_10551);
and U13763 (N_13763,N_11512,N_10898);
xor U13764 (N_13764,N_7823,N_9581);
nor U13765 (N_13765,N_9576,N_10427);
and U13766 (N_13766,N_8963,N_9570);
xor U13767 (N_13767,N_7723,N_11500);
nand U13768 (N_13768,N_9201,N_6325);
nand U13769 (N_13769,N_11861,N_7815);
xor U13770 (N_13770,N_6921,N_9037);
nor U13771 (N_13771,N_9214,N_6515);
nand U13772 (N_13772,N_11185,N_8297);
or U13773 (N_13773,N_7171,N_6839);
xnor U13774 (N_13774,N_9971,N_6409);
xor U13775 (N_13775,N_10178,N_9720);
xor U13776 (N_13776,N_8417,N_9291);
xnor U13777 (N_13777,N_10911,N_7141);
nor U13778 (N_13778,N_10133,N_8869);
xnor U13779 (N_13779,N_7094,N_7270);
xnor U13780 (N_13780,N_11696,N_11224);
or U13781 (N_13781,N_7181,N_11063);
nor U13782 (N_13782,N_9966,N_9682);
nand U13783 (N_13783,N_9133,N_10190);
or U13784 (N_13784,N_10933,N_8584);
or U13785 (N_13785,N_6677,N_7923);
xnor U13786 (N_13786,N_10097,N_7454);
and U13787 (N_13787,N_11592,N_7903);
xor U13788 (N_13788,N_7539,N_7938);
and U13789 (N_13789,N_10843,N_9525);
or U13790 (N_13790,N_8243,N_8917);
nor U13791 (N_13791,N_6521,N_6487);
nand U13792 (N_13792,N_6924,N_8152);
and U13793 (N_13793,N_9689,N_9846);
or U13794 (N_13794,N_8776,N_9209);
nor U13795 (N_13795,N_10522,N_12275);
xnor U13796 (N_13796,N_12353,N_11806);
nand U13797 (N_13797,N_6384,N_11201);
nor U13798 (N_13798,N_12430,N_7466);
nand U13799 (N_13799,N_8899,N_6835);
or U13800 (N_13800,N_12436,N_10980);
or U13801 (N_13801,N_10985,N_10660);
xor U13802 (N_13802,N_8718,N_9781);
or U13803 (N_13803,N_11684,N_11126);
nor U13804 (N_13804,N_6799,N_7551);
or U13805 (N_13805,N_8643,N_10388);
or U13806 (N_13806,N_9764,N_11983);
or U13807 (N_13807,N_10034,N_12359);
nor U13808 (N_13808,N_11811,N_7085);
xnor U13809 (N_13809,N_7106,N_8239);
or U13810 (N_13810,N_8209,N_10877);
xor U13811 (N_13811,N_8078,N_8765);
or U13812 (N_13812,N_9057,N_10205);
xor U13813 (N_13813,N_7866,N_7396);
and U13814 (N_13814,N_10165,N_10837);
nor U13815 (N_13815,N_8481,N_12362);
and U13816 (N_13816,N_11118,N_10535);
or U13817 (N_13817,N_12065,N_6351);
or U13818 (N_13818,N_7944,N_9747);
xor U13819 (N_13819,N_9995,N_10817);
and U13820 (N_13820,N_9688,N_9411);
xor U13821 (N_13821,N_12387,N_6395);
xor U13822 (N_13822,N_11160,N_7831);
nor U13823 (N_13823,N_12068,N_9054);
or U13824 (N_13824,N_9164,N_9090);
or U13825 (N_13825,N_11557,N_9507);
nor U13826 (N_13826,N_8443,N_10617);
nor U13827 (N_13827,N_7222,N_9882);
xnor U13828 (N_13828,N_6823,N_11236);
and U13829 (N_13829,N_11032,N_12336);
or U13830 (N_13830,N_6746,N_11098);
and U13831 (N_13831,N_11465,N_12048);
and U13832 (N_13832,N_8011,N_9192);
nand U13833 (N_13833,N_8165,N_8296);
nor U13834 (N_13834,N_11127,N_8439);
nand U13835 (N_13835,N_9191,N_11226);
nor U13836 (N_13836,N_6483,N_7191);
xnor U13837 (N_13837,N_9231,N_6364);
nor U13838 (N_13838,N_12103,N_7398);
or U13839 (N_13839,N_11005,N_11920);
or U13840 (N_13840,N_11524,N_7631);
nor U13841 (N_13841,N_8428,N_10220);
nor U13842 (N_13842,N_8097,N_12280);
nor U13843 (N_13843,N_6683,N_6573);
xnor U13844 (N_13844,N_10235,N_9597);
xnor U13845 (N_13845,N_12302,N_11047);
nand U13846 (N_13846,N_6342,N_11827);
nand U13847 (N_13847,N_8665,N_6934);
xnor U13848 (N_13848,N_9330,N_9805);
nor U13849 (N_13849,N_9255,N_8833);
nand U13850 (N_13850,N_11358,N_9007);
xor U13851 (N_13851,N_10253,N_7526);
xor U13852 (N_13852,N_9908,N_10703);
or U13853 (N_13853,N_9532,N_8533);
nor U13854 (N_13854,N_7644,N_8400);
nor U13855 (N_13855,N_6529,N_7632);
xor U13856 (N_13856,N_10716,N_6809);
or U13857 (N_13857,N_6556,N_11649);
xnor U13858 (N_13858,N_8376,N_9692);
or U13859 (N_13859,N_12235,N_7383);
and U13860 (N_13860,N_10185,N_8368);
nor U13861 (N_13861,N_10966,N_7269);
xnor U13862 (N_13862,N_9879,N_9754);
xor U13863 (N_13863,N_11767,N_6875);
and U13864 (N_13864,N_7016,N_9343);
or U13865 (N_13865,N_8277,N_7799);
and U13866 (N_13866,N_11615,N_8600);
or U13867 (N_13867,N_9858,N_6906);
or U13868 (N_13868,N_6503,N_10139);
or U13869 (N_13869,N_9254,N_7818);
or U13870 (N_13870,N_11975,N_11865);
and U13871 (N_13871,N_11766,N_9585);
or U13872 (N_13872,N_11858,N_12460);
and U13873 (N_13873,N_11225,N_7381);
nand U13874 (N_13874,N_7926,N_11441);
xor U13875 (N_13875,N_7144,N_12046);
xnor U13876 (N_13876,N_6414,N_6723);
nor U13877 (N_13877,N_8856,N_7453);
or U13878 (N_13878,N_9465,N_9939);
xnor U13879 (N_13879,N_7306,N_6328);
and U13880 (N_13880,N_10946,N_8032);
and U13881 (N_13881,N_12042,N_9671);
xor U13882 (N_13882,N_10774,N_6520);
xnor U13883 (N_13883,N_7485,N_8143);
nor U13884 (N_13884,N_12097,N_7101);
nor U13885 (N_13885,N_9921,N_12143);
and U13886 (N_13886,N_6519,N_7549);
or U13887 (N_13887,N_10204,N_12312);
nand U13888 (N_13888,N_11395,N_7469);
nor U13889 (N_13889,N_10807,N_7205);
or U13890 (N_13890,N_8873,N_6273);
and U13891 (N_13891,N_8614,N_11913);
and U13892 (N_13892,N_8727,N_6662);
or U13893 (N_13893,N_6444,N_8666);
nor U13894 (N_13894,N_11672,N_10328);
nor U13895 (N_13895,N_8364,N_7096);
and U13896 (N_13896,N_8224,N_12200);
and U13897 (N_13897,N_6612,N_10834);
nand U13898 (N_13898,N_6338,N_9820);
nor U13899 (N_13899,N_10908,N_6814);
or U13900 (N_13900,N_8106,N_12215);
nor U13901 (N_13901,N_11578,N_7955);
and U13902 (N_13902,N_7710,N_7212);
xor U13903 (N_13903,N_11315,N_7189);
xor U13904 (N_13904,N_10446,N_9076);
xnor U13905 (N_13905,N_6621,N_7792);
nor U13906 (N_13906,N_10223,N_6461);
xnor U13907 (N_13907,N_10196,N_9558);
nor U13908 (N_13908,N_7400,N_10061);
nand U13909 (N_13909,N_11470,N_11365);
nand U13910 (N_13910,N_9117,N_9641);
nor U13911 (N_13911,N_6509,N_12345);
nor U13912 (N_13912,N_7858,N_9769);
xnor U13913 (N_13913,N_8893,N_9647);
or U13914 (N_13914,N_7490,N_10115);
and U13915 (N_13915,N_7207,N_6567);
and U13916 (N_13916,N_9701,N_7428);
and U13917 (N_13917,N_9205,N_7732);
nand U13918 (N_13918,N_12346,N_8923);
or U13919 (N_13919,N_6534,N_11083);
xnor U13920 (N_13920,N_12300,N_7759);
xnor U13921 (N_13921,N_10077,N_11554);
xor U13922 (N_13922,N_11764,N_9393);
or U13923 (N_13923,N_6972,N_10648);
nand U13924 (N_13924,N_10403,N_12456);
and U13925 (N_13925,N_8501,N_7173);
xnor U13926 (N_13926,N_12486,N_9549);
nand U13927 (N_13927,N_8935,N_12004);
xor U13928 (N_13928,N_11900,N_7023);
nor U13929 (N_13929,N_10181,N_8322);
xnor U13930 (N_13930,N_6671,N_10810);
and U13931 (N_13931,N_11317,N_7157);
xor U13932 (N_13932,N_7929,N_8367);
and U13933 (N_13933,N_7585,N_10917);
or U13934 (N_13934,N_10255,N_7015);
nand U13935 (N_13935,N_8110,N_8432);
nand U13936 (N_13936,N_10874,N_11974);
and U13937 (N_13937,N_11195,N_11909);
nand U13938 (N_13938,N_8150,N_6942);
xor U13939 (N_13939,N_6707,N_12314);
or U13940 (N_13940,N_12405,N_9433);
and U13941 (N_13941,N_7456,N_7760);
nand U13942 (N_13942,N_9602,N_10184);
nor U13943 (N_13943,N_7350,N_11771);
nor U13944 (N_13944,N_9973,N_10507);
and U13945 (N_13945,N_8163,N_10637);
or U13946 (N_13946,N_7885,N_12388);
and U13947 (N_13947,N_8876,N_8402);
or U13948 (N_13948,N_10714,N_9025);
xnor U13949 (N_13949,N_11244,N_11657);
nand U13950 (N_13950,N_12329,N_10867);
and U13951 (N_13951,N_9337,N_7586);
and U13952 (N_13952,N_7936,N_7900);
xnor U13953 (N_13953,N_10423,N_10855);
nand U13954 (N_13954,N_11364,N_7475);
and U13955 (N_13955,N_10540,N_11075);
or U13956 (N_13956,N_10262,N_9547);
nor U13957 (N_13957,N_11136,N_6953);
xnor U13958 (N_13958,N_7794,N_12147);
nand U13959 (N_13959,N_9027,N_8323);
or U13960 (N_13960,N_12361,N_11095);
nor U13961 (N_13961,N_9953,N_10746);
xnor U13962 (N_13962,N_8015,N_9213);
or U13963 (N_13963,N_8098,N_8821);
xnor U13964 (N_13964,N_10454,N_12239);
xnor U13965 (N_13965,N_11589,N_11496);
and U13966 (N_13966,N_11417,N_12179);
and U13967 (N_13967,N_9534,N_11590);
or U13968 (N_13968,N_12064,N_7685);
xnor U13969 (N_13969,N_10876,N_10785);
xnor U13970 (N_13970,N_9543,N_8318);
or U13971 (N_13971,N_7392,N_11480);
nand U13972 (N_13972,N_11245,N_11804);
xor U13973 (N_13973,N_8274,N_6753);
or U13974 (N_13974,N_6299,N_10900);
nor U13975 (N_13975,N_12174,N_6550);
and U13976 (N_13976,N_7442,N_10498);
nor U13977 (N_13977,N_7330,N_10788);
nor U13978 (N_13978,N_6613,N_6572);
and U13979 (N_13979,N_9221,N_12295);
xor U13980 (N_13980,N_11862,N_8820);
and U13981 (N_13981,N_12171,N_6742);
nand U13982 (N_13982,N_8307,N_10151);
and U13983 (N_13983,N_7796,N_6878);
nor U13984 (N_13984,N_8319,N_7649);
nor U13985 (N_13985,N_12146,N_6845);
or U13986 (N_13986,N_6531,N_9439);
nand U13987 (N_13987,N_10229,N_12307);
and U13988 (N_13988,N_11012,N_11605);
xnor U13989 (N_13989,N_8121,N_11923);
or U13990 (N_13990,N_7417,N_7434);
and U13991 (N_13991,N_7209,N_6276);
or U13992 (N_13992,N_7509,N_7019);
nor U13993 (N_13993,N_10371,N_9287);
nor U13994 (N_13994,N_7881,N_9026);
nor U13995 (N_13995,N_11664,N_11555);
or U13996 (N_13996,N_10221,N_8331);
nor U13997 (N_13997,N_9981,N_11946);
nor U13998 (N_13998,N_8779,N_10451);
nor U13999 (N_13999,N_12263,N_10377);
or U14000 (N_14000,N_10269,N_11939);
and U14001 (N_14001,N_10004,N_10699);
or U14002 (N_14002,N_8523,N_9363);
and U14003 (N_14003,N_10073,N_9610);
nand U14004 (N_14004,N_8621,N_8258);
nand U14005 (N_14005,N_8160,N_11949);
or U14006 (N_14006,N_12228,N_6445);
nor U14007 (N_14007,N_10231,N_7412);
nor U14008 (N_14008,N_7856,N_9035);
and U14009 (N_14009,N_8176,N_8570);
and U14010 (N_14010,N_8369,N_10350);
xor U14011 (N_14011,N_6793,N_12281);
or U14012 (N_14012,N_10203,N_9478);
xor U14013 (N_14013,N_12085,N_10725);
and U14014 (N_14014,N_11173,N_6803);
nor U14015 (N_14015,N_10334,N_7014);
nand U14016 (N_14016,N_7482,N_11941);
xnor U14017 (N_14017,N_11298,N_10710);
nand U14018 (N_14018,N_11740,N_12196);
nor U14019 (N_14019,N_6907,N_11544);
nor U14020 (N_14020,N_9982,N_10465);
nor U14021 (N_14021,N_11553,N_10475);
and U14022 (N_14022,N_7660,N_7984);
nand U14023 (N_14023,N_8141,N_9332);
or U14024 (N_14024,N_7324,N_10794);
and U14025 (N_14025,N_6651,N_10243);
nand U14026 (N_14026,N_8558,N_7122);
nor U14027 (N_14027,N_7614,N_6336);
or U14028 (N_14028,N_12037,N_9141);
xor U14029 (N_14029,N_6477,N_8119);
xor U14030 (N_14030,N_6557,N_7525);
nand U14031 (N_14031,N_8401,N_10518);
or U14032 (N_14032,N_7249,N_11276);
or U14033 (N_14033,N_6825,N_6933);
nand U14034 (N_14034,N_7030,N_10560);
xnor U14035 (N_14035,N_7746,N_10389);
and U14036 (N_14036,N_10923,N_11842);
or U14037 (N_14037,N_7070,N_9614);
and U14038 (N_14038,N_10428,N_7489);
and U14039 (N_14039,N_8338,N_9013);
nand U14040 (N_14040,N_6960,N_10833);
nand U14041 (N_14041,N_8293,N_11625);
and U14042 (N_14042,N_7560,N_9733);
xnor U14043 (N_14043,N_10719,N_7718);
nor U14044 (N_14044,N_8290,N_9385);
xor U14045 (N_14045,N_12370,N_6394);
or U14046 (N_14046,N_7616,N_9193);
nor U14047 (N_14047,N_10217,N_9470);
nand U14048 (N_14048,N_9776,N_8653);
xnor U14049 (N_14049,N_10265,N_9162);
nand U14050 (N_14050,N_9537,N_8240);
nor U14051 (N_14051,N_9294,N_6450);
nand U14052 (N_14052,N_6635,N_6535);
xor U14053 (N_14053,N_9217,N_11197);
or U14054 (N_14054,N_10691,N_8810);
xor U14055 (N_14055,N_7980,N_8329);
nand U14056 (N_14056,N_11426,N_11346);
nand U14057 (N_14057,N_12380,N_10605);
or U14058 (N_14058,N_8839,N_12176);
or U14059 (N_14059,N_8906,N_8268);
nand U14060 (N_14060,N_7665,N_7050);
xnor U14061 (N_14061,N_8627,N_11138);
xnor U14062 (N_14062,N_12023,N_10382);
xnor U14063 (N_14063,N_6512,N_9722);
nor U14064 (N_14064,N_7814,N_6356);
nor U14065 (N_14065,N_7754,N_9785);
nand U14066 (N_14066,N_12457,N_9796);
xor U14067 (N_14067,N_6598,N_9046);
xor U14068 (N_14068,N_11730,N_9333);
and U14069 (N_14069,N_8377,N_10544);
nand U14070 (N_14070,N_10194,N_12257);
nor U14071 (N_14071,N_12170,N_6920);
or U14072 (N_14072,N_6455,N_8464);
nand U14073 (N_14073,N_8885,N_7789);
nand U14074 (N_14074,N_8414,N_7842);
or U14075 (N_14075,N_11303,N_10360);
nor U14076 (N_14076,N_6947,N_6525);
nand U14077 (N_14077,N_9047,N_9211);
nand U14078 (N_14078,N_8559,N_11930);
nand U14079 (N_14079,N_7411,N_6608);
or U14080 (N_14080,N_9497,N_6410);
xor U14081 (N_14081,N_10623,N_10901);
and U14082 (N_14082,N_10276,N_8264);
or U14083 (N_14083,N_9018,N_10961);
nor U14084 (N_14084,N_12438,N_12195);
nand U14085 (N_14085,N_11598,N_10473);
nor U14086 (N_14086,N_10916,N_11655);
and U14087 (N_14087,N_11250,N_7397);
or U14088 (N_14088,N_12491,N_7706);
nor U14089 (N_14089,N_9660,N_7830);
and U14090 (N_14090,N_11377,N_11616);
or U14091 (N_14091,N_12451,N_8113);
nor U14092 (N_14092,N_10163,N_9190);
or U14093 (N_14093,N_7953,N_6810);
and U14094 (N_14094,N_11331,N_9303);
nand U14095 (N_14095,N_7348,N_10944);
or U14096 (N_14096,N_8663,N_11405);
xnor U14097 (N_14097,N_9084,N_9990);
and U14098 (N_14098,N_9743,N_11905);
or U14099 (N_14099,N_12449,N_8333);
or U14100 (N_14100,N_6943,N_10250);
xnor U14101 (N_14101,N_11155,N_9809);
and U14102 (N_14102,N_11871,N_7775);
xnor U14103 (N_14103,N_6310,N_11144);
nor U14104 (N_14104,N_7177,N_9767);
nor U14105 (N_14105,N_10850,N_7939);
nor U14106 (N_14106,N_8366,N_12031);
and U14107 (N_14107,N_11971,N_8922);
xor U14108 (N_14108,N_7092,N_10851);
nand U14109 (N_14109,N_11289,N_8610);
xor U14110 (N_14110,N_11897,N_6334);
and U14111 (N_14111,N_6432,N_11761);
xnor U14112 (N_14112,N_11107,N_7989);
and U14113 (N_14113,N_10153,N_9297);
nor U14114 (N_14114,N_10150,N_10533);
nand U14115 (N_14115,N_9716,N_7134);
and U14116 (N_14116,N_8933,N_9030);
and U14117 (N_14117,N_7206,N_7378);
nor U14118 (N_14118,N_10607,N_11830);
xnor U14119 (N_14119,N_9683,N_6494);
and U14120 (N_14120,N_7168,N_10005);
nand U14121 (N_14121,N_12052,N_8313);
xnor U14122 (N_14122,N_11916,N_7049);
nor U14123 (N_14123,N_7554,N_6527);
nand U14124 (N_14124,N_8731,N_6987);
nand U14125 (N_14125,N_11685,N_12245);
nand U14126 (N_14126,N_8473,N_10996);
nor U14127 (N_14127,N_6601,N_8189);
or U14128 (N_14128,N_9775,N_10020);
nor U14129 (N_14129,N_9724,N_9267);
and U14130 (N_14130,N_12234,N_9111);
or U14131 (N_14131,N_11291,N_10160);
and U14132 (N_14132,N_7232,N_8868);
xor U14133 (N_14133,N_6888,N_12406);
xor U14134 (N_14134,N_7204,N_10494);
nand U14135 (N_14135,N_6602,N_7032);
nand U14136 (N_14136,N_7567,N_11116);
and U14137 (N_14137,N_9587,N_11836);
or U14138 (N_14138,N_6674,N_10939);
xor U14139 (N_14139,N_12320,N_11177);
and U14140 (N_14140,N_7907,N_8309);
xnor U14141 (N_14141,N_6579,N_9826);
nand U14142 (N_14142,N_11319,N_9392);
or U14143 (N_14143,N_11254,N_10056);
xor U14144 (N_14144,N_11349,N_10381);
and U14145 (N_14145,N_11817,N_10634);
or U14146 (N_14146,N_6939,N_8903);
xor U14147 (N_14147,N_9077,N_12480);
xor U14148 (N_14148,N_12175,N_8476);
nand U14149 (N_14149,N_11283,N_7426);
nand U14150 (N_14150,N_10890,N_7542);
nor U14151 (N_14151,N_9358,N_8070);
xor U14152 (N_14152,N_11938,N_11760);
and U14153 (N_14153,N_7820,N_10770);
nor U14154 (N_14154,N_8844,N_10694);
nor U14155 (N_14155,N_11396,N_11332);
or U14156 (N_14156,N_9204,N_10326);
xnor U14157 (N_14157,N_11309,N_12327);
xnor U14158 (N_14158,N_7236,N_8288);
nand U14159 (N_14159,N_9821,N_10780);
xor U14160 (N_14160,N_9548,N_10653);
xnor U14161 (N_14161,N_8499,N_6584);
xor U14162 (N_14162,N_10536,N_8411);
and U14163 (N_14163,N_10285,N_12201);
nand U14164 (N_14164,N_6419,N_7915);
xnor U14165 (N_14165,N_7740,N_7540);
nor U14166 (N_14166,N_7163,N_10720);
xor U14167 (N_14167,N_7444,N_10832);
xnor U14168 (N_14168,N_8532,N_11626);
xnor U14169 (N_14169,N_7670,N_10701);
or U14170 (N_14170,N_10057,N_10766);
nor U14171 (N_14171,N_7713,N_11488);
nand U14172 (N_14172,N_6722,N_7773);
or U14173 (N_14173,N_6629,N_6882);
or U14174 (N_14174,N_7506,N_8424);
nand U14175 (N_14175,N_7193,N_8359);
nand U14176 (N_14176,N_12408,N_9502);
and U14177 (N_14177,N_9055,N_7675);
nand U14178 (N_14178,N_11023,N_8427);
and U14179 (N_14179,N_10935,N_10392);
nand U14180 (N_14180,N_6826,N_8787);
nor U14181 (N_14181,N_10314,N_12461);
nand U14182 (N_14182,N_6435,N_6588);
nand U14183 (N_14183,N_9609,N_8118);
xor U14184 (N_14184,N_10826,N_9234);
nor U14185 (N_14185,N_6708,N_6747);
xor U14186 (N_14186,N_6836,N_12127);
and U14187 (N_14187,N_6504,N_8278);
nor U14188 (N_14188,N_7772,N_11307);
xnor U14189 (N_14189,N_9998,N_10924);
xor U14190 (N_14190,N_9398,N_6930);
xnor U14191 (N_14191,N_8548,N_6641);
and U14192 (N_14192,N_10124,N_11306);
nand U14193 (N_14193,N_7960,N_6491);
and U14194 (N_14194,N_9362,N_10143);
nor U14195 (N_14195,N_10669,N_8042);
or U14196 (N_14196,N_9501,N_8371);
nor U14197 (N_14197,N_10805,N_7441);
and U14198 (N_14198,N_7075,N_10579);
nor U14199 (N_14199,N_12313,N_12233);
or U14200 (N_14200,N_10563,N_11044);
nand U14201 (N_14201,N_11189,N_9875);
nand U14202 (N_14202,N_11513,N_10485);
and U14203 (N_14203,N_8125,N_7046);
nand U14204 (N_14204,N_8842,N_7867);
nand U14205 (N_14205,N_9230,N_8546);
nor U14206 (N_14206,N_10656,N_9202);
and U14207 (N_14207,N_6383,N_9130);
xnor U14208 (N_14208,N_11145,N_9041);
xnor U14209 (N_14209,N_7422,N_9110);
nand U14210 (N_14210,N_9594,N_8976);
nor U14211 (N_14211,N_6316,N_11255);
nor U14212 (N_14212,N_6736,N_6689);
nand U14213 (N_14213,N_8134,N_7361);
nor U14214 (N_14214,N_12240,N_11603);
or U14215 (N_14215,N_11527,N_11178);
xor U14216 (N_14216,N_6768,N_11758);
or U14217 (N_14217,N_8023,N_8327);
nand U14218 (N_14218,N_10749,N_6543);
nor U14219 (N_14219,N_7544,N_11190);
or U14220 (N_14220,N_7527,N_7187);
and U14221 (N_14221,N_10661,N_7118);
or U14222 (N_14222,N_8940,N_10110);
nor U14223 (N_14223,N_11092,N_6292);
xnor U14224 (N_14224,N_11181,N_9898);
and U14225 (N_14225,N_12088,N_10556);
and U14226 (N_14226,N_6640,N_7562);
and U14227 (N_14227,N_8009,N_9887);
xor U14228 (N_14228,N_7563,N_11414);
nor U14229 (N_14229,N_12024,N_11693);
and U14230 (N_14230,N_9408,N_11081);
or U14231 (N_14231,N_9493,N_6880);
nor U14232 (N_14232,N_10207,N_12355);
or U14233 (N_14233,N_7777,N_9812);
nor U14234 (N_14234,N_6919,N_8952);
nor U14235 (N_14235,N_10022,N_10878);
nor U14236 (N_14236,N_10013,N_11917);
nor U14237 (N_14237,N_12189,N_10904);
nand U14238 (N_14238,N_7536,N_7664);
xnor U14239 (N_14239,N_8375,N_9739);
and U14240 (N_14240,N_7645,N_12340);
or U14241 (N_14241,N_8835,N_9819);
xor U14242 (N_14242,N_6774,N_8356);
xnor U14243 (N_14243,N_8677,N_6717);
and U14244 (N_14244,N_7394,N_10801);
xor U14245 (N_14245,N_10858,N_9269);
nor U14246 (N_14246,N_11141,N_9967);
nand U14247 (N_14247,N_9292,N_10134);
and U14248 (N_14248,N_9006,N_7429);
nor U14249 (N_14249,N_10478,N_6327);
and U14250 (N_14250,N_11409,N_8228);
or U14251 (N_14251,N_8813,N_9902);
and U14252 (N_14252,N_9400,N_7558);
nor U14253 (N_14253,N_10273,N_6984);
nor U14254 (N_14254,N_10903,N_8087);
nand U14255 (N_14255,N_7243,N_9388);
xor U14256 (N_14256,N_10881,N_10587);
or U14257 (N_14257,N_6282,N_11756);
xnor U14258 (N_14258,N_6442,N_8182);
and U14259 (N_14259,N_10432,N_10028);
nor U14260 (N_14260,N_7638,N_8488);
or U14261 (N_14261,N_7941,N_11481);
nand U14262 (N_14262,N_10313,N_12045);
and U14263 (N_14263,N_8673,N_10209);
xor U14264 (N_14264,N_8219,N_11537);
nor U14265 (N_14265,N_11184,N_9905);
nand U14266 (N_14266,N_6363,N_7906);
or U14267 (N_14267,N_10177,N_8622);
nand U14268 (N_14268,N_12094,N_11709);
nand U14269 (N_14269,N_11697,N_9510);
xor U14270 (N_14270,N_10421,N_12154);
nand U14271 (N_14271,N_10418,N_11887);
nor U14272 (N_14272,N_11312,N_8075);
nor U14273 (N_14273,N_11534,N_12054);
or U14274 (N_14274,N_10846,N_12296);
nor U14275 (N_14275,N_10155,N_6495);
or U14276 (N_14276,N_6536,N_7292);
xnor U14277 (N_14277,N_7040,N_11427);
xor U14278 (N_14278,N_7704,N_8479);
nand U14279 (N_14279,N_8341,N_11878);
nand U14280 (N_14280,N_9752,N_8509);
nand U14281 (N_14281,N_9128,N_9938);
xor U14282 (N_14282,N_8334,N_7119);
xnor U14283 (N_14283,N_10487,N_9452);
and U14284 (N_14284,N_11484,N_10895);
and U14285 (N_14285,N_8092,N_10084);
nor U14286 (N_14286,N_9484,N_6370);
and U14287 (N_14287,N_7334,N_8669);
and U14288 (N_14288,N_8951,N_8857);
nor U14289 (N_14289,N_9698,N_11743);
nor U14290 (N_14290,N_12128,N_6716);
nor U14291 (N_14291,N_9365,N_8577);
nand U14292 (N_14292,N_7595,N_10215);
nand U14293 (N_14293,N_7828,N_10517);
xor U14294 (N_14294,N_7438,N_9360);
nor U14295 (N_14295,N_7946,N_10909);
nor U14296 (N_14296,N_7203,N_7195);
nand U14297 (N_14297,N_11028,N_11943);
and U14298 (N_14298,N_7656,N_9421);
or U14299 (N_14299,N_9838,N_10468);
nand U14300 (N_14300,N_10131,N_10297);
nor U14301 (N_14301,N_6577,N_10953);
or U14302 (N_14302,N_10087,N_7060);
nor U14303 (N_14303,N_7837,N_11925);
nor U14304 (N_14304,N_11794,N_9448);
and U14305 (N_14305,N_7612,N_7964);
nor U14306 (N_14306,N_8829,N_9382);
and U14307 (N_14307,N_9872,N_11460);
nor U14308 (N_14308,N_11987,N_11548);
and U14309 (N_14309,N_11154,N_8640);
or U14310 (N_14310,N_8303,N_10435);
or U14311 (N_14311,N_7079,N_9108);
and U14312 (N_14312,N_10321,N_7894);
and U14313 (N_14313,N_7896,N_8618);
nand U14314 (N_14314,N_11230,N_11437);
nor U14315 (N_14315,N_10082,N_10951);
nand U14316 (N_14316,N_10047,N_7800);
and U14317 (N_14317,N_12458,N_11182);
xor U14318 (N_14318,N_6448,N_8461);
and U14319 (N_14319,N_12184,N_8492);
or U14320 (N_14320,N_11478,N_9489);
nand U14321 (N_14321,N_9896,N_9252);
nand U14322 (N_14322,N_10977,N_7838);
nor U14323 (N_14323,N_8300,N_12416);
or U14324 (N_14324,N_9512,N_6980);
and U14325 (N_14325,N_11690,N_8920);
or U14326 (N_14326,N_7501,N_8583);
nand U14327 (N_14327,N_7954,N_7114);
or U14328 (N_14328,N_10502,N_11741);
nand U14329 (N_14329,N_7666,N_6898);
nand U14330 (N_14330,N_7695,N_8538);
nor U14331 (N_14331,N_11232,N_8167);
or U14332 (N_14332,N_7990,N_8477);
nand U14333 (N_14333,N_6831,N_8230);
and U14334 (N_14334,N_12291,N_10452);
and U14335 (N_14335,N_11310,N_8321);
xor U14336 (N_14336,N_12027,N_11768);
xor U14337 (N_14337,N_8749,N_7669);
or U14338 (N_14338,N_7449,N_7994);
xnor U14339 (N_14339,N_9779,N_11105);
xor U14340 (N_14340,N_9347,N_9364);
or U14341 (N_14341,N_10687,N_11591);
nor U14342 (N_14342,N_9565,N_12140);
nand U14343 (N_14343,N_6842,N_9240);
nor U14344 (N_14344,N_10937,N_9955);
and U14345 (N_14345,N_10991,N_8947);
xor U14346 (N_14346,N_7757,N_7561);
and U14347 (N_14347,N_10284,N_7893);
or U14348 (N_14348,N_10107,N_11566);
xnor U14349 (N_14349,N_10599,N_9323);
nor U14350 (N_14350,N_9676,N_9199);
nand U14351 (N_14351,N_8037,N_9247);
nand U14352 (N_14352,N_10914,N_9886);
xnor U14353 (N_14353,N_9469,N_11286);
nand U14354 (N_14354,N_8756,N_12301);
xnor U14355 (N_14355,N_10697,N_8272);
or U14356 (N_14356,N_9924,N_12259);
or U14357 (N_14357,N_11376,N_11203);
and U14358 (N_14358,N_9653,N_10945);
nand U14359 (N_14359,N_7897,N_6265);
and U14360 (N_14360,N_7780,N_10078);
xnor U14361 (N_14361,N_7336,N_11097);
nand U14362 (N_14362,N_10705,N_7829);
xor U14363 (N_14363,N_11228,N_7159);
and U14364 (N_14364,N_10349,N_6252);
or U14365 (N_14365,N_6881,N_9646);
and U14366 (N_14366,N_12075,N_7045);
nand U14367 (N_14367,N_9353,N_10611);
xor U14368 (N_14368,N_9099,N_6425);
and U14369 (N_14369,N_7305,N_11646);
nor U14370 (N_14370,N_11448,N_9088);
and U14371 (N_14371,N_8848,N_9719);
and U14372 (N_14372,N_12155,N_6725);
nand U14373 (N_14373,N_9083,N_11989);
and U14374 (N_14374,N_8127,N_7024);
and U14375 (N_14375,N_10001,N_9301);
xor U14376 (N_14376,N_8860,N_9096);
nand U14377 (N_14377,N_10940,N_10148);
nor U14378 (N_14378,N_10106,N_8034);
xor U14379 (N_14379,N_10844,N_7991);
nand U14380 (N_14380,N_9067,N_8216);
nand U14381 (N_14381,N_8054,N_11139);
nand U14382 (N_14382,N_8740,N_11213);
nor U14383 (N_14383,N_11357,N_12397);
nand U14384 (N_14384,N_7979,N_7985);
nand U14385 (N_14385,N_11234,N_9105);
or U14386 (N_14386,N_10330,N_7663);
nor U14387 (N_14387,N_11679,N_7186);
nor U14388 (N_14388,N_8988,N_6405);
nand U14389 (N_14389,N_6938,N_8452);
xnor U14390 (N_14390,N_6918,N_9203);
xor U14391 (N_14391,N_7480,N_9259);
or U14392 (N_14392,N_6653,N_7839);
xor U14393 (N_14393,N_8580,N_11209);
or U14394 (N_14394,N_9575,N_7139);
nor U14395 (N_14395,N_8573,N_10375);
nand U14396 (N_14396,N_6514,N_7132);
and U14397 (N_14397,N_11507,N_10758);
and U14398 (N_14398,N_10429,N_11045);
nor U14399 (N_14399,N_10481,N_12426);
nand U14400 (N_14400,N_11084,N_8448);
xnor U14401 (N_14401,N_11599,N_11191);
nand U14402 (N_14402,N_6871,N_12481);
nand U14403 (N_14403,N_7432,N_8292);
nor U14404 (N_14404,N_7229,N_8232);
xnor U14405 (N_14405,N_7403,N_9892);
nor U14406 (N_14406,N_8723,N_10496);
or U14407 (N_14407,N_9109,N_11610);
nor U14408 (N_14408,N_9416,N_12194);
or U14409 (N_14409,N_7117,N_10467);
or U14410 (N_14410,N_6570,N_9674);
xnor U14411 (N_14411,N_9748,N_11435);
or U14412 (N_14412,N_6407,N_8244);
xor U14413 (N_14413,N_10132,N_10140);
nor U14414 (N_14414,N_11710,N_7587);
nor U14415 (N_14415,N_9666,N_6306);
or U14416 (N_14416,N_11115,N_6581);
and U14417 (N_14417,N_6630,N_12399);
nor U14418 (N_14418,N_8927,N_12476);
xnor U14419 (N_14419,N_11305,N_11874);
or U14420 (N_14420,N_10657,N_10280);
or U14421 (N_14421,N_11370,N_11328);
nor U14422 (N_14422,N_8535,N_12258);
nand U14423 (N_14423,N_7607,N_9381);
or U14424 (N_14424,N_12117,N_8470);
nand U14425 (N_14425,N_10525,N_10915);
nor U14426 (N_14426,N_7932,N_8155);
xor U14427 (N_14427,N_11894,N_7199);
and U14428 (N_14428,N_6470,N_11108);
or U14429 (N_14429,N_11137,N_6773);
or U14430 (N_14430,N_11985,N_12108);
and U14431 (N_14431,N_9064,N_12057);
or U14432 (N_14432,N_6475,N_9593);
nor U14433 (N_14433,N_10000,N_9974);
nand U14434 (N_14434,N_8853,N_12063);
xnor U14435 (N_14435,N_9424,N_10242);
xnor U14436 (N_14436,N_7265,N_12420);
nand U14437 (N_14437,N_10919,N_11780);
or U14438 (N_14438,N_12268,N_8620);
and U14439 (N_14439,N_6965,N_10192);
and U14440 (N_14440,N_7367,N_10721);
or U14441 (N_14441,N_11541,N_8804);
nand U14442 (N_14442,N_7568,N_10011);
xnor U14443 (N_14443,N_7078,N_8782);
and U14444 (N_14444,N_8335,N_7972);
or U14445 (N_14445,N_12186,N_10311);
nand U14446 (N_14446,N_11356,N_10767);
and U14447 (N_14447,N_6732,N_11652);
or U14448 (N_14448,N_10406,N_9986);
nand U14449 (N_14449,N_11412,N_12192);
or U14450 (N_14450,N_7643,N_7786);
and U14451 (N_14451,N_9249,N_10103);
nand U14452 (N_14452,N_7197,N_10397);
or U14453 (N_14453,N_8129,N_8468);
xor U14454 (N_14454,N_8567,N_10306);
nor U14455 (N_14455,N_8814,N_6704);
nand U14456 (N_14456,N_7847,N_11381);
or U14457 (N_14457,N_7743,N_6728);
or U14458 (N_14458,N_9947,N_6821);
and U14459 (N_14459,N_10322,N_6684);
and U14460 (N_14460,N_6686,N_7410);
or U14461 (N_14461,N_11875,N_7121);
nor U14462 (N_14462,N_8430,N_11833);
xnor U14463 (N_14463,N_9220,N_11459);
nand U14464 (N_14464,N_10266,N_10344);
xnor U14465 (N_14465,N_7653,N_9000);
or U14466 (N_14466,N_12254,N_10754);
xnor U14467 (N_14467,N_6663,N_11716);
or U14468 (N_14468,N_7192,N_6913);
and U14469 (N_14469,N_6565,N_10251);
nor U14470 (N_14470,N_8575,N_11455);
or U14471 (N_14471,N_11048,N_8238);
xor U14472 (N_14472,N_11809,N_7714);
nor U14473 (N_14473,N_10967,N_7448);
nor U14474 (N_14474,N_10813,N_10730);
or U14475 (N_14475,N_9014,N_7384);
or U14476 (N_14476,N_9153,N_11820);
and U14477 (N_14477,N_8056,N_9598);
xnor U14478 (N_14478,N_7904,N_12012);
nor U14479 (N_14479,N_10414,N_9630);
xnor U14480 (N_14480,N_10442,N_12319);
nand U14481 (N_14481,N_7077,N_10600);
nor U14482 (N_14482,N_11452,N_10959);
and U14483 (N_14483,N_9183,N_12182);
nor U14484 (N_14484,N_11745,N_9519);
xor U14485 (N_14485,N_8090,N_11708);
xnor U14486 (N_14486,N_8190,N_7875);
xor U14487 (N_14487,N_12153,N_6317);
nand U14488 (N_14488,N_11112,N_12452);
nor U14489 (N_14489,N_9952,N_8788);
xnor U14490 (N_14490,N_8822,N_10216);
and U14491 (N_14491,N_12498,N_10042);
nor U14492 (N_14492,N_6468,N_9677);
nor U14493 (N_14493,N_10542,N_7655);
or U14494 (N_14494,N_11483,N_12190);
and U14495 (N_14495,N_9925,N_10430);
nand U14496 (N_14496,N_7933,N_12119);
nand U14497 (N_14497,N_7513,N_10614);
or U14498 (N_14498,N_9765,N_8204);
or U14499 (N_14499,N_10305,N_7458);
xnor U14500 (N_14500,N_7379,N_10244);
xor U14501 (N_14501,N_11175,N_8817);
xor U14502 (N_14502,N_8193,N_11497);
and U14503 (N_14503,N_8281,N_9893);
xor U14504 (N_14504,N_9778,N_8710);
or U14505 (N_14505,N_12032,N_9395);
nand U14506 (N_14506,N_9862,N_10711);
xnor U14507 (N_14507,N_10064,N_11981);
or U14508 (N_14508,N_6962,N_11628);
or U14509 (N_14509,N_8816,N_11980);
nor U14510 (N_14510,N_7147,N_9638);
and U14511 (N_14511,N_8658,N_9011);
and U14512 (N_14512,N_8884,N_7012);
nor U14513 (N_14513,N_7724,N_6377);
nor U14514 (N_14514,N_7808,N_10121);
nor U14515 (N_14515,N_9406,N_6713);
nand U14516 (N_14516,N_6944,N_11373);
nor U14517 (N_14517,N_12142,N_10172);
xnor U14518 (N_14518,N_8139,N_7299);
and U14519 (N_14519,N_11665,N_12010);
nor U14520 (N_14520,N_11280,N_6262);
nor U14521 (N_14521,N_8948,N_12131);
and U14522 (N_14522,N_7116,N_6905);
and U14523 (N_14523,N_9466,N_12404);
and U14524 (N_14524,N_12090,N_12168);
xnor U14525 (N_14525,N_7528,N_11882);
nor U14526 (N_14526,N_8266,N_8317);
nand U14527 (N_14527,N_9319,N_10553);
or U14528 (N_14528,N_10989,N_10355);
nor U14529 (N_14529,N_11866,N_12386);
or U14530 (N_14530,N_7351,N_11813);
nor U14531 (N_14531,N_9607,N_8437);
xnor U14532 (N_14532,N_9662,N_11363);
nor U14533 (N_14533,N_6374,N_7200);
nor U14534 (N_14534,N_7111,N_10857);
nand U14535 (N_14535,N_7455,N_7673);
and U14536 (N_14536,N_8063,N_12082);
xor U14537 (N_14537,N_11901,N_8911);
or U14538 (N_14538,N_9215,N_6545);
nand U14539 (N_14539,N_12011,N_12124);
nor U14540 (N_14540,N_8529,N_6832);
nor U14541 (N_14541,N_10894,N_6900);
nand U14542 (N_14542,N_11562,N_10315);
and U14543 (N_14543,N_9232,N_9978);
and U14544 (N_14544,N_12187,N_11339);
and U14545 (N_14545,N_8551,N_8115);
or U14546 (N_14546,N_9341,N_11325);
xor U14547 (N_14547,N_6619,N_11757);
xnor U14548 (N_14548,N_11219,N_11660);
nand U14549 (N_14549,N_7811,N_8471);
nor U14550 (N_14550,N_6381,N_10537);
xnor U14551 (N_14551,N_9589,N_11620);
xnor U14552 (N_14552,N_9094,N_12093);
or U14553 (N_14553,N_10167,N_10869);
nand U14554 (N_14554,N_7690,N_12372);
or U14555 (N_14555,N_11835,N_8065);
nor U14556 (N_14556,N_11563,N_9841);
xor U14557 (N_14557,N_10955,N_7347);
or U14558 (N_14558,N_9912,N_10201);
nor U14559 (N_14559,N_8336,N_12286);
or U14560 (N_14560,N_12007,N_12442);
or U14561 (N_14561,N_8283,N_8052);
nor U14562 (N_14562,N_10638,N_7508);
nor U14563 (N_14563,N_6343,N_8793);
nor U14564 (N_14564,N_9508,N_12448);
nand U14565 (N_14565,N_7416,N_11807);
or U14566 (N_14566,N_7027,N_6903);
nor U14567 (N_14567,N_6586,N_6781);
nand U14568 (N_14568,N_11220,N_8691);
nand U14569 (N_14569,N_6687,N_7319);
xor U14570 (N_14570,N_11420,N_7328);
nand U14571 (N_14571,N_8137,N_8361);
nor U14572 (N_14572,N_8668,N_7447);
and U14573 (N_14573,N_8599,N_11438);
and U14574 (N_14574,N_6580,N_9186);
nand U14575 (N_14575,N_10175,N_9367);
xor U14576 (N_14576,N_8057,N_6297);
nor U14577 (N_14577,N_10416,N_10092);
and U14578 (N_14578,N_6542,N_8431);
and U14579 (N_14579,N_7679,N_11073);
or U14580 (N_14580,N_7238,N_6284);
nand U14581 (N_14581,N_12255,N_10555);
and U14582 (N_14582,N_11161,N_7474);
nand U14583 (N_14583,N_7940,N_7700);
and U14584 (N_14584,N_11847,N_6721);
and U14585 (N_14585,N_10437,N_7029);
and U14586 (N_14586,N_7887,N_7824);
or U14587 (N_14587,N_8956,N_9629);
nand U14588 (N_14588,N_7274,N_6977);
or U14589 (N_14589,N_11021,N_8346);
and U14590 (N_14590,N_12328,N_12471);
nand U14591 (N_14591,N_6315,N_8124);
and U14592 (N_14592,N_6673,N_7011);
nor U14593 (N_14593,N_9640,N_11838);
or U14594 (N_14594,N_9176,N_7339);
and U14595 (N_14595,N_9699,N_8350);
nor U14596 (N_14596,N_9635,N_7230);
or U14597 (N_14597,N_8851,N_6675);
nor U14598 (N_14598,N_8062,N_9907);
xor U14599 (N_14599,N_12211,N_12356);
or U14600 (N_14600,N_7321,N_11802);
nand U14601 (N_14601,N_11361,N_6314);
nand U14602 (N_14602,N_12041,N_9181);
and U14603 (N_14603,N_6818,N_9144);
xnor U14604 (N_14604,N_11055,N_8180);
or U14605 (N_14605,N_7566,N_10872);
nand U14606 (N_14606,N_10233,N_11094);
xor U14607 (N_14607,N_7952,N_9004);
and U14608 (N_14608,N_11067,N_11036);
xnor U14609 (N_14609,N_7472,N_10513);
nor U14610 (N_14610,N_9608,N_7523);
nor U14611 (N_14611,N_11575,N_9871);
nor U14612 (N_14612,N_11629,N_8280);
xor U14613 (N_14613,N_10413,N_12401);
nand U14614 (N_14614,N_11198,N_8086);
and U14615 (N_14615,N_8036,N_10973);
and U14616 (N_14616,N_9188,N_12269);
nand U14617 (N_14617,N_12412,N_8802);
nor U14618 (N_14618,N_10356,N_10224);
nand U14619 (N_14619,N_10053,N_11111);
or U14620 (N_14620,N_8545,N_6738);
and U14621 (N_14621,N_12087,N_11961);
and U14622 (N_14622,N_8846,N_9707);
xor U14623 (N_14623,N_7507,N_9471);
nor U14624 (N_14624,N_8603,N_11781);
nor U14625 (N_14625,N_10870,N_8513);
xnor U14626 (N_14626,N_9777,N_10170);
or U14627 (N_14627,N_7280,N_11973);
and U14628 (N_14628,N_7795,N_6287);
xor U14629 (N_14629,N_8746,N_12242);
or U14630 (N_14630,N_12389,N_10046);
or U14631 (N_14631,N_8074,N_8785);
nand U14632 (N_14632,N_12450,N_11601);
or U14633 (N_14633,N_7735,N_11970);
and U14634 (N_14634,N_7268,N_7304);
or U14635 (N_14635,N_8619,N_8738);
xnor U14636 (N_14636,N_9143,N_11068);
nor U14637 (N_14637,N_10792,N_11217);
xor U14638 (N_14638,N_10752,N_11604);
nand U14639 (N_14639,N_9043,N_6453);
xnor U14640 (N_14640,N_9741,N_7286);
and U14641 (N_14641,N_9949,N_6765);
xor U14642 (N_14642,N_9289,N_11001);
or U14643 (N_14643,N_8024,N_11595);
or U14644 (N_14644,N_8986,N_10968);
nor U14645 (N_14645,N_10021,N_10527);
or U14646 (N_14646,N_8960,N_12305);
xnor U14647 (N_14647,N_8014,N_11218);
xor U14648 (N_14648,N_11844,N_8946);
or U14649 (N_14649,N_10928,N_9479);
and U14650 (N_14650,N_7910,N_11568);
or U14651 (N_14651,N_6530,N_6782);
nand U14652 (N_14652,N_8049,N_8578);
nand U14653 (N_14653,N_8025,N_12335);
nand U14654 (N_14654,N_10290,N_7997);
nor U14655 (N_14655,N_7257,N_6983);
nand U14656 (N_14656,N_9980,N_9184);
xor U14657 (N_14657,N_7500,N_7307);
nand U14658 (N_14658,N_11850,N_11152);
nand U14659 (N_14659,N_11688,N_9273);
nand U14660 (N_14660,N_11640,N_10195);
nand U14661 (N_14661,N_9563,N_10278);
xnor U14662 (N_14662,N_7716,N_8169);
nor U14663 (N_14663,N_12039,N_12454);
and U14664 (N_14664,N_8142,N_7497);
nand U14665 (N_14665,N_12413,N_11773);
and U14666 (N_14666,N_7555,N_12193);
and U14667 (N_14667,N_7927,N_11025);
and U14668 (N_14668,N_11526,N_11421);
or U14669 (N_14669,N_10713,N_6851);
and U14670 (N_14670,N_12276,N_6429);
or U14671 (N_14671,N_6744,N_9622);
xnor U14672 (N_14672,N_12172,N_10549);
and U14673 (N_14673,N_11839,N_8260);
and U14674 (N_14674,N_11479,N_10006);
or U14675 (N_14675,N_10245,N_10019);
nor U14676 (N_14676,N_12114,N_12347);
nand U14677 (N_14677,N_8955,N_11192);
and U14678 (N_14678,N_6755,N_11148);
or U14679 (N_14679,N_6999,N_7064);
or U14680 (N_14680,N_11402,N_10146);
nor U14681 (N_14681,N_11531,N_7516);
and U14682 (N_14682,N_11410,N_6754);
nand U14683 (N_14683,N_11171,N_10798);
and U14684 (N_14684,N_9070,N_10581);
and U14685 (N_14685,N_12151,N_6599);
nand U14686 (N_14686,N_6404,N_6371);
and U14687 (N_14687,N_8934,N_11292);
xor U14688 (N_14688,N_12091,N_11163);
or U14689 (N_14689,N_8662,N_12078);
and U14690 (N_14690,N_9050,N_7039);
xor U14691 (N_14691,N_6446,N_8101);
or U14692 (N_14692,N_8082,N_10927);
nor U14693 (N_14693,N_8764,N_10237);
xnor U14694 (N_14694,N_10166,N_7919);
or U14695 (N_14695,N_11992,N_9399);
nor U14696 (N_14696,N_7854,N_7816);
nand U14697 (N_14697,N_9727,N_10385);
xnor U14698 (N_14698,N_11602,N_6968);
and U14699 (N_14699,N_7658,N_11430);
and U14700 (N_14700,N_9555,N_10041);
xor U14701 (N_14701,N_8812,N_10954);
nor U14702 (N_14702,N_6633,N_7756);
nand U14703 (N_14703,N_9038,N_7871);
nand U14704 (N_14704,N_8910,N_11988);
or U14705 (N_14705,N_8689,N_11183);
nor U14706 (N_14706,N_11499,N_7237);
nor U14707 (N_14707,N_9972,N_10602);
and U14708 (N_14708,N_10543,N_7692);
and U14709 (N_14709,N_6762,N_8667);
or U14710 (N_14710,N_6486,N_7603);
and U14711 (N_14711,N_7037,N_9962);
or U14712 (N_14712,N_6957,N_8587);
or U14713 (N_14713,N_9320,N_10590);
nand U14714 (N_14714,N_9396,N_9342);
nor U14715 (N_14715,N_12148,N_9062);
and U14716 (N_14716,N_9272,N_7214);
and U14717 (N_14717,N_11508,N_9446);
or U14718 (N_14718,N_12089,N_9086);
xnor U14719 (N_14719,N_10979,N_10635);
nand U14720 (N_14720,N_12005,N_8353);
xor U14721 (N_14721,N_8188,N_11822);
nand U14722 (N_14722,N_7545,N_12101);
nand U14723 (N_14723,N_7855,N_8047);
nor U14724 (N_14724,N_11931,N_8644);
or U14725 (N_14725,N_10261,N_8186);
xnor U14726 (N_14726,N_7922,N_11157);
and U14727 (N_14727,N_7172,N_8695);
nor U14728 (N_14728,N_10753,N_9304);
nor U14729 (N_14729,N_7617,N_8686);
nor U14730 (N_14730,N_9315,N_8202);
nand U14731 (N_14731,N_9847,N_11940);
nor U14732 (N_14732,N_11587,N_10277);
and U14733 (N_14733,N_12306,N_7620);
and U14734 (N_14734,N_10806,N_7924);
xor U14735 (N_14735,N_8574,N_11491);
nor U14736 (N_14736,N_8626,N_11695);
xor U14737 (N_14737,N_11574,N_9729);
and U14738 (N_14738,N_10179,N_8391);
xnor U14739 (N_14739,N_7178,N_9177);
nand U14740 (N_14740,N_9087,N_11070);
and U14741 (N_14741,N_11248,N_10039);
xor U14742 (N_14742,N_6366,N_8709);
nor U14743 (N_14743,N_9180,N_8168);
or U14744 (N_14744,N_11831,N_10761);
nor U14745 (N_14745,N_11187,N_9335);
and U14746 (N_14746,N_8002,N_7110);
nand U14747 (N_14747,N_7496,N_8937);
nand U14748 (N_14748,N_12482,N_10992);
nor U14749 (N_14749,N_11490,N_10931);
xor U14750 (N_14750,N_12178,N_7264);
xor U14751 (N_14751,N_9127,N_8493);
xnor U14752 (N_14752,N_10578,N_6463);
nand U14753 (N_14753,N_10365,N_12264);
nor U14754 (N_14754,N_8041,N_10208);
nor U14755 (N_14755,N_7356,N_11506);
nand U14756 (N_14756,N_6456,N_12278);
or U14757 (N_14757,N_9611,N_10065);
nor U14758 (N_14758,N_8711,N_9712);
and U14759 (N_14759,N_9721,N_11785);
nor U14760 (N_14760,N_7873,N_8104);
xor U14761 (N_14761,N_10268,N_12224);
nand U14762 (N_14762,N_8592,N_6443);
nor U14763 (N_14763,N_8654,N_12002);
nand U14764 (N_14764,N_7872,N_10501);
or U14765 (N_14765,N_7521,N_9124);
and U14766 (N_14766,N_7731,N_6472);
xor U14767 (N_14767,N_12149,N_10632);
nand U14768 (N_14768,N_7880,N_6638);
nor U14769 (N_14769,N_6731,N_11474);
nor U14770 (N_14770,N_11211,N_11843);
and U14771 (N_14771,N_10631,N_6910);
xnor U14772 (N_14772,N_6822,N_9970);
and U14773 (N_14773,N_7495,N_7771);
nor U14774 (N_14774,N_9080,N_8046);
nor U14775 (N_14775,N_7677,N_12485);
or U14776 (N_14776,N_8996,N_6893);
nand U14777 (N_14777,N_9900,N_11170);
or U14778 (N_14778,N_7102,N_7308);
and U14779 (N_14779,N_8534,N_9239);
nor U14780 (N_14780,N_11648,N_8651);
or U14781 (N_14781,N_10420,N_9578);
xnor U14782 (N_14782,N_8801,N_8398);
xnor U14783 (N_14783,N_11104,N_11954);
nand U14784 (N_14784,N_11798,N_9693);
nor U14785 (N_14785,N_8229,N_10930);
or U14786 (N_14786,N_6975,N_6267);
and U14787 (N_14787,N_6866,N_11269);
nand U14788 (N_14788,N_8001,N_11880);
or U14789 (N_14789,N_12464,N_8674);
nand U14790 (N_14790,N_7345,N_10585);
or U14791 (N_14791,N_7169,N_7327);
nor U14792 (N_14792,N_8112,N_8122);
and U14793 (N_14793,N_9218,N_8623);
or U14794 (N_14794,N_8221,N_12469);
or U14795 (N_14795,N_8200,N_9784);
xor U14796 (N_14796,N_10147,N_9618);
or U14797 (N_14797,N_7368,N_8998);
nand U14798 (N_14798,N_11020,N_10351);
or U14799 (N_14799,N_8732,N_9171);
xnor U14800 (N_14800,N_6787,N_9596);
nor U14801 (N_14801,N_7654,N_8877);
xnor U14802 (N_14802,N_6281,N_11431);
or U14803 (N_14803,N_7821,N_11714);
or U14804 (N_14804,N_12441,N_6678);
or U14805 (N_14805,N_9123,N_12363);
xor U14806 (N_14806,N_8719,N_7219);
nor U14807 (N_14807,N_11725,N_9475);
or U14808 (N_14808,N_11643,N_8466);
xnor U14809 (N_14809,N_9378,N_11678);
nor U14810 (N_14810,N_8035,N_9518);
or U14811 (N_14811,N_11428,N_7180);
or U14812 (N_14812,N_7711,N_8763);
nor U14813 (N_14813,N_11342,N_9453);
nor U14814 (N_14814,N_7546,N_12205);
and U14815 (N_14815,N_8003,N_9036);
xor U14816 (N_14816,N_10300,N_9815);
nand U14817 (N_14817,N_6309,N_6915);
xor U14818 (N_14818,N_11801,N_9999);
or U14819 (N_14819,N_12009,N_7902);
xor U14820 (N_14820,N_12341,N_10353);
xor U14821 (N_14821,N_7228,N_12135);
xor U14822 (N_14822,N_8326,N_11498);
and U14823 (N_14823,N_8207,N_8465);
xor U14824 (N_14824,N_12400,N_12277);
and U14825 (N_14825,N_12163,N_10331);
or U14826 (N_14826,N_10329,N_8682);
nor U14827 (N_14827,N_11582,N_10279);
and U14828 (N_14828,N_9045,N_9010);
and U14829 (N_14829,N_11689,N_11960);
nand U14830 (N_14830,N_6967,N_10693);
or U14831 (N_14831,N_8647,N_10327);
and U14832 (N_14832,N_8836,N_9293);
nor U14833 (N_14833,N_6806,N_10298);
nand U14834 (N_14834,N_12303,N_9530);
and U14835 (N_14835,N_6449,N_11984);
xnor U14836 (N_14836,N_6670,N_7812);
and U14837 (N_14837,N_7642,N_11069);
and U14838 (N_14838,N_10081,N_9051);
nand U14839 (N_14839,N_11019,N_11088);
and U14840 (N_14840,N_7073,N_6340);
xor U14841 (N_14841,N_11567,N_8390);
nor U14842 (N_14842,N_11564,N_8064);
xor U14843 (N_14843,N_10436,N_11413);
nor U14844 (N_14844,N_9989,N_11445);
and U14845 (N_14845,N_6950,N_10704);
nand U14846 (N_14846,N_10188,N_11131);
and U14847 (N_14847,N_10287,N_8328);
or U14848 (N_14848,N_11352,N_10568);
nand U14849 (N_14849,N_9650,N_6275);
nor U14850 (N_14850,N_8164,N_9718);
or U14851 (N_14851,N_8222,N_7591);
nand U14852 (N_14852,N_12226,N_10755);
and U14853 (N_14853,N_9317,N_8451);
nand U14854 (N_14854,N_9605,N_9621);
nand U14855 (N_14855,N_6295,N_12473);
xnor U14856 (N_14856,N_8083,N_7981);
and U14857 (N_14857,N_10654,N_6669);
xnor U14858 (N_14858,N_11326,N_11252);
nor U14859 (N_14859,N_10312,N_6280);
xnor U14860 (N_14860,N_9237,N_10083);
xor U14861 (N_14861,N_9402,N_10564);
nand U14862 (N_14862,N_10674,N_10453);
or U14863 (N_14863,N_7087,N_10316);
or U14864 (N_14864,N_11384,N_10712);
xnor U14865 (N_14865,N_12120,N_9409);
nand U14866 (N_14866,N_7387,N_11800);
nand U14867 (N_14867,N_8913,N_11327);
xnor U14868 (N_14868,N_9486,N_7401);
or U14869 (N_14869,N_8043,N_11632);
or U14870 (N_14870,N_7294,N_12283);
nand U14871 (N_14871,N_6847,N_8516);
nand U14872 (N_14872,N_6795,N_6447);
nor U14873 (N_14873,N_12077,N_11113);
nor U14874 (N_14874,N_10771,N_8508);
nor U14875 (N_14875,N_9414,N_10164);
nor U14876 (N_14876,N_7707,N_10744);
xnor U14877 (N_14877,N_10094,N_10822);
nand U14878 (N_14878,N_10445,N_10663);
nor U14879 (N_14879,N_11919,N_7682);
and U14880 (N_14880,N_6459,N_11398);
nor U14881 (N_14881,N_7779,N_7763);
or U14882 (N_14882,N_11627,N_6300);
nor U14883 (N_14883,N_7863,N_7259);
and U14884 (N_14884,N_9814,N_11397);
nand U14885 (N_14885,N_7124,N_7223);
and U14886 (N_14886,N_12470,N_6269);
nor U14887 (N_14887,N_9060,N_8123);
nor U14888 (N_14888,N_12191,N_11962);
nor U14889 (N_14889,N_8409,N_8498);
nand U14890 (N_14890,N_11261,N_8707);
or U14891 (N_14891,N_6460,N_7708);
and U14892 (N_14892,N_7056,N_11440);
nand U14893 (N_14893,N_10128,N_12468);
or U14894 (N_14894,N_9516,N_8166);
xor U14895 (N_14895,N_10252,N_7817);
or U14896 (N_14896,N_9151,N_6993);
nand U14897 (N_14897,N_7993,N_8607);
nand U14898 (N_14898,N_9024,N_6427);
or U14899 (N_14899,N_9468,N_11296);
and U14900 (N_14900,N_12230,N_10239);
or U14901 (N_14901,N_12130,N_7190);
nand U14902 (N_14902,N_10824,N_8918);
nand U14903 (N_14903,N_10091,N_11814);
nand U14904 (N_14904,N_8855,N_10379);
xnor U14905 (N_14905,N_8841,N_7325);
xor U14906 (N_14906,N_10552,N_12434);
or U14907 (N_14907,N_8706,N_7198);
or U14908 (N_14908,N_7625,N_8850);
xnor U14909 (N_14909,N_11369,N_7862);
or U14910 (N_14910,N_12453,N_8739);
and U14911 (N_14911,N_7499,N_10816);
or U14912 (N_14912,N_10777,N_6562);
xnor U14913 (N_14913,N_7709,N_6876);
nand U14914 (N_14914,N_10491,N_7402);
nand U14915 (N_14915,N_9302,N_11026);
and U14916 (N_14916,N_8881,N_9828);
nor U14917 (N_14917,N_6879,N_7749);
nor U14918 (N_14918,N_11275,N_9256);
xor U14919 (N_14919,N_8863,N_6887);
and U14920 (N_14920,N_9536,N_11473);
and U14921 (N_14921,N_10295,N_11260);
or U14922 (N_14922,N_9107,N_8044);
and U14923 (N_14923,N_9834,N_8598);
xor U14924 (N_14924,N_9490,N_11815);
nor U14925 (N_14925,N_8909,N_6935);
nor U14926 (N_14926,N_11846,N_10018);
or U14927 (N_14927,N_10706,N_6660);
or U14928 (N_14928,N_9394,N_7303);
or U14929 (N_14929,N_10887,N_8434);
or U14930 (N_14930,N_10823,N_9387);
nand U14931 (N_14931,N_7504,N_8571);
and U14932 (N_14932,N_7552,N_6506);
xnor U14933 (N_14933,N_9620,N_7806);
or U14934 (N_14934,N_8425,N_6870);
and U14935 (N_14935,N_9850,N_6346);
or U14936 (N_14936,N_8299,N_6258);
nand U14937 (N_14937,N_12447,N_11636);
and U14938 (N_14938,N_8363,N_10685);
xnor U14939 (N_14939,N_6583,N_10859);
and U14940 (N_14940,N_9566,N_8828);
or U14941 (N_14941,N_9357,N_9817);
and U14942 (N_14942,N_9975,N_11424);
nand U14943 (N_14943,N_7245,N_9348);
and U14944 (N_14944,N_11778,N_7995);
or U14945 (N_14945,N_10002,N_6283);
or U14946 (N_14946,N_8690,N_8514);
or U14947 (N_14947,N_12157,N_7534);
xor U14948 (N_14948,N_11103,N_6290);
and U14949 (N_14949,N_10905,N_11013);
and U14950 (N_14950,N_7764,N_6253);
nand U14951 (N_14951,N_7052,N_12440);
nor U14952 (N_14952,N_7217,N_7408);
nand U14953 (N_14953,N_7067,N_7377);
or U14954 (N_14954,N_6250,N_6890);
and U14955 (N_14955,N_12274,N_10120);
xor U14956 (N_14956,N_11439,N_8149);
xnor U14957 (N_14957,N_6802,N_7373);
nand U14958 (N_14958,N_8099,N_10854);
nor U14959 (N_14959,N_10698,N_9072);
nand U14960 (N_14960,N_11383,N_10988);
nand U14961 (N_14961,N_10618,N_9179);
nand U14962 (N_14962,N_11422,N_10173);
xor U14963 (N_14963,N_10492,N_8680);
nor U14964 (N_14964,N_8108,N_10157);
and U14965 (N_14965,N_8572,N_8019);
nand U14966 (N_14966,N_8897,N_9485);
nand U14967 (N_14967,N_6424,N_7170);
or U14968 (N_14968,N_12260,N_8120);
nor U14969 (N_14969,N_8657,N_8100);
nor U14970 (N_14970,N_9945,N_9800);
and U14971 (N_14971,N_10842,N_9103);
nor U14972 (N_14972,N_8637,N_10476);
nor U14973 (N_14973,N_11132,N_10812);
or U14974 (N_14974,N_7317,N_12478);
and U14975 (N_14975,N_9331,N_7937);
xnor U14976 (N_14976,N_7287,N_7293);
or U14977 (N_14977,N_11787,N_6502);
and U14978 (N_14978,N_9420,N_7502);
nand U14979 (N_14979,N_11550,N_11638);
nor U14980 (N_14980,N_6886,N_10477);
or U14981 (N_14981,N_11109,N_6789);
or U14982 (N_14982,N_11613,N_11854);
and U14983 (N_14983,N_11552,N_7975);
or U14984 (N_14984,N_10198,N_12407);
and U14985 (N_14985,N_11775,N_10831);
and U14986 (N_14986,N_8945,N_7279);
and U14987 (N_14987,N_7998,N_7805);
or U14988 (N_14988,N_6544,N_11281);
or U14989 (N_14989,N_8872,N_9545);
and U14990 (N_14990,N_9873,N_11457);
and U14991 (N_14991,N_9760,N_9979);
xor U14992 (N_14992,N_7001,N_11135);
nor U14993 (N_14993,N_7826,N_7564);
and U14994 (N_14994,N_6578,N_10668);
and U14995 (N_14995,N_6715,N_9245);
nand U14996 (N_14996,N_10994,N_8521);
nand U14997 (N_14997,N_11547,N_7611);
xnor U14998 (N_14998,N_6518,N_12287);
and U14999 (N_14999,N_8670,N_8017);
nor U15000 (N_15000,N_9326,N_11446);
nand U15001 (N_15001,N_7623,N_10963);
nand U15002 (N_15002,N_9075,N_12467);
or U15003 (N_15003,N_10848,N_9544);
and U15004 (N_15004,N_9049,N_12123);
xnor U15005 (N_15005,N_12059,N_9370);
and U15006 (N_15006,N_10393,N_7928);
or U15007 (N_15007,N_10246,N_11928);
or U15008 (N_15008,N_8823,N_11493);
nor U15009 (N_15009,N_11033,N_9233);
or U15010 (N_15010,N_12126,N_8726);
xor U15011 (N_15011,N_10982,N_7622);
xor U15012 (N_15012,N_8735,N_7104);
xor U15013 (N_15013,N_11374,N_11792);
nor U15014 (N_15014,N_12463,N_7160);
nor U15015 (N_15015,N_8704,N_8773);
and U15016 (N_15016,N_10144,N_10372);
or U15017 (N_15017,N_10052,N_10136);
xnor U15018 (N_15018,N_7315,N_7803);
nor U15019 (N_15019,N_6970,N_10970);
xor U15020 (N_15020,N_12284,N_6743);
or U15021 (N_15021,N_10483,N_8256);
nand U15022 (N_15022,N_6682,N_11053);
nor U15023 (N_15023,N_12137,N_6277);
nor U15024 (N_15024,N_7978,N_8625);
and U15025 (N_15025,N_8907,N_9706);
nor U15026 (N_15026,N_11461,N_10015);
nor U15027 (N_15027,N_11279,N_9823);
nor U15028 (N_15028,N_6990,N_8324);
nand U15029 (N_15029,N_7329,N_8095);
nand U15030 (N_15030,N_11958,N_7912);
xor U15031 (N_15031,N_7231,N_11471);
or U15032 (N_15032,N_10646,N_9795);
and U15033 (N_15033,N_10472,N_11618);
nand U15034 (N_15034,N_8659,N_8294);
or U15035 (N_15035,N_9389,N_11522);
nand U15036 (N_15036,N_7570,N_12427);
nand U15037 (N_15037,N_12487,N_8724);
xor U15038 (N_15038,N_11642,N_9626);
nor U15039 (N_15039,N_8525,N_8980);
nand U15040 (N_15040,N_9628,N_9340);
nand U15041 (N_15041,N_11834,N_11523);
and U15042 (N_15042,N_7575,N_9306);
or U15043 (N_15043,N_7684,N_12019);
or U15044 (N_15044,N_12360,N_9855);
or U15045 (N_15045,N_9009,N_11359);
nor U15046 (N_15046,N_10776,N_11731);
or U15047 (N_15047,N_7288,N_11704);
or U15048 (N_15048,N_8287,N_12299);
nor U15049 (N_15049,N_7959,N_9624);
nand U15050 (N_15050,N_10342,N_9869);
nor U15051 (N_15051,N_9933,N_11273);
and U15052 (N_15052,N_10808,N_11571);
xnor U15053 (N_15053,N_12071,N_9467);
and U15054 (N_15054,N_10620,N_11722);
nor U15055 (N_15055,N_8154,N_6699);
nor U15056 (N_15056,N_8722,N_10384);
xnor U15057 (N_15057,N_10346,N_6691);
nand U15058 (N_15058,N_6396,N_11130);
and U15059 (N_15059,N_10214,N_10682);
xnor U15060 (N_15060,N_10724,N_10333);
xnor U15061 (N_15061,N_9114,N_7091);
nor U15062 (N_15062,N_10696,N_7041);
and U15063 (N_15063,N_11380,N_9147);
nor U15064 (N_15064,N_12080,N_9451);
or U15065 (N_15065,N_12056,N_8556);
nand U15066 (N_15066,N_10096,N_8483);
nor U15067 (N_15067,N_12167,N_6256);
xnor U15068 (N_15068,N_8485,N_7576);
or U15069 (N_15069,N_11907,N_9648);
nand U15070 (N_15070,N_11142,N_11058);
xnor U15071 (N_15071,N_12366,N_11519);
nor U15072 (N_15072,N_6293,N_8989);
and U15073 (N_15073,N_7460,N_10686);
nor U15074 (N_15074,N_10069,N_7436);
nand U15075 (N_15075,N_9443,N_9937);
nand U15076 (N_15076,N_9564,N_6624);
xor U15077 (N_15077,N_7255,N_11864);
nor U15078 (N_15078,N_7254,N_8636);
xor U15079 (N_15079,N_10161,N_6278);
xnor U15080 (N_15080,N_9813,N_7483);
xor U15081 (N_15081,N_8389,N_11738);
xnor U15082 (N_15082,N_9219,N_9454);
xnor U15083 (N_15083,N_11525,N_9197);
and U15084 (N_15084,N_11056,N_9019);
and U15085 (N_15085,N_11039,N_10247);
nand U15086 (N_15086,N_8630,N_9854);
and U15087 (N_15087,N_7825,N_6353);
and U15088 (N_15088,N_8541,N_8629);
or U15089 (N_15089,N_12055,N_7167);
nor U15090 (N_15090,N_7948,N_8147);
nand U15091 (N_15091,N_10591,N_6559);
and U15092 (N_15092,N_9625,N_11258);
and U15093 (N_15093,N_10742,N_6591);
xor U15094 (N_15094,N_9822,N_8276);
nand U15095 (N_15095,N_11074,N_7832);
or U15096 (N_15096,N_12290,N_12164);
or U15097 (N_15097,N_11630,N_7956);
nand U15098 (N_15098,N_7481,N_7338);
xor U15099 (N_15099,N_9194,N_11623);
or U15100 (N_15100,N_7911,N_7533);
nand U15101 (N_15101,N_8870,N_7901);
nor U15102 (N_15102,N_7809,N_11060);
nor U15103 (N_15103,N_10626,N_7849);
and U15104 (N_15104,N_10521,N_8345);
or U15105 (N_15105,N_10800,N_7284);
nor U15106 (N_15106,N_10676,N_12058);
nand U15107 (N_15107,N_7156,N_12437);
and U15108 (N_15108,N_10309,N_7609);
xor U15109 (N_15109,N_9770,N_6788);
or U15110 (N_15110,N_12203,N_10514);
or U15111 (N_15111,N_6590,N_12202);
nor U15112 (N_15112,N_9865,N_10616);
and U15113 (N_15113,N_10962,N_8426);
or U15114 (N_15114,N_9636,N_10258);
nor U15115 (N_15115,N_11090,N_6439);
nand U15116 (N_15116,N_8045,N_8289);
xor U15117 (N_15117,N_10158,N_6807);
or U15118 (N_15118,N_6323,N_11399);
xor U15119 (N_15119,N_10060,N_10059);
or U15120 (N_15120,N_9863,N_7687);
nand U15121 (N_15121,N_8586,N_11290);
or U15122 (N_15122,N_8972,N_8246);
and U15123 (N_15123,N_8027,N_10189);
and U15124 (N_15124,N_9003,N_9928);
nand U15125 (N_15125,N_7836,N_8339);
nor U15126 (N_15126,N_12145,N_6976);
xor U15127 (N_15127,N_6260,N_6320);
and U15128 (N_15128,N_7080,N_7621);
nand U15129 (N_15129,N_8162,N_12445);
and U15130 (N_15130,N_6480,N_6418);
or U15131 (N_15131,N_12073,N_8604);
and U15132 (N_15132,N_7835,N_12022);
and U15133 (N_15133,N_6508,N_6969);
nor U15134 (N_15134,N_9738,N_10601);
nor U15135 (N_15135,N_7158,N_11379);
or U15136 (N_15136,N_7843,N_9307);
nand U15137 (N_15137,N_9681,N_10338);
and U15138 (N_15138,N_9216,N_6537);
xor U15139 (N_15139,N_7289,N_11926);
and U15140 (N_15140,N_8962,N_11174);
xor U15141 (N_15141,N_11631,N_9379);
and U15142 (N_15142,N_6973,N_11259);
nand U15143 (N_15143,N_7571,N_11540);
xnor U15144 (N_15144,N_6862,N_10027);
or U15145 (N_15145,N_7125,N_6361);
xnor U15146 (N_15146,N_6628,N_10762);
xnor U15147 (N_15147,N_6517,N_6901);
nand U15148 (N_15148,N_11881,N_10074);
nand U15149 (N_15149,N_12081,N_9243);
xor U15150 (N_15150,N_9016,N_11929);
nand U15151 (N_15151,N_7313,N_10836);
nand U15152 (N_15152,N_7112,N_11271);
nand U15153 (N_15153,N_7511,N_10510);
and U15154 (N_15154,N_7865,N_11805);
xor U15155 (N_15155,N_6952,N_8392);
or U15156 (N_15156,N_7813,N_12000);
nand U15157 (N_15157,N_8867,N_9782);
and U15158 (N_15158,N_11463,N_8175);
nor U15159 (N_15159,N_10238,N_8349);
and U15160 (N_15160,N_6413,N_8968);
xnor U15161 (N_15161,N_10731,N_6533);
or U15162 (N_15162,N_6695,N_6490);
or U15163 (N_15163,N_8396,N_8650);
nand U15164 (N_15164,N_7247,N_9223);
nor U15165 (N_15165,N_10868,N_8449);
and U15166 (N_15166,N_11037,N_7057);
xnor U15167 (N_15167,N_6701,N_12197);
or U15168 (N_15168,N_12432,N_9789);
nand U15169 (N_15169,N_7969,N_10779);
and U15170 (N_15170,N_7541,N_11569);
nand U15171 (N_15171,N_6593,N_6843);
and U15172 (N_15172,N_12220,N_11502);
nor U15173 (N_15173,N_9286,N_11091);
nor U15174 (N_15174,N_9745,N_7220);
nand U15175 (N_15175,N_8382,N_12369);
nand U15176 (N_15176,N_12246,N_9788);
or U15177 (N_15177,N_9412,N_7446);
and U15178 (N_15178,N_7983,N_8315);
nor U15179 (N_15179,N_11338,N_7674);
xnor U15180 (N_15180,N_11167,N_11193);
or U15181 (N_15181,N_6416,N_7651);
nor U15182 (N_15182,N_10769,N_11606);
and U15183 (N_15183,N_7531,N_8579);
or U15184 (N_15184,N_8010,N_6329);
and U15185 (N_15185,N_6492,N_10645);
xnor U15186 (N_15186,N_12243,N_9386);
and U15187 (N_15187,N_8444,N_10584);
or U15188 (N_15188,N_10787,N_12072);
xnor U15189 (N_15189,N_10763,N_9472);
or U15190 (N_15190,N_9513,N_10835);
and U15191 (N_15191,N_9361,N_9932);
nand U15192 (N_15192,N_9119,N_9142);
and U15193 (N_15193,N_10075,N_8091);
or U15194 (N_15194,N_10726,N_12158);
nand U15195 (N_15195,N_8241,N_8978);
and U15196 (N_15196,N_10440,N_8522);
and U15197 (N_15197,N_9668,N_8456);
xnor U15198 (N_15198,N_6560,N_10738);
nand U15199 (N_15199,N_11240,N_8883);
nor U15200 (N_15200,N_8736,N_6259);
nand U15201 (N_15201,N_10604,N_9462);
nand U15202 (N_15202,N_6623,N_11494);
xor U15203 (N_15203,N_7726,N_6995);
xnor U15204 (N_15204,N_9637,N_7035);
or U15205 (N_15205,N_9506,N_7120);
and U15206 (N_15206,N_7522,N_11080);
nand U15207 (N_15207,N_9491,N_6700);
nand U15208 (N_15208,N_8347,N_6335);
or U15209 (N_15209,N_11059,N_10830);
or U15210 (N_15210,N_8581,N_6540);
and U15211 (N_15211,N_8606,N_10571);
nor U15212 (N_15212,N_6592,N_10014);
or U15213 (N_15213,N_7712,N_6711);
and U15214 (N_15214,N_12188,N_7108);
nand U15215 (N_15215,N_7889,N_10336);
or U15216 (N_15216,N_9226,N_11558);
and U15217 (N_15217,N_8582,N_8026);
xnor U15218 (N_15218,N_12373,N_8316);
nor U15219 (N_15219,N_12125,N_6511);
nand U15220 (N_15220,N_9950,N_11841);
or U15221 (N_15221,N_12376,N_6388);
nor U15222 (N_15222,N_10723,N_11392);
xnor U15223 (N_15223,N_7273,N_11717);
nor U15224 (N_15224,N_11222,N_10952);
xnor U15225 (N_15225,N_9375,N_10799);
nor U15226 (N_15226,N_9065,N_9251);
nand U15227 (N_15227,N_8491,N_9095);
nand U15228 (N_15228,N_7913,N_10493);
xor U15229 (N_15229,N_7476,N_10756);
xnor U15230 (N_15230,N_10783,N_11164);
or U15231 (N_15231,N_7626,N_9487);
nand U15232 (N_15232,N_8005,N_7868);
xnor U15233 (N_15233,N_11935,N_9313);
nor U15234 (N_15234,N_10789,N_12156);
or U15235 (N_15235,N_10879,N_7068);
xnor U15236 (N_15236,N_9787,N_11406);
and U15237 (N_15237,N_8688,N_11821);
xnor U15238 (N_15238,N_9295,N_7427);
and U15239 (N_15239,N_11408,N_11375);
or U15240 (N_15240,N_9444,N_7768);
and U15241 (N_15241,N_7883,N_6603);
or U15242 (N_15242,N_7042,N_10670);
and U15243 (N_15243,N_11119,N_10433);
or U15244 (N_15244,N_11264,N_8950);
nand U15245 (N_15245,N_7694,N_9827);
xor U15246 (N_15246,N_11034,N_7179);
or U15247 (N_15247,N_8205,N_8932);
and U15248 (N_15248,N_10234,N_10772);
and U15249 (N_15249,N_8825,N_6815);
nor U15250 (N_15250,N_10615,N_11593);
or U15251 (N_15251,N_6496,N_9714);
xnor U15252 (N_15252,N_8171,N_8896);
or U15253 (N_15253,N_9157,N_6626);
xnor U15254 (N_15254,N_9702,N_6408);
nand U15255 (N_15255,N_10983,N_12351);
or U15256 (N_15256,N_7277,N_6632);
and U15257 (N_15257,N_10906,N_8126);
or U15258 (N_15258,N_9665,N_11770);
nand U15259 (N_15259,N_7851,N_7947);
or U15260 (N_15260,N_6917,N_10033);
xnor U15261 (N_15261,N_8482,N_8248);
nor U15262 (N_15262,N_10497,N_11194);
xnor U15263 (N_15263,N_7235,N_7376);
and U15264 (N_15264,N_10183,N_9599);
nand U15265 (N_15265,N_10847,N_8975);
xor U15266 (N_15266,N_6352,N_10026);
nor U15267 (N_15267,N_6688,N_10865);
or U15268 (N_15268,N_10524,N_12393);
nor U15269 (N_15269,N_11585,N_10218);
or U15270 (N_15270,N_11968,N_11739);
and U15271 (N_15271,N_11845,N_11411);
xnor U15272 (N_15272,N_8994,N_8769);
and U15273 (N_15273,N_6941,N_11266);
nor U15274 (N_15274,N_11169,N_6423);
xor U15275 (N_15275,N_12396,N_10675);
or U15276 (N_15276,N_6403,N_6961);
xnor U15277 (N_15277,N_11509,N_10838);
xor U15278 (N_15278,N_9039,N_9735);
nand U15279 (N_15279,N_9571,N_10987);
nand U15280 (N_15280,N_9708,N_8214);
nand U15281 (N_15281,N_10739,N_9418);
or U15282 (N_15282,N_11667,N_10609);
nor U15283 (N_15283,N_7473,N_9112);
nand U15284 (N_15284,N_9583,N_6760);
and U15285 (N_15285,N_10152,N_6936);
or U15286 (N_15286,N_7785,N_10672);
xor U15287 (N_15287,N_12365,N_12433);
xor U15288 (N_15288,N_6575,N_10819);
xnor U15289 (N_15289,N_11719,N_7137);
or U15290 (N_15290,N_6458,N_10640);
and U15291 (N_15291,N_11671,N_9790);
nand U15292 (N_15292,N_9669,N_7271);
nand U15293 (N_15293,N_7594,N_6595);
and U15294 (N_15294,N_6856,N_10302);
or U15295 (N_15295,N_7423,N_10736);
and U15296 (N_15296,N_6462,N_12136);
nor U15297 (N_15297,N_11150,N_11065);
or U15298 (N_15298,N_7548,N_7372);
or U15299 (N_15299,N_9783,N_11826);
and U15300 (N_15300,N_10459,N_6291);
or U15301 (N_15301,N_8974,N_10757);
and U15302 (N_15302,N_9899,N_10969);
xnor U15303 (N_15303,N_6759,N_7353);
xnor U15304 (N_15304,N_10902,N_9859);
xnor U15305 (N_15305,N_6676,N_7335);
or U15306 (N_15306,N_12382,N_6794);
and U15307 (N_15307,N_6528,N_6597);
nand U15308 (N_15308,N_6656,N_6841);
nand U15309 (N_15309,N_11751,N_7498);
and U15310 (N_15310,N_11936,N_10101);
or U15311 (N_15311,N_12034,N_9709);
or U15312 (N_15312,N_11477,N_10241);
nor U15313 (N_15313,N_9934,N_6345);
and U15314 (N_15314,N_9461,N_7342);
and U15315 (N_15315,N_10051,N_6428);
nor U15316 (N_15316,N_8900,N_6302);
and U15317 (N_15317,N_11737,N_10260);
or U15318 (N_15318,N_7864,N_7730);
nor U15319 (N_15319,N_10024,N_10759);
or U15320 (N_15320,N_9270,N_8393);
or U15321 (N_15321,N_12199,N_8733);
xor U15322 (N_15322,N_8218,N_8815);
and U15323 (N_15323,N_6693,N_12377);
or U15324 (N_15324,N_10873,N_9802);
nor U15325 (N_15325,N_8531,N_7543);
xnor U15326 (N_15326,N_6697,N_7781);
or U15327 (N_15327,N_10947,N_9959);
and U15328 (N_15328,N_7165,N_7728);
xor U15329 (N_15329,N_10677,N_8641);
nand U15330 (N_15330,N_12368,N_9523);
and U15331 (N_15331,N_7033,N_8279);
nor U15332 (N_15332,N_11318,N_11752);
nor U15333 (N_15333,N_8675,N_7468);
nor U15334 (N_15334,N_6568,N_10275);
xor U15335 (N_15335,N_6354,N_11639);
or U15336 (N_15336,N_6776,N_8871);
and U15337 (N_15337,N_10561,N_8459);
nand U15338 (N_15338,N_7930,N_7451);
xor U15339 (N_15339,N_11872,N_8864);
nand U15340 (N_15340,N_11682,N_11888);
or U15341 (N_15341,N_7945,N_9710);
or U15342 (N_15342,N_10950,N_11007);
nand U15343 (N_15343,N_8713,N_10345);
and U15344 (N_15344,N_7659,N_11335);
nor U15345 (N_15345,N_12028,N_11950);
and U15346 (N_15346,N_7028,N_8211);
nand U15347 (N_15347,N_10680,N_7464);
or U15348 (N_15348,N_8969,N_10689);
nor U15349 (N_15349,N_6769,N_10412);
and U15350 (N_15350,N_10727,N_9473);
and U15351 (N_15351,N_8415,N_12297);
xnor U15352 (N_15352,N_11879,N_11257);
or U15353 (N_15353,N_9874,N_11049);
nor U15354 (N_15354,N_9619,N_6311);
or U15355 (N_15355,N_11129,N_11419);
or U15356 (N_15356,N_12338,N_8696);
nor U15357 (N_15357,N_10673,N_9957);
nand U15358 (N_15358,N_8480,N_7484);
xnor U15359 (N_15359,N_9397,N_10803);
nor U15360 (N_15360,N_8467,N_7729);
or U15361 (N_15361,N_6417,N_12273);
xor U15362 (N_15362,N_12014,N_9431);
nor U15363 (N_15363,N_6563,N_11311);
or U15364 (N_15364,N_9182,N_8660);
or U15365 (N_15365,N_9426,N_9798);
xor U15366 (N_15366,N_11205,N_8257);
and U15367 (N_15367,N_7153,N_11293);
xor U15368 (N_15368,N_9436,N_10357);
nand U15369 (N_15369,N_9377,N_12223);
and U15370 (N_15370,N_7751,N_11362);
nand U15371 (N_15371,N_11151,N_7753);
nand U15372 (N_15372,N_8170,N_10505);
nand U15373 (N_15373,N_7691,N_10400);
or U15374 (N_15374,N_12016,N_6855);
xor U15375 (N_15375,N_7352,N_11853);
nand U15376 (N_15376,N_9852,N_9580);
nor U15377 (N_15377,N_6585,N_11746);
nand U15378 (N_15378,N_10458,N_6541);
nand U15379 (N_15379,N_8021,N_8540);
and U15380 (N_15380,N_8388,N_12049);
xnor U15381 (N_15381,N_10547,N_6392);
xor U15382 (N_15382,N_10532,N_8463);
or U15383 (N_15383,N_9455,N_8217);
and U15384 (N_15384,N_8929,N_7145);
or U15385 (N_15385,N_9149,N_10325);
or U15386 (N_15386,N_11824,N_9334);
nor U15387 (N_15387,N_10880,N_8949);
nor U15388 (N_15388,N_7639,N_10863);
nor U15389 (N_15389,N_6307,N_7840);
or U15390 (N_15390,N_6499,N_7097);
and U15391 (N_15391,N_8226,N_10187);
nor U15392 (N_15392,N_10470,N_8068);
nand U15393 (N_15393,N_9730,N_6926);
xor U15394 (N_15394,N_6840,N_8085);
xor U15395 (N_15395,N_10162,N_12115);
nand U15396 (N_15396,N_9639,N_7556);
xor U15397 (N_15397,N_9174,N_10751);
and U15398 (N_15398,N_10230,N_9810);
and U15399 (N_15399,N_8800,N_12222);
xnor U15400 (N_15400,N_7386,N_8543);
and U15401 (N_15401,N_9250,N_9225);
and U15402 (N_15402,N_6811,N_11579);
or U15403 (N_15403,N_10647,N_6908);
or U15404 (N_15404,N_8325,N_12492);
nand U15405 (N_15405,N_11516,N_7943);
nor U15406 (N_15406,N_10882,N_9844);
xor U15407 (N_15407,N_7492,N_8007);
xnor U15408 (N_15408,N_11867,N_10709);
nand U15409 (N_15409,N_9799,N_9097);
and U15410 (N_15410,N_8441,N_10206);
or U15411 (N_15411,N_11123,N_9322);
nor U15412 (N_15412,N_8184,N_11367);
nand U15413 (N_15413,N_12323,N_9691);
nor U15414 (N_15414,N_9836,N_6861);
nand U15415 (N_15415,N_6465,N_11996);
nor U15416 (N_15416,N_7437,N_7013);
xnor U15417 (N_15417,N_6421,N_10748);
xnor U15418 (N_15418,N_10572,N_9930);
nor U15419 (N_15419,N_9651,N_10603);
and U15420 (N_15420,N_10821,N_11146);
or U15421 (N_15421,N_10232,N_11661);
xor U15422 (N_15422,N_6959,N_8827);
xnor U15423 (N_15423,N_6379,N_11686);
or U15424 (N_15424,N_11166,N_12484);
and U15425 (N_15425,N_10627,N_8875);
xnor U15426 (N_15426,N_8895,N_8908);
nand U15427 (N_15427,N_9198,N_9044);
nor U15428 (N_15428,N_12493,N_9344);
or U15429 (N_15429,N_11278,N_11852);
and U15430 (N_15430,N_8433,N_7055);
xor U15431 (N_15431,N_10456,N_6752);
or U15432 (N_15432,N_6489,N_11797);
and U15433 (N_15433,N_7431,N_8979);
and U15434 (N_15434,N_6380,N_8874);
nor U15435 (N_15435,N_11125,N_6784);
and U15436 (N_15436,N_8515,N_10319);
nor U15437 (N_15437,N_6358,N_10829);
nand U15438 (N_15438,N_12110,N_7239);
and U15439 (N_15439,N_10119,N_8656);
or U15440 (N_15440,N_11206,N_8528);
xnor U15441 (N_15441,N_12111,N_8458);
nor U15442 (N_15442,N_10023,N_12459);
or U15443 (N_15443,N_10728,N_9742);
xor U15444 (N_15444,N_7366,N_9623);
or U15445 (N_15445,N_12317,N_11212);
xnor U15446 (N_15446,N_8984,N_8904);
nand U15447 (N_15447,N_6484,N_9655);
nor U15448 (N_15448,N_10186,N_11143);
and U15449 (N_15449,N_10936,N_6668);
nand U15450 (N_15450,N_7318,N_11921);
nand U15451 (N_15451,N_10912,N_8720);
xor U15452 (N_15452,N_9222,N_7323);
nor U15453 (N_15453,N_7925,N_6386);
and U15454 (N_15454,N_7337,N_8751);
or U15455 (N_15455,N_7676,N_9568);
nand U15456 (N_15456,N_6685,N_7491);
nor U15457 (N_15457,N_11658,N_11650);
or U15458 (N_15458,N_6615,N_11082);
nor U15459 (N_15459,N_9492,N_7105);
xor U15460 (N_15460,N_8397,N_7150);
nand U15461 (N_15461,N_10784,N_11087);
nand U15462 (N_15462,N_11538,N_9658);
and U15463 (N_15463,N_7061,N_7251);
xnor U15464 (N_15464,N_6680,N_8616);
nand U15465 (N_15465,N_12333,N_7615);
or U15466 (N_15466,N_7488,N_7009);
xor U15467 (N_15467,N_10548,N_9574);
nand U15468 (N_15468,N_7260,N_7174);
nand U15469 (N_15469,N_7357,N_11485);
nor U15470 (N_15470,N_8838,N_8442);
xnor U15471 (N_15471,N_9994,N_8008);
and U15472 (N_15472,N_9242,N_7493);
nand U15473 (N_15473,N_7518,N_7725);
and U15474 (N_15474,N_11086,N_9325);
xnor U15475 (N_15475,N_9056,N_7630);
or U15476 (N_15476,N_9965,N_8797);
or U15477 (N_15477,N_8213,N_12241);
and U15478 (N_15478,N_7461,N_8013);
nor U15479 (N_15479,N_11462,N_6523);
xor U15480 (N_15480,N_8537,N_6391);
or U15481 (N_15481,N_9459,N_10624);
xnor U15482 (N_15482,N_11515,N_7136);
and U15483 (N_15483,N_8144,N_10378);
and U15484 (N_15484,N_8954,N_9807);
xor U15485 (N_15485,N_8502,N_11172);
nand U15486 (N_15486,N_6571,N_7647);
xor U15487 (N_15487,N_10079,N_11432);
or U15488 (N_15488,N_8987,N_9715);
xnor U15489 (N_15489,N_7421,N_6319);
nand U15490 (N_15490,N_10070,N_8197);
xnor U15491 (N_15491,N_10030,N_6750);
nand U15492 (N_15492,N_9442,N_6914);
and U15493 (N_15493,N_10934,N_10861);
or U15494 (N_15494,N_7445,N_12378);
or U15495 (N_15495,N_7021,N_7184);
xnor U15496 (N_15496,N_10461,N_11849);
xor U15497 (N_15497,N_8273,N_8386);
or U15498 (N_15498,N_12271,N_6526);
nor U15499 (N_15499,N_9457,N_8146);
xnor U15500 (N_15500,N_7382,N_12006);
xnor U15501 (N_15501,N_8778,N_9753);
nor U15502 (N_15502,N_11072,N_10370);
xnor U15503 (N_15503,N_6631,N_8791);
nand U15504 (N_15504,N_11772,N_10957);
nor U15505 (N_15505,N_9100,N_7344);
nand U15506 (N_15506,N_6955,N_11458);
or U15507 (N_15507,N_9032,N_8748);
nand U15508 (N_15508,N_7065,N_6849);
and U15509 (N_15509,N_8728,N_6761);
and U15510 (N_15510,N_11677,N_8694);
and U15511 (N_15511,N_10764,N_9296);
nor U15512 (N_15512,N_10156,N_12308);
and U15513 (N_15513,N_10404,N_11022);
or U15514 (N_15514,N_11263,N_9390);
xor U15515 (N_15515,N_9627,N_8103);
or U15516 (N_15516,N_9464,N_9678);
xnor U15517 (N_15517,N_6627,N_10035);
nor U15518 (N_15518,N_9435,N_10176);
nor U15519 (N_15519,N_7018,N_8826);
nor U15520 (N_15520,N_7208,N_10080);
nor U15521 (N_15521,N_10592,N_8212);
nor U15522 (N_15522,N_8530,N_9661);
nand U15523 (N_15523,N_11729,N_10913);
and U15524 (N_15524,N_11906,N_11869);
nand U15525 (N_15525,N_10995,N_7311);
or U15526 (N_15526,N_7316,N_9713);
nor U15527 (N_15527,N_10045,N_7600);
or U15528 (N_15528,N_6777,N_12415);
nand U15529 (N_15529,N_8880,N_9913);
nor U15530 (N_15530,N_8750,N_8320);
nand U15531 (N_15531,N_9115,N_9756);
nor U15532 (N_15532,N_7734,N_8834);
and U15533 (N_15533,N_7375,N_11877);
and U15534 (N_15534,N_10641,N_9600);
nand U15535 (N_15535,N_11433,N_7827);
xor U15536 (N_15536,N_11085,N_9438);
or U15537 (N_15537,N_6672,N_10441);
and U15538 (N_15538,N_8088,N_7774);
or U15539 (N_15539,N_6868,N_9413);
nand U15540 (N_15540,N_10197,N_7462);
nor U15541 (N_15541,N_8039,N_6694);
nand U15542 (N_15542,N_10324,N_6872);
nand U15543 (N_15543,N_8286,N_11041);
nor U15544 (N_15544,N_8304,N_9134);
or U15545 (N_15545,N_11388,N_7263);
xor U15546 (N_15546,N_10135,N_10642);
nor U15547 (N_15547,N_12248,N_9883);
nand U15548 (N_15548,N_8362,N_6951);
or U15549 (N_15549,N_10566,N_9017);
nand U15550 (N_15550,N_8985,N_8652);
xor U15551 (N_15551,N_9158,N_8330);
nand U15552 (N_15552,N_8901,N_8894);
and U15553 (N_15553,N_10032,N_9766);
and U15554 (N_15554,N_8360,N_11221);
and U15555 (N_15555,N_11886,N_10256);
nor U15556 (N_15556,N_6289,N_12402);
or U15557 (N_15557,N_6312,N_11683);
nor U15558 (N_15558,N_7788,N_7086);
nand U15559 (N_15559,N_8006,N_10608);
nor U15560 (N_15560,N_11803,N_9279);
nor U15561 (N_15561,N_11449,N_8889);
xor U15562 (N_15562,N_9612,N_9780);
and U15563 (N_15563,N_12166,N_11533);
xnor U15564 (N_15564,N_9595,N_9321);
nor U15565 (N_15565,N_7515,N_8676);
and U15566 (N_15566,N_11503,N_11239);
xor U15567 (N_15567,N_11256,N_9212);
xnor U15568 (N_15568,N_6681,N_9499);
nor U15569 (N_15569,N_6719,N_6982);
or U15570 (N_15570,N_8370,N_11675);
nand U15571 (N_15571,N_10508,N_7966);
nand U15572 (N_15572,N_11986,N_7951);
nor U15573 (N_15573,N_7130,N_6801);
nor U15574 (N_15574,N_11528,N_6783);
xnor U15575 (N_15575,N_12109,N_7762);
xor U15576 (N_15576,N_10577,N_12322);
nand U15577 (N_15577,N_8497,N_8602);
or U15578 (N_15578,N_10582,N_12462);
nand U15579 (N_15579,N_12076,N_11691);
or U15580 (N_15580,N_11641,N_6547);
and U15581 (N_15581,N_12251,N_6666);
or U15582 (N_15582,N_6873,N_8156);
and U15583 (N_15583,N_9763,N_9146);
and U15584 (N_15584,N_11711,N_7905);
xnor U15585 (N_15585,N_10815,N_8747);
nand U15586 (N_15586,N_10814,N_8254);
nand U15587 (N_15587,N_7802,N_7069);
nand U15588 (N_15588,N_10407,N_11188);
or U15589 (N_15589,N_9195,N_12288);
xor U15590 (N_15590,N_12444,N_8138);
xnor U15591 (N_15591,N_6263,N_12001);
and U15592 (N_15592,N_8250,N_7974);
nand U15593 (N_15593,N_7505,N_7722);
nor U15594 (N_15594,N_8311,N_10956);
and U15595 (N_15595,N_6385,N_11336);
nand U15596 (N_15596,N_6493,N_7285);
xnor U15597 (N_15597,N_10281,N_12021);
xnor U15598 (N_15598,N_11294,N_9368);
nor U15599 (N_15599,N_9554,N_10348);
or U15600 (N_15600,N_7090,N_9135);
and U15601 (N_15601,N_11314,N_9922);
or U15602 (N_15602,N_10464,N_10012);
nor U15603 (N_15603,N_11017,N_12418);
nand U15604 (N_15604,N_6897,N_10809);
xor U15605 (N_15605,N_10786,N_8140);
nand U15606 (N_15606,N_7225,N_10104);
xnor U15607 (N_15607,N_8861,N_9509);
or U15608 (N_15608,N_6931,N_11057);
xnor U15609 (N_15609,N_9352,N_10369);
xnor U15610 (N_15610,N_8547,N_10741);
nor U15611 (N_15611,N_9700,N_12429);
nand U15612 (N_15612,N_11723,N_8410);
nand U15613 (N_15613,N_12403,N_12053);
or U15614 (N_15614,N_11495,N_9020);
and U15615 (N_15615,N_8072,N_7752);
and U15616 (N_15616,N_6804,N_11334);
nand U15617 (N_15617,N_6664,N_11076);
nand U15618 (N_15618,N_12435,N_11504);
and U15619 (N_15619,N_7211,N_9601);
xnor U15620 (N_15620,N_10426,N_9588);
and U15621 (N_15621,N_8157,N_11324);
nand U15622 (N_15622,N_11117,N_7332);
nor U15623 (N_15623,N_10613,N_9290);
nand U15624 (N_15624,N_11889,N_10734);
or U15625 (N_15625,N_6890,N_6781);
nand U15626 (N_15626,N_9046,N_10757);
or U15627 (N_15627,N_9972,N_10231);
nand U15628 (N_15628,N_7803,N_7136);
nand U15629 (N_15629,N_8622,N_9567);
nor U15630 (N_15630,N_8250,N_10371);
or U15631 (N_15631,N_12240,N_8239);
nor U15632 (N_15632,N_8365,N_7843);
or U15633 (N_15633,N_6739,N_10323);
and U15634 (N_15634,N_6285,N_10088);
and U15635 (N_15635,N_10205,N_11249);
or U15636 (N_15636,N_10822,N_10009);
nor U15637 (N_15637,N_8573,N_10874);
nor U15638 (N_15638,N_12224,N_6546);
nand U15639 (N_15639,N_8761,N_9592);
xor U15640 (N_15640,N_9432,N_7777);
xor U15641 (N_15641,N_9991,N_8371);
and U15642 (N_15642,N_7879,N_11174);
nand U15643 (N_15643,N_9023,N_9784);
and U15644 (N_15644,N_10856,N_6970);
nor U15645 (N_15645,N_12198,N_7599);
or U15646 (N_15646,N_7772,N_9916);
nor U15647 (N_15647,N_7261,N_10410);
or U15648 (N_15648,N_10694,N_7791);
nor U15649 (N_15649,N_10594,N_10235);
nor U15650 (N_15650,N_11692,N_11664);
nor U15651 (N_15651,N_10680,N_8406);
and U15652 (N_15652,N_11792,N_9354);
or U15653 (N_15653,N_8599,N_7167);
and U15654 (N_15654,N_10734,N_8397);
or U15655 (N_15655,N_8355,N_9388);
and U15656 (N_15656,N_9547,N_9766);
nor U15657 (N_15657,N_6373,N_7672);
or U15658 (N_15658,N_8702,N_10444);
nand U15659 (N_15659,N_7366,N_8555);
xnor U15660 (N_15660,N_12370,N_9875);
and U15661 (N_15661,N_7934,N_8778);
or U15662 (N_15662,N_7588,N_11806);
nor U15663 (N_15663,N_7224,N_9819);
xor U15664 (N_15664,N_7096,N_9165);
xor U15665 (N_15665,N_10087,N_7519);
or U15666 (N_15666,N_6471,N_12206);
nand U15667 (N_15667,N_10476,N_6434);
nand U15668 (N_15668,N_9041,N_6879);
nand U15669 (N_15669,N_9087,N_11198);
nor U15670 (N_15670,N_8842,N_10938);
or U15671 (N_15671,N_8636,N_8358);
and U15672 (N_15672,N_10639,N_7453);
and U15673 (N_15673,N_9619,N_12229);
and U15674 (N_15674,N_11036,N_7430);
nand U15675 (N_15675,N_10473,N_10292);
xnor U15676 (N_15676,N_12071,N_12253);
nor U15677 (N_15677,N_11025,N_9808);
nand U15678 (N_15678,N_12014,N_8038);
or U15679 (N_15679,N_6530,N_11616);
xnor U15680 (N_15680,N_10584,N_10359);
nor U15681 (N_15681,N_10075,N_8964);
xnor U15682 (N_15682,N_8925,N_10738);
xor U15683 (N_15683,N_11734,N_8608);
or U15684 (N_15684,N_7183,N_8976);
and U15685 (N_15685,N_9240,N_10609);
or U15686 (N_15686,N_12322,N_9947);
or U15687 (N_15687,N_7284,N_11741);
or U15688 (N_15688,N_11881,N_8623);
or U15689 (N_15689,N_7839,N_12496);
nand U15690 (N_15690,N_8852,N_12140);
nand U15691 (N_15691,N_6453,N_10085);
nor U15692 (N_15692,N_10098,N_11689);
xnor U15693 (N_15693,N_6425,N_10764);
xnor U15694 (N_15694,N_6870,N_7156);
nand U15695 (N_15695,N_11964,N_10276);
xnor U15696 (N_15696,N_6433,N_12137);
xor U15697 (N_15697,N_9013,N_9702);
and U15698 (N_15698,N_7778,N_11568);
nor U15699 (N_15699,N_10700,N_8484);
xnor U15700 (N_15700,N_8949,N_7390);
and U15701 (N_15701,N_7384,N_11535);
and U15702 (N_15702,N_7038,N_8161);
nor U15703 (N_15703,N_9798,N_11270);
or U15704 (N_15704,N_6764,N_8282);
and U15705 (N_15705,N_11320,N_11587);
or U15706 (N_15706,N_9993,N_8591);
nor U15707 (N_15707,N_9982,N_8087);
xnor U15708 (N_15708,N_12332,N_8932);
or U15709 (N_15709,N_11034,N_11935);
or U15710 (N_15710,N_6501,N_11675);
xor U15711 (N_15711,N_6918,N_6263);
nor U15712 (N_15712,N_10690,N_10706);
and U15713 (N_15713,N_12479,N_6827);
nand U15714 (N_15714,N_7120,N_10189);
or U15715 (N_15715,N_6298,N_9010);
or U15716 (N_15716,N_7677,N_9140);
nand U15717 (N_15717,N_8854,N_6813);
or U15718 (N_15718,N_11172,N_11330);
xnor U15719 (N_15719,N_9475,N_7016);
nand U15720 (N_15720,N_11659,N_10340);
or U15721 (N_15721,N_6882,N_6801);
and U15722 (N_15722,N_10993,N_7273);
xnor U15723 (N_15723,N_6818,N_10491);
xnor U15724 (N_15724,N_9590,N_9771);
or U15725 (N_15725,N_7589,N_10666);
xnor U15726 (N_15726,N_6941,N_11697);
nand U15727 (N_15727,N_8581,N_9831);
xor U15728 (N_15728,N_12125,N_7281);
or U15729 (N_15729,N_6879,N_8155);
or U15730 (N_15730,N_7422,N_10568);
or U15731 (N_15731,N_10211,N_11809);
or U15732 (N_15732,N_9605,N_7370);
nor U15733 (N_15733,N_10242,N_10641);
nand U15734 (N_15734,N_6924,N_11824);
and U15735 (N_15735,N_9466,N_7351);
nor U15736 (N_15736,N_10419,N_11687);
nand U15737 (N_15737,N_11710,N_6322);
nor U15738 (N_15738,N_7545,N_7846);
xnor U15739 (N_15739,N_11479,N_6975);
nor U15740 (N_15740,N_7169,N_12144);
xor U15741 (N_15741,N_10826,N_6909);
nor U15742 (N_15742,N_10116,N_8719);
xnor U15743 (N_15743,N_10745,N_10681);
nor U15744 (N_15744,N_8600,N_11544);
xor U15745 (N_15745,N_9106,N_6259);
and U15746 (N_15746,N_8696,N_9406);
xnor U15747 (N_15747,N_12084,N_12315);
and U15748 (N_15748,N_10888,N_7905);
and U15749 (N_15749,N_7537,N_8211);
nand U15750 (N_15750,N_6252,N_12322);
xor U15751 (N_15751,N_10236,N_12458);
or U15752 (N_15752,N_8244,N_9608);
or U15753 (N_15753,N_10738,N_11997);
and U15754 (N_15754,N_7905,N_10120);
or U15755 (N_15755,N_7839,N_8965);
nand U15756 (N_15756,N_8029,N_8117);
or U15757 (N_15757,N_7954,N_11647);
or U15758 (N_15758,N_6423,N_11093);
xor U15759 (N_15759,N_10567,N_10293);
nand U15760 (N_15760,N_7672,N_6951);
xor U15761 (N_15761,N_11442,N_10900);
nand U15762 (N_15762,N_11004,N_8357);
nor U15763 (N_15763,N_9526,N_12343);
and U15764 (N_15764,N_8644,N_9954);
nor U15765 (N_15765,N_11492,N_6613);
or U15766 (N_15766,N_10916,N_6331);
nor U15767 (N_15767,N_9692,N_11769);
xor U15768 (N_15768,N_9294,N_11735);
and U15769 (N_15769,N_11011,N_8333);
and U15770 (N_15770,N_9997,N_10330);
nand U15771 (N_15771,N_7169,N_11607);
or U15772 (N_15772,N_9439,N_12159);
or U15773 (N_15773,N_12312,N_10248);
nand U15774 (N_15774,N_12207,N_12492);
xor U15775 (N_15775,N_12094,N_11438);
xnor U15776 (N_15776,N_10262,N_7212);
nand U15777 (N_15777,N_11631,N_6346);
nor U15778 (N_15778,N_11599,N_9673);
and U15779 (N_15779,N_10938,N_7054);
and U15780 (N_15780,N_7423,N_8247);
xnor U15781 (N_15781,N_7029,N_10936);
xnor U15782 (N_15782,N_9170,N_12166);
nand U15783 (N_15783,N_10912,N_10165);
xnor U15784 (N_15784,N_10421,N_11259);
or U15785 (N_15785,N_7502,N_10749);
nand U15786 (N_15786,N_11349,N_7408);
nor U15787 (N_15787,N_7512,N_10635);
nand U15788 (N_15788,N_12111,N_8114);
nand U15789 (N_15789,N_8663,N_7354);
and U15790 (N_15790,N_10479,N_6787);
xnor U15791 (N_15791,N_10479,N_9112);
xnor U15792 (N_15792,N_8960,N_8720);
nor U15793 (N_15793,N_9901,N_10123);
xor U15794 (N_15794,N_8628,N_8383);
and U15795 (N_15795,N_10998,N_11233);
or U15796 (N_15796,N_8667,N_11352);
and U15797 (N_15797,N_6930,N_8907);
and U15798 (N_15798,N_8904,N_7204);
xnor U15799 (N_15799,N_11442,N_11093);
xnor U15800 (N_15800,N_8682,N_9074);
nand U15801 (N_15801,N_8900,N_8157);
nand U15802 (N_15802,N_8528,N_9772);
and U15803 (N_15803,N_10264,N_7807);
and U15804 (N_15804,N_6798,N_7585);
or U15805 (N_15805,N_6876,N_10150);
nand U15806 (N_15806,N_9077,N_8424);
and U15807 (N_15807,N_8346,N_10564);
nor U15808 (N_15808,N_7246,N_12064);
nand U15809 (N_15809,N_11158,N_12288);
or U15810 (N_15810,N_7745,N_11462);
nand U15811 (N_15811,N_10972,N_9069);
nor U15812 (N_15812,N_6849,N_9385);
nor U15813 (N_15813,N_6686,N_8533);
or U15814 (N_15814,N_8216,N_11916);
nand U15815 (N_15815,N_9113,N_9659);
and U15816 (N_15816,N_9869,N_7839);
xnor U15817 (N_15817,N_11521,N_6656);
or U15818 (N_15818,N_8306,N_6919);
nor U15819 (N_15819,N_11518,N_8658);
xnor U15820 (N_15820,N_11572,N_8578);
nand U15821 (N_15821,N_10936,N_8858);
nand U15822 (N_15822,N_12224,N_7895);
nand U15823 (N_15823,N_8769,N_10645);
and U15824 (N_15824,N_9433,N_9269);
xnor U15825 (N_15825,N_6378,N_9406);
or U15826 (N_15826,N_12209,N_7089);
xnor U15827 (N_15827,N_9472,N_7904);
and U15828 (N_15828,N_8079,N_9486);
and U15829 (N_15829,N_7696,N_10762);
nor U15830 (N_15830,N_11142,N_9323);
nor U15831 (N_15831,N_6945,N_12220);
nor U15832 (N_15832,N_10063,N_12067);
or U15833 (N_15833,N_7633,N_8756);
nor U15834 (N_15834,N_9759,N_10858);
or U15835 (N_15835,N_7746,N_12355);
xnor U15836 (N_15836,N_10259,N_12330);
and U15837 (N_15837,N_10383,N_10001);
xor U15838 (N_15838,N_7752,N_8045);
nand U15839 (N_15839,N_12125,N_6932);
nor U15840 (N_15840,N_11180,N_10367);
nand U15841 (N_15841,N_11279,N_6384);
nand U15842 (N_15842,N_6526,N_11217);
nor U15843 (N_15843,N_10419,N_6422);
and U15844 (N_15844,N_11170,N_7448);
and U15845 (N_15845,N_10005,N_11716);
nand U15846 (N_15846,N_7415,N_11284);
and U15847 (N_15847,N_6859,N_12378);
and U15848 (N_15848,N_8503,N_9153);
or U15849 (N_15849,N_11103,N_10291);
nand U15850 (N_15850,N_11057,N_8009);
xnor U15851 (N_15851,N_7256,N_10031);
xnor U15852 (N_15852,N_12336,N_12089);
or U15853 (N_15853,N_8706,N_12230);
xnor U15854 (N_15854,N_6358,N_9123);
xnor U15855 (N_15855,N_11758,N_11804);
or U15856 (N_15856,N_8268,N_9600);
nor U15857 (N_15857,N_7683,N_11070);
xnor U15858 (N_15858,N_11200,N_11397);
nor U15859 (N_15859,N_9402,N_9080);
nor U15860 (N_15860,N_8680,N_9106);
xor U15861 (N_15861,N_12387,N_12205);
nand U15862 (N_15862,N_6554,N_9298);
nand U15863 (N_15863,N_12148,N_9828);
and U15864 (N_15864,N_8797,N_11205);
nand U15865 (N_15865,N_9578,N_9611);
xnor U15866 (N_15866,N_9539,N_7831);
nand U15867 (N_15867,N_7237,N_9952);
or U15868 (N_15868,N_6431,N_6898);
and U15869 (N_15869,N_6648,N_12289);
nor U15870 (N_15870,N_7104,N_11426);
nor U15871 (N_15871,N_9125,N_11865);
xor U15872 (N_15872,N_7920,N_11852);
or U15873 (N_15873,N_10586,N_7783);
nor U15874 (N_15874,N_9869,N_11954);
and U15875 (N_15875,N_10789,N_8577);
nand U15876 (N_15876,N_10485,N_10478);
and U15877 (N_15877,N_11912,N_8582);
nand U15878 (N_15878,N_10015,N_9707);
nand U15879 (N_15879,N_11225,N_9938);
xnor U15880 (N_15880,N_10657,N_9519);
or U15881 (N_15881,N_6339,N_8882);
or U15882 (N_15882,N_11450,N_8895);
nor U15883 (N_15883,N_7993,N_9476);
nand U15884 (N_15884,N_6307,N_7313);
nand U15885 (N_15885,N_7408,N_8444);
xnor U15886 (N_15886,N_11419,N_8145);
or U15887 (N_15887,N_7362,N_11653);
and U15888 (N_15888,N_10918,N_10590);
or U15889 (N_15889,N_7432,N_6261);
nor U15890 (N_15890,N_7940,N_12095);
and U15891 (N_15891,N_10363,N_8824);
xnor U15892 (N_15892,N_6309,N_8680);
and U15893 (N_15893,N_10027,N_11476);
and U15894 (N_15894,N_7234,N_9488);
and U15895 (N_15895,N_6415,N_6761);
and U15896 (N_15896,N_11245,N_7048);
or U15897 (N_15897,N_6486,N_11972);
or U15898 (N_15898,N_8032,N_11600);
nor U15899 (N_15899,N_7657,N_12204);
and U15900 (N_15900,N_7788,N_8161);
xor U15901 (N_15901,N_7148,N_7440);
and U15902 (N_15902,N_6441,N_11511);
xor U15903 (N_15903,N_10182,N_10029);
nand U15904 (N_15904,N_8376,N_10432);
nor U15905 (N_15905,N_11964,N_12294);
nor U15906 (N_15906,N_10528,N_10900);
or U15907 (N_15907,N_8091,N_8816);
and U15908 (N_15908,N_7563,N_6724);
nor U15909 (N_15909,N_11980,N_11734);
nand U15910 (N_15910,N_10641,N_9772);
nor U15911 (N_15911,N_7074,N_6301);
nor U15912 (N_15912,N_7349,N_12040);
nand U15913 (N_15913,N_10598,N_9082);
nand U15914 (N_15914,N_10508,N_12179);
nand U15915 (N_15915,N_11973,N_10350);
or U15916 (N_15916,N_7508,N_8978);
nor U15917 (N_15917,N_8010,N_11722);
and U15918 (N_15918,N_11165,N_11291);
xor U15919 (N_15919,N_9785,N_7742);
nor U15920 (N_15920,N_8967,N_12076);
and U15921 (N_15921,N_7147,N_12382);
or U15922 (N_15922,N_8126,N_9898);
nand U15923 (N_15923,N_10098,N_11819);
and U15924 (N_15924,N_12009,N_10647);
or U15925 (N_15925,N_6892,N_8178);
and U15926 (N_15926,N_12004,N_10057);
and U15927 (N_15927,N_7104,N_7817);
and U15928 (N_15928,N_11424,N_11988);
nand U15929 (N_15929,N_7151,N_10151);
or U15930 (N_15930,N_11796,N_12368);
or U15931 (N_15931,N_8330,N_11679);
xnor U15932 (N_15932,N_8580,N_8660);
nand U15933 (N_15933,N_7016,N_12181);
xor U15934 (N_15934,N_6996,N_11126);
nand U15935 (N_15935,N_6345,N_11519);
nor U15936 (N_15936,N_11004,N_6691);
or U15937 (N_15937,N_6718,N_7177);
nand U15938 (N_15938,N_10777,N_11854);
nor U15939 (N_15939,N_8782,N_12253);
xnor U15940 (N_15940,N_9276,N_9643);
nor U15941 (N_15941,N_8680,N_9155);
nor U15942 (N_15942,N_9824,N_10708);
and U15943 (N_15943,N_10160,N_10800);
xor U15944 (N_15944,N_7287,N_11598);
nor U15945 (N_15945,N_7235,N_11025);
nor U15946 (N_15946,N_12273,N_10620);
xnor U15947 (N_15947,N_9603,N_8323);
nor U15948 (N_15948,N_12071,N_8551);
nand U15949 (N_15949,N_6940,N_9987);
or U15950 (N_15950,N_10145,N_6629);
xnor U15951 (N_15951,N_7957,N_11122);
or U15952 (N_15952,N_10269,N_6565);
or U15953 (N_15953,N_11368,N_11001);
or U15954 (N_15954,N_7034,N_8440);
and U15955 (N_15955,N_7625,N_9592);
nor U15956 (N_15956,N_8831,N_9306);
nor U15957 (N_15957,N_8940,N_11601);
nor U15958 (N_15958,N_10901,N_8133);
xor U15959 (N_15959,N_9746,N_8430);
or U15960 (N_15960,N_10065,N_10943);
and U15961 (N_15961,N_11650,N_10865);
or U15962 (N_15962,N_11236,N_9048);
or U15963 (N_15963,N_8193,N_6876);
xnor U15964 (N_15964,N_11088,N_10487);
xor U15965 (N_15965,N_10726,N_12269);
nand U15966 (N_15966,N_7505,N_8840);
and U15967 (N_15967,N_11889,N_11733);
nand U15968 (N_15968,N_9006,N_9076);
or U15969 (N_15969,N_9068,N_7379);
nor U15970 (N_15970,N_12478,N_9589);
nand U15971 (N_15971,N_9556,N_9567);
or U15972 (N_15972,N_7522,N_8858);
xnor U15973 (N_15973,N_9734,N_11109);
and U15974 (N_15974,N_8985,N_10384);
nor U15975 (N_15975,N_7655,N_8764);
or U15976 (N_15976,N_11538,N_8776);
or U15977 (N_15977,N_9990,N_10687);
nand U15978 (N_15978,N_7220,N_10588);
or U15979 (N_15979,N_9169,N_7467);
or U15980 (N_15980,N_8186,N_6336);
xor U15981 (N_15981,N_9660,N_11288);
or U15982 (N_15982,N_11918,N_8369);
nor U15983 (N_15983,N_10103,N_8760);
and U15984 (N_15984,N_8427,N_6751);
nor U15985 (N_15985,N_11640,N_11381);
nand U15986 (N_15986,N_7074,N_7688);
xnor U15987 (N_15987,N_10941,N_9115);
nor U15988 (N_15988,N_7438,N_10587);
nand U15989 (N_15989,N_8577,N_11813);
nor U15990 (N_15990,N_12279,N_11892);
nor U15991 (N_15991,N_7833,N_7086);
xnor U15992 (N_15992,N_9976,N_6940);
and U15993 (N_15993,N_10854,N_12191);
nand U15994 (N_15994,N_7845,N_11530);
nor U15995 (N_15995,N_12488,N_11504);
and U15996 (N_15996,N_12206,N_11628);
xor U15997 (N_15997,N_10132,N_7932);
xnor U15998 (N_15998,N_6823,N_7252);
or U15999 (N_15999,N_11675,N_7158);
nor U16000 (N_16000,N_9582,N_9729);
and U16001 (N_16001,N_10280,N_7712);
xor U16002 (N_16002,N_11904,N_11681);
xor U16003 (N_16003,N_9874,N_7491);
nor U16004 (N_16004,N_10338,N_10459);
or U16005 (N_16005,N_12151,N_9582);
nor U16006 (N_16006,N_7376,N_11581);
and U16007 (N_16007,N_7208,N_10146);
and U16008 (N_16008,N_12403,N_9114);
and U16009 (N_16009,N_7670,N_8792);
nor U16010 (N_16010,N_11385,N_6316);
nor U16011 (N_16011,N_11733,N_11547);
nand U16012 (N_16012,N_6440,N_12408);
nor U16013 (N_16013,N_6651,N_9058);
xor U16014 (N_16014,N_10326,N_7988);
nor U16015 (N_16015,N_11358,N_10034);
nand U16016 (N_16016,N_10898,N_7427);
or U16017 (N_16017,N_6435,N_8576);
xnor U16018 (N_16018,N_9777,N_10479);
or U16019 (N_16019,N_11304,N_8295);
nand U16020 (N_16020,N_6516,N_10520);
or U16021 (N_16021,N_8281,N_11801);
nor U16022 (N_16022,N_8035,N_7108);
and U16023 (N_16023,N_6405,N_6477);
and U16024 (N_16024,N_10619,N_12393);
nand U16025 (N_16025,N_7469,N_7765);
nand U16026 (N_16026,N_9982,N_9570);
nor U16027 (N_16027,N_12295,N_8002);
xor U16028 (N_16028,N_11942,N_8452);
or U16029 (N_16029,N_9271,N_11263);
and U16030 (N_16030,N_9535,N_7501);
or U16031 (N_16031,N_10700,N_9860);
xnor U16032 (N_16032,N_7747,N_8084);
xor U16033 (N_16033,N_8610,N_9730);
or U16034 (N_16034,N_7919,N_7674);
nor U16035 (N_16035,N_12053,N_11057);
xnor U16036 (N_16036,N_10854,N_12075);
nand U16037 (N_16037,N_7497,N_9066);
xnor U16038 (N_16038,N_7972,N_11349);
or U16039 (N_16039,N_6711,N_6493);
or U16040 (N_16040,N_6864,N_7681);
or U16041 (N_16041,N_6740,N_11340);
xnor U16042 (N_16042,N_10698,N_7644);
and U16043 (N_16043,N_10264,N_8979);
and U16044 (N_16044,N_7568,N_7057);
and U16045 (N_16045,N_12359,N_7911);
xnor U16046 (N_16046,N_9516,N_10767);
nand U16047 (N_16047,N_12469,N_10239);
or U16048 (N_16048,N_10274,N_6929);
nand U16049 (N_16049,N_8512,N_7473);
xor U16050 (N_16050,N_7888,N_7929);
nand U16051 (N_16051,N_10244,N_8392);
nor U16052 (N_16052,N_10662,N_7024);
or U16053 (N_16053,N_8477,N_9891);
xnor U16054 (N_16054,N_7214,N_10456);
or U16055 (N_16055,N_8182,N_9407);
or U16056 (N_16056,N_9976,N_7800);
nand U16057 (N_16057,N_8515,N_12084);
nand U16058 (N_16058,N_6600,N_8629);
xnor U16059 (N_16059,N_10324,N_12128);
and U16060 (N_16060,N_8113,N_8024);
nor U16061 (N_16061,N_6325,N_11560);
or U16062 (N_16062,N_9994,N_10562);
nand U16063 (N_16063,N_9960,N_6699);
and U16064 (N_16064,N_10213,N_7139);
xor U16065 (N_16065,N_8953,N_8286);
nand U16066 (N_16066,N_7466,N_8583);
xnor U16067 (N_16067,N_8399,N_6522);
xnor U16068 (N_16068,N_8541,N_12290);
and U16069 (N_16069,N_9847,N_11872);
and U16070 (N_16070,N_11752,N_9902);
xnor U16071 (N_16071,N_9625,N_7588);
xnor U16072 (N_16072,N_7970,N_9285);
nor U16073 (N_16073,N_11262,N_10548);
nand U16074 (N_16074,N_7549,N_8680);
nor U16075 (N_16075,N_9651,N_11489);
and U16076 (N_16076,N_6525,N_8555);
nor U16077 (N_16077,N_11000,N_11267);
nand U16078 (N_16078,N_10620,N_8549);
and U16079 (N_16079,N_12436,N_7626);
and U16080 (N_16080,N_6885,N_9170);
or U16081 (N_16081,N_6995,N_10975);
nand U16082 (N_16082,N_10170,N_6450);
or U16083 (N_16083,N_6441,N_8013);
or U16084 (N_16084,N_9787,N_11036);
nand U16085 (N_16085,N_8027,N_10589);
and U16086 (N_16086,N_11237,N_11739);
and U16087 (N_16087,N_8746,N_11889);
xor U16088 (N_16088,N_6467,N_10282);
or U16089 (N_16089,N_9189,N_12400);
nor U16090 (N_16090,N_9327,N_6421);
nor U16091 (N_16091,N_12414,N_8271);
xnor U16092 (N_16092,N_8951,N_10894);
xnor U16093 (N_16093,N_9008,N_9982);
nor U16094 (N_16094,N_10636,N_10504);
and U16095 (N_16095,N_10771,N_6437);
xnor U16096 (N_16096,N_9511,N_8042);
xnor U16097 (N_16097,N_11790,N_12285);
nor U16098 (N_16098,N_8763,N_9374);
nor U16099 (N_16099,N_11742,N_10325);
nor U16100 (N_16100,N_7633,N_8769);
xnor U16101 (N_16101,N_6592,N_9081);
or U16102 (N_16102,N_10703,N_11984);
or U16103 (N_16103,N_7997,N_9741);
or U16104 (N_16104,N_10571,N_10517);
nand U16105 (N_16105,N_6721,N_6941);
or U16106 (N_16106,N_9117,N_10629);
xor U16107 (N_16107,N_8788,N_10383);
or U16108 (N_16108,N_6382,N_9930);
xor U16109 (N_16109,N_10867,N_11500);
or U16110 (N_16110,N_6711,N_10061);
or U16111 (N_16111,N_12352,N_11038);
or U16112 (N_16112,N_6672,N_12261);
xnor U16113 (N_16113,N_9441,N_11540);
or U16114 (N_16114,N_11421,N_8203);
nand U16115 (N_16115,N_11587,N_7424);
or U16116 (N_16116,N_7875,N_9535);
nor U16117 (N_16117,N_11336,N_9307);
or U16118 (N_16118,N_11375,N_10696);
nor U16119 (N_16119,N_6580,N_12229);
nand U16120 (N_16120,N_11562,N_6961);
or U16121 (N_16121,N_7940,N_7108);
nand U16122 (N_16122,N_10162,N_11926);
nand U16123 (N_16123,N_9876,N_9417);
nor U16124 (N_16124,N_10720,N_8687);
nor U16125 (N_16125,N_12361,N_6929);
or U16126 (N_16126,N_6276,N_10479);
nor U16127 (N_16127,N_9067,N_12405);
xor U16128 (N_16128,N_9748,N_6902);
xnor U16129 (N_16129,N_11062,N_12066);
nand U16130 (N_16130,N_8245,N_12136);
nand U16131 (N_16131,N_8609,N_11351);
nand U16132 (N_16132,N_6373,N_7017);
nor U16133 (N_16133,N_6571,N_8732);
nor U16134 (N_16134,N_11598,N_7883);
or U16135 (N_16135,N_9392,N_9059);
and U16136 (N_16136,N_7558,N_10436);
xor U16137 (N_16137,N_10942,N_8178);
and U16138 (N_16138,N_7880,N_9245);
or U16139 (N_16139,N_10641,N_6976);
and U16140 (N_16140,N_11536,N_9565);
xnor U16141 (N_16141,N_10764,N_12390);
nand U16142 (N_16142,N_11542,N_10592);
and U16143 (N_16143,N_8041,N_12124);
and U16144 (N_16144,N_7776,N_7915);
nor U16145 (N_16145,N_7982,N_8206);
xnor U16146 (N_16146,N_9325,N_7071);
nand U16147 (N_16147,N_8886,N_7557);
nor U16148 (N_16148,N_9475,N_8888);
nand U16149 (N_16149,N_10638,N_10555);
and U16150 (N_16150,N_9814,N_7882);
or U16151 (N_16151,N_8462,N_7402);
or U16152 (N_16152,N_11194,N_9888);
xnor U16153 (N_16153,N_9889,N_9817);
xnor U16154 (N_16154,N_6774,N_12319);
nand U16155 (N_16155,N_11801,N_9032);
and U16156 (N_16156,N_8113,N_8214);
or U16157 (N_16157,N_10222,N_9684);
nor U16158 (N_16158,N_7793,N_7926);
or U16159 (N_16159,N_10862,N_6666);
nand U16160 (N_16160,N_9406,N_10463);
nand U16161 (N_16161,N_8491,N_12166);
nor U16162 (N_16162,N_12478,N_9040);
nor U16163 (N_16163,N_11689,N_6763);
nor U16164 (N_16164,N_9357,N_6809);
nand U16165 (N_16165,N_12325,N_9768);
nor U16166 (N_16166,N_7691,N_7718);
or U16167 (N_16167,N_10474,N_12273);
and U16168 (N_16168,N_10256,N_9891);
nor U16169 (N_16169,N_10270,N_7216);
and U16170 (N_16170,N_11544,N_9199);
nand U16171 (N_16171,N_9195,N_10338);
nor U16172 (N_16172,N_9764,N_11926);
and U16173 (N_16173,N_12040,N_8431);
and U16174 (N_16174,N_10012,N_6430);
nor U16175 (N_16175,N_10352,N_6740);
and U16176 (N_16176,N_11801,N_10916);
xor U16177 (N_16177,N_10696,N_11655);
and U16178 (N_16178,N_7693,N_12264);
xor U16179 (N_16179,N_10953,N_11682);
xor U16180 (N_16180,N_8744,N_8681);
nor U16181 (N_16181,N_11931,N_11155);
xor U16182 (N_16182,N_10020,N_7650);
xnor U16183 (N_16183,N_11151,N_7787);
nor U16184 (N_16184,N_8568,N_7381);
nor U16185 (N_16185,N_12020,N_10994);
nand U16186 (N_16186,N_10357,N_7962);
nand U16187 (N_16187,N_7424,N_8019);
xnor U16188 (N_16188,N_8106,N_9708);
nand U16189 (N_16189,N_12236,N_12329);
nor U16190 (N_16190,N_10183,N_9336);
nor U16191 (N_16191,N_8370,N_6938);
nor U16192 (N_16192,N_8152,N_8300);
or U16193 (N_16193,N_11076,N_12485);
xnor U16194 (N_16194,N_10169,N_7699);
xnor U16195 (N_16195,N_8916,N_9753);
or U16196 (N_16196,N_8745,N_6859);
nor U16197 (N_16197,N_7092,N_11628);
nand U16198 (N_16198,N_9799,N_6400);
xnor U16199 (N_16199,N_9449,N_11547);
nand U16200 (N_16200,N_9609,N_6792);
or U16201 (N_16201,N_12242,N_6410);
or U16202 (N_16202,N_8567,N_9746);
nor U16203 (N_16203,N_6392,N_10812);
or U16204 (N_16204,N_10723,N_9847);
xor U16205 (N_16205,N_10236,N_9549);
nand U16206 (N_16206,N_9068,N_8360);
xor U16207 (N_16207,N_8496,N_6727);
xor U16208 (N_16208,N_9978,N_7253);
nand U16209 (N_16209,N_7052,N_7179);
or U16210 (N_16210,N_11716,N_11269);
nor U16211 (N_16211,N_10815,N_11321);
and U16212 (N_16212,N_12219,N_11065);
and U16213 (N_16213,N_10801,N_10328);
xor U16214 (N_16214,N_10382,N_10906);
or U16215 (N_16215,N_12279,N_6841);
or U16216 (N_16216,N_10749,N_11040);
nand U16217 (N_16217,N_8829,N_7290);
or U16218 (N_16218,N_12047,N_7276);
xnor U16219 (N_16219,N_7807,N_10362);
nand U16220 (N_16220,N_11743,N_9301);
nand U16221 (N_16221,N_9429,N_12025);
or U16222 (N_16222,N_10086,N_9477);
nor U16223 (N_16223,N_11632,N_10373);
xor U16224 (N_16224,N_8368,N_6543);
xnor U16225 (N_16225,N_10542,N_9844);
nand U16226 (N_16226,N_9267,N_6660);
nor U16227 (N_16227,N_11748,N_7311);
or U16228 (N_16228,N_11437,N_7117);
or U16229 (N_16229,N_9158,N_6934);
or U16230 (N_16230,N_11188,N_9961);
xnor U16231 (N_16231,N_7727,N_11681);
nand U16232 (N_16232,N_10621,N_8695);
nand U16233 (N_16233,N_11566,N_8350);
nor U16234 (N_16234,N_7277,N_8508);
xnor U16235 (N_16235,N_7463,N_10574);
nand U16236 (N_16236,N_8535,N_8311);
xnor U16237 (N_16237,N_8081,N_10101);
nand U16238 (N_16238,N_9832,N_9138);
nor U16239 (N_16239,N_7308,N_7900);
nand U16240 (N_16240,N_10012,N_12123);
nor U16241 (N_16241,N_11927,N_6287);
nand U16242 (N_16242,N_7603,N_10301);
xor U16243 (N_16243,N_10549,N_12049);
xor U16244 (N_16244,N_11444,N_10906);
xnor U16245 (N_16245,N_7508,N_11924);
nor U16246 (N_16246,N_8160,N_12034);
nand U16247 (N_16247,N_12310,N_8098);
or U16248 (N_16248,N_7834,N_7309);
xnor U16249 (N_16249,N_8713,N_11096);
or U16250 (N_16250,N_7773,N_8712);
or U16251 (N_16251,N_11652,N_10949);
or U16252 (N_16252,N_12330,N_6568);
nor U16253 (N_16253,N_8166,N_6795);
xnor U16254 (N_16254,N_6622,N_10294);
nor U16255 (N_16255,N_7272,N_7235);
nand U16256 (N_16256,N_8590,N_11514);
nor U16257 (N_16257,N_11970,N_9884);
nor U16258 (N_16258,N_9682,N_8115);
and U16259 (N_16259,N_6797,N_11602);
nand U16260 (N_16260,N_11190,N_6662);
xnor U16261 (N_16261,N_8158,N_12117);
xor U16262 (N_16262,N_11685,N_6878);
nand U16263 (N_16263,N_8694,N_7724);
or U16264 (N_16264,N_10303,N_9964);
and U16265 (N_16265,N_8111,N_8604);
nand U16266 (N_16266,N_12207,N_10582);
or U16267 (N_16267,N_11034,N_11611);
xor U16268 (N_16268,N_7404,N_6958);
and U16269 (N_16269,N_7457,N_9259);
nand U16270 (N_16270,N_10612,N_7312);
nor U16271 (N_16271,N_9655,N_12028);
nor U16272 (N_16272,N_12377,N_11987);
or U16273 (N_16273,N_6486,N_8556);
and U16274 (N_16274,N_12171,N_10966);
nor U16275 (N_16275,N_10013,N_9346);
or U16276 (N_16276,N_7073,N_12322);
or U16277 (N_16277,N_6473,N_8316);
and U16278 (N_16278,N_8212,N_11185);
or U16279 (N_16279,N_6844,N_9612);
and U16280 (N_16280,N_6787,N_11989);
xnor U16281 (N_16281,N_11407,N_11916);
xnor U16282 (N_16282,N_10657,N_10053);
xnor U16283 (N_16283,N_9111,N_8316);
nor U16284 (N_16284,N_10045,N_9748);
nand U16285 (N_16285,N_8260,N_10776);
xor U16286 (N_16286,N_11399,N_6295);
or U16287 (N_16287,N_8269,N_8665);
nor U16288 (N_16288,N_9985,N_10592);
or U16289 (N_16289,N_8371,N_6537);
xor U16290 (N_16290,N_11061,N_8816);
and U16291 (N_16291,N_8504,N_7777);
and U16292 (N_16292,N_9985,N_10981);
nor U16293 (N_16293,N_10199,N_11433);
nand U16294 (N_16294,N_10622,N_9378);
or U16295 (N_16295,N_10999,N_11102);
or U16296 (N_16296,N_6824,N_10569);
nand U16297 (N_16297,N_11543,N_9083);
and U16298 (N_16298,N_7617,N_9428);
or U16299 (N_16299,N_7683,N_11825);
nor U16300 (N_16300,N_7404,N_10929);
and U16301 (N_16301,N_9495,N_8180);
and U16302 (N_16302,N_11115,N_8530);
and U16303 (N_16303,N_9378,N_8207);
nand U16304 (N_16304,N_12058,N_10482);
nand U16305 (N_16305,N_12133,N_12372);
nor U16306 (N_16306,N_9739,N_7746);
nand U16307 (N_16307,N_11579,N_9844);
or U16308 (N_16308,N_10604,N_11983);
nand U16309 (N_16309,N_9671,N_6898);
or U16310 (N_16310,N_7533,N_10918);
nor U16311 (N_16311,N_9448,N_9112);
and U16312 (N_16312,N_9273,N_10754);
nand U16313 (N_16313,N_11889,N_10296);
or U16314 (N_16314,N_7275,N_7660);
or U16315 (N_16315,N_9365,N_12361);
xor U16316 (N_16316,N_7165,N_11718);
nor U16317 (N_16317,N_7152,N_9731);
and U16318 (N_16318,N_9154,N_6389);
nand U16319 (N_16319,N_8027,N_7178);
nor U16320 (N_16320,N_8994,N_9609);
nor U16321 (N_16321,N_8037,N_11393);
or U16322 (N_16322,N_6945,N_11209);
and U16323 (N_16323,N_11286,N_11631);
and U16324 (N_16324,N_10913,N_6367);
nand U16325 (N_16325,N_6961,N_7919);
and U16326 (N_16326,N_10318,N_8022);
or U16327 (N_16327,N_9739,N_12207);
and U16328 (N_16328,N_7318,N_12045);
or U16329 (N_16329,N_11608,N_8818);
nand U16330 (N_16330,N_11466,N_9123);
nor U16331 (N_16331,N_8691,N_8216);
nand U16332 (N_16332,N_7521,N_6759);
nand U16333 (N_16333,N_7594,N_7434);
xor U16334 (N_16334,N_7779,N_12036);
xnor U16335 (N_16335,N_9504,N_9469);
nand U16336 (N_16336,N_9996,N_9017);
or U16337 (N_16337,N_8095,N_7386);
nor U16338 (N_16338,N_6910,N_11653);
nor U16339 (N_16339,N_9380,N_9029);
nor U16340 (N_16340,N_10507,N_8852);
nor U16341 (N_16341,N_6330,N_6995);
and U16342 (N_16342,N_8810,N_9026);
and U16343 (N_16343,N_7131,N_11168);
and U16344 (N_16344,N_6884,N_11795);
nand U16345 (N_16345,N_7320,N_6268);
nand U16346 (N_16346,N_10892,N_7771);
or U16347 (N_16347,N_12336,N_9435);
or U16348 (N_16348,N_7212,N_8044);
xor U16349 (N_16349,N_9386,N_10206);
or U16350 (N_16350,N_10933,N_9986);
xor U16351 (N_16351,N_8458,N_7225);
nand U16352 (N_16352,N_9909,N_9194);
nor U16353 (N_16353,N_8717,N_11542);
nor U16354 (N_16354,N_8843,N_9584);
and U16355 (N_16355,N_7925,N_7560);
nand U16356 (N_16356,N_7186,N_11987);
or U16357 (N_16357,N_6632,N_9008);
nor U16358 (N_16358,N_7679,N_8108);
or U16359 (N_16359,N_6363,N_8415);
and U16360 (N_16360,N_8572,N_10944);
and U16361 (N_16361,N_12216,N_8459);
and U16362 (N_16362,N_8742,N_9086);
or U16363 (N_16363,N_8246,N_7434);
xor U16364 (N_16364,N_6537,N_6707);
nor U16365 (N_16365,N_7454,N_12032);
and U16366 (N_16366,N_7575,N_12212);
xor U16367 (N_16367,N_8385,N_7921);
and U16368 (N_16368,N_8490,N_11012);
xnor U16369 (N_16369,N_8842,N_6264);
nand U16370 (N_16370,N_11267,N_7044);
or U16371 (N_16371,N_8200,N_8553);
or U16372 (N_16372,N_7297,N_10005);
nor U16373 (N_16373,N_11917,N_11717);
and U16374 (N_16374,N_8009,N_11733);
or U16375 (N_16375,N_8681,N_7632);
nand U16376 (N_16376,N_12212,N_11181);
nand U16377 (N_16377,N_9922,N_8423);
nor U16378 (N_16378,N_7845,N_8810);
xnor U16379 (N_16379,N_10017,N_10966);
nand U16380 (N_16380,N_9370,N_11322);
nor U16381 (N_16381,N_11409,N_6486);
nor U16382 (N_16382,N_7528,N_9957);
and U16383 (N_16383,N_9572,N_10373);
nand U16384 (N_16384,N_10882,N_7917);
xnor U16385 (N_16385,N_10850,N_11111);
or U16386 (N_16386,N_10608,N_12083);
and U16387 (N_16387,N_8698,N_9032);
or U16388 (N_16388,N_8946,N_11122);
nand U16389 (N_16389,N_9337,N_8013);
or U16390 (N_16390,N_7283,N_7156);
and U16391 (N_16391,N_7319,N_6910);
xnor U16392 (N_16392,N_7473,N_8332);
or U16393 (N_16393,N_9352,N_6892);
or U16394 (N_16394,N_7517,N_6918);
or U16395 (N_16395,N_7428,N_9658);
nor U16396 (N_16396,N_11560,N_6396);
xnor U16397 (N_16397,N_9899,N_11872);
nand U16398 (N_16398,N_10608,N_6957);
nand U16399 (N_16399,N_8253,N_10537);
or U16400 (N_16400,N_9865,N_9391);
and U16401 (N_16401,N_11864,N_11178);
nand U16402 (N_16402,N_10217,N_10320);
nand U16403 (N_16403,N_8318,N_8992);
nor U16404 (N_16404,N_11964,N_9960);
and U16405 (N_16405,N_6536,N_11517);
nor U16406 (N_16406,N_9638,N_12491);
nor U16407 (N_16407,N_7472,N_6795);
and U16408 (N_16408,N_8916,N_6897);
nor U16409 (N_16409,N_8524,N_12306);
nand U16410 (N_16410,N_12328,N_9985);
nand U16411 (N_16411,N_9315,N_6602);
and U16412 (N_16412,N_10363,N_7141);
and U16413 (N_16413,N_7660,N_6849);
nor U16414 (N_16414,N_6466,N_9192);
nand U16415 (N_16415,N_6899,N_6801);
and U16416 (N_16416,N_8868,N_10947);
and U16417 (N_16417,N_10297,N_8959);
or U16418 (N_16418,N_10305,N_7559);
xor U16419 (N_16419,N_9181,N_10940);
nor U16420 (N_16420,N_7949,N_8415);
and U16421 (N_16421,N_12062,N_9841);
nor U16422 (N_16422,N_6948,N_7739);
or U16423 (N_16423,N_10785,N_11676);
or U16424 (N_16424,N_11630,N_12233);
or U16425 (N_16425,N_7587,N_10239);
or U16426 (N_16426,N_8788,N_10943);
and U16427 (N_16427,N_11081,N_7379);
nand U16428 (N_16428,N_6825,N_9958);
nor U16429 (N_16429,N_10946,N_10650);
xor U16430 (N_16430,N_10467,N_11154);
or U16431 (N_16431,N_10392,N_9883);
xor U16432 (N_16432,N_8027,N_10036);
nor U16433 (N_16433,N_10244,N_9115);
or U16434 (N_16434,N_10786,N_7565);
and U16435 (N_16435,N_8144,N_7930);
nor U16436 (N_16436,N_7199,N_11356);
or U16437 (N_16437,N_11597,N_11128);
nand U16438 (N_16438,N_10914,N_9507);
and U16439 (N_16439,N_11242,N_9076);
nor U16440 (N_16440,N_7384,N_10379);
nor U16441 (N_16441,N_7343,N_9893);
nand U16442 (N_16442,N_11346,N_6688);
or U16443 (N_16443,N_7172,N_9916);
nand U16444 (N_16444,N_8266,N_12208);
xnor U16445 (N_16445,N_6686,N_12137);
xnor U16446 (N_16446,N_7690,N_7319);
nand U16447 (N_16447,N_9811,N_8186);
or U16448 (N_16448,N_11801,N_11642);
nand U16449 (N_16449,N_9627,N_12441);
nor U16450 (N_16450,N_9919,N_10911);
xnor U16451 (N_16451,N_10820,N_10016);
and U16452 (N_16452,N_8740,N_8061);
xnor U16453 (N_16453,N_9094,N_11023);
nand U16454 (N_16454,N_10262,N_10515);
nor U16455 (N_16455,N_12210,N_10493);
or U16456 (N_16456,N_10004,N_6816);
nor U16457 (N_16457,N_10226,N_10696);
nor U16458 (N_16458,N_6374,N_7373);
and U16459 (N_16459,N_6932,N_10162);
nand U16460 (N_16460,N_11337,N_11300);
and U16461 (N_16461,N_9359,N_8509);
or U16462 (N_16462,N_7811,N_9884);
nor U16463 (N_16463,N_10582,N_7562);
nor U16464 (N_16464,N_11125,N_11284);
xor U16465 (N_16465,N_9594,N_11893);
or U16466 (N_16466,N_12033,N_7545);
nand U16467 (N_16467,N_11488,N_11124);
nand U16468 (N_16468,N_8413,N_12220);
nor U16469 (N_16469,N_10392,N_11649);
nand U16470 (N_16470,N_10162,N_9036);
or U16471 (N_16471,N_9890,N_11933);
nor U16472 (N_16472,N_9258,N_7390);
nand U16473 (N_16473,N_9648,N_10762);
and U16474 (N_16474,N_6359,N_10723);
nand U16475 (N_16475,N_9291,N_7889);
nor U16476 (N_16476,N_9032,N_8996);
xnor U16477 (N_16477,N_8159,N_11783);
and U16478 (N_16478,N_9636,N_11590);
nor U16479 (N_16479,N_8585,N_11773);
nor U16480 (N_16480,N_9508,N_7577);
and U16481 (N_16481,N_8717,N_6626);
xor U16482 (N_16482,N_8358,N_6418);
nand U16483 (N_16483,N_6391,N_9828);
nor U16484 (N_16484,N_6319,N_7422);
nand U16485 (N_16485,N_10232,N_11015);
nand U16486 (N_16486,N_8412,N_6945);
xor U16487 (N_16487,N_11084,N_9103);
nand U16488 (N_16488,N_9799,N_8443);
and U16489 (N_16489,N_6926,N_7356);
nor U16490 (N_16490,N_9399,N_7879);
or U16491 (N_16491,N_9628,N_9133);
or U16492 (N_16492,N_12022,N_12142);
and U16493 (N_16493,N_8861,N_12147);
or U16494 (N_16494,N_7180,N_7276);
nor U16495 (N_16495,N_10861,N_10662);
and U16496 (N_16496,N_11553,N_9005);
and U16497 (N_16497,N_9388,N_6286);
nor U16498 (N_16498,N_9722,N_9885);
nand U16499 (N_16499,N_11452,N_11128);
and U16500 (N_16500,N_7676,N_12399);
xnor U16501 (N_16501,N_8597,N_8468);
nand U16502 (N_16502,N_8550,N_8547);
or U16503 (N_16503,N_12041,N_9006);
nor U16504 (N_16504,N_6412,N_8833);
and U16505 (N_16505,N_6605,N_9262);
and U16506 (N_16506,N_11923,N_9011);
or U16507 (N_16507,N_6541,N_9138);
nor U16508 (N_16508,N_8365,N_11513);
and U16509 (N_16509,N_10702,N_7991);
or U16510 (N_16510,N_6583,N_11194);
nand U16511 (N_16511,N_11835,N_7659);
and U16512 (N_16512,N_10608,N_8419);
or U16513 (N_16513,N_7536,N_7303);
nor U16514 (N_16514,N_10869,N_11301);
nor U16515 (N_16515,N_11536,N_9115);
and U16516 (N_16516,N_8091,N_10820);
nand U16517 (N_16517,N_10991,N_10707);
nand U16518 (N_16518,N_11686,N_9065);
nand U16519 (N_16519,N_6293,N_7934);
or U16520 (N_16520,N_11309,N_10348);
nand U16521 (N_16521,N_6333,N_8243);
or U16522 (N_16522,N_6577,N_7640);
or U16523 (N_16523,N_6676,N_7506);
or U16524 (N_16524,N_10462,N_7521);
nand U16525 (N_16525,N_9859,N_9486);
and U16526 (N_16526,N_7884,N_7450);
xor U16527 (N_16527,N_6656,N_7699);
or U16528 (N_16528,N_7433,N_10133);
and U16529 (N_16529,N_10771,N_10083);
nand U16530 (N_16530,N_6261,N_9157);
and U16531 (N_16531,N_12341,N_9196);
or U16532 (N_16532,N_6682,N_10269);
or U16533 (N_16533,N_12463,N_8057);
nor U16534 (N_16534,N_12121,N_10334);
nor U16535 (N_16535,N_7175,N_11012);
nor U16536 (N_16536,N_6966,N_7753);
nand U16537 (N_16537,N_11661,N_8249);
nor U16538 (N_16538,N_6349,N_7086);
or U16539 (N_16539,N_8382,N_6396);
and U16540 (N_16540,N_12222,N_8912);
nor U16541 (N_16541,N_9953,N_11997);
or U16542 (N_16542,N_11469,N_11648);
nor U16543 (N_16543,N_10373,N_11429);
or U16544 (N_16544,N_7487,N_6568);
nor U16545 (N_16545,N_6628,N_10733);
nand U16546 (N_16546,N_10054,N_9391);
or U16547 (N_16547,N_11922,N_11297);
or U16548 (N_16548,N_6363,N_12499);
or U16549 (N_16549,N_11901,N_11946);
nand U16550 (N_16550,N_9545,N_6298);
nor U16551 (N_16551,N_8015,N_9715);
xor U16552 (N_16552,N_6408,N_11754);
nor U16553 (N_16553,N_7462,N_10698);
and U16554 (N_16554,N_7168,N_9679);
nand U16555 (N_16555,N_11816,N_10353);
nor U16556 (N_16556,N_6378,N_9213);
or U16557 (N_16557,N_7971,N_8757);
nand U16558 (N_16558,N_8887,N_9842);
or U16559 (N_16559,N_7078,N_11062);
or U16560 (N_16560,N_8934,N_10232);
nand U16561 (N_16561,N_7234,N_10655);
nor U16562 (N_16562,N_8053,N_9431);
or U16563 (N_16563,N_12253,N_11871);
or U16564 (N_16564,N_6710,N_9187);
nand U16565 (N_16565,N_11594,N_11041);
nor U16566 (N_16566,N_11123,N_10428);
nand U16567 (N_16567,N_10531,N_7002);
xnor U16568 (N_16568,N_7855,N_8084);
nand U16569 (N_16569,N_9719,N_10588);
nor U16570 (N_16570,N_11695,N_10497);
nand U16571 (N_16571,N_10543,N_12064);
and U16572 (N_16572,N_7230,N_9284);
nor U16573 (N_16573,N_7262,N_11094);
nor U16574 (N_16574,N_7829,N_8930);
xor U16575 (N_16575,N_12482,N_8687);
xnor U16576 (N_16576,N_10026,N_7826);
xnor U16577 (N_16577,N_10592,N_12489);
xnor U16578 (N_16578,N_8324,N_7503);
xor U16579 (N_16579,N_10064,N_11844);
xnor U16580 (N_16580,N_6431,N_9084);
nand U16581 (N_16581,N_11772,N_10211);
xor U16582 (N_16582,N_12364,N_7532);
nor U16583 (N_16583,N_8344,N_6445);
nor U16584 (N_16584,N_6846,N_11992);
or U16585 (N_16585,N_9263,N_11738);
or U16586 (N_16586,N_9985,N_9909);
nand U16587 (N_16587,N_10195,N_12119);
nand U16588 (N_16588,N_12092,N_11130);
and U16589 (N_16589,N_10142,N_9386);
xor U16590 (N_16590,N_12457,N_11637);
nand U16591 (N_16591,N_11943,N_7572);
nor U16592 (N_16592,N_10797,N_8238);
nand U16593 (N_16593,N_8744,N_9556);
xnor U16594 (N_16594,N_9295,N_7973);
or U16595 (N_16595,N_10421,N_10305);
xor U16596 (N_16596,N_8422,N_8310);
xor U16597 (N_16597,N_8821,N_9145);
xor U16598 (N_16598,N_6382,N_10518);
and U16599 (N_16599,N_12199,N_9034);
nor U16600 (N_16600,N_6586,N_11093);
nor U16601 (N_16601,N_6862,N_9907);
nand U16602 (N_16602,N_8648,N_10711);
xnor U16603 (N_16603,N_9792,N_8769);
nor U16604 (N_16604,N_11448,N_7338);
xnor U16605 (N_16605,N_10417,N_10971);
nand U16606 (N_16606,N_8557,N_11370);
nand U16607 (N_16607,N_8612,N_9957);
nand U16608 (N_16608,N_8326,N_10946);
xor U16609 (N_16609,N_8028,N_7931);
and U16610 (N_16610,N_8828,N_10882);
xor U16611 (N_16611,N_11453,N_9278);
and U16612 (N_16612,N_10310,N_11120);
xor U16613 (N_16613,N_10580,N_6407);
nand U16614 (N_16614,N_10170,N_9376);
nand U16615 (N_16615,N_8203,N_7134);
nor U16616 (N_16616,N_6291,N_7451);
and U16617 (N_16617,N_8903,N_8270);
or U16618 (N_16618,N_6644,N_12022);
and U16619 (N_16619,N_8482,N_6844);
nand U16620 (N_16620,N_7499,N_8145);
nand U16621 (N_16621,N_11627,N_9838);
nand U16622 (N_16622,N_9236,N_6290);
and U16623 (N_16623,N_7630,N_8089);
or U16624 (N_16624,N_8467,N_8585);
xor U16625 (N_16625,N_11294,N_8657);
nand U16626 (N_16626,N_11691,N_7436);
xnor U16627 (N_16627,N_6824,N_9326);
nand U16628 (N_16628,N_9303,N_9808);
xnor U16629 (N_16629,N_12425,N_6457);
and U16630 (N_16630,N_10626,N_8581);
or U16631 (N_16631,N_7481,N_7577);
nand U16632 (N_16632,N_11251,N_10733);
or U16633 (N_16633,N_10729,N_12183);
and U16634 (N_16634,N_7087,N_7732);
and U16635 (N_16635,N_9882,N_12367);
xnor U16636 (N_16636,N_6908,N_8048);
nor U16637 (N_16637,N_9837,N_6517);
nand U16638 (N_16638,N_7776,N_12242);
or U16639 (N_16639,N_6990,N_8434);
xnor U16640 (N_16640,N_10395,N_10339);
or U16641 (N_16641,N_8906,N_10102);
nor U16642 (N_16642,N_8749,N_8411);
and U16643 (N_16643,N_8960,N_9611);
and U16644 (N_16644,N_6876,N_11743);
nor U16645 (N_16645,N_10056,N_7423);
or U16646 (N_16646,N_12368,N_7647);
xnor U16647 (N_16647,N_8195,N_7347);
xnor U16648 (N_16648,N_8988,N_8117);
xor U16649 (N_16649,N_6304,N_9806);
nor U16650 (N_16650,N_7569,N_7973);
or U16651 (N_16651,N_9459,N_6484);
xnor U16652 (N_16652,N_7798,N_11732);
nor U16653 (N_16653,N_10877,N_11597);
nor U16654 (N_16654,N_12226,N_12394);
nor U16655 (N_16655,N_11488,N_6675);
and U16656 (N_16656,N_11053,N_10947);
and U16657 (N_16657,N_11478,N_7540);
and U16658 (N_16658,N_8320,N_8562);
and U16659 (N_16659,N_11789,N_7327);
or U16660 (N_16660,N_6794,N_8877);
nand U16661 (N_16661,N_6838,N_10705);
xnor U16662 (N_16662,N_8209,N_10698);
nand U16663 (N_16663,N_6811,N_8302);
xor U16664 (N_16664,N_10913,N_7138);
and U16665 (N_16665,N_12022,N_8913);
and U16666 (N_16666,N_9099,N_10748);
nor U16667 (N_16667,N_12486,N_10044);
xor U16668 (N_16668,N_10773,N_11175);
or U16669 (N_16669,N_10437,N_7382);
xnor U16670 (N_16670,N_10635,N_7207);
nor U16671 (N_16671,N_9250,N_6528);
xnor U16672 (N_16672,N_11256,N_6328);
xor U16673 (N_16673,N_6482,N_11563);
nand U16674 (N_16674,N_7204,N_9679);
nor U16675 (N_16675,N_10119,N_10955);
xor U16676 (N_16676,N_8422,N_6706);
and U16677 (N_16677,N_8101,N_9209);
or U16678 (N_16678,N_6373,N_11509);
or U16679 (N_16679,N_6265,N_6943);
nor U16680 (N_16680,N_12064,N_11546);
xor U16681 (N_16681,N_10955,N_12352);
nand U16682 (N_16682,N_9103,N_11580);
nand U16683 (N_16683,N_11204,N_7304);
xor U16684 (N_16684,N_7662,N_9246);
nor U16685 (N_16685,N_10907,N_9183);
xor U16686 (N_16686,N_7456,N_8354);
and U16687 (N_16687,N_11398,N_7753);
and U16688 (N_16688,N_7570,N_10612);
nand U16689 (N_16689,N_11498,N_6341);
and U16690 (N_16690,N_10055,N_11316);
xor U16691 (N_16691,N_8013,N_9943);
or U16692 (N_16692,N_10822,N_6256);
nor U16693 (N_16693,N_10626,N_6995);
nand U16694 (N_16694,N_10766,N_7082);
nor U16695 (N_16695,N_7926,N_8428);
or U16696 (N_16696,N_12268,N_7616);
or U16697 (N_16697,N_11796,N_6618);
or U16698 (N_16698,N_12145,N_8578);
xnor U16699 (N_16699,N_7600,N_9455);
nand U16700 (N_16700,N_7287,N_7235);
nor U16701 (N_16701,N_11198,N_9407);
and U16702 (N_16702,N_12095,N_10638);
xor U16703 (N_16703,N_11164,N_10250);
and U16704 (N_16704,N_9283,N_9711);
or U16705 (N_16705,N_10887,N_10063);
xnor U16706 (N_16706,N_6765,N_6698);
nand U16707 (N_16707,N_11195,N_7169);
and U16708 (N_16708,N_12160,N_11025);
nand U16709 (N_16709,N_7803,N_9471);
xnor U16710 (N_16710,N_8350,N_6560);
or U16711 (N_16711,N_10375,N_10371);
xor U16712 (N_16712,N_12365,N_10742);
xor U16713 (N_16713,N_8661,N_11477);
xnor U16714 (N_16714,N_8539,N_7916);
nand U16715 (N_16715,N_7922,N_8177);
nor U16716 (N_16716,N_7568,N_6379);
nor U16717 (N_16717,N_8789,N_10489);
xor U16718 (N_16718,N_10028,N_11003);
nand U16719 (N_16719,N_6781,N_7514);
or U16720 (N_16720,N_7802,N_7560);
and U16721 (N_16721,N_11674,N_6749);
nor U16722 (N_16722,N_9831,N_10849);
and U16723 (N_16723,N_7782,N_7993);
xnor U16724 (N_16724,N_12126,N_8032);
or U16725 (N_16725,N_9102,N_11088);
and U16726 (N_16726,N_8019,N_8150);
nand U16727 (N_16727,N_8751,N_7391);
nor U16728 (N_16728,N_6872,N_11997);
and U16729 (N_16729,N_10944,N_8637);
nor U16730 (N_16730,N_8903,N_6993);
nor U16731 (N_16731,N_8894,N_9934);
and U16732 (N_16732,N_8119,N_6811);
or U16733 (N_16733,N_10339,N_9113);
and U16734 (N_16734,N_10273,N_11337);
xnor U16735 (N_16735,N_10031,N_11178);
nand U16736 (N_16736,N_8723,N_10434);
or U16737 (N_16737,N_11560,N_10870);
xor U16738 (N_16738,N_11504,N_11139);
xor U16739 (N_16739,N_11787,N_9068);
or U16740 (N_16740,N_7155,N_12382);
and U16741 (N_16741,N_12170,N_11287);
nor U16742 (N_16742,N_11224,N_7288);
nor U16743 (N_16743,N_10551,N_7595);
or U16744 (N_16744,N_10444,N_8897);
xor U16745 (N_16745,N_12172,N_10360);
or U16746 (N_16746,N_7275,N_10166);
or U16747 (N_16747,N_9695,N_11846);
xnor U16748 (N_16748,N_9628,N_7778);
and U16749 (N_16749,N_8531,N_12098);
nor U16750 (N_16750,N_11021,N_6675);
and U16751 (N_16751,N_10961,N_7092);
nand U16752 (N_16752,N_7411,N_11227);
and U16753 (N_16753,N_10494,N_11673);
and U16754 (N_16754,N_7278,N_9583);
or U16755 (N_16755,N_10835,N_12245);
nand U16756 (N_16756,N_6454,N_11427);
nor U16757 (N_16757,N_6295,N_11525);
xor U16758 (N_16758,N_8239,N_11357);
and U16759 (N_16759,N_10353,N_6881);
and U16760 (N_16760,N_11484,N_7033);
nor U16761 (N_16761,N_9366,N_9149);
and U16762 (N_16762,N_10549,N_6874);
xnor U16763 (N_16763,N_7240,N_10350);
nor U16764 (N_16764,N_9751,N_10424);
nor U16765 (N_16765,N_6803,N_8832);
and U16766 (N_16766,N_9863,N_12211);
xnor U16767 (N_16767,N_10288,N_10789);
or U16768 (N_16768,N_9310,N_8292);
or U16769 (N_16769,N_8010,N_7952);
and U16770 (N_16770,N_7847,N_8064);
nand U16771 (N_16771,N_10709,N_10547);
and U16772 (N_16772,N_12106,N_7407);
nor U16773 (N_16773,N_10493,N_12291);
xor U16774 (N_16774,N_9534,N_7546);
nor U16775 (N_16775,N_7338,N_6875);
or U16776 (N_16776,N_7067,N_8868);
nand U16777 (N_16777,N_12419,N_11168);
nand U16778 (N_16778,N_12311,N_9123);
nand U16779 (N_16779,N_12044,N_6676);
nor U16780 (N_16780,N_9705,N_8456);
nor U16781 (N_16781,N_7509,N_6453);
nand U16782 (N_16782,N_8518,N_11107);
xor U16783 (N_16783,N_6572,N_12105);
or U16784 (N_16784,N_6575,N_11390);
nand U16785 (N_16785,N_9171,N_9784);
or U16786 (N_16786,N_10712,N_8649);
xnor U16787 (N_16787,N_8978,N_7307);
nand U16788 (N_16788,N_9932,N_9043);
and U16789 (N_16789,N_7649,N_10875);
xor U16790 (N_16790,N_8932,N_6929);
or U16791 (N_16791,N_11755,N_7979);
and U16792 (N_16792,N_9325,N_6907);
nor U16793 (N_16793,N_9159,N_10398);
and U16794 (N_16794,N_7581,N_10077);
nor U16795 (N_16795,N_8325,N_9503);
nand U16796 (N_16796,N_6722,N_10993);
or U16797 (N_16797,N_10993,N_9061);
nor U16798 (N_16798,N_8830,N_11882);
xor U16799 (N_16799,N_12235,N_11937);
nor U16800 (N_16800,N_6765,N_9079);
nand U16801 (N_16801,N_10945,N_12150);
nand U16802 (N_16802,N_7767,N_10929);
nor U16803 (N_16803,N_10784,N_10080);
nand U16804 (N_16804,N_7009,N_7594);
or U16805 (N_16805,N_10382,N_7429);
or U16806 (N_16806,N_8579,N_12393);
xor U16807 (N_16807,N_9879,N_6649);
nand U16808 (N_16808,N_8534,N_10455);
and U16809 (N_16809,N_9184,N_6364);
or U16810 (N_16810,N_10952,N_8739);
nor U16811 (N_16811,N_9944,N_7852);
xnor U16812 (N_16812,N_9183,N_9735);
xnor U16813 (N_16813,N_9057,N_11260);
and U16814 (N_16814,N_8016,N_10570);
xnor U16815 (N_16815,N_10920,N_8930);
or U16816 (N_16816,N_12355,N_10126);
or U16817 (N_16817,N_10062,N_9308);
nand U16818 (N_16818,N_8806,N_8368);
or U16819 (N_16819,N_8836,N_11040);
nand U16820 (N_16820,N_9913,N_8454);
xor U16821 (N_16821,N_9337,N_11123);
and U16822 (N_16822,N_7882,N_8100);
nand U16823 (N_16823,N_8406,N_6707);
and U16824 (N_16824,N_9424,N_7807);
and U16825 (N_16825,N_12196,N_7316);
or U16826 (N_16826,N_6519,N_10417);
nor U16827 (N_16827,N_7521,N_8166);
nor U16828 (N_16828,N_9366,N_8896);
or U16829 (N_16829,N_7906,N_8213);
nor U16830 (N_16830,N_9485,N_11511);
or U16831 (N_16831,N_7994,N_6534);
nor U16832 (N_16832,N_8132,N_9618);
xor U16833 (N_16833,N_8993,N_7160);
xnor U16834 (N_16834,N_6649,N_9702);
or U16835 (N_16835,N_10808,N_9461);
xor U16836 (N_16836,N_8634,N_12350);
nor U16837 (N_16837,N_7032,N_7134);
xor U16838 (N_16838,N_7326,N_10701);
nand U16839 (N_16839,N_8400,N_10002);
and U16840 (N_16840,N_12078,N_9924);
nor U16841 (N_16841,N_8892,N_9283);
and U16842 (N_16842,N_6782,N_9063);
xor U16843 (N_16843,N_11268,N_8386);
xor U16844 (N_16844,N_11518,N_10609);
nor U16845 (N_16845,N_10223,N_7647);
or U16846 (N_16846,N_7958,N_8921);
or U16847 (N_16847,N_12146,N_9218);
or U16848 (N_16848,N_9419,N_9933);
nor U16849 (N_16849,N_6874,N_10289);
nand U16850 (N_16850,N_11362,N_9951);
xnor U16851 (N_16851,N_7451,N_9766);
nor U16852 (N_16852,N_10397,N_7311);
nand U16853 (N_16853,N_6703,N_11336);
nor U16854 (N_16854,N_12318,N_7226);
xnor U16855 (N_16855,N_9781,N_6329);
nand U16856 (N_16856,N_9287,N_10048);
nor U16857 (N_16857,N_8760,N_10011);
and U16858 (N_16858,N_8191,N_10091);
nand U16859 (N_16859,N_7351,N_11464);
or U16860 (N_16860,N_11786,N_8776);
xor U16861 (N_16861,N_10359,N_9515);
nor U16862 (N_16862,N_9910,N_6647);
nor U16863 (N_16863,N_6835,N_12064);
and U16864 (N_16864,N_6932,N_11592);
and U16865 (N_16865,N_12348,N_10773);
nand U16866 (N_16866,N_6593,N_7632);
xnor U16867 (N_16867,N_12340,N_8380);
nor U16868 (N_16868,N_6355,N_10413);
nand U16869 (N_16869,N_9560,N_11730);
and U16870 (N_16870,N_8001,N_8183);
and U16871 (N_16871,N_7166,N_7369);
and U16872 (N_16872,N_8046,N_11599);
nand U16873 (N_16873,N_10401,N_12069);
or U16874 (N_16874,N_10352,N_6947);
nor U16875 (N_16875,N_10855,N_6255);
nor U16876 (N_16876,N_8757,N_11807);
nand U16877 (N_16877,N_8761,N_12414);
xor U16878 (N_16878,N_11139,N_7500);
nand U16879 (N_16879,N_7779,N_12331);
and U16880 (N_16880,N_6621,N_10547);
or U16881 (N_16881,N_12264,N_10893);
nand U16882 (N_16882,N_7161,N_8985);
nor U16883 (N_16883,N_7425,N_6447);
xor U16884 (N_16884,N_7361,N_7866);
nor U16885 (N_16885,N_11820,N_8237);
nor U16886 (N_16886,N_11644,N_10657);
or U16887 (N_16887,N_12210,N_12056);
and U16888 (N_16888,N_11748,N_8955);
nor U16889 (N_16889,N_10807,N_11822);
or U16890 (N_16890,N_8774,N_6496);
or U16891 (N_16891,N_12387,N_8582);
nor U16892 (N_16892,N_10390,N_12473);
nand U16893 (N_16893,N_9823,N_11796);
nor U16894 (N_16894,N_10472,N_10339);
nor U16895 (N_16895,N_11066,N_6931);
xnor U16896 (N_16896,N_9051,N_6515);
and U16897 (N_16897,N_10083,N_6726);
and U16898 (N_16898,N_11120,N_10788);
nand U16899 (N_16899,N_8038,N_8241);
or U16900 (N_16900,N_6578,N_10541);
or U16901 (N_16901,N_8765,N_9628);
nand U16902 (N_16902,N_9987,N_10465);
nand U16903 (N_16903,N_11560,N_6809);
nor U16904 (N_16904,N_6856,N_10106);
or U16905 (N_16905,N_6580,N_7088);
or U16906 (N_16906,N_7937,N_10908);
xor U16907 (N_16907,N_12333,N_10221);
xnor U16908 (N_16908,N_9256,N_8998);
nand U16909 (N_16909,N_10656,N_6943);
and U16910 (N_16910,N_8899,N_9071);
or U16911 (N_16911,N_9652,N_9121);
xor U16912 (N_16912,N_9472,N_7714);
and U16913 (N_16913,N_10133,N_10690);
nor U16914 (N_16914,N_9238,N_9186);
nor U16915 (N_16915,N_11408,N_6325);
xnor U16916 (N_16916,N_11008,N_8862);
nand U16917 (N_16917,N_9542,N_9009);
and U16918 (N_16918,N_12045,N_7495);
nand U16919 (N_16919,N_10127,N_6864);
and U16920 (N_16920,N_12387,N_8080);
and U16921 (N_16921,N_11815,N_11373);
nand U16922 (N_16922,N_6828,N_7975);
nand U16923 (N_16923,N_12018,N_7665);
nand U16924 (N_16924,N_7961,N_6422);
nand U16925 (N_16925,N_10215,N_6274);
nor U16926 (N_16926,N_8979,N_7832);
nor U16927 (N_16927,N_7657,N_8316);
nor U16928 (N_16928,N_8114,N_9589);
nand U16929 (N_16929,N_10323,N_8146);
nor U16930 (N_16930,N_11989,N_9640);
nand U16931 (N_16931,N_6402,N_7436);
and U16932 (N_16932,N_10717,N_9286);
and U16933 (N_16933,N_7574,N_7947);
nor U16934 (N_16934,N_12339,N_8892);
nor U16935 (N_16935,N_10108,N_8408);
nand U16936 (N_16936,N_7042,N_10160);
and U16937 (N_16937,N_7368,N_8077);
nor U16938 (N_16938,N_11671,N_10513);
nor U16939 (N_16939,N_10937,N_7741);
and U16940 (N_16940,N_10554,N_6477);
nand U16941 (N_16941,N_8969,N_8734);
nand U16942 (N_16942,N_8992,N_11355);
nor U16943 (N_16943,N_9786,N_12019);
xor U16944 (N_16944,N_7199,N_10331);
nor U16945 (N_16945,N_7371,N_9411);
and U16946 (N_16946,N_9237,N_8553);
or U16947 (N_16947,N_6534,N_9986);
or U16948 (N_16948,N_7724,N_6887);
or U16949 (N_16949,N_6627,N_11536);
nor U16950 (N_16950,N_12201,N_12318);
and U16951 (N_16951,N_7385,N_8367);
xor U16952 (N_16952,N_6413,N_8829);
and U16953 (N_16953,N_8512,N_12435);
and U16954 (N_16954,N_7136,N_7124);
and U16955 (N_16955,N_9457,N_12146);
or U16956 (N_16956,N_9769,N_11948);
xnor U16957 (N_16957,N_6898,N_7289);
or U16958 (N_16958,N_8532,N_10405);
nand U16959 (N_16959,N_10727,N_9833);
nand U16960 (N_16960,N_7764,N_11672);
or U16961 (N_16961,N_10912,N_9839);
and U16962 (N_16962,N_12187,N_9274);
nand U16963 (N_16963,N_11079,N_8986);
nor U16964 (N_16964,N_9365,N_6641);
nand U16965 (N_16965,N_8655,N_6831);
nand U16966 (N_16966,N_12367,N_7165);
or U16967 (N_16967,N_8573,N_7674);
xnor U16968 (N_16968,N_10537,N_10356);
and U16969 (N_16969,N_10245,N_7630);
xor U16970 (N_16970,N_9823,N_7905);
or U16971 (N_16971,N_9312,N_12393);
or U16972 (N_16972,N_11080,N_8293);
or U16973 (N_16973,N_7805,N_6381);
or U16974 (N_16974,N_10868,N_9482);
and U16975 (N_16975,N_10363,N_6534);
and U16976 (N_16976,N_6489,N_6336);
and U16977 (N_16977,N_7948,N_7739);
nor U16978 (N_16978,N_8651,N_8771);
nand U16979 (N_16979,N_8757,N_11265);
or U16980 (N_16980,N_11019,N_9617);
and U16981 (N_16981,N_10679,N_10095);
nor U16982 (N_16982,N_10569,N_9637);
xnor U16983 (N_16983,N_11627,N_6399);
xor U16984 (N_16984,N_10930,N_7787);
and U16985 (N_16985,N_7662,N_12303);
nor U16986 (N_16986,N_8287,N_12279);
xor U16987 (N_16987,N_10303,N_12225);
nor U16988 (N_16988,N_11553,N_6379);
xnor U16989 (N_16989,N_8128,N_9574);
or U16990 (N_16990,N_10519,N_7464);
or U16991 (N_16991,N_12066,N_7883);
nand U16992 (N_16992,N_7684,N_10433);
xnor U16993 (N_16993,N_9086,N_9518);
or U16994 (N_16994,N_9261,N_11898);
xor U16995 (N_16995,N_9974,N_7418);
and U16996 (N_16996,N_9229,N_6737);
or U16997 (N_16997,N_8604,N_8797);
and U16998 (N_16998,N_8817,N_7490);
nand U16999 (N_16999,N_11369,N_11794);
nand U17000 (N_17000,N_12385,N_8337);
nand U17001 (N_17001,N_10112,N_8782);
nor U17002 (N_17002,N_11622,N_9724);
nand U17003 (N_17003,N_7964,N_12464);
or U17004 (N_17004,N_8171,N_9516);
xor U17005 (N_17005,N_11387,N_9262);
nor U17006 (N_17006,N_7898,N_7762);
xor U17007 (N_17007,N_12191,N_11320);
xor U17008 (N_17008,N_8276,N_11966);
nand U17009 (N_17009,N_11488,N_8247);
or U17010 (N_17010,N_9259,N_11511);
and U17011 (N_17011,N_6369,N_11856);
nand U17012 (N_17012,N_7234,N_6264);
or U17013 (N_17013,N_8645,N_8835);
nor U17014 (N_17014,N_10654,N_6339);
nand U17015 (N_17015,N_12066,N_7612);
nand U17016 (N_17016,N_8730,N_9470);
or U17017 (N_17017,N_11774,N_9600);
xor U17018 (N_17018,N_8746,N_10838);
or U17019 (N_17019,N_11805,N_9243);
and U17020 (N_17020,N_11971,N_6328);
nand U17021 (N_17021,N_7809,N_9892);
nor U17022 (N_17022,N_11700,N_7875);
xnor U17023 (N_17023,N_7937,N_10897);
and U17024 (N_17024,N_7514,N_7631);
and U17025 (N_17025,N_8703,N_10951);
nor U17026 (N_17026,N_8239,N_6656);
nor U17027 (N_17027,N_7024,N_12108);
xnor U17028 (N_17028,N_10035,N_11514);
xnor U17029 (N_17029,N_7068,N_8056);
or U17030 (N_17030,N_8629,N_9213);
xnor U17031 (N_17031,N_11788,N_9236);
nor U17032 (N_17032,N_11885,N_7444);
nand U17033 (N_17033,N_7884,N_7645);
nand U17034 (N_17034,N_10606,N_10694);
and U17035 (N_17035,N_12294,N_7342);
nand U17036 (N_17036,N_10484,N_8738);
nand U17037 (N_17037,N_11535,N_8166);
xnor U17038 (N_17038,N_12052,N_6583);
nor U17039 (N_17039,N_10453,N_6980);
and U17040 (N_17040,N_10484,N_10055);
xnor U17041 (N_17041,N_8287,N_12095);
nor U17042 (N_17042,N_12394,N_8649);
nand U17043 (N_17043,N_9651,N_10206);
nor U17044 (N_17044,N_11176,N_9353);
xnor U17045 (N_17045,N_8410,N_10501);
or U17046 (N_17046,N_12133,N_8084);
xnor U17047 (N_17047,N_8652,N_6969);
nor U17048 (N_17048,N_6323,N_10031);
nor U17049 (N_17049,N_7366,N_8191);
xor U17050 (N_17050,N_12499,N_7537);
nor U17051 (N_17051,N_6414,N_9834);
or U17052 (N_17052,N_6941,N_9713);
nor U17053 (N_17053,N_10166,N_9091);
nand U17054 (N_17054,N_7467,N_10168);
xor U17055 (N_17055,N_10794,N_9743);
nor U17056 (N_17056,N_7342,N_10227);
and U17057 (N_17057,N_7045,N_12314);
nor U17058 (N_17058,N_9779,N_6997);
or U17059 (N_17059,N_11405,N_10186);
xnor U17060 (N_17060,N_7976,N_12055);
nor U17061 (N_17061,N_7159,N_9880);
xnor U17062 (N_17062,N_12330,N_6711);
nand U17063 (N_17063,N_6465,N_6346);
xor U17064 (N_17064,N_10137,N_11039);
nand U17065 (N_17065,N_12393,N_8223);
xor U17066 (N_17066,N_12272,N_7056);
and U17067 (N_17067,N_12398,N_10848);
or U17068 (N_17068,N_7191,N_8976);
xor U17069 (N_17069,N_10378,N_6871);
nor U17070 (N_17070,N_8992,N_9579);
nor U17071 (N_17071,N_11072,N_7290);
and U17072 (N_17072,N_7076,N_12332);
nor U17073 (N_17073,N_11955,N_10536);
or U17074 (N_17074,N_6726,N_7838);
or U17075 (N_17075,N_11898,N_6410);
and U17076 (N_17076,N_9917,N_7660);
and U17077 (N_17077,N_12278,N_7232);
nor U17078 (N_17078,N_10289,N_6798);
nor U17079 (N_17079,N_8883,N_7176);
nor U17080 (N_17080,N_6758,N_11821);
or U17081 (N_17081,N_8326,N_10108);
and U17082 (N_17082,N_6346,N_10015);
nand U17083 (N_17083,N_7274,N_7295);
or U17084 (N_17084,N_10277,N_8790);
xnor U17085 (N_17085,N_10645,N_10179);
and U17086 (N_17086,N_7883,N_8987);
or U17087 (N_17087,N_9347,N_11449);
nand U17088 (N_17088,N_6706,N_12091);
nand U17089 (N_17089,N_7327,N_6776);
nor U17090 (N_17090,N_7623,N_8699);
or U17091 (N_17091,N_8930,N_10862);
nor U17092 (N_17092,N_12229,N_8964);
nand U17093 (N_17093,N_10448,N_11957);
nand U17094 (N_17094,N_6255,N_9342);
xnor U17095 (N_17095,N_11599,N_9818);
and U17096 (N_17096,N_8513,N_12319);
or U17097 (N_17097,N_9329,N_10478);
or U17098 (N_17098,N_8430,N_9774);
and U17099 (N_17099,N_6394,N_7897);
and U17100 (N_17100,N_11020,N_11688);
nand U17101 (N_17101,N_10966,N_8152);
nor U17102 (N_17102,N_6826,N_7709);
and U17103 (N_17103,N_11129,N_11183);
nor U17104 (N_17104,N_6904,N_10763);
nand U17105 (N_17105,N_10578,N_11623);
and U17106 (N_17106,N_10852,N_11552);
nand U17107 (N_17107,N_9631,N_9906);
or U17108 (N_17108,N_8748,N_9681);
nor U17109 (N_17109,N_8063,N_8622);
nand U17110 (N_17110,N_7480,N_7148);
and U17111 (N_17111,N_7409,N_12400);
and U17112 (N_17112,N_9831,N_8844);
xor U17113 (N_17113,N_7784,N_8219);
nor U17114 (N_17114,N_6692,N_11948);
or U17115 (N_17115,N_6435,N_8438);
nand U17116 (N_17116,N_7815,N_11549);
nor U17117 (N_17117,N_8601,N_8504);
nor U17118 (N_17118,N_7721,N_12187);
and U17119 (N_17119,N_7745,N_9845);
xnor U17120 (N_17120,N_12209,N_8063);
and U17121 (N_17121,N_9311,N_10160);
xor U17122 (N_17122,N_9546,N_7409);
nor U17123 (N_17123,N_12255,N_10093);
nand U17124 (N_17124,N_9125,N_12091);
nand U17125 (N_17125,N_10322,N_12438);
or U17126 (N_17126,N_10174,N_7380);
and U17127 (N_17127,N_8116,N_9379);
and U17128 (N_17128,N_12457,N_8998);
nand U17129 (N_17129,N_9812,N_6606);
and U17130 (N_17130,N_10321,N_9816);
xor U17131 (N_17131,N_11977,N_6817);
xor U17132 (N_17132,N_8924,N_7185);
xnor U17133 (N_17133,N_9769,N_7090);
nand U17134 (N_17134,N_10313,N_8840);
or U17135 (N_17135,N_6476,N_7826);
nand U17136 (N_17136,N_6849,N_7392);
nor U17137 (N_17137,N_6428,N_7984);
and U17138 (N_17138,N_9847,N_8619);
nand U17139 (N_17139,N_9858,N_11178);
xor U17140 (N_17140,N_10415,N_10681);
xnor U17141 (N_17141,N_10835,N_8191);
xor U17142 (N_17142,N_9253,N_11559);
nor U17143 (N_17143,N_10953,N_11434);
nor U17144 (N_17144,N_6414,N_6443);
nor U17145 (N_17145,N_6922,N_10886);
nand U17146 (N_17146,N_11746,N_10684);
nor U17147 (N_17147,N_9253,N_10475);
xnor U17148 (N_17148,N_7427,N_8262);
nor U17149 (N_17149,N_10942,N_8981);
and U17150 (N_17150,N_10058,N_6957);
nand U17151 (N_17151,N_9948,N_10890);
xnor U17152 (N_17152,N_10200,N_11499);
or U17153 (N_17153,N_9904,N_8581);
or U17154 (N_17154,N_11602,N_10755);
xnor U17155 (N_17155,N_10761,N_12079);
xor U17156 (N_17156,N_9256,N_11086);
xnor U17157 (N_17157,N_6407,N_7501);
and U17158 (N_17158,N_7506,N_10363);
xor U17159 (N_17159,N_11706,N_9622);
xor U17160 (N_17160,N_10873,N_6373);
nand U17161 (N_17161,N_12007,N_10023);
nand U17162 (N_17162,N_11231,N_8729);
nand U17163 (N_17163,N_9423,N_9280);
nor U17164 (N_17164,N_7722,N_8921);
nor U17165 (N_17165,N_8197,N_8551);
nor U17166 (N_17166,N_12180,N_10950);
and U17167 (N_17167,N_10693,N_10436);
xnor U17168 (N_17168,N_7862,N_9550);
and U17169 (N_17169,N_10566,N_7046);
and U17170 (N_17170,N_7708,N_11162);
nand U17171 (N_17171,N_7461,N_11546);
xor U17172 (N_17172,N_12311,N_7773);
nand U17173 (N_17173,N_7300,N_9074);
nand U17174 (N_17174,N_7331,N_11183);
or U17175 (N_17175,N_12271,N_8830);
nor U17176 (N_17176,N_7330,N_6258);
and U17177 (N_17177,N_6631,N_10366);
nor U17178 (N_17178,N_7518,N_10947);
and U17179 (N_17179,N_11879,N_8161);
xor U17180 (N_17180,N_9112,N_8640);
nor U17181 (N_17181,N_8036,N_6577);
and U17182 (N_17182,N_9257,N_7236);
and U17183 (N_17183,N_10061,N_10446);
and U17184 (N_17184,N_6908,N_11602);
and U17185 (N_17185,N_6440,N_12474);
xnor U17186 (N_17186,N_9093,N_6354);
nand U17187 (N_17187,N_8367,N_9263);
xor U17188 (N_17188,N_7847,N_8818);
and U17189 (N_17189,N_6624,N_6977);
or U17190 (N_17190,N_7384,N_7107);
nor U17191 (N_17191,N_9896,N_7752);
xor U17192 (N_17192,N_11202,N_10117);
nor U17193 (N_17193,N_6909,N_11404);
and U17194 (N_17194,N_8928,N_11384);
nor U17195 (N_17195,N_8826,N_6331);
nand U17196 (N_17196,N_11779,N_12148);
nor U17197 (N_17197,N_9686,N_8038);
or U17198 (N_17198,N_7935,N_8869);
xor U17199 (N_17199,N_10029,N_6998);
nand U17200 (N_17200,N_8868,N_12470);
xor U17201 (N_17201,N_8664,N_8621);
or U17202 (N_17202,N_11264,N_6523);
and U17203 (N_17203,N_9049,N_10941);
xor U17204 (N_17204,N_11587,N_11827);
xor U17205 (N_17205,N_11617,N_11848);
nand U17206 (N_17206,N_10225,N_6984);
or U17207 (N_17207,N_10029,N_6250);
nor U17208 (N_17208,N_11739,N_10836);
and U17209 (N_17209,N_7983,N_10208);
and U17210 (N_17210,N_7567,N_7336);
nand U17211 (N_17211,N_9699,N_9526);
nand U17212 (N_17212,N_11845,N_6504);
nand U17213 (N_17213,N_6579,N_9889);
nor U17214 (N_17214,N_9194,N_12259);
nand U17215 (N_17215,N_10646,N_12172);
and U17216 (N_17216,N_7543,N_9874);
and U17217 (N_17217,N_10746,N_9354);
and U17218 (N_17218,N_6313,N_12035);
or U17219 (N_17219,N_9551,N_11814);
nand U17220 (N_17220,N_12048,N_11338);
xnor U17221 (N_17221,N_12220,N_6739);
nand U17222 (N_17222,N_11952,N_10982);
and U17223 (N_17223,N_7036,N_9903);
xnor U17224 (N_17224,N_10129,N_9336);
or U17225 (N_17225,N_7626,N_8067);
xor U17226 (N_17226,N_11552,N_6433);
or U17227 (N_17227,N_7559,N_7148);
or U17228 (N_17228,N_9718,N_7836);
and U17229 (N_17229,N_7701,N_10686);
nand U17230 (N_17230,N_8288,N_9451);
nand U17231 (N_17231,N_7144,N_6830);
xor U17232 (N_17232,N_9542,N_11747);
nor U17233 (N_17233,N_10802,N_7763);
nand U17234 (N_17234,N_6655,N_6364);
nand U17235 (N_17235,N_9957,N_10766);
or U17236 (N_17236,N_8194,N_9451);
or U17237 (N_17237,N_10699,N_8775);
and U17238 (N_17238,N_11906,N_8133);
nand U17239 (N_17239,N_8858,N_6729);
or U17240 (N_17240,N_7665,N_7977);
or U17241 (N_17241,N_7737,N_8552);
nor U17242 (N_17242,N_6611,N_8988);
and U17243 (N_17243,N_11333,N_8850);
xnor U17244 (N_17244,N_11819,N_11551);
nand U17245 (N_17245,N_10061,N_6309);
nor U17246 (N_17246,N_7859,N_11474);
and U17247 (N_17247,N_10539,N_6278);
nor U17248 (N_17248,N_10395,N_11338);
and U17249 (N_17249,N_9314,N_10320);
and U17250 (N_17250,N_10922,N_7738);
nand U17251 (N_17251,N_12272,N_10977);
xnor U17252 (N_17252,N_8938,N_11398);
nand U17253 (N_17253,N_12272,N_6941);
or U17254 (N_17254,N_7520,N_10488);
and U17255 (N_17255,N_6469,N_9388);
or U17256 (N_17256,N_9372,N_7205);
xor U17257 (N_17257,N_6414,N_11186);
nand U17258 (N_17258,N_7587,N_9008);
xnor U17259 (N_17259,N_7873,N_7814);
and U17260 (N_17260,N_6442,N_7217);
nor U17261 (N_17261,N_7052,N_7434);
nor U17262 (N_17262,N_10113,N_12346);
and U17263 (N_17263,N_6706,N_7601);
or U17264 (N_17264,N_11428,N_7539);
and U17265 (N_17265,N_8134,N_11251);
xor U17266 (N_17266,N_12139,N_10069);
nor U17267 (N_17267,N_8158,N_11807);
xor U17268 (N_17268,N_12156,N_10658);
or U17269 (N_17269,N_9593,N_7552);
nor U17270 (N_17270,N_7720,N_8277);
xnor U17271 (N_17271,N_8666,N_11011);
nor U17272 (N_17272,N_12079,N_12393);
nor U17273 (N_17273,N_7201,N_6684);
nand U17274 (N_17274,N_7011,N_8795);
nor U17275 (N_17275,N_7367,N_7166);
and U17276 (N_17276,N_7857,N_6978);
xnor U17277 (N_17277,N_10982,N_9742);
or U17278 (N_17278,N_7990,N_6328);
or U17279 (N_17279,N_10518,N_11482);
or U17280 (N_17280,N_10588,N_9339);
or U17281 (N_17281,N_6962,N_11835);
or U17282 (N_17282,N_10618,N_12443);
nand U17283 (N_17283,N_7996,N_12185);
or U17284 (N_17284,N_10380,N_10627);
nor U17285 (N_17285,N_8267,N_7690);
nand U17286 (N_17286,N_11779,N_9784);
nand U17287 (N_17287,N_9840,N_7451);
and U17288 (N_17288,N_8991,N_8380);
and U17289 (N_17289,N_6688,N_7851);
nand U17290 (N_17290,N_10039,N_12470);
or U17291 (N_17291,N_8222,N_12025);
nor U17292 (N_17292,N_10251,N_6421);
and U17293 (N_17293,N_10398,N_8584);
or U17294 (N_17294,N_9485,N_11686);
nor U17295 (N_17295,N_12491,N_7912);
and U17296 (N_17296,N_9728,N_6299);
nor U17297 (N_17297,N_8015,N_9772);
and U17298 (N_17298,N_9934,N_7181);
xor U17299 (N_17299,N_6269,N_9569);
xor U17300 (N_17300,N_12171,N_11399);
or U17301 (N_17301,N_7629,N_10120);
nor U17302 (N_17302,N_9333,N_6571);
xnor U17303 (N_17303,N_7136,N_10858);
nand U17304 (N_17304,N_7780,N_8458);
nor U17305 (N_17305,N_12461,N_8595);
xor U17306 (N_17306,N_8308,N_7306);
xor U17307 (N_17307,N_8423,N_8063);
or U17308 (N_17308,N_11545,N_6860);
nand U17309 (N_17309,N_11147,N_8138);
and U17310 (N_17310,N_10233,N_9782);
or U17311 (N_17311,N_6372,N_10855);
or U17312 (N_17312,N_9751,N_9612);
and U17313 (N_17313,N_10072,N_7458);
nor U17314 (N_17314,N_10625,N_6711);
nand U17315 (N_17315,N_11914,N_8680);
and U17316 (N_17316,N_12377,N_8656);
nand U17317 (N_17317,N_6340,N_12452);
and U17318 (N_17318,N_11911,N_10001);
xnor U17319 (N_17319,N_11227,N_8011);
xnor U17320 (N_17320,N_11766,N_10095);
and U17321 (N_17321,N_8809,N_9602);
or U17322 (N_17322,N_12463,N_9212);
or U17323 (N_17323,N_9256,N_11734);
or U17324 (N_17324,N_12055,N_7995);
and U17325 (N_17325,N_8153,N_7558);
or U17326 (N_17326,N_10565,N_7787);
nor U17327 (N_17327,N_8481,N_10561);
or U17328 (N_17328,N_9833,N_12355);
nor U17329 (N_17329,N_8659,N_9841);
or U17330 (N_17330,N_8436,N_9998);
or U17331 (N_17331,N_8424,N_10938);
xnor U17332 (N_17332,N_6303,N_7405);
nand U17333 (N_17333,N_10303,N_12447);
nand U17334 (N_17334,N_11798,N_6551);
and U17335 (N_17335,N_7690,N_11330);
nand U17336 (N_17336,N_9758,N_11048);
or U17337 (N_17337,N_12107,N_8796);
nor U17338 (N_17338,N_9586,N_11103);
nor U17339 (N_17339,N_11313,N_7947);
nand U17340 (N_17340,N_7244,N_6658);
and U17341 (N_17341,N_11588,N_10907);
xor U17342 (N_17342,N_8322,N_11645);
or U17343 (N_17343,N_7211,N_8380);
or U17344 (N_17344,N_7331,N_6651);
nor U17345 (N_17345,N_11258,N_9872);
nand U17346 (N_17346,N_9964,N_8361);
and U17347 (N_17347,N_11732,N_7381);
or U17348 (N_17348,N_11031,N_9396);
or U17349 (N_17349,N_6784,N_11946);
xnor U17350 (N_17350,N_6899,N_11724);
nand U17351 (N_17351,N_12369,N_8812);
and U17352 (N_17352,N_10218,N_7224);
nand U17353 (N_17353,N_11738,N_7436);
nor U17354 (N_17354,N_8378,N_6442);
nand U17355 (N_17355,N_10360,N_7821);
xor U17356 (N_17356,N_7070,N_11209);
nand U17357 (N_17357,N_8797,N_9005);
nand U17358 (N_17358,N_11763,N_11028);
xnor U17359 (N_17359,N_10378,N_10604);
and U17360 (N_17360,N_10230,N_10437);
nor U17361 (N_17361,N_9682,N_9713);
or U17362 (N_17362,N_6796,N_9077);
nand U17363 (N_17363,N_8675,N_10381);
or U17364 (N_17364,N_6296,N_10149);
nor U17365 (N_17365,N_6419,N_8747);
nand U17366 (N_17366,N_7049,N_7564);
and U17367 (N_17367,N_6948,N_7559);
xor U17368 (N_17368,N_8007,N_10856);
and U17369 (N_17369,N_7179,N_10028);
nor U17370 (N_17370,N_11694,N_9637);
xor U17371 (N_17371,N_11732,N_10977);
xnor U17372 (N_17372,N_8604,N_11321);
nand U17373 (N_17373,N_8405,N_12381);
nand U17374 (N_17374,N_8299,N_10003);
nor U17375 (N_17375,N_10494,N_7478);
nand U17376 (N_17376,N_6361,N_9788);
nor U17377 (N_17377,N_6520,N_10140);
xnor U17378 (N_17378,N_8030,N_7498);
nor U17379 (N_17379,N_11504,N_10918);
xor U17380 (N_17380,N_7479,N_6415);
nand U17381 (N_17381,N_7392,N_12221);
nor U17382 (N_17382,N_7001,N_6947);
nor U17383 (N_17383,N_10727,N_9574);
nor U17384 (N_17384,N_9441,N_10875);
nor U17385 (N_17385,N_9956,N_7891);
and U17386 (N_17386,N_6628,N_12056);
xnor U17387 (N_17387,N_8184,N_11652);
or U17388 (N_17388,N_10656,N_9602);
nand U17389 (N_17389,N_10692,N_9555);
nor U17390 (N_17390,N_7796,N_6269);
and U17391 (N_17391,N_6745,N_8774);
and U17392 (N_17392,N_9540,N_7868);
and U17393 (N_17393,N_6592,N_9253);
xor U17394 (N_17394,N_9435,N_8701);
and U17395 (N_17395,N_6786,N_8232);
xor U17396 (N_17396,N_11819,N_7664);
and U17397 (N_17397,N_11955,N_8616);
nor U17398 (N_17398,N_12184,N_8269);
nor U17399 (N_17399,N_12219,N_9687);
nand U17400 (N_17400,N_11384,N_6378);
nand U17401 (N_17401,N_8866,N_7857);
nand U17402 (N_17402,N_10197,N_6293);
and U17403 (N_17403,N_11734,N_12224);
nand U17404 (N_17404,N_12496,N_9855);
nor U17405 (N_17405,N_11787,N_7151);
and U17406 (N_17406,N_7445,N_6643);
nor U17407 (N_17407,N_6400,N_10627);
nand U17408 (N_17408,N_11287,N_11838);
or U17409 (N_17409,N_9215,N_6781);
or U17410 (N_17410,N_8655,N_7498);
nor U17411 (N_17411,N_7507,N_8985);
nand U17412 (N_17412,N_11517,N_7657);
nand U17413 (N_17413,N_9366,N_8840);
nand U17414 (N_17414,N_8076,N_8487);
or U17415 (N_17415,N_10150,N_8842);
xnor U17416 (N_17416,N_11923,N_8144);
xnor U17417 (N_17417,N_10246,N_8820);
or U17418 (N_17418,N_9703,N_8354);
or U17419 (N_17419,N_10367,N_7361);
and U17420 (N_17420,N_8229,N_8447);
nand U17421 (N_17421,N_11193,N_9073);
and U17422 (N_17422,N_6546,N_7484);
and U17423 (N_17423,N_11425,N_6312);
or U17424 (N_17424,N_7664,N_7696);
and U17425 (N_17425,N_7269,N_10055);
and U17426 (N_17426,N_6398,N_7231);
xor U17427 (N_17427,N_7550,N_12454);
nor U17428 (N_17428,N_12205,N_6796);
xnor U17429 (N_17429,N_9544,N_11387);
or U17430 (N_17430,N_10227,N_12483);
nand U17431 (N_17431,N_8151,N_8570);
nor U17432 (N_17432,N_9106,N_9091);
nor U17433 (N_17433,N_11251,N_10741);
nand U17434 (N_17434,N_6332,N_9994);
xnor U17435 (N_17435,N_10383,N_10167);
xor U17436 (N_17436,N_9344,N_6730);
nand U17437 (N_17437,N_7512,N_9988);
nor U17438 (N_17438,N_8404,N_9353);
xor U17439 (N_17439,N_11407,N_6912);
or U17440 (N_17440,N_12016,N_8530);
or U17441 (N_17441,N_6753,N_6295);
nor U17442 (N_17442,N_6596,N_7846);
xor U17443 (N_17443,N_10196,N_10964);
or U17444 (N_17444,N_12334,N_7884);
and U17445 (N_17445,N_9741,N_8311);
or U17446 (N_17446,N_8776,N_7157);
nand U17447 (N_17447,N_9273,N_8292);
or U17448 (N_17448,N_11873,N_9693);
xor U17449 (N_17449,N_8511,N_11708);
nor U17450 (N_17450,N_8799,N_8707);
nand U17451 (N_17451,N_9598,N_12216);
and U17452 (N_17452,N_9063,N_8034);
or U17453 (N_17453,N_11070,N_8733);
xnor U17454 (N_17454,N_8248,N_10204);
or U17455 (N_17455,N_7285,N_7710);
or U17456 (N_17456,N_7709,N_9430);
or U17457 (N_17457,N_10434,N_9818);
nand U17458 (N_17458,N_11609,N_11630);
xnor U17459 (N_17459,N_11685,N_6769);
nand U17460 (N_17460,N_10707,N_8747);
nand U17461 (N_17461,N_11544,N_8856);
or U17462 (N_17462,N_8369,N_9495);
and U17463 (N_17463,N_8173,N_11351);
nor U17464 (N_17464,N_8309,N_9976);
or U17465 (N_17465,N_10833,N_8248);
or U17466 (N_17466,N_8924,N_7270);
nor U17467 (N_17467,N_11012,N_10179);
xor U17468 (N_17468,N_11166,N_9119);
and U17469 (N_17469,N_8842,N_11980);
and U17470 (N_17470,N_7150,N_9606);
and U17471 (N_17471,N_8650,N_9891);
nor U17472 (N_17472,N_8558,N_11016);
nor U17473 (N_17473,N_7611,N_9391);
or U17474 (N_17474,N_10491,N_11577);
xnor U17475 (N_17475,N_10040,N_8983);
nand U17476 (N_17476,N_7477,N_8878);
xnor U17477 (N_17477,N_10823,N_6716);
xnor U17478 (N_17478,N_12044,N_9965);
nor U17479 (N_17479,N_8434,N_12079);
and U17480 (N_17480,N_7029,N_9178);
or U17481 (N_17481,N_9743,N_8809);
and U17482 (N_17482,N_10407,N_9996);
nor U17483 (N_17483,N_6900,N_8479);
and U17484 (N_17484,N_6738,N_7246);
and U17485 (N_17485,N_6507,N_9493);
xor U17486 (N_17486,N_6843,N_6978);
nor U17487 (N_17487,N_11990,N_9321);
nand U17488 (N_17488,N_6430,N_7599);
nor U17489 (N_17489,N_11497,N_7242);
xnor U17490 (N_17490,N_11508,N_6330);
or U17491 (N_17491,N_7892,N_11551);
nand U17492 (N_17492,N_9517,N_11682);
or U17493 (N_17493,N_11320,N_11335);
nand U17494 (N_17494,N_7624,N_8473);
or U17495 (N_17495,N_6936,N_8876);
nand U17496 (N_17496,N_8246,N_7345);
nor U17497 (N_17497,N_7704,N_8744);
xnor U17498 (N_17498,N_9134,N_9241);
and U17499 (N_17499,N_6599,N_9153);
or U17500 (N_17500,N_6645,N_6978);
nor U17501 (N_17501,N_7476,N_10520);
nor U17502 (N_17502,N_11061,N_8613);
nand U17503 (N_17503,N_11933,N_9751);
nor U17504 (N_17504,N_11956,N_11051);
and U17505 (N_17505,N_7065,N_12318);
or U17506 (N_17506,N_6338,N_10911);
xnor U17507 (N_17507,N_9997,N_7884);
nand U17508 (N_17508,N_8426,N_11667);
or U17509 (N_17509,N_8075,N_6987);
xor U17510 (N_17510,N_7446,N_11797);
nand U17511 (N_17511,N_11808,N_9857);
nor U17512 (N_17512,N_7984,N_6283);
xnor U17513 (N_17513,N_9072,N_10685);
and U17514 (N_17514,N_10467,N_6471);
or U17515 (N_17515,N_8060,N_11301);
and U17516 (N_17516,N_10044,N_8034);
nor U17517 (N_17517,N_10140,N_7582);
xor U17518 (N_17518,N_9435,N_8794);
nand U17519 (N_17519,N_7086,N_12140);
or U17520 (N_17520,N_10097,N_6376);
nand U17521 (N_17521,N_6642,N_6286);
nor U17522 (N_17522,N_8739,N_8907);
or U17523 (N_17523,N_11893,N_11203);
and U17524 (N_17524,N_8488,N_12244);
nor U17525 (N_17525,N_6714,N_7429);
or U17526 (N_17526,N_8762,N_8604);
or U17527 (N_17527,N_7814,N_8068);
xor U17528 (N_17528,N_11639,N_8531);
xor U17529 (N_17529,N_9352,N_10605);
nand U17530 (N_17530,N_7988,N_7370);
nor U17531 (N_17531,N_9454,N_10707);
and U17532 (N_17532,N_11613,N_8929);
nand U17533 (N_17533,N_10437,N_7002);
nand U17534 (N_17534,N_8872,N_11664);
or U17535 (N_17535,N_8160,N_6399);
and U17536 (N_17536,N_9191,N_11641);
xnor U17537 (N_17537,N_8222,N_8086);
nor U17538 (N_17538,N_8299,N_8516);
nand U17539 (N_17539,N_9700,N_8026);
nand U17540 (N_17540,N_7993,N_7202);
and U17541 (N_17541,N_9621,N_8062);
nor U17542 (N_17542,N_7656,N_11460);
xnor U17543 (N_17543,N_12021,N_10634);
nor U17544 (N_17544,N_7454,N_7339);
or U17545 (N_17545,N_12484,N_10066);
nor U17546 (N_17546,N_8670,N_9812);
nand U17547 (N_17547,N_6914,N_7214);
or U17548 (N_17548,N_9865,N_10932);
or U17549 (N_17549,N_7302,N_10306);
and U17550 (N_17550,N_8861,N_7762);
nor U17551 (N_17551,N_7305,N_10106);
or U17552 (N_17552,N_8728,N_10827);
and U17553 (N_17553,N_11959,N_6998);
and U17554 (N_17554,N_7916,N_11640);
and U17555 (N_17555,N_6301,N_12224);
and U17556 (N_17556,N_7193,N_8526);
or U17557 (N_17557,N_11348,N_10699);
and U17558 (N_17558,N_11281,N_8458);
and U17559 (N_17559,N_7170,N_11312);
or U17560 (N_17560,N_10154,N_10237);
nor U17561 (N_17561,N_10980,N_10672);
nand U17562 (N_17562,N_10596,N_6551);
and U17563 (N_17563,N_10221,N_9664);
and U17564 (N_17564,N_10418,N_12007);
xnor U17565 (N_17565,N_9988,N_7784);
xnor U17566 (N_17566,N_8117,N_10363);
nor U17567 (N_17567,N_11842,N_8369);
nor U17568 (N_17568,N_8010,N_9936);
or U17569 (N_17569,N_8793,N_11547);
or U17570 (N_17570,N_6786,N_7607);
nor U17571 (N_17571,N_9501,N_8714);
or U17572 (N_17572,N_11576,N_7224);
xnor U17573 (N_17573,N_6819,N_11151);
xnor U17574 (N_17574,N_10673,N_6376);
or U17575 (N_17575,N_10040,N_9213);
or U17576 (N_17576,N_11658,N_9192);
nand U17577 (N_17577,N_6301,N_6512);
nor U17578 (N_17578,N_9330,N_9399);
or U17579 (N_17579,N_11746,N_12216);
and U17580 (N_17580,N_9490,N_7093);
or U17581 (N_17581,N_8965,N_10721);
xor U17582 (N_17582,N_10248,N_10062);
or U17583 (N_17583,N_8609,N_11915);
xor U17584 (N_17584,N_7994,N_7778);
nand U17585 (N_17585,N_12225,N_10573);
xnor U17586 (N_17586,N_11900,N_11182);
nand U17587 (N_17587,N_12304,N_10956);
nand U17588 (N_17588,N_8431,N_6839);
or U17589 (N_17589,N_6606,N_11886);
and U17590 (N_17590,N_9589,N_7598);
xnor U17591 (N_17591,N_10508,N_10850);
nor U17592 (N_17592,N_12203,N_11946);
or U17593 (N_17593,N_10153,N_10971);
or U17594 (N_17594,N_9713,N_10897);
or U17595 (N_17595,N_7318,N_7377);
or U17596 (N_17596,N_11197,N_9432);
nand U17597 (N_17597,N_9225,N_8405);
xor U17598 (N_17598,N_8340,N_11025);
or U17599 (N_17599,N_7932,N_9757);
nor U17600 (N_17600,N_7565,N_10315);
or U17601 (N_17601,N_9531,N_12335);
nor U17602 (N_17602,N_7881,N_7141);
nor U17603 (N_17603,N_8462,N_12264);
and U17604 (N_17604,N_9048,N_11704);
and U17605 (N_17605,N_10223,N_12126);
xnor U17606 (N_17606,N_8635,N_9629);
nor U17607 (N_17607,N_9307,N_9044);
nand U17608 (N_17608,N_7855,N_7056);
or U17609 (N_17609,N_8466,N_11343);
xor U17610 (N_17610,N_8808,N_7847);
xor U17611 (N_17611,N_9756,N_8820);
or U17612 (N_17612,N_12169,N_12121);
and U17613 (N_17613,N_11670,N_9358);
xor U17614 (N_17614,N_11614,N_8643);
and U17615 (N_17615,N_7943,N_9088);
or U17616 (N_17616,N_7851,N_8627);
nand U17617 (N_17617,N_9372,N_6517);
xor U17618 (N_17618,N_9323,N_7895);
nor U17619 (N_17619,N_9191,N_11937);
or U17620 (N_17620,N_11350,N_11216);
and U17621 (N_17621,N_9758,N_6396);
nand U17622 (N_17622,N_10867,N_6988);
or U17623 (N_17623,N_6789,N_9239);
or U17624 (N_17624,N_11401,N_7498);
nor U17625 (N_17625,N_7016,N_9647);
nand U17626 (N_17626,N_6315,N_8518);
or U17627 (N_17627,N_7462,N_9569);
nand U17628 (N_17628,N_11342,N_12369);
and U17629 (N_17629,N_6738,N_10832);
nor U17630 (N_17630,N_7422,N_11699);
xor U17631 (N_17631,N_9321,N_9888);
nor U17632 (N_17632,N_9212,N_6649);
or U17633 (N_17633,N_10626,N_10361);
and U17634 (N_17634,N_12333,N_7580);
or U17635 (N_17635,N_12474,N_10778);
and U17636 (N_17636,N_9030,N_8761);
xor U17637 (N_17637,N_9472,N_9205);
and U17638 (N_17638,N_10957,N_11986);
or U17639 (N_17639,N_9473,N_8569);
nand U17640 (N_17640,N_6643,N_10426);
nor U17641 (N_17641,N_7539,N_11197);
or U17642 (N_17642,N_8834,N_12110);
or U17643 (N_17643,N_8047,N_12051);
nor U17644 (N_17644,N_8633,N_9911);
and U17645 (N_17645,N_11715,N_10149);
nor U17646 (N_17646,N_9921,N_7599);
nand U17647 (N_17647,N_6686,N_11222);
and U17648 (N_17648,N_6349,N_11979);
xor U17649 (N_17649,N_7742,N_12066);
nor U17650 (N_17650,N_7224,N_11623);
and U17651 (N_17651,N_11435,N_11481);
nand U17652 (N_17652,N_11375,N_8002);
and U17653 (N_17653,N_7746,N_10945);
xor U17654 (N_17654,N_11471,N_8032);
nand U17655 (N_17655,N_6890,N_11148);
or U17656 (N_17656,N_8806,N_7416);
and U17657 (N_17657,N_11882,N_6559);
and U17658 (N_17658,N_11606,N_10708);
xor U17659 (N_17659,N_8959,N_8509);
and U17660 (N_17660,N_11983,N_10061);
nor U17661 (N_17661,N_7672,N_10692);
or U17662 (N_17662,N_8781,N_7443);
or U17663 (N_17663,N_10385,N_11627);
xor U17664 (N_17664,N_11131,N_7656);
nor U17665 (N_17665,N_8551,N_10133);
xnor U17666 (N_17666,N_7032,N_8023);
nand U17667 (N_17667,N_9644,N_11035);
and U17668 (N_17668,N_11990,N_10289);
nor U17669 (N_17669,N_9700,N_7383);
or U17670 (N_17670,N_7498,N_11813);
or U17671 (N_17671,N_11513,N_12233);
xor U17672 (N_17672,N_7026,N_9947);
nor U17673 (N_17673,N_7174,N_6674);
nor U17674 (N_17674,N_8600,N_8307);
xnor U17675 (N_17675,N_12478,N_9852);
nor U17676 (N_17676,N_10879,N_10310);
and U17677 (N_17677,N_11930,N_10991);
and U17678 (N_17678,N_12142,N_8637);
nor U17679 (N_17679,N_10702,N_6321);
nor U17680 (N_17680,N_6610,N_6852);
nor U17681 (N_17681,N_9212,N_7252);
or U17682 (N_17682,N_9690,N_8081);
and U17683 (N_17683,N_7575,N_10229);
or U17684 (N_17684,N_6712,N_11971);
or U17685 (N_17685,N_10620,N_7842);
nor U17686 (N_17686,N_8076,N_7326);
xor U17687 (N_17687,N_8658,N_10904);
and U17688 (N_17688,N_11384,N_9987);
and U17689 (N_17689,N_11691,N_12373);
xor U17690 (N_17690,N_12196,N_12164);
xnor U17691 (N_17691,N_12076,N_9350);
xnor U17692 (N_17692,N_12441,N_8871);
and U17693 (N_17693,N_11538,N_12012);
nor U17694 (N_17694,N_7696,N_10240);
or U17695 (N_17695,N_9612,N_8168);
or U17696 (N_17696,N_9130,N_10977);
and U17697 (N_17697,N_10425,N_10465);
nand U17698 (N_17698,N_8206,N_7606);
nor U17699 (N_17699,N_9369,N_10701);
nand U17700 (N_17700,N_6449,N_9316);
or U17701 (N_17701,N_9838,N_7594);
and U17702 (N_17702,N_12070,N_11457);
and U17703 (N_17703,N_7445,N_10147);
xnor U17704 (N_17704,N_7481,N_10564);
xnor U17705 (N_17705,N_10070,N_9086);
or U17706 (N_17706,N_9696,N_11892);
nand U17707 (N_17707,N_11672,N_11188);
and U17708 (N_17708,N_9614,N_7502);
nand U17709 (N_17709,N_6389,N_6551);
or U17710 (N_17710,N_8119,N_9162);
or U17711 (N_17711,N_9629,N_6269);
nand U17712 (N_17712,N_7204,N_11606);
or U17713 (N_17713,N_8894,N_8211);
nor U17714 (N_17714,N_8900,N_12051);
nor U17715 (N_17715,N_8457,N_11220);
nand U17716 (N_17716,N_10429,N_8342);
or U17717 (N_17717,N_11366,N_7722);
xor U17718 (N_17718,N_7109,N_8961);
nand U17719 (N_17719,N_12102,N_9100);
nor U17720 (N_17720,N_7021,N_6507);
nand U17721 (N_17721,N_6392,N_12179);
or U17722 (N_17722,N_7094,N_8464);
nor U17723 (N_17723,N_6931,N_9789);
or U17724 (N_17724,N_11110,N_7156);
nor U17725 (N_17725,N_11808,N_9929);
nand U17726 (N_17726,N_10350,N_8093);
nand U17727 (N_17727,N_10415,N_12021);
and U17728 (N_17728,N_11868,N_8475);
and U17729 (N_17729,N_9037,N_9650);
and U17730 (N_17730,N_9827,N_7253);
or U17731 (N_17731,N_7533,N_9502);
nor U17732 (N_17732,N_8627,N_7848);
xor U17733 (N_17733,N_11648,N_7154);
xor U17734 (N_17734,N_11090,N_10127);
xnor U17735 (N_17735,N_8710,N_6917);
nand U17736 (N_17736,N_6893,N_11265);
or U17737 (N_17737,N_9267,N_7746);
nand U17738 (N_17738,N_10386,N_12232);
xor U17739 (N_17739,N_9642,N_12013);
or U17740 (N_17740,N_9610,N_11438);
xor U17741 (N_17741,N_7281,N_7926);
xor U17742 (N_17742,N_8225,N_12373);
or U17743 (N_17743,N_10421,N_6743);
or U17744 (N_17744,N_7275,N_7310);
nor U17745 (N_17745,N_6804,N_10287);
nor U17746 (N_17746,N_8866,N_10284);
xor U17747 (N_17747,N_9384,N_8852);
or U17748 (N_17748,N_8174,N_9471);
nand U17749 (N_17749,N_9983,N_12450);
or U17750 (N_17750,N_11915,N_11813);
or U17751 (N_17751,N_11185,N_8304);
and U17752 (N_17752,N_8624,N_8753);
xnor U17753 (N_17753,N_6690,N_9598);
nand U17754 (N_17754,N_7305,N_7942);
and U17755 (N_17755,N_8251,N_8116);
nand U17756 (N_17756,N_7320,N_7139);
nand U17757 (N_17757,N_10767,N_10023);
xor U17758 (N_17758,N_7350,N_8700);
nand U17759 (N_17759,N_11334,N_11652);
and U17760 (N_17760,N_6502,N_10054);
or U17761 (N_17761,N_10316,N_6575);
nor U17762 (N_17762,N_6260,N_9600);
or U17763 (N_17763,N_9350,N_8044);
nor U17764 (N_17764,N_10536,N_6509);
nand U17765 (N_17765,N_12467,N_6342);
nand U17766 (N_17766,N_8884,N_7678);
and U17767 (N_17767,N_7497,N_10451);
nand U17768 (N_17768,N_8448,N_9658);
and U17769 (N_17769,N_10716,N_10470);
xnor U17770 (N_17770,N_6976,N_10464);
nor U17771 (N_17771,N_11473,N_11908);
xnor U17772 (N_17772,N_9543,N_8175);
nor U17773 (N_17773,N_8379,N_9510);
or U17774 (N_17774,N_8918,N_8954);
and U17775 (N_17775,N_7650,N_12417);
and U17776 (N_17776,N_7336,N_6418);
xor U17777 (N_17777,N_7284,N_6757);
xor U17778 (N_17778,N_8436,N_10699);
nand U17779 (N_17779,N_11047,N_10257);
or U17780 (N_17780,N_10811,N_8877);
xor U17781 (N_17781,N_8365,N_7434);
and U17782 (N_17782,N_9727,N_10005);
nor U17783 (N_17783,N_11624,N_9857);
xor U17784 (N_17784,N_10826,N_6621);
nand U17785 (N_17785,N_7282,N_9420);
nor U17786 (N_17786,N_10352,N_6450);
and U17787 (N_17787,N_7564,N_12018);
nand U17788 (N_17788,N_11354,N_9488);
xnor U17789 (N_17789,N_7255,N_8798);
xor U17790 (N_17790,N_8496,N_7086);
and U17791 (N_17791,N_7006,N_11279);
nor U17792 (N_17792,N_12368,N_10210);
nor U17793 (N_17793,N_11329,N_7538);
and U17794 (N_17794,N_12287,N_9948);
or U17795 (N_17795,N_6490,N_7327);
nor U17796 (N_17796,N_10938,N_8252);
nand U17797 (N_17797,N_6591,N_7863);
and U17798 (N_17798,N_7674,N_8893);
xnor U17799 (N_17799,N_11294,N_8415);
nand U17800 (N_17800,N_11394,N_9261);
nor U17801 (N_17801,N_10586,N_7607);
nor U17802 (N_17802,N_7498,N_8608);
nor U17803 (N_17803,N_6694,N_10038);
or U17804 (N_17804,N_7725,N_11846);
xnor U17805 (N_17805,N_8183,N_12317);
and U17806 (N_17806,N_12430,N_7688);
nand U17807 (N_17807,N_9698,N_7035);
and U17808 (N_17808,N_6412,N_6380);
xor U17809 (N_17809,N_11969,N_6701);
and U17810 (N_17810,N_10892,N_12494);
nor U17811 (N_17811,N_8962,N_10437);
nand U17812 (N_17812,N_7890,N_11573);
nor U17813 (N_17813,N_8988,N_9369);
or U17814 (N_17814,N_8709,N_10907);
and U17815 (N_17815,N_7039,N_6341);
or U17816 (N_17816,N_11593,N_8049);
or U17817 (N_17817,N_10734,N_6428);
nor U17818 (N_17818,N_9301,N_7190);
xor U17819 (N_17819,N_6601,N_8545);
nor U17820 (N_17820,N_9128,N_11056);
or U17821 (N_17821,N_12338,N_6846);
nor U17822 (N_17822,N_11966,N_9564);
or U17823 (N_17823,N_7859,N_10791);
nand U17824 (N_17824,N_8956,N_10993);
nand U17825 (N_17825,N_6979,N_12395);
xor U17826 (N_17826,N_8244,N_6716);
xnor U17827 (N_17827,N_8841,N_11999);
xor U17828 (N_17828,N_7398,N_6962);
and U17829 (N_17829,N_7618,N_11331);
nor U17830 (N_17830,N_8313,N_11065);
nand U17831 (N_17831,N_6772,N_12342);
nand U17832 (N_17832,N_10662,N_10315);
nor U17833 (N_17833,N_10562,N_10970);
nor U17834 (N_17834,N_8384,N_7719);
or U17835 (N_17835,N_11110,N_7454);
nor U17836 (N_17836,N_10020,N_7531);
xnor U17837 (N_17837,N_8761,N_10627);
xor U17838 (N_17838,N_9079,N_8546);
or U17839 (N_17839,N_12267,N_6661);
nand U17840 (N_17840,N_8979,N_10500);
nand U17841 (N_17841,N_11596,N_9488);
and U17842 (N_17842,N_11174,N_8408);
xnor U17843 (N_17843,N_6693,N_7159);
nor U17844 (N_17844,N_12286,N_12389);
xor U17845 (N_17845,N_11154,N_10256);
and U17846 (N_17846,N_8613,N_6285);
xnor U17847 (N_17847,N_8664,N_7082);
or U17848 (N_17848,N_9469,N_7414);
nor U17849 (N_17849,N_8274,N_8375);
xor U17850 (N_17850,N_9362,N_8605);
or U17851 (N_17851,N_9017,N_6361);
and U17852 (N_17852,N_9275,N_8759);
nor U17853 (N_17853,N_10697,N_12296);
and U17854 (N_17854,N_11482,N_6499);
nor U17855 (N_17855,N_6461,N_9886);
xor U17856 (N_17856,N_7373,N_11246);
and U17857 (N_17857,N_11519,N_9039);
xor U17858 (N_17858,N_7380,N_8172);
and U17859 (N_17859,N_9169,N_9044);
xor U17860 (N_17860,N_10306,N_9042);
nand U17861 (N_17861,N_10646,N_7620);
nor U17862 (N_17862,N_6865,N_11640);
nand U17863 (N_17863,N_10383,N_12368);
and U17864 (N_17864,N_11157,N_8713);
nor U17865 (N_17865,N_9706,N_6327);
xor U17866 (N_17866,N_7762,N_8150);
xnor U17867 (N_17867,N_10393,N_9059);
xor U17868 (N_17868,N_9186,N_8361);
nor U17869 (N_17869,N_11199,N_11893);
and U17870 (N_17870,N_6973,N_10508);
and U17871 (N_17871,N_9638,N_9230);
nand U17872 (N_17872,N_9388,N_6775);
or U17873 (N_17873,N_10847,N_9760);
xor U17874 (N_17874,N_7200,N_7813);
or U17875 (N_17875,N_9578,N_7282);
nor U17876 (N_17876,N_11102,N_11873);
and U17877 (N_17877,N_7784,N_8037);
xor U17878 (N_17878,N_12185,N_10630);
nor U17879 (N_17879,N_10439,N_9635);
nor U17880 (N_17880,N_7948,N_11746);
nand U17881 (N_17881,N_11494,N_9253);
xor U17882 (N_17882,N_9854,N_9126);
and U17883 (N_17883,N_10511,N_8054);
nor U17884 (N_17884,N_12059,N_12160);
or U17885 (N_17885,N_8619,N_10735);
and U17886 (N_17886,N_9089,N_9935);
or U17887 (N_17887,N_11370,N_9436);
nand U17888 (N_17888,N_7602,N_9868);
or U17889 (N_17889,N_11057,N_11814);
or U17890 (N_17890,N_11589,N_11859);
nand U17891 (N_17891,N_12037,N_7502);
and U17892 (N_17892,N_6327,N_7438);
xor U17893 (N_17893,N_10114,N_11585);
nand U17894 (N_17894,N_8193,N_12052);
or U17895 (N_17895,N_10421,N_8366);
nor U17896 (N_17896,N_11238,N_12356);
xor U17897 (N_17897,N_7835,N_6848);
nand U17898 (N_17898,N_10581,N_8462);
and U17899 (N_17899,N_7053,N_11249);
or U17900 (N_17900,N_8965,N_10900);
and U17901 (N_17901,N_9185,N_12127);
or U17902 (N_17902,N_11990,N_12111);
and U17903 (N_17903,N_7947,N_10043);
or U17904 (N_17904,N_6666,N_10986);
and U17905 (N_17905,N_10461,N_9591);
xnor U17906 (N_17906,N_10796,N_12335);
or U17907 (N_17907,N_7406,N_6806);
nand U17908 (N_17908,N_9516,N_9225);
or U17909 (N_17909,N_8355,N_11723);
or U17910 (N_17910,N_9615,N_7169);
and U17911 (N_17911,N_10946,N_7582);
nand U17912 (N_17912,N_11435,N_6320);
nand U17913 (N_17913,N_8155,N_10432);
nor U17914 (N_17914,N_7770,N_7756);
nor U17915 (N_17915,N_10986,N_7226);
or U17916 (N_17916,N_7585,N_9073);
nor U17917 (N_17917,N_7807,N_10817);
nand U17918 (N_17918,N_6295,N_10738);
xnor U17919 (N_17919,N_9092,N_7511);
nor U17920 (N_17920,N_8586,N_9153);
nor U17921 (N_17921,N_9812,N_9905);
nand U17922 (N_17922,N_9124,N_11858);
or U17923 (N_17923,N_8126,N_6447);
and U17924 (N_17924,N_11731,N_11349);
and U17925 (N_17925,N_10503,N_11105);
nand U17926 (N_17926,N_8067,N_12152);
or U17927 (N_17927,N_11121,N_9259);
xnor U17928 (N_17928,N_8183,N_8597);
nand U17929 (N_17929,N_11771,N_8863);
nor U17930 (N_17930,N_7580,N_11157);
and U17931 (N_17931,N_9233,N_7449);
xnor U17932 (N_17932,N_7057,N_8560);
and U17933 (N_17933,N_12440,N_9392);
nor U17934 (N_17934,N_8153,N_6632);
or U17935 (N_17935,N_11389,N_7672);
and U17936 (N_17936,N_11652,N_9012);
xor U17937 (N_17937,N_12306,N_10142);
nor U17938 (N_17938,N_9384,N_12013);
xor U17939 (N_17939,N_7980,N_9641);
xor U17940 (N_17940,N_10999,N_7591);
or U17941 (N_17941,N_7368,N_8968);
and U17942 (N_17942,N_12062,N_12269);
nand U17943 (N_17943,N_12229,N_8687);
and U17944 (N_17944,N_8639,N_6577);
or U17945 (N_17945,N_9679,N_7781);
nor U17946 (N_17946,N_6577,N_7803);
nand U17947 (N_17947,N_9171,N_10035);
nor U17948 (N_17948,N_10616,N_9610);
or U17949 (N_17949,N_7232,N_10292);
nand U17950 (N_17950,N_12068,N_10378);
nand U17951 (N_17951,N_10273,N_11985);
nor U17952 (N_17952,N_11313,N_11432);
xnor U17953 (N_17953,N_8770,N_8274);
or U17954 (N_17954,N_7161,N_6911);
nor U17955 (N_17955,N_7555,N_12408);
xnor U17956 (N_17956,N_11256,N_11275);
nand U17957 (N_17957,N_6612,N_7012);
nor U17958 (N_17958,N_9505,N_10699);
nor U17959 (N_17959,N_9027,N_7186);
or U17960 (N_17960,N_12455,N_7183);
nand U17961 (N_17961,N_9291,N_7458);
and U17962 (N_17962,N_7862,N_7214);
nand U17963 (N_17963,N_9021,N_10918);
and U17964 (N_17964,N_9005,N_10451);
and U17965 (N_17965,N_8745,N_8293);
nor U17966 (N_17966,N_9975,N_10693);
or U17967 (N_17967,N_8857,N_11797);
and U17968 (N_17968,N_11951,N_6305);
and U17969 (N_17969,N_7573,N_10474);
nand U17970 (N_17970,N_10890,N_6748);
nor U17971 (N_17971,N_6399,N_10249);
nand U17972 (N_17972,N_8966,N_8156);
or U17973 (N_17973,N_12053,N_6534);
xor U17974 (N_17974,N_10937,N_7068);
nand U17975 (N_17975,N_9855,N_11327);
and U17976 (N_17976,N_6609,N_6422);
and U17977 (N_17977,N_10811,N_6416);
nand U17978 (N_17978,N_9146,N_7390);
nand U17979 (N_17979,N_7147,N_7733);
nor U17980 (N_17980,N_8081,N_6844);
xor U17981 (N_17981,N_7429,N_9547);
nor U17982 (N_17982,N_11241,N_8365);
nand U17983 (N_17983,N_10699,N_6744);
nor U17984 (N_17984,N_9627,N_12068);
nor U17985 (N_17985,N_11563,N_10444);
xnor U17986 (N_17986,N_10371,N_8841);
and U17987 (N_17987,N_6900,N_8281);
nand U17988 (N_17988,N_10136,N_11094);
nand U17989 (N_17989,N_7854,N_7258);
or U17990 (N_17990,N_10060,N_11346);
xnor U17991 (N_17991,N_10084,N_7573);
xnor U17992 (N_17992,N_8430,N_10588);
xor U17993 (N_17993,N_10448,N_9807);
nor U17994 (N_17994,N_8477,N_11273);
xnor U17995 (N_17995,N_6575,N_9919);
or U17996 (N_17996,N_11300,N_11383);
xor U17997 (N_17997,N_11264,N_8640);
nand U17998 (N_17998,N_8195,N_9250);
or U17999 (N_17999,N_12239,N_7399);
and U18000 (N_18000,N_10400,N_9323);
or U18001 (N_18001,N_7085,N_9280);
and U18002 (N_18002,N_10724,N_7500);
nand U18003 (N_18003,N_9053,N_11958);
or U18004 (N_18004,N_7961,N_6414);
and U18005 (N_18005,N_12095,N_11185);
or U18006 (N_18006,N_8351,N_11473);
nand U18007 (N_18007,N_11497,N_10056);
and U18008 (N_18008,N_10111,N_11130);
nor U18009 (N_18009,N_10166,N_6944);
nand U18010 (N_18010,N_11944,N_9445);
nand U18011 (N_18011,N_7679,N_10687);
nor U18012 (N_18012,N_11748,N_8377);
nor U18013 (N_18013,N_7681,N_12303);
or U18014 (N_18014,N_12025,N_11563);
nor U18015 (N_18015,N_8686,N_10067);
or U18016 (N_18016,N_6418,N_10060);
nand U18017 (N_18017,N_7790,N_11905);
or U18018 (N_18018,N_8038,N_12305);
nand U18019 (N_18019,N_7865,N_8704);
xor U18020 (N_18020,N_7722,N_11230);
or U18021 (N_18021,N_8061,N_8147);
or U18022 (N_18022,N_12016,N_8871);
nor U18023 (N_18023,N_9830,N_11637);
nor U18024 (N_18024,N_6387,N_9516);
and U18025 (N_18025,N_10495,N_7598);
xnor U18026 (N_18026,N_9726,N_8417);
nor U18027 (N_18027,N_10580,N_7938);
or U18028 (N_18028,N_10700,N_8707);
nand U18029 (N_18029,N_11823,N_9984);
and U18030 (N_18030,N_12190,N_8791);
nor U18031 (N_18031,N_7551,N_7215);
nor U18032 (N_18032,N_9890,N_12137);
nand U18033 (N_18033,N_6459,N_7580);
nor U18034 (N_18034,N_10106,N_9282);
nor U18035 (N_18035,N_6979,N_8321);
xor U18036 (N_18036,N_7498,N_11155);
xnor U18037 (N_18037,N_10458,N_8354);
or U18038 (N_18038,N_6597,N_9475);
nor U18039 (N_18039,N_7267,N_9553);
xor U18040 (N_18040,N_12411,N_11981);
and U18041 (N_18041,N_8745,N_9036);
nor U18042 (N_18042,N_8429,N_11418);
or U18043 (N_18043,N_12297,N_6753);
nor U18044 (N_18044,N_10350,N_7790);
nand U18045 (N_18045,N_10425,N_12416);
and U18046 (N_18046,N_7568,N_11996);
nor U18047 (N_18047,N_11770,N_8129);
and U18048 (N_18048,N_12387,N_9784);
nor U18049 (N_18049,N_10775,N_12050);
xnor U18050 (N_18050,N_9148,N_9044);
and U18051 (N_18051,N_12075,N_10593);
or U18052 (N_18052,N_11000,N_11282);
or U18053 (N_18053,N_11945,N_6459);
and U18054 (N_18054,N_8528,N_9224);
and U18055 (N_18055,N_10377,N_8511);
and U18056 (N_18056,N_6481,N_10778);
xnor U18057 (N_18057,N_6659,N_11111);
or U18058 (N_18058,N_10181,N_6465);
or U18059 (N_18059,N_12167,N_11376);
nand U18060 (N_18060,N_7214,N_10587);
nand U18061 (N_18061,N_9025,N_9669);
nand U18062 (N_18062,N_10694,N_10091);
or U18063 (N_18063,N_9785,N_12139);
xor U18064 (N_18064,N_11055,N_11001);
xnor U18065 (N_18065,N_7247,N_8980);
and U18066 (N_18066,N_9657,N_12040);
xnor U18067 (N_18067,N_7583,N_7772);
xor U18068 (N_18068,N_12054,N_7250);
nor U18069 (N_18069,N_8506,N_9778);
nor U18070 (N_18070,N_8411,N_9846);
and U18071 (N_18071,N_11070,N_10570);
xor U18072 (N_18072,N_6494,N_9337);
or U18073 (N_18073,N_11549,N_9948);
xor U18074 (N_18074,N_8102,N_12348);
xor U18075 (N_18075,N_10874,N_11815);
xnor U18076 (N_18076,N_10744,N_10522);
nand U18077 (N_18077,N_7142,N_7824);
xnor U18078 (N_18078,N_12172,N_11941);
and U18079 (N_18079,N_8065,N_9695);
nor U18080 (N_18080,N_10448,N_9974);
nor U18081 (N_18081,N_10685,N_11043);
xor U18082 (N_18082,N_9687,N_11782);
or U18083 (N_18083,N_9585,N_10466);
xnor U18084 (N_18084,N_7577,N_11586);
and U18085 (N_18085,N_9724,N_11832);
nand U18086 (N_18086,N_11557,N_9260);
xnor U18087 (N_18087,N_11561,N_8391);
nor U18088 (N_18088,N_8679,N_7095);
nor U18089 (N_18089,N_6275,N_10730);
xor U18090 (N_18090,N_9644,N_11218);
nand U18091 (N_18091,N_9954,N_12166);
or U18092 (N_18092,N_10574,N_7892);
nand U18093 (N_18093,N_11549,N_9825);
and U18094 (N_18094,N_9019,N_12131);
or U18095 (N_18095,N_11331,N_11903);
xor U18096 (N_18096,N_10700,N_7335);
nor U18097 (N_18097,N_11350,N_11289);
nand U18098 (N_18098,N_11118,N_7970);
and U18099 (N_18099,N_8725,N_10405);
nor U18100 (N_18100,N_11169,N_11496);
or U18101 (N_18101,N_9158,N_11145);
xnor U18102 (N_18102,N_7181,N_8616);
and U18103 (N_18103,N_7332,N_10330);
nand U18104 (N_18104,N_11054,N_6262);
nor U18105 (N_18105,N_9167,N_10105);
nand U18106 (N_18106,N_6788,N_6442);
and U18107 (N_18107,N_8353,N_10836);
or U18108 (N_18108,N_12451,N_10357);
and U18109 (N_18109,N_11383,N_11255);
nor U18110 (N_18110,N_10588,N_11748);
and U18111 (N_18111,N_11130,N_8440);
xor U18112 (N_18112,N_7911,N_10858);
nor U18113 (N_18113,N_7586,N_11753);
and U18114 (N_18114,N_8676,N_11938);
or U18115 (N_18115,N_10477,N_12304);
nor U18116 (N_18116,N_10494,N_10357);
or U18117 (N_18117,N_7444,N_8803);
or U18118 (N_18118,N_8331,N_11769);
nor U18119 (N_18119,N_12005,N_9860);
and U18120 (N_18120,N_8454,N_10200);
nand U18121 (N_18121,N_7198,N_12113);
nor U18122 (N_18122,N_9129,N_10853);
and U18123 (N_18123,N_6461,N_10859);
or U18124 (N_18124,N_10478,N_12083);
or U18125 (N_18125,N_6946,N_8634);
nor U18126 (N_18126,N_6530,N_7272);
xnor U18127 (N_18127,N_9360,N_7374);
xnor U18128 (N_18128,N_10858,N_10589);
or U18129 (N_18129,N_9606,N_12436);
nand U18130 (N_18130,N_6454,N_6363);
or U18131 (N_18131,N_11158,N_8664);
nand U18132 (N_18132,N_11979,N_8390);
xnor U18133 (N_18133,N_9497,N_10644);
or U18134 (N_18134,N_10310,N_11431);
nand U18135 (N_18135,N_8970,N_10574);
or U18136 (N_18136,N_11434,N_11097);
nand U18137 (N_18137,N_7054,N_11093);
or U18138 (N_18138,N_10181,N_8483);
or U18139 (N_18139,N_11072,N_12080);
nor U18140 (N_18140,N_9692,N_7635);
xor U18141 (N_18141,N_12490,N_11906);
xnor U18142 (N_18142,N_6947,N_11517);
nor U18143 (N_18143,N_9019,N_9817);
nor U18144 (N_18144,N_8469,N_8594);
xnor U18145 (N_18145,N_12311,N_9786);
xor U18146 (N_18146,N_12213,N_11925);
nor U18147 (N_18147,N_11448,N_10318);
or U18148 (N_18148,N_11679,N_6828);
xor U18149 (N_18149,N_6768,N_10755);
nor U18150 (N_18150,N_10655,N_8444);
nor U18151 (N_18151,N_11704,N_10235);
nand U18152 (N_18152,N_7683,N_11146);
nand U18153 (N_18153,N_11996,N_11647);
nor U18154 (N_18154,N_8047,N_10331);
nor U18155 (N_18155,N_7103,N_12168);
xnor U18156 (N_18156,N_10746,N_11151);
nor U18157 (N_18157,N_8384,N_10064);
nor U18158 (N_18158,N_9353,N_10378);
nand U18159 (N_18159,N_6697,N_6814);
nand U18160 (N_18160,N_10570,N_11339);
xnor U18161 (N_18161,N_8025,N_7274);
or U18162 (N_18162,N_6491,N_11763);
xnor U18163 (N_18163,N_9769,N_9972);
and U18164 (N_18164,N_8953,N_8592);
and U18165 (N_18165,N_10078,N_9952);
nor U18166 (N_18166,N_8448,N_12252);
and U18167 (N_18167,N_8384,N_7795);
and U18168 (N_18168,N_6957,N_9146);
xor U18169 (N_18169,N_7860,N_11007);
xor U18170 (N_18170,N_10760,N_9517);
nor U18171 (N_18171,N_9493,N_11012);
nand U18172 (N_18172,N_11913,N_9975);
nor U18173 (N_18173,N_8756,N_7308);
nor U18174 (N_18174,N_11174,N_7118);
or U18175 (N_18175,N_6531,N_8443);
or U18176 (N_18176,N_9087,N_7591);
and U18177 (N_18177,N_11889,N_9121);
xor U18178 (N_18178,N_9313,N_8318);
or U18179 (N_18179,N_12150,N_7949);
nand U18180 (N_18180,N_8530,N_8180);
nand U18181 (N_18181,N_10846,N_9339);
or U18182 (N_18182,N_7697,N_8654);
nand U18183 (N_18183,N_8047,N_11867);
nor U18184 (N_18184,N_7113,N_11124);
nand U18185 (N_18185,N_8140,N_8569);
or U18186 (N_18186,N_12474,N_7407);
nand U18187 (N_18187,N_8345,N_8763);
and U18188 (N_18188,N_7024,N_9300);
or U18189 (N_18189,N_10988,N_7176);
xnor U18190 (N_18190,N_10974,N_9166);
and U18191 (N_18191,N_11913,N_7657);
nand U18192 (N_18192,N_9471,N_9194);
nor U18193 (N_18193,N_7365,N_10024);
xor U18194 (N_18194,N_10457,N_8238);
or U18195 (N_18195,N_9393,N_8073);
nor U18196 (N_18196,N_10140,N_8884);
xor U18197 (N_18197,N_10101,N_6728);
xor U18198 (N_18198,N_11916,N_7287);
nand U18199 (N_18199,N_12035,N_10057);
nor U18200 (N_18200,N_10658,N_8783);
and U18201 (N_18201,N_9036,N_8261);
xnor U18202 (N_18202,N_11098,N_6353);
nor U18203 (N_18203,N_10619,N_8343);
xor U18204 (N_18204,N_7310,N_7685);
nand U18205 (N_18205,N_12412,N_9959);
nor U18206 (N_18206,N_9234,N_7201);
nor U18207 (N_18207,N_9124,N_9660);
xor U18208 (N_18208,N_7830,N_12483);
and U18209 (N_18209,N_8511,N_9053);
nand U18210 (N_18210,N_12121,N_8119);
xnor U18211 (N_18211,N_9654,N_9092);
xor U18212 (N_18212,N_7338,N_8314);
and U18213 (N_18213,N_10542,N_10461);
nand U18214 (N_18214,N_6810,N_6794);
nand U18215 (N_18215,N_10195,N_9230);
nor U18216 (N_18216,N_7633,N_8779);
nand U18217 (N_18217,N_6295,N_11034);
nand U18218 (N_18218,N_6749,N_9560);
nand U18219 (N_18219,N_7404,N_9129);
xor U18220 (N_18220,N_6592,N_7514);
and U18221 (N_18221,N_8850,N_7893);
nand U18222 (N_18222,N_6946,N_9812);
nor U18223 (N_18223,N_8903,N_6992);
nor U18224 (N_18224,N_12009,N_7732);
or U18225 (N_18225,N_7418,N_11504);
nor U18226 (N_18226,N_12395,N_11724);
nor U18227 (N_18227,N_8691,N_11842);
nor U18228 (N_18228,N_8522,N_9703);
nor U18229 (N_18229,N_10433,N_10990);
nand U18230 (N_18230,N_6875,N_6589);
nand U18231 (N_18231,N_7755,N_7582);
or U18232 (N_18232,N_7193,N_10008);
xor U18233 (N_18233,N_8469,N_9346);
xnor U18234 (N_18234,N_10729,N_9974);
or U18235 (N_18235,N_7883,N_10780);
and U18236 (N_18236,N_10558,N_9812);
nor U18237 (N_18237,N_10788,N_8507);
nor U18238 (N_18238,N_10623,N_8109);
nand U18239 (N_18239,N_11706,N_12469);
or U18240 (N_18240,N_12425,N_8915);
nor U18241 (N_18241,N_8777,N_9393);
and U18242 (N_18242,N_6926,N_10880);
nor U18243 (N_18243,N_6615,N_8374);
xnor U18244 (N_18244,N_8722,N_10858);
nand U18245 (N_18245,N_10980,N_9259);
nor U18246 (N_18246,N_11293,N_10512);
xnor U18247 (N_18247,N_12324,N_12366);
or U18248 (N_18248,N_10821,N_10217);
or U18249 (N_18249,N_9569,N_8088);
nor U18250 (N_18250,N_10928,N_9811);
nor U18251 (N_18251,N_9888,N_10864);
nor U18252 (N_18252,N_10053,N_9917);
xor U18253 (N_18253,N_10957,N_9861);
xor U18254 (N_18254,N_9666,N_6325);
or U18255 (N_18255,N_9245,N_11646);
nor U18256 (N_18256,N_7151,N_12261);
nand U18257 (N_18257,N_6338,N_7600);
nor U18258 (N_18258,N_6938,N_11359);
or U18259 (N_18259,N_8551,N_6729);
xnor U18260 (N_18260,N_7471,N_12175);
nand U18261 (N_18261,N_10444,N_10539);
xor U18262 (N_18262,N_10352,N_8342);
and U18263 (N_18263,N_7220,N_10308);
or U18264 (N_18264,N_7403,N_8670);
nor U18265 (N_18265,N_7337,N_9835);
nor U18266 (N_18266,N_6940,N_12307);
nand U18267 (N_18267,N_12430,N_6355);
or U18268 (N_18268,N_8415,N_10910);
nor U18269 (N_18269,N_9688,N_9860);
nor U18270 (N_18270,N_7432,N_12479);
nand U18271 (N_18271,N_9004,N_9017);
or U18272 (N_18272,N_8957,N_7218);
nor U18273 (N_18273,N_10318,N_12015);
and U18274 (N_18274,N_7849,N_10870);
xor U18275 (N_18275,N_11933,N_6929);
or U18276 (N_18276,N_9382,N_10224);
xnor U18277 (N_18277,N_6687,N_6862);
xnor U18278 (N_18278,N_11538,N_6312);
and U18279 (N_18279,N_6373,N_10472);
nand U18280 (N_18280,N_6395,N_11038);
or U18281 (N_18281,N_9870,N_8066);
nor U18282 (N_18282,N_10157,N_6845);
or U18283 (N_18283,N_10795,N_11270);
nand U18284 (N_18284,N_9327,N_12319);
nand U18285 (N_18285,N_12434,N_10199);
and U18286 (N_18286,N_6313,N_6459);
or U18287 (N_18287,N_11552,N_11558);
nor U18288 (N_18288,N_10338,N_6938);
xor U18289 (N_18289,N_10461,N_6615);
xnor U18290 (N_18290,N_9415,N_10060);
and U18291 (N_18291,N_8924,N_6850);
xnor U18292 (N_18292,N_11627,N_11035);
xor U18293 (N_18293,N_10770,N_6526);
nor U18294 (N_18294,N_11340,N_9806);
and U18295 (N_18295,N_7951,N_6852);
nor U18296 (N_18296,N_11484,N_12088);
and U18297 (N_18297,N_7643,N_6276);
or U18298 (N_18298,N_11406,N_7201);
nand U18299 (N_18299,N_11121,N_12096);
or U18300 (N_18300,N_6558,N_11815);
and U18301 (N_18301,N_9022,N_8288);
nor U18302 (N_18302,N_7799,N_11612);
or U18303 (N_18303,N_10393,N_7098);
nand U18304 (N_18304,N_10393,N_10556);
nor U18305 (N_18305,N_10641,N_10653);
or U18306 (N_18306,N_9773,N_7057);
nor U18307 (N_18307,N_11905,N_7268);
nand U18308 (N_18308,N_9822,N_10716);
nor U18309 (N_18309,N_6965,N_9817);
or U18310 (N_18310,N_11708,N_7492);
and U18311 (N_18311,N_8827,N_8318);
or U18312 (N_18312,N_10616,N_11446);
xnor U18313 (N_18313,N_10496,N_8932);
or U18314 (N_18314,N_8121,N_10729);
or U18315 (N_18315,N_6861,N_8445);
xor U18316 (N_18316,N_8488,N_12474);
and U18317 (N_18317,N_12129,N_11913);
nand U18318 (N_18318,N_11607,N_12070);
xnor U18319 (N_18319,N_10138,N_8832);
and U18320 (N_18320,N_8442,N_12053);
xor U18321 (N_18321,N_9531,N_11389);
and U18322 (N_18322,N_12182,N_9585);
xnor U18323 (N_18323,N_7074,N_6580);
nand U18324 (N_18324,N_9078,N_8818);
or U18325 (N_18325,N_7037,N_11861);
nor U18326 (N_18326,N_12234,N_10353);
nand U18327 (N_18327,N_11905,N_7537);
and U18328 (N_18328,N_8603,N_10694);
and U18329 (N_18329,N_8748,N_11443);
and U18330 (N_18330,N_6830,N_11704);
nand U18331 (N_18331,N_8749,N_12113);
nand U18332 (N_18332,N_10367,N_6762);
or U18333 (N_18333,N_7188,N_6265);
nand U18334 (N_18334,N_10338,N_12101);
or U18335 (N_18335,N_8155,N_8511);
xor U18336 (N_18336,N_10864,N_11483);
nand U18337 (N_18337,N_9280,N_7927);
xor U18338 (N_18338,N_6256,N_7948);
and U18339 (N_18339,N_9795,N_9136);
or U18340 (N_18340,N_10124,N_8997);
nand U18341 (N_18341,N_7567,N_6786);
and U18342 (N_18342,N_9001,N_11897);
nand U18343 (N_18343,N_8605,N_6717);
xnor U18344 (N_18344,N_11547,N_9642);
xnor U18345 (N_18345,N_9114,N_11810);
nor U18346 (N_18346,N_6522,N_11936);
and U18347 (N_18347,N_11463,N_10842);
or U18348 (N_18348,N_9392,N_10052);
nand U18349 (N_18349,N_6969,N_6798);
nor U18350 (N_18350,N_8882,N_12241);
xnor U18351 (N_18351,N_11338,N_6974);
nor U18352 (N_18352,N_11023,N_9591);
or U18353 (N_18353,N_6250,N_10557);
xnor U18354 (N_18354,N_10906,N_10523);
or U18355 (N_18355,N_9658,N_11082);
nor U18356 (N_18356,N_12275,N_7219);
xor U18357 (N_18357,N_8272,N_7005);
and U18358 (N_18358,N_10591,N_11664);
or U18359 (N_18359,N_8524,N_6949);
xnor U18360 (N_18360,N_8746,N_7728);
and U18361 (N_18361,N_6318,N_8135);
nand U18362 (N_18362,N_11434,N_8328);
xnor U18363 (N_18363,N_7830,N_11727);
and U18364 (N_18364,N_7701,N_8595);
or U18365 (N_18365,N_10975,N_12008);
or U18366 (N_18366,N_10090,N_10027);
nor U18367 (N_18367,N_9408,N_6425);
or U18368 (N_18368,N_8192,N_10505);
nor U18369 (N_18369,N_7052,N_6836);
or U18370 (N_18370,N_6497,N_8753);
xnor U18371 (N_18371,N_11133,N_6715);
nand U18372 (N_18372,N_6310,N_8261);
and U18373 (N_18373,N_9406,N_12323);
xnor U18374 (N_18374,N_7226,N_12129);
nor U18375 (N_18375,N_12156,N_7180);
xor U18376 (N_18376,N_8819,N_7222);
nand U18377 (N_18377,N_10725,N_10798);
nand U18378 (N_18378,N_6682,N_10810);
nor U18379 (N_18379,N_10411,N_10152);
xnor U18380 (N_18380,N_8612,N_8088);
and U18381 (N_18381,N_11744,N_9886);
nor U18382 (N_18382,N_11034,N_7440);
xor U18383 (N_18383,N_12342,N_8580);
xor U18384 (N_18384,N_9842,N_11597);
and U18385 (N_18385,N_8614,N_8960);
xnor U18386 (N_18386,N_10081,N_11206);
or U18387 (N_18387,N_10021,N_10963);
nand U18388 (N_18388,N_11256,N_11213);
nand U18389 (N_18389,N_11329,N_9701);
or U18390 (N_18390,N_9940,N_11835);
nand U18391 (N_18391,N_7530,N_11372);
and U18392 (N_18392,N_7301,N_7581);
xnor U18393 (N_18393,N_11283,N_8608);
nand U18394 (N_18394,N_11063,N_7984);
xnor U18395 (N_18395,N_9358,N_7407);
and U18396 (N_18396,N_7134,N_6364);
and U18397 (N_18397,N_12325,N_11891);
or U18398 (N_18398,N_8205,N_10210);
nand U18399 (N_18399,N_8756,N_11741);
xnor U18400 (N_18400,N_8302,N_8631);
or U18401 (N_18401,N_10340,N_6867);
and U18402 (N_18402,N_9359,N_7620);
nand U18403 (N_18403,N_6577,N_7810);
and U18404 (N_18404,N_9999,N_11815);
nor U18405 (N_18405,N_11856,N_11383);
xor U18406 (N_18406,N_9659,N_10354);
and U18407 (N_18407,N_11684,N_7033);
nor U18408 (N_18408,N_7103,N_10819);
nor U18409 (N_18409,N_8642,N_10473);
and U18410 (N_18410,N_11748,N_9556);
nand U18411 (N_18411,N_8154,N_6458);
or U18412 (N_18412,N_10086,N_8472);
nand U18413 (N_18413,N_11081,N_6981);
or U18414 (N_18414,N_9947,N_9315);
or U18415 (N_18415,N_12318,N_10403);
xnor U18416 (N_18416,N_11527,N_7098);
and U18417 (N_18417,N_6653,N_7990);
or U18418 (N_18418,N_9021,N_12482);
nand U18419 (N_18419,N_9212,N_8511);
nand U18420 (N_18420,N_8935,N_10134);
and U18421 (N_18421,N_7356,N_7414);
nand U18422 (N_18422,N_11481,N_6574);
nor U18423 (N_18423,N_10066,N_9802);
nand U18424 (N_18424,N_8897,N_6661);
nand U18425 (N_18425,N_12201,N_7360);
and U18426 (N_18426,N_11236,N_11032);
and U18427 (N_18427,N_9947,N_6281);
nor U18428 (N_18428,N_6738,N_10365);
or U18429 (N_18429,N_8673,N_11149);
and U18430 (N_18430,N_8218,N_7109);
nor U18431 (N_18431,N_11336,N_7278);
nand U18432 (N_18432,N_11862,N_10230);
and U18433 (N_18433,N_8065,N_11490);
xnor U18434 (N_18434,N_10764,N_6806);
and U18435 (N_18435,N_11047,N_8628);
nor U18436 (N_18436,N_6635,N_9365);
xor U18437 (N_18437,N_11518,N_8033);
nor U18438 (N_18438,N_11273,N_11987);
nor U18439 (N_18439,N_8138,N_11952);
xnor U18440 (N_18440,N_6977,N_10127);
and U18441 (N_18441,N_8574,N_8486);
nor U18442 (N_18442,N_9076,N_12276);
nor U18443 (N_18443,N_11383,N_11095);
xnor U18444 (N_18444,N_10701,N_7432);
nand U18445 (N_18445,N_6264,N_12159);
nor U18446 (N_18446,N_11987,N_10313);
or U18447 (N_18447,N_11323,N_7383);
nand U18448 (N_18448,N_7554,N_6735);
nor U18449 (N_18449,N_9692,N_11507);
and U18450 (N_18450,N_9939,N_7750);
nand U18451 (N_18451,N_10100,N_7339);
xnor U18452 (N_18452,N_10163,N_7873);
or U18453 (N_18453,N_6714,N_11604);
nor U18454 (N_18454,N_8056,N_7720);
xor U18455 (N_18455,N_10849,N_12396);
xor U18456 (N_18456,N_8633,N_11093);
and U18457 (N_18457,N_11565,N_9180);
and U18458 (N_18458,N_10614,N_8044);
nand U18459 (N_18459,N_8332,N_7007);
nor U18460 (N_18460,N_10798,N_6644);
xor U18461 (N_18461,N_8194,N_6475);
xnor U18462 (N_18462,N_8543,N_11199);
nor U18463 (N_18463,N_10946,N_7398);
xor U18464 (N_18464,N_7596,N_11803);
and U18465 (N_18465,N_10201,N_9359);
xnor U18466 (N_18466,N_7716,N_7873);
nand U18467 (N_18467,N_6420,N_11046);
nand U18468 (N_18468,N_7263,N_11706);
nand U18469 (N_18469,N_7633,N_6722);
nand U18470 (N_18470,N_11048,N_12121);
xor U18471 (N_18471,N_10569,N_8502);
nor U18472 (N_18472,N_10748,N_8269);
xnor U18473 (N_18473,N_8885,N_8038);
xnor U18474 (N_18474,N_7378,N_7803);
nand U18475 (N_18475,N_7959,N_7802);
xnor U18476 (N_18476,N_7414,N_7406);
nor U18477 (N_18477,N_10034,N_11143);
nor U18478 (N_18478,N_7777,N_7123);
and U18479 (N_18479,N_7056,N_7005);
nor U18480 (N_18480,N_9201,N_7599);
or U18481 (N_18481,N_9157,N_8973);
nor U18482 (N_18482,N_6989,N_6452);
xor U18483 (N_18483,N_11224,N_7238);
xor U18484 (N_18484,N_11460,N_10160);
or U18485 (N_18485,N_10089,N_11288);
or U18486 (N_18486,N_8653,N_9062);
and U18487 (N_18487,N_10894,N_9331);
and U18488 (N_18488,N_10928,N_11426);
or U18489 (N_18489,N_10356,N_7723);
or U18490 (N_18490,N_7060,N_10884);
and U18491 (N_18491,N_8108,N_8659);
nor U18492 (N_18492,N_9988,N_10270);
nor U18493 (N_18493,N_7273,N_9477);
and U18494 (N_18494,N_10466,N_10985);
nand U18495 (N_18495,N_8586,N_10387);
xor U18496 (N_18496,N_8486,N_8478);
xnor U18497 (N_18497,N_8743,N_8035);
and U18498 (N_18498,N_9931,N_7001);
nand U18499 (N_18499,N_6456,N_10443);
and U18500 (N_18500,N_11490,N_7763);
or U18501 (N_18501,N_10439,N_10730);
nor U18502 (N_18502,N_6574,N_9330);
nand U18503 (N_18503,N_10938,N_11165);
nor U18504 (N_18504,N_12399,N_11787);
nand U18505 (N_18505,N_11359,N_8887);
nand U18506 (N_18506,N_12020,N_11056);
nor U18507 (N_18507,N_7251,N_8171);
xnor U18508 (N_18508,N_6512,N_12343);
nand U18509 (N_18509,N_7925,N_7603);
or U18510 (N_18510,N_7092,N_7626);
xnor U18511 (N_18511,N_6686,N_7832);
or U18512 (N_18512,N_11220,N_10677);
nand U18513 (N_18513,N_7175,N_11557);
nand U18514 (N_18514,N_8762,N_10587);
nor U18515 (N_18515,N_7061,N_11972);
and U18516 (N_18516,N_12269,N_8743);
nand U18517 (N_18517,N_6377,N_6819);
or U18518 (N_18518,N_11922,N_9474);
nor U18519 (N_18519,N_10327,N_8986);
xor U18520 (N_18520,N_8467,N_7256);
nor U18521 (N_18521,N_8676,N_11180);
or U18522 (N_18522,N_8232,N_8572);
and U18523 (N_18523,N_9281,N_7631);
nand U18524 (N_18524,N_6467,N_7460);
nor U18525 (N_18525,N_10140,N_7100);
or U18526 (N_18526,N_11028,N_8118);
nand U18527 (N_18527,N_7028,N_8748);
xnor U18528 (N_18528,N_9692,N_7657);
nand U18529 (N_18529,N_6518,N_11437);
xor U18530 (N_18530,N_8139,N_10816);
nor U18531 (N_18531,N_6857,N_11933);
xor U18532 (N_18532,N_8107,N_12415);
and U18533 (N_18533,N_9017,N_11909);
xnor U18534 (N_18534,N_6289,N_8963);
or U18535 (N_18535,N_11071,N_9201);
nand U18536 (N_18536,N_8440,N_9235);
nor U18537 (N_18537,N_11565,N_8845);
and U18538 (N_18538,N_7659,N_7945);
or U18539 (N_18539,N_8181,N_7699);
nand U18540 (N_18540,N_11641,N_11931);
nor U18541 (N_18541,N_10572,N_11714);
or U18542 (N_18542,N_8286,N_7048);
nand U18543 (N_18543,N_11308,N_7329);
nand U18544 (N_18544,N_8786,N_8143);
nor U18545 (N_18545,N_7707,N_8484);
xnor U18546 (N_18546,N_7565,N_12274);
and U18547 (N_18547,N_9608,N_7319);
nor U18548 (N_18548,N_8824,N_8221);
and U18549 (N_18549,N_10520,N_8230);
nor U18550 (N_18550,N_10472,N_8501);
or U18551 (N_18551,N_6760,N_11512);
or U18552 (N_18552,N_6400,N_11898);
or U18553 (N_18553,N_11365,N_9345);
and U18554 (N_18554,N_9507,N_8797);
and U18555 (N_18555,N_9061,N_11053);
and U18556 (N_18556,N_7417,N_9178);
xor U18557 (N_18557,N_10998,N_12079);
xnor U18558 (N_18558,N_8311,N_6696);
nor U18559 (N_18559,N_6891,N_11387);
xnor U18560 (N_18560,N_11852,N_7472);
nor U18561 (N_18561,N_9515,N_6551);
xnor U18562 (N_18562,N_7353,N_6924);
and U18563 (N_18563,N_6778,N_9054);
xnor U18564 (N_18564,N_7115,N_8535);
nor U18565 (N_18565,N_7692,N_7533);
xor U18566 (N_18566,N_8219,N_7905);
xor U18567 (N_18567,N_11776,N_12166);
nor U18568 (N_18568,N_11462,N_10351);
xor U18569 (N_18569,N_9948,N_9524);
or U18570 (N_18570,N_11924,N_7162);
and U18571 (N_18571,N_7245,N_11652);
and U18572 (N_18572,N_8769,N_6902);
or U18573 (N_18573,N_10722,N_6606);
nor U18574 (N_18574,N_10645,N_11549);
nor U18575 (N_18575,N_12133,N_8584);
or U18576 (N_18576,N_7049,N_12233);
and U18577 (N_18577,N_11056,N_8393);
nand U18578 (N_18578,N_9064,N_9009);
nor U18579 (N_18579,N_11863,N_8859);
or U18580 (N_18580,N_9785,N_9902);
nor U18581 (N_18581,N_12314,N_6742);
nand U18582 (N_18582,N_8595,N_6618);
nor U18583 (N_18583,N_9765,N_9004);
and U18584 (N_18584,N_7351,N_9043);
nand U18585 (N_18585,N_7319,N_9711);
xnor U18586 (N_18586,N_10937,N_9653);
or U18587 (N_18587,N_12075,N_6901);
nor U18588 (N_18588,N_12069,N_11758);
nand U18589 (N_18589,N_12199,N_8628);
or U18590 (N_18590,N_11398,N_6950);
nand U18591 (N_18591,N_12231,N_8015);
or U18592 (N_18592,N_10524,N_11290);
xor U18593 (N_18593,N_6630,N_8295);
and U18594 (N_18594,N_11967,N_6367);
or U18595 (N_18595,N_8905,N_8249);
nand U18596 (N_18596,N_9963,N_11247);
and U18597 (N_18597,N_12300,N_12140);
or U18598 (N_18598,N_11899,N_10552);
nor U18599 (N_18599,N_8665,N_8038);
or U18600 (N_18600,N_7274,N_10202);
and U18601 (N_18601,N_10300,N_12265);
and U18602 (N_18602,N_10633,N_8626);
nor U18603 (N_18603,N_10648,N_11354);
or U18604 (N_18604,N_11524,N_11303);
nor U18605 (N_18605,N_8288,N_12192);
nand U18606 (N_18606,N_12463,N_7383);
nor U18607 (N_18607,N_8411,N_6428);
xnor U18608 (N_18608,N_11290,N_12236);
and U18609 (N_18609,N_8162,N_9878);
or U18610 (N_18610,N_6477,N_10005);
or U18611 (N_18611,N_11700,N_9670);
nand U18612 (N_18612,N_9030,N_11145);
or U18613 (N_18613,N_8085,N_9369);
or U18614 (N_18614,N_11614,N_10627);
nor U18615 (N_18615,N_11910,N_6988);
nand U18616 (N_18616,N_8372,N_9263);
and U18617 (N_18617,N_8712,N_9710);
and U18618 (N_18618,N_7465,N_6825);
nand U18619 (N_18619,N_8186,N_11039);
or U18620 (N_18620,N_10001,N_10800);
nor U18621 (N_18621,N_8332,N_6710);
and U18622 (N_18622,N_9099,N_11042);
xor U18623 (N_18623,N_11268,N_12326);
nor U18624 (N_18624,N_8684,N_11158);
xor U18625 (N_18625,N_8276,N_6721);
or U18626 (N_18626,N_7596,N_12480);
nor U18627 (N_18627,N_10186,N_8056);
nor U18628 (N_18628,N_6685,N_6439);
nand U18629 (N_18629,N_8413,N_9554);
xor U18630 (N_18630,N_6416,N_12375);
or U18631 (N_18631,N_10360,N_10469);
xor U18632 (N_18632,N_9975,N_8010);
nor U18633 (N_18633,N_11604,N_11200);
nor U18634 (N_18634,N_6923,N_7223);
nor U18635 (N_18635,N_6563,N_11886);
nor U18636 (N_18636,N_12147,N_12152);
nor U18637 (N_18637,N_8247,N_11090);
xor U18638 (N_18638,N_9034,N_11867);
and U18639 (N_18639,N_10581,N_9764);
xor U18640 (N_18640,N_11149,N_12247);
nand U18641 (N_18641,N_12329,N_10021);
and U18642 (N_18642,N_7703,N_10077);
or U18643 (N_18643,N_10684,N_11526);
nor U18644 (N_18644,N_10167,N_11965);
and U18645 (N_18645,N_8803,N_6863);
or U18646 (N_18646,N_8991,N_8323);
xor U18647 (N_18647,N_7853,N_7576);
and U18648 (N_18648,N_11462,N_11001);
or U18649 (N_18649,N_10035,N_8292);
xnor U18650 (N_18650,N_12114,N_12086);
and U18651 (N_18651,N_8629,N_8077);
nor U18652 (N_18652,N_8204,N_11178);
or U18653 (N_18653,N_8821,N_9020);
and U18654 (N_18654,N_10883,N_12300);
or U18655 (N_18655,N_9983,N_8128);
nor U18656 (N_18656,N_9553,N_10459);
or U18657 (N_18657,N_12377,N_9963);
nor U18658 (N_18658,N_12081,N_8492);
nor U18659 (N_18659,N_10968,N_9255);
and U18660 (N_18660,N_10781,N_7125);
or U18661 (N_18661,N_10218,N_6604);
xor U18662 (N_18662,N_10035,N_10058);
xnor U18663 (N_18663,N_11909,N_11401);
or U18664 (N_18664,N_11153,N_10817);
xor U18665 (N_18665,N_9762,N_8954);
or U18666 (N_18666,N_11660,N_10457);
nand U18667 (N_18667,N_11637,N_7450);
nand U18668 (N_18668,N_12225,N_7812);
or U18669 (N_18669,N_11360,N_8727);
and U18670 (N_18670,N_9209,N_9156);
nor U18671 (N_18671,N_11836,N_9130);
nor U18672 (N_18672,N_8387,N_11252);
and U18673 (N_18673,N_6538,N_8878);
nand U18674 (N_18674,N_6392,N_12048);
xor U18675 (N_18675,N_9490,N_8675);
xnor U18676 (N_18676,N_7384,N_11470);
nor U18677 (N_18677,N_9588,N_11684);
or U18678 (N_18678,N_8830,N_9294);
or U18679 (N_18679,N_8620,N_10160);
nand U18680 (N_18680,N_8050,N_8134);
nor U18681 (N_18681,N_11016,N_6808);
and U18682 (N_18682,N_12477,N_10340);
nor U18683 (N_18683,N_12450,N_8876);
xor U18684 (N_18684,N_12174,N_6349);
nand U18685 (N_18685,N_10244,N_6288);
nor U18686 (N_18686,N_9603,N_11489);
xnor U18687 (N_18687,N_6322,N_10244);
xnor U18688 (N_18688,N_9445,N_10608);
nand U18689 (N_18689,N_10833,N_12222);
nand U18690 (N_18690,N_10588,N_11468);
or U18691 (N_18691,N_9510,N_7767);
and U18692 (N_18692,N_8474,N_6864);
or U18693 (N_18693,N_6497,N_11532);
nand U18694 (N_18694,N_7754,N_12183);
nand U18695 (N_18695,N_6975,N_11028);
xor U18696 (N_18696,N_7846,N_8521);
nor U18697 (N_18697,N_11538,N_9645);
nor U18698 (N_18698,N_7554,N_6515);
and U18699 (N_18699,N_8007,N_11511);
xnor U18700 (N_18700,N_11349,N_11777);
nor U18701 (N_18701,N_7281,N_6377);
xor U18702 (N_18702,N_11194,N_7155);
or U18703 (N_18703,N_6533,N_7007);
or U18704 (N_18704,N_10750,N_9657);
and U18705 (N_18705,N_11605,N_11371);
and U18706 (N_18706,N_7307,N_6451);
and U18707 (N_18707,N_8006,N_8320);
xnor U18708 (N_18708,N_9086,N_11752);
xor U18709 (N_18709,N_8136,N_10916);
and U18710 (N_18710,N_11021,N_8002);
xor U18711 (N_18711,N_12022,N_6554);
nand U18712 (N_18712,N_8077,N_6608);
or U18713 (N_18713,N_6422,N_9776);
and U18714 (N_18714,N_7042,N_7744);
and U18715 (N_18715,N_12135,N_7605);
or U18716 (N_18716,N_6972,N_9944);
xor U18717 (N_18717,N_11679,N_10062);
xnor U18718 (N_18718,N_11264,N_6829);
nand U18719 (N_18719,N_9133,N_10747);
and U18720 (N_18720,N_9454,N_9171);
or U18721 (N_18721,N_10867,N_7382);
nor U18722 (N_18722,N_11642,N_7619);
nor U18723 (N_18723,N_7965,N_7828);
and U18724 (N_18724,N_11881,N_10449);
nor U18725 (N_18725,N_6295,N_11481);
or U18726 (N_18726,N_6631,N_10423);
or U18727 (N_18727,N_11444,N_6815);
or U18728 (N_18728,N_10466,N_8877);
xor U18729 (N_18729,N_10872,N_7407);
nand U18730 (N_18730,N_8553,N_6993);
nand U18731 (N_18731,N_8094,N_12188);
and U18732 (N_18732,N_8788,N_10681);
or U18733 (N_18733,N_9988,N_8714);
nor U18734 (N_18734,N_10577,N_11398);
and U18735 (N_18735,N_6251,N_8046);
xnor U18736 (N_18736,N_8341,N_10069);
and U18737 (N_18737,N_9815,N_10743);
and U18738 (N_18738,N_12028,N_11897);
nand U18739 (N_18739,N_10571,N_11090);
nand U18740 (N_18740,N_9453,N_8525);
and U18741 (N_18741,N_8344,N_6822);
xnor U18742 (N_18742,N_8223,N_11848);
xnor U18743 (N_18743,N_11973,N_9449);
or U18744 (N_18744,N_10685,N_9608);
nand U18745 (N_18745,N_8483,N_7497);
nor U18746 (N_18746,N_9113,N_11622);
nor U18747 (N_18747,N_12083,N_6293);
or U18748 (N_18748,N_12026,N_9968);
nand U18749 (N_18749,N_9765,N_10559);
or U18750 (N_18750,N_17566,N_16122);
and U18751 (N_18751,N_17919,N_15404);
nor U18752 (N_18752,N_12930,N_12617);
nand U18753 (N_18753,N_16038,N_12910);
nand U18754 (N_18754,N_13436,N_18319);
xor U18755 (N_18755,N_15441,N_14411);
nand U18756 (N_18756,N_14425,N_15369);
or U18757 (N_18757,N_15266,N_15499);
and U18758 (N_18758,N_18190,N_14816);
nor U18759 (N_18759,N_15148,N_13810);
nand U18760 (N_18760,N_15246,N_17656);
and U18761 (N_18761,N_15541,N_14243);
nand U18762 (N_18762,N_17140,N_12662);
nor U18763 (N_18763,N_17973,N_16286);
or U18764 (N_18764,N_18539,N_17003);
nor U18765 (N_18765,N_12935,N_13169);
nor U18766 (N_18766,N_13207,N_13924);
nand U18767 (N_18767,N_16535,N_17519);
and U18768 (N_18768,N_17520,N_16448);
or U18769 (N_18769,N_17905,N_17830);
and U18770 (N_18770,N_17210,N_13718);
and U18771 (N_18771,N_13748,N_13601);
or U18772 (N_18772,N_15718,N_14636);
nor U18773 (N_18773,N_15245,N_17080);
and U18774 (N_18774,N_15019,N_14619);
nor U18775 (N_18775,N_14678,N_16229);
xnor U18776 (N_18776,N_15547,N_17365);
nand U18777 (N_18777,N_17804,N_13253);
nor U18778 (N_18778,N_17768,N_15176);
and U18779 (N_18779,N_13906,N_13671);
nor U18780 (N_18780,N_16208,N_15443);
or U18781 (N_18781,N_15039,N_13248);
or U18782 (N_18782,N_16377,N_18710);
or U18783 (N_18783,N_17009,N_18010);
nand U18784 (N_18784,N_16248,N_16846);
nand U18785 (N_18785,N_14118,N_17828);
xnor U18786 (N_18786,N_17840,N_15109);
nand U18787 (N_18787,N_12561,N_13491);
nor U18788 (N_18788,N_13649,N_13648);
and U18789 (N_18789,N_13123,N_17655);
nand U18790 (N_18790,N_15239,N_14149);
or U18791 (N_18791,N_14763,N_16776);
and U18792 (N_18792,N_13614,N_14585);
xnor U18793 (N_18793,N_15159,N_15200);
or U18794 (N_18794,N_18729,N_18631);
and U18795 (N_18795,N_12801,N_16689);
or U18796 (N_18796,N_15611,N_16268);
xor U18797 (N_18797,N_18000,N_18193);
or U18798 (N_18798,N_14008,N_16727);
nor U18799 (N_18799,N_17067,N_17879);
or U18800 (N_18800,N_16271,N_12555);
and U18801 (N_18801,N_16064,N_13930);
xor U18802 (N_18802,N_18153,N_16210);
and U18803 (N_18803,N_16033,N_13866);
nand U18804 (N_18804,N_15069,N_13558);
nand U18805 (N_18805,N_15225,N_18115);
or U18806 (N_18806,N_17562,N_14163);
or U18807 (N_18807,N_17676,N_15784);
or U18808 (N_18808,N_13826,N_12905);
xor U18809 (N_18809,N_15213,N_15324);
nor U18810 (N_18810,N_18154,N_18095);
or U18811 (N_18811,N_17025,N_15495);
nor U18812 (N_18812,N_15865,N_13816);
nand U18813 (N_18813,N_16372,N_16432);
nor U18814 (N_18814,N_14203,N_17426);
or U18815 (N_18815,N_18464,N_15994);
nand U18816 (N_18816,N_17068,N_12677);
and U18817 (N_18817,N_15998,N_12945);
nor U18818 (N_18818,N_12749,N_14230);
nand U18819 (N_18819,N_16241,N_16990);
and U18820 (N_18820,N_13499,N_13894);
and U18821 (N_18821,N_13607,N_17273);
nor U18822 (N_18822,N_13783,N_16476);
nand U18823 (N_18823,N_12894,N_14086);
or U18824 (N_18824,N_16669,N_15306);
nor U18825 (N_18825,N_17586,N_16013);
xor U18826 (N_18826,N_18648,N_18224);
and U18827 (N_18827,N_13322,N_14604);
nand U18828 (N_18828,N_13680,N_16109);
and U18829 (N_18829,N_12719,N_17991);
nand U18830 (N_18830,N_15861,N_13070);
xor U18831 (N_18831,N_13953,N_17268);
xnor U18832 (N_18832,N_14434,N_17423);
and U18833 (N_18833,N_16879,N_17002);
and U18834 (N_18834,N_14233,N_18284);
or U18835 (N_18835,N_18503,N_16808);
nor U18836 (N_18836,N_17685,N_17231);
xnor U18837 (N_18837,N_17375,N_14238);
or U18838 (N_18838,N_14896,N_16779);
and U18839 (N_18839,N_12873,N_18655);
and U18840 (N_18840,N_16339,N_17459);
and U18841 (N_18841,N_17578,N_18024);
xor U18842 (N_18842,N_13781,N_12861);
and U18843 (N_18843,N_12881,N_15501);
nor U18844 (N_18844,N_14364,N_17042);
nor U18845 (N_18845,N_14525,N_12667);
or U18846 (N_18846,N_18666,N_12536);
and U18847 (N_18847,N_17189,N_16207);
nand U18848 (N_18848,N_16747,N_14354);
and U18849 (N_18849,N_16265,N_14644);
nand U18850 (N_18850,N_16561,N_13732);
or U18851 (N_18851,N_17922,N_15626);
and U18852 (N_18852,N_13703,N_14491);
and U18853 (N_18853,N_16955,N_13747);
or U18854 (N_18854,N_13466,N_12526);
or U18855 (N_18855,N_17441,N_14812);
xnor U18856 (N_18856,N_14251,N_13398);
xnor U18857 (N_18857,N_17616,N_12712);
or U18858 (N_18858,N_17248,N_16507);
nor U18859 (N_18859,N_16550,N_17324);
nor U18860 (N_18860,N_18717,N_18704);
nand U18861 (N_18861,N_15568,N_14863);
nand U18862 (N_18862,N_14710,N_15424);
nor U18863 (N_18863,N_17601,N_14949);
nor U18864 (N_18864,N_12598,N_18350);
xnor U18865 (N_18865,N_16503,N_14642);
nor U18866 (N_18866,N_14805,N_16181);
or U18867 (N_18867,N_14563,N_18113);
or U18868 (N_18868,N_16970,N_12838);
xor U18869 (N_18869,N_16802,N_14299);
xnor U18870 (N_18870,N_15919,N_15842);
or U18871 (N_18871,N_14240,N_17865);
xor U18872 (N_18872,N_14482,N_17201);
or U18873 (N_18873,N_13009,N_15941);
nor U18874 (N_18874,N_14090,N_18070);
and U18875 (N_18875,N_12682,N_15248);
nand U18876 (N_18876,N_17075,N_14503);
nor U18877 (N_18877,N_12521,N_18584);
nor U18878 (N_18878,N_14249,N_13201);
or U18879 (N_18879,N_13175,N_14134);
nand U18880 (N_18880,N_16478,N_13298);
xnor U18881 (N_18881,N_13561,N_15112);
and U18882 (N_18882,N_13042,N_13834);
nand U18883 (N_18883,N_17502,N_17598);
nor U18884 (N_18884,N_15824,N_18199);
and U18885 (N_18885,N_12740,N_15691);
nor U18886 (N_18886,N_18291,N_15769);
xor U18887 (N_18887,N_17953,N_16831);
nor U18888 (N_18888,N_17449,N_15223);
nand U18889 (N_18889,N_16330,N_14036);
or U18890 (N_18890,N_16934,N_15577);
and U18891 (N_18891,N_15191,N_12824);
xnor U18892 (N_18892,N_17594,N_16782);
nand U18893 (N_18893,N_17928,N_14576);
or U18894 (N_18894,N_13069,N_16393);
or U18895 (N_18895,N_14392,N_12781);
xor U18896 (N_18896,N_17698,N_13758);
nor U18897 (N_18897,N_17305,N_15733);
nand U18898 (N_18898,N_13210,N_13545);
xnor U18899 (N_18899,N_13712,N_18116);
xor U18900 (N_18900,N_15182,N_16678);
xor U18901 (N_18901,N_16646,N_17439);
xnor U18902 (N_18902,N_13777,N_15338);
nor U18903 (N_18903,N_15567,N_16405);
xor U18904 (N_18904,N_15863,N_18678);
or U18905 (N_18905,N_16088,N_17710);
xor U18906 (N_18906,N_17795,N_13922);
nor U18907 (N_18907,N_17577,N_15599);
xnor U18908 (N_18908,N_15821,N_15360);
or U18909 (N_18909,N_18501,N_14511);
nor U18910 (N_18910,N_16410,N_13774);
nor U18911 (N_18911,N_13563,N_13048);
nand U18912 (N_18912,N_17455,N_16847);
xnor U18913 (N_18913,N_13590,N_16750);
nor U18914 (N_18914,N_16166,N_18743);
nor U18915 (N_18915,N_16982,N_16605);
nor U18916 (N_18916,N_13650,N_14999);
nand U18917 (N_18917,N_12643,N_13572);
and U18918 (N_18918,N_18490,N_16517);
or U18919 (N_18919,N_14773,N_18593);
and U18920 (N_18920,N_15202,N_14941);
or U18921 (N_18921,N_13245,N_12967);
nand U18922 (N_18922,N_13976,N_15509);
nor U18923 (N_18923,N_15931,N_15767);
nand U18924 (N_18924,N_16200,N_15811);
nor U18925 (N_18925,N_15737,N_14154);
and U18926 (N_18926,N_13219,N_17670);
nand U18927 (N_18927,N_15725,N_17334);
or U18928 (N_18928,N_18201,N_15988);
and U18929 (N_18929,N_17274,N_12603);
xnor U18930 (N_18930,N_14599,N_14138);
nand U18931 (N_18931,N_12618,N_15673);
xor U18932 (N_18932,N_12636,N_17505);
or U18933 (N_18933,N_13991,N_15703);
nor U18934 (N_18934,N_17348,N_14860);
and U18935 (N_18935,N_13634,N_13222);
nor U18936 (N_18936,N_13497,N_16839);
nand U18937 (N_18937,N_15634,N_14869);
xor U18938 (N_18938,N_18128,N_15234);
or U18939 (N_18939,N_16409,N_15397);
or U18940 (N_18940,N_12944,N_17155);
or U18941 (N_18941,N_15074,N_14779);
and U18942 (N_18942,N_15799,N_18042);
and U18943 (N_18943,N_18724,N_16105);
and U18944 (N_18944,N_14685,N_14332);
nor U18945 (N_18945,N_13531,N_16145);
nand U18946 (N_18946,N_16039,N_14955);
or U18947 (N_18947,N_12853,N_17366);
and U18948 (N_18948,N_12898,N_14435);
nand U18949 (N_18949,N_14419,N_13768);
nand U18950 (N_18950,N_16568,N_14423);
or U18951 (N_18951,N_17216,N_15760);
and U18952 (N_18952,N_14510,N_14232);
xor U18953 (N_18953,N_15578,N_15518);
xnor U18954 (N_18954,N_15834,N_15292);
or U18955 (N_18955,N_18719,N_17667);
xor U18956 (N_18956,N_14880,N_17633);
and U18957 (N_18957,N_16770,N_16278);
xor U18958 (N_18958,N_18004,N_13603);
nor U18959 (N_18959,N_16518,N_13710);
xnor U18960 (N_18960,N_13327,N_18058);
nand U18961 (N_18961,N_16665,N_12735);
and U18962 (N_18962,N_13237,N_16653);
and U18963 (N_18963,N_15910,N_15620);
nor U18964 (N_18964,N_17557,N_15484);
and U18965 (N_18965,N_13293,N_16856);
nor U18966 (N_18966,N_17385,N_14554);
and U18967 (N_18967,N_14104,N_14991);
or U18968 (N_18968,N_17895,N_12730);
and U18969 (N_18969,N_15043,N_17653);
xnor U18970 (N_18970,N_15692,N_15381);
and U18971 (N_18971,N_14506,N_13141);
and U18972 (N_18972,N_13181,N_16301);
xor U18973 (N_18973,N_17010,N_18516);
nand U18974 (N_18974,N_16163,N_14729);
or U18975 (N_18975,N_14975,N_17389);
nor U18976 (N_18976,N_18415,N_14798);
and U18977 (N_18977,N_12939,N_14326);
nand U18978 (N_18978,N_14033,N_13092);
xnor U18979 (N_18979,N_14460,N_16259);
or U18980 (N_18980,N_12810,N_15220);
and U18981 (N_18981,N_14566,N_14442);
and U18982 (N_18982,N_16975,N_17356);
xnor U18983 (N_18983,N_13557,N_15029);
nand U18984 (N_18984,N_18151,N_15339);
xnor U18985 (N_18985,N_17877,N_16918);
nor U18986 (N_18986,N_12543,N_18212);
or U18987 (N_18987,N_12835,N_18407);
xor U18988 (N_18988,N_18345,N_14744);
and U18989 (N_18989,N_18585,N_16801);
xnor U18990 (N_18990,N_14106,N_15340);
nand U18991 (N_18991,N_18394,N_17885);
or U18992 (N_18992,N_15370,N_17948);
xor U18993 (N_18993,N_14409,N_17647);
nand U18994 (N_18994,N_14140,N_18705);
or U18995 (N_18995,N_13011,N_16269);
or U18996 (N_18996,N_16754,N_18209);
and U18997 (N_18997,N_14914,N_14221);
nor U18998 (N_18998,N_17171,N_12866);
and U18999 (N_18999,N_17051,N_18304);
or U19000 (N_19000,N_16910,N_16713);
nor U19001 (N_19001,N_17143,N_15859);
or U19002 (N_19002,N_16637,N_18281);
and U19003 (N_19003,N_15560,N_16688);
xor U19004 (N_19004,N_13884,N_16641);
nand U19005 (N_19005,N_18688,N_15482);
and U19006 (N_19006,N_13278,N_14217);
nand U19007 (N_19007,N_15034,N_15832);
or U19008 (N_19008,N_16319,N_12863);
nor U19009 (N_19009,N_16051,N_13445);
xnor U19010 (N_19010,N_15506,N_12778);
or U19011 (N_19011,N_16686,N_13112);
and U19012 (N_19012,N_12796,N_16498);
nand U19013 (N_19013,N_15089,N_16971);
nand U19014 (N_19014,N_16866,N_17026);
nand U19015 (N_19015,N_17965,N_13525);
or U19016 (N_19016,N_17541,N_16819);
nor U19017 (N_19017,N_18351,N_18700);
nand U19018 (N_19018,N_13336,N_16472);
or U19019 (N_19019,N_14751,N_15476);
nand U19020 (N_19020,N_14595,N_17161);
nand U19021 (N_19021,N_18340,N_13211);
and U19022 (N_19022,N_14671,N_18522);
xor U19023 (N_19023,N_17821,N_18545);
nor U19024 (N_19024,N_15804,N_12761);
nand U19025 (N_19025,N_17343,N_17465);
xnor U19026 (N_19026,N_13297,N_16826);
nor U19027 (N_19027,N_16923,N_14899);
xor U19028 (N_19028,N_15709,N_16891);
xnor U19029 (N_19029,N_12868,N_14341);
xnor U19030 (N_19030,N_16935,N_18438);
and U19031 (N_19031,N_18448,N_15285);
nand U19032 (N_19032,N_17517,N_15001);
nand U19033 (N_19033,N_14723,N_16395);
and U19034 (N_19034,N_18061,N_13326);
and U19035 (N_19035,N_18337,N_13346);
nand U19036 (N_19036,N_14325,N_18441);
and U19037 (N_19037,N_18382,N_17607);
or U19038 (N_19038,N_14100,N_17311);
nor U19039 (N_19039,N_14564,N_16896);
xor U19040 (N_19040,N_14205,N_16621);
nor U19041 (N_19041,N_13138,N_17748);
and U19042 (N_19042,N_18371,N_17309);
nand U19043 (N_19043,N_16362,N_14550);
or U19044 (N_19044,N_14837,N_17336);
nand U19045 (N_19045,N_15759,N_17294);
nand U19046 (N_19046,N_17117,N_16916);
xor U19047 (N_19047,N_15907,N_18094);
nor U19048 (N_19048,N_14822,N_18478);
or U19049 (N_19049,N_15014,N_14903);
xnor U19050 (N_19050,N_13877,N_14150);
xor U19051 (N_19051,N_15674,N_15696);
nor U19052 (N_19052,N_16807,N_14388);
and U19053 (N_19053,N_15918,N_17071);
or U19054 (N_19054,N_16461,N_14547);
and U19055 (N_19055,N_15520,N_17509);
and U19056 (N_19056,N_12797,N_17634);
or U19057 (N_19057,N_13527,N_14730);
or U19058 (N_19058,N_18472,N_16315);
or U19059 (N_19059,N_13337,N_17695);
or U19060 (N_19060,N_18624,N_15473);
xnor U19061 (N_19061,N_13532,N_17875);
and U19062 (N_19062,N_15592,N_13999);
nor U19063 (N_19063,N_17668,N_16187);
nand U19064 (N_19064,N_16592,N_14324);
and U19065 (N_19065,N_13799,N_16499);
nor U19066 (N_19066,N_18426,N_16930);
nor U19067 (N_19067,N_18656,N_17611);
or U19068 (N_19068,N_16387,N_14142);
nand U19069 (N_19069,N_14818,N_17891);
and U19070 (N_19070,N_13630,N_12644);
nor U19071 (N_19071,N_12726,N_16912);
and U19072 (N_19072,N_13931,N_17024);
and U19073 (N_19073,N_17226,N_17062);
nand U19074 (N_19074,N_17107,N_15664);
nand U19075 (N_19075,N_16717,N_14709);
nand U19076 (N_19076,N_17864,N_12785);
xnor U19077 (N_19077,N_17779,N_16093);
nor U19078 (N_19078,N_14436,N_15735);
or U19079 (N_19079,N_12833,N_15395);
or U19080 (N_19080,N_16277,N_17408);
nor U19081 (N_19081,N_13895,N_15550);
nor U19082 (N_19082,N_16570,N_13909);
and U19083 (N_19083,N_13269,N_13031);
and U19084 (N_19084,N_15704,N_13421);
xnor U19085 (N_19085,N_13679,N_17976);
xor U19086 (N_19086,N_13980,N_15399);
nor U19087 (N_19087,N_17418,N_15050);
and U19088 (N_19088,N_18587,N_17416);
nand U19089 (N_19089,N_13414,N_14174);
xnor U19090 (N_19090,N_13870,N_14950);
xnor U19091 (N_19091,N_17013,N_16977);
nand U19092 (N_19092,N_15479,N_14276);
xnor U19093 (N_19093,N_13890,N_18099);
xor U19094 (N_19094,N_14697,N_17192);
nor U19095 (N_19095,N_17193,N_17632);
xnor U19096 (N_19096,N_13734,N_13394);
or U19097 (N_19097,N_14030,N_13691);
nor U19098 (N_19098,N_14126,N_13104);
and U19099 (N_19099,N_14987,N_13083);
xor U19100 (N_19100,N_17224,N_14897);
nand U19101 (N_19101,N_15556,N_14707);
xor U19102 (N_19102,N_12988,N_12586);
xnor U19103 (N_19103,N_14791,N_17850);
nand U19104 (N_19104,N_15900,N_16142);
xnor U19105 (N_19105,N_13541,N_14942);
xor U19106 (N_19106,N_14328,N_12685);
xor U19107 (N_19107,N_17745,N_15584);
nor U19108 (N_19108,N_13964,N_17512);
nor U19109 (N_19109,N_12856,N_15287);
nor U19110 (N_19110,N_18707,N_18366);
or U19111 (N_19111,N_16467,N_17243);
nand U19112 (N_19112,N_14045,N_16823);
xor U19113 (N_19113,N_13157,N_17453);
and U19114 (N_19114,N_16731,N_14193);
nor U19115 (N_19115,N_17829,N_18687);
and U19116 (N_19116,N_15321,N_13389);
and U19117 (N_19117,N_14979,N_17751);
nor U19118 (N_19118,N_18258,N_12753);
and U19119 (N_19119,N_12906,N_16441);
xnor U19120 (N_19120,N_17979,N_14873);
and U19121 (N_19121,N_13625,N_12897);
or U19122 (N_19122,N_13736,N_17338);
xnor U19123 (N_19123,N_12931,N_12874);
and U19124 (N_19124,N_12963,N_18053);
or U19125 (N_19125,N_17587,N_16594);
xor U19126 (N_19126,N_13153,N_13285);
nand U19127 (N_19127,N_16716,N_17472);
and U19128 (N_19128,N_12537,N_15921);
or U19129 (N_19129,N_16483,N_17741);
and U19130 (N_19130,N_13978,N_18264);
and U19131 (N_19131,N_15688,N_14429);
nand U19132 (N_19132,N_14750,N_17691);
xor U19133 (N_19133,N_14353,N_15978);
nor U19134 (N_19134,N_13459,N_13893);
nor U19135 (N_19135,N_13613,N_17128);
nand U19136 (N_19136,N_17733,N_13496);
or U19137 (N_19137,N_12693,N_14626);
xnor U19138 (N_19138,N_16791,N_14057);
nand U19139 (N_19139,N_16877,N_13638);
nand U19140 (N_19140,N_16470,N_17456);
nand U19141 (N_19141,N_15985,N_18012);
nand U19142 (N_19142,N_16001,N_15197);
xor U19143 (N_19143,N_17360,N_16000);
nor U19144 (N_19144,N_14405,N_12772);
and U19145 (N_19145,N_14129,N_13687);
nand U19146 (N_19146,N_14611,N_17136);
or U19147 (N_19147,N_18747,N_14139);
and U19148 (N_19148,N_16338,N_16378);
xnor U19149 (N_19149,N_15357,N_18402);
or U19150 (N_19150,N_16950,N_15425);
and U19151 (N_19151,N_16397,N_16789);
nand U19152 (N_19152,N_13849,N_16020);
nor U19153 (N_19153,N_14404,N_16575);
and U19154 (N_19154,N_14242,N_18450);
xnor U19155 (N_19155,N_17835,N_15107);
or U19156 (N_19156,N_17575,N_16160);
nand U19157 (N_19157,N_16588,N_14124);
xor U19158 (N_19158,N_14080,N_16543);
and U19159 (N_19159,N_18699,N_16421);
xor U19160 (N_19160,N_13760,N_13698);
nor U19161 (N_19161,N_16243,N_13822);
and U19162 (N_19162,N_14147,N_18542);
xnor U19163 (N_19163,N_14652,N_14358);
nor U19164 (N_19164,N_13837,N_16625);
xnor U19165 (N_19165,N_15435,N_15401);
nand U19166 (N_19166,N_18006,N_13560);
or U19167 (N_19167,N_16564,N_16041);
or U19168 (N_19168,N_13144,N_15969);
nor U19169 (N_19169,N_16164,N_17568);
nor U19170 (N_19170,N_16199,N_13514);
nand U19171 (N_19171,N_17551,N_12843);
nand U19172 (N_19172,N_16548,N_13086);
and U19173 (N_19173,N_13038,N_13988);
nor U19174 (N_19174,N_13160,N_18228);
or U19175 (N_19175,N_13908,N_14262);
nand U19176 (N_19176,N_16673,N_16071);
nand U19177 (N_19177,N_17728,N_13187);
xnor U19178 (N_19178,N_13959,N_18092);
xor U19179 (N_19179,N_16723,N_17776);
and U19180 (N_19180,N_17532,N_17582);
or U19181 (N_19181,N_17183,N_12878);
nand U19182 (N_19182,N_16018,N_15575);
nand U19183 (N_19183,N_14911,N_18100);
and U19184 (N_19184,N_15117,N_13936);
nor U19185 (N_19185,N_15031,N_12591);
or U19186 (N_19186,N_17901,N_13072);
xor U19187 (N_19187,N_12571,N_12996);
or U19188 (N_19188,N_14708,N_14451);
and U19189 (N_19189,N_16995,N_14743);
nand U19190 (N_19190,N_17629,N_15820);
or U19191 (N_19191,N_18214,N_15666);
nand U19192 (N_19192,N_12922,N_15668);
or U19193 (N_19193,N_13666,N_15152);
xor U19194 (N_19194,N_16585,N_15937);
nand U19195 (N_19195,N_17490,N_18566);
nor U19196 (N_19196,N_12793,N_13667);
or U19197 (N_19197,N_13199,N_17933);
and U19198 (N_19198,N_12524,N_15650);
xnor U19199 (N_19199,N_15408,N_16932);
nand U19200 (N_19200,N_16009,N_13244);
or U19201 (N_19201,N_15817,N_15719);
nand U19202 (N_19202,N_15440,N_17176);
and U19203 (N_19203,N_17109,N_16600);
nand U19204 (N_19204,N_16340,N_16814);
nor U19205 (N_19205,N_15894,N_17152);
nor U19206 (N_19206,N_16103,N_15235);
xnor U19207 (N_19207,N_14214,N_13343);
or U19208 (N_19208,N_12582,N_18709);
and U19209 (N_19209,N_13746,N_18018);
nand U19210 (N_19210,N_14314,N_15858);
nand U19211 (N_19211,N_14895,N_13766);
and U19212 (N_19212,N_13958,N_17537);
xnor U19213 (N_19213,N_13861,N_17618);
and U19214 (N_19214,N_18148,N_18417);
nor U19215 (N_19215,N_15742,N_12558);
or U19216 (N_19216,N_17282,N_14971);
xor U19217 (N_19217,N_12901,N_17157);
xnor U19218 (N_19218,N_17106,N_18627);
nor U19219 (N_19219,N_14518,N_15012);
nand U19220 (N_19220,N_16872,N_15571);
nand U19221 (N_19221,N_16549,N_15415);
nor U19222 (N_19222,N_17581,N_15079);
xor U19223 (N_19223,N_17208,N_16416);
or U19224 (N_19224,N_12828,N_15946);
xor U19225 (N_19225,N_14884,N_13657);
nand U19226 (N_19226,N_17605,N_18654);
xor U19227 (N_19227,N_18287,N_13681);
or U19228 (N_19228,N_18663,N_16254);
and U19229 (N_19229,N_13252,N_18181);
and U19230 (N_19230,N_16440,N_16250);
nand U19231 (N_19231,N_14938,N_13200);
xor U19232 (N_19232,N_16171,N_18505);
or U19233 (N_19233,N_14614,N_13110);
nor U19234 (N_19234,N_17099,N_12933);
or U19235 (N_19235,N_13473,N_16859);
and U19236 (N_19236,N_14716,N_15876);
nand U19237 (N_19237,N_16659,N_15980);
and U19238 (N_19238,N_16974,N_16464);
or U19239 (N_19239,N_13982,N_12530);
xor U19240 (N_19240,N_16050,N_18680);
xnor U19241 (N_19241,N_14637,N_14391);
nor U19242 (N_19242,N_18436,N_17163);
and U19243 (N_19243,N_14630,N_17495);
xnor U19244 (N_19244,N_17823,N_16374);
xor U19245 (N_19245,N_12698,N_17049);
nor U19246 (N_19246,N_13275,N_14463);
or U19247 (N_19247,N_16817,N_15629);
nand U19248 (N_19248,N_13889,N_17015);
nor U19249 (N_19249,N_18497,N_12563);
or U19250 (N_19250,N_13963,N_13790);
nor U19251 (N_19251,N_13440,N_17384);
nand U19252 (N_19252,N_16459,N_17079);
nand U19253 (N_19253,N_12849,N_14018);
xnor U19254 (N_19254,N_13063,N_17686);
nor U19255 (N_19255,N_18456,N_13972);
or U19256 (N_19256,N_15713,N_12700);
or U19257 (N_19257,N_15485,N_16897);
xnor U19258 (N_19258,N_18574,N_18137);
nor U19259 (N_19259,N_17145,N_15414);
nor U19260 (N_19260,N_16322,N_12633);
and U19261 (N_19261,N_14196,N_16155);
nor U19262 (N_19262,N_15032,N_17129);
xnor U19263 (N_19263,N_13324,N_15290);
xor U19264 (N_19264,N_15334,N_13221);
nor U19265 (N_19265,N_17569,N_14956);
xor U19266 (N_19266,N_13378,N_18052);
nand U19267 (N_19267,N_12953,N_17630);
or U19268 (N_19268,N_13279,N_14281);
nor U19269 (N_19269,N_18535,N_17564);
nand U19270 (N_19270,N_16246,N_14963);
or U19271 (N_19271,N_17848,N_17332);
and U19272 (N_19272,N_16712,N_14091);
nor U19273 (N_19273,N_16094,N_14499);
and U19274 (N_19274,N_13905,N_14162);
nor U19275 (N_19275,N_17083,N_16218);
nand U19276 (N_19276,N_18636,N_15648);
or U19277 (N_19277,N_17711,N_17046);
and U19278 (N_19278,N_16255,N_17241);
nor U19279 (N_19279,N_13356,N_13665);
xnor U19280 (N_19280,N_16956,N_12547);
or U19281 (N_19281,N_15512,N_18028);
and U19282 (N_19282,N_15371,N_13508);
nand U19283 (N_19283,N_18347,N_14504);
nand U19284 (N_19284,N_15715,N_14159);
and U19285 (N_19285,N_16446,N_14137);
xnor U19286 (N_19286,N_12973,N_12814);
nor U19287 (N_19287,N_17787,N_13587);
xor U19288 (N_19288,N_12805,N_18484);
nor U19289 (N_19289,N_18132,N_14622);
xnor U19290 (N_19290,N_17882,N_17424);
or U19291 (N_19291,N_14878,N_16080);
and U19292 (N_19292,N_16272,N_12768);
nand U19293 (N_19293,N_16466,N_14272);
or U19294 (N_19294,N_17341,N_13154);
and U19295 (N_19295,N_17287,N_14254);
nand U19296 (N_19296,N_16540,N_14133);
xnor U19297 (N_19297,N_18510,N_12597);
and U19298 (N_19298,N_17797,N_13411);
nor U19299 (N_19299,N_15645,N_15749);
or U19300 (N_19300,N_13957,N_12612);
nand U19301 (N_19301,N_15474,N_13850);
nand U19302 (N_19302,N_13548,N_13661);
or U19303 (N_19303,N_16045,N_16597);
nor U19304 (N_19304,N_13302,N_13651);
and U19305 (N_19305,N_17436,N_14165);
nand U19306 (N_19306,N_12692,N_13787);
or U19307 (N_19307,N_17286,N_14748);
nand U19308 (N_19308,N_18271,N_13984);
nand U19309 (N_19309,N_17681,N_16417);
xor U19310 (N_19310,N_16674,N_13475);
nor U19311 (N_19311,N_17744,N_18701);
xnor U19312 (N_19312,N_17386,N_14902);
or U19313 (N_19313,N_16328,N_13139);
xnor U19314 (N_19314,N_14224,N_15388);
and U19315 (N_19315,N_17089,N_18473);
or U19316 (N_19316,N_13464,N_12554);
xnor U19317 (N_19317,N_15925,N_14948);
or U19318 (N_19318,N_15956,N_13163);
xor U19319 (N_19319,N_16253,N_14122);
nand U19320 (N_19320,N_18486,N_14649);
nor U19321 (N_19321,N_17964,N_15930);
and U19322 (N_19322,N_18198,N_18698);
nor U19323 (N_19323,N_14635,N_14790);
or U19324 (N_19324,N_17806,N_14803);
and U19325 (N_19325,N_13956,N_12875);
nand U19326 (N_19326,N_15218,N_12671);
and U19327 (N_19327,N_14185,N_13920);
nor U19328 (N_19328,N_17159,N_16346);
or U19329 (N_19329,N_15544,N_16353);
and U19330 (N_19330,N_13420,N_15377);
xor U19331 (N_19331,N_16141,N_18289);
xnor U19332 (N_19332,N_15752,N_14345);
or U19333 (N_19333,N_16987,N_13494);
xnor U19334 (N_19334,N_17606,N_17281);
nor U19335 (N_19335,N_15705,N_17120);
or U19336 (N_19336,N_13299,N_17263);
or U19337 (N_19337,N_16501,N_16149);
xor U19338 (N_19338,N_18040,N_18076);
nor U19339 (N_19339,N_17956,N_14919);
and U19340 (N_19340,N_16758,N_15264);
or U19341 (N_19341,N_17934,N_12714);
nand U19342 (N_19342,N_12896,N_17648);
nand U19343 (N_19343,N_17296,N_16493);
xor U19344 (N_19344,N_13852,N_15699);
nand U19345 (N_19345,N_18540,N_13241);
nand U19346 (N_19346,N_17086,N_18568);
or U19347 (N_19347,N_15563,N_12915);
nor U19348 (N_19348,N_14810,N_13053);
nor U19349 (N_19349,N_15376,N_14390);
xnor U19350 (N_19350,N_14173,N_14918);
nand U19351 (N_19351,N_16765,N_13755);
nor U19352 (N_19352,N_12800,N_18273);
and U19353 (N_19353,N_17525,N_16902);
or U19354 (N_19354,N_14983,N_17038);
and U19355 (N_19355,N_16709,N_14146);
or U19356 (N_19356,N_16903,N_15261);
nand U19357 (N_19357,N_14540,N_15378);
or U19358 (N_19358,N_17177,N_12859);
and U19359 (N_19359,N_16870,N_12891);
nor U19360 (N_19360,N_15426,N_17029);
or U19361 (N_19361,N_14721,N_16683);
xor U19362 (N_19362,N_13595,N_17697);
nand U19363 (N_19363,N_15935,N_14155);
and U19364 (N_19364,N_15623,N_13775);
xnor U19365 (N_19365,N_15761,N_14889);
and U19366 (N_19366,N_14766,N_15896);
xor U19367 (N_19367,N_14718,N_15593);
or U19368 (N_19368,N_17218,N_17220);
xnor U19369 (N_19369,N_12903,N_15954);
xor U19370 (N_19370,N_14014,N_17799);
and U19371 (N_19371,N_16833,N_16030);
nor U19372 (N_19372,N_12770,N_16333);
or U19373 (N_19373,N_14407,N_15275);
or U19374 (N_19374,N_17205,N_16204);
and U19375 (N_19375,N_15616,N_12836);
or U19376 (N_19376,N_13090,N_17927);
or U19377 (N_19377,N_16893,N_13105);
xnor U19378 (N_19378,N_13730,N_17794);
nor U19379 (N_19379,N_15483,N_12920);
or U19380 (N_19380,N_16595,N_14973);
nor U19381 (N_19381,N_18395,N_18507);
or U19382 (N_19382,N_17331,N_13006);
and U19383 (N_19383,N_16703,N_17912);
nor U19384 (N_19384,N_15826,N_14327);
nand U19385 (N_19385,N_15707,N_15642);
xor U19386 (N_19386,N_15273,N_16004);
xnor U19387 (N_19387,N_16941,N_16394);
or U19388 (N_19388,N_14688,N_15406);
xor U19389 (N_19389,N_16952,N_14777);
or U19390 (N_19390,N_12925,N_12837);
nor U19391 (N_19391,N_13949,N_13631);
nand U19392 (N_19392,N_16002,N_15678);
xnor U19393 (N_19393,N_12995,N_16305);
xnor U19394 (N_19394,N_15746,N_12775);
xor U19395 (N_19395,N_17563,N_17346);
or U19396 (N_19396,N_14857,N_16947);
nor U19397 (N_19397,N_13762,N_12993);
nor U19398 (N_19398,N_12816,N_18459);
or U19399 (N_19399,N_14447,N_17405);
xnor U19400 (N_19400,N_16044,N_17373);
nor U19401 (N_19401,N_16586,N_16324);
xnor U19402 (N_19402,N_16144,N_13064);
xor U19403 (N_19403,N_13345,N_13693);
nand U19404 (N_19404,N_18163,N_18243);
nand U19405 (N_19405,N_18625,N_14444);
nor U19406 (N_19406,N_14362,N_13773);
nor U19407 (N_19407,N_15794,N_16424);
nand U19408 (N_19408,N_15316,N_13642);
or U19409 (N_19409,N_16792,N_16107);
xor U19410 (N_19410,N_13402,N_12754);
nand U19411 (N_19411,N_13156,N_16345);
and U19412 (N_19412,N_14613,N_15265);
or U19413 (N_19413,N_16825,N_13772);
or U19414 (N_19414,N_16373,N_13675);
or U19415 (N_19415,N_12943,N_14820);
and U19416 (N_19416,N_16168,N_17211);
or U19417 (N_19417,N_15466,N_17662);
xor U19418 (N_19418,N_16924,N_15652);
nand U19419 (N_19419,N_15885,N_16677);
nor U19420 (N_19420,N_13183,N_16282);
xor U19421 (N_19421,N_16858,N_18005);
and U19422 (N_19422,N_18396,N_14143);
xnor U19423 (N_19423,N_15839,N_13863);
xnor U19424 (N_19424,N_18159,N_17621);
xnor U19425 (N_19425,N_17983,N_14038);
and U19426 (N_19426,N_14487,N_17288);
xnor U19427 (N_19427,N_18676,N_13381);
xnor U19428 (N_19428,N_12703,N_17721);
or U19429 (N_19429,N_16165,N_14625);
xor U19430 (N_19430,N_14278,N_13249);
or U19431 (N_19431,N_13907,N_12653);
or U19432 (N_19432,N_18658,N_14998);
nand U19433 (N_19433,N_16816,N_16436);
or U19434 (N_19434,N_14359,N_13556);
xnor U19435 (N_19435,N_14592,N_16386);
xnor U19436 (N_19436,N_13050,N_17054);
or U19437 (N_19437,N_18210,N_17330);
nand U19438 (N_19438,N_17397,N_17347);
xnor U19439 (N_19439,N_15046,N_14670);
xor U19440 (N_19440,N_15132,N_17043);
xnor U19441 (N_19441,N_18420,N_12622);
or U19442 (N_19442,N_12817,N_18220);
nand U19443 (N_19443,N_15229,N_16124);
and U19444 (N_19444,N_13342,N_17937);
xnor U19445 (N_19445,N_18629,N_16577);
xnor U19446 (N_19446,N_16420,N_16146);
or U19447 (N_19447,N_13859,N_12802);
xor U19448 (N_19448,N_17715,N_16921);
nor U19449 (N_19449,N_14226,N_16314);
nand U19450 (N_19450,N_14157,N_15906);
nand U19451 (N_19451,N_15188,N_15127);
nor U19452 (N_19452,N_14831,N_12825);
xor U19453 (N_19453,N_15891,N_16607);
and U19454 (N_19454,N_15497,N_13582);
and U19455 (N_19455,N_16862,N_12907);
and U19456 (N_19456,N_16704,N_16881);
or U19457 (N_19457,N_17212,N_17101);
nand U19458 (N_19458,N_15622,N_13793);
nand U19459 (N_19459,N_14235,N_15331);
nand U19460 (N_19460,N_12979,N_14197);
nor U19461 (N_19461,N_16293,N_16120);
nand U19462 (N_19462,N_16635,N_13868);
and U19463 (N_19463,N_13047,N_14826);
and U19464 (N_19464,N_14584,N_16739);
xnor U19465 (N_19465,N_12553,N_14283);
and U19466 (N_19466,N_13130,N_18089);
and U19467 (N_19467,N_18621,N_18668);
and U19468 (N_19468,N_14158,N_15135);
and U19469 (N_19469,N_14178,N_14523);
or U19470 (N_19470,N_17207,N_13362);
and U19471 (N_19471,N_13380,N_13896);
nor U19472 (N_19472,N_13576,N_17946);
nor U19473 (N_19473,N_17476,N_12674);
nand U19474 (N_19474,N_17319,N_16837);
nand U19475 (N_19475,N_17918,N_13430);
or U19476 (N_19476,N_12917,N_15352);
nor U19477 (N_19477,N_17726,N_13258);
xnor U19478 (N_19478,N_15822,N_14212);
nor U19479 (N_19479,N_15288,N_18002);
nand U19480 (N_19480,N_13379,N_16384);
or U19481 (N_19481,N_13478,N_15807);
nand U19482 (N_19482,N_17061,N_18630);
xor U19483 (N_19483,N_14257,N_14994);
nor U19484 (N_19484,N_12535,N_18213);
nand U19485 (N_19485,N_15828,N_16062);
nor U19486 (N_19486,N_15914,N_17209);
and U19487 (N_19487,N_13733,N_15916);
and U19488 (N_19488,N_13805,N_17675);
or U19489 (N_19489,N_17672,N_18408);
and U19490 (N_19490,N_12615,N_15274);
nand U19491 (N_19491,N_18504,N_12619);
or U19492 (N_19492,N_18601,N_13434);
or U19493 (N_19493,N_16306,N_18476);
xnor U19494 (N_19494,N_13348,N_16647);
xor U19495 (N_19495,N_15566,N_17513);
nor U19496 (N_19496,N_17527,N_17497);
or U19497 (N_19497,N_15216,N_13552);
nand U19498 (N_19498,N_15534,N_13301);
nand U19499 (N_19499,N_12600,N_16634);
xnor U19500 (N_19500,N_13507,N_17955);
and U19501 (N_19501,N_15597,N_14934);
or U19502 (N_19502,N_18679,N_12929);
nand U19503 (N_19503,N_17230,N_15304);
nor U19504 (N_19504,N_14556,N_16626);
xor U19505 (N_19505,N_14567,N_15208);
and U19506 (N_19506,N_16358,N_18231);
nand U19507 (N_19507,N_14220,N_17732);
or U19508 (N_19508,N_15687,N_15282);
and U19509 (N_19509,N_16929,N_15337);
nor U19510 (N_19510,N_12803,N_15270);
nor U19511 (N_19511,N_16900,N_15180);
nand U19512 (N_19512,N_13373,N_16108);
or U19513 (N_19513,N_13966,N_13318);
xnor U19514 (N_19514,N_13272,N_14501);
xor U19515 (N_19515,N_15133,N_16718);
xor U19516 (N_19516,N_14852,N_16492);
or U19517 (N_19517,N_14285,N_15895);
nand U19518 (N_19518,N_17492,N_14148);
and U19519 (N_19519,N_15809,N_17342);
and U19520 (N_19520,N_12504,N_16256);
and U19521 (N_19521,N_15181,N_18410);
xnor U19522 (N_19522,N_13453,N_16161);
xor U19523 (N_19523,N_18423,N_15893);
or U19524 (N_19524,N_13314,N_13695);
xnor U19525 (N_19525,N_17876,N_14207);
xor U19526 (N_19526,N_14200,N_18696);
nand U19527 (N_19527,N_17935,N_18105);
nor U19528 (N_19528,N_14758,N_12938);
nor U19529 (N_19529,N_13812,N_18176);
xor U19530 (N_19530,N_15646,N_15244);
nor U19531 (N_19531,N_15528,N_14912);
and U19532 (N_19532,N_18008,N_16230);
or U19533 (N_19533,N_13469,N_16349);
xor U19534 (N_19534,N_16102,N_16662);
xnor U19535 (N_19535,N_13711,N_17508);
nand U19536 (N_19536,N_13087,N_14422);
nand U19537 (N_19537,N_13454,N_13670);
nand U19538 (N_19538,N_17197,N_13602);
and U19539 (N_19539,N_18626,N_14856);
and U19540 (N_19540,N_17333,N_17350);
and U19541 (N_19541,N_17831,N_14769);
nand U19542 (N_19542,N_15461,N_16402);
and U19543 (N_19543,N_17415,N_14535);
and U19544 (N_19544,N_15953,N_14719);
and U19545 (N_19545,N_17464,N_16313);
nand U19546 (N_19546,N_15962,N_14638);
and U19547 (N_19547,N_15536,N_13610);
or U19548 (N_19548,N_12767,N_17368);
and U19549 (N_19549,N_12911,N_17781);
or U19550 (N_19550,N_14078,N_17654);
or U19551 (N_19551,N_12738,N_14333);
or U19552 (N_19552,N_17008,N_16958);
nand U19553 (N_19553,N_17467,N_12812);
xor U19554 (N_19554,N_16931,N_17134);
or U19555 (N_19555,N_16236,N_12912);
and U19556 (N_19556,N_14530,N_17175);
nor U19557 (N_19557,N_12766,N_16389);
nor U19558 (N_19558,N_12737,N_16805);
and U19559 (N_19559,N_18563,N_18596);
or U19560 (N_19560,N_18288,N_16925);
xor U19561 (N_19561,N_16655,N_16832);
nor U19562 (N_19562,N_15394,N_13372);
or U19563 (N_19563,N_17265,N_18362);
nand U19564 (N_19564,N_14059,N_16672);
xor U19565 (N_19565,N_16106,N_18275);
nor U19566 (N_19566,N_16761,N_15755);
or U19567 (N_19567,N_12694,N_12882);
nor U19568 (N_19568,N_13814,N_13182);
xnor U19569 (N_19569,N_13442,N_18114);
and U19570 (N_19570,N_17921,N_15530);
nand U19571 (N_19571,N_15231,N_17290);
xor U19572 (N_19572,N_17339,N_12628);
xor U19573 (N_19573,N_16334,N_13231);
nand U19574 (N_19574,N_18741,N_15351);
and U19575 (N_19575,N_14483,N_17153);
or U19576 (N_19576,N_16945,N_13830);
xor U19577 (N_19577,N_13172,N_18429);
or U19578 (N_19578,N_18695,N_16428);
or U19579 (N_19579,N_18614,N_15055);
xor U19580 (N_19580,N_12876,N_15469);
nor U19581 (N_19581,N_13965,N_14075);
and U19582 (N_19582,N_15094,N_18435);
or U19583 (N_19583,N_14529,N_18653);
nand U19584 (N_19584,N_12734,N_12679);
nand U19585 (N_19585,N_13292,N_18318);
or U19586 (N_19586,N_14572,N_12921);
and U19587 (N_19587,N_15867,N_14123);
xnor U19588 (N_19588,N_14865,N_13451);
nand U19589 (N_19589,N_13408,N_14633);
or U19590 (N_19590,N_12724,N_14959);
or U19591 (N_19591,N_13490,N_15600);
and U19592 (N_19592,N_14706,N_17597);
and U19593 (N_19593,N_13981,N_15054);
nor U19594 (N_19594,N_13328,N_15753);
and U19595 (N_19595,N_15047,N_13547);
nand U19596 (N_19596,N_17514,N_15960);
xor U19597 (N_19597,N_18606,N_14534);
and U19598 (N_19598,N_15601,N_12799);
nor U19599 (N_19599,N_17412,N_15048);
xor U19600 (N_19600,N_14765,N_13288);
and U19601 (N_19601,N_12517,N_13538);
nor U19602 (N_19602,N_17402,N_13776);
nand U19603 (N_19603,N_17023,N_16220);
or U19604 (N_19604,N_14609,N_15237);
nor U19605 (N_19605,N_17432,N_14046);
or U19606 (N_19606,N_17031,N_13323);
nand U19607 (N_19607,N_15860,N_14308);
and U19608 (N_19608,N_13708,N_15902);
and U19609 (N_19609,N_17549,N_18623);
nand U19610 (N_19610,N_18694,N_18245);
nand U19611 (N_19611,N_15085,N_17404);
xnor U19612 (N_19612,N_14318,N_17814);
xnor U19613 (N_19613,N_13137,N_17609);
nand U19614 (N_19614,N_15052,N_18016);
nand U19615 (N_19615,N_13100,N_14690);
or U19616 (N_19616,N_16276,N_17734);
or U19617 (N_19617,N_16211,N_12947);
or U19618 (N_19618,N_15711,N_17716);
nor U19619 (N_19619,N_12789,N_13683);
xor U19620 (N_19620,N_13874,N_15137);
xor U19621 (N_19621,N_14290,N_14047);
nor U19622 (N_19622,N_17841,N_12968);
nor U19623 (N_19623,N_14793,N_15106);
or U19624 (N_19624,N_12720,N_16027);
and U19625 (N_19625,N_13986,N_15576);
nor U19626 (N_19626,N_12959,N_14119);
nor U19627 (N_19627,N_12762,N_14992);
or U19628 (N_19628,N_14594,N_13427);
nand U19629 (N_19629,N_16827,N_16297);
nor U19630 (N_19630,N_16668,N_14042);
nand U19631 (N_19631,N_17862,N_16006);
xnor U19632 (N_19632,N_13745,N_13417);
and U19633 (N_19633,N_18236,N_15952);
or U19634 (N_19634,N_15016,N_14172);
nand U19635 (N_19635,N_18328,N_14795);
and U19636 (N_19636,N_12977,N_16292);
nor U19637 (N_19637,N_13195,N_12572);
or U19638 (N_19638,N_12872,N_13317);
xnor U19639 (N_19639,N_18553,N_13753);
nand U19640 (N_19640,N_18141,N_17815);
and U19641 (N_19641,N_15697,N_12739);
nand U19642 (N_19642,N_16407,N_16580);
and U19643 (N_19643,N_13127,N_16104);
and U19644 (N_19644,N_13888,N_13605);
nor U19645 (N_19645,N_18586,N_15833);
nand U19646 (N_19646,N_13054,N_18254);
nor U19647 (N_19647,N_15336,N_17301);
nand U19648 (N_19648,N_14647,N_16512);
nor U19649 (N_19649,N_14457,N_13264);
nor U19650 (N_19650,N_15307,N_14930);
or U19651 (N_19651,N_13366,N_14120);
xor U19652 (N_19652,N_14578,N_13045);
nor U19653 (N_19653,N_15736,N_17714);
and U19654 (N_19654,N_18262,N_15359);
nor U19655 (N_19655,N_16569,N_14229);
xor U19656 (N_19656,N_12658,N_17240);
nor U19657 (N_19657,N_17552,N_15877);
and U19658 (N_19658,N_18453,N_17838);
nand U19659 (N_19659,N_14520,N_17421);
xnor U19660 (N_19660,N_17369,N_14746);
or U19661 (N_19661,N_13283,N_14548);
nand U19662 (N_19662,N_15432,N_16615);
or U19663 (N_19663,N_13640,N_14297);
and U19664 (N_19664,N_12638,N_17910);
nand U19665 (N_19665,N_14519,N_13276);
and U19666 (N_19666,N_18577,N_12567);
xnor U19667 (N_19667,N_16465,N_15856);
xnor U19668 (N_19668,N_13882,N_16434);
and U19669 (N_19669,N_12528,N_15615);
xor U19670 (N_19670,N_16291,N_16460);
xor U19671 (N_19671,N_14844,N_15384);
nor U19672 (N_19672,N_15036,N_15975);
nand U19673 (N_19673,N_16491,N_16012);
and U19674 (N_19674,N_14432,N_13842);
xor U19675 (N_19675,N_15638,N_14677);
or U19676 (N_19676,N_13242,N_12702);
or U19677 (N_19677,N_12952,N_18363);
xor U19678 (N_19678,N_15177,N_15810);
xor U19679 (N_19679,N_13516,N_15214);
and U19680 (N_19680,N_13886,N_15454);
xnor U19681 (N_19681,N_15587,N_15573);
nor U19682 (N_19682,N_14368,N_13618);
or U19683 (N_19683,N_13194,N_15553);
nand U19684 (N_19684,N_15452,N_12549);
and U19685 (N_19685,N_13586,N_15478);
and U19686 (N_19686,N_17798,N_14702);
nor U19687 (N_19687,N_15347,N_16121);
or U19688 (N_19688,N_14093,N_14687);
nor U19689 (N_19689,N_17027,N_15457);
and U19690 (N_19690,N_13566,N_12981);
or U19691 (N_19691,N_17297,N_15904);
and U19692 (N_19692,N_16751,N_15092);
and U19693 (N_19693,N_15765,N_14258);
and U19694 (N_19694,N_12642,N_14069);
or U19695 (N_19695,N_18567,N_13113);
nand U19696 (N_19696,N_15149,N_17753);
or U19697 (N_19697,N_16959,N_13570);
nand U19698 (N_19698,N_18014,N_17030);
or U19699 (N_19699,N_16016,N_13744);
and U19700 (N_19700,N_15490,N_15350);
and U19701 (N_19701,N_18267,N_13939);
nand U19702 (N_19702,N_13872,N_14680);
xnor U19703 (N_19703,N_17604,N_18182);
xnor U19704 (N_19704,N_14537,N_15004);
nand U19705 (N_19705,N_18292,N_15038);
and U19706 (N_19706,N_14533,N_13161);
nor U19707 (N_19707,N_17847,N_16993);
nand U19708 (N_19708,N_12501,N_17925);
and U19709 (N_19709,N_14542,N_15346);
or U19710 (N_19710,N_15621,N_17306);
or U19711 (N_19711,N_14367,N_12691);
nor U19712 (N_19712,N_15653,N_18608);
or U19713 (N_19713,N_13095,N_17314);
nor U19714 (N_19714,N_14201,N_16984);
and U19715 (N_19715,N_16909,N_13528);
nor U19716 (N_19716,N_16771,N_16183);
nor U19717 (N_19717,N_16661,N_14374);
and U19718 (N_19718,N_16486,N_14679);
and U19719 (N_19719,N_17022,N_14408);
xnor U19720 (N_19720,N_17574,N_16863);
xor U19721 (N_19721,N_15186,N_15450);
nor U19722 (N_19722,N_18276,N_14321);
nor U19723 (N_19723,N_18147,N_18573);
or U19724 (N_19724,N_15557,N_15153);
and U19725 (N_19725,N_15932,N_18515);
or U19726 (N_19726,N_16755,N_15714);
xor U19727 (N_19727,N_12519,N_14464);
or U19728 (N_19728,N_15948,N_15301);
or U19729 (N_19729,N_18649,N_17693);
xnor U19730 (N_19730,N_15968,N_15184);
xnor U19731 (N_19731,N_15236,N_16201);
xnor U19732 (N_19732,N_14960,N_16400);
and U19733 (N_19733,N_17981,N_16612);
xnor U19734 (N_19734,N_17321,N_17447);
nor U19735 (N_19735,N_15105,N_15104);
nor U19736 (N_19736,N_14772,N_18009);
or U19737 (N_19737,N_17275,N_13875);
xnor U19738 (N_19738,N_17626,N_13358);
or U19739 (N_19739,N_15446,N_12786);
nand U19740 (N_19740,N_15516,N_14521);
nand U19741 (N_19741,N_15455,N_12681);
or U19742 (N_19742,N_14128,N_12661);
xor U19743 (N_19743,N_13904,N_16777);
nor U19744 (N_19744,N_15850,N_16922);
or U19745 (N_19745,N_17765,N_13854);
xnor U19746 (N_19746,N_14947,N_14917);
xnor U19747 (N_19747,N_18123,N_16509);
xor U19748 (N_19748,N_15777,N_14005);
xor U19749 (N_19749,N_13498,N_15183);
nand U19750 (N_19750,N_18015,N_15951);
nor U19751 (N_19751,N_18111,N_16042);
or U19752 (N_19752,N_14565,N_17954);
nand U19753 (N_19753,N_15958,N_12900);
xnor U19754 (N_19754,N_16125,N_18702);
nor U19755 (N_19755,N_13375,N_17649);
nor U19756 (N_19756,N_17554,N_12832);
nand U19757 (N_19757,N_17199,N_13520);
or U19758 (N_19758,N_17929,N_13057);
xor U19759 (N_19759,N_15430,N_13715);
and U19760 (N_19760,N_15419,N_15591);
nand U19761 (N_19761,N_14579,N_18582);
or U19762 (N_19762,N_16237,N_12969);
xor U19763 (N_19763,N_16772,N_12989);
nand U19764 (N_19764,N_15976,N_14377);
and U19765 (N_19765,N_17496,N_13425);
nand U19766 (N_19766,N_13947,N_13205);
nand U19767 (N_19767,N_18558,N_13639);
or U19768 (N_19768,N_15217,N_18298);
xor U19769 (N_19769,N_14828,N_12635);
and U19770 (N_19770,N_14549,N_17820);
xnor U19771 (N_19771,N_13795,N_15487);
nor U19772 (N_19772,N_14761,N_15021);
nand U19773 (N_19773,N_13079,N_12926);
nor U19774 (N_19774,N_13992,N_15525);
and U19775 (N_19775,N_15993,N_16079);
and U19776 (N_19776,N_15402,N_14039);
xor U19777 (N_19777,N_17754,N_15481);
nand U19778 (N_19778,N_16043,N_16954);
or U19779 (N_19779,N_18736,N_15924);
and U19780 (N_19780,N_14373,N_17018);
or U19781 (N_19781,N_17942,N_15837);
nand U19782 (N_19782,N_14672,N_16380);
and U19783 (N_19783,N_18165,N_16495);
and U19784 (N_19784,N_18177,N_15561);
and U19785 (N_19785,N_14337,N_17978);
nor U19786 (N_19786,N_18690,N_12718);
nor U19787 (N_19787,N_17589,N_13209);
xor U19788 (N_19788,N_14344,N_13612);
nor U19789 (N_19789,N_16767,N_13014);
nand U19790 (N_19790,N_14349,N_16186);
xor U19791 (N_19791,N_18066,N_17545);
and U19792 (N_19792,N_17899,N_16762);
nand U19793 (N_19793,N_15996,N_14551);
xnor U19794 (N_19794,N_15639,N_16841);
or U19795 (N_19795,N_14271,N_15257);
xnor U19796 (N_19796,N_17791,N_16601);
nand U19797 (N_19797,N_15818,N_18072);
and U19798 (N_19798,N_13019,N_18470);
and U19799 (N_19799,N_18122,N_14894);
nor U19800 (N_19800,N_14062,N_17470);
xor U19801 (N_19801,N_15174,N_15433);
xnor U19802 (N_19802,N_16724,N_12531);
xor U19803 (N_19803,N_17775,N_16917);
xnor U19804 (N_19804,N_18216,N_17091);
nor U19805 (N_19805,N_14190,N_17151);
nand U19806 (N_19806,N_14294,N_15788);
xor U19807 (N_19807,N_12566,N_17730);
or U19808 (N_19808,N_16235,N_17718);
nand U19809 (N_19809,N_14342,N_17064);
and U19810 (N_19810,N_14302,N_14049);
nor U19811 (N_19811,N_16262,N_13915);
or U19812 (N_19812,N_14010,N_18025);
or U19813 (N_19813,N_16511,N_15963);
nand U19814 (N_19814,N_18411,N_18021);
and U19815 (N_19815,N_14870,N_13165);
or U19816 (N_19816,N_18591,N_13023);
or U19817 (N_19817,N_15727,N_18667);
nand U19818 (N_19818,N_17962,N_13626);
xor U19819 (N_19819,N_16005,N_15332);
or U19820 (N_19820,N_17289,N_18133);
and U19821 (N_19821,N_12713,N_16602);
nand U19822 (N_19822,N_13012,N_13722);
and U19823 (N_19823,N_14872,N_18344);
or U19824 (N_19824,N_15100,N_15468);
nand U19825 (N_19825,N_16290,N_13066);
or U19826 (N_19826,N_18054,N_15572);
xnor U19827 (N_19827,N_16737,N_17692);
or U19828 (N_19828,N_17700,N_18738);
xor U19829 (N_19829,N_14117,N_17788);
or U19830 (N_19830,N_17039,N_16126);
nand U19831 (N_19831,N_13851,N_17530);
xor U19832 (N_19832,N_17112,N_14784);
nor U19833 (N_19833,N_18665,N_16736);
nor U19834 (N_19834,N_18514,N_15141);
or U19835 (N_19835,N_15607,N_14101);
nand U19836 (N_19836,N_17312,N_18599);
nand U19837 (N_19837,N_18433,N_12630);
nand U19838 (N_19838,N_15493,N_13941);
or U19839 (N_19839,N_12821,N_13131);
xnor U19840 (N_19840,N_16766,N_16835);
nor U19841 (N_19841,N_16335,N_18145);
or U19842 (N_19842,N_15315,N_15238);
nand U19843 (N_19843,N_17790,N_15500);
or U19844 (N_19844,N_14040,N_14573);
or U19845 (N_19845,N_14239,N_15302);
nor U19846 (N_19846,N_14631,N_13786);
and U19847 (N_19847,N_17673,N_14713);
nor U19848 (N_19848,N_12711,N_14854);
nor U19849 (N_19849,N_16017,N_12654);
nand U19850 (N_19850,N_14569,N_15665);
nand U19851 (N_19851,N_17097,N_12791);
or U19852 (N_19852,N_14259,N_16231);
and U19853 (N_19853,N_12680,N_16488);
xor U19854 (N_19854,N_12834,N_13974);
nand U19855 (N_19855,N_15739,N_18170);
xnor U19856 (N_19856,N_15920,N_16957);
and U19857 (N_19857,N_17326,N_16830);
nor U19858 (N_19858,N_16184,N_16266);
and U19859 (N_19859,N_14066,N_13405);
nand U19860 (N_19860,N_13869,N_13644);
xor U19861 (N_19861,N_12746,N_16245);
xor U19862 (N_19862,N_15310,N_18728);
xor U19863 (N_19863,N_18342,N_18247);
and U19864 (N_19864,N_16616,N_17202);
or U19865 (N_19865,N_15027,N_12794);
or U19866 (N_19866,N_12721,N_16973);
nor U19867 (N_19867,N_15716,N_18528);
xnor U19868 (N_19868,N_14598,N_13797);
and U19869 (N_19869,N_17826,N_12990);
or U19870 (N_19870,N_17204,N_18520);
xnor U19871 (N_19871,N_16515,N_15087);
and U19872 (N_19872,N_16799,N_12913);
xnor U19873 (N_19873,N_14800,N_17736);
nand U19874 (N_19874,N_14180,N_14832);
nand U19875 (N_19875,N_17627,N_16011);
and U19876 (N_19876,N_13985,N_16860);
xor U19877 (N_19877,N_13103,N_12858);
nor U19878 (N_19878,N_12557,N_12971);
xor U19879 (N_19879,N_17378,N_16438);
and U19880 (N_19880,N_17471,N_17987);
nand U19881 (N_19881,N_14990,N_15552);
and U19882 (N_19882,N_14393,N_16252);
and U19883 (N_19883,N_18479,N_18090);
xnor U19884 (N_19884,N_13443,N_16620);
or U19885 (N_19885,N_18266,N_15706);
and U19886 (N_19886,N_16978,N_16562);
xnor U19887 (N_19887,N_15464,N_13764);
or U19888 (N_19888,N_15740,N_16216);
nor U19889 (N_19889,N_13973,N_14989);
nor U19890 (N_19890,N_14485,N_13653);
nand U19891 (N_19891,N_18299,N_16342);
nand U19892 (N_19892,N_16157,N_16178);
nand U19893 (N_19893,N_16453,N_16323);
xor U19894 (N_19894,N_17028,N_12846);
and U19895 (N_19895,N_18499,N_16652);
xor U19896 (N_19896,N_16388,N_18353);
xor U19897 (N_19897,N_13228,N_14583);
or U19898 (N_19898,N_13617,N_12884);
xnor U19899 (N_19899,N_13627,N_15915);
nor U19900 (N_19900,N_16173,N_17995);
nand U19901 (N_19901,N_14851,N_18246);
or U19902 (N_19902,N_16508,N_17315);
or U19903 (N_19903,N_16190,N_16536);
and U19904 (N_19904,N_18491,N_12675);
xnor U19905 (N_19905,N_13455,N_15846);
and U19906 (N_19906,N_17165,N_15748);
nor U19907 (N_19907,N_18638,N_15654);
xnor U19908 (N_19908,N_14156,N_14277);
and U19909 (N_19909,N_15355,N_17102);
and U19910 (N_19910,N_17507,N_14043);
and U19911 (N_19911,N_17390,N_13967);
nor U19912 (N_19912,N_16551,N_18118);
nor U19913 (N_19913,N_15456,N_13780);
xnor U19914 (N_19914,N_18715,N_16908);
and U19915 (N_19915,N_16261,N_18269);
nor U19916 (N_19916,N_14413,N_17249);
and U19917 (N_19917,N_14406,N_18037);
nor U19918 (N_19918,N_15142,N_13771);
xor U19919 (N_19919,N_16599,N_13948);
nand U19920 (N_19920,N_14829,N_16247);
and U19921 (N_19921,N_18418,N_18488);
and U19922 (N_19922,N_14898,N_18650);
or U19923 (N_19923,N_12909,N_18681);
nor U19924 (N_19924,N_16205,N_13136);
nand U19925 (N_19925,N_15379,N_14350);
nor U19926 (N_19926,N_16224,N_13429);
nand U19927 (N_19927,N_17643,N_18238);
nand U19928 (N_19928,N_16084,N_14717);
nand U19929 (N_19929,N_17072,N_15942);
xor U19930 (N_19930,N_15647,N_14188);
or U19931 (N_19931,N_14026,N_14753);
xor U19932 (N_19932,N_12560,N_18445);
nor U19933 (N_19933,N_18661,N_16650);
and U19934 (N_19934,N_18487,N_18483);
or U19935 (N_19935,N_15944,N_16888);
nor U19936 (N_19936,N_15698,N_18730);
nand U19937 (N_19937,N_17904,N_14821);
or U19938 (N_19938,N_15318,N_14152);
or U19939 (N_19939,N_15222,N_13655);
or U19940 (N_19940,N_16883,N_14313);
or U19941 (N_19941,N_18384,N_13910);
and U19942 (N_19942,N_14234,N_18671);
nor U19943 (N_19943,N_16354,N_14489);
and U19944 (N_19944,N_15965,N_12733);
xnor U19945 (N_19945,N_15294,N_13969);
or U19946 (N_19946,N_13114,N_16026);
nor U19947 (N_19947,N_12889,N_16836);
xor U19948 (N_19948,N_17100,N_17221);
and U19949 (N_19949,N_15502,N_15296);
xnor U19950 (N_19950,N_15901,N_17110);
nor U19951 (N_19951,N_13522,N_15289);
nor U19952 (N_19952,N_18307,N_12806);
xnor U19953 (N_19953,N_18257,N_15844);
nand U19954 (N_19954,N_14684,N_15504);
and U19955 (N_19955,N_13065,N_16695);
nor U19956 (N_19956,N_17917,N_18098);
or U19957 (N_19957,N_13565,N_14365);
nor U19958 (N_19958,N_13034,N_12741);
and U19959 (N_19959,N_12723,N_18091);
nand U19960 (N_19960,N_18521,N_17533);
nor U19961 (N_19961,N_12788,N_12736);
nor U19962 (N_19962,N_13725,N_17548);
and U19963 (N_19963,N_17986,N_18179);
xnor U19964 (N_19964,N_14945,N_15470);
or U19965 (N_19965,N_14570,N_13233);
xor U19966 (N_19966,N_14824,N_15796);
nor U19967 (N_19967,N_13433,N_14977);
xor U19968 (N_19968,N_15606,N_14023);
nand U19969 (N_19969,N_15326,N_18640);
or U19970 (N_19970,N_16325,N_15588);
nand U19971 (N_19971,N_13214,N_17303);
xor U19972 (N_19972,N_16496,N_13598);
nor U19973 (N_19973,N_14053,N_13919);
nand U19974 (N_19974,N_13267,N_14470);
nor U19975 (N_19975,N_18047,N_16469);
nand U19976 (N_19976,N_17251,N_13641);
or U19977 (N_19977,N_13347,N_18711);
nand U19978 (N_19978,N_17154,N_15201);
or U19979 (N_19979,N_17801,N_16985);
nor U19980 (N_19980,N_14524,N_16528);
and U19981 (N_19981,N_14640,N_15328);
xor U19982 (N_19982,N_16757,N_18530);
xor U19983 (N_19983,N_16719,N_17669);
nand U19984 (N_19984,N_14974,N_15409);
or U19985 (N_19985,N_16060,N_13284);
and U19986 (N_19986,N_16656,N_13311);
nand U19987 (N_19987,N_16895,N_13813);
and U19988 (N_19988,N_15543,N_14752);
and U19989 (N_19989,N_14166,N_14738);
or U19990 (N_19990,N_17712,N_18431);
nor U19991 (N_19991,N_15685,N_18048);
and U19992 (N_19992,N_12577,N_15178);
nand U19993 (N_19993,N_18001,N_16228);
nand U19994 (N_19994,N_16948,N_16019);
nand U19995 (N_19995,N_15071,N_17355);
and U19996 (N_19996,N_12976,N_17073);
or U19997 (N_19997,N_17264,N_17256);
nand U19998 (N_19998,N_14228,N_16632);
nor U19999 (N_19999,N_14130,N_13960);
xor U20000 (N_20000,N_17680,N_15080);
nand U20001 (N_20001,N_13990,N_17438);
nand U20002 (N_20002,N_12500,N_14446);
and U20003 (N_20003,N_14002,N_14092);
nor U20004 (N_20004,N_16015,N_18131);
nand U20005 (N_20005,N_13833,N_17560);
or U20006 (N_20006,N_17283,N_13484);
and U20007 (N_20007,N_14867,N_12763);
nor U20008 (N_20008,N_16273,N_14722);
or U20009 (N_20009,N_13802,N_14762);
or U20010 (N_20010,N_12759,N_18404);
nand U20011 (N_20011,N_18444,N_12565);
nand U20012 (N_20012,N_17699,N_17635);
or U20013 (N_20013,N_12855,N_18635);
xnor U20014 (N_20014,N_17460,N_13867);
xor U20015 (N_20015,N_16418,N_12624);
xnor U20016 (N_20016,N_18117,N_12776);
xnor U20017 (N_20017,N_18713,N_13129);
nor U20018 (N_20018,N_13526,N_18127);
xnor U20019 (N_20019,N_17878,N_16047);
xor U20020 (N_20020,N_13251,N_15134);
nor U20021 (N_20021,N_18357,N_12928);
and U20022 (N_20022,N_13186,N_13259);
or U20023 (N_20023,N_14877,N_14891);
xor U20024 (N_20024,N_13594,N_14256);
nor U20025 (N_20025,N_15816,N_13032);
and U20026 (N_20026,N_17292,N_15108);
nand U20027 (N_20027,N_12960,N_16901);
or U20028 (N_20028,N_15010,N_16593);
nor U20029 (N_20029,N_13955,N_15847);
nand U20030 (N_20030,N_16367,N_18428);
nor U20031 (N_20031,N_17816,N_16618);
nand U20032 (N_20032,N_17353,N_13391);
or U20033 (N_20033,N_13546,N_14369);
and U20034 (N_20034,N_16850,N_17825);
or U20035 (N_20035,N_17285,N_17727);
or U20036 (N_20036,N_14607,N_18422);
nor U20037 (N_20037,N_17679,N_15670);
nand U20038 (N_20038,N_17284,N_15800);
nand U20039 (N_20039,N_13944,N_12659);
xnor U20040 (N_20040,N_18527,N_16760);
or U20041 (N_20041,N_13458,N_16177);
and U20042 (N_20042,N_16521,N_12637);
and U20043 (N_20043,N_15407,N_13133);
and U20044 (N_20044,N_17752,N_14808);
and U20045 (N_20045,N_15732,N_13470);
or U20046 (N_20046,N_15734,N_18235);
or U20047 (N_20047,N_14691,N_17478);
nor U20048 (N_20048,N_13825,N_17593);
nor U20049 (N_20049,N_16660,N_15836);
xor U20050 (N_20050,N_13240,N_13363);
or U20051 (N_20051,N_12522,N_15277);
or U20052 (N_20052,N_16573,N_13663);
xor U20053 (N_20053,N_16357,N_13353);
nor U20054 (N_20054,N_17186,N_15185);
xor U20055 (N_20055,N_14336,N_17094);
or U20056 (N_20056,N_15701,N_16824);
xnor U20057 (N_20057,N_15115,N_17920);
and U20058 (N_20058,N_16851,N_13798);
nor U20059 (N_20059,N_16443,N_15617);
xnor U20060 (N_20060,N_15772,N_12829);
or U20061 (N_20061,N_17567,N_14629);
xnor U20062 (N_20062,N_15312,N_14015);
nand U20063 (N_20063,N_15671,N_16442);
and U20064 (N_20064,N_18498,N_17837);
nor U20065 (N_20065,N_16951,N_15814);
or U20066 (N_20066,N_14456,N_13060);
nand U20067 (N_20067,N_17214,N_12962);
and U20068 (N_20068,N_13820,N_14643);
and U20069 (N_20069,N_14673,N_16869);
nand U20070 (N_20070,N_13592,N_17345);
and U20071 (N_20071,N_13268,N_16559);
or U20072 (N_20072,N_12757,N_18642);
and U20073 (N_20073,N_13481,N_15984);
and U20074 (N_20074,N_17394,N_12809);
nor U20075 (N_20075,N_17770,N_16820);
nand U20076 (N_20076,N_18581,N_17547);
or U20077 (N_20077,N_17191,N_14927);
xnor U20078 (N_20078,N_14861,N_18164);
xnor U20079 (N_20079,N_18377,N_15632);
or U20080 (N_20080,N_13335,N_17111);
nand U20081 (N_20081,N_15416,N_13678);
nor U20082 (N_20082,N_14850,N_15000);
or U20083 (N_20083,N_16936,N_18330);
xor U20084 (N_20084,N_17255,N_13349);
or U20085 (N_20085,N_16096,N_18628);
or U20086 (N_20086,N_17487,N_17361);
nand U20087 (N_20087,N_13519,N_16609);
nor U20088 (N_20088,N_17335,N_17579);
xnor U20089 (N_20089,N_17322,N_13227);
and U20090 (N_20090,N_17158,N_18306);
xnor U20091 (N_20091,N_12961,N_16745);
and U20092 (N_20092,N_17855,N_17498);
nor U20093 (N_20093,N_16711,N_13913);
nand U20094 (N_20094,N_15779,N_17146);
nand U20095 (N_20095,N_14836,N_13933);
or U20096 (N_20096,N_17223,N_13390);
xnor U20097 (N_20097,N_13446,N_16623);
nand U20098 (N_20098,N_16099,N_16730);
nand U20099 (N_20099,N_14734,N_15730);
and U20100 (N_20100,N_17475,N_16298);
nor U20101 (N_20101,N_13235,N_16590);
and U20102 (N_20102,N_16034,N_13355);
or U20103 (N_20103,N_15065,N_15187);
nor U20104 (N_20104,N_17377,N_13699);
nor U20105 (N_20105,N_18686,N_15922);
nor U20106 (N_20106,N_16963,N_14031);
nand U20107 (N_20107,N_15787,N_17069);
xnor U20108 (N_20108,N_18481,N_13512);
xor U20109 (N_20109,N_15110,N_12954);
xnor U20110 (N_20110,N_14651,N_14459);
and U20111 (N_20111,N_17376,N_18191);
nand U20112 (N_20112,N_17474,N_18294);
xnor U20113 (N_20113,N_17689,N_16986);
or U20114 (N_20114,N_15936,N_18538);
nand U20115 (N_20115,N_14135,N_16768);
and U20116 (N_20116,N_15524,N_14590);
or U20117 (N_20117,N_12895,N_14376);
nor U20118 (N_20118,N_13903,N_13185);
nor U20119 (N_20119,N_12562,N_15196);
and U20120 (N_20120,N_17190,N_13855);
and U20121 (N_20121,N_18218,N_18322);
and U20122 (N_20122,N_17115,N_14694);
nand U20123 (N_20123,N_15785,N_18250);
nor U20124 (N_20124,N_17694,N_14712);
and U20125 (N_20125,N_16326,N_14111);
nor U20126 (N_20126,N_16871,N_17299);
and U20127 (N_20127,N_13515,N_14029);
nand U20128 (N_20128,N_15120,N_18068);
and U20129 (N_20129,N_17259,N_17150);
nor U20130 (N_20130,N_12986,N_15840);
xnor U20131 (N_20131,N_18607,N_13503);
or U20132 (N_20132,N_12845,N_12783);
and U20133 (N_20133,N_18745,N_17890);
or U20134 (N_20134,N_14571,N_17381);
xor U20135 (N_20135,N_18617,N_12690);
xor U20136 (N_20136,N_18589,N_13584);
and U20137 (N_20137,N_18576,N_13168);
nand U20138 (N_20138,N_16232,N_13261);
xor U20139 (N_20139,N_12538,N_18129);
or U20140 (N_20140,N_13571,N_13001);
nand U20141 (N_20141,N_16821,N_18496);
xor U20142 (N_20142,N_16783,N_15655);
nor U20143 (N_20143,N_15156,N_17494);
and U20144 (N_20144,N_14164,N_14351);
or U20145 (N_20145,N_16556,N_12606);
xnor U20146 (N_20146,N_14381,N_18664);
nor U20147 (N_20147,N_18720,N_14965);
nand U20148 (N_20148,N_16321,N_16558);
or U20149 (N_20149,N_13435,N_13010);
or U20150 (N_20150,N_13562,N_14811);
nand U20151 (N_20151,N_13055,N_13357);
and U20152 (N_20152,N_15199,N_14866);
or U20153 (N_20153,N_18167,N_18460);
xnor U20154 (N_20154,N_12992,N_13128);
nor U20155 (N_20155,N_14764,N_12715);
nor U20156 (N_20156,N_15308,N_16545);
nand U20157 (N_20157,N_13339,N_16502);
and U20158 (N_20158,N_17127,N_13583);
and U20159 (N_20159,N_13099,N_16542);
nor U20160 (N_20160,N_16705,N_14532);
or U20161 (N_20161,N_17050,N_17631);
or U20162 (N_20162,N_17466,N_18219);
nand U20163 (N_20163,N_13533,N_17419);
nand U20164 (N_20164,N_13438,N_16749);
and U20165 (N_20165,N_16366,N_16969);
xnor U20166 (N_20166,N_14621,N_14835);
and U20167 (N_20167,N_16722,N_14961);
nor U20168 (N_20168,N_13763,N_15298);
xnor U20169 (N_20169,N_15375,N_17526);
and U20170 (N_20170,N_14496,N_17884);
xor U20171 (N_20171,N_15170,N_14946);
nor U20172 (N_20172,N_14624,N_16967);
nand U20173 (N_20173,N_17595,N_18677);
nand U20174 (N_20174,N_18139,N_14304);
nor U20175 (N_20175,N_13174,N_15793);
or U20176 (N_20176,N_16855,N_17489);
or U20177 (N_20177,N_13171,N_17388);
or U20178 (N_20178,N_15605,N_17235);
or U20179 (N_20179,N_12955,N_14731);
nor U20180 (N_20180,N_18253,N_17674);
and U20181 (N_20181,N_15558,N_12941);
or U20182 (N_20182,N_13581,N_15667);
nor U20183 (N_20183,N_14908,N_13476);
nor U20184 (N_20184,N_18083,N_13310);
nand U20185 (N_20185,N_12857,N_16195);
xnor U20186 (N_20186,N_13996,N_13509);
xor U20187 (N_20187,N_13815,N_13262);
nand U20188 (N_20188,N_16746,N_12601);
or U20189 (N_20189,N_17229,N_13836);
xor U20190 (N_20190,N_13002,N_14653);
or U20191 (N_20191,N_12583,N_15694);
and U20192 (N_20192,N_17066,N_15053);
nor U20193 (N_20193,N_16920,N_12985);
nor U20194 (N_20194,N_14806,N_17852);
xor U20195 (N_20195,N_14817,N_14454);
nor U20196 (N_20196,N_17625,N_18383);
and U20197 (N_20197,N_17778,N_17357);
and U20198 (N_20198,N_18364,N_14352);
and U20199 (N_20199,N_13794,N_16066);
xor U20200 (N_20200,N_12623,N_18124);
xor U20201 (N_20201,N_15507,N_16078);
nand U20202 (N_20202,N_17081,N_14855);
xnor U20203 (N_20203,N_13589,N_17636);
nand U20204 (N_20204,N_15929,N_15866);
nor U20205 (N_20205,N_18546,N_14319);
nor U20206 (N_20206,N_12807,N_15438);
nor U20207 (N_20207,N_12936,N_13274);
xor U20208 (N_20208,N_17731,N_14703);
xor U20209 (N_20209,N_17769,N_17510);
xnor U20210 (N_20210,N_12854,N_17713);
nand U20211 (N_20211,N_15630,N_17903);
nand U20212 (N_20212,N_14252,N_14347);
or U20213 (N_20213,N_16213,N_17608);
and U20214 (N_20214,N_17897,N_13524);
nand U20215 (N_20215,N_15077,N_13821);
xnor U20216 (N_20216,N_16462,N_17750);
xnor U20217 (N_20217,N_17735,N_17665);
xor U20218 (N_20218,N_13028,N_12987);
nor U20219 (N_20219,N_17880,N_13492);
xnor U20220 (N_20220,N_16706,N_15771);
and U20221 (N_20221,N_17481,N_14479);
nor U20222 (N_20222,N_17234,N_12852);
nand U20223 (N_20223,N_16734,N_18332);
or U20224 (N_20224,N_17805,N_17278);
and U20225 (N_20225,N_12627,N_13422);
or U20226 (N_20226,N_16793,N_16189);
xor U20227 (N_20227,N_18026,N_17603);
nor U20228 (N_20228,N_17488,N_12748);
nor U20229 (N_20229,N_15548,N_13709);
or U20230 (N_20230,N_13067,N_16425);
and U20231 (N_20231,N_16036,N_13191);
and U20232 (N_20232,N_13569,N_16191);
and U20233 (N_20233,N_15421,N_16880);
or U20234 (N_20234,N_14398,N_18475);
or U20235 (N_20235,N_14016,N_18185);
nor U20236 (N_20236,N_16414,N_15013);
nor U20237 (N_20237,N_17660,N_17755);
and U20238 (N_20238,N_15488,N_17057);
xor U20239 (N_20239,N_15072,N_17406);
nor U20240 (N_20240,N_12648,N_15207);
xor U20241 (N_20241,N_15624,N_12569);
nor U20242 (N_20242,N_13860,N_17291);
xnor U20243 (N_20243,N_14664,N_18712);
nand U20244 (N_20244,N_18575,N_16193);
xor U20245 (N_20245,N_17164,N_15708);
xnor U20246 (N_20246,N_12629,N_12927);
xor U20247 (N_20247,N_18207,N_13843);
or U20248 (N_20248,N_16999,N_16132);
nor U20249 (N_20249,N_18060,N_14169);
or U20250 (N_20250,N_18057,N_13371);
or U20251 (N_20251,N_16307,N_18343);
xor U20252 (N_20252,N_14654,N_17446);
nand U20253 (N_20253,N_13668,N_14183);
nand U20254 (N_20254,N_13109,N_16907);
xor U20255 (N_20255,N_16732,N_17784);
or U20256 (N_20256,N_12592,N_12590);
nand U20257 (N_20257,N_16076,N_16197);
or U20258 (N_20258,N_18560,N_14787);
or U20259 (N_20259,N_13505,N_18149);
and U20260 (N_20260,N_17886,N_17738);
and U20261 (N_20261,N_13148,N_13597);
and U20262 (N_20262,N_16489,N_12660);
nand U20263 (N_20263,N_12842,N_16864);
and U20264 (N_20264,N_13887,N_12646);
xnor U20265 (N_20265,N_16886,N_18107);
xnor U20266 (N_20266,N_15581,N_13074);
nand U20267 (N_20267,N_16433,N_13116);
xor U20268 (N_20268,N_17907,N_17893);
nand U20269 (N_20269,N_16172,N_12908);
and U20270 (N_20270,N_16310,N_15413);
xor U20271 (N_20271,N_17540,N_14387);
xor U20272 (N_20272,N_17055,N_15987);
nand U20273 (N_20273,N_15546,N_12934);
xnor U20274 (N_20274,N_16848,N_14475);
xor U20275 (N_20275,N_12890,N_14704);
or U20276 (N_20276,N_15167,N_16702);
or U20277 (N_20277,N_14658,N_14700);
or U20278 (N_20278,N_13004,N_14195);
nor U20279 (N_20279,N_15025,N_13697);
and U20280 (N_20280,N_16657,N_17572);
or U20281 (N_20281,N_17657,N_13831);
or U20282 (N_20282,N_18726,N_16904);
and U20283 (N_20283,N_14455,N_18309);
xnor U20284 (N_20284,N_14410,N_17887);
and U20285 (N_20285,N_16919,N_16679);
nor U20286 (N_20286,N_14083,N_14648);
nand U20287 (N_20287,N_18365,N_14473);
and U20288 (N_20288,N_18508,N_16457);
or U20289 (N_20289,N_17704,N_14915);
nand U20290 (N_20290,N_15436,N_12640);
nand U20291 (N_20291,N_16889,N_16274);
or U20292 (N_20292,N_17522,N_17011);
nor U20293 (N_20293,N_13623,N_18049);
or U20294 (N_20294,N_14901,N_16167);
xor U20295 (N_20295,N_13553,N_12508);
or U20296 (N_20296,N_15097,N_15364);
nor U20297 (N_20297,N_16795,N_18259);
xnor U20298 (N_20298,N_18685,N_13767);
nand U20299 (N_20299,N_13544,N_15555);
and U20300 (N_20300,N_14236,N_18670);
or U20301 (N_20301,N_14615,N_12602);
nor U20302 (N_20302,N_15093,N_14182);
or U20303 (N_20303,N_13857,N_18714);
or U20304 (N_20304,N_15841,N_17364);
nor U20305 (N_20305,N_13912,N_14846);
or U20306 (N_20306,N_16914,N_18511);
nor U20307 (N_20307,N_14645,N_16720);
nand U20308 (N_20308,N_14097,N_18278);
and U20309 (N_20309,N_15815,N_15243);
nor U20310 (N_20310,N_14003,N_17469);
nand U20311 (N_20311,N_13397,N_15886);
and U20312 (N_20312,N_18375,N_15078);
nand U20313 (N_20313,N_13839,N_16219);
nor U20314 (N_20314,N_17473,N_14480);
xnor U20315 (N_20315,N_15330,N_18731);
nor U20316 (N_20316,N_17705,N_13529);
nand U20317 (N_20317,N_14546,N_16403);
and U20318 (N_20318,N_13041,N_15146);
nand U20319 (N_20319,N_18618,N_15747);
and U20320 (N_20320,N_14995,N_13068);
nor U20321 (N_20321,N_17162,N_17538);
or U20322 (N_20322,N_18356,N_13504);
xor U20323 (N_20323,N_13361,N_13876);
or U20324 (N_20324,N_17764,N_16364);
and U20325 (N_20325,N_12958,N_18391);
nand U20326 (N_20326,N_12645,N_17898);
and U20327 (N_20327,N_15574,N_14623);
or U20328 (N_20328,N_13883,N_16960);
nor U20329 (N_20329,N_17395,N_14082);
nand U20330 (N_20330,N_16032,N_15023);
and U20331 (N_20331,N_12625,N_14618);
nor U20332 (N_20332,N_18380,N_14476);
or U20333 (N_20333,N_16865,N_17966);
xnor U20334 (N_20334,N_17869,N_16140);
and U20335 (N_20335,N_17004,N_18032);
or U20336 (N_20336,N_13942,N_15773);
and U20337 (N_20337,N_18742,N_12756);
nand U20338 (N_20338,N_12545,N_13782);
and U20339 (N_20339,N_15582,N_17585);
and U20340 (N_20340,N_14883,N_18327);
nor U20341 (N_20341,N_18029,N_12879);
and U20342 (N_20342,N_17950,N_14507);
or U20343 (N_20343,N_16743,N_14301);
xor U20344 (N_20344,N_17440,N_18525);
xor U20345 (N_20345,N_14792,N_18430);
or U20346 (N_20346,N_17126,N_16007);
nor U20347 (N_20347,N_17269,N_14073);
or U20348 (N_20348,N_18166,N_17391);
and U20349 (N_20349,N_17195,N_18215);
nand U20350 (N_20350,N_15150,N_14287);
or U20351 (N_20351,N_14329,N_17462);
nand U20352 (N_20352,N_14034,N_18432);
nand U20353 (N_20353,N_13118,N_15658);
or U20354 (N_20354,N_14248,N_15603);
nor U20355 (N_20355,N_16913,N_17093);
and U20356 (N_20356,N_15618,N_14293);
or U20357 (N_20357,N_15598,N_18652);
or U20358 (N_20358,N_15460,N_15982);
or U20359 (N_20359,N_15467,N_16452);
nor U20360 (N_20360,N_18552,N_14668);
xor U20361 (N_20361,N_15024,N_17945);
nand U20362 (N_20362,N_18452,N_17036);
or U20363 (N_20363,N_14027,N_15299);
or U20364 (N_20364,N_17180,N_13729);
xnor U20365 (N_20365,N_15986,N_17793);
xor U20366 (N_20366,N_13159,N_12923);
xor U20367 (N_20367,N_17602,N_12613);
or U20368 (N_20368,N_15911,N_18669);
and U20369 (N_20369,N_15212,N_14581);
nor U20370 (N_20370,N_17851,N_18493);
xnor U20371 (N_20371,N_13197,N_17035);
or U20372 (N_20372,N_18419,N_16304);
and U20373 (N_20373,N_18078,N_15609);
and U20374 (N_20374,N_15136,N_15060);
xnor U20375 (N_20375,N_17056,N_14982);
nand U20376 (N_20376,N_15128,N_15068);
or U20377 (N_20377,N_12862,N_15099);
and U20378 (N_20378,N_17088,N_17853);
or U20379 (N_20379,N_14403,N_15006);
nand U20380 (N_20380,N_15015,N_15798);
nor U20381 (N_20381,N_17749,N_15657);
nand U20382 (N_20382,N_15278,N_14552);
xor U20383 (N_20383,N_14084,N_16072);
nand U20384 (N_20384,N_14267,N_14316);
nand U20385 (N_20385,N_13579,N_13593);
or U20386 (N_20386,N_17352,N_14593);
xnor U20387 (N_20387,N_12699,N_15539);
xnor U20388 (N_20388,N_13714,N_14650);
and U20389 (N_20389,N_17431,N_18295);
and U20390 (N_20390,N_13862,N_14580);
and U20391 (N_20391,N_14089,N_14853);
nor U20392 (N_20392,N_14215,N_15594);
nor U20393 (N_20393,N_13140,N_18555);
nand U20394 (N_20394,N_15221,N_17729);
and U20395 (N_20395,N_15554,N_18189);
or U20396 (N_20396,N_13720,N_13289);
nand U20397 (N_20397,N_18202,N_15007);
nor U20398 (N_20398,N_12666,N_16101);
and U20399 (N_20399,N_17994,N_16151);
and U20400 (N_20400,N_14041,N_18221);
or U20401 (N_20401,N_18320,N_13629);
xnor U20402 (N_20402,N_13462,N_13840);
xnor U20403 (N_20403,N_12790,N_16415);
nand U20404 (N_20404,N_17254,N_15923);
or U20405 (N_20405,N_16014,N_13740);
xor U20406 (N_20406,N_12651,N_14125);
and U20407 (N_20407,N_16312,N_14920);
or U20408 (N_20408,N_14441,N_12594);
nor U20409 (N_20409,N_15999,N_12541);
nor U20410 (N_20410,N_14063,N_12752);
nor U20411 (N_20411,N_16454,N_15738);
and U20412 (N_20412,N_15565,N_17902);
and U20413 (N_20413,N_18598,N_13164);
nor U20414 (N_20414,N_17615,N_14132);
nand U20415 (N_20415,N_15215,N_13900);
nand U20416 (N_20416,N_18641,N_12684);
or U20417 (N_20417,N_14208,N_17642);
nor U20418 (N_20418,N_15636,N_13620);
xnor U20419 (N_20419,N_18482,N_15938);
and U20420 (N_20420,N_14602,N_13089);
and U20421 (N_20421,N_18138,N_14206);
xnor U20422 (N_20422,N_14017,N_16379);
nor U20423 (N_20423,N_12751,N_18660);
and U20424 (N_20424,N_14682,N_14726);
or U20425 (N_20425,N_14055,N_13824);
nand U20426 (N_20426,N_12518,N_18749);
xor U20427 (N_20427,N_17047,N_16938);
nand U20428 (N_20428,N_15026,N_14771);
nor U20429 (N_20429,N_17516,N_17639);
and U20430 (N_20430,N_14657,N_14587);
nand U20431 (N_20431,N_13155,N_17543);
xor U20432 (N_20432,N_15640,N_12764);
nor U20433 (N_20433,N_18265,N_17016);
nand U20434 (N_20434,N_15661,N_15792);
and U20435 (N_20435,N_17620,N_14978);
and U20436 (N_20436,N_13881,N_14001);
nand U20437 (N_20437,N_16239,N_16445);
and U20438 (N_20438,N_18039,N_13270);
and U20439 (N_20439,N_16447,N_12965);
or U20440 (N_20440,N_12710,N_18043);
xor U20441 (N_20441,N_13488,N_13039);
or U20442 (N_20442,N_18732,N_18397);
and U20443 (N_20443,N_14492,N_18249);
and U20444 (N_20444,N_13940,N_18609);
nand U20445 (N_20445,N_14168,N_17351);
xor U20446 (N_20446,N_14639,N_12975);
and U20447 (N_20447,N_13265,N_15123);
nand U20448 (N_20448,N_13788,N_12932);
nand U20449 (N_20449,N_16175,N_12683);
or U20450 (N_20450,N_13208,N_13431);
nor U20451 (N_20451,N_12546,N_15465);
nor U20452 (N_20452,N_18270,N_17302);
and U20453 (N_20453,N_16100,N_13467);
nor U20454 (N_20454,N_18604,N_15684);
xnor U20455 (N_20455,N_12506,N_15649);
nor U20456 (N_20456,N_15018,N_14449);
and U20457 (N_20457,N_16426,N_12650);
nand U20458 (N_20458,N_17958,N_16455);
and U20459 (N_20459,N_15879,N_16937);
or U20460 (N_20460,N_17074,N_16946);
xnor U20461 (N_20461,N_12773,N_15585);
xor U20462 (N_20462,N_17411,N_17573);
nand U20463 (N_20463,N_13203,N_18045);
and U20464 (N_20464,N_16844,N_15972);
nand U20465 (N_20465,N_16117,N_14827);
xnor U20466 (N_20466,N_12705,N_15912);
nand U20467 (N_20467,N_14545,N_17881);
and U20468 (N_20468,N_14887,N_13384);
nor U20469 (N_20469,N_15075,N_18462);
xor U20470 (N_20470,N_15873,N_16352);
nor U20471 (N_20471,N_14591,N_17982);
nand U20472 (N_20472,N_13452,N_18280);
and U20473 (N_20473,N_13403,N_15139);
nor U20474 (N_20474,N_15943,N_18173);
nor U20475 (N_20475,N_14937,N_16666);
nand U20476 (N_20476,N_16332,N_17187);
nand U20477 (N_20477,N_14025,N_16049);
and U20478 (N_20478,N_14210,N_14659);
xor U20479 (N_20479,N_17717,N_13537);
nor U20480 (N_20480,N_15037,N_13848);
nor U20481 (N_20481,N_12552,N_13506);
and U20482 (N_20482,N_14009,N_13858);
nor U20483 (N_20483,N_16383,N_18305);
xor U20484 (N_20484,N_12599,N_12596);
or U20485 (N_20485,N_17414,N_16608);
nand U20486 (N_20486,N_15961,N_14060);
and U20487 (N_20487,N_16174,N_13989);
nor U20488 (N_20488,N_17434,N_15681);
xnor U20489 (N_20489,N_17491,N_16843);
nor U20490 (N_20490,N_16347,N_15392);
nor U20491 (N_20491,N_16225,N_17565);
or U20492 (N_20492,N_18155,N_16714);
xnor U20493 (N_20493,N_16707,N_17596);
nand U20494 (N_20494,N_14462,N_13588);
and U20495 (N_20495,N_17813,N_14926);
xor U20496 (N_20496,N_15878,N_12887);
nor U20497 (N_20497,N_15813,N_14601);
nor U20498 (N_20498,N_12722,N_15903);
or U20499 (N_20499,N_16063,N_12745);
or U20500 (N_20500,N_16861,N_18379);
xor U20501 (N_20501,N_16533,N_13543);
or U20502 (N_20502,N_16690,N_16778);
nand U20503 (N_20503,N_15489,N_16437);
nor U20504 (N_20504,N_17724,N_12813);
or U20505 (N_20505,N_14662,N_16697);
nand U20506 (N_20506,N_14954,N_15682);
nand U20507 (N_20507,N_15625,N_14343);
nand U20508 (N_20508,N_13096,N_15280);
or U20509 (N_20509,N_14322,N_15365);
xnor U20510 (N_20510,N_12568,N_18106);
xor U20511 (N_20511,N_18017,N_15869);
nor U20512 (N_20512,N_18081,N_15173);
and U20513 (N_20513,N_13750,N_16557);
or U20514 (N_20514,N_15400,N_12964);
or U20515 (N_20515,N_13135,N_16764);
nand U20516 (N_20516,N_15160,N_18349);
nor U20517 (N_20517,N_17340,N_18409);
xor U20518 (N_20518,N_18036,N_16566);
or U20519 (N_20519,N_13117,N_17228);
and U20520 (N_20520,N_16123,N_17131);
nor U20521 (N_20521,N_13819,N_18360);
and U20522 (N_20522,N_17650,N_13835);
nand U20523 (N_20523,N_14689,N_12539);
xor U20524 (N_20524,N_13878,N_18268);
xnor U20525 (N_20525,N_15175,N_17277);
or U20526 (N_20526,N_15604,N_12548);
nand U20527 (N_20527,N_15676,N_13426);
nor U20528 (N_20528,N_16089,N_14968);
or U20529 (N_20529,N_16885,N_13365);
and U20530 (N_20530,N_13419,N_15633);
nor U20531 (N_20531,N_12515,N_13193);
nand U20532 (N_20532,N_17709,N_13071);
or U20533 (N_20533,N_17971,N_15522);
or U20534 (N_20534,N_18602,N_14932);
xor U20535 (N_20535,N_17952,N_17923);
or U20536 (N_20536,N_13277,N_18334);
nand U20537 (N_20537,N_17534,N_15757);
xnor U20538 (N_20538,N_14371,N_16939);
xor U20539 (N_20539,N_18632,N_14858);
and U20540 (N_20540,N_13724,N_14414);
and U20541 (N_20541,N_17181,N_12687);
nand U20542 (N_20542,N_17939,N_14363);
and U20543 (N_20543,N_13827,N_14261);
nand U20544 (N_20544,N_14184,N_13865);
and U20545 (N_20545,N_13418,N_14906);
or U20546 (N_20546,N_18556,N_16150);
and U20547 (N_20547,N_17906,N_16613);
nor U20548 (N_20548,N_17092,N_18597);
or U20549 (N_20549,N_14871,N_12540);
nand U20550 (N_20550,N_17135,N_14114);
nand U20551 (N_20551,N_13792,N_16058);
nor U20552 (N_20552,N_14255,N_13818);
xor U20553 (N_20553,N_16520,N_13669);
or U20554 (N_20554,N_16794,N_16209);
xnor U20555 (N_20555,N_18447,N_16867);
and U20556 (N_20556,N_16887,N_18279);
xnor U20557 (N_20557,N_12550,N_16890);
nand U20558 (N_20558,N_16118,N_13025);
xnor U20559 (N_20559,N_12902,N_12652);
nand U20560 (N_20560,N_16147,N_14809);
nor U20561 (N_20561,N_13463,N_17957);
nand U20562 (N_20562,N_15327,N_16399);
and U20563 (N_20563,N_13026,N_14024);
nor U20564 (N_20564,N_17166,N_13847);
or U20565 (N_20565,N_13202,N_17182);
nand U20566 (N_20566,N_13701,N_13652);
nand U20567 (N_20567,N_13555,N_17320);
nand U20568 (N_20568,N_17757,N_16983);
nor U20569 (N_20569,N_16112,N_13717);
and U20570 (N_20570,N_14241,N_14065);
nand U20571 (N_20571,N_16853,N_13809);
or U20572 (N_20572,N_17222,N_17664);
nand U20573 (N_20573,N_14179,N_16223);
xor U20574 (N_20574,N_14448,N_16287);
and U20575 (N_20575,N_17763,N_14876);
nand U20576 (N_20576,N_12970,N_13051);
nand U20577 (N_20577,N_16998,N_18737);
and U20578 (N_20578,N_15122,N_18675);
nand U20579 (N_20579,N_18746,N_18346);
nor U20580 (N_20580,N_17619,N_14577);
and U20581 (N_20581,N_14186,N_14610);
nand U20582 (N_20582,N_15042,N_15144);
and U20583 (N_20583,N_13700,N_15672);
nor U20584 (N_20584,N_13654,N_15206);
nor U20585 (N_20585,N_15854,N_13551);
xnor U20586 (N_20586,N_16475,N_15549);
nand U20587 (N_20587,N_14574,N_14103);
and U20588 (N_20588,N_18403,N_12815);
nand U20589 (N_20589,N_14568,N_13577);
nand U20590 (N_20590,N_12830,N_14088);
or U20591 (N_20591,N_13993,N_15195);
or U20592 (N_20592,N_15689,N_13934);
xor U20593 (N_20593,N_16082,N_16359);
nand U20594 (N_20594,N_12774,N_18446);
xnor U20595 (N_20595,N_16785,N_14279);
and U20596 (N_20596,N_14665,N_16643);
nand U20597 (N_20597,N_16320,N_14044);
xnor U20598 (N_20598,N_17792,N_12689);
nor U20599 (N_20599,N_16667,N_18622);
nor U20600 (N_20600,N_15073,N_14789);
nand U20601 (N_20601,N_17846,N_15444);
xor U20602 (N_20602,N_18234,N_18455);
or U20603 (N_20603,N_15102,N_14176);
or U20604 (N_20604,N_13081,N_18073);
and U20605 (N_20605,N_14397,N_18615);
nor U20606 (N_20606,N_16774,N_13676);
and U20607 (N_20607,N_15659,N_13493);
nand U20608 (N_20608,N_16685,N_15889);
and U20609 (N_20609,N_18708,N_16074);
xnor U20610 (N_20610,N_14265,N_18414);
and U20611 (N_20611,N_17909,N_14616);
or U20612 (N_20612,N_14231,N_13898);
nor U20613 (N_20613,N_16529,N_17941);
xor U20614 (N_20614,N_14560,N_14776);
nor U20615 (N_20615,N_13845,N_16143);
or U20616 (N_20616,N_17947,N_15551);
and U20617 (N_20617,N_14669,N_14589);
nand U20618 (N_20618,N_16696,N_18449);
and U20619 (N_20619,N_14291,N_17988);
nor U20620 (N_20620,N_13521,N_13377);
or U20621 (N_20621,N_17980,N_16052);
or U20622 (N_20622,N_18643,N_15838);
nor U20623 (N_20623,N_14582,N_14559);
nor U20624 (N_20624,N_17703,N_16381);
xor U20625 (N_20625,N_16962,N_14136);
xor U20626 (N_20626,N_14698,N_15131);
xnor U20627 (N_20627,N_17861,N_15595);
nor U20628 (N_20628,N_13178,N_13035);
nor U20629 (N_20629,N_18398,N_17760);
or U20630 (N_20630,N_15669,N_16115);
nor U20631 (N_20631,N_15163,N_14074);
and U20632 (N_20632,N_13784,N_14964);
nand U20633 (N_20633,N_18085,N_18194);
nor U20634 (N_20634,N_16991,N_14785);
nor U20635 (N_20635,N_15082,N_16989);
or U20636 (N_20636,N_15437,N_13769);
nand U20637 (N_20637,N_14539,N_12892);
and U20638 (N_20638,N_15391,N_16479);
nand U20639 (N_20639,N_13923,N_17550);
nor U20640 (N_20640,N_14742,N_14115);
nor U20641 (N_20641,N_13018,N_16627);
nor U20642 (N_20642,N_15260,N_16244);
or U20643 (N_20643,N_16401,N_14054);
nor U20644 (N_20644,N_16260,N_13917);
or U20645 (N_20645,N_15267,N_17811);
nand U20646 (N_20646,N_16203,N_15249);
and U20647 (N_20647,N_14845,N_14543);
xnor U20648 (N_20648,N_14720,N_17832);
nor U20649 (N_20649,N_12701,N_15786);
and U20650 (N_20650,N_12918,N_13334);
nor U20651 (N_20651,N_13817,N_15637);
and U20652 (N_20652,N_15230,N_13616);
or U20653 (N_20653,N_15643,N_18011);
nand U20654 (N_20654,N_15242,N_16532);
xor U20655 (N_20655,N_15890,N_14269);
and U20656 (N_20656,N_14814,N_17843);
or U20657 (N_20657,N_17908,N_18385);
or U20658 (N_20658,N_13167,N_12610);
nor U20659 (N_20659,N_15003,N_13479);
xor U20660 (N_20660,N_16368,N_17468);
nand U20661 (N_20661,N_16281,N_17889);
nor U20662 (N_20662,N_15933,N_18485);
nor U20663 (N_20663,N_16110,N_18633);
or U20664 (N_20664,N_14794,N_16031);
and U20665 (N_20665,N_17936,N_13622);
and U20666 (N_20666,N_18506,N_15750);
xnor U20667 (N_20667,N_14094,N_14076);
nor U20668 (N_20668,N_17539,N_15113);
and U20669 (N_20669,N_14928,N_16263);
or U20670 (N_20670,N_17260,N_12864);
or U20671 (N_20671,N_17959,N_17802);
nand U20672 (N_20672,N_15731,N_14628);
xor U20673 (N_20673,N_12595,N_13485);
xor U20674 (N_20674,N_13918,N_17803);
xor U20675 (N_20675,N_18437,N_14141);
and U20676 (N_20676,N_13196,N_17561);
nand U20677 (N_20677,N_15422,N_16682);
nor U20678 (N_20678,N_13386,N_16311);
xnor U20679 (N_20679,N_15888,N_15088);
nor U20680 (N_20680,N_14484,N_13754);
and U20681 (N_20681,N_13688,N_17800);
nand U20682 (N_20682,N_12523,N_13600);
and U20683 (N_20683,N_16510,N_13325);
and U20684 (N_20684,N_13951,N_12556);
xnor U20685 (N_20685,N_15717,N_16698);
or U20686 (N_20686,N_14151,N_15663);
nand U20687 (N_20687,N_13447,N_14997);
xor U20688 (N_20688,N_17213,N_15033);
nor U20689 (N_20689,N_15198,N_15880);
and U20690 (N_20690,N_14274,N_15205);
or U20691 (N_20691,N_17132,N_16728);
xnor U20692 (N_20692,N_17179,N_13472);
nand U20693 (N_20693,N_16234,N_14715);
nor U20694 (N_20694,N_17452,N_17174);
xnor U20695 (N_20695,N_14962,N_17104);
nor U20696 (N_20696,N_12893,N_12844);
or U20697 (N_20697,N_15227,N_15145);
xor U20698 (N_20698,N_15204,N_13664);
xnor U20699 (N_20699,N_16892,N_17420);
and U20700 (N_20700,N_13213,N_16294);
or U20701 (N_20701,N_14661,N_15268);
and U20702 (N_20702,N_14840,N_14338);
xor U20703 (N_20703,N_15076,N_15700);
nor U20704 (N_20704,N_15766,N_13158);
or U20705 (N_20705,N_18502,N_17782);
or U20706 (N_20706,N_13152,N_18195);
xor U20707 (N_20707,N_12670,N_12732);
or U20708 (N_20708,N_14330,N_18317);
or U20709 (N_20709,N_12867,N_13027);
or U20710 (N_20710,N_13232,N_14340);
xor U20711 (N_20711,N_13950,N_15418);
and U20712 (N_20712,N_14617,N_13294);
xnor U20713 (N_20713,N_15240,N_12707);
xnor U20714 (N_20714,N_12994,N_16687);
and U20715 (N_20715,N_16046,N_12880);
xor U20716 (N_20716,N_13217,N_16285);
nor U20717 (N_20717,N_16487,N_18277);
and U20718 (N_20718,N_14813,N_18208);
nor U20719 (N_20719,N_16640,N_18600);
nand U20720 (N_20720,N_17096,N_13223);
or U20721 (N_20721,N_14170,N_18171);
xor U20722 (N_20722,N_15067,N_13460);
and U20723 (N_20723,N_16840,N_18489);
nor U20724 (N_20724,N_18492,N_14384);
nand U20725 (N_20725,N_13647,N_17337);
nand U20726 (N_20726,N_13351,N_17747);
xnor U20727 (N_20727,N_13879,N_17323);
nand U20728 (N_20728,N_17250,N_16539);
or U20729 (N_20729,N_14028,N_17084);
nor U20730 (N_20730,N_16300,N_18526);
xnor U20731 (N_20731,N_16759,N_18547);
nand U20732 (N_20732,N_16849,N_13465);
xnor U20733 (N_20733,N_17661,N_16431);
and U20734 (N_20734,N_12823,N_17951);
xor U20735 (N_20735,N_14004,N_15209);
xnor U20736 (N_20736,N_16217,N_15724);
xnor U20737 (N_20737,N_14531,N_18374);
nand U20738 (N_20738,N_14461,N_14841);
xor U20739 (N_20739,N_13037,N_17990);
nor U20740 (N_20740,N_14006,N_13395);
xnor U20741 (N_20741,N_18378,N_18178);
xor U20742 (N_20742,N_18121,N_15035);
nand U20743 (N_20743,N_15151,N_14204);
and U20744 (N_20744,N_16994,N_15380);
or U20745 (N_20745,N_15354,N_15030);
xor U20746 (N_20746,N_18748,N_14733);
or U20747 (N_20747,N_16176,N_13534);
nand U20748 (N_20748,N_13052,N_13542);
and U20749 (N_20749,N_14699,N_18263);
or U20750 (N_20750,N_18324,N_16059);
and U20751 (N_20751,N_17531,N_13383);
nand U20752 (N_20752,N_18023,N_12589);
xnor U20753 (N_20753,N_14013,N_12747);
and U20754 (N_20754,N_12784,N_13673);
nand U20755 (N_20755,N_14471,N_14420);
nor U20756 (N_20756,N_12620,N_15462);
nor U20757 (N_20757,N_18469,N_13111);
nand U20758 (N_20758,N_14634,N_13549);
or U20759 (N_20759,N_14849,N_14177);
nor U20760 (N_20760,N_16283,N_15096);
and U20761 (N_20761,N_13536,N_13559);
nor U20762 (N_20762,N_15897,N_15641);
nor U20763 (N_20763,N_18672,N_13043);
and U20764 (N_20764,N_13970,N_16538);
and U20765 (N_20765,N_18619,N_13330);
nor U20766 (N_20766,N_13998,N_13281);
nor U20767 (N_20767,N_16158,N_15955);
xor U20768 (N_20768,N_18013,N_14780);
xor U20769 (N_20769,N_13901,N_14843);
and U20770 (N_20770,N_13550,N_15977);
nand U20771 (N_20771,N_15722,N_14922);
nor U20772 (N_20772,N_18035,N_14799);
nor U20773 (N_20773,N_13932,N_13719);
xnor U20774 (N_20774,N_15686,N_15449);
nand U20775 (N_20775,N_14605,N_17169);
or U20776 (N_20776,N_13899,N_16185);
nand U20777 (N_20777,N_18050,N_15991);
or U20778 (N_20778,N_17591,N_14655);
nand U20779 (N_20779,N_18471,N_17571);
and U20780 (N_20780,N_12588,N_15405);
xnor U20781 (N_20781,N_13286,N_15675);
nor U20782 (N_20782,N_16003,N_13591);
and U20783 (N_20783,N_14309,N_14940);
or U20784 (N_20784,N_16882,N_15805);
and U20785 (N_20785,N_16873,N_17624);
nor U20786 (N_20786,N_15949,N_12584);
nor U20787 (N_20787,N_14415,N_16135);
and U20788 (N_20788,N_17141,N_12604);
or U20789 (N_20789,N_13396,N_17932);
and U20790 (N_20790,N_14198,N_15101);
nor U20791 (N_20791,N_13291,N_15387);
and U20792 (N_20792,N_17014,N_15651);
nor U20793 (N_20793,N_17379,N_12503);
nor U20794 (N_20794,N_16829,N_14885);
nor U20795 (N_20795,N_16138,N_16797);
and U20796 (N_20796,N_16972,N_15983);
and U20797 (N_20797,N_14656,N_17637);
or U20798 (N_20798,N_14394,N_13928);
xnor U20799 (N_20799,N_16680,N_15385);
and U20800 (N_20800,N_18109,N_13692);
nor U20801 (N_20801,N_17232,N_18192);
and U20802 (N_20802,N_15780,N_12804);
nand U20803 (N_20803,N_16522,N_17570);
nand U20804 (N_20804,N_15989,N_16818);
nor U20805 (N_20805,N_16068,N_18038);
xor U20806 (N_20806,N_18120,N_13721);
nor U20807 (N_20807,N_15995,N_18564);
xnor U20808 (N_20808,N_17430,N_16131);
xnor U20809 (N_20809,N_16800,N_13024);
or U20810 (N_20810,N_14555,N_12851);
nand U20811 (N_20811,N_15228,N_16622);
xnor U20812 (N_20812,N_14848,N_15171);
or U20813 (N_20813,N_12869,N_17772);
and U20814 (N_20814,N_17425,N_16303);
nor U20815 (N_20815,N_18381,N_13564);
or U20816 (N_20816,N_17622,N_15909);
or U20817 (N_20817,N_16514,N_14366);
or U20818 (N_20818,N_15061,N_17807);
nor U20819 (N_20819,N_18637,N_15905);
and U20820 (N_20820,N_14888,N_14417);
and U20821 (N_20821,N_14253,N_17535);
xor U20822 (N_20822,N_18369,N_18657);
xnor U20823 (N_20823,N_13611,N_14467);
or U20824 (N_20824,N_13246,N_13468);
nor U20825 (N_20825,N_16740,N_16944);
xor U20826 (N_20826,N_15898,N_17588);
nor U20827 (N_20827,N_18184,N_17486);
or U20828 (N_20828,N_18739,N_13808);
nand U20829 (N_20829,N_17329,N_12811);
nor U20830 (N_20830,N_12708,N_12529);
nand U20831 (N_20831,N_16721,N_15966);
or U20832 (N_20832,N_14077,N_16857);
nor U20833 (N_20833,N_17483,N_16061);
or U20834 (N_20834,N_16406,N_13413);
nor U20835 (N_20835,N_14250,N_17417);
xor U20836 (N_20836,N_16473,N_17720);
xor U20837 (N_20837,N_16091,N_12877);
nor U20838 (N_20838,N_14396,N_18152);
nor U20839 (N_20839,N_18509,N_13635);
xor U20840 (N_20840,N_12765,N_14925);
nor U20841 (N_20841,N_16365,N_18744);
nand U20842 (N_20842,N_12870,N_15219);
nand U20843 (N_20843,N_13393,N_18241);
nand U20844 (N_20844,N_17701,N_16404);
xnor U20845 (N_20845,N_14112,N_18237);
nand U20846 (N_20846,N_15189,N_18174);
nand U20847 (N_20847,N_14264,N_15417);
nand U20848 (N_20848,N_17989,N_18716);
nand U20849 (N_20849,N_12534,N_18400);
nor U20850 (N_20850,N_14495,N_12847);
or U20851 (N_20851,N_18427,N_13685);
or U20852 (N_20852,N_15899,N_15628);
or U20853 (N_20853,N_18125,N_15412);
xnor U20854 (N_20854,N_14061,N_18071);
xnor U20855 (N_20855,N_15420,N_14674);
and U20856 (N_20856,N_17280,N_13107);
or U20857 (N_20857,N_13599,N_15590);
nor U20858 (N_20858,N_16748,N_15526);
or U20859 (N_20859,N_15314,N_12980);
and U20860 (N_20860,N_15143,N_16726);
xor U20861 (N_20861,N_14379,N_18313);
and U20862 (N_20862,N_14300,N_18569);
nand U20863 (N_20863,N_17943,N_17771);
xnor U20864 (N_20864,N_14311,N_15169);
and U20865 (N_20865,N_14348,N_15155);
xor U20866 (N_20866,N_14099,N_13578);
xnor U20867 (N_20867,N_14050,N_13108);
and U20868 (N_20868,N_13015,N_12983);
and U20869 (N_20869,N_15439,N_15271);
and U20870 (N_20870,N_15158,N_16806);
nor U20871 (N_20871,N_15313,N_17870);
and U20872 (N_20872,N_14527,N_17203);
nand U20873 (N_20873,N_16480,N_12575);
and U20874 (N_20874,N_12822,N_17584);
and U20875 (N_20875,N_17316,N_13975);
nand U20876 (N_20876,N_13170,N_15656);
nand U20877 (N_20877,N_18533,N_13864);
xnor U20878 (N_20878,N_14775,N_16376);
nand U20879 (N_20879,N_14175,N_15335);
or U20880 (N_20880,N_17044,N_16343);
or U20881 (N_20881,N_17367,N_17354);
and U20882 (N_20882,N_14890,N_16390);
nand U20883 (N_20883,N_15723,N_18150);
or U20884 (N_20884,N_17448,N_17033);
xnor U20885 (N_20885,N_14292,N_15790);
nor U20886 (N_20886,N_13333,N_14468);
xor U20887 (N_20887,N_16341,N_17267);
nor U20888 (N_20888,N_14383,N_14312);
nand U20889 (N_20889,N_12578,N_17238);
and U20890 (N_20890,N_14418,N_16638);
and U20891 (N_20891,N_12672,N_18421);
xnor U20892 (N_20892,N_12580,N_18300);
or U20893 (N_20893,N_13765,N_16675);
and U20894 (N_20894,N_16077,N_16583);
and U20895 (N_20895,N_17859,N_17188);
and U20896 (N_20896,N_15781,N_16497);
or U20897 (N_20897,N_18674,N_17998);
or U20898 (N_20898,N_13926,N_17125);
nand U20899 (N_20899,N_15857,N_15510);
and U20900 (N_20900,N_15494,N_18534);
xnor U20901 (N_20901,N_13707,N_15081);
or U20902 (N_20902,N_13308,N_15644);
nand U20903 (N_20903,N_16524,N_17844);
nor U20904 (N_20904,N_17827,N_17493);
xor U20905 (N_20905,N_17723,N_13801);
and U20906 (N_20906,N_18518,N_14108);
or U20907 (N_20907,N_15614,N_16180);
or U20908 (N_20908,N_14900,N_17678);
or U20909 (N_20909,N_17317,N_18282);
and U20910 (N_20910,N_15086,N_16361);
nor U20911 (N_20911,N_17374,N_16257);
nand U20912 (N_20912,N_13188,N_14303);
or U20913 (N_20913,N_15882,N_12649);
xnor U20914 (N_20914,N_17433,N_18134);
xor U20915 (N_20915,N_14728,N_12655);
and U20916 (N_20916,N_13416,N_16811);
and U20917 (N_20917,N_17786,N_18722);
nor U20918 (N_20918,N_15848,N_18605);
nor U20919 (N_20919,N_12728,N_18297);
or U20920 (N_20920,N_17121,N_12686);
xor U20921 (N_20921,N_15390,N_16651);
nor U20922 (N_20922,N_17623,N_15990);
nor U20923 (N_20923,N_14711,N_16095);
and U20924 (N_20924,N_16192,N_16813);
and U20925 (N_20925,N_13082,N_13713);
or U20926 (N_20926,N_15579,N_16681);
nor U20927 (N_20927,N_16787,N_18541);
and U20928 (N_20928,N_15118,N_12950);
and U20929 (N_20929,N_15322,N_13914);
or U20930 (N_20930,N_16427,N_17451);
xor U20931 (N_20931,N_17429,N_16029);
and U20932 (N_20932,N_13094,N_15498);
nand U20933 (N_20933,N_16327,N_14676);
nand U20934 (N_20934,N_13682,N_17445);
or U20935 (N_20935,N_15232,N_14875);
nand U20936 (N_20936,N_15084,N_15726);
xor U20937 (N_20937,N_15283,N_16128);
and U20938 (N_20938,N_15162,N_17114);
nor U20939 (N_20939,N_15540,N_15887);
xnor U20940 (N_20940,N_12839,N_18197);
nor U20941 (N_20941,N_16788,N_16828);
and U20942 (N_20942,N_13412,N_16348);
and U20943 (N_20943,N_14453,N_12626);
nor U20944 (N_20944,N_12669,N_16113);
xnor U20945 (N_20945,N_14882,N_14450);
or U20946 (N_20946,N_13315,N_12559);
and U20947 (N_20947,N_17725,N_16382);
and U20948 (N_20948,N_17558,N_14701);
and U20949 (N_20949,N_18126,N_14781);
nand U20950 (N_20950,N_13406,N_18130);
nor U20951 (N_20951,N_16606,N_13609);
nand U20952 (N_20952,N_18367,N_13806);
and U20953 (N_20953,N_13662,N_13040);
nor U20954 (N_20954,N_17006,N_16316);
nor U20955 (N_20955,N_14317,N_15157);
and U20956 (N_20956,N_14513,N_14988);
nand U20957 (N_20957,N_12991,N_18161);
and U20958 (N_20958,N_18578,N_18316);
xor U20959 (N_20959,N_15610,N_13093);
nand U20960 (N_20960,N_13856,N_18562);
nor U20961 (N_20961,N_15602,N_13756);
or U20962 (N_20962,N_14469,N_13360);
xnor U20963 (N_20963,N_15154,N_18610);
or U20964 (N_20964,N_16617,N_12725);
xor U20965 (N_20965,N_12678,N_18595);
nor U20966 (N_20966,N_16159,N_14879);
nand U20967 (N_20967,N_14725,N_17842);
xor U20968 (N_20968,N_17883,N_13404);
nand U20969 (N_20969,N_14905,N_13300);
or U20970 (N_20970,N_18144,N_16355);
nor U20971 (N_20971,N_16527,N_17168);
xor U20972 (N_20972,N_12616,N_18683);
nand U20973 (N_20973,N_15348,N_13332);
nor U20974 (N_20974,N_15743,N_15802);
and U20975 (N_20975,N_15305,N_17809);
or U20976 (N_20976,N_14830,N_15849);
and U20977 (N_20977,N_16148,N_17528);
nor U20978 (N_20978,N_15491,N_13000);
xnor U20979 (N_20979,N_13316,N_13016);
nor U20980 (N_20980,N_18101,N_16633);
xor U20981 (N_20981,N_15161,N_13480);
or U20982 (N_20982,N_16604,N_14087);
nor U20983 (N_20983,N_17863,N_13749);
xor U20984 (N_20984,N_15403,N_16928);
and U20985 (N_20985,N_16526,N_14289);
nor U20986 (N_20986,N_18217,N_14953);
or U20987 (N_20987,N_17658,N_16221);
and U20988 (N_20988,N_15589,N_16796);
or U20989 (N_20989,N_17076,N_16130);
nor U20990 (N_20990,N_17444,N_17926);
and U20991 (N_20991,N_16202,N_15521);
and U20992 (N_20992,N_18693,N_14747);
or U20993 (N_20993,N_14909,N_13234);
xnor U20994 (N_20994,N_15363,N_15451);
or U20995 (N_20995,N_16504,N_18067);
and U20996 (N_20996,N_17783,N_13770);
or U20997 (N_20997,N_18634,N_16572);
and U20998 (N_20998,N_16534,N_15255);
xnor U20999 (N_20999,N_15883,N_13359);
nand U21000 (N_21000,N_17985,N_13540);
xor U21001 (N_21001,N_18413,N_18721);
xor U21002 (N_21002,N_13943,N_13225);
nand U21003 (N_21003,N_16092,N_16852);
nand U21004 (N_21004,N_13352,N_16996);
xor U21005 (N_21005,N_15758,N_12899);
and U21006 (N_21006,N_18477,N_13530);
nor U21007 (N_21007,N_13250,N_14494);
and U21008 (N_21008,N_17271,N_12634);
xnor U21009 (N_21009,N_15596,N_14993);
nand U21010 (N_21010,N_13145,N_13575);
nor U21011 (N_21011,N_12516,N_18310);
nand U21012 (N_21012,N_13704,N_13751);
nor U21013 (N_21013,N_12542,N_13173);
nand U21014 (N_21014,N_13690,N_15341);
or U21015 (N_21015,N_14596,N_13672);
xor U21016 (N_21016,N_16299,N_16876);
xnor U21017 (N_21017,N_16127,N_13271);
xor U21018 (N_21018,N_14167,N_15997);
xor U21019 (N_21019,N_15533,N_18272);
nand U21020 (N_21020,N_17053,N_17477);
nand U21021 (N_21021,N_13176,N_15317);
xnor U21022 (N_21022,N_13273,N_14346);
or U21023 (N_21023,N_14802,N_18256);
nor U21024 (N_21024,N_13778,N_12605);
nand U21025 (N_21025,N_16701,N_16942);
nor U21026 (N_21026,N_15580,N_16513);
and U21027 (N_21027,N_16284,N_14474);
nand U21028 (N_21028,N_13483,N_15165);
nand U21029 (N_21029,N_14361,N_16065);
nand U21030 (N_21030,N_18019,N_17900);
or U21031 (N_21031,N_14996,N_13716);
nand U21032 (N_21032,N_16451,N_13885);
or U21033 (N_21033,N_16603,N_15423);
or U21034 (N_21034,N_13080,N_14426);
or U21035 (N_21035,N_14395,N_14160);
or U21036 (N_21036,N_13658,N_15950);
xnor U21037 (N_21037,N_18027,N_16854);
nand U21038 (N_21038,N_16024,N_17617);
nor U21039 (N_21039,N_14244,N_13615);
xnor U21040 (N_21040,N_17777,N_14481);
nor U21041 (N_21041,N_16251,N_14923);
nand U21042 (N_21042,N_17144,N_13296);
and U21043 (N_21043,N_15680,N_18156);
and U21044 (N_21044,N_17722,N_15926);
nor U21045 (N_21045,N_15583,N_14181);
and U21046 (N_21046,N_13791,N_18056);
nor U21047 (N_21047,N_16139,N_16129);
or U21048 (N_21048,N_14355,N_13523);
or U21049 (N_21049,N_14666,N_15210);
xor U21050 (N_21050,N_16894,N_12957);
nand U21051 (N_21051,N_13256,N_16516);
xor U21052 (N_21052,N_15041,N_18046);
xor U21053 (N_21053,N_12631,N_17407);
and U21054 (N_21054,N_14749,N_16040);
and U21055 (N_21055,N_14171,N_14693);
or U21056 (N_21056,N_12505,N_14443);
xor U21057 (N_21057,N_14939,N_17295);
nand U21058 (N_21058,N_13752,N_13785);
and U21059 (N_21059,N_18323,N_15523);
nor U21060 (N_21060,N_12848,N_13757);
nand U21061 (N_21061,N_14105,N_16898);
or U21062 (N_21062,N_13216,N_16471);
xnor U21063 (N_21063,N_12579,N_17868);
or U21064 (N_21064,N_18386,N_15256);
nor U21065 (N_21065,N_16587,N_17706);
xor U21066 (N_21066,N_16136,N_13401);
and U21067 (N_21067,N_14245,N_14976);
or U21068 (N_21068,N_12949,N_17515);
nand U21069 (N_21069,N_18007,N_17065);
or U21070 (N_21070,N_12609,N_13387);
xor U21071 (N_21071,N_18519,N_13424);
nand U21072 (N_21072,N_13309,N_13439);
or U21073 (N_21073,N_13759,N_15147);
xor U21074 (N_21074,N_18169,N_13190);
or U21075 (N_21075,N_12656,N_17628);
nand U21076 (N_21076,N_15028,N_17756);
nand U21077 (N_21077,N_14847,N_13633);
nor U21078 (N_21078,N_15250,N_14227);
or U21079 (N_21079,N_16198,N_17328);
or U21080 (N_21080,N_15934,N_14098);
nand U21081 (N_21081,N_15830,N_14736);
or U21082 (N_21082,N_16196,N_15241);
and U21083 (N_21083,N_14161,N_18373);
xnor U21084 (N_21084,N_18204,N_17362);
or U21085 (N_21085,N_15529,N_12808);
and U21086 (N_21086,N_12826,N_15049);
nor U21087 (N_21087,N_17683,N_12525);
nand U21088 (N_21088,N_16226,N_12574);
xnor U21089 (N_21089,N_13304,N_15559);
nor U21090 (N_21090,N_13078,N_17236);
nor U21091 (N_21091,N_17644,N_13997);
nand U21092 (N_21092,N_17590,N_15517);
and U21093 (N_21093,N_17172,N_15562);
nor U21094 (N_21094,N_18157,N_17555);
and U21095 (N_21095,N_17396,N_13204);
nand U21096 (N_21096,N_14295,N_13621);
or U21097 (N_21097,N_12593,N_15095);
nand U21098 (N_21098,N_14692,N_15262);
nand U21099 (N_21099,N_14199,N_16392);
or U21100 (N_21100,N_17105,N_13101);
or U21101 (N_21101,N_14958,N_15411);
xnor U21102 (N_21102,N_16742,N_12742);
nand U21103 (N_21103,N_17511,N_16484);
nand U21104 (N_21104,N_17938,N_16073);
nand U21105 (N_21105,N_17007,N_18592);
and U21106 (N_21106,N_15116,N_17484);
and U21107 (N_21107,N_13149,N_13061);
and U21108 (N_21108,N_14686,N_17442);
nor U21109 (N_21109,N_13702,N_18703);
nand U21110 (N_21110,N_13971,N_16786);
xnor U21111 (N_21111,N_18697,N_14310);
nand U21112 (N_21112,N_12704,N_16926);
or U21113 (N_21113,N_15002,N_17410);
xor U21114 (N_21114,N_14588,N_16834);
and U21115 (N_21115,N_13313,N_13368);
or U21116 (N_21116,N_13929,N_15535);
or U21117 (N_21117,N_16598,N_14116);
nor U21118 (N_21118,N_15480,N_16048);
or U21119 (N_21119,N_16648,N_14323);
nand U21120 (N_21120,N_15279,N_13062);
nand U21121 (N_21121,N_17671,N_17663);
or U21122 (N_21122,N_13761,N_12888);
or U21123 (N_21123,N_15254,N_12512);
and U21124 (N_21124,N_15098,N_13180);
or U21125 (N_21125,N_13319,N_18616);
and U21126 (N_21126,N_15974,N_17969);
and U21127 (N_21127,N_13120,N_14037);
and U21128 (N_21128,N_17521,N_14737);
and U21129 (N_21129,N_13119,N_13126);
or U21130 (N_21130,N_16238,N_17944);
xor U21131 (N_21131,N_18242,N_15751);
xnor U21132 (N_21132,N_15973,N_15917);
nand U21133 (N_21133,N_17178,N_16961);
or U21134 (N_21134,N_13457,N_17503);
xnor U21135 (N_21135,N_12904,N_18088);
xnor U21136 (N_21136,N_14458,N_18311);
nor U21137 (N_21137,N_16803,N_18252);
nor U21138 (N_21138,N_14335,N_17707);
nand U21139 (N_21139,N_16981,N_18274);
and U21140 (N_21140,N_12883,N_14081);
or U21141 (N_21141,N_13088,N_12587);
nand U21142 (N_21142,N_16153,N_18466);
nand U21143 (N_21143,N_13106,N_16725);
nor U21144 (N_21144,N_17393,N_18354);
nand U21145 (N_21145,N_16591,N_17246);
or U21146 (N_21146,N_14951,N_13044);
and U21147 (N_21147,N_13844,N_13684);
or U21148 (N_21148,N_15373,N_18338);
or U21149 (N_21149,N_15871,N_13677);
xor U21150 (N_21150,N_16905,N_12782);
or U21151 (N_21151,N_16085,N_15190);
nor U21152 (N_21152,N_15193,N_14874);
xor U21153 (N_21153,N_14096,N_17894);
or U21154 (N_21154,N_18003,N_17833);
xnor U21155 (N_21155,N_17266,N_13229);
or U21156 (N_21156,N_18326,N_13637);
xnor U21157 (N_21157,N_13689,N_18524);
nor U21158 (N_21158,N_18230,N_13257);
xor U21159 (N_21159,N_14886,N_12946);
xor U21160 (N_21160,N_18296,N_13823);
xor U21161 (N_21161,N_17999,N_14735);
nor U21162 (N_21162,N_14754,N_14218);
nand U21163 (N_21163,N_17359,N_14334);
nor U21164 (N_21164,N_18733,N_14833);
or U21165 (N_21165,N_17327,N_14375);
nand U21166 (N_21166,N_16170,N_12676);
xnor U21167 (N_21167,N_17599,N_18033);
nand U21168 (N_21168,N_14759,N_18523);
nand U21169 (N_21169,N_12937,N_15819);
and U21170 (N_21170,N_16070,N_14739);
nand U21171 (N_21171,N_13604,N_13220);
and U21172 (N_21172,N_17856,N_17984);
nor U21173 (N_21173,N_18064,N_13995);
nand U21174 (N_21174,N_17708,N_17300);
and U21175 (N_21175,N_13036,N_13502);
xnor U21176 (N_21176,N_17651,N_13871);
or U21177 (N_21177,N_18579,N_17767);
or U21178 (N_21178,N_13448,N_17974);
nor U21179 (N_21179,N_17524,N_13370);
or U21180 (N_21180,N_17858,N_18439);
xnor U21181 (N_21181,N_17742,N_17762);
nand U21182 (N_21182,N_13192,N_15702);
nor U21183 (N_21183,N_15295,N_12502);
nand U21184 (N_21184,N_12573,N_18096);
nand U21185 (N_21185,N_12999,N_15851);
nor U21186 (N_21186,N_13338,N_18302);
nand U21187 (N_21187,N_14972,N_14967);
nand U21188 (N_21188,N_12841,N_15741);
or U21189 (N_21189,N_12611,N_12827);
nor U21190 (N_21190,N_18022,N_15374);
nor U21191 (N_21191,N_18119,N_18612);
and U21192 (N_21192,N_16619,N_18572);
xor U21193 (N_21193,N_16554,N_18331);
or U21194 (N_21194,N_15635,N_14223);
nor U21195 (N_21195,N_16267,N_13303);
xnor U21196 (N_21196,N_13477,N_17457);
nand U21197 (N_21197,N_15853,N_15226);
and U21198 (N_21198,N_15827,N_17696);
or U21199 (N_21199,N_18457,N_18673);
nor U21200 (N_21200,N_16684,N_16289);
xor U21201 (N_21201,N_16763,N_14452);
nor U21202 (N_21202,N_12948,N_18303);
nor U21203 (N_21203,N_14370,N_13456);
xnor U21204 (N_21204,N_16578,N_16582);
xnor U21205 (N_21205,N_13321,N_17997);
xor U21206 (N_21206,N_17363,N_18341);
nand U21207 (N_21207,N_17138,N_13146);
nor U21208 (N_21208,N_15129,N_14505);
xnor U21209 (N_21209,N_15329,N_18355);
or U21210 (N_21210,N_18314,N_17108);
nor U21211 (N_21211,N_15252,N_17546);
xnor U21212 (N_21212,N_12514,N_17085);
nand U21213 (N_21213,N_18639,N_16968);
or U21214 (N_21214,N_15693,N_17098);
or U21215 (N_21215,N_18651,N_15356);
and U21216 (N_21216,N_13902,N_14296);
nand U21217 (N_21217,N_18416,N_17215);
nor U21218 (N_21218,N_18093,N_16351);
or U21219 (N_21219,N_16134,N_12668);
nand U21220 (N_21220,N_16949,N_18550);
and U21221 (N_21221,N_17996,N_12919);
xnor U21222 (N_21222,N_14935,N_13968);
xor U21223 (N_21223,N_17196,N_17687);
nand U21224 (N_21224,N_12860,N_16295);
and U21225 (N_21225,N_16875,N_16086);
and U21226 (N_21226,N_14019,N_17427);
and U21227 (N_21227,N_12695,N_17684);
nor U21228 (N_21228,N_12972,N_15508);
or U21229 (N_21229,N_15140,N_14465);
nor U21230 (N_21230,N_13367,N_12513);
and U21231 (N_21231,N_17677,N_14986);
xor U21232 (N_21232,N_14237,N_13198);
or U21233 (N_21233,N_14981,N_13838);
and U21234 (N_21234,N_15797,N_17600);
nor U21235 (N_21235,N_18329,N_13236);
xor U21236 (N_21236,N_13811,N_12798);
and U21237 (N_21237,N_13596,N_12510);
nand U21238 (N_21238,N_14399,N_17501);
xor U21239 (N_21239,N_16976,N_18725);
nand U21240 (N_21240,N_14189,N_15683);
xnor U21241 (N_21241,N_14575,N_17048);
xnor U21242 (N_21242,N_13077,N_18512);
nor U21243 (N_21243,N_17244,N_18186);
or U21244 (N_21244,N_12886,N_12632);
or U21245 (N_21245,N_17576,N_17422);
xnor U21246 (N_21246,N_16270,N_16456);
nand U21247 (N_21247,N_17913,N_15496);
or U21248 (N_21248,N_18570,N_16214);
or U21249 (N_21249,N_18611,N_15434);
and U21250 (N_21250,N_16419,N_17087);
and U21251 (N_21251,N_15939,N_16992);
nor U21252 (N_21252,N_15806,N_17217);
nand U21253 (N_21253,N_14957,N_13645);
xor U21254 (N_21254,N_13280,N_16025);
nand U21255 (N_21255,N_16422,N_16581);
xnor U21256 (N_21256,N_13873,N_15008);
or U21257 (N_21257,N_15458,N_17824);
and U21258 (N_21258,N_12997,N_15981);
and U21259 (N_21259,N_14660,N_13539);
xnor U21260 (N_21260,N_14431,N_17613);
xor U21261 (N_21261,N_13935,N_15383);
and U21262 (N_21262,N_15179,N_14929);
nand U21263 (N_21263,N_16565,N_17836);
nor U21264 (N_21264,N_14127,N_12564);
xnor U21265 (N_21265,N_15774,N_13832);
or U21266 (N_21266,N_13029,N_14904);
nand U21267 (N_21267,N_18142,N_14921);
or U21268 (N_21268,N_16966,N_12831);
and U21269 (N_21269,N_18691,N_16371);
or U21270 (N_21270,N_13255,N_15782);
and U21271 (N_21271,N_13880,N_13482);
xor U21272 (N_21272,N_18055,N_12758);
and U21273 (N_21273,N_15503,N_17137);
or U21274 (N_21274,N_15320,N_13075);
or U21275 (N_21275,N_18684,N_13743);
nor U21276 (N_21276,N_13723,N_16429);
nand U21277 (N_21277,N_15775,N_17968);
nor U21278 (N_21278,N_18348,N_17113);
nand U21279 (N_21279,N_16692,N_14072);
xor U21280 (N_21280,N_12647,N_14306);
or U21281 (N_21281,N_13295,N_15103);
xor U21282 (N_21282,N_14056,N_17960);
nand U21283 (N_21283,N_14012,N_12956);
and U21284 (N_21284,N_14714,N_16997);
nor U21285 (N_21285,N_17184,N_14213);
and U21286 (N_21286,N_17766,N_14782);
xor U21287 (N_21287,N_17659,N_14696);
or U21288 (N_21288,N_15970,N_18723);
or U21289 (N_21289,N_16075,N_18102);
nand U21290 (N_21290,N_17740,N_17200);
xor U21291 (N_21291,N_18536,N_16008);
and U21292 (N_21292,N_14305,N_15044);
and U21293 (N_21293,N_18205,N_14020);
nand U21294 (N_21294,N_18454,N_18465);
nor U21295 (N_21295,N_17839,N_13189);
and U21296 (N_21296,N_16264,N_13624);
nand U21297 (N_21297,N_14219,N_16798);
xnor U21298 (N_21298,N_12760,N_18308);
nor U21299 (N_21299,N_16611,N_15872);
or U21300 (N_21300,N_16884,N_14558);
or U21301 (N_21301,N_13423,N_18434);
nor U21302 (N_21302,N_14121,N_16965);
nand U21303 (N_21303,N_17304,N_12871);
or U21304 (N_21304,N_15660,N_17133);
xnor U21305 (N_21305,N_15253,N_13841);
nor U21306 (N_21306,N_14107,N_15475);
or U21307 (N_21307,N_18662,N_17435);
or U21308 (N_21308,N_18461,N_13097);
nand U21309 (N_21309,N_16733,N_16023);
nor U21310 (N_21310,N_13510,N_16468);
nand U21311 (N_21311,N_15513,N_13987);
nor U21312 (N_21312,N_15166,N_18162);
nand U21313 (N_21313,N_14756,N_13263);
and U21314 (N_21314,N_14804,N_13059);
or U21315 (N_21315,N_17403,N_18335);
and U21316 (N_21316,N_16911,N_15532);
xor U21317 (N_21317,N_17690,N_17500);
and U21318 (N_21318,N_13573,N_14627);
and U21319 (N_21319,N_15386,N_17759);
nand U21320 (N_21320,N_16258,N_15677);
xnor U21321 (N_21321,N_17559,N_15967);
and U21322 (N_21322,N_15045,N_12697);
xor U21323 (N_21323,N_13020,N_18543);
nor U21324 (N_21324,N_16988,N_17401);
nand U21325 (N_21325,N_18358,N_17931);
nand U21326 (N_21326,N_14268,N_16553);
or U21327 (N_21327,N_15537,N_14102);
and U21328 (N_21328,N_16523,N_15908);
xnor U21329 (N_21329,N_17463,N_18041);
nor U21330 (N_21330,N_13437,N_16943);
xor U21331 (N_21331,N_15959,N_14385);
xor U21332 (N_21332,N_12777,N_16645);
nand U21333 (N_21333,N_14517,N_13517);
xor U21334 (N_21334,N_15319,N_15362);
or U21335 (N_21335,N_17536,N_14608);
xor U21336 (N_21336,N_15531,N_16642);
xnor U21337 (N_21337,N_13320,N_17911);
and U21338 (N_21338,N_15538,N_17479);
nand U21339 (N_21339,N_13238,N_14187);
nor U21340 (N_21340,N_14211,N_14757);
or U21341 (N_21341,N_13287,N_14064);
xor U21342 (N_21342,N_14943,N_17638);
nand U21343 (N_21343,N_16081,N_15258);
and U21344 (N_21344,N_17458,N_12696);
or U21345 (N_21345,N_16317,N_15564);
xnor U21346 (N_21346,N_17398,N_15928);
nor U21347 (N_21347,N_14815,N_14868);
nor U21348 (N_21348,N_13739,N_18077);
and U21349 (N_21349,N_14378,N_13162);
nor U21350 (N_21350,N_16693,N_14675);
nand U21351 (N_21351,N_13151,N_16663);
xor U21352 (N_21352,N_13007,N_16838);
and U21353 (N_21353,N_18260,N_14497);
xnor U21354 (N_21354,N_12744,N_15349);
nor U21355 (N_21355,N_16537,N_17454);
or U21356 (N_21356,N_14430,N_14705);
and U21357 (N_21357,N_12743,N_15874);
nor U21358 (N_21358,N_14544,N_13450);
or U21359 (N_21359,N_16037,N_17400);
nand U21360 (N_21360,N_16631,N_15309);
nor U21361 (N_21361,N_17148,N_12607);
and U21362 (N_21362,N_12795,N_18557);
nand U21363 (N_21363,N_17743,N_17298);
nand U21364 (N_21364,N_18561,N_15368);
nor U21365 (N_21365,N_15119,N_16182);
nor U21366 (N_21366,N_17544,N_16188);
or U21367 (N_21367,N_13354,N_13804);
and U21368 (N_21368,N_15126,N_14646);
xor U21369 (N_21369,N_14307,N_15754);
or U21370 (N_21370,N_18074,N_12729);
xnor U21371 (N_21371,N_17005,N_17307);
or U21372 (N_21372,N_16098,N_15396);
xnor U21373 (N_21373,N_16485,N_16398);
or U21374 (N_21374,N_18442,N_18376);
and U21375 (N_21375,N_13741,N_17614);
or U21376 (N_21376,N_17198,N_14606);
xnor U21377 (N_21377,N_12984,N_14035);
nand U21378 (N_21378,N_13350,N_17737);
xor U21379 (N_21379,N_14273,N_14192);
and U21380 (N_21380,N_18388,N_16408);
nor U21381 (N_21381,N_13049,N_15511);
or U21382 (N_21382,N_18044,N_16980);
or U21383 (N_21383,N_12706,N_13921);
and U21384 (N_21384,N_14286,N_17037);
xnor U21385 (N_21385,N_17523,N_17774);
xor U21386 (N_21386,N_15344,N_17253);
nand U21387 (N_21387,N_15057,N_14360);
or U21388 (N_21388,N_14048,N_15286);
and U21389 (N_21389,N_13005,N_13742);
or U21390 (N_21390,N_18551,N_15269);
nand U21391 (N_21391,N_13853,N_15868);
or U21392 (N_21392,N_18248,N_17812);
or U21393 (N_21393,N_14421,N_16396);
or U21394 (N_21394,N_14724,N_14557);
nand U21395 (N_21395,N_14825,N_16391);
and U21396 (N_21396,N_15763,N_15957);
or U21397 (N_21397,N_18468,N_13828);
nand U21398 (N_21398,N_16119,N_16654);
and U21399 (N_21399,N_17206,N_18286);
nor U21400 (N_21400,N_17237,N_14768);
nand U21401 (N_21401,N_14597,N_15756);
nor U21402 (N_21402,N_17873,N_17817);
or U21403 (N_21403,N_13500,N_15300);
and U21404 (N_21404,N_13892,N_13230);
nor U21405 (N_21405,N_16370,N_13073);
and U21406 (N_21406,N_15345,N_17409);
xor U21407 (N_21407,N_17682,N_14740);
nand U21408 (N_21408,N_17556,N_17845);
and U21409 (N_21409,N_17090,N_13306);
nand U21410 (N_21410,N_12885,N_14131);
and U21411 (N_21411,N_16302,N_18312);
nand U21412 (N_21412,N_13728,N_13124);
nand U21413 (N_21413,N_14834,N_18293);
and U21414 (N_21414,N_16067,N_16179);
nand U21415 (N_21415,N_13091,N_17499);
or U21416 (N_21416,N_17610,N_16363);
or U21417 (N_21417,N_18740,N_17170);
nand U21418 (N_21418,N_17646,N_15855);
nand U21419 (N_21419,N_12621,N_17383);
nor U21420 (N_21420,N_17871,N_13017);
or U21421 (N_21421,N_15263,N_14401);
nand U21422 (N_21422,N_12865,N_17233);
nand U21423 (N_21423,N_15051,N_18689);
xor U21424 (N_21424,N_18401,N_15164);
nor U21425 (N_21425,N_13489,N_14209);
and U21426 (N_21426,N_18075,N_15789);
or U21427 (N_21427,N_18146,N_13574);
or U21428 (N_21428,N_13312,N_18222);
or U21429 (N_21429,N_17819,N_13409);
nor U21430 (N_21430,N_15323,N_16375);
nor U21431 (N_21431,N_12507,N_12850);
and U21432 (N_21432,N_18571,N_14907);
or U21433 (N_21433,N_15631,N_14382);
xor U21434 (N_21434,N_17344,N_16691);
nand U21435 (N_21435,N_15343,N_14222);
nand U21436 (N_21436,N_14144,N_15884);
or U21437 (N_21437,N_13415,N_13392);
or U21438 (N_21438,N_18735,N_16242);
and U21439 (N_21439,N_13927,N_17719);
and U21440 (N_21440,N_16664,N_16671);
xnor U21441 (N_21441,N_17078,N_15472);
and U21442 (N_21442,N_13399,N_12940);
and U21443 (N_21443,N_13254,N_14356);
nand U21444 (N_21444,N_14924,N_16589);
nand U21445 (N_21445,N_13224,N_13779);
and U21446 (N_21446,N_17257,N_16114);
and U21447 (N_21447,N_18187,N_14486);
or U21448 (N_21448,N_13215,N_18474);
and U21449 (N_21449,N_17156,N_16630);
and U21450 (N_21450,N_16699,N_14516);
xor U21451 (N_21451,N_13282,N_14007);
xnor U21452 (N_21452,N_13305,N_18451);
nor U21453 (N_21453,N_16423,N_17242);
nand U21454 (N_21454,N_13983,N_12509);
nand U21455 (N_21455,N_15303,N_16206);
nand U21456 (N_21456,N_18112,N_13102);
nor U21457 (N_21457,N_17021,N_17017);
nand U21458 (N_21458,N_15586,N_15745);
nor U21459 (N_21459,N_18706,N_12608);
nand U21460 (N_21460,N_17308,N_15366);
nand U21461 (N_21461,N_17461,N_16054);
or U21462 (N_21462,N_13726,N_14000);
or U21463 (N_21463,N_16090,N_16715);
nor U21464 (N_21464,N_16035,N_13803);
nand U21465 (N_21465,N_16162,N_16964);
or U21466 (N_21466,N_17872,N_16133);
xor U21467 (N_21467,N_16222,N_15259);
nand U21468 (N_21468,N_14966,N_15062);
nor U21469 (N_21469,N_18188,N_16494);
nand U21470 (N_21470,N_15720,N_13030);
nand U21471 (N_21471,N_17041,N_17185);
and U21472 (N_21472,N_18206,N_16812);
nand U21473 (N_21473,N_15764,N_16481);
xnor U21474 (N_21474,N_13937,N_14051);
xor U21475 (N_21475,N_13487,N_13994);
nand U21476 (N_21476,N_16344,N_13184);
and U21477 (N_21477,N_17480,N_17975);
nor U21478 (N_21478,N_12641,N_15744);
or U21479 (N_21479,N_18203,N_15519);
or U21480 (N_21480,N_14600,N_18544);
or U21481 (N_21481,N_15342,N_14952);
nand U21482 (N_21482,N_18135,N_15358);
or U21483 (N_21483,N_17641,N_16412);
xor U21484 (N_21484,N_16057,N_13125);
or U21485 (N_21485,N_15124,N_14478);
nand U21486 (N_21486,N_13441,N_18063);
nand U21487 (N_21487,N_16309,N_12916);
nand U21488 (N_21488,N_18285,N_15056);
or U21489 (N_21489,N_13735,N_18517);
or U21490 (N_21490,N_18160,N_16842);
nand U21491 (N_21491,N_17789,N_16369);
xor U21492 (N_21492,N_18425,N_18315);
nor U21493 (N_21493,N_16694,N_15429);
or U21494 (N_21494,N_14284,N_17542);
xor U21495 (N_21495,N_18368,N_17040);
nor U21496 (N_21496,N_15459,N_18480);
and U21497 (N_21497,N_18580,N_16413);
nor U21498 (N_21498,N_17993,N_16552);
xnor U21499 (N_21499,N_17371,N_18390);
nand U21500 (N_21500,N_16563,N_18594);
and U21501 (N_21501,N_14389,N_16490);
nand U21502 (N_21502,N_15453,N_16784);
or U21503 (N_21503,N_18172,N_15505);
nor U21504 (N_21504,N_15090,N_18140);
or U21505 (N_21505,N_15083,N_16933);
nand U21506 (N_21506,N_15835,N_15875);
nand U21507 (N_21507,N_16152,N_17019);
and U21508 (N_21508,N_16212,N_15515);
xnor U21509 (N_21509,N_17261,N_13344);
and U21510 (N_21510,N_14612,N_18393);
and U21511 (N_21511,N_18226,N_16670);
or U21512 (N_21512,N_18065,N_16240);
or U21513 (N_21513,N_14745,N_14288);
or U21514 (N_21514,N_13428,N_12665);
nor U21515 (N_21515,N_13800,N_17116);
or U21516 (N_21516,N_18339,N_18412);
and U21517 (N_21517,N_13085,N_13568);
and U21518 (N_21518,N_16194,N_14788);
nand U21519 (N_21519,N_15251,N_14819);
or U21520 (N_21520,N_13535,N_17780);
and U21521 (N_21521,N_18494,N_16649);
and U21522 (N_21522,N_17149,N_15892);
or U21523 (N_21523,N_13407,N_16087);
and U21524 (N_21524,N_17822,N_16280);
nor U21525 (N_21525,N_17914,N_18554);
and U21526 (N_21526,N_16308,N_12818);
xor U21527 (N_21527,N_14515,N_13660);
xnor U21528 (N_21528,N_15695,N_15448);
or U21529 (N_21529,N_17413,N_16571);
nand U21530 (N_21530,N_15913,N_17758);
and U21531 (N_21531,N_15091,N_13142);
or U21532 (N_21532,N_13727,N_13656);
xnor U21533 (N_21533,N_15247,N_16028);
nand U21534 (N_21534,N_13807,N_13212);
nand U21535 (N_21535,N_16979,N_17272);
nand U21536 (N_21536,N_14153,N_15843);
xor U21537 (N_21537,N_16360,N_14969);
xnor U21538 (N_21538,N_13643,N_17252);
nand U21539 (N_21539,N_12576,N_14247);
xor U21540 (N_21540,N_13796,N_18211);
xnor U21541 (N_21541,N_18559,N_15852);
xor U21542 (N_21542,N_14439,N_14807);
nand U21543 (N_21543,N_15233,N_12755);
nand U21544 (N_21544,N_16097,N_15492);
and U21545 (N_21545,N_18031,N_17896);
or U21546 (N_21546,N_13632,N_16624);
and U21547 (N_21547,N_14522,N_17173);
xor U21548 (N_21548,N_14488,N_18532);
and U21549 (N_21549,N_14493,N_17652);
nand U21550 (N_21550,N_13606,N_14067);
xnor U21551 (N_21551,N_14440,N_14021);
and U21552 (N_21552,N_17318,N_13166);
and U21553 (N_21553,N_14970,N_13979);
nand U21554 (N_21554,N_13608,N_14145);
nand U21555 (N_21555,N_17583,N_16629);
xnor U21556 (N_21556,N_15812,N_15284);
and U21557 (N_21557,N_13226,N_16275);
xor U21558 (N_21558,N_17142,N_13382);
xor U21559 (N_21559,N_13486,N_15211);
nor U21560 (N_21560,N_13115,N_14514);
nor U21561 (N_21561,N_15823,N_17666);
nor U21562 (N_21562,N_18233,N_12792);
and U21563 (N_21563,N_18565,N_15063);
and U21564 (N_21564,N_18389,N_17785);
xnor U21565 (N_21565,N_15203,N_18051);
nand U21566 (N_21566,N_18108,N_13076);
nand U21567 (N_21567,N_14032,N_15662);
and U21568 (N_21568,N_12820,N_15022);
nor U21569 (N_21569,N_15005,N_14298);
nand U21570 (N_21570,N_12974,N_16752);
xor U21571 (N_21571,N_15712,N_17518);
nor U21572 (N_21572,N_15808,N_16756);
or U21573 (N_21573,N_17262,N_16708);
nand U21574 (N_21574,N_17167,N_16915);
and U21575 (N_21575,N_18244,N_13432);
nand U21576 (N_21576,N_15427,N_13385);
xnor U21577 (N_21577,N_12551,N_16331);
and U21578 (N_21578,N_15125,N_15367);
or U21579 (N_21579,N_15009,N_16530);
and U21580 (N_21580,N_18659,N_18692);
and U21581 (N_21581,N_15111,N_16055);
and U21582 (N_21582,N_16636,N_15992);
or U21583 (N_21583,N_16555,N_18405);
nor U21584 (N_21584,N_17963,N_14913);
xor U21585 (N_21585,N_16735,N_17866);
nand U21586 (N_21586,N_17052,N_16505);
xor U21587 (N_21587,N_17854,N_14508);
nand U21588 (N_21588,N_16337,N_12779);
xor U21589 (N_21589,N_13738,N_15608);
xnor U21590 (N_21590,N_17077,N_14603);
and U21591 (N_21591,N_16574,N_16435);
nor U21592 (N_21592,N_14859,N_16525);
nand U21593 (N_21593,N_13307,N_17103);
xor U21594 (N_21594,N_15389,N_15831);
or U21595 (N_21595,N_13218,N_12769);
nand U21596 (N_21596,N_16579,N_13628);
nor U21597 (N_21597,N_16056,N_15121);
nand U21598 (N_21598,N_15829,N_15272);
nor U21599 (N_21599,N_16940,N_15619);
nor U21600 (N_21600,N_15864,N_13374);
or U21601 (N_21601,N_17450,N_14681);
xnor U21602 (N_21602,N_13449,N_18590);
xor U21603 (N_21603,N_13410,N_14910);
nand U21604 (N_21604,N_15947,N_16010);
xnor U21605 (N_21605,N_16700,N_16560);
nand U21606 (N_21606,N_13938,N_18513);
and U21607 (N_21607,N_12673,N_17032);
nand U21608 (N_21608,N_14490,N_13132);
nor U21609 (N_21609,N_16753,N_17063);
nor U21610 (N_21610,N_15795,N_18352);
nor U21611 (N_21611,N_13846,N_16906);
nor U21612 (N_21612,N_16639,N_13962);
and U21613 (N_21613,N_17553,N_12581);
xor U21614 (N_21614,N_17247,N_17270);
xnor U21615 (N_21615,N_13916,N_17967);
and U21616 (N_21616,N_18080,N_13925);
and U21617 (N_21617,N_15192,N_15570);
nor U21618 (N_21618,N_17992,N_14498);
and U21619 (N_21619,N_12520,N_16288);
and U21620 (N_21620,N_17310,N_18500);
or U21621 (N_21621,N_13444,N_17276);
xnor U21622 (N_21622,N_18424,N_16804);
nand U21623 (N_21623,N_12664,N_14477);
xnor U21624 (N_21624,N_14755,N_14732);
nor U21625 (N_21625,N_17123,N_18196);
nor U21626 (N_21626,N_17645,N_16547);
and U21627 (N_21627,N_17915,N_13143);
nand U21628 (N_21628,N_16596,N_17194);
nand U21629 (N_21629,N_14741,N_18104);
or U21630 (N_21630,N_17045,N_17977);
or U21631 (N_21631,N_16444,N_15783);
nand U21632 (N_21632,N_15881,N_16781);
or U21633 (N_21633,N_18467,N_12771);
nand U21634 (N_21634,N_16336,N_16584);
nor U21635 (N_21635,N_17867,N_16477);
nand U21636 (N_21636,N_14541,N_17892);
xor U21637 (N_21637,N_14933,N_16156);
and U21638 (N_21638,N_17857,N_13290);
nand U21639 (N_21639,N_18261,N_17640);
or U21640 (N_21640,N_15945,N_12819);
or U21641 (N_21641,N_13056,N_13021);
or U21642 (N_21642,N_17924,N_17147);
or U21643 (N_21643,N_16296,N_15870);
nand U21644 (N_21644,N_17874,N_16809);
nand U21645 (N_21645,N_14071,N_12914);
xnor U21646 (N_21646,N_15058,N_17761);
xnor U21647 (N_21647,N_17058,N_16430);
and U21648 (N_21648,N_17095,N_13518);
nor U21649 (N_21649,N_14936,N_17118);
nor U21650 (N_21650,N_17225,N_14985);
nand U21651 (N_21651,N_16053,N_16385);
nand U21652 (N_21652,N_15463,N_18255);
or U21653 (N_21653,N_14113,N_12570);
nor U21654 (N_21654,N_18321,N_15613);
xnor U21655 (N_21655,N_13003,N_12978);
xor U21656 (N_21656,N_14070,N_17001);
nor U21657 (N_21657,N_14331,N_17940);
nand U21658 (N_21658,N_15393,N_16769);
and U21659 (N_21659,N_12924,N_18069);
nand U21660 (N_21660,N_17849,N_13341);
xnor U21661 (N_21661,N_13636,N_16775);
nand U21662 (N_21662,N_16576,N_15011);
xor U21663 (N_21663,N_14400,N_15971);
xnor U21664 (N_21664,N_15542,N_12840);
or U21665 (N_21665,N_15020,N_16822);
nand U21666 (N_21666,N_14270,N_13340);
nor U21667 (N_21667,N_14263,N_12966);
and U21668 (N_21668,N_14797,N_17370);
xor U21669 (N_21669,N_15447,N_17239);
nand U21670 (N_21670,N_16519,N_16878);
nor U21671 (N_21671,N_15291,N_15361);
or U21672 (N_21672,N_18059,N_14109);
xnor U21673 (N_21673,N_18229,N_14838);
nand U21674 (N_21674,N_16953,N_17612);
nand U21675 (N_21675,N_14427,N_15431);
nand U21676 (N_21676,N_17119,N_15130);
nor U21677 (N_21677,N_18225,N_14412);
xnor U21678 (N_21678,N_18232,N_13977);
nand U21679 (N_21679,N_15477,N_17972);
and U21680 (N_21680,N_13058,N_14194);
xor U21681 (N_21681,N_18183,N_14778);
and U21682 (N_21682,N_17888,N_16815);
xnor U21683 (N_21683,N_12780,N_17688);
and U21684 (N_21684,N_13737,N_17258);
nor U21685 (N_21685,N_14068,N_15679);
nand U21686 (N_21686,N_14085,N_16482);
xnor U21687 (N_21687,N_12716,N_16463);
and U21688 (N_21688,N_15066,N_17834);
and U21689 (N_21689,N_13897,N_17796);
nand U21690 (N_21690,N_14402,N_15729);
nor U21691 (N_21691,N_17392,N_14561);
nand U21692 (N_21692,N_15728,N_16021);
and U21693 (N_21693,N_13554,N_16169);
nand U21694 (N_21694,N_16546,N_14770);
xor U21695 (N_21695,N_14372,N_16614);
xnor U21696 (N_21696,N_15778,N_15801);
nand U21697 (N_21697,N_13891,N_14472);
nor U21698 (N_21698,N_18086,N_13147);
nor U21699 (N_21699,N_16137,N_13013);
xor U21700 (N_21700,N_14786,N_12663);
or U21701 (N_21701,N_17961,N_13511);
or U21702 (N_21702,N_13513,N_18359);
nand U21703 (N_21703,N_14509,N_14500);
and U21704 (N_21704,N_15325,N_18251);
nor U21705 (N_21705,N_13008,N_15612);
nor U21706 (N_21706,N_14641,N_12511);
nor U21707 (N_21707,N_12657,N_13329);
nor U21708 (N_21708,N_13206,N_16874);
xnor U21709 (N_21709,N_18620,N_17810);
nand U21710 (N_21710,N_16899,N_13098);
xnor U21711 (N_21711,N_15293,N_15333);
or U21712 (N_21712,N_15690,N_12951);
and U21713 (N_21713,N_13659,N_16350);
or U21714 (N_21714,N_15979,N_14632);
or U21715 (N_21715,N_15445,N_14437);
nor U21716 (N_21716,N_16233,N_12731);
and U21717 (N_21717,N_13829,N_14881);
nand U21718 (N_21718,N_16154,N_13567);
or U21719 (N_21719,N_16411,N_18646);
xnor U21720 (N_21720,N_13266,N_17349);
xnor U21721 (N_21721,N_13388,N_15017);
xnor U21722 (N_21722,N_16773,N_13474);
nand U21723 (N_21723,N_17082,N_13247);
or U21724 (N_21724,N_17428,N_16439);
and U21725 (N_21725,N_12750,N_16249);
nand U21726 (N_21726,N_17580,N_12787);
or U21727 (N_21727,N_14502,N_14727);
xnor U21728 (N_21728,N_18087,N_17219);
xnor U21729 (N_21729,N_13134,N_14058);
nor U21730 (N_21730,N_14428,N_14386);
and U21731 (N_21731,N_17592,N_14246);
and U21732 (N_21732,N_18082,N_16215);
xor U21733 (N_21733,N_16658,N_14862);
nand U21734 (N_21734,N_16227,N_17529);
or U21735 (N_21735,N_18168,N_14538);
or U21736 (N_21736,N_18223,N_14864);
and U21737 (N_21737,N_14980,N_14893);
nand U21738 (N_21738,N_15070,N_15791);
xor U21739 (N_21739,N_18283,N_15353);
nor U21740 (N_21740,N_16506,N_17060);
or U21741 (N_21741,N_18392,N_18079);
nand U21742 (N_21742,N_14339,N_17818);
nor U21743 (N_21743,N_13400,N_18718);
or U21744 (N_21744,N_18458,N_17358);
or U21745 (N_21745,N_15398,N_17020);
nor U21746 (N_21746,N_14586,N_13495);
xor U21747 (N_21747,N_13696,N_12639);
and U21748 (N_21748,N_14796,N_14695);
or U21749 (N_21749,N_15372,N_14553);
nand U21750 (N_21750,N_17313,N_18588);
nand U21751 (N_21751,N_13789,N_17139);
xor U21752 (N_21752,N_18030,N_17482);
nor U21753 (N_21753,N_14380,N_15627);
xor U21754 (N_21754,N_15442,N_12727);
or U21755 (N_21755,N_15297,N_17437);
or U21756 (N_21756,N_14225,N_18548);
xor U21757 (N_21757,N_14916,N_14767);
or U21758 (N_21758,N_14931,N_14052);
nand U21759 (N_21759,N_16729,N_13946);
nor U21760 (N_21760,N_18549,N_15940);
nand U21761 (N_21761,N_13580,N_15382);
nor U21762 (N_21762,N_13471,N_13084);
nor U21763 (N_21763,N_16474,N_13705);
and U21764 (N_21764,N_13239,N_18361);
and U21765 (N_21765,N_14620,N_13150);
nor U21766 (N_21766,N_18443,N_18034);
or U21767 (N_21767,N_14562,N_15845);
or U21768 (N_21768,N_13260,N_16744);
or U21769 (N_21769,N_15825,N_15545);
and U21770 (N_21770,N_15194,N_12614);
nand U21771 (N_21771,N_14260,N_14424);
nand U21772 (N_21772,N_18336,N_13952);
nor U21773 (N_21773,N_13674,N_18110);
nand U21774 (N_21774,N_13686,N_16741);
and U21775 (N_21775,N_14357,N_17916);
nand U21776 (N_21776,N_18301,N_12998);
or U21777 (N_21777,N_18613,N_13243);
and U21778 (N_21778,N_14683,N_13022);
nand U21779 (N_21779,N_18240,N_17443);
nor U21780 (N_21780,N_16541,N_17773);
and U21781 (N_21781,N_18175,N_15311);
nand U21782 (N_21782,N_14022,N_13961);
or U21783 (N_21783,N_17970,N_12709);
and U21784 (N_21784,N_18325,N_13179);
xnor U21785 (N_21785,N_14944,N_17387);
xor U21786 (N_21786,N_14526,N_18103);
xor U21787 (N_21787,N_14892,N_18463);
nor U21788 (N_21788,N_17059,N_18529);
nand U21789 (N_21789,N_15762,N_14774);
nor U21790 (N_21790,N_14663,N_17702);
xor U21791 (N_21791,N_17860,N_13369);
nand U21792 (N_21792,N_15138,N_16738);
nor U21793 (N_21793,N_13376,N_16022);
or U21794 (N_21794,N_13033,N_12532);
xor U21795 (N_21795,N_14801,N_13694);
or U21796 (N_21796,N_15514,N_13945);
xor U21797 (N_21797,N_14445,N_18136);
and U21798 (N_21798,N_14216,N_12717);
xor U21799 (N_21799,N_16500,N_14536);
and U21800 (N_21800,N_15224,N_15776);
nor U21801 (N_21801,N_18603,N_12942);
or U21802 (N_21802,N_18645,N_15862);
nand U21803 (N_21803,N_15527,N_16083);
xor U21804 (N_21804,N_14760,N_14823);
xnor U21805 (N_21805,N_15710,N_14438);
nor U21806 (N_21806,N_14266,N_17808);
nand U21807 (N_21807,N_15059,N_15803);
xor U21808 (N_21808,N_18227,N_18387);
or U21809 (N_21809,N_16868,N_14783);
xor U21810 (N_21810,N_17506,N_15964);
nor U21811 (N_21811,N_18647,N_15410);
nand U21812 (N_21812,N_18644,N_14280);
or U21813 (N_21813,N_18333,N_17739);
xnor U21814 (N_21814,N_18062,N_17746);
and U21815 (N_21815,N_16610,N_14512);
xor U21816 (N_21816,N_14667,N_18537);
and U21817 (N_21817,N_15168,N_16676);
nand U21818 (N_21818,N_17382,N_18143);
nor U21819 (N_21819,N_15486,N_13619);
xor U21820 (N_21820,N_18495,N_17949);
nor U21821 (N_21821,N_18583,N_13731);
xor U21822 (N_21822,N_18239,N_17930);
nor U21823 (N_21823,N_12533,N_16279);
nand U21824 (N_21824,N_16544,N_18734);
nand U21825 (N_21825,N_18158,N_12688);
and U21826 (N_21826,N_14466,N_13911);
nand U21827 (N_21827,N_13364,N_14011);
and U21828 (N_21828,N_14079,N_13501);
or U21829 (N_21829,N_16318,N_18290);
nand U21830 (N_21830,N_18084,N_13706);
nor U21831 (N_21831,N_16329,N_16531);
and U21832 (N_21832,N_13121,N_18727);
nor U21833 (N_21833,N_12544,N_17485);
and U21834 (N_21834,N_18200,N_14202);
and U21835 (N_21835,N_17160,N_13585);
and U21836 (N_21836,N_16927,N_16567);
and U21837 (N_21837,N_17000,N_16356);
and U21838 (N_21838,N_14282,N_15172);
nand U21839 (N_21839,N_13046,N_16449);
and U21840 (N_21840,N_17012,N_14416);
nand U21841 (N_21841,N_17293,N_12585);
xor U21842 (N_21842,N_16845,N_17124);
nand U21843 (N_21843,N_13646,N_16069);
nand U21844 (N_21844,N_15064,N_14528);
nand U21845 (N_21845,N_13331,N_18531);
nand U21846 (N_21846,N_15040,N_16116);
and U21847 (N_21847,N_14842,N_14839);
and U21848 (N_21848,N_14320,N_15927);
or U21849 (N_21849,N_16450,N_12527);
or U21850 (N_21850,N_16780,N_17122);
nor U21851 (N_21851,N_15721,N_17130);
nor U21852 (N_21852,N_17504,N_15569);
xnor U21853 (N_21853,N_16628,N_16790);
nand U21854 (N_21854,N_12982,N_18406);
and U21855 (N_21855,N_14433,N_18399);
and U21856 (N_21856,N_16710,N_17245);
xnor U21857 (N_21857,N_14315,N_18682);
nor U21858 (N_21858,N_15281,N_14191);
or U21859 (N_21859,N_15276,N_17325);
nor U21860 (N_21860,N_14095,N_18180);
and U21861 (N_21861,N_16111,N_18440);
and U21862 (N_21862,N_13177,N_17372);
or U21863 (N_21863,N_17399,N_16644);
and U21864 (N_21864,N_15770,N_17227);
xor U21865 (N_21865,N_18370,N_17380);
and U21866 (N_21866,N_15768,N_13461);
nand U21867 (N_21867,N_18097,N_18020);
or U21868 (N_21868,N_16810,N_17279);
xnor U21869 (N_21869,N_15471,N_13122);
and U21870 (N_21870,N_13954,N_16458);
and U21871 (N_21871,N_15114,N_15428);
nand U21872 (N_21872,N_14984,N_17034);
or U21873 (N_21873,N_14275,N_18372);
nand U21874 (N_21874,N_17070,N_14110);
xnor U21875 (N_21875,N_15553,N_18331);
xor U21876 (N_21876,N_18263,N_13495);
xor U21877 (N_21877,N_12847,N_13503);
or U21878 (N_21878,N_15085,N_15524);
xnor U21879 (N_21879,N_16831,N_14599);
or U21880 (N_21880,N_12543,N_16200);
nand U21881 (N_21881,N_14605,N_14659);
or U21882 (N_21882,N_18597,N_16640);
nand U21883 (N_21883,N_17535,N_18335);
and U21884 (N_21884,N_18168,N_14224);
xor U21885 (N_21885,N_13659,N_15301);
or U21886 (N_21886,N_18492,N_14772);
xnor U21887 (N_21887,N_18466,N_15297);
or U21888 (N_21888,N_13151,N_14532);
and U21889 (N_21889,N_15752,N_14183);
nand U21890 (N_21890,N_14228,N_17420);
and U21891 (N_21891,N_13373,N_17947);
nor U21892 (N_21892,N_17201,N_14478);
xnor U21893 (N_21893,N_14662,N_15880);
xor U21894 (N_21894,N_18015,N_17649);
or U21895 (N_21895,N_18368,N_18524);
nor U21896 (N_21896,N_13500,N_15606);
xnor U21897 (N_21897,N_12951,N_17955);
nor U21898 (N_21898,N_16114,N_15418);
nand U21899 (N_21899,N_13036,N_15679);
xor U21900 (N_21900,N_17147,N_16491);
and U21901 (N_21901,N_17043,N_16745);
nand U21902 (N_21902,N_17697,N_17939);
nand U21903 (N_21903,N_13365,N_17399);
nor U21904 (N_21904,N_16072,N_12710);
nand U21905 (N_21905,N_13315,N_18487);
or U21906 (N_21906,N_16783,N_18466);
or U21907 (N_21907,N_17357,N_15200);
and U21908 (N_21908,N_12908,N_14353);
nand U21909 (N_21909,N_15519,N_16096);
or U21910 (N_21910,N_13470,N_17022);
nand U21911 (N_21911,N_13257,N_14296);
xnor U21912 (N_21912,N_15485,N_14783);
nor U21913 (N_21913,N_14730,N_16857);
nand U21914 (N_21914,N_13041,N_13214);
or U21915 (N_21915,N_14781,N_12641);
or U21916 (N_21916,N_18157,N_12611);
nor U21917 (N_21917,N_13026,N_14031);
nand U21918 (N_21918,N_12579,N_18631);
nand U21919 (N_21919,N_14422,N_18234);
nor U21920 (N_21920,N_14133,N_13717);
or U21921 (N_21921,N_17611,N_17280);
nor U21922 (N_21922,N_15172,N_12727);
nor U21923 (N_21923,N_13208,N_16417);
or U21924 (N_21924,N_16809,N_12730);
and U21925 (N_21925,N_13512,N_17347);
xor U21926 (N_21926,N_12989,N_18073);
or U21927 (N_21927,N_15418,N_15095);
xnor U21928 (N_21928,N_13143,N_12525);
nand U21929 (N_21929,N_13640,N_16440);
nor U21930 (N_21930,N_16394,N_15212);
nand U21931 (N_21931,N_17611,N_18580);
nand U21932 (N_21932,N_12727,N_14660);
or U21933 (N_21933,N_13159,N_13064);
nor U21934 (N_21934,N_17999,N_16462);
or U21935 (N_21935,N_18248,N_14978);
or U21936 (N_21936,N_16809,N_16072);
nor U21937 (N_21937,N_13247,N_17022);
and U21938 (N_21938,N_15883,N_13538);
nand U21939 (N_21939,N_13836,N_16674);
nand U21940 (N_21940,N_17352,N_15704);
nor U21941 (N_21941,N_17159,N_17119);
and U21942 (N_21942,N_15681,N_13850);
xor U21943 (N_21943,N_14516,N_13408);
nor U21944 (N_21944,N_17098,N_13165);
nor U21945 (N_21945,N_17296,N_13499);
nor U21946 (N_21946,N_14893,N_15945);
or U21947 (N_21947,N_12917,N_14275);
and U21948 (N_21948,N_18641,N_15299);
and U21949 (N_21949,N_13218,N_12822);
nand U21950 (N_21950,N_17841,N_18067);
nor U21951 (N_21951,N_12769,N_13219);
or U21952 (N_21952,N_17273,N_13941);
or U21953 (N_21953,N_13022,N_15875);
xor U21954 (N_21954,N_15797,N_18115);
and U21955 (N_21955,N_13436,N_17507);
or U21956 (N_21956,N_13857,N_16494);
xor U21957 (N_21957,N_16437,N_13910);
xor U21958 (N_21958,N_16923,N_18207);
xor U21959 (N_21959,N_16335,N_16303);
nand U21960 (N_21960,N_15836,N_13358);
or U21961 (N_21961,N_14310,N_12582);
and U21962 (N_21962,N_14507,N_18342);
nand U21963 (N_21963,N_17922,N_15528);
nand U21964 (N_21964,N_13685,N_16732);
or U21965 (N_21965,N_12860,N_17114);
xnor U21966 (N_21966,N_16694,N_17899);
and U21967 (N_21967,N_14819,N_15438);
xnor U21968 (N_21968,N_14984,N_17144);
nand U21969 (N_21969,N_15073,N_12929);
xnor U21970 (N_21970,N_14046,N_15006);
nand U21971 (N_21971,N_14439,N_13409);
xor U21972 (N_21972,N_14282,N_16970);
xnor U21973 (N_21973,N_16288,N_15396);
and U21974 (N_21974,N_13386,N_12968);
nand U21975 (N_21975,N_16408,N_16330);
nand U21976 (N_21976,N_17728,N_15452);
nand U21977 (N_21977,N_17887,N_17745);
nand U21978 (N_21978,N_18548,N_14051);
and U21979 (N_21979,N_17060,N_17723);
and U21980 (N_21980,N_16334,N_13814);
and U21981 (N_21981,N_16560,N_16083);
nand U21982 (N_21982,N_14056,N_14826);
nand U21983 (N_21983,N_14305,N_15333);
xor U21984 (N_21984,N_18339,N_17793);
xnor U21985 (N_21985,N_14743,N_16380);
nor U21986 (N_21986,N_18569,N_15306);
nand U21987 (N_21987,N_16082,N_18537);
or U21988 (N_21988,N_14395,N_16375);
and U21989 (N_21989,N_14350,N_16323);
nor U21990 (N_21990,N_16804,N_15461);
or U21991 (N_21991,N_13583,N_17295);
nand U21992 (N_21992,N_14984,N_18089);
or U21993 (N_21993,N_13374,N_15396);
nor U21994 (N_21994,N_15627,N_17832);
nor U21995 (N_21995,N_17671,N_17356);
nand U21996 (N_21996,N_14567,N_14396);
or U21997 (N_21997,N_18219,N_13694);
nand U21998 (N_21998,N_13577,N_18548);
xnor U21999 (N_21999,N_15112,N_16742);
nor U22000 (N_22000,N_14379,N_18206);
xnor U22001 (N_22001,N_17682,N_15615);
nor U22002 (N_22002,N_14067,N_13582);
nand U22003 (N_22003,N_17376,N_14602);
nor U22004 (N_22004,N_18137,N_15810);
xnor U22005 (N_22005,N_16857,N_13396);
nand U22006 (N_22006,N_12964,N_14431);
or U22007 (N_22007,N_14641,N_13271);
nor U22008 (N_22008,N_12715,N_17599);
xor U22009 (N_22009,N_17138,N_18714);
xnor U22010 (N_22010,N_16241,N_12964);
or U22011 (N_22011,N_14958,N_13096);
and U22012 (N_22012,N_18139,N_14538);
xor U22013 (N_22013,N_16875,N_17512);
or U22014 (N_22014,N_18707,N_16953);
and U22015 (N_22015,N_15137,N_18150);
xor U22016 (N_22016,N_15639,N_14608);
and U22017 (N_22017,N_16559,N_15244);
xnor U22018 (N_22018,N_15701,N_14722);
and U22019 (N_22019,N_13887,N_14527);
and U22020 (N_22020,N_13715,N_12604);
nor U22021 (N_22021,N_16103,N_17465);
nor U22022 (N_22022,N_16872,N_16935);
xor U22023 (N_22023,N_12611,N_13781);
or U22024 (N_22024,N_14883,N_16898);
xor U22025 (N_22025,N_13231,N_15542);
nor U22026 (N_22026,N_16520,N_16764);
nor U22027 (N_22027,N_14647,N_15682);
xor U22028 (N_22028,N_15861,N_12573);
xnor U22029 (N_22029,N_17528,N_13567);
and U22030 (N_22030,N_14291,N_12682);
xor U22031 (N_22031,N_18319,N_13126);
nand U22032 (N_22032,N_17758,N_16367);
or U22033 (N_22033,N_14699,N_18675);
or U22034 (N_22034,N_13699,N_15343);
nand U22035 (N_22035,N_14262,N_15873);
nand U22036 (N_22036,N_14343,N_17695);
or U22037 (N_22037,N_12737,N_17539);
xnor U22038 (N_22038,N_18194,N_17312);
and U22039 (N_22039,N_15030,N_16135);
or U22040 (N_22040,N_13830,N_16750);
nand U22041 (N_22041,N_12709,N_14377);
and U22042 (N_22042,N_17055,N_18335);
nand U22043 (N_22043,N_15345,N_17711);
nand U22044 (N_22044,N_17568,N_13920);
or U22045 (N_22045,N_14446,N_17329);
xor U22046 (N_22046,N_14260,N_15553);
or U22047 (N_22047,N_12718,N_17353);
nand U22048 (N_22048,N_17339,N_14819);
nand U22049 (N_22049,N_18649,N_18416);
and U22050 (N_22050,N_18087,N_16281);
and U22051 (N_22051,N_14971,N_16877);
and U22052 (N_22052,N_16525,N_15598);
xor U22053 (N_22053,N_16586,N_12650);
or U22054 (N_22054,N_17062,N_14399);
nand U22055 (N_22055,N_16595,N_13173);
nand U22056 (N_22056,N_17436,N_14160);
and U22057 (N_22057,N_16687,N_14500);
nand U22058 (N_22058,N_15857,N_17102);
xnor U22059 (N_22059,N_15970,N_14151);
and U22060 (N_22060,N_16070,N_16631);
nor U22061 (N_22061,N_17939,N_15236);
nand U22062 (N_22062,N_18281,N_17440);
xor U22063 (N_22063,N_15358,N_18625);
nand U22064 (N_22064,N_17011,N_16004);
or U22065 (N_22065,N_12855,N_13148);
nor U22066 (N_22066,N_17850,N_15263);
nand U22067 (N_22067,N_17105,N_16365);
nor U22068 (N_22068,N_15793,N_12646);
and U22069 (N_22069,N_18214,N_16714);
and U22070 (N_22070,N_18337,N_13971);
or U22071 (N_22071,N_18181,N_14262);
and U22072 (N_22072,N_18612,N_16202);
nor U22073 (N_22073,N_13838,N_17832);
and U22074 (N_22074,N_12943,N_15671);
nand U22075 (N_22075,N_14801,N_16835);
or U22076 (N_22076,N_17963,N_12785);
nor U22077 (N_22077,N_13123,N_17753);
nor U22078 (N_22078,N_15067,N_17874);
nand U22079 (N_22079,N_14768,N_18535);
nand U22080 (N_22080,N_14351,N_14861);
nor U22081 (N_22081,N_14137,N_14196);
nand U22082 (N_22082,N_12907,N_15455);
nor U22083 (N_22083,N_14103,N_14925);
nor U22084 (N_22084,N_13984,N_13725);
nor U22085 (N_22085,N_18059,N_18702);
and U22086 (N_22086,N_12991,N_15366);
nand U22087 (N_22087,N_17570,N_17095);
and U22088 (N_22088,N_18725,N_16297);
nand U22089 (N_22089,N_16350,N_13434);
xnor U22090 (N_22090,N_15137,N_15286);
xor U22091 (N_22091,N_13482,N_15093);
xnor U22092 (N_22092,N_12798,N_17308);
and U22093 (N_22093,N_12627,N_14372);
and U22094 (N_22094,N_16176,N_16289);
or U22095 (N_22095,N_12751,N_15747);
or U22096 (N_22096,N_16778,N_14049);
and U22097 (N_22097,N_18499,N_18028);
nor U22098 (N_22098,N_16432,N_12516);
nor U22099 (N_22099,N_12723,N_18312);
or U22100 (N_22100,N_18639,N_16325);
nor U22101 (N_22101,N_14387,N_17727);
or U22102 (N_22102,N_13267,N_18180);
or U22103 (N_22103,N_16800,N_14290);
nand U22104 (N_22104,N_13387,N_16530);
and U22105 (N_22105,N_13615,N_15033);
nor U22106 (N_22106,N_17882,N_13861);
or U22107 (N_22107,N_15989,N_13145);
or U22108 (N_22108,N_14556,N_18196);
xor U22109 (N_22109,N_17798,N_17034);
and U22110 (N_22110,N_16233,N_14350);
and U22111 (N_22111,N_15508,N_13616);
or U22112 (N_22112,N_13991,N_16056);
nand U22113 (N_22113,N_13586,N_13821);
nand U22114 (N_22114,N_14254,N_14512);
or U22115 (N_22115,N_15277,N_18526);
xnor U22116 (N_22116,N_17156,N_16620);
nor U22117 (N_22117,N_12848,N_14630);
or U22118 (N_22118,N_16028,N_14720);
and U22119 (N_22119,N_13353,N_17194);
nand U22120 (N_22120,N_15073,N_15181);
nor U22121 (N_22121,N_17822,N_14369);
or U22122 (N_22122,N_13599,N_13392);
xnor U22123 (N_22123,N_16331,N_18317);
and U22124 (N_22124,N_18130,N_17345);
and U22125 (N_22125,N_15925,N_17968);
or U22126 (N_22126,N_15716,N_12741);
and U22127 (N_22127,N_14247,N_18678);
nor U22128 (N_22128,N_13312,N_13229);
nor U22129 (N_22129,N_15911,N_18342);
and U22130 (N_22130,N_17450,N_15175);
nor U22131 (N_22131,N_15125,N_16424);
xor U22132 (N_22132,N_17417,N_14452);
and U22133 (N_22133,N_18354,N_12999);
or U22134 (N_22134,N_15884,N_18595);
nor U22135 (N_22135,N_14733,N_18025);
and U22136 (N_22136,N_15732,N_15447);
nor U22137 (N_22137,N_14148,N_17545);
and U22138 (N_22138,N_14327,N_13226);
or U22139 (N_22139,N_15507,N_18132);
nor U22140 (N_22140,N_15334,N_14100);
nor U22141 (N_22141,N_17098,N_16736);
or U22142 (N_22142,N_16070,N_15225);
nand U22143 (N_22143,N_13630,N_16121);
xnor U22144 (N_22144,N_16222,N_12713);
xnor U22145 (N_22145,N_13388,N_18022);
and U22146 (N_22146,N_13806,N_14301);
and U22147 (N_22147,N_15889,N_15470);
or U22148 (N_22148,N_16198,N_14724);
nor U22149 (N_22149,N_15371,N_14620);
xnor U22150 (N_22150,N_18229,N_15455);
or U22151 (N_22151,N_15944,N_14778);
xor U22152 (N_22152,N_18609,N_15659);
nand U22153 (N_22153,N_17760,N_14020);
nand U22154 (N_22154,N_17569,N_17717);
nor U22155 (N_22155,N_16782,N_17172);
nor U22156 (N_22156,N_12778,N_18496);
and U22157 (N_22157,N_17537,N_13896);
xnor U22158 (N_22158,N_18374,N_12713);
nand U22159 (N_22159,N_13045,N_14174);
or U22160 (N_22160,N_13511,N_12858);
and U22161 (N_22161,N_13116,N_14078);
nand U22162 (N_22162,N_16068,N_16239);
and U22163 (N_22163,N_14194,N_17401);
and U22164 (N_22164,N_16452,N_15913);
nor U22165 (N_22165,N_18603,N_16546);
or U22166 (N_22166,N_18657,N_15992);
or U22167 (N_22167,N_18719,N_15077);
nand U22168 (N_22168,N_15938,N_14221);
or U22169 (N_22169,N_16611,N_15458);
or U22170 (N_22170,N_14889,N_18521);
or U22171 (N_22171,N_16221,N_17042);
and U22172 (N_22172,N_16853,N_14554);
nor U22173 (N_22173,N_17767,N_13744);
xor U22174 (N_22174,N_18090,N_14273);
nor U22175 (N_22175,N_18109,N_14457);
and U22176 (N_22176,N_17632,N_15148);
and U22177 (N_22177,N_12585,N_17269);
and U22178 (N_22178,N_18533,N_16012);
nor U22179 (N_22179,N_18574,N_14741);
xor U22180 (N_22180,N_12511,N_14289);
xor U22181 (N_22181,N_12714,N_14165);
xnor U22182 (N_22182,N_14775,N_13683);
or U22183 (N_22183,N_18559,N_15033);
and U22184 (N_22184,N_17924,N_18403);
nor U22185 (N_22185,N_15229,N_18246);
and U22186 (N_22186,N_12883,N_18249);
and U22187 (N_22187,N_14551,N_13132);
nand U22188 (N_22188,N_14344,N_14912);
or U22189 (N_22189,N_17826,N_17158);
xnor U22190 (N_22190,N_18585,N_13125);
xor U22191 (N_22191,N_13799,N_15824);
nand U22192 (N_22192,N_14977,N_15580);
nor U22193 (N_22193,N_15245,N_13490);
and U22194 (N_22194,N_12915,N_17287);
nor U22195 (N_22195,N_15553,N_13439);
and U22196 (N_22196,N_16839,N_17682);
or U22197 (N_22197,N_16467,N_12787);
and U22198 (N_22198,N_17893,N_17741);
and U22199 (N_22199,N_13110,N_12980);
or U22200 (N_22200,N_13856,N_13150);
nand U22201 (N_22201,N_17387,N_13944);
or U22202 (N_22202,N_13507,N_14335);
xnor U22203 (N_22203,N_14352,N_15839);
nor U22204 (N_22204,N_16402,N_12804);
nand U22205 (N_22205,N_13592,N_17918);
or U22206 (N_22206,N_14828,N_17694);
nor U22207 (N_22207,N_16669,N_13145);
nor U22208 (N_22208,N_14900,N_14907);
and U22209 (N_22209,N_12750,N_12608);
nand U22210 (N_22210,N_14879,N_14872);
nor U22211 (N_22211,N_14172,N_13675);
nand U22212 (N_22212,N_15261,N_16038);
and U22213 (N_22213,N_16496,N_16407);
nor U22214 (N_22214,N_13222,N_17448);
nor U22215 (N_22215,N_16447,N_17024);
and U22216 (N_22216,N_18437,N_17389);
nand U22217 (N_22217,N_17453,N_13708);
xor U22218 (N_22218,N_14678,N_13221);
and U22219 (N_22219,N_15137,N_12967);
nor U22220 (N_22220,N_16674,N_15307);
or U22221 (N_22221,N_16476,N_13439);
and U22222 (N_22222,N_15174,N_14211);
xor U22223 (N_22223,N_15044,N_18313);
and U22224 (N_22224,N_13937,N_18021);
and U22225 (N_22225,N_17495,N_13471);
nand U22226 (N_22226,N_15978,N_18471);
xnor U22227 (N_22227,N_13919,N_15751);
xnor U22228 (N_22228,N_15481,N_13128);
xor U22229 (N_22229,N_14465,N_15200);
or U22230 (N_22230,N_14923,N_15619);
and U22231 (N_22231,N_16053,N_14228);
xnor U22232 (N_22232,N_17138,N_12848);
nor U22233 (N_22233,N_15735,N_18543);
and U22234 (N_22234,N_16797,N_14779);
nand U22235 (N_22235,N_14815,N_17054);
nor U22236 (N_22236,N_17440,N_17067);
or U22237 (N_22237,N_16647,N_18618);
nor U22238 (N_22238,N_18682,N_14422);
nor U22239 (N_22239,N_14019,N_13206);
or U22240 (N_22240,N_16427,N_18463);
nand U22241 (N_22241,N_13042,N_13225);
xnor U22242 (N_22242,N_17807,N_14309);
nor U22243 (N_22243,N_15876,N_15303);
xor U22244 (N_22244,N_17409,N_18069);
xor U22245 (N_22245,N_16310,N_13533);
nand U22246 (N_22246,N_14740,N_15432);
nand U22247 (N_22247,N_16858,N_15417);
nor U22248 (N_22248,N_15694,N_12736);
and U22249 (N_22249,N_17265,N_15127);
nand U22250 (N_22250,N_15370,N_14596);
nand U22251 (N_22251,N_15350,N_13861);
nor U22252 (N_22252,N_14051,N_15328);
xnor U22253 (N_22253,N_14158,N_13369);
nor U22254 (N_22254,N_18675,N_14923);
nor U22255 (N_22255,N_14166,N_16317);
or U22256 (N_22256,N_18063,N_18349);
nor U22257 (N_22257,N_15151,N_14353);
and U22258 (N_22258,N_15784,N_14127);
nor U22259 (N_22259,N_13808,N_17357);
nor U22260 (N_22260,N_13022,N_17630);
nor U22261 (N_22261,N_15965,N_17586);
and U22262 (N_22262,N_13245,N_14700);
xor U22263 (N_22263,N_15552,N_13005);
or U22264 (N_22264,N_14078,N_16171);
and U22265 (N_22265,N_15855,N_16304);
or U22266 (N_22266,N_13844,N_13146);
and U22267 (N_22267,N_15389,N_14945);
and U22268 (N_22268,N_15202,N_16937);
nor U22269 (N_22269,N_16981,N_16474);
and U22270 (N_22270,N_16857,N_15443);
nor U22271 (N_22271,N_16625,N_15894);
or U22272 (N_22272,N_16395,N_17773);
nand U22273 (N_22273,N_14620,N_13408);
nor U22274 (N_22274,N_17645,N_15232);
xnor U22275 (N_22275,N_14030,N_14897);
nor U22276 (N_22276,N_13385,N_15363);
and U22277 (N_22277,N_18427,N_15916);
xor U22278 (N_22278,N_13934,N_15972);
or U22279 (N_22279,N_17099,N_18723);
nor U22280 (N_22280,N_13037,N_12814);
or U22281 (N_22281,N_13395,N_16817);
nor U22282 (N_22282,N_18200,N_18674);
nand U22283 (N_22283,N_17700,N_12615);
or U22284 (N_22284,N_18127,N_15760);
nand U22285 (N_22285,N_16843,N_15248);
nor U22286 (N_22286,N_17675,N_15142);
nand U22287 (N_22287,N_13590,N_13891);
nor U22288 (N_22288,N_16087,N_15264);
or U22289 (N_22289,N_16467,N_14997);
nor U22290 (N_22290,N_17345,N_15863);
nand U22291 (N_22291,N_13082,N_16266);
xnor U22292 (N_22292,N_18697,N_17071);
nand U22293 (N_22293,N_16975,N_17611);
and U22294 (N_22294,N_14304,N_13906);
nor U22295 (N_22295,N_15875,N_16667);
nor U22296 (N_22296,N_15942,N_18518);
nand U22297 (N_22297,N_12749,N_18034);
and U22298 (N_22298,N_17483,N_17501);
nor U22299 (N_22299,N_18120,N_17126);
nand U22300 (N_22300,N_17643,N_14105);
nand U22301 (N_22301,N_12516,N_15689);
and U22302 (N_22302,N_14167,N_18511);
xor U22303 (N_22303,N_17767,N_14197);
and U22304 (N_22304,N_15198,N_17424);
nand U22305 (N_22305,N_17618,N_13867);
or U22306 (N_22306,N_13032,N_16875);
or U22307 (N_22307,N_18247,N_13436);
xnor U22308 (N_22308,N_15004,N_17733);
xor U22309 (N_22309,N_15024,N_18235);
nor U22310 (N_22310,N_18031,N_15286);
and U22311 (N_22311,N_16989,N_16484);
nor U22312 (N_22312,N_18102,N_15314);
xnor U22313 (N_22313,N_17515,N_13694);
or U22314 (N_22314,N_13641,N_14514);
nor U22315 (N_22315,N_13477,N_12834);
and U22316 (N_22316,N_17863,N_14343);
xor U22317 (N_22317,N_17131,N_15523);
nand U22318 (N_22318,N_16993,N_18166);
nor U22319 (N_22319,N_12581,N_12627);
and U22320 (N_22320,N_15855,N_12903);
nand U22321 (N_22321,N_13006,N_13638);
and U22322 (N_22322,N_13165,N_15813);
nor U22323 (N_22323,N_18664,N_13998);
and U22324 (N_22324,N_18643,N_15986);
or U22325 (N_22325,N_12985,N_12516);
xnor U22326 (N_22326,N_16334,N_14121);
and U22327 (N_22327,N_14648,N_16990);
nand U22328 (N_22328,N_14154,N_13174);
nor U22329 (N_22329,N_14490,N_16533);
xor U22330 (N_22330,N_17796,N_17509);
and U22331 (N_22331,N_12533,N_17135);
or U22332 (N_22332,N_12569,N_15479);
nand U22333 (N_22333,N_13478,N_15073);
nand U22334 (N_22334,N_13117,N_14485);
or U22335 (N_22335,N_15735,N_14751);
nand U22336 (N_22336,N_16468,N_14551);
xnor U22337 (N_22337,N_15622,N_17264);
nor U22338 (N_22338,N_18053,N_13069);
xnor U22339 (N_22339,N_15698,N_18549);
and U22340 (N_22340,N_18117,N_17941);
or U22341 (N_22341,N_15537,N_14667);
xor U22342 (N_22342,N_12558,N_12898);
xnor U22343 (N_22343,N_14043,N_17177);
nor U22344 (N_22344,N_16663,N_15105);
xnor U22345 (N_22345,N_15718,N_16507);
and U22346 (N_22346,N_12826,N_17049);
or U22347 (N_22347,N_16273,N_13364);
nor U22348 (N_22348,N_15715,N_16396);
nand U22349 (N_22349,N_17143,N_15204);
and U22350 (N_22350,N_13229,N_12537);
nor U22351 (N_22351,N_14053,N_17389);
nand U22352 (N_22352,N_16166,N_15531);
xor U22353 (N_22353,N_14089,N_14373);
and U22354 (N_22354,N_16790,N_14421);
nand U22355 (N_22355,N_14281,N_12785);
nor U22356 (N_22356,N_16488,N_13770);
or U22357 (N_22357,N_15700,N_18109);
nor U22358 (N_22358,N_14055,N_17318);
nand U22359 (N_22359,N_13005,N_15657);
and U22360 (N_22360,N_15822,N_16235);
nor U22361 (N_22361,N_15593,N_16128);
or U22362 (N_22362,N_14701,N_14015);
xnor U22363 (N_22363,N_16863,N_18349);
nand U22364 (N_22364,N_17581,N_13627);
or U22365 (N_22365,N_17833,N_18131);
nand U22366 (N_22366,N_14204,N_18739);
nand U22367 (N_22367,N_14943,N_18484);
nand U22368 (N_22368,N_18297,N_16247);
nand U22369 (N_22369,N_14954,N_13462);
nor U22370 (N_22370,N_13660,N_14197);
and U22371 (N_22371,N_17869,N_17264);
or U22372 (N_22372,N_17254,N_13014);
or U22373 (N_22373,N_17156,N_16180);
and U22374 (N_22374,N_12925,N_16471);
xor U22375 (N_22375,N_15104,N_14683);
nor U22376 (N_22376,N_18632,N_15745);
nand U22377 (N_22377,N_17010,N_13517);
or U22378 (N_22378,N_15829,N_13667);
or U22379 (N_22379,N_15847,N_13538);
nand U22380 (N_22380,N_17734,N_16729);
or U22381 (N_22381,N_18441,N_13971);
and U22382 (N_22382,N_16572,N_16967);
nor U22383 (N_22383,N_16150,N_15941);
nor U22384 (N_22384,N_18618,N_16779);
nor U22385 (N_22385,N_13211,N_15206);
and U22386 (N_22386,N_13181,N_12551);
and U22387 (N_22387,N_17582,N_18614);
xor U22388 (N_22388,N_17359,N_16398);
nor U22389 (N_22389,N_17829,N_16229);
and U22390 (N_22390,N_18421,N_14348);
and U22391 (N_22391,N_12712,N_13507);
and U22392 (N_22392,N_18345,N_14126);
xnor U22393 (N_22393,N_18579,N_18061);
nor U22394 (N_22394,N_17333,N_13708);
nor U22395 (N_22395,N_17446,N_17136);
nor U22396 (N_22396,N_16510,N_15525);
nor U22397 (N_22397,N_13542,N_18198);
xor U22398 (N_22398,N_14573,N_16747);
nor U22399 (N_22399,N_16640,N_16802);
and U22400 (N_22400,N_15722,N_12805);
xor U22401 (N_22401,N_17677,N_18220);
or U22402 (N_22402,N_17182,N_12827);
nor U22403 (N_22403,N_14168,N_17998);
and U22404 (N_22404,N_14688,N_12888);
xor U22405 (N_22405,N_16050,N_16218);
or U22406 (N_22406,N_17587,N_14651);
or U22407 (N_22407,N_18563,N_18113);
and U22408 (N_22408,N_14300,N_14731);
xor U22409 (N_22409,N_17028,N_18734);
and U22410 (N_22410,N_14815,N_17267);
nor U22411 (N_22411,N_14268,N_15170);
nor U22412 (N_22412,N_17846,N_15243);
or U22413 (N_22413,N_13752,N_14698);
and U22414 (N_22414,N_16884,N_18330);
and U22415 (N_22415,N_12693,N_15654);
nor U22416 (N_22416,N_13050,N_12796);
nor U22417 (N_22417,N_18379,N_14485);
or U22418 (N_22418,N_18704,N_16025);
or U22419 (N_22419,N_16725,N_12553);
xnor U22420 (N_22420,N_13957,N_16595);
nand U22421 (N_22421,N_17260,N_13251);
nor U22422 (N_22422,N_17789,N_16432);
nor U22423 (N_22423,N_17793,N_14755);
and U22424 (N_22424,N_13523,N_17929);
or U22425 (N_22425,N_15998,N_15109);
or U22426 (N_22426,N_17541,N_12807);
nor U22427 (N_22427,N_15364,N_16367);
nand U22428 (N_22428,N_13135,N_15376);
and U22429 (N_22429,N_14847,N_15020);
or U22430 (N_22430,N_12618,N_18290);
nor U22431 (N_22431,N_17313,N_12738);
nand U22432 (N_22432,N_18329,N_13983);
nand U22433 (N_22433,N_16798,N_12882);
nand U22434 (N_22434,N_16903,N_18222);
or U22435 (N_22435,N_16399,N_12971);
nor U22436 (N_22436,N_13190,N_16237);
nand U22437 (N_22437,N_15065,N_12932);
nor U22438 (N_22438,N_16898,N_13912);
nor U22439 (N_22439,N_17789,N_16128);
nor U22440 (N_22440,N_12846,N_13448);
nor U22441 (N_22441,N_15567,N_16468);
or U22442 (N_22442,N_17726,N_12860);
xnor U22443 (N_22443,N_13062,N_13420);
or U22444 (N_22444,N_17362,N_15722);
nand U22445 (N_22445,N_12908,N_15719);
and U22446 (N_22446,N_16986,N_16428);
nor U22447 (N_22447,N_17451,N_13126);
or U22448 (N_22448,N_16567,N_18242);
nor U22449 (N_22449,N_14452,N_16984);
or U22450 (N_22450,N_16595,N_13609);
or U22451 (N_22451,N_13320,N_17218);
and U22452 (N_22452,N_18622,N_17680);
xnor U22453 (N_22453,N_17357,N_16715);
nand U22454 (N_22454,N_18181,N_18081);
xnor U22455 (N_22455,N_13895,N_15047);
nand U22456 (N_22456,N_16060,N_14162);
or U22457 (N_22457,N_18383,N_17636);
nor U22458 (N_22458,N_13303,N_12720);
nor U22459 (N_22459,N_17944,N_18716);
or U22460 (N_22460,N_15016,N_16118);
and U22461 (N_22461,N_16398,N_16818);
nand U22462 (N_22462,N_12842,N_14053);
nor U22463 (N_22463,N_17146,N_17813);
xor U22464 (N_22464,N_18331,N_15234);
xor U22465 (N_22465,N_18006,N_12508);
xor U22466 (N_22466,N_17407,N_16104);
or U22467 (N_22467,N_18574,N_17196);
xor U22468 (N_22468,N_13929,N_15028);
and U22469 (N_22469,N_12610,N_15993);
nor U22470 (N_22470,N_18606,N_15912);
and U22471 (N_22471,N_15692,N_13870);
and U22472 (N_22472,N_16548,N_18745);
and U22473 (N_22473,N_17526,N_18113);
and U22474 (N_22474,N_13639,N_15438);
xor U22475 (N_22475,N_14330,N_15891);
or U22476 (N_22476,N_13121,N_16947);
and U22477 (N_22477,N_13472,N_17303);
nor U22478 (N_22478,N_13012,N_13480);
and U22479 (N_22479,N_15816,N_14213);
nor U22480 (N_22480,N_16411,N_13894);
nand U22481 (N_22481,N_13675,N_14192);
nand U22482 (N_22482,N_16076,N_14761);
nand U22483 (N_22483,N_16873,N_14827);
nand U22484 (N_22484,N_16208,N_14238);
nand U22485 (N_22485,N_14222,N_16525);
nor U22486 (N_22486,N_13717,N_13838);
nor U22487 (N_22487,N_14546,N_13852);
or U22488 (N_22488,N_13769,N_14188);
nand U22489 (N_22489,N_14905,N_15604);
nor U22490 (N_22490,N_14511,N_16107);
or U22491 (N_22491,N_18178,N_13645);
nand U22492 (N_22492,N_13209,N_16531);
nand U22493 (N_22493,N_14047,N_17175);
xnor U22494 (N_22494,N_13082,N_15313);
and U22495 (N_22495,N_14136,N_14629);
nand U22496 (N_22496,N_14754,N_16608);
and U22497 (N_22497,N_14786,N_18297);
xnor U22498 (N_22498,N_13040,N_17865);
nor U22499 (N_22499,N_13745,N_17306);
nor U22500 (N_22500,N_16040,N_13225);
nand U22501 (N_22501,N_18413,N_12655);
and U22502 (N_22502,N_14738,N_14437);
xor U22503 (N_22503,N_12658,N_13477);
and U22504 (N_22504,N_18160,N_17548);
or U22505 (N_22505,N_13859,N_18680);
xnor U22506 (N_22506,N_12636,N_14896);
or U22507 (N_22507,N_13698,N_17097);
and U22508 (N_22508,N_13485,N_17053);
xnor U22509 (N_22509,N_18214,N_17652);
nand U22510 (N_22510,N_14146,N_14917);
nor U22511 (N_22511,N_14335,N_15493);
and U22512 (N_22512,N_14136,N_18494);
xnor U22513 (N_22513,N_17520,N_15634);
nand U22514 (N_22514,N_16687,N_12828);
or U22515 (N_22515,N_14021,N_14202);
or U22516 (N_22516,N_13248,N_18560);
xor U22517 (N_22517,N_16027,N_15201);
xnor U22518 (N_22518,N_15257,N_16153);
or U22519 (N_22519,N_16416,N_13199);
nand U22520 (N_22520,N_13565,N_14287);
nor U22521 (N_22521,N_17418,N_12788);
xnor U22522 (N_22522,N_16511,N_17781);
nand U22523 (N_22523,N_16662,N_16291);
xnor U22524 (N_22524,N_12536,N_18562);
xnor U22525 (N_22525,N_18495,N_12683);
and U22526 (N_22526,N_16975,N_17748);
xor U22527 (N_22527,N_17367,N_12752);
or U22528 (N_22528,N_13637,N_16135);
and U22529 (N_22529,N_14299,N_18457);
xnor U22530 (N_22530,N_16082,N_13337);
nor U22531 (N_22531,N_17754,N_13637);
nor U22532 (N_22532,N_16518,N_17734);
nor U22533 (N_22533,N_17811,N_13285);
nand U22534 (N_22534,N_13820,N_17359);
xnor U22535 (N_22535,N_15450,N_15307);
nand U22536 (N_22536,N_17097,N_16220);
nor U22537 (N_22537,N_15225,N_16588);
and U22538 (N_22538,N_15858,N_16506);
xor U22539 (N_22539,N_15642,N_15208);
and U22540 (N_22540,N_16697,N_18490);
or U22541 (N_22541,N_14628,N_14161);
or U22542 (N_22542,N_17402,N_13926);
or U22543 (N_22543,N_13548,N_14643);
nand U22544 (N_22544,N_17575,N_14533);
or U22545 (N_22545,N_16476,N_14535);
and U22546 (N_22546,N_17988,N_15586);
xnor U22547 (N_22547,N_17210,N_14691);
or U22548 (N_22548,N_14173,N_15101);
nor U22549 (N_22549,N_14695,N_12680);
or U22550 (N_22550,N_18736,N_18157);
nor U22551 (N_22551,N_17535,N_13541);
nor U22552 (N_22552,N_14026,N_18310);
or U22553 (N_22553,N_18491,N_14370);
and U22554 (N_22554,N_13802,N_16993);
xor U22555 (N_22555,N_17366,N_13362);
nand U22556 (N_22556,N_17135,N_13355);
or U22557 (N_22557,N_17562,N_17612);
xor U22558 (N_22558,N_13303,N_17437);
and U22559 (N_22559,N_16320,N_14360);
and U22560 (N_22560,N_13425,N_13368);
nor U22561 (N_22561,N_17353,N_13379);
xnor U22562 (N_22562,N_14836,N_16727);
or U22563 (N_22563,N_17810,N_14463);
or U22564 (N_22564,N_14304,N_16414);
nor U22565 (N_22565,N_14625,N_17885);
and U22566 (N_22566,N_14857,N_14832);
xnor U22567 (N_22567,N_15707,N_14577);
and U22568 (N_22568,N_13206,N_18312);
nor U22569 (N_22569,N_15858,N_17087);
and U22570 (N_22570,N_16718,N_18743);
and U22571 (N_22571,N_16689,N_14384);
or U22572 (N_22572,N_16721,N_16318);
and U22573 (N_22573,N_16511,N_12552);
xnor U22574 (N_22574,N_14761,N_13938);
xor U22575 (N_22575,N_15797,N_14232);
nor U22576 (N_22576,N_15653,N_14753);
and U22577 (N_22577,N_17486,N_14574);
nor U22578 (N_22578,N_16685,N_14079);
or U22579 (N_22579,N_12887,N_14016);
nand U22580 (N_22580,N_15898,N_16780);
nand U22581 (N_22581,N_15269,N_16476);
xnor U22582 (N_22582,N_18231,N_16445);
and U22583 (N_22583,N_17652,N_15966);
nor U22584 (N_22584,N_14138,N_13536);
nor U22585 (N_22585,N_15847,N_13341);
nor U22586 (N_22586,N_18622,N_16828);
and U22587 (N_22587,N_13926,N_16065);
xor U22588 (N_22588,N_14882,N_13441);
nor U22589 (N_22589,N_12975,N_12611);
nor U22590 (N_22590,N_17190,N_15012);
xnor U22591 (N_22591,N_15947,N_15910);
nor U22592 (N_22592,N_13944,N_17997);
nor U22593 (N_22593,N_14981,N_16607);
or U22594 (N_22594,N_16823,N_15381);
and U22595 (N_22595,N_18081,N_14325);
and U22596 (N_22596,N_16789,N_15848);
or U22597 (N_22597,N_12654,N_15621);
or U22598 (N_22598,N_15753,N_16959);
nor U22599 (N_22599,N_18440,N_18047);
xor U22600 (N_22600,N_16981,N_18282);
nand U22601 (N_22601,N_13293,N_14486);
xnor U22602 (N_22602,N_15120,N_17646);
nor U22603 (N_22603,N_16272,N_16012);
xor U22604 (N_22604,N_16646,N_15598);
and U22605 (N_22605,N_14777,N_18157);
nand U22606 (N_22606,N_16397,N_18383);
xnor U22607 (N_22607,N_16472,N_12838);
or U22608 (N_22608,N_16832,N_17350);
nor U22609 (N_22609,N_16147,N_16713);
xnor U22610 (N_22610,N_16060,N_14471);
and U22611 (N_22611,N_15567,N_17025);
xnor U22612 (N_22612,N_16902,N_18215);
nor U22613 (N_22613,N_15607,N_17987);
nand U22614 (N_22614,N_15812,N_17066);
xor U22615 (N_22615,N_17521,N_17562);
xor U22616 (N_22616,N_13458,N_18622);
and U22617 (N_22617,N_15489,N_16273);
nand U22618 (N_22618,N_15929,N_14017);
or U22619 (N_22619,N_13212,N_15462);
or U22620 (N_22620,N_17510,N_16759);
nor U22621 (N_22621,N_15475,N_15829);
nand U22622 (N_22622,N_17409,N_14802);
and U22623 (N_22623,N_16594,N_17759);
or U22624 (N_22624,N_16469,N_16920);
nor U22625 (N_22625,N_18542,N_17496);
and U22626 (N_22626,N_17110,N_17705);
xnor U22627 (N_22627,N_17330,N_14891);
or U22628 (N_22628,N_18039,N_13715);
or U22629 (N_22629,N_17688,N_17254);
and U22630 (N_22630,N_16305,N_15383);
nor U22631 (N_22631,N_15842,N_12566);
nor U22632 (N_22632,N_16831,N_15086);
xor U22633 (N_22633,N_14460,N_15352);
and U22634 (N_22634,N_17698,N_18493);
nand U22635 (N_22635,N_15944,N_16642);
nand U22636 (N_22636,N_13053,N_12923);
and U22637 (N_22637,N_13218,N_15597);
nor U22638 (N_22638,N_14642,N_13838);
nand U22639 (N_22639,N_14706,N_17407);
nand U22640 (N_22640,N_14131,N_15585);
nor U22641 (N_22641,N_13848,N_15742);
and U22642 (N_22642,N_13456,N_18743);
or U22643 (N_22643,N_13714,N_12956);
or U22644 (N_22644,N_17939,N_17331);
and U22645 (N_22645,N_16308,N_12766);
and U22646 (N_22646,N_15475,N_18172);
xor U22647 (N_22647,N_16521,N_15027);
xnor U22648 (N_22648,N_13601,N_12996);
nor U22649 (N_22649,N_13192,N_18050);
nor U22650 (N_22650,N_17692,N_17616);
nand U22651 (N_22651,N_17778,N_18649);
or U22652 (N_22652,N_16108,N_18081);
or U22653 (N_22653,N_14482,N_13939);
and U22654 (N_22654,N_12899,N_18154);
nand U22655 (N_22655,N_16256,N_17961);
and U22656 (N_22656,N_15399,N_18195);
or U22657 (N_22657,N_16854,N_17489);
and U22658 (N_22658,N_18244,N_15022);
nor U22659 (N_22659,N_16342,N_17044);
xnor U22660 (N_22660,N_15432,N_13808);
and U22661 (N_22661,N_15347,N_18008);
nor U22662 (N_22662,N_15321,N_16581);
nor U22663 (N_22663,N_18177,N_16088);
and U22664 (N_22664,N_18724,N_14032);
xor U22665 (N_22665,N_14940,N_13567);
nor U22666 (N_22666,N_17582,N_16880);
and U22667 (N_22667,N_15941,N_15969);
xnor U22668 (N_22668,N_14058,N_16118);
and U22669 (N_22669,N_13755,N_16121);
nand U22670 (N_22670,N_14662,N_18623);
xor U22671 (N_22671,N_16892,N_16577);
nand U22672 (N_22672,N_15701,N_15645);
or U22673 (N_22673,N_16544,N_14681);
nor U22674 (N_22674,N_17819,N_18704);
xnor U22675 (N_22675,N_15839,N_14896);
nand U22676 (N_22676,N_14056,N_15342);
nand U22677 (N_22677,N_17981,N_14510);
nand U22678 (N_22678,N_15063,N_17840);
and U22679 (N_22679,N_15574,N_13907);
and U22680 (N_22680,N_14053,N_14360);
nor U22681 (N_22681,N_14070,N_15587);
nor U22682 (N_22682,N_17529,N_17758);
nand U22683 (N_22683,N_13307,N_16721);
xnor U22684 (N_22684,N_18202,N_14682);
nand U22685 (N_22685,N_17364,N_13075);
and U22686 (N_22686,N_18739,N_18256);
nand U22687 (N_22687,N_14969,N_16065);
nand U22688 (N_22688,N_17881,N_16229);
or U22689 (N_22689,N_12571,N_15296);
xor U22690 (N_22690,N_13566,N_16105);
or U22691 (N_22691,N_15449,N_17292);
nor U22692 (N_22692,N_12718,N_15931);
nor U22693 (N_22693,N_14332,N_13287);
and U22694 (N_22694,N_13701,N_18261);
nor U22695 (N_22695,N_18721,N_14072);
nor U22696 (N_22696,N_16482,N_17489);
and U22697 (N_22697,N_14846,N_17750);
or U22698 (N_22698,N_13975,N_17886);
and U22699 (N_22699,N_14255,N_18302);
nand U22700 (N_22700,N_15655,N_12727);
and U22701 (N_22701,N_17975,N_15047);
xnor U22702 (N_22702,N_16820,N_13445);
nand U22703 (N_22703,N_12592,N_17219);
nand U22704 (N_22704,N_14342,N_12914);
and U22705 (N_22705,N_13757,N_17555);
nand U22706 (N_22706,N_13592,N_15486);
nor U22707 (N_22707,N_13790,N_12780);
and U22708 (N_22708,N_13719,N_13246);
nand U22709 (N_22709,N_12582,N_18212);
nor U22710 (N_22710,N_18143,N_12909);
nor U22711 (N_22711,N_18205,N_15759);
nand U22712 (N_22712,N_18113,N_16210);
nand U22713 (N_22713,N_13973,N_15591);
or U22714 (N_22714,N_13428,N_15441);
nor U22715 (N_22715,N_15377,N_13607);
and U22716 (N_22716,N_14284,N_18737);
nor U22717 (N_22717,N_13831,N_17525);
or U22718 (N_22718,N_18535,N_18267);
nand U22719 (N_22719,N_18343,N_17550);
xor U22720 (N_22720,N_12602,N_15406);
and U22721 (N_22721,N_12700,N_18314);
nand U22722 (N_22722,N_12964,N_18417);
or U22723 (N_22723,N_17766,N_15476);
xnor U22724 (N_22724,N_18255,N_13622);
xnor U22725 (N_22725,N_13612,N_12674);
nor U22726 (N_22726,N_15866,N_15933);
and U22727 (N_22727,N_17261,N_12648);
xor U22728 (N_22728,N_18081,N_12525);
and U22729 (N_22729,N_16492,N_17959);
nand U22730 (N_22730,N_17586,N_16438);
nor U22731 (N_22731,N_16136,N_14746);
and U22732 (N_22732,N_13878,N_13437);
or U22733 (N_22733,N_13976,N_14723);
nor U22734 (N_22734,N_13457,N_15936);
nor U22735 (N_22735,N_13104,N_13095);
xnor U22736 (N_22736,N_17864,N_14248);
nand U22737 (N_22737,N_15429,N_13874);
xor U22738 (N_22738,N_14123,N_14651);
nor U22739 (N_22739,N_13978,N_13429);
xnor U22740 (N_22740,N_17839,N_18489);
xor U22741 (N_22741,N_18460,N_12554);
or U22742 (N_22742,N_13412,N_13745);
nand U22743 (N_22743,N_14184,N_15489);
nor U22744 (N_22744,N_17237,N_18245);
nand U22745 (N_22745,N_15616,N_14429);
nand U22746 (N_22746,N_17317,N_14129);
nor U22747 (N_22747,N_12654,N_13382);
nand U22748 (N_22748,N_17426,N_15622);
nor U22749 (N_22749,N_16263,N_13060);
nor U22750 (N_22750,N_17240,N_16485);
and U22751 (N_22751,N_12963,N_13198);
or U22752 (N_22752,N_16383,N_12819);
and U22753 (N_22753,N_14120,N_17232);
and U22754 (N_22754,N_18573,N_13612);
nand U22755 (N_22755,N_15258,N_18142);
nor U22756 (N_22756,N_14078,N_17973);
xnor U22757 (N_22757,N_18383,N_13088);
nor U22758 (N_22758,N_14522,N_17084);
xor U22759 (N_22759,N_15405,N_12521);
nor U22760 (N_22760,N_13784,N_16815);
nand U22761 (N_22761,N_14795,N_15601);
xnor U22762 (N_22762,N_13176,N_18004);
or U22763 (N_22763,N_15327,N_12644);
and U22764 (N_22764,N_12821,N_18572);
or U22765 (N_22765,N_13688,N_13133);
and U22766 (N_22766,N_16482,N_15381);
xnor U22767 (N_22767,N_16038,N_13408);
and U22768 (N_22768,N_18535,N_17494);
or U22769 (N_22769,N_13874,N_15320);
xnor U22770 (N_22770,N_15046,N_16484);
nand U22771 (N_22771,N_18184,N_14271);
and U22772 (N_22772,N_13730,N_15121);
nor U22773 (N_22773,N_13077,N_14685);
or U22774 (N_22774,N_13618,N_18253);
and U22775 (N_22775,N_16931,N_15160);
xnor U22776 (N_22776,N_14093,N_14750);
or U22777 (N_22777,N_12856,N_13748);
xnor U22778 (N_22778,N_14965,N_14019);
nand U22779 (N_22779,N_17682,N_17433);
and U22780 (N_22780,N_13317,N_16172);
or U22781 (N_22781,N_14090,N_14510);
and U22782 (N_22782,N_14313,N_12995);
xor U22783 (N_22783,N_14351,N_12696);
and U22784 (N_22784,N_13350,N_17115);
and U22785 (N_22785,N_14256,N_15931);
nor U22786 (N_22786,N_13782,N_17258);
nor U22787 (N_22787,N_14530,N_16079);
and U22788 (N_22788,N_18257,N_17624);
xnor U22789 (N_22789,N_15591,N_12764);
xnor U22790 (N_22790,N_13518,N_17082);
nand U22791 (N_22791,N_18186,N_12910);
nand U22792 (N_22792,N_18292,N_17216);
or U22793 (N_22793,N_18086,N_16741);
nor U22794 (N_22794,N_18209,N_12756);
or U22795 (N_22795,N_18027,N_17621);
xor U22796 (N_22796,N_16723,N_17302);
xor U22797 (N_22797,N_14055,N_15425);
or U22798 (N_22798,N_16186,N_18085);
or U22799 (N_22799,N_14407,N_16054);
nand U22800 (N_22800,N_16456,N_14470);
nor U22801 (N_22801,N_14350,N_15760);
xor U22802 (N_22802,N_16785,N_14153);
nor U22803 (N_22803,N_13907,N_13373);
nor U22804 (N_22804,N_14951,N_18065);
or U22805 (N_22805,N_18565,N_16649);
and U22806 (N_22806,N_18709,N_18051);
nor U22807 (N_22807,N_17294,N_17672);
or U22808 (N_22808,N_17783,N_13235);
nand U22809 (N_22809,N_15159,N_14903);
nor U22810 (N_22810,N_18485,N_14966);
xor U22811 (N_22811,N_13952,N_12707);
and U22812 (N_22812,N_14490,N_16420);
nand U22813 (N_22813,N_14023,N_15535);
and U22814 (N_22814,N_15879,N_16653);
xnor U22815 (N_22815,N_12893,N_13676);
nand U22816 (N_22816,N_15994,N_15279);
nand U22817 (N_22817,N_14585,N_14962);
and U22818 (N_22818,N_13422,N_14201);
nor U22819 (N_22819,N_12730,N_13364);
xnor U22820 (N_22820,N_15860,N_18678);
nand U22821 (N_22821,N_15856,N_16823);
or U22822 (N_22822,N_13205,N_17325);
or U22823 (N_22823,N_17038,N_17579);
nand U22824 (N_22824,N_17638,N_14549);
xnor U22825 (N_22825,N_12792,N_15113);
and U22826 (N_22826,N_15442,N_18040);
xnor U22827 (N_22827,N_16745,N_18036);
or U22828 (N_22828,N_16938,N_15704);
xnor U22829 (N_22829,N_16848,N_15795);
or U22830 (N_22830,N_18628,N_16825);
xnor U22831 (N_22831,N_14184,N_16880);
nand U22832 (N_22832,N_17350,N_17206);
or U22833 (N_22833,N_18564,N_12703);
xnor U22834 (N_22834,N_14333,N_14586);
nor U22835 (N_22835,N_12995,N_14985);
nand U22836 (N_22836,N_17915,N_15072);
xor U22837 (N_22837,N_14390,N_17522);
or U22838 (N_22838,N_17928,N_14006);
nand U22839 (N_22839,N_17147,N_17870);
xor U22840 (N_22840,N_13633,N_14329);
xor U22841 (N_22841,N_13678,N_12705);
nor U22842 (N_22842,N_12791,N_17152);
and U22843 (N_22843,N_16883,N_17120);
and U22844 (N_22844,N_17205,N_15491);
or U22845 (N_22845,N_14299,N_15643);
nand U22846 (N_22846,N_13311,N_13544);
xor U22847 (N_22847,N_17407,N_13515);
nor U22848 (N_22848,N_14261,N_14201);
nand U22849 (N_22849,N_14191,N_13963);
and U22850 (N_22850,N_12886,N_14286);
nand U22851 (N_22851,N_12940,N_14001);
or U22852 (N_22852,N_17392,N_12660);
xor U22853 (N_22853,N_16473,N_14376);
nand U22854 (N_22854,N_18160,N_17739);
nor U22855 (N_22855,N_17762,N_16312);
or U22856 (N_22856,N_14711,N_17893);
xnor U22857 (N_22857,N_15446,N_15670);
nand U22858 (N_22858,N_13892,N_17100);
xor U22859 (N_22859,N_15391,N_14759);
or U22860 (N_22860,N_18615,N_17659);
xnor U22861 (N_22861,N_15194,N_16507);
nor U22862 (N_22862,N_18577,N_15201);
xnor U22863 (N_22863,N_16422,N_16060);
nor U22864 (N_22864,N_15855,N_13714);
nand U22865 (N_22865,N_17591,N_14977);
xor U22866 (N_22866,N_15313,N_13767);
xnor U22867 (N_22867,N_17209,N_12789);
xor U22868 (N_22868,N_17791,N_15273);
nor U22869 (N_22869,N_17805,N_17751);
and U22870 (N_22870,N_15743,N_16903);
nand U22871 (N_22871,N_15834,N_16343);
or U22872 (N_22872,N_16958,N_17974);
nor U22873 (N_22873,N_16728,N_12920);
nor U22874 (N_22874,N_15403,N_16389);
nor U22875 (N_22875,N_14279,N_16377);
xnor U22876 (N_22876,N_13945,N_16090);
xor U22877 (N_22877,N_16862,N_17916);
or U22878 (N_22878,N_12602,N_14856);
or U22879 (N_22879,N_18110,N_15848);
nand U22880 (N_22880,N_15261,N_14752);
and U22881 (N_22881,N_18043,N_14381);
nand U22882 (N_22882,N_18474,N_18197);
nand U22883 (N_22883,N_17116,N_15920);
nand U22884 (N_22884,N_17776,N_18089);
xnor U22885 (N_22885,N_17080,N_14624);
xnor U22886 (N_22886,N_13167,N_14376);
or U22887 (N_22887,N_13738,N_14640);
and U22888 (N_22888,N_17632,N_14839);
and U22889 (N_22889,N_17512,N_14824);
and U22890 (N_22890,N_13286,N_12601);
nor U22891 (N_22891,N_16211,N_14637);
nor U22892 (N_22892,N_12511,N_13647);
and U22893 (N_22893,N_13283,N_18624);
and U22894 (N_22894,N_13027,N_16292);
nor U22895 (N_22895,N_18502,N_13695);
or U22896 (N_22896,N_17715,N_13589);
nor U22897 (N_22897,N_14887,N_18460);
or U22898 (N_22898,N_13839,N_18600);
or U22899 (N_22899,N_13292,N_14507);
xnor U22900 (N_22900,N_18362,N_12946);
and U22901 (N_22901,N_13729,N_16480);
and U22902 (N_22902,N_15940,N_15629);
nand U22903 (N_22903,N_17489,N_17349);
or U22904 (N_22904,N_15715,N_17943);
nor U22905 (N_22905,N_14403,N_17855);
nand U22906 (N_22906,N_14022,N_15356);
or U22907 (N_22907,N_16209,N_13796);
nor U22908 (N_22908,N_15407,N_13871);
or U22909 (N_22909,N_16142,N_15256);
xor U22910 (N_22910,N_18211,N_15530);
nand U22911 (N_22911,N_14936,N_16865);
and U22912 (N_22912,N_16715,N_12864);
or U22913 (N_22913,N_16897,N_13736);
or U22914 (N_22914,N_18404,N_14494);
or U22915 (N_22915,N_15740,N_16468);
and U22916 (N_22916,N_13649,N_14323);
xnor U22917 (N_22917,N_18041,N_13291);
xnor U22918 (N_22918,N_13930,N_17279);
xor U22919 (N_22919,N_16586,N_17333);
nand U22920 (N_22920,N_15049,N_14130);
nand U22921 (N_22921,N_14557,N_17005);
nor U22922 (N_22922,N_16941,N_16874);
xor U22923 (N_22923,N_14808,N_16764);
or U22924 (N_22924,N_12590,N_12767);
xnor U22925 (N_22925,N_17435,N_13945);
nand U22926 (N_22926,N_16304,N_16966);
or U22927 (N_22927,N_14588,N_14917);
nor U22928 (N_22928,N_18367,N_12647);
or U22929 (N_22929,N_15762,N_17556);
or U22930 (N_22930,N_17021,N_14863);
xnor U22931 (N_22931,N_16241,N_16995);
nor U22932 (N_22932,N_15647,N_17564);
and U22933 (N_22933,N_18205,N_15740);
nand U22934 (N_22934,N_12983,N_14977);
xor U22935 (N_22935,N_14913,N_15965);
and U22936 (N_22936,N_18241,N_13216);
xnor U22937 (N_22937,N_14212,N_15452);
nor U22938 (N_22938,N_18441,N_16381);
nor U22939 (N_22939,N_14536,N_15871);
or U22940 (N_22940,N_18491,N_14848);
and U22941 (N_22941,N_18515,N_15582);
nand U22942 (N_22942,N_12514,N_14983);
xnor U22943 (N_22943,N_12705,N_17206);
nand U22944 (N_22944,N_16287,N_16774);
and U22945 (N_22945,N_13870,N_13586);
nand U22946 (N_22946,N_15973,N_16999);
nand U22947 (N_22947,N_14652,N_14087);
nand U22948 (N_22948,N_12833,N_14183);
nand U22949 (N_22949,N_13513,N_15890);
nand U22950 (N_22950,N_13105,N_16076);
or U22951 (N_22951,N_17762,N_18276);
and U22952 (N_22952,N_15807,N_14931);
nand U22953 (N_22953,N_16332,N_13942);
nor U22954 (N_22954,N_14111,N_18471);
nor U22955 (N_22955,N_13360,N_16512);
nor U22956 (N_22956,N_15852,N_16568);
xnor U22957 (N_22957,N_12595,N_15056);
nand U22958 (N_22958,N_15120,N_15594);
or U22959 (N_22959,N_14751,N_12840);
or U22960 (N_22960,N_16857,N_14838);
nand U22961 (N_22961,N_15429,N_16760);
xnor U22962 (N_22962,N_18713,N_15224);
and U22963 (N_22963,N_16423,N_14081);
nand U22964 (N_22964,N_14618,N_16813);
and U22965 (N_22965,N_15245,N_15537);
nand U22966 (N_22966,N_15486,N_12835);
xnor U22967 (N_22967,N_14763,N_16593);
or U22968 (N_22968,N_17722,N_14657);
and U22969 (N_22969,N_13913,N_18432);
nand U22970 (N_22970,N_17673,N_17735);
and U22971 (N_22971,N_14433,N_13830);
and U22972 (N_22972,N_15687,N_14733);
nand U22973 (N_22973,N_14453,N_17500);
and U22974 (N_22974,N_17258,N_14746);
nand U22975 (N_22975,N_17657,N_15487);
nand U22976 (N_22976,N_12831,N_13136);
or U22977 (N_22977,N_15993,N_12919);
nor U22978 (N_22978,N_17824,N_17785);
nor U22979 (N_22979,N_15211,N_13121);
or U22980 (N_22980,N_14025,N_18420);
xor U22981 (N_22981,N_13629,N_12838);
xor U22982 (N_22982,N_15381,N_15451);
or U22983 (N_22983,N_16553,N_18132);
nand U22984 (N_22984,N_12535,N_12959);
or U22985 (N_22985,N_18396,N_14785);
and U22986 (N_22986,N_12731,N_13349);
nand U22987 (N_22987,N_17495,N_16260);
and U22988 (N_22988,N_15235,N_16247);
and U22989 (N_22989,N_17904,N_15776);
xor U22990 (N_22990,N_14247,N_15373);
and U22991 (N_22991,N_17229,N_18370);
nor U22992 (N_22992,N_17507,N_17388);
and U22993 (N_22993,N_13720,N_13618);
or U22994 (N_22994,N_15070,N_16119);
nor U22995 (N_22995,N_14516,N_16286);
nor U22996 (N_22996,N_15566,N_15375);
xnor U22997 (N_22997,N_16892,N_13958);
nor U22998 (N_22998,N_14947,N_16330);
and U22999 (N_22999,N_16516,N_13007);
or U23000 (N_23000,N_12746,N_17390);
nor U23001 (N_23001,N_12639,N_14133);
nand U23002 (N_23002,N_17385,N_17020);
nor U23003 (N_23003,N_16766,N_15428);
nand U23004 (N_23004,N_17867,N_17717);
or U23005 (N_23005,N_16035,N_16744);
nor U23006 (N_23006,N_17655,N_14948);
and U23007 (N_23007,N_16363,N_14902);
or U23008 (N_23008,N_14742,N_17215);
or U23009 (N_23009,N_17977,N_15529);
nor U23010 (N_23010,N_13077,N_14321);
or U23011 (N_23011,N_18235,N_12785);
and U23012 (N_23012,N_15717,N_13265);
nand U23013 (N_23013,N_15105,N_12752);
and U23014 (N_23014,N_18459,N_15522);
xnor U23015 (N_23015,N_14010,N_15352);
nand U23016 (N_23016,N_15314,N_15392);
nand U23017 (N_23017,N_16548,N_17083);
nor U23018 (N_23018,N_13061,N_14129);
or U23019 (N_23019,N_17008,N_13004);
nand U23020 (N_23020,N_15390,N_14720);
and U23021 (N_23021,N_16462,N_17491);
or U23022 (N_23022,N_16656,N_13016);
nand U23023 (N_23023,N_12901,N_14638);
xor U23024 (N_23024,N_17367,N_17181);
or U23025 (N_23025,N_16569,N_15667);
and U23026 (N_23026,N_16741,N_16983);
and U23027 (N_23027,N_13608,N_15627);
xor U23028 (N_23028,N_14732,N_15241);
nand U23029 (N_23029,N_18348,N_16041);
xnor U23030 (N_23030,N_17891,N_15249);
and U23031 (N_23031,N_15086,N_17904);
and U23032 (N_23032,N_16432,N_18669);
or U23033 (N_23033,N_17034,N_13708);
xor U23034 (N_23034,N_13635,N_16925);
xnor U23035 (N_23035,N_14723,N_17748);
or U23036 (N_23036,N_15709,N_15108);
or U23037 (N_23037,N_15498,N_17647);
nand U23038 (N_23038,N_18358,N_16060);
or U23039 (N_23039,N_15935,N_14141);
and U23040 (N_23040,N_15263,N_14734);
nand U23041 (N_23041,N_16381,N_14755);
nor U23042 (N_23042,N_16124,N_13071);
nor U23043 (N_23043,N_15758,N_15413);
nor U23044 (N_23044,N_15328,N_15998);
and U23045 (N_23045,N_18182,N_13898);
nor U23046 (N_23046,N_14026,N_13527);
nand U23047 (N_23047,N_14057,N_14431);
nor U23048 (N_23048,N_17886,N_18688);
and U23049 (N_23049,N_16469,N_13977);
or U23050 (N_23050,N_14212,N_12553);
nor U23051 (N_23051,N_16515,N_13888);
nor U23052 (N_23052,N_17248,N_15986);
xnor U23053 (N_23053,N_13583,N_13227);
nand U23054 (N_23054,N_13921,N_17775);
nand U23055 (N_23055,N_15510,N_17472);
xnor U23056 (N_23056,N_16628,N_14848);
nand U23057 (N_23057,N_18512,N_17666);
or U23058 (N_23058,N_16549,N_16561);
and U23059 (N_23059,N_17299,N_17838);
nor U23060 (N_23060,N_15043,N_17619);
nand U23061 (N_23061,N_14945,N_12914);
nor U23062 (N_23062,N_18409,N_13934);
and U23063 (N_23063,N_15153,N_16493);
nand U23064 (N_23064,N_16573,N_12952);
and U23065 (N_23065,N_18460,N_17407);
or U23066 (N_23066,N_13212,N_18410);
nand U23067 (N_23067,N_16669,N_17733);
and U23068 (N_23068,N_13403,N_16268);
nor U23069 (N_23069,N_13860,N_14387);
and U23070 (N_23070,N_15527,N_14958);
nor U23071 (N_23071,N_15461,N_16297);
and U23072 (N_23072,N_17494,N_15932);
nand U23073 (N_23073,N_13803,N_17381);
xor U23074 (N_23074,N_14591,N_14263);
nor U23075 (N_23075,N_15236,N_16501);
or U23076 (N_23076,N_15222,N_18402);
and U23077 (N_23077,N_13370,N_14922);
xnor U23078 (N_23078,N_13464,N_14285);
nor U23079 (N_23079,N_14252,N_15515);
xor U23080 (N_23080,N_17715,N_12585);
xnor U23081 (N_23081,N_14098,N_15426);
xnor U23082 (N_23082,N_13404,N_12555);
nand U23083 (N_23083,N_14128,N_16423);
and U23084 (N_23084,N_14387,N_16136);
nor U23085 (N_23085,N_16679,N_17751);
nor U23086 (N_23086,N_15204,N_14544);
and U23087 (N_23087,N_12925,N_18482);
xnor U23088 (N_23088,N_17157,N_14674);
xnor U23089 (N_23089,N_18531,N_18576);
nor U23090 (N_23090,N_18131,N_16319);
or U23091 (N_23091,N_14720,N_17678);
or U23092 (N_23092,N_18203,N_13030);
nand U23093 (N_23093,N_13508,N_15730);
or U23094 (N_23094,N_17857,N_16029);
and U23095 (N_23095,N_16067,N_17263);
and U23096 (N_23096,N_17645,N_18366);
nor U23097 (N_23097,N_16639,N_17309);
nor U23098 (N_23098,N_14337,N_18562);
or U23099 (N_23099,N_17845,N_14153);
nand U23100 (N_23100,N_15855,N_12907);
and U23101 (N_23101,N_15069,N_15404);
nor U23102 (N_23102,N_14356,N_14131);
xor U23103 (N_23103,N_12708,N_12841);
or U23104 (N_23104,N_16121,N_12638);
nand U23105 (N_23105,N_18234,N_13235);
nand U23106 (N_23106,N_13179,N_16626);
nor U23107 (N_23107,N_13494,N_15898);
nand U23108 (N_23108,N_12667,N_18066);
nand U23109 (N_23109,N_14464,N_18669);
or U23110 (N_23110,N_16085,N_14563);
or U23111 (N_23111,N_18203,N_12587);
nand U23112 (N_23112,N_14810,N_12512);
nand U23113 (N_23113,N_18316,N_16066);
or U23114 (N_23114,N_15980,N_15241);
nand U23115 (N_23115,N_12642,N_18612);
nor U23116 (N_23116,N_18439,N_16582);
nor U23117 (N_23117,N_13576,N_15937);
or U23118 (N_23118,N_14582,N_12730);
nor U23119 (N_23119,N_18355,N_16664);
nand U23120 (N_23120,N_14490,N_17720);
and U23121 (N_23121,N_15371,N_16754);
nand U23122 (N_23122,N_16807,N_17328);
xnor U23123 (N_23123,N_16442,N_14662);
or U23124 (N_23124,N_13654,N_13671);
xor U23125 (N_23125,N_17515,N_15284);
or U23126 (N_23126,N_14308,N_15640);
or U23127 (N_23127,N_15298,N_14743);
and U23128 (N_23128,N_17371,N_15363);
nand U23129 (N_23129,N_15390,N_14863);
and U23130 (N_23130,N_15715,N_14347);
or U23131 (N_23131,N_18671,N_13132);
and U23132 (N_23132,N_17368,N_17088);
or U23133 (N_23133,N_16291,N_17240);
xnor U23134 (N_23134,N_13542,N_15153);
xnor U23135 (N_23135,N_18052,N_15390);
xor U23136 (N_23136,N_18011,N_17174);
nand U23137 (N_23137,N_12764,N_18476);
nand U23138 (N_23138,N_15456,N_17760);
nor U23139 (N_23139,N_16566,N_16421);
nor U23140 (N_23140,N_16974,N_14581);
or U23141 (N_23141,N_16116,N_15986);
or U23142 (N_23142,N_15002,N_14040);
or U23143 (N_23143,N_15856,N_14252);
nand U23144 (N_23144,N_16061,N_17434);
nor U23145 (N_23145,N_16761,N_14555);
or U23146 (N_23146,N_16637,N_18009);
xor U23147 (N_23147,N_15778,N_15512);
xnor U23148 (N_23148,N_17434,N_15628);
or U23149 (N_23149,N_12882,N_12854);
and U23150 (N_23150,N_16973,N_18002);
nand U23151 (N_23151,N_15568,N_18625);
or U23152 (N_23152,N_18119,N_17195);
xnor U23153 (N_23153,N_17407,N_15968);
nor U23154 (N_23154,N_14284,N_12867);
and U23155 (N_23155,N_12786,N_13932);
nor U23156 (N_23156,N_17962,N_17582);
xor U23157 (N_23157,N_12787,N_15681);
nor U23158 (N_23158,N_12738,N_15535);
nand U23159 (N_23159,N_16216,N_18471);
nand U23160 (N_23160,N_14899,N_12501);
or U23161 (N_23161,N_15740,N_13495);
nor U23162 (N_23162,N_15157,N_12904);
and U23163 (N_23163,N_15056,N_16590);
xnor U23164 (N_23164,N_13551,N_12856);
or U23165 (N_23165,N_15037,N_16227);
nor U23166 (N_23166,N_12502,N_12946);
nor U23167 (N_23167,N_13836,N_13591);
nor U23168 (N_23168,N_17593,N_14711);
xor U23169 (N_23169,N_14238,N_17496);
or U23170 (N_23170,N_13257,N_13199);
nor U23171 (N_23171,N_13631,N_14299);
or U23172 (N_23172,N_14713,N_13637);
or U23173 (N_23173,N_15919,N_14759);
or U23174 (N_23174,N_18145,N_13006);
and U23175 (N_23175,N_16672,N_16099);
xor U23176 (N_23176,N_12756,N_16485);
and U23177 (N_23177,N_16526,N_13520);
or U23178 (N_23178,N_18529,N_14449);
xnor U23179 (N_23179,N_18552,N_16402);
nor U23180 (N_23180,N_16765,N_15940);
nor U23181 (N_23181,N_15422,N_13785);
and U23182 (N_23182,N_18123,N_12772);
xnor U23183 (N_23183,N_17491,N_14785);
or U23184 (N_23184,N_13755,N_15712);
nor U23185 (N_23185,N_17459,N_13211);
and U23186 (N_23186,N_12942,N_12925);
nor U23187 (N_23187,N_12922,N_16749);
nor U23188 (N_23188,N_16906,N_12876);
or U23189 (N_23189,N_14288,N_18150);
nor U23190 (N_23190,N_17573,N_13316);
xnor U23191 (N_23191,N_16585,N_13948);
nor U23192 (N_23192,N_17672,N_17535);
and U23193 (N_23193,N_14270,N_17038);
xor U23194 (N_23194,N_16713,N_14666);
and U23195 (N_23195,N_12815,N_14345);
xnor U23196 (N_23196,N_17196,N_14923);
or U23197 (N_23197,N_13448,N_13275);
nor U23198 (N_23198,N_17716,N_16847);
nand U23199 (N_23199,N_12704,N_13839);
nand U23200 (N_23200,N_12787,N_17423);
and U23201 (N_23201,N_15997,N_12540);
or U23202 (N_23202,N_17666,N_13235);
or U23203 (N_23203,N_15760,N_12798);
and U23204 (N_23204,N_14368,N_13632);
nor U23205 (N_23205,N_17994,N_18312);
nor U23206 (N_23206,N_18323,N_15439);
xor U23207 (N_23207,N_15204,N_13639);
nor U23208 (N_23208,N_13950,N_12554);
and U23209 (N_23209,N_16753,N_13148);
or U23210 (N_23210,N_18223,N_17119);
nor U23211 (N_23211,N_13357,N_16011);
and U23212 (N_23212,N_15418,N_13504);
xor U23213 (N_23213,N_14330,N_14956);
xnor U23214 (N_23214,N_13741,N_15192);
nor U23215 (N_23215,N_15349,N_18261);
or U23216 (N_23216,N_16920,N_13003);
nand U23217 (N_23217,N_17070,N_12912);
xor U23218 (N_23218,N_15777,N_12795);
xnor U23219 (N_23219,N_17673,N_15891);
xnor U23220 (N_23220,N_14711,N_17802);
nor U23221 (N_23221,N_14510,N_17940);
nand U23222 (N_23222,N_17926,N_12619);
or U23223 (N_23223,N_16395,N_17065);
nand U23224 (N_23224,N_17993,N_14138);
nor U23225 (N_23225,N_15557,N_12641);
nor U23226 (N_23226,N_14839,N_15387);
nor U23227 (N_23227,N_17642,N_17955);
nor U23228 (N_23228,N_14173,N_13097);
or U23229 (N_23229,N_18194,N_15690);
xor U23230 (N_23230,N_15171,N_14992);
or U23231 (N_23231,N_13599,N_16839);
and U23232 (N_23232,N_15874,N_13694);
nor U23233 (N_23233,N_16411,N_16244);
or U23234 (N_23234,N_14874,N_16644);
xor U23235 (N_23235,N_16944,N_16358);
nor U23236 (N_23236,N_18214,N_14671);
or U23237 (N_23237,N_17541,N_17445);
or U23238 (N_23238,N_18413,N_16619);
xor U23239 (N_23239,N_14861,N_17283);
nor U23240 (N_23240,N_14066,N_13583);
nor U23241 (N_23241,N_15622,N_16573);
nand U23242 (N_23242,N_13286,N_17461);
xor U23243 (N_23243,N_14730,N_14689);
nand U23244 (N_23244,N_13555,N_14646);
and U23245 (N_23245,N_16290,N_15344);
or U23246 (N_23246,N_15389,N_16526);
nor U23247 (N_23247,N_15668,N_14779);
and U23248 (N_23248,N_16905,N_14379);
nor U23249 (N_23249,N_14264,N_14568);
xor U23250 (N_23250,N_12701,N_12537);
or U23251 (N_23251,N_16151,N_13060);
and U23252 (N_23252,N_15828,N_14972);
nand U23253 (N_23253,N_16528,N_16810);
nor U23254 (N_23254,N_12881,N_14685);
xnor U23255 (N_23255,N_16364,N_13759);
or U23256 (N_23256,N_14570,N_15673);
and U23257 (N_23257,N_12760,N_15492);
or U23258 (N_23258,N_18648,N_12837);
or U23259 (N_23259,N_14700,N_18733);
xor U23260 (N_23260,N_15635,N_14798);
or U23261 (N_23261,N_18735,N_14587);
nor U23262 (N_23262,N_15834,N_16066);
and U23263 (N_23263,N_15071,N_17236);
nor U23264 (N_23264,N_12735,N_17645);
xnor U23265 (N_23265,N_18281,N_13205);
or U23266 (N_23266,N_18522,N_13300);
nor U23267 (N_23267,N_17703,N_17337);
xnor U23268 (N_23268,N_18685,N_15206);
nor U23269 (N_23269,N_17337,N_16026);
xor U23270 (N_23270,N_17771,N_15098);
nor U23271 (N_23271,N_14778,N_16825);
nor U23272 (N_23272,N_14366,N_14202);
nor U23273 (N_23273,N_17188,N_18659);
nand U23274 (N_23274,N_15047,N_12599);
nand U23275 (N_23275,N_18487,N_15966);
xnor U23276 (N_23276,N_17089,N_18142);
xor U23277 (N_23277,N_16872,N_18645);
nor U23278 (N_23278,N_18651,N_16982);
xnor U23279 (N_23279,N_14350,N_13815);
and U23280 (N_23280,N_16962,N_13939);
nand U23281 (N_23281,N_12685,N_14196);
xnor U23282 (N_23282,N_13903,N_13892);
nand U23283 (N_23283,N_15981,N_15419);
nor U23284 (N_23284,N_18317,N_15591);
or U23285 (N_23285,N_15216,N_17248);
nand U23286 (N_23286,N_15000,N_12559);
nor U23287 (N_23287,N_12597,N_14151);
or U23288 (N_23288,N_15708,N_14048);
and U23289 (N_23289,N_15536,N_17978);
nor U23290 (N_23290,N_17586,N_18600);
xor U23291 (N_23291,N_13878,N_17506);
nor U23292 (N_23292,N_12529,N_12830);
or U23293 (N_23293,N_17153,N_17044);
xnor U23294 (N_23294,N_15302,N_16440);
nand U23295 (N_23295,N_16195,N_14082);
nor U23296 (N_23296,N_17970,N_18610);
or U23297 (N_23297,N_17027,N_16419);
and U23298 (N_23298,N_16098,N_12780);
nor U23299 (N_23299,N_15017,N_18634);
nor U23300 (N_23300,N_13958,N_18441);
and U23301 (N_23301,N_12808,N_13300);
or U23302 (N_23302,N_16272,N_18036);
nand U23303 (N_23303,N_17215,N_14038);
nand U23304 (N_23304,N_16942,N_12934);
or U23305 (N_23305,N_18080,N_14215);
nor U23306 (N_23306,N_14383,N_17211);
or U23307 (N_23307,N_17536,N_17616);
or U23308 (N_23308,N_13260,N_15172);
nor U23309 (N_23309,N_12597,N_18621);
nand U23310 (N_23310,N_14640,N_13364);
or U23311 (N_23311,N_13307,N_12608);
xor U23312 (N_23312,N_15463,N_15470);
and U23313 (N_23313,N_17112,N_16379);
xnor U23314 (N_23314,N_15372,N_18123);
nand U23315 (N_23315,N_12572,N_18531);
or U23316 (N_23316,N_13957,N_17257);
nand U23317 (N_23317,N_14264,N_18419);
nand U23318 (N_23318,N_14498,N_17943);
xor U23319 (N_23319,N_16429,N_14340);
nand U23320 (N_23320,N_14620,N_16201);
xnor U23321 (N_23321,N_13991,N_13559);
nand U23322 (N_23322,N_15909,N_14780);
or U23323 (N_23323,N_14595,N_16533);
or U23324 (N_23324,N_14993,N_18304);
or U23325 (N_23325,N_13355,N_15534);
nand U23326 (N_23326,N_14191,N_13267);
xor U23327 (N_23327,N_16082,N_14216);
nor U23328 (N_23328,N_17400,N_14237);
and U23329 (N_23329,N_17421,N_13433);
and U23330 (N_23330,N_15176,N_12966);
nand U23331 (N_23331,N_18528,N_14948);
and U23332 (N_23332,N_15378,N_16047);
or U23333 (N_23333,N_16817,N_16265);
nand U23334 (N_23334,N_16096,N_18508);
xor U23335 (N_23335,N_13201,N_13947);
and U23336 (N_23336,N_15365,N_15656);
and U23337 (N_23337,N_12759,N_12806);
xnor U23338 (N_23338,N_16679,N_17769);
or U23339 (N_23339,N_12858,N_14665);
and U23340 (N_23340,N_15152,N_14491);
nand U23341 (N_23341,N_14720,N_18584);
nor U23342 (N_23342,N_13092,N_18446);
or U23343 (N_23343,N_13581,N_16525);
nor U23344 (N_23344,N_17910,N_16912);
or U23345 (N_23345,N_14114,N_12551);
xor U23346 (N_23346,N_16248,N_16010);
and U23347 (N_23347,N_18529,N_14102);
or U23348 (N_23348,N_13282,N_14045);
nor U23349 (N_23349,N_13775,N_17675);
nor U23350 (N_23350,N_15050,N_15949);
xnor U23351 (N_23351,N_16970,N_18178);
nand U23352 (N_23352,N_13912,N_13402);
nand U23353 (N_23353,N_16323,N_12922);
and U23354 (N_23354,N_15020,N_16217);
and U23355 (N_23355,N_13306,N_13515);
and U23356 (N_23356,N_15587,N_12993);
nand U23357 (N_23357,N_17725,N_14448);
and U23358 (N_23358,N_13223,N_15190);
xnor U23359 (N_23359,N_14505,N_15851);
or U23360 (N_23360,N_14999,N_15213);
nor U23361 (N_23361,N_16142,N_13383);
xor U23362 (N_23362,N_12677,N_15065);
nor U23363 (N_23363,N_15922,N_16882);
or U23364 (N_23364,N_14633,N_16322);
xor U23365 (N_23365,N_14906,N_12649);
nand U23366 (N_23366,N_15243,N_12661);
and U23367 (N_23367,N_17764,N_17716);
nand U23368 (N_23368,N_18727,N_18000);
nor U23369 (N_23369,N_16814,N_16862);
and U23370 (N_23370,N_13988,N_16484);
nor U23371 (N_23371,N_14243,N_17963);
xor U23372 (N_23372,N_14136,N_13624);
or U23373 (N_23373,N_17210,N_17164);
xnor U23374 (N_23374,N_13881,N_13515);
nor U23375 (N_23375,N_18563,N_16211);
nor U23376 (N_23376,N_14758,N_18277);
nor U23377 (N_23377,N_16097,N_15276);
and U23378 (N_23378,N_15769,N_12572);
xor U23379 (N_23379,N_16109,N_13666);
or U23380 (N_23380,N_15214,N_14279);
xor U23381 (N_23381,N_18161,N_14804);
and U23382 (N_23382,N_13597,N_18526);
nor U23383 (N_23383,N_12868,N_15293);
and U23384 (N_23384,N_13704,N_16723);
xor U23385 (N_23385,N_14754,N_13711);
nand U23386 (N_23386,N_18031,N_17669);
nand U23387 (N_23387,N_16604,N_13587);
nand U23388 (N_23388,N_13589,N_17793);
nor U23389 (N_23389,N_13856,N_15734);
and U23390 (N_23390,N_18050,N_13154);
or U23391 (N_23391,N_15152,N_18331);
and U23392 (N_23392,N_16094,N_17287);
nor U23393 (N_23393,N_16440,N_14598);
and U23394 (N_23394,N_17187,N_18232);
or U23395 (N_23395,N_14328,N_17122);
nor U23396 (N_23396,N_17456,N_15562);
or U23397 (N_23397,N_15401,N_14660);
and U23398 (N_23398,N_18368,N_16279);
and U23399 (N_23399,N_12681,N_13944);
nand U23400 (N_23400,N_14836,N_16121);
xor U23401 (N_23401,N_17327,N_17975);
nor U23402 (N_23402,N_18600,N_15609);
nor U23403 (N_23403,N_15599,N_13653);
or U23404 (N_23404,N_16703,N_17202);
nand U23405 (N_23405,N_15539,N_14328);
nand U23406 (N_23406,N_17856,N_14266);
nor U23407 (N_23407,N_15452,N_14624);
and U23408 (N_23408,N_17127,N_17800);
xor U23409 (N_23409,N_17653,N_13272);
nand U23410 (N_23410,N_14247,N_13880);
nor U23411 (N_23411,N_16610,N_17591);
nand U23412 (N_23412,N_13018,N_17095);
xnor U23413 (N_23413,N_17371,N_17612);
and U23414 (N_23414,N_13587,N_17025);
and U23415 (N_23415,N_17718,N_15509);
xnor U23416 (N_23416,N_13865,N_13814);
nand U23417 (N_23417,N_14592,N_17091);
nand U23418 (N_23418,N_15355,N_16237);
or U23419 (N_23419,N_16819,N_16457);
or U23420 (N_23420,N_17049,N_14326);
nor U23421 (N_23421,N_16443,N_14235);
xor U23422 (N_23422,N_16680,N_16144);
xnor U23423 (N_23423,N_14490,N_17394);
and U23424 (N_23424,N_12619,N_13001);
xnor U23425 (N_23425,N_16198,N_13286);
nor U23426 (N_23426,N_16634,N_13057);
and U23427 (N_23427,N_15911,N_16070);
nor U23428 (N_23428,N_16237,N_15375);
and U23429 (N_23429,N_13603,N_13527);
and U23430 (N_23430,N_15928,N_12939);
and U23431 (N_23431,N_15508,N_16568);
and U23432 (N_23432,N_13215,N_18318);
and U23433 (N_23433,N_13788,N_13494);
and U23434 (N_23434,N_17997,N_14565);
xnor U23435 (N_23435,N_18129,N_14917);
nand U23436 (N_23436,N_14499,N_13772);
or U23437 (N_23437,N_16340,N_17070);
and U23438 (N_23438,N_15361,N_14029);
nand U23439 (N_23439,N_13546,N_12571);
xnor U23440 (N_23440,N_15780,N_14112);
or U23441 (N_23441,N_13217,N_18638);
nor U23442 (N_23442,N_15438,N_16146);
nor U23443 (N_23443,N_17634,N_16878);
and U23444 (N_23444,N_14945,N_14433);
and U23445 (N_23445,N_16342,N_16212);
nand U23446 (N_23446,N_13656,N_17246);
nand U23447 (N_23447,N_14942,N_18136);
or U23448 (N_23448,N_17633,N_14859);
nand U23449 (N_23449,N_14492,N_14545);
and U23450 (N_23450,N_17734,N_18637);
nor U23451 (N_23451,N_15505,N_14999);
nand U23452 (N_23452,N_15503,N_16519);
or U23453 (N_23453,N_16944,N_13631);
or U23454 (N_23454,N_18415,N_15867);
nor U23455 (N_23455,N_13745,N_17220);
nand U23456 (N_23456,N_17551,N_15742);
nor U23457 (N_23457,N_14472,N_14065);
and U23458 (N_23458,N_13507,N_17956);
or U23459 (N_23459,N_17242,N_16869);
xor U23460 (N_23460,N_12698,N_17256);
and U23461 (N_23461,N_15674,N_15997);
nand U23462 (N_23462,N_18136,N_15584);
or U23463 (N_23463,N_15310,N_17478);
nand U23464 (N_23464,N_15116,N_18570);
nor U23465 (N_23465,N_14491,N_17049);
nand U23466 (N_23466,N_18174,N_16377);
nand U23467 (N_23467,N_17920,N_13707);
nand U23468 (N_23468,N_14129,N_15159);
nor U23469 (N_23469,N_15129,N_18608);
nand U23470 (N_23470,N_18596,N_15080);
nand U23471 (N_23471,N_18628,N_18178);
nand U23472 (N_23472,N_15120,N_16989);
and U23473 (N_23473,N_17661,N_16740);
nor U23474 (N_23474,N_15749,N_18697);
and U23475 (N_23475,N_14779,N_14280);
and U23476 (N_23476,N_16147,N_17005);
xor U23477 (N_23477,N_12776,N_13280);
nand U23478 (N_23478,N_14682,N_12632);
or U23479 (N_23479,N_17636,N_15185);
or U23480 (N_23480,N_14183,N_17362);
and U23481 (N_23481,N_18405,N_13861);
xnor U23482 (N_23482,N_12749,N_16913);
xnor U23483 (N_23483,N_18048,N_13942);
xor U23484 (N_23484,N_15475,N_18684);
nor U23485 (N_23485,N_14229,N_13498);
and U23486 (N_23486,N_14252,N_16081);
and U23487 (N_23487,N_15688,N_13511);
and U23488 (N_23488,N_12538,N_16154);
xor U23489 (N_23489,N_14294,N_13778);
xnor U23490 (N_23490,N_15528,N_18585);
nand U23491 (N_23491,N_18517,N_18470);
or U23492 (N_23492,N_16312,N_18372);
or U23493 (N_23493,N_13764,N_13429);
nor U23494 (N_23494,N_15152,N_14412);
nand U23495 (N_23495,N_17130,N_14176);
and U23496 (N_23496,N_14220,N_13071);
and U23497 (N_23497,N_14274,N_16454);
nor U23498 (N_23498,N_15751,N_17123);
or U23499 (N_23499,N_14193,N_15695);
xnor U23500 (N_23500,N_16533,N_13672);
and U23501 (N_23501,N_15156,N_14568);
or U23502 (N_23502,N_17495,N_18611);
and U23503 (N_23503,N_13887,N_15536);
or U23504 (N_23504,N_17598,N_18327);
nand U23505 (N_23505,N_14429,N_14160);
or U23506 (N_23506,N_12957,N_17064);
xor U23507 (N_23507,N_13943,N_16222);
or U23508 (N_23508,N_12795,N_17445);
xor U23509 (N_23509,N_15825,N_16821);
xnor U23510 (N_23510,N_13945,N_17093);
and U23511 (N_23511,N_15107,N_17525);
nand U23512 (N_23512,N_16999,N_16707);
nor U23513 (N_23513,N_16866,N_17958);
nor U23514 (N_23514,N_14021,N_18310);
or U23515 (N_23515,N_15514,N_18250);
and U23516 (N_23516,N_18588,N_18532);
or U23517 (N_23517,N_13069,N_16819);
and U23518 (N_23518,N_14382,N_13047);
or U23519 (N_23519,N_16920,N_17040);
xor U23520 (N_23520,N_16913,N_17103);
nor U23521 (N_23521,N_18446,N_15650);
nand U23522 (N_23522,N_16464,N_16034);
xor U23523 (N_23523,N_16221,N_16814);
and U23524 (N_23524,N_17883,N_13668);
xor U23525 (N_23525,N_14268,N_13548);
and U23526 (N_23526,N_13489,N_17788);
xor U23527 (N_23527,N_14553,N_17950);
or U23528 (N_23528,N_15122,N_17205);
nand U23529 (N_23529,N_13453,N_17912);
nand U23530 (N_23530,N_12587,N_13248);
nor U23531 (N_23531,N_16525,N_13807);
nand U23532 (N_23532,N_14356,N_16868);
nand U23533 (N_23533,N_15808,N_12746);
nor U23534 (N_23534,N_15212,N_17692);
xnor U23535 (N_23535,N_17025,N_17333);
nand U23536 (N_23536,N_17491,N_13722);
or U23537 (N_23537,N_14304,N_15341);
xor U23538 (N_23538,N_17823,N_16891);
xor U23539 (N_23539,N_13856,N_15331);
xnor U23540 (N_23540,N_13064,N_14532);
or U23541 (N_23541,N_13731,N_14916);
and U23542 (N_23542,N_14048,N_13907);
or U23543 (N_23543,N_16588,N_17170);
nor U23544 (N_23544,N_16740,N_15663);
or U23545 (N_23545,N_15788,N_16348);
xor U23546 (N_23546,N_18139,N_15576);
nand U23547 (N_23547,N_14020,N_14257);
nor U23548 (N_23548,N_13693,N_17905);
or U23549 (N_23549,N_16934,N_17980);
nor U23550 (N_23550,N_16138,N_14304);
and U23551 (N_23551,N_14446,N_14715);
nor U23552 (N_23552,N_15528,N_13052);
or U23553 (N_23553,N_17452,N_17145);
or U23554 (N_23554,N_13725,N_17419);
nor U23555 (N_23555,N_14156,N_14971);
nand U23556 (N_23556,N_18243,N_15046);
xor U23557 (N_23557,N_16001,N_13855);
xnor U23558 (N_23558,N_12863,N_17751);
nand U23559 (N_23559,N_18575,N_14596);
nor U23560 (N_23560,N_13206,N_12988);
or U23561 (N_23561,N_16828,N_18294);
or U23562 (N_23562,N_15926,N_13305);
nand U23563 (N_23563,N_17791,N_16140);
and U23564 (N_23564,N_15817,N_15176);
and U23565 (N_23565,N_17831,N_18581);
and U23566 (N_23566,N_17598,N_16462);
nand U23567 (N_23567,N_14189,N_18024);
or U23568 (N_23568,N_13352,N_18042);
xnor U23569 (N_23569,N_15603,N_18199);
and U23570 (N_23570,N_12807,N_13126);
nand U23571 (N_23571,N_15665,N_15016);
nor U23572 (N_23572,N_15503,N_13098);
nand U23573 (N_23573,N_14310,N_15833);
nand U23574 (N_23574,N_12597,N_16787);
or U23575 (N_23575,N_12829,N_14598);
nand U23576 (N_23576,N_15355,N_12546);
nand U23577 (N_23577,N_13994,N_16322);
xor U23578 (N_23578,N_13484,N_18424);
or U23579 (N_23579,N_16580,N_14695);
nor U23580 (N_23580,N_18034,N_18308);
nor U23581 (N_23581,N_17042,N_17876);
and U23582 (N_23582,N_14438,N_18187);
nand U23583 (N_23583,N_13948,N_13674);
or U23584 (N_23584,N_18157,N_16464);
nand U23585 (N_23585,N_16812,N_15909);
nor U23586 (N_23586,N_15621,N_15864);
or U23587 (N_23587,N_17826,N_14881);
nor U23588 (N_23588,N_15006,N_17216);
nand U23589 (N_23589,N_15548,N_12641);
and U23590 (N_23590,N_15801,N_18082);
xor U23591 (N_23591,N_16871,N_18698);
nand U23592 (N_23592,N_18152,N_13926);
xnor U23593 (N_23593,N_18741,N_14627);
xor U23594 (N_23594,N_14054,N_15229);
nand U23595 (N_23595,N_14430,N_18250);
and U23596 (N_23596,N_16228,N_13238);
or U23597 (N_23597,N_16943,N_18604);
and U23598 (N_23598,N_13615,N_12884);
and U23599 (N_23599,N_18540,N_15530);
nand U23600 (N_23600,N_13101,N_15797);
nor U23601 (N_23601,N_15411,N_18728);
or U23602 (N_23602,N_17177,N_17477);
xnor U23603 (N_23603,N_12613,N_18718);
nor U23604 (N_23604,N_12552,N_16738);
or U23605 (N_23605,N_17798,N_14170);
and U23606 (N_23606,N_12837,N_15041);
xor U23607 (N_23607,N_17195,N_16907);
xnor U23608 (N_23608,N_16868,N_16007);
or U23609 (N_23609,N_17882,N_16414);
nor U23610 (N_23610,N_16827,N_18644);
nor U23611 (N_23611,N_14704,N_13645);
nor U23612 (N_23612,N_17659,N_14947);
nand U23613 (N_23613,N_17213,N_16725);
nand U23614 (N_23614,N_15661,N_14105);
xnor U23615 (N_23615,N_12659,N_14697);
xnor U23616 (N_23616,N_18489,N_16409);
xnor U23617 (N_23617,N_12676,N_13408);
and U23618 (N_23618,N_15971,N_17445);
and U23619 (N_23619,N_13824,N_18529);
xnor U23620 (N_23620,N_16883,N_12610);
or U23621 (N_23621,N_15413,N_17083);
nand U23622 (N_23622,N_17924,N_12988);
or U23623 (N_23623,N_16452,N_16345);
nor U23624 (N_23624,N_14212,N_17414);
nor U23625 (N_23625,N_18669,N_14450);
xnor U23626 (N_23626,N_15476,N_14739);
nand U23627 (N_23627,N_16251,N_17120);
nand U23628 (N_23628,N_13506,N_12551);
or U23629 (N_23629,N_17763,N_18100);
or U23630 (N_23630,N_16637,N_17187);
and U23631 (N_23631,N_13223,N_14192);
or U23632 (N_23632,N_16453,N_15499);
xnor U23633 (N_23633,N_13564,N_16369);
xor U23634 (N_23634,N_17151,N_13816);
or U23635 (N_23635,N_17414,N_16273);
nand U23636 (N_23636,N_18101,N_18741);
and U23637 (N_23637,N_17146,N_13993);
nand U23638 (N_23638,N_14865,N_16239);
xor U23639 (N_23639,N_13575,N_15106);
and U23640 (N_23640,N_17687,N_18743);
nor U23641 (N_23641,N_17963,N_15559);
nor U23642 (N_23642,N_15054,N_13443);
and U23643 (N_23643,N_13175,N_18346);
nand U23644 (N_23644,N_13722,N_18337);
or U23645 (N_23645,N_17348,N_14395);
nor U23646 (N_23646,N_15743,N_17234);
nand U23647 (N_23647,N_16412,N_18539);
and U23648 (N_23648,N_16542,N_16379);
or U23649 (N_23649,N_16521,N_13116);
nor U23650 (N_23650,N_16044,N_14025);
xor U23651 (N_23651,N_15690,N_13329);
and U23652 (N_23652,N_14420,N_17807);
or U23653 (N_23653,N_17098,N_15360);
and U23654 (N_23654,N_18545,N_15994);
xor U23655 (N_23655,N_14508,N_14319);
and U23656 (N_23656,N_14156,N_12914);
or U23657 (N_23657,N_17051,N_14107);
nand U23658 (N_23658,N_15019,N_17640);
nand U23659 (N_23659,N_12958,N_16966);
nand U23660 (N_23660,N_13633,N_16662);
or U23661 (N_23661,N_13802,N_14532);
xnor U23662 (N_23662,N_16286,N_17898);
and U23663 (N_23663,N_14842,N_14379);
or U23664 (N_23664,N_12508,N_13665);
xnor U23665 (N_23665,N_14428,N_14744);
or U23666 (N_23666,N_15508,N_17601);
and U23667 (N_23667,N_18401,N_15259);
or U23668 (N_23668,N_17011,N_15109);
xor U23669 (N_23669,N_14927,N_18080);
or U23670 (N_23670,N_13205,N_17170);
or U23671 (N_23671,N_15394,N_15171);
and U23672 (N_23672,N_17562,N_14866);
xor U23673 (N_23673,N_18637,N_15966);
nor U23674 (N_23674,N_18339,N_13465);
and U23675 (N_23675,N_15840,N_17954);
xnor U23676 (N_23676,N_17946,N_14426);
or U23677 (N_23677,N_18093,N_18327);
or U23678 (N_23678,N_12544,N_17146);
or U23679 (N_23679,N_15217,N_15681);
nor U23680 (N_23680,N_17367,N_13189);
xor U23681 (N_23681,N_15188,N_18635);
or U23682 (N_23682,N_15227,N_16759);
nor U23683 (N_23683,N_16782,N_16065);
xor U23684 (N_23684,N_14013,N_13632);
or U23685 (N_23685,N_12961,N_18236);
and U23686 (N_23686,N_15939,N_14823);
or U23687 (N_23687,N_14506,N_12901);
xor U23688 (N_23688,N_18380,N_14524);
nor U23689 (N_23689,N_18570,N_16838);
and U23690 (N_23690,N_17363,N_12765);
xnor U23691 (N_23691,N_14815,N_18610);
xor U23692 (N_23692,N_15136,N_16227);
xnor U23693 (N_23693,N_14043,N_18102);
xnor U23694 (N_23694,N_18482,N_17409);
or U23695 (N_23695,N_18440,N_16340);
nor U23696 (N_23696,N_14988,N_15842);
nor U23697 (N_23697,N_17051,N_13482);
nand U23698 (N_23698,N_13570,N_14771);
xor U23699 (N_23699,N_17166,N_12907);
and U23700 (N_23700,N_17734,N_18728);
nor U23701 (N_23701,N_12579,N_18348);
or U23702 (N_23702,N_17288,N_15837);
and U23703 (N_23703,N_17132,N_14844);
and U23704 (N_23704,N_14425,N_12790);
xnor U23705 (N_23705,N_12533,N_18067);
nand U23706 (N_23706,N_17472,N_13876);
and U23707 (N_23707,N_14706,N_18434);
and U23708 (N_23708,N_18423,N_16553);
nor U23709 (N_23709,N_16049,N_16402);
or U23710 (N_23710,N_14401,N_13288);
nand U23711 (N_23711,N_14922,N_16439);
nor U23712 (N_23712,N_12908,N_15582);
or U23713 (N_23713,N_15519,N_16552);
or U23714 (N_23714,N_12952,N_14743);
nor U23715 (N_23715,N_13323,N_13421);
and U23716 (N_23716,N_15842,N_14324);
xor U23717 (N_23717,N_18399,N_12920);
or U23718 (N_23718,N_18076,N_15467);
nor U23719 (N_23719,N_14181,N_12760);
and U23720 (N_23720,N_15532,N_16775);
xor U23721 (N_23721,N_14652,N_13413);
xnor U23722 (N_23722,N_12702,N_14366);
nand U23723 (N_23723,N_15984,N_17833);
nand U23724 (N_23724,N_14275,N_13927);
nor U23725 (N_23725,N_16219,N_17592);
and U23726 (N_23726,N_17863,N_18273);
nor U23727 (N_23727,N_17966,N_16193);
nor U23728 (N_23728,N_13445,N_13547);
nand U23729 (N_23729,N_18007,N_15378);
xnor U23730 (N_23730,N_17455,N_17678);
xnor U23731 (N_23731,N_16527,N_16242);
and U23732 (N_23732,N_12744,N_13552);
nor U23733 (N_23733,N_14071,N_17802);
and U23734 (N_23734,N_13646,N_17120);
and U23735 (N_23735,N_17207,N_16435);
nand U23736 (N_23736,N_18055,N_16142);
and U23737 (N_23737,N_15326,N_15081);
or U23738 (N_23738,N_14302,N_14642);
nor U23739 (N_23739,N_13643,N_16870);
xor U23740 (N_23740,N_15183,N_15749);
xnor U23741 (N_23741,N_15596,N_17108);
nor U23742 (N_23742,N_13031,N_16164);
or U23743 (N_23743,N_17912,N_15785);
nor U23744 (N_23744,N_16563,N_16203);
and U23745 (N_23745,N_17810,N_18095);
or U23746 (N_23746,N_15171,N_16652);
nor U23747 (N_23747,N_14017,N_14774);
nor U23748 (N_23748,N_14149,N_17488);
or U23749 (N_23749,N_12960,N_18516);
and U23750 (N_23750,N_14749,N_12785);
nor U23751 (N_23751,N_13441,N_17683);
xor U23752 (N_23752,N_17010,N_14167);
or U23753 (N_23753,N_13107,N_14941);
xnor U23754 (N_23754,N_15654,N_18116);
nand U23755 (N_23755,N_18627,N_15429);
nor U23756 (N_23756,N_12544,N_16480);
xor U23757 (N_23757,N_17707,N_14367);
nor U23758 (N_23758,N_15670,N_15666);
nor U23759 (N_23759,N_14161,N_12833);
and U23760 (N_23760,N_16673,N_14494);
xnor U23761 (N_23761,N_15604,N_12900);
xnor U23762 (N_23762,N_16298,N_13594);
nand U23763 (N_23763,N_14838,N_17926);
xor U23764 (N_23764,N_13926,N_13220);
xor U23765 (N_23765,N_17047,N_15843);
xnor U23766 (N_23766,N_14156,N_18246);
nor U23767 (N_23767,N_16868,N_15449);
or U23768 (N_23768,N_14946,N_16211);
and U23769 (N_23769,N_15970,N_14918);
and U23770 (N_23770,N_16101,N_12901);
and U23771 (N_23771,N_15032,N_12669);
or U23772 (N_23772,N_14767,N_18133);
xor U23773 (N_23773,N_12534,N_13909);
xor U23774 (N_23774,N_15126,N_16865);
and U23775 (N_23775,N_18614,N_16659);
xnor U23776 (N_23776,N_14085,N_13178);
or U23777 (N_23777,N_16698,N_14125);
nor U23778 (N_23778,N_17010,N_14299);
nor U23779 (N_23779,N_17872,N_17017);
nand U23780 (N_23780,N_18088,N_13023);
or U23781 (N_23781,N_12566,N_15078);
xor U23782 (N_23782,N_13112,N_14474);
nand U23783 (N_23783,N_17238,N_13560);
or U23784 (N_23784,N_14001,N_17210);
and U23785 (N_23785,N_16430,N_13628);
and U23786 (N_23786,N_13601,N_18616);
or U23787 (N_23787,N_16136,N_17327);
and U23788 (N_23788,N_16187,N_13767);
nor U23789 (N_23789,N_18458,N_17304);
or U23790 (N_23790,N_14078,N_15988);
and U23791 (N_23791,N_13727,N_17187);
nor U23792 (N_23792,N_18687,N_16426);
and U23793 (N_23793,N_14936,N_17842);
nor U23794 (N_23794,N_13718,N_17168);
nand U23795 (N_23795,N_13771,N_18224);
nand U23796 (N_23796,N_14851,N_13045);
and U23797 (N_23797,N_16526,N_17492);
or U23798 (N_23798,N_14320,N_13795);
and U23799 (N_23799,N_13870,N_18395);
xor U23800 (N_23800,N_16218,N_17087);
or U23801 (N_23801,N_15799,N_17455);
nor U23802 (N_23802,N_14931,N_16990);
nand U23803 (N_23803,N_14327,N_18196);
xor U23804 (N_23804,N_18260,N_14192);
nand U23805 (N_23805,N_17192,N_16751);
nor U23806 (N_23806,N_13010,N_13232);
nor U23807 (N_23807,N_13162,N_16513);
and U23808 (N_23808,N_14808,N_17250);
or U23809 (N_23809,N_17525,N_14645);
or U23810 (N_23810,N_17184,N_13628);
and U23811 (N_23811,N_13630,N_14004);
and U23812 (N_23812,N_17198,N_14992);
nor U23813 (N_23813,N_15093,N_18622);
or U23814 (N_23814,N_15428,N_17108);
nand U23815 (N_23815,N_15188,N_12955);
nor U23816 (N_23816,N_15002,N_14640);
and U23817 (N_23817,N_16663,N_14122);
or U23818 (N_23818,N_14017,N_14495);
and U23819 (N_23819,N_14136,N_15127);
or U23820 (N_23820,N_13755,N_12795);
nand U23821 (N_23821,N_18610,N_15391);
nor U23822 (N_23822,N_16218,N_13668);
nor U23823 (N_23823,N_14498,N_18658);
nor U23824 (N_23824,N_16456,N_15271);
nand U23825 (N_23825,N_15917,N_18424);
or U23826 (N_23826,N_16447,N_15181);
nand U23827 (N_23827,N_16687,N_15233);
and U23828 (N_23828,N_16876,N_15565);
or U23829 (N_23829,N_17136,N_15272);
or U23830 (N_23830,N_14486,N_18201);
nand U23831 (N_23831,N_12979,N_16794);
and U23832 (N_23832,N_13548,N_18326);
nor U23833 (N_23833,N_16602,N_14585);
xor U23834 (N_23834,N_16706,N_13964);
nand U23835 (N_23835,N_13448,N_18661);
and U23836 (N_23836,N_16023,N_13799);
or U23837 (N_23837,N_17555,N_17521);
xor U23838 (N_23838,N_14102,N_14924);
or U23839 (N_23839,N_17994,N_17026);
nor U23840 (N_23840,N_14978,N_12979);
xnor U23841 (N_23841,N_15922,N_18371);
nand U23842 (N_23842,N_17588,N_18224);
and U23843 (N_23843,N_13953,N_18185);
nor U23844 (N_23844,N_16358,N_16739);
and U23845 (N_23845,N_18394,N_14079);
or U23846 (N_23846,N_14063,N_15212);
nand U23847 (N_23847,N_15697,N_13031);
nand U23848 (N_23848,N_14342,N_14413);
nor U23849 (N_23849,N_16483,N_13468);
nand U23850 (N_23850,N_16581,N_12921);
and U23851 (N_23851,N_14648,N_14161);
xor U23852 (N_23852,N_15573,N_14242);
xnor U23853 (N_23853,N_17386,N_14236);
nor U23854 (N_23854,N_18075,N_15406);
nor U23855 (N_23855,N_16419,N_14922);
xnor U23856 (N_23856,N_15383,N_14077);
xor U23857 (N_23857,N_17923,N_16378);
nor U23858 (N_23858,N_13857,N_13355);
and U23859 (N_23859,N_14314,N_15193);
nor U23860 (N_23860,N_18475,N_16759);
or U23861 (N_23861,N_17138,N_15423);
or U23862 (N_23862,N_14911,N_14470);
nand U23863 (N_23863,N_14980,N_15766);
nand U23864 (N_23864,N_16409,N_17853);
xor U23865 (N_23865,N_15485,N_14156);
and U23866 (N_23866,N_12713,N_16610);
xnor U23867 (N_23867,N_16743,N_13361);
nor U23868 (N_23868,N_13344,N_14969);
and U23869 (N_23869,N_15631,N_13978);
xor U23870 (N_23870,N_16347,N_17769);
nor U23871 (N_23871,N_17885,N_14208);
xnor U23872 (N_23872,N_16278,N_13057);
nand U23873 (N_23873,N_16459,N_15849);
xnor U23874 (N_23874,N_13674,N_18017);
or U23875 (N_23875,N_13434,N_16510);
xor U23876 (N_23876,N_13223,N_13390);
and U23877 (N_23877,N_13734,N_18647);
and U23878 (N_23878,N_17565,N_13033);
or U23879 (N_23879,N_18099,N_13467);
xnor U23880 (N_23880,N_12557,N_16230);
or U23881 (N_23881,N_12824,N_13798);
nor U23882 (N_23882,N_15682,N_12513);
and U23883 (N_23883,N_16486,N_14568);
or U23884 (N_23884,N_16853,N_13811);
nand U23885 (N_23885,N_12615,N_17009);
nand U23886 (N_23886,N_17646,N_13779);
nand U23887 (N_23887,N_13586,N_16982);
nor U23888 (N_23888,N_16818,N_15891);
or U23889 (N_23889,N_12909,N_17175);
xnor U23890 (N_23890,N_13924,N_15876);
and U23891 (N_23891,N_16148,N_12926);
nand U23892 (N_23892,N_16979,N_17270);
nand U23893 (N_23893,N_14026,N_18214);
and U23894 (N_23894,N_12679,N_13345);
and U23895 (N_23895,N_15330,N_12781);
or U23896 (N_23896,N_17146,N_13533);
or U23897 (N_23897,N_16435,N_16983);
nand U23898 (N_23898,N_16312,N_12813);
nand U23899 (N_23899,N_17659,N_17207);
and U23900 (N_23900,N_13122,N_17636);
xor U23901 (N_23901,N_14651,N_17547);
nor U23902 (N_23902,N_13510,N_15978);
or U23903 (N_23903,N_13519,N_14497);
xor U23904 (N_23904,N_13218,N_14241);
and U23905 (N_23905,N_17128,N_13599);
nand U23906 (N_23906,N_16135,N_13611);
xor U23907 (N_23907,N_15893,N_16494);
or U23908 (N_23908,N_12601,N_13653);
or U23909 (N_23909,N_16036,N_17510);
xor U23910 (N_23910,N_15140,N_18701);
xor U23911 (N_23911,N_13114,N_16483);
nand U23912 (N_23912,N_17439,N_13686);
or U23913 (N_23913,N_14967,N_16499);
xor U23914 (N_23914,N_14993,N_15378);
or U23915 (N_23915,N_12698,N_13033);
nand U23916 (N_23916,N_18593,N_14240);
xnor U23917 (N_23917,N_13858,N_14539);
or U23918 (N_23918,N_15853,N_14414);
nor U23919 (N_23919,N_18454,N_16533);
and U23920 (N_23920,N_17762,N_13012);
or U23921 (N_23921,N_15576,N_16093);
or U23922 (N_23922,N_14166,N_14878);
nor U23923 (N_23923,N_16329,N_14005);
or U23924 (N_23924,N_16048,N_14064);
nand U23925 (N_23925,N_18030,N_15558);
xnor U23926 (N_23926,N_15903,N_14387);
nand U23927 (N_23927,N_14713,N_17504);
and U23928 (N_23928,N_13025,N_16554);
and U23929 (N_23929,N_14535,N_14184);
nor U23930 (N_23930,N_13939,N_16898);
or U23931 (N_23931,N_12681,N_18143);
xnor U23932 (N_23932,N_18167,N_17736);
xor U23933 (N_23933,N_13465,N_16765);
and U23934 (N_23934,N_16446,N_15620);
nand U23935 (N_23935,N_15037,N_13121);
or U23936 (N_23936,N_13758,N_15811);
nand U23937 (N_23937,N_14840,N_16785);
or U23938 (N_23938,N_18366,N_14671);
xor U23939 (N_23939,N_18290,N_15303);
nor U23940 (N_23940,N_13431,N_13919);
nand U23941 (N_23941,N_17256,N_18031);
xor U23942 (N_23942,N_14025,N_14531);
xnor U23943 (N_23943,N_14718,N_13893);
nand U23944 (N_23944,N_17803,N_15416);
xnor U23945 (N_23945,N_13108,N_15891);
nor U23946 (N_23946,N_17022,N_16724);
and U23947 (N_23947,N_18276,N_16839);
and U23948 (N_23948,N_17993,N_16649);
nor U23949 (N_23949,N_18184,N_16913);
or U23950 (N_23950,N_13029,N_14229);
xor U23951 (N_23951,N_13326,N_13061);
nand U23952 (N_23952,N_13515,N_14489);
xor U23953 (N_23953,N_12933,N_17480);
and U23954 (N_23954,N_18339,N_13369);
and U23955 (N_23955,N_17372,N_16910);
nor U23956 (N_23956,N_16296,N_17961);
xnor U23957 (N_23957,N_13640,N_17048);
nor U23958 (N_23958,N_12845,N_13509);
nor U23959 (N_23959,N_17266,N_16702);
or U23960 (N_23960,N_13649,N_12804);
nand U23961 (N_23961,N_18039,N_16756);
nand U23962 (N_23962,N_12841,N_14245);
and U23963 (N_23963,N_12908,N_12737);
nand U23964 (N_23964,N_15933,N_14419);
or U23965 (N_23965,N_15439,N_14345);
or U23966 (N_23966,N_12892,N_13339);
nor U23967 (N_23967,N_13810,N_15240);
nor U23968 (N_23968,N_18016,N_18338);
nand U23969 (N_23969,N_12876,N_15424);
and U23970 (N_23970,N_18335,N_12642);
or U23971 (N_23971,N_14663,N_13803);
and U23972 (N_23972,N_12510,N_15737);
nor U23973 (N_23973,N_17408,N_13068);
nand U23974 (N_23974,N_16338,N_17761);
and U23975 (N_23975,N_12707,N_14103);
and U23976 (N_23976,N_16519,N_13107);
nand U23977 (N_23977,N_15499,N_15488);
xor U23978 (N_23978,N_17684,N_14415);
nand U23979 (N_23979,N_14539,N_14598);
nor U23980 (N_23980,N_16861,N_16284);
nand U23981 (N_23981,N_13716,N_13203);
xnor U23982 (N_23982,N_15028,N_15324);
or U23983 (N_23983,N_12685,N_12665);
and U23984 (N_23984,N_13522,N_14595);
xor U23985 (N_23985,N_17302,N_15828);
xnor U23986 (N_23986,N_13973,N_14256);
nor U23987 (N_23987,N_15281,N_18732);
xor U23988 (N_23988,N_17118,N_14592);
xnor U23989 (N_23989,N_14343,N_12511);
xor U23990 (N_23990,N_14052,N_14095);
nor U23991 (N_23991,N_15561,N_14403);
nor U23992 (N_23992,N_17963,N_13846);
or U23993 (N_23993,N_13891,N_18406);
xnor U23994 (N_23994,N_12722,N_14290);
xnor U23995 (N_23995,N_18110,N_15441);
or U23996 (N_23996,N_18187,N_12954);
and U23997 (N_23997,N_14434,N_13008);
or U23998 (N_23998,N_12646,N_15727);
and U23999 (N_23999,N_13773,N_15228);
xor U24000 (N_24000,N_18531,N_14242);
nand U24001 (N_24001,N_16746,N_15223);
xnor U24002 (N_24002,N_16023,N_17750);
or U24003 (N_24003,N_12740,N_14135);
nor U24004 (N_24004,N_17548,N_14346);
and U24005 (N_24005,N_18028,N_16205);
nor U24006 (N_24006,N_15554,N_16026);
nand U24007 (N_24007,N_16160,N_15421);
nor U24008 (N_24008,N_15020,N_16621);
or U24009 (N_24009,N_15016,N_14756);
nand U24010 (N_24010,N_14662,N_13706);
nand U24011 (N_24011,N_12681,N_13402);
and U24012 (N_24012,N_18323,N_13030);
and U24013 (N_24013,N_16698,N_16874);
or U24014 (N_24014,N_17651,N_15006);
nand U24015 (N_24015,N_17475,N_14610);
xor U24016 (N_24016,N_14526,N_15407);
xor U24017 (N_24017,N_18636,N_14111);
or U24018 (N_24018,N_15721,N_17408);
and U24019 (N_24019,N_15320,N_15900);
nand U24020 (N_24020,N_13324,N_17587);
nand U24021 (N_24021,N_12553,N_13770);
xor U24022 (N_24022,N_13476,N_18288);
nand U24023 (N_24023,N_14676,N_18477);
nand U24024 (N_24024,N_15563,N_14068);
nand U24025 (N_24025,N_18106,N_13170);
or U24026 (N_24026,N_12787,N_18025);
or U24027 (N_24027,N_14609,N_15457);
nand U24028 (N_24028,N_14391,N_18540);
and U24029 (N_24029,N_17493,N_18395);
and U24030 (N_24030,N_16808,N_14735);
nor U24031 (N_24031,N_14137,N_17878);
xor U24032 (N_24032,N_12840,N_17077);
nand U24033 (N_24033,N_14727,N_12553);
nand U24034 (N_24034,N_13200,N_14297);
xor U24035 (N_24035,N_17095,N_13479);
xor U24036 (N_24036,N_14753,N_17533);
and U24037 (N_24037,N_16017,N_16666);
and U24038 (N_24038,N_15996,N_18574);
nor U24039 (N_24039,N_16057,N_14048);
xnor U24040 (N_24040,N_14467,N_14148);
xor U24041 (N_24041,N_15425,N_18313);
nor U24042 (N_24042,N_17434,N_18430);
or U24043 (N_24043,N_13635,N_13518);
xor U24044 (N_24044,N_16125,N_15412);
or U24045 (N_24045,N_16369,N_17962);
nand U24046 (N_24046,N_17461,N_14518);
nor U24047 (N_24047,N_16942,N_15152);
and U24048 (N_24048,N_14776,N_15807);
nor U24049 (N_24049,N_15285,N_14065);
xnor U24050 (N_24050,N_16375,N_14179);
xor U24051 (N_24051,N_15124,N_18307);
xnor U24052 (N_24052,N_18269,N_14323);
and U24053 (N_24053,N_15333,N_15805);
nand U24054 (N_24054,N_14861,N_16214);
nand U24055 (N_24055,N_14596,N_16860);
nor U24056 (N_24056,N_15433,N_13182);
and U24057 (N_24057,N_14507,N_17760);
nor U24058 (N_24058,N_17944,N_13600);
nand U24059 (N_24059,N_13236,N_15599);
and U24060 (N_24060,N_13911,N_15502);
nand U24061 (N_24061,N_18051,N_16071);
nor U24062 (N_24062,N_15511,N_13891);
and U24063 (N_24063,N_16775,N_17416);
xor U24064 (N_24064,N_12799,N_16641);
or U24065 (N_24065,N_16230,N_13343);
or U24066 (N_24066,N_14144,N_18689);
or U24067 (N_24067,N_18309,N_15601);
nor U24068 (N_24068,N_17347,N_18682);
nor U24069 (N_24069,N_16894,N_16546);
nor U24070 (N_24070,N_18232,N_13373);
xor U24071 (N_24071,N_16604,N_15799);
and U24072 (N_24072,N_13591,N_18098);
xnor U24073 (N_24073,N_17702,N_13428);
or U24074 (N_24074,N_13495,N_16225);
xnor U24075 (N_24075,N_14462,N_17651);
nand U24076 (N_24076,N_13758,N_13331);
nand U24077 (N_24077,N_15165,N_16204);
and U24078 (N_24078,N_18292,N_14075);
or U24079 (N_24079,N_18287,N_18396);
nor U24080 (N_24080,N_16238,N_18166);
nand U24081 (N_24081,N_14144,N_14768);
and U24082 (N_24082,N_16506,N_16774);
xor U24083 (N_24083,N_14003,N_16288);
or U24084 (N_24084,N_14824,N_15248);
nor U24085 (N_24085,N_15219,N_18236);
nand U24086 (N_24086,N_14748,N_17057);
xnor U24087 (N_24087,N_15833,N_15602);
nor U24088 (N_24088,N_14705,N_16126);
or U24089 (N_24089,N_18599,N_16645);
and U24090 (N_24090,N_14002,N_13979);
or U24091 (N_24091,N_18351,N_13935);
xnor U24092 (N_24092,N_15455,N_15631);
nand U24093 (N_24093,N_13542,N_16323);
xnor U24094 (N_24094,N_13060,N_15657);
xnor U24095 (N_24095,N_18556,N_14181);
nand U24096 (N_24096,N_13768,N_12715);
or U24097 (N_24097,N_16893,N_14916);
and U24098 (N_24098,N_16769,N_13541);
nor U24099 (N_24099,N_14425,N_16637);
and U24100 (N_24100,N_17235,N_17963);
or U24101 (N_24101,N_17635,N_13806);
nand U24102 (N_24102,N_18020,N_18617);
xnor U24103 (N_24103,N_13466,N_16018);
or U24104 (N_24104,N_18546,N_17341);
xnor U24105 (N_24105,N_13078,N_15898);
nor U24106 (N_24106,N_18699,N_17316);
nor U24107 (N_24107,N_13454,N_15204);
xnor U24108 (N_24108,N_12724,N_18146);
or U24109 (N_24109,N_15871,N_16695);
or U24110 (N_24110,N_14921,N_15858);
and U24111 (N_24111,N_17027,N_15613);
nand U24112 (N_24112,N_13706,N_17052);
xor U24113 (N_24113,N_17087,N_13137);
or U24114 (N_24114,N_14554,N_15411);
and U24115 (N_24115,N_16069,N_16631);
nand U24116 (N_24116,N_14662,N_12829);
or U24117 (N_24117,N_15187,N_17665);
nor U24118 (N_24118,N_14592,N_18069);
xnor U24119 (N_24119,N_14291,N_14511);
nand U24120 (N_24120,N_17464,N_13516);
xor U24121 (N_24121,N_17526,N_17554);
xor U24122 (N_24122,N_14730,N_18438);
and U24123 (N_24123,N_14929,N_14700);
nand U24124 (N_24124,N_14991,N_18315);
nor U24125 (N_24125,N_18348,N_15316);
nor U24126 (N_24126,N_15489,N_17605);
and U24127 (N_24127,N_12623,N_18209);
nor U24128 (N_24128,N_17671,N_14211);
or U24129 (N_24129,N_17277,N_14703);
nand U24130 (N_24130,N_17705,N_13202);
or U24131 (N_24131,N_18636,N_14989);
and U24132 (N_24132,N_12800,N_17885);
or U24133 (N_24133,N_15041,N_16089);
and U24134 (N_24134,N_15830,N_13410);
nand U24135 (N_24135,N_14256,N_15521);
and U24136 (N_24136,N_13479,N_15851);
nand U24137 (N_24137,N_13729,N_16441);
nand U24138 (N_24138,N_15482,N_17000);
nor U24139 (N_24139,N_18055,N_13096);
nor U24140 (N_24140,N_12838,N_18590);
xor U24141 (N_24141,N_13123,N_15909);
or U24142 (N_24142,N_15099,N_13637);
nor U24143 (N_24143,N_16180,N_14432);
nand U24144 (N_24144,N_14010,N_17727);
and U24145 (N_24145,N_12618,N_18141);
nor U24146 (N_24146,N_15079,N_16355);
and U24147 (N_24147,N_18336,N_15926);
nor U24148 (N_24148,N_17928,N_16685);
nor U24149 (N_24149,N_17335,N_14615);
xnor U24150 (N_24150,N_17537,N_14053);
and U24151 (N_24151,N_16787,N_17481);
or U24152 (N_24152,N_18022,N_16297);
nor U24153 (N_24153,N_15121,N_18618);
xnor U24154 (N_24154,N_15161,N_15169);
nand U24155 (N_24155,N_16484,N_17155);
xor U24156 (N_24156,N_17156,N_16297);
or U24157 (N_24157,N_18191,N_13468);
nand U24158 (N_24158,N_13579,N_15775);
xnor U24159 (N_24159,N_13400,N_16997);
and U24160 (N_24160,N_13345,N_18561);
and U24161 (N_24161,N_16007,N_13919);
and U24162 (N_24162,N_12686,N_17120);
or U24163 (N_24163,N_14348,N_14003);
nor U24164 (N_24164,N_15488,N_15788);
nand U24165 (N_24165,N_17939,N_15392);
xor U24166 (N_24166,N_17650,N_18391);
and U24167 (N_24167,N_12935,N_17884);
nand U24168 (N_24168,N_15801,N_13038);
nand U24169 (N_24169,N_17569,N_14210);
or U24170 (N_24170,N_18218,N_13377);
xnor U24171 (N_24171,N_13704,N_13948);
nor U24172 (N_24172,N_13092,N_18369);
xnor U24173 (N_24173,N_15477,N_13418);
nor U24174 (N_24174,N_13855,N_14047);
xnor U24175 (N_24175,N_15042,N_13544);
and U24176 (N_24176,N_14681,N_16300);
or U24177 (N_24177,N_13525,N_14391);
nor U24178 (N_24178,N_13102,N_14586);
nand U24179 (N_24179,N_18027,N_12656);
xnor U24180 (N_24180,N_17946,N_18149);
and U24181 (N_24181,N_16135,N_16599);
or U24182 (N_24182,N_13166,N_14064);
or U24183 (N_24183,N_17231,N_17672);
nand U24184 (N_24184,N_16427,N_16266);
nor U24185 (N_24185,N_16820,N_13767);
and U24186 (N_24186,N_13799,N_14423);
or U24187 (N_24187,N_16367,N_17502);
or U24188 (N_24188,N_12531,N_16747);
or U24189 (N_24189,N_17378,N_16782);
nor U24190 (N_24190,N_14130,N_17366);
or U24191 (N_24191,N_16128,N_18071);
xnor U24192 (N_24192,N_17020,N_14626);
nand U24193 (N_24193,N_17540,N_15062);
nand U24194 (N_24194,N_15542,N_18346);
xor U24195 (N_24195,N_18516,N_13536);
or U24196 (N_24196,N_13740,N_14400);
nor U24197 (N_24197,N_13079,N_18324);
xor U24198 (N_24198,N_16117,N_13999);
nand U24199 (N_24199,N_18198,N_18087);
xnor U24200 (N_24200,N_18299,N_16300);
nor U24201 (N_24201,N_16546,N_16441);
and U24202 (N_24202,N_15715,N_17565);
xnor U24203 (N_24203,N_14518,N_16063);
or U24204 (N_24204,N_12867,N_13896);
nor U24205 (N_24205,N_14626,N_17102);
nand U24206 (N_24206,N_18552,N_17455);
nor U24207 (N_24207,N_13570,N_13747);
and U24208 (N_24208,N_13230,N_16155);
xor U24209 (N_24209,N_15874,N_14547);
xnor U24210 (N_24210,N_17838,N_14055);
and U24211 (N_24211,N_15475,N_17713);
nor U24212 (N_24212,N_14336,N_12706);
xnor U24213 (N_24213,N_15052,N_17627);
and U24214 (N_24214,N_18013,N_15449);
and U24215 (N_24215,N_13348,N_13812);
nand U24216 (N_24216,N_14397,N_13849);
nor U24217 (N_24217,N_18267,N_15975);
nor U24218 (N_24218,N_16060,N_12681);
nor U24219 (N_24219,N_13578,N_13375);
nor U24220 (N_24220,N_17411,N_14473);
or U24221 (N_24221,N_18277,N_16316);
nor U24222 (N_24222,N_13614,N_17641);
nand U24223 (N_24223,N_17228,N_13245);
xnor U24224 (N_24224,N_18712,N_15973);
or U24225 (N_24225,N_16933,N_13987);
or U24226 (N_24226,N_14141,N_17714);
or U24227 (N_24227,N_17873,N_15584);
xnor U24228 (N_24228,N_15829,N_15562);
nor U24229 (N_24229,N_15307,N_12568);
xnor U24230 (N_24230,N_14844,N_14596);
xnor U24231 (N_24231,N_13618,N_12783);
nor U24232 (N_24232,N_13062,N_18566);
xnor U24233 (N_24233,N_16217,N_16052);
or U24234 (N_24234,N_18161,N_15394);
xor U24235 (N_24235,N_14958,N_18462);
xor U24236 (N_24236,N_13102,N_14482);
nor U24237 (N_24237,N_15509,N_13930);
and U24238 (N_24238,N_16482,N_12706);
nand U24239 (N_24239,N_13579,N_18638);
nor U24240 (N_24240,N_14614,N_16167);
and U24241 (N_24241,N_12508,N_13871);
and U24242 (N_24242,N_14437,N_15059);
and U24243 (N_24243,N_16599,N_12880);
and U24244 (N_24244,N_17771,N_14734);
nand U24245 (N_24245,N_17808,N_16948);
nor U24246 (N_24246,N_15971,N_15061);
or U24247 (N_24247,N_15295,N_15192);
and U24248 (N_24248,N_13937,N_18426);
nor U24249 (N_24249,N_16545,N_15627);
nand U24250 (N_24250,N_13046,N_17661);
nor U24251 (N_24251,N_14888,N_15736);
nor U24252 (N_24252,N_13565,N_16435);
and U24253 (N_24253,N_15931,N_13386);
and U24254 (N_24254,N_16388,N_17979);
nor U24255 (N_24255,N_15492,N_15080);
or U24256 (N_24256,N_15590,N_14358);
nand U24257 (N_24257,N_13927,N_13515);
xnor U24258 (N_24258,N_13861,N_16517);
nor U24259 (N_24259,N_17670,N_13548);
xnor U24260 (N_24260,N_15388,N_13303);
and U24261 (N_24261,N_14027,N_17739);
xor U24262 (N_24262,N_14107,N_14621);
xor U24263 (N_24263,N_18312,N_16756);
nand U24264 (N_24264,N_13144,N_17311);
xnor U24265 (N_24265,N_18682,N_18188);
nor U24266 (N_24266,N_13787,N_13104);
xor U24267 (N_24267,N_13363,N_14920);
and U24268 (N_24268,N_14464,N_14257);
nand U24269 (N_24269,N_18202,N_16328);
nand U24270 (N_24270,N_13533,N_15704);
nand U24271 (N_24271,N_16287,N_16309);
or U24272 (N_24272,N_17287,N_14453);
and U24273 (N_24273,N_16983,N_14160);
nor U24274 (N_24274,N_12591,N_16788);
or U24275 (N_24275,N_14214,N_16472);
nor U24276 (N_24276,N_15445,N_15911);
or U24277 (N_24277,N_12658,N_14905);
xor U24278 (N_24278,N_15864,N_13361);
nor U24279 (N_24279,N_16716,N_17232);
or U24280 (N_24280,N_17157,N_16003);
nor U24281 (N_24281,N_15116,N_15319);
nand U24282 (N_24282,N_16260,N_18238);
and U24283 (N_24283,N_14285,N_17698);
nor U24284 (N_24284,N_13832,N_17547);
and U24285 (N_24285,N_18045,N_16602);
nor U24286 (N_24286,N_17486,N_15939);
xor U24287 (N_24287,N_18469,N_14798);
nand U24288 (N_24288,N_13177,N_13221);
nor U24289 (N_24289,N_13645,N_16476);
and U24290 (N_24290,N_16788,N_14967);
nand U24291 (N_24291,N_14800,N_13462);
nand U24292 (N_24292,N_14226,N_15807);
and U24293 (N_24293,N_17835,N_12610);
or U24294 (N_24294,N_13813,N_17033);
or U24295 (N_24295,N_16692,N_18333);
nand U24296 (N_24296,N_17211,N_18649);
nand U24297 (N_24297,N_15153,N_16450);
xnor U24298 (N_24298,N_16983,N_13508);
or U24299 (N_24299,N_15502,N_16195);
or U24300 (N_24300,N_13203,N_15403);
xor U24301 (N_24301,N_17478,N_12772);
nor U24302 (N_24302,N_17088,N_16840);
nand U24303 (N_24303,N_13273,N_14353);
nand U24304 (N_24304,N_16296,N_16455);
nand U24305 (N_24305,N_14879,N_18217);
and U24306 (N_24306,N_15142,N_13522);
or U24307 (N_24307,N_16380,N_16306);
nand U24308 (N_24308,N_12863,N_18374);
xor U24309 (N_24309,N_12728,N_14267);
or U24310 (N_24310,N_13829,N_18250);
nor U24311 (N_24311,N_16027,N_14099);
and U24312 (N_24312,N_17449,N_15485);
nand U24313 (N_24313,N_12526,N_18416);
nor U24314 (N_24314,N_16391,N_14277);
or U24315 (N_24315,N_18066,N_16677);
nand U24316 (N_24316,N_17152,N_13944);
nor U24317 (N_24317,N_16185,N_13286);
or U24318 (N_24318,N_17213,N_18158);
nand U24319 (N_24319,N_15197,N_18311);
xnor U24320 (N_24320,N_13394,N_13859);
and U24321 (N_24321,N_18264,N_15997);
xor U24322 (N_24322,N_16725,N_15915);
nor U24323 (N_24323,N_18010,N_18033);
and U24324 (N_24324,N_12765,N_14996);
nor U24325 (N_24325,N_17178,N_15889);
or U24326 (N_24326,N_17628,N_13414);
nor U24327 (N_24327,N_15902,N_13094);
xnor U24328 (N_24328,N_16450,N_12847);
nand U24329 (N_24329,N_17925,N_15591);
nor U24330 (N_24330,N_17796,N_12568);
nand U24331 (N_24331,N_15012,N_18124);
nand U24332 (N_24332,N_14745,N_12524);
nor U24333 (N_24333,N_16068,N_16960);
or U24334 (N_24334,N_18688,N_16598);
or U24335 (N_24335,N_16381,N_16780);
or U24336 (N_24336,N_14492,N_16680);
nand U24337 (N_24337,N_17497,N_14496);
xnor U24338 (N_24338,N_14697,N_16285);
and U24339 (N_24339,N_18073,N_16793);
nand U24340 (N_24340,N_15656,N_14731);
and U24341 (N_24341,N_18372,N_12709);
or U24342 (N_24342,N_14890,N_15030);
and U24343 (N_24343,N_16816,N_14450);
xor U24344 (N_24344,N_15629,N_13452);
xnor U24345 (N_24345,N_13383,N_15774);
xnor U24346 (N_24346,N_18075,N_17992);
nor U24347 (N_24347,N_12909,N_15461);
or U24348 (N_24348,N_14241,N_13635);
nand U24349 (N_24349,N_16800,N_16579);
xnor U24350 (N_24350,N_15828,N_14971);
nor U24351 (N_24351,N_17661,N_15542);
nor U24352 (N_24352,N_14549,N_14136);
nand U24353 (N_24353,N_15847,N_16437);
and U24354 (N_24354,N_14542,N_14789);
or U24355 (N_24355,N_18203,N_16537);
nor U24356 (N_24356,N_18159,N_16446);
nor U24357 (N_24357,N_18227,N_15691);
or U24358 (N_24358,N_17544,N_17091);
or U24359 (N_24359,N_14119,N_13529);
or U24360 (N_24360,N_15321,N_16447);
xor U24361 (N_24361,N_13092,N_13653);
and U24362 (N_24362,N_12551,N_15199);
xnor U24363 (N_24363,N_15627,N_15316);
xnor U24364 (N_24364,N_14843,N_15323);
nor U24365 (N_24365,N_16975,N_15730);
nand U24366 (N_24366,N_17313,N_18366);
nand U24367 (N_24367,N_13213,N_18004);
xnor U24368 (N_24368,N_15226,N_13004);
nor U24369 (N_24369,N_16920,N_16763);
or U24370 (N_24370,N_13311,N_16300);
and U24371 (N_24371,N_14938,N_12854);
or U24372 (N_24372,N_17471,N_17123);
or U24373 (N_24373,N_16297,N_15242);
nor U24374 (N_24374,N_18655,N_17649);
xor U24375 (N_24375,N_16707,N_16779);
or U24376 (N_24376,N_15034,N_14378);
and U24377 (N_24377,N_12974,N_15487);
and U24378 (N_24378,N_15123,N_16313);
xor U24379 (N_24379,N_17781,N_16140);
nand U24380 (N_24380,N_13167,N_16884);
nor U24381 (N_24381,N_17492,N_18642);
xnor U24382 (N_24382,N_12948,N_18332);
xnor U24383 (N_24383,N_16923,N_17651);
and U24384 (N_24384,N_14476,N_18145);
and U24385 (N_24385,N_17395,N_14743);
and U24386 (N_24386,N_14806,N_13511);
or U24387 (N_24387,N_14113,N_14872);
nand U24388 (N_24388,N_18320,N_16943);
xnor U24389 (N_24389,N_13124,N_15378);
xor U24390 (N_24390,N_15219,N_15610);
or U24391 (N_24391,N_13242,N_12614);
and U24392 (N_24392,N_15366,N_17389);
nand U24393 (N_24393,N_15914,N_15053);
and U24394 (N_24394,N_14917,N_16993);
or U24395 (N_24395,N_16954,N_15098);
or U24396 (N_24396,N_15071,N_18471);
xnor U24397 (N_24397,N_12679,N_18244);
nor U24398 (N_24398,N_18457,N_18285);
or U24399 (N_24399,N_18598,N_15688);
and U24400 (N_24400,N_17762,N_16147);
xor U24401 (N_24401,N_15461,N_14039);
nor U24402 (N_24402,N_15068,N_13004);
or U24403 (N_24403,N_15661,N_16446);
nand U24404 (N_24404,N_12696,N_14821);
or U24405 (N_24405,N_16053,N_12616);
or U24406 (N_24406,N_17554,N_13905);
nor U24407 (N_24407,N_17855,N_17595);
or U24408 (N_24408,N_18703,N_18156);
nor U24409 (N_24409,N_18319,N_16872);
xnor U24410 (N_24410,N_17418,N_13331);
xor U24411 (N_24411,N_15251,N_13718);
nor U24412 (N_24412,N_14652,N_12838);
nand U24413 (N_24413,N_14259,N_15248);
and U24414 (N_24414,N_15802,N_14735);
or U24415 (N_24415,N_18696,N_16737);
or U24416 (N_24416,N_14289,N_15494);
nor U24417 (N_24417,N_13777,N_16850);
nand U24418 (N_24418,N_15646,N_18023);
and U24419 (N_24419,N_12896,N_17085);
or U24420 (N_24420,N_16874,N_14605);
nor U24421 (N_24421,N_17730,N_15267);
xnor U24422 (N_24422,N_18408,N_18410);
xor U24423 (N_24423,N_14853,N_13203);
nor U24424 (N_24424,N_18717,N_17552);
and U24425 (N_24425,N_12873,N_13685);
nand U24426 (N_24426,N_15618,N_16063);
and U24427 (N_24427,N_12975,N_13619);
nand U24428 (N_24428,N_14808,N_12924);
xnor U24429 (N_24429,N_16166,N_16078);
xnor U24430 (N_24430,N_13265,N_13032);
xnor U24431 (N_24431,N_16391,N_15276);
xnor U24432 (N_24432,N_15141,N_17753);
nand U24433 (N_24433,N_18129,N_12878);
or U24434 (N_24434,N_12636,N_17659);
and U24435 (N_24435,N_17773,N_13529);
nand U24436 (N_24436,N_15581,N_18261);
nand U24437 (N_24437,N_18074,N_15059);
or U24438 (N_24438,N_16539,N_16275);
or U24439 (N_24439,N_13469,N_14643);
nor U24440 (N_24440,N_13766,N_15457);
xnor U24441 (N_24441,N_14151,N_15768);
xor U24442 (N_24442,N_16037,N_14659);
nor U24443 (N_24443,N_13228,N_14790);
or U24444 (N_24444,N_17427,N_16417);
nor U24445 (N_24445,N_12667,N_15569);
xor U24446 (N_24446,N_16775,N_15965);
nor U24447 (N_24447,N_18278,N_13236);
xnor U24448 (N_24448,N_16851,N_17608);
nand U24449 (N_24449,N_18741,N_13769);
or U24450 (N_24450,N_17695,N_13273);
xnor U24451 (N_24451,N_18218,N_15512);
xnor U24452 (N_24452,N_13730,N_15014);
xor U24453 (N_24453,N_18557,N_16845);
nand U24454 (N_24454,N_15508,N_15939);
nor U24455 (N_24455,N_15562,N_15887);
nand U24456 (N_24456,N_13155,N_15831);
or U24457 (N_24457,N_16727,N_14192);
or U24458 (N_24458,N_13696,N_15980);
nand U24459 (N_24459,N_13891,N_14753);
and U24460 (N_24460,N_13438,N_12672);
nor U24461 (N_24461,N_15658,N_16205);
or U24462 (N_24462,N_15295,N_14340);
nand U24463 (N_24463,N_17926,N_17106);
xor U24464 (N_24464,N_18407,N_17417);
nor U24465 (N_24465,N_15369,N_17935);
and U24466 (N_24466,N_15580,N_16754);
nor U24467 (N_24467,N_16447,N_13835);
nor U24468 (N_24468,N_14710,N_14239);
or U24469 (N_24469,N_14454,N_17524);
and U24470 (N_24470,N_13522,N_13475);
and U24471 (N_24471,N_12510,N_12661);
nand U24472 (N_24472,N_14482,N_17938);
and U24473 (N_24473,N_16599,N_16288);
or U24474 (N_24474,N_15730,N_16254);
xor U24475 (N_24475,N_17293,N_14390);
xnor U24476 (N_24476,N_13288,N_13223);
xor U24477 (N_24477,N_15802,N_15166);
and U24478 (N_24478,N_14848,N_17786);
and U24479 (N_24479,N_16743,N_17286);
xor U24480 (N_24480,N_14523,N_16234);
nor U24481 (N_24481,N_13323,N_17319);
xor U24482 (N_24482,N_17330,N_16516);
nor U24483 (N_24483,N_13386,N_16499);
or U24484 (N_24484,N_15167,N_15379);
xor U24485 (N_24485,N_14216,N_14491);
and U24486 (N_24486,N_17978,N_14006);
nor U24487 (N_24487,N_16604,N_17468);
and U24488 (N_24488,N_14002,N_15433);
xnor U24489 (N_24489,N_16495,N_14520);
nand U24490 (N_24490,N_14705,N_18279);
nor U24491 (N_24491,N_14060,N_12797);
and U24492 (N_24492,N_13743,N_15617);
nor U24493 (N_24493,N_14404,N_17930);
xor U24494 (N_24494,N_15011,N_18639);
or U24495 (N_24495,N_13931,N_17784);
xnor U24496 (N_24496,N_16201,N_13984);
nor U24497 (N_24497,N_14928,N_13003);
or U24498 (N_24498,N_15719,N_15387);
nand U24499 (N_24499,N_17021,N_18055);
nand U24500 (N_24500,N_14571,N_14877);
nand U24501 (N_24501,N_16098,N_18554);
nand U24502 (N_24502,N_18432,N_15844);
and U24503 (N_24503,N_15269,N_18686);
xor U24504 (N_24504,N_17971,N_13356);
xor U24505 (N_24505,N_14979,N_16937);
or U24506 (N_24506,N_17136,N_16973);
nand U24507 (N_24507,N_15026,N_13662);
xnor U24508 (N_24508,N_17895,N_15726);
or U24509 (N_24509,N_15025,N_18375);
nand U24510 (N_24510,N_14296,N_16856);
xnor U24511 (N_24511,N_17791,N_18739);
nor U24512 (N_24512,N_14034,N_15597);
or U24513 (N_24513,N_12548,N_14760);
or U24514 (N_24514,N_17915,N_17799);
and U24515 (N_24515,N_15943,N_16603);
or U24516 (N_24516,N_18710,N_17317);
nor U24517 (N_24517,N_15114,N_16838);
nor U24518 (N_24518,N_14429,N_12962);
or U24519 (N_24519,N_18712,N_13413);
nor U24520 (N_24520,N_18135,N_16683);
nand U24521 (N_24521,N_15563,N_16493);
and U24522 (N_24522,N_12708,N_14225);
nor U24523 (N_24523,N_16631,N_16879);
nor U24524 (N_24524,N_18645,N_14499);
xor U24525 (N_24525,N_13028,N_14857);
or U24526 (N_24526,N_17085,N_13755);
and U24527 (N_24527,N_17915,N_15139);
and U24528 (N_24528,N_16434,N_16559);
nand U24529 (N_24529,N_17229,N_15000);
nand U24530 (N_24530,N_13912,N_18490);
nand U24531 (N_24531,N_14513,N_14333);
or U24532 (N_24532,N_17946,N_14537);
nand U24533 (N_24533,N_16600,N_12744);
and U24534 (N_24534,N_15257,N_15038);
nand U24535 (N_24535,N_17898,N_16468);
nor U24536 (N_24536,N_18567,N_14786);
and U24537 (N_24537,N_14739,N_16733);
and U24538 (N_24538,N_15841,N_14443);
nor U24539 (N_24539,N_13908,N_18162);
nand U24540 (N_24540,N_15118,N_15528);
or U24541 (N_24541,N_12727,N_12836);
xor U24542 (N_24542,N_14357,N_17349);
and U24543 (N_24543,N_16368,N_15645);
nand U24544 (N_24544,N_18368,N_15009);
nand U24545 (N_24545,N_14408,N_17830);
nor U24546 (N_24546,N_12687,N_13123);
nand U24547 (N_24547,N_12827,N_13481);
or U24548 (N_24548,N_12909,N_13877);
and U24549 (N_24549,N_12983,N_16316);
and U24550 (N_24550,N_18629,N_15666);
nor U24551 (N_24551,N_15845,N_14288);
or U24552 (N_24552,N_18649,N_13314);
nand U24553 (N_24553,N_13616,N_16214);
nor U24554 (N_24554,N_14967,N_17937);
nand U24555 (N_24555,N_14169,N_17955);
and U24556 (N_24556,N_14174,N_15065);
xnor U24557 (N_24557,N_16150,N_17585);
nand U24558 (N_24558,N_17692,N_16308);
or U24559 (N_24559,N_13716,N_13688);
or U24560 (N_24560,N_18529,N_13992);
or U24561 (N_24561,N_14550,N_16190);
nand U24562 (N_24562,N_16994,N_13409);
and U24563 (N_24563,N_14025,N_12856);
xnor U24564 (N_24564,N_15498,N_15256);
or U24565 (N_24565,N_17050,N_17252);
or U24566 (N_24566,N_13675,N_12981);
and U24567 (N_24567,N_14188,N_14292);
nor U24568 (N_24568,N_15852,N_13692);
nand U24569 (N_24569,N_15054,N_16705);
or U24570 (N_24570,N_16793,N_13445);
or U24571 (N_24571,N_16114,N_12952);
or U24572 (N_24572,N_14805,N_14996);
xor U24573 (N_24573,N_12656,N_13805);
and U24574 (N_24574,N_13674,N_15632);
xor U24575 (N_24575,N_18545,N_13728);
and U24576 (N_24576,N_12924,N_15059);
nand U24577 (N_24577,N_17285,N_13955);
xnor U24578 (N_24578,N_13525,N_13429);
xor U24579 (N_24579,N_14559,N_12665);
nor U24580 (N_24580,N_14974,N_15886);
nor U24581 (N_24581,N_13329,N_18558);
nor U24582 (N_24582,N_13728,N_14515);
xor U24583 (N_24583,N_16036,N_17569);
nand U24584 (N_24584,N_17514,N_18164);
and U24585 (N_24585,N_14862,N_16325);
nor U24586 (N_24586,N_15916,N_16599);
xor U24587 (N_24587,N_17623,N_16445);
and U24588 (N_24588,N_15962,N_15705);
and U24589 (N_24589,N_16046,N_12793);
and U24590 (N_24590,N_17055,N_15966);
or U24591 (N_24591,N_16462,N_15917);
nand U24592 (N_24592,N_13759,N_14224);
or U24593 (N_24593,N_13823,N_14941);
or U24594 (N_24594,N_16068,N_16852);
xnor U24595 (N_24595,N_17267,N_18627);
nand U24596 (N_24596,N_16659,N_18682);
and U24597 (N_24597,N_15732,N_14166);
xnor U24598 (N_24598,N_12536,N_18142);
or U24599 (N_24599,N_17218,N_13230);
nor U24600 (N_24600,N_18477,N_15925);
xnor U24601 (N_24601,N_13281,N_13880);
nand U24602 (N_24602,N_17212,N_13311);
and U24603 (N_24603,N_13905,N_18037);
or U24604 (N_24604,N_15495,N_14901);
nand U24605 (N_24605,N_13030,N_17141);
or U24606 (N_24606,N_18055,N_17780);
nand U24607 (N_24607,N_14766,N_13223);
xor U24608 (N_24608,N_14528,N_15668);
nand U24609 (N_24609,N_13063,N_18638);
or U24610 (N_24610,N_17827,N_18441);
xnor U24611 (N_24611,N_14268,N_14005);
nand U24612 (N_24612,N_16316,N_13233);
nand U24613 (N_24613,N_15381,N_15440);
nor U24614 (N_24614,N_14270,N_13755);
nand U24615 (N_24615,N_17286,N_13976);
or U24616 (N_24616,N_12960,N_13171);
and U24617 (N_24617,N_16307,N_13284);
nor U24618 (N_24618,N_12630,N_12519);
and U24619 (N_24619,N_12945,N_18692);
nor U24620 (N_24620,N_13664,N_16195);
nor U24621 (N_24621,N_15545,N_13264);
nand U24622 (N_24622,N_16517,N_15065);
and U24623 (N_24623,N_17414,N_18334);
or U24624 (N_24624,N_16250,N_16612);
and U24625 (N_24625,N_18085,N_15749);
xor U24626 (N_24626,N_16602,N_12585);
or U24627 (N_24627,N_17219,N_14395);
nor U24628 (N_24628,N_16791,N_13344);
or U24629 (N_24629,N_15589,N_16157);
and U24630 (N_24630,N_15350,N_16081);
nand U24631 (N_24631,N_15375,N_17455);
or U24632 (N_24632,N_13666,N_13906);
and U24633 (N_24633,N_15400,N_16280);
and U24634 (N_24634,N_13688,N_15302);
nand U24635 (N_24635,N_12764,N_16470);
or U24636 (N_24636,N_18650,N_16908);
nor U24637 (N_24637,N_17381,N_12921);
nor U24638 (N_24638,N_15569,N_18431);
and U24639 (N_24639,N_16872,N_13937);
and U24640 (N_24640,N_13995,N_12829);
or U24641 (N_24641,N_16668,N_16459);
nor U24642 (N_24642,N_18007,N_14074);
and U24643 (N_24643,N_14475,N_12973);
nand U24644 (N_24644,N_14439,N_13518);
nand U24645 (N_24645,N_14599,N_12595);
xnor U24646 (N_24646,N_14639,N_14068);
nand U24647 (N_24647,N_12580,N_16404);
and U24648 (N_24648,N_18711,N_18495);
xor U24649 (N_24649,N_16476,N_14234);
or U24650 (N_24650,N_13091,N_14581);
and U24651 (N_24651,N_17665,N_16707);
xnor U24652 (N_24652,N_12606,N_15433);
or U24653 (N_24653,N_14495,N_18641);
xor U24654 (N_24654,N_17890,N_18612);
and U24655 (N_24655,N_15305,N_15715);
xnor U24656 (N_24656,N_18708,N_15688);
or U24657 (N_24657,N_14668,N_15476);
nand U24658 (N_24658,N_16872,N_15282);
or U24659 (N_24659,N_17442,N_17094);
nand U24660 (N_24660,N_13467,N_18108);
nor U24661 (N_24661,N_16176,N_16656);
and U24662 (N_24662,N_13600,N_15950);
and U24663 (N_24663,N_12844,N_13457);
and U24664 (N_24664,N_15367,N_15249);
and U24665 (N_24665,N_14871,N_17793);
or U24666 (N_24666,N_17171,N_13203);
nand U24667 (N_24667,N_12937,N_14484);
xnor U24668 (N_24668,N_17380,N_14214);
nand U24669 (N_24669,N_13178,N_17056);
and U24670 (N_24670,N_17348,N_17385);
nand U24671 (N_24671,N_17677,N_16614);
and U24672 (N_24672,N_17259,N_16995);
or U24673 (N_24673,N_17918,N_13024);
nor U24674 (N_24674,N_15924,N_17496);
xor U24675 (N_24675,N_13596,N_18032);
xnor U24676 (N_24676,N_17028,N_13821);
and U24677 (N_24677,N_13513,N_16293);
nor U24678 (N_24678,N_12621,N_15342);
or U24679 (N_24679,N_13839,N_14704);
and U24680 (N_24680,N_18014,N_17333);
xor U24681 (N_24681,N_17593,N_12799);
xor U24682 (N_24682,N_18486,N_14519);
nand U24683 (N_24683,N_17540,N_12994);
xnor U24684 (N_24684,N_13155,N_16605);
xnor U24685 (N_24685,N_16126,N_15240);
nand U24686 (N_24686,N_17998,N_15358);
xnor U24687 (N_24687,N_17059,N_13239);
or U24688 (N_24688,N_16345,N_16853);
and U24689 (N_24689,N_13548,N_14475);
xnor U24690 (N_24690,N_14343,N_17992);
or U24691 (N_24691,N_15162,N_15436);
and U24692 (N_24692,N_16375,N_14964);
or U24693 (N_24693,N_14501,N_17546);
nand U24694 (N_24694,N_13195,N_14561);
and U24695 (N_24695,N_18600,N_15606);
or U24696 (N_24696,N_14599,N_17511);
nand U24697 (N_24697,N_18448,N_16802);
xor U24698 (N_24698,N_13288,N_17684);
nand U24699 (N_24699,N_16273,N_12629);
nand U24700 (N_24700,N_13269,N_15447);
or U24701 (N_24701,N_15250,N_18716);
nand U24702 (N_24702,N_17848,N_13242);
and U24703 (N_24703,N_17681,N_17867);
and U24704 (N_24704,N_17963,N_12509);
or U24705 (N_24705,N_13000,N_13053);
nand U24706 (N_24706,N_17756,N_16485);
xor U24707 (N_24707,N_13383,N_17364);
and U24708 (N_24708,N_17810,N_15589);
xnor U24709 (N_24709,N_13554,N_14223);
xor U24710 (N_24710,N_16046,N_16407);
nor U24711 (N_24711,N_18170,N_12669);
xor U24712 (N_24712,N_17703,N_13430);
nand U24713 (N_24713,N_18186,N_12517);
nand U24714 (N_24714,N_14656,N_14669);
or U24715 (N_24715,N_14773,N_18466);
nand U24716 (N_24716,N_18100,N_17752);
xnor U24717 (N_24717,N_13426,N_12665);
nand U24718 (N_24718,N_16633,N_16535);
xnor U24719 (N_24719,N_14526,N_12771);
xor U24720 (N_24720,N_16292,N_14880);
nand U24721 (N_24721,N_17734,N_13982);
xnor U24722 (N_24722,N_14528,N_12881);
nor U24723 (N_24723,N_16590,N_13537);
and U24724 (N_24724,N_17340,N_12943);
nor U24725 (N_24725,N_15034,N_17256);
or U24726 (N_24726,N_14472,N_17183);
xor U24727 (N_24727,N_17053,N_15572);
and U24728 (N_24728,N_14434,N_17037);
xor U24729 (N_24729,N_13209,N_17720);
or U24730 (N_24730,N_12966,N_14586);
and U24731 (N_24731,N_18095,N_18487);
or U24732 (N_24732,N_16838,N_17514);
or U24733 (N_24733,N_16083,N_12765);
nand U24734 (N_24734,N_13525,N_16934);
nor U24735 (N_24735,N_17045,N_14128);
nor U24736 (N_24736,N_15678,N_15686);
and U24737 (N_24737,N_15319,N_15092);
and U24738 (N_24738,N_15870,N_16846);
nand U24739 (N_24739,N_15601,N_18046);
xor U24740 (N_24740,N_15442,N_18577);
xnor U24741 (N_24741,N_18353,N_15100);
nand U24742 (N_24742,N_13025,N_16000);
and U24743 (N_24743,N_15211,N_16422);
nor U24744 (N_24744,N_18567,N_17570);
xor U24745 (N_24745,N_17482,N_16392);
nand U24746 (N_24746,N_15393,N_17586);
and U24747 (N_24747,N_13476,N_13581);
or U24748 (N_24748,N_14744,N_17601);
xor U24749 (N_24749,N_12740,N_16194);
and U24750 (N_24750,N_17558,N_13176);
and U24751 (N_24751,N_14384,N_13536);
or U24752 (N_24752,N_13666,N_17550);
xor U24753 (N_24753,N_12575,N_15586);
nor U24754 (N_24754,N_15848,N_15172);
nor U24755 (N_24755,N_14312,N_16656);
or U24756 (N_24756,N_17412,N_17085);
xnor U24757 (N_24757,N_16529,N_13433);
or U24758 (N_24758,N_14733,N_13044);
or U24759 (N_24759,N_12687,N_17704);
or U24760 (N_24760,N_14275,N_17878);
xor U24761 (N_24761,N_15556,N_17492);
xor U24762 (N_24762,N_13468,N_14509);
and U24763 (N_24763,N_17777,N_13919);
and U24764 (N_24764,N_13528,N_16228);
nor U24765 (N_24765,N_18433,N_16119);
or U24766 (N_24766,N_18423,N_14160);
nand U24767 (N_24767,N_12757,N_12591);
nand U24768 (N_24768,N_15427,N_16527);
xor U24769 (N_24769,N_17220,N_17275);
or U24770 (N_24770,N_17036,N_13114);
or U24771 (N_24771,N_18597,N_13971);
and U24772 (N_24772,N_16823,N_13058);
nand U24773 (N_24773,N_12844,N_15879);
nor U24774 (N_24774,N_15935,N_16354);
xor U24775 (N_24775,N_15450,N_15804);
nand U24776 (N_24776,N_14019,N_17659);
nand U24777 (N_24777,N_17590,N_14523);
xnor U24778 (N_24778,N_14370,N_15710);
or U24779 (N_24779,N_14800,N_14500);
nand U24780 (N_24780,N_15681,N_17419);
nand U24781 (N_24781,N_16869,N_18706);
nor U24782 (N_24782,N_14471,N_17741);
nand U24783 (N_24783,N_17109,N_12555);
nor U24784 (N_24784,N_15627,N_16442);
or U24785 (N_24785,N_17960,N_14473);
nand U24786 (N_24786,N_14734,N_15555);
and U24787 (N_24787,N_18674,N_12538);
xnor U24788 (N_24788,N_12841,N_14290);
xnor U24789 (N_24789,N_14307,N_12694);
or U24790 (N_24790,N_13076,N_13928);
xnor U24791 (N_24791,N_17896,N_15253);
nand U24792 (N_24792,N_14317,N_12995);
and U24793 (N_24793,N_16313,N_12929);
xor U24794 (N_24794,N_15890,N_16924);
nor U24795 (N_24795,N_13058,N_15411);
xor U24796 (N_24796,N_16544,N_17764);
xnor U24797 (N_24797,N_17985,N_17683);
nor U24798 (N_24798,N_14009,N_13747);
xor U24799 (N_24799,N_18118,N_14624);
and U24800 (N_24800,N_17164,N_17128);
nor U24801 (N_24801,N_14211,N_18693);
nor U24802 (N_24802,N_13206,N_15829);
nor U24803 (N_24803,N_17749,N_18508);
or U24804 (N_24804,N_16624,N_18506);
or U24805 (N_24805,N_14879,N_17499);
xor U24806 (N_24806,N_13730,N_15145);
nor U24807 (N_24807,N_16522,N_16362);
nand U24808 (N_24808,N_15274,N_18382);
xor U24809 (N_24809,N_14879,N_12822);
and U24810 (N_24810,N_18387,N_18465);
xnor U24811 (N_24811,N_17658,N_17578);
nor U24812 (N_24812,N_12632,N_14334);
xnor U24813 (N_24813,N_17752,N_18568);
xor U24814 (N_24814,N_17864,N_14916);
xor U24815 (N_24815,N_16667,N_15461);
xnor U24816 (N_24816,N_18635,N_13661);
and U24817 (N_24817,N_15225,N_17476);
nand U24818 (N_24818,N_18468,N_17993);
xor U24819 (N_24819,N_16642,N_17213);
or U24820 (N_24820,N_14837,N_15337);
nand U24821 (N_24821,N_13683,N_13477);
xor U24822 (N_24822,N_18008,N_15125);
and U24823 (N_24823,N_17867,N_14186);
xor U24824 (N_24824,N_14592,N_13076);
xor U24825 (N_24825,N_13668,N_18117);
nor U24826 (N_24826,N_14402,N_17407);
xnor U24827 (N_24827,N_14616,N_14697);
xor U24828 (N_24828,N_15609,N_14114);
nor U24829 (N_24829,N_17905,N_17267);
or U24830 (N_24830,N_13694,N_17119);
and U24831 (N_24831,N_17096,N_13732);
or U24832 (N_24832,N_17736,N_15801);
nand U24833 (N_24833,N_16342,N_13656);
nand U24834 (N_24834,N_16852,N_14186);
nor U24835 (N_24835,N_16920,N_14894);
nor U24836 (N_24836,N_13682,N_17934);
nand U24837 (N_24837,N_15145,N_18747);
or U24838 (N_24838,N_12861,N_13969);
and U24839 (N_24839,N_16428,N_18147);
nor U24840 (N_24840,N_18622,N_16758);
and U24841 (N_24841,N_12778,N_13497);
nor U24842 (N_24842,N_18582,N_16097);
or U24843 (N_24843,N_17501,N_12821);
xnor U24844 (N_24844,N_15432,N_18294);
and U24845 (N_24845,N_15192,N_18057);
xor U24846 (N_24846,N_18484,N_17559);
xor U24847 (N_24847,N_14123,N_15894);
and U24848 (N_24848,N_14705,N_16285);
nor U24849 (N_24849,N_16206,N_14955);
nor U24850 (N_24850,N_17156,N_18153);
and U24851 (N_24851,N_18732,N_13763);
nor U24852 (N_24852,N_17293,N_15654);
xnor U24853 (N_24853,N_13629,N_17445);
nor U24854 (N_24854,N_13044,N_18128);
xor U24855 (N_24855,N_15675,N_13138);
or U24856 (N_24856,N_12947,N_16944);
xnor U24857 (N_24857,N_18728,N_15115);
and U24858 (N_24858,N_14003,N_16270);
nor U24859 (N_24859,N_17701,N_13931);
nor U24860 (N_24860,N_18043,N_15074);
and U24861 (N_24861,N_15486,N_18608);
nand U24862 (N_24862,N_13789,N_16268);
and U24863 (N_24863,N_13326,N_13200);
and U24864 (N_24864,N_16651,N_16009);
nand U24865 (N_24865,N_14040,N_17582);
nor U24866 (N_24866,N_18519,N_16736);
nor U24867 (N_24867,N_17210,N_17291);
xnor U24868 (N_24868,N_12954,N_18134);
nor U24869 (N_24869,N_12745,N_13688);
nor U24870 (N_24870,N_18405,N_14213);
nand U24871 (N_24871,N_18193,N_14271);
nand U24872 (N_24872,N_15843,N_14921);
nor U24873 (N_24873,N_17336,N_13886);
nand U24874 (N_24874,N_18099,N_17455);
nor U24875 (N_24875,N_14142,N_16814);
xnor U24876 (N_24876,N_18071,N_14654);
or U24877 (N_24877,N_14846,N_16910);
or U24878 (N_24878,N_16987,N_18519);
nand U24879 (N_24879,N_13211,N_12833);
and U24880 (N_24880,N_18158,N_13781);
or U24881 (N_24881,N_18250,N_18538);
and U24882 (N_24882,N_15372,N_13200);
nor U24883 (N_24883,N_12553,N_15983);
or U24884 (N_24884,N_15287,N_16322);
or U24885 (N_24885,N_17388,N_18536);
nor U24886 (N_24886,N_14354,N_16715);
or U24887 (N_24887,N_16995,N_18478);
nor U24888 (N_24888,N_15073,N_13097);
xnor U24889 (N_24889,N_18545,N_17997);
or U24890 (N_24890,N_16083,N_17141);
and U24891 (N_24891,N_14832,N_17300);
and U24892 (N_24892,N_16000,N_16570);
nor U24893 (N_24893,N_18007,N_12628);
nor U24894 (N_24894,N_15967,N_17133);
nand U24895 (N_24895,N_14640,N_14713);
or U24896 (N_24896,N_15299,N_16531);
and U24897 (N_24897,N_17396,N_18420);
or U24898 (N_24898,N_15935,N_15473);
nand U24899 (N_24899,N_14318,N_14558);
nand U24900 (N_24900,N_15243,N_18083);
xnor U24901 (N_24901,N_14634,N_14123);
and U24902 (N_24902,N_18706,N_13845);
nand U24903 (N_24903,N_18056,N_12523);
and U24904 (N_24904,N_15658,N_15890);
xor U24905 (N_24905,N_14312,N_13077);
xor U24906 (N_24906,N_14635,N_15665);
and U24907 (N_24907,N_12806,N_14848);
nor U24908 (N_24908,N_17257,N_15529);
nor U24909 (N_24909,N_15087,N_14569);
and U24910 (N_24910,N_13203,N_13752);
nand U24911 (N_24911,N_16030,N_16417);
nor U24912 (N_24912,N_14682,N_16485);
and U24913 (N_24913,N_17081,N_14284);
or U24914 (N_24914,N_18234,N_16196);
nand U24915 (N_24915,N_17146,N_12994);
or U24916 (N_24916,N_15943,N_17794);
nand U24917 (N_24917,N_12931,N_16217);
nor U24918 (N_24918,N_16467,N_17416);
xnor U24919 (N_24919,N_13438,N_15480);
xnor U24920 (N_24920,N_13625,N_15172);
nor U24921 (N_24921,N_14674,N_12855);
xnor U24922 (N_24922,N_16758,N_18397);
or U24923 (N_24923,N_18529,N_15209);
or U24924 (N_24924,N_13562,N_13650);
nand U24925 (N_24925,N_13901,N_15726);
nand U24926 (N_24926,N_15511,N_12672);
and U24927 (N_24927,N_13467,N_15931);
or U24928 (N_24928,N_17286,N_15835);
nand U24929 (N_24929,N_14856,N_15093);
nor U24930 (N_24930,N_18524,N_16527);
nor U24931 (N_24931,N_14195,N_18439);
nand U24932 (N_24932,N_17258,N_12934);
nand U24933 (N_24933,N_18579,N_14432);
xnor U24934 (N_24934,N_15360,N_18429);
nand U24935 (N_24935,N_13001,N_15194);
and U24936 (N_24936,N_15341,N_12618);
nand U24937 (N_24937,N_15897,N_14061);
nor U24938 (N_24938,N_16627,N_16637);
nor U24939 (N_24939,N_14642,N_14747);
or U24940 (N_24940,N_17994,N_13350);
nor U24941 (N_24941,N_17566,N_15110);
and U24942 (N_24942,N_12794,N_16586);
and U24943 (N_24943,N_12677,N_18446);
nand U24944 (N_24944,N_13414,N_16378);
nor U24945 (N_24945,N_16709,N_17085);
or U24946 (N_24946,N_16656,N_16848);
nand U24947 (N_24947,N_15475,N_16592);
or U24948 (N_24948,N_14442,N_13947);
nand U24949 (N_24949,N_18083,N_15455);
nand U24950 (N_24950,N_13353,N_14424);
xnor U24951 (N_24951,N_16806,N_17722);
and U24952 (N_24952,N_18607,N_16084);
nor U24953 (N_24953,N_14887,N_17177);
nand U24954 (N_24954,N_13284,N_17856);
nor U24955 (N_24955,N_15990,N_15540);
or U24956 (N_24956,N_13022,N_13772);
nand U24957 (N_24957,N_12682,N_12898);
or U24958 (N_24958,N_13585,N_16388);
and U24959 (N_24959,N_18378,N_13341);
nor U24960 (N_24960,N_14125,N_14409);
nand U24961 (N_24961,N_14008,N_17624);
or U24962 (N_24962,N_14454,N_14404);
nand U24963 (N_24963,N_18500,N_18661);
or U24964 (N_24964,N_16031,N_16619);
or U24965 (N_24965,N_15930,N_13257);
or U24966 (N_24966,N_17128,N_18349);
or U24967 (N_24967,N_15615,N_16519);
nand U24968 (N_24968,N_15721,N_12809);
and U24969 (N_24969,N_17555,N_17377);
or U24970 (N_24970,N_18620,N_18626);
nor U24971 (N_24971,N_16822,N_14451);
nand U24972 (N_24972,N_17871,N_13984);
xor U24973 (N_24973,N_13550,N_17087);
xor U24974 (N_24974,N_12907,N_15011);
and U24975 (N_24975,N_15512,N_17657);
nand U24976 (N_24976,N_17050,N_13976);
nor U24977 (N_24977,N_18038,N_13976);
nand U24978 (N_24978,N_13064,N_14509);
xor U24979 (N_24979,N_14291,N_17007);
xnor U24980 (N_24980,N_14880,N_13774);
nor U24981 (N_24981,N_13134,N_13808);
xor U24982 (N_24982,N_18439,N_13880);
and U24983 (N_24983,N_12691,N_13036);
nor U24984 (N_24984,N_17153,N_13958);
or U24985 (N_24985,N_15140,N_15866);
and U24986 (N_24986,N_17067,N_13121);
nor U24987 (N_24987,N_13404,N_12690);
xnor U24988 (N_24988,N_18403,N_18619);
xor U24989 (N_24989,N_16946,N_17793);
and U24990 (N_24990,N_18368,N_17097);
nor U24991 (N_24991,N_13204,N_15079);
nand U24992 (N_24992,N_14430,N_13311);
or U24993 (N_24993,N_16924,N_18425);
and U24994 (N_24994,N_16011,N_18050);
nor U24995 (N_24995,N_13835,N_13004);
nor U24996 (N_24996,N_16659,N_17926);
xnor U24997 (N_24997,N_17371,N_13227);
and U24998 (N_24998,N_18623,N_16859);
nor U24999 (N_24999,N_14394,N_18427);
nor UO_0 (O_0,N_21074,N_21656);
or UO_1 (O_1,N_19134,N_22901);
nor UO_2 (O_2,N_22259,N_24801);
nor UO_3 (O_3,N_23387,N_20344);
nor UO_4 (O_4,N_23444,N_19995);
xnor UO_5 (O_5,N_19268,N_23980);
nor UO_6 (O_6,N_22119,N_23479);
xor UO_7 (O_7,N_23393,N_21321);
nand UO_8 (O_8,N_19262,N_24146);
nor UO_9 (O_9,N_19867,N_20969);
xnor UO_10 (O_10,N_22862,N_21243);
nor UO_11 (O_11,N_22617,N_19812);
or UO_12 (O_12,N_20657,N_24860);
xor UO_13 (O_13,N_21118,N_22662);
xnor UO_14 (O_14,N_23965,N_23260);
nor UO_15 (O_15,N_23414,N_21883);
nor UO_16 (O_16,N_24498,N_21290);
nor UO_17 (O_17,N_20175,N_23610);
nand UO_18 (O_18,N_20961,N_20474);
or UO_19 (O_19,N_22017,N_23937);
nand UO_20 (O_20,N_19880,N_23793);
xor UO_21 (O_21,N_23033,N_20566);
and UO_22 (O_22,N_23231,N_22312);
nor UO_23 (O_23,N_21623,N_24506);
or UO_24 (O_24,N_24272,N_19331);
nor UO_25 (O_25,N_19640,N_21050);
nor UO_26 (O_26,N_24776,N_21414);
or UO_27 (O_27,N_23014,N_20311);
xor UO_28 (O_28,N_23295,N_20430);
nand UO_29 (O_29,N_24172,N_23357);
or UO_30 (O_30,N_21943,N_21419);
or UO_31 (O_31,N_21671,N_21087);
nor UO_32 (O_32,N_19754,N_22347);
xnor UO_33 (O_33,N_19090,N_24986);
and UO_34 (O_34,N_19939,N_24923);
nand UO_35 (O_35,N_20431,N_19267);
nand UO_36 (O_36,N_24931,N_23091);
or UO_37 (O_37,N_20504,N_20329);
and UO_38 (O_38,N_24675,N_24846);
nand UO_39 (O_39,N_23591,N_23878);
nor UO_40 (O_40,N_23476,N_23163);
and UO_41 (O_41,N_21319,N_19479);
and UO_42 (O_42,N_19361,N_22613);
nand UO_43 (O_43,N_23145,N_24190);
xor UO_44 (O_44,N_22827,N_18769);
xnor UO_45 (O_45,N_22116,N_22291);
nor UO_46 (O_46,N_21689,N_24067);
nor UO_47 (O_47,N_24589,N_18959);
xor UO_48 (O_48,N_23485,N_21484);
or UO_49 (O_49,N_23528,N_19504);
nand UO_50 (O_50,N_19150,N_23283);
xnor UO_51 (O_51,N_23885,N_20509);
and UO_52 (O_52,N_21665,N_20692);
nor UO_53 (O_53,N_20390,N_24118);
nor UO_54 (O_54,N_24399,N_21455);
and UO_55 (O_55,N_20007,N_24501);
xnor UO_56 (O_56,N_22595,N_23077);
xor UO_57 (O_57,N_21744,N_23988);
nor UO_58 (O_58,N_24549,N_23266);
or UO_59 (O_59,N_21864,N_21352);
nor UO_60 (O_60,N_22389,N_24401);
or UO_61 (O_61,N_20499,N_21724);
nor UO_62 (O_62,N_22885,N_20744);
nor UO_63 (O_63,N_20859,N_19818);
and UO_64 (O_64,N_23820,N_21487);
or UO_65 (O_65,N_19299,N_20507);
or UO_66 (O_66,N_20642,N_20716);
xnor UO_67 (O_67,N_20035,N_23042);
xor UO_68 (O_68,N_22205,N_22311);
nor UO_69 (O_69,N_20876,N_21501);
nor UO_70 (O_70,N_19056,N_19355);
and UO_71 (O_71,N_20972,N_18817);
or UO_72 (O_72,N_21509,N_21267);
or UO_73 (O_73,N_21706,N_23380);
or UO_74 (O_74,N_21497,N_21170);
and UO_75 (O_75,N_24220,N_20325);
nor UO_76 (O_76,N_22697,N_19254);
xnor UO_77 (O_77,N_24640,N_23092);
and UO_78 (O_78,N_22274,N_22674);
or UO_79 (O_79,N_24936,N_23707);
or UO_80 (O_80,N_19264,N_20619);
nand UO_81 (O_81,N_24041,N_20111);
and UO_82 (O_82,N_20239,N_23970);
or UO_83 (O_83,N_19684,N_23105);
xnor UO_84 (O_84,N_21451,N_19656);
nor UO_85 (O_85,N_24376,N_20373);
or UO_86 (O_86,N_20779,N_21088);
nor UO_87 (O_87,N_24817,N_22063);
xnor UO_88 (O_88,N_22546,N_21466);
nor UO_89 (O_89,N_20124,N_22607);
and UO_90 (O_90,N_21098,N_24750);
xnor UO_91 (O_91,N_24449,N_19742);
xor UO_92 (O_92,N_21990,N_20277);
nor UO_93 (O_93,N_19289,N_19310);
and UO_94 (O_94,N_21475,N_21401);
nor UO_95 (O_95,N_22496,N_23178);
xor UO_96 (O_96,N_18983,N_24875);
nor UO_97 (O_97,N_21651,N_20603);
nand UO_98 (O_98,N_23730,N_24641);
or UO_99 (O_99,N_20490,N_24322);
nor UO_100 (O_100,N_18879,N_21531);
or UO_101 (O_101,N_24264,N_22949);
xor UO_102 (O_102,N_22603,N_19883);
or UO_103 (O_103,N_21412,N_19788);
and UO_104 (O_104,N_23358,N_24335);
nand UO_105 (O_105,N_23764,N_24344);
or UO_106 (O_106,N_19165,N_22791);
xnor UO_107 (O_107,N_24767,N_22399);
and UO_108 (O_108,N_20608,N_22764);
xnor UO_109 (O_109,N_23397,N_20655);
and UO_110 (O_110,N_22393,N_20511);
nand UO_111 (O_111,N_24310,N_22130);
xor UO_112 (O_112,N_24325,N_23902);
and UO_113 (O_113,N_23676,N_20717);
or UO_114 (O_114,N_18981,N_21722);
nor UO_115 (O_115,N_23087,N_19723);
xor UO_116 (O_116,N_19367,N_19810);
nor UO_117 (O_117,N_22372,N_20123);
xnor UO_118 (O_118,N_20061,N_24574);
nor UO_119 (O_119,N_19138,N_19458);
or UO_120 (O_120,N_24351,N_18904);
and UO_121 (O_121,N_20117,N_19392);
nand UO_122 (O_122,N_24983,N_19382);
nand UO_123 (O_123,N_24929,N_23931);
xnor UO_124 (O_124,N_20081,N_19647);
nand UO_125 (O_125,N_23149,N_20886);
and UO_126 (O_126,N_23616,N_23951);
or UO_127 (O_127,N_19193,N_22933);
or UO_128 (O_128,N_23119,N_23169);
xor UO_129 (O_129,N_22159,N_23705);
or UO_130 (O_130,N_23983,N_19916);
and UO_131 (O_131,N_23964,N_21546);
or UO_132 (O_132,N_20918,N_24160);
or UO_133 (O_133,N_21700,N_22763);
or UO_134 (O_134,N_20863,N_24063);
nor UO_135 (O_135,N_18913,N_18860);
or UO_136 (O_136,N_21095,N_24511);
or UO_137 (O_137,N_19119,N_21986);
nand UO_138 (O_138,N_24466,N_20354);
nor UO_139 (O_139,N_20898,N_24505);
or UO_140 (O_140,N_18935,N_19046);
and UO_141 (O_141,N_24768,N_21370);
xnor UO_142 (O_142,N_24763,N_22362);
or UO_143 (O_143,N_19806,N_22436);
xnor UO_144 (O_144,N_20467,N_22925);
and UO_145 (O_145,N_22792,N_20633);
nor UO_146 (O_146,N_19461,N_20183);
nor UO_147 (O_147,N_20729,N_24033);
nand UO_148 (O_148,N_23636,N_21933);
nor UO_149 (O_149,N_21849,N_20451);
nor UO_150 (O_150,N_23689,N_24142);
xor UO_151 (O_151,N_22295,N_21355);
or UO_152 (O_152,N_23767,N_24785);
xor UO_153 (O_153,N_21038,N_22958);
and UO_154 (O_154,N_20809,N_23121);
xnor UO_155 (O_155,N_21175,N_22637);
nand UO_156 (O_156,N_23870,N_23760);
or UO_157 (O_157,N_19120,N_24577);
nand UO_158 (O_158,N_19739,N_21131);
nor UO_159 (O_159,N_21174,N_22369);
or UO_160 (O_160,N_23113,N_24550);
or UO_161 (O_161,N_24567,N_19368);
nor UO_162 (O_162,N_20556,N_21931);
nand UO_163 (O_163,N_22175,N_19437);
or UO_164 (O_164,N_24448,N_19650);
nand UO_165 (O_165,N_21900,N_23976);
xnor UO_166 (O_166,N_20500,N_22066);
xor UO_167 (O_167,N_20101,N_20588);
xnor UO_168 (O_168,N_22745,N_20181);
and UO_169 (O_169,N_21379,N_22518);
and UO_170 (O_170,N_20418,N_24321);
or UO_171 (O_171,N_21029,N_19335);
nor UO_172 (O_172,N_18875,N_21291);
xor UO_173 (O_173,N_21720,N_23401);
and UO_174 (O_174,N_24676,N_22582);
or UO_175 (O_175,N_19843,N_21371);
and UO_176 (O_176,N_21664,N_22927);
or UO_177 (O_177,N_20502,N_23913);
or UO_178 (O_178,N_22672,N_21042);
and UO_179 (O_179,N_23316,N_21279);
or UO_180 (O_180,N_23122,N_19982);
nor UO_181 (O_181,N_22472,N_22869);
or UO_182 (O_182,N_22442,N_22330);
nand UO_183 (O_183,N_21333,N_21113);
nand UO_184 (O_184,N_19936,N_24833);
and UO_185 (O_185,N_21498,N_20468);
and UO_186 (O_186,N_24704,N_21168);
or UO_187 (O_187,N_23765,N_20133);
nor UO_188 (O_188,N_19620,N_21912);
xnor UO_189 (O_189,N_18869,N_21181);
nand UO_190 (O_190,N_22645,N_20552);
or UO_191 (O_191,N_23047,N_22848);
and UO_192 (O_192,N_21397,N_23425);
xnor UO_193 (O_193,N_22811,N_20766);
nand UO_194 (O_194,N_24495,N_21879);
nand UO_195 (O_195,N_21364,N_24114);
nor UO_196 (O_196,N_22267,N_23018);
nor UO_197 (O_197,N_24665,N_21732);
nand UO_198 (O_198,N_21630,N_23439);
xor UO_199 (O_199,N_21874,N_22826);
or UO_200 (O_200,N_18826,N_21597);
or UO_201 (O_201,N_20911,N_24420);
nor UO_202 (O_202,N_19817,N_24112);
nor UO_203 (O_203,N_22984,N_21235);
nor UO_204 (O_204,N_24475,N_20414);
or UO_205 (O_205,N_18903,N_21872);
and UO_206 (O_206,N_22386,N_21821);
nor UO_207 (O_207,N_22029,N_22887);
nand UO_208 (O_208,N_21640,N_19468);
nor UO_209 (O_209,N_20360,N_23867);
xnor UO_210 (O_210,N_20108,N_22693);
nand UO_211 (O_211,N_21791,N_20607);
and UO_212 (O_212,N_20539,N_24513);
nand UO_213 (O_213,N_24065,N_24944);
and UO_214 (O_214,N_23146,N_20030);
or UO_215 (O_215,N_19233,N_19763);
and UO_216 (O_216,N_23265,N_23621);
or UO_217 (O_217,N_23207,N_19644);
or UO_218 (O_218,N_18809,N_20764);
xor UO_219 (O_219,N_21491,N_20113);
or UO_220 (O_220,N_22810,N_23673);
xnor UO_221 (O_221,N_22303,N_20463);
or UO_222 (O_222,N_23906,N_24880);
nand UO_223 (O_223,N_19433,N_23667);
and UO_224 (O_224,N_21992,N_19885);
nand UO_225 (O_225,N_19702,N_22584);
nor UO_226 (O_226,N_20562,N_19309);
or UO_227 (O_227,N_20204,N_23461);
xnor UO_228 (O_228,N_21737,N_23829);
and UO_229 (O_229,N_21457,N_24965);
or UO_230 (O_230,N_22707,N_19703);
and UO_231 (O_231,N_19799,N_22247);
or UO_232 (O_232,N_20601,N_22860);
xnor UO_233 (O_233,N_21756,N_23477);
and UO_234 (O_234,N_19607,N_22153);
xnor UO_235 (O_235,N_19615,N_19339);
nor UO_236 (O_236,N_23398,N_21081);
or UO_237 (O_237,N_20096,N_23194);
nand UO_238 (O_238,N_20709,N_23889);
and UO_239 (O_239,N_23935,N_23454);
and UO_240 (O_240,N_24761,N_20217);
nor UO_241 (O_241,N_21406,N_20284);
or UO_242 (O_242,N_19016,N_21767);
xor UO_243 (O_243,N_24618,N_21408);
nand UO_244 (O_244,N_23487,N_24056);
or UO_245 (O_245,N_24298,N_20212);
and UO_246 (O_246,N_21760,N_19213);
nor UO_247 (O_247,N_21729,N_24612);
nand UO_248 (O_248,N_22000,N_24836);
or UO_249 (O_249,N_24997,N_21776);
and UO_250 (O_250,N_19876,N_21749);
nor UO_251 (O_251,N_23865,N_19553);
and UO_252 (O_252,N_22398,N_20921);
xnor UO_253 (O_253,N_20236,N_22755);
nor UO_254 (O_254,N_18772,N_19899);
and UO_255 (O_255,N_20524,N_24650);
nand UO_256 (O_256,N_23108,N_20027);
or UO_257 (O_257,N_23144,N_23921);
nor UO_258 (O_258,N_20651,N_22015);
nor UO_259 (O_259,N_22454,N_20658);
and UO_260 (O_260,N_20094,N_21218);
or UO_261 (O_261,N_24843,N_23589);
and UO_262 (O_262,N_22475,N_22986);
xor UO_263 (O_263,N_20713,N_24708);
or UO_264 (O_264,N_20760,N_24167);
xnor UO_265 (O_265,N_19265,N_21053);
nor UO_266 (O_266,N_24547,N_19466);
or UO_267 (O_267,N_21748,N_19135);
nand UO_268 (O_268,N_21367,N_20997);
nand UO_269 (O_269,N_20924,N_24855);
xnor UO_270 (O_270,N_22052,N_23185);
or UO_271 (O_271,N_22028,N_21194);
xor UO_272 (O_272,N_23566,N_23781);
or UO_273 (O_273,N_20115,N_18885);
and UO_274 (O_274,N_19825,N_19263);
or UO_275 (O_275,N_24425,N_21479);
or UO_276 (O_276,N_23232,N_22642);
nor UO_277 (O_277,N_22985,N_21676);
xnor UO_278 (O_278,N_21153,N_24955);
xor UO_279 (O_279,N_21985,N_22906);
nor UO_280 (O_280,N_24392,N_24598);
nand UO_281 (O_281,N_22676,N_19243);
or UO_282 (O_282,N_22950,N_20333);
and UO_283 (O_283,N_24862,N_20148);
nor UO_284 (O_284,N_20477,N_19049);
nand UO_285 (O_285,N_23432,N_23275);
nor UO_286 (O_286,N_22675,N_22337);
or UO_287 (O_287,N_23737,N_23949);
nor UO_288 (O_288,N_20410,N_19029);
and UO_289 (O_289,N_22018,N_23235);
and UO_290 (O_290,N_24473,N_20627);
nor UO_291 (O_291,N_21616,N_22344);
nand UO_292 (O_292,N_22233,N_22075);
and UO_293 (O_293,N_24367,N_19646);
nor UO_294 (O_294,N_22979,N_22004);
or UO_295 (O_295,N_18861,N_24897);
xnor UO_296 (O_296,N_21137,N_21921);
nor UO_297 (O_297,N_23056,N_21890);
or UO_298 (O_298,N_18964,N_23143);
and UO_299 (O_299,N_19002,N_19215);
nor UO_300 (O_300,N_22717,N_21505);
and UO_301 (O_301,N_24611,N_21499);
and UO_302 (O_302,N_23173,N_23202);
and UO_303 (O_303,N_20806,N_24820);
xnor UO_304 (O_304,N_20084,N_23218);
or UO_305 (O_305,N_21507,N_19140);
or UO_306 (O_306,N_23972,N_23986);
or UO_307 (O_307,N_22356,N_23456);
nand UO_308 (O_308,N_23597,N_19168);
xor UO_309 (O_309,N_21984,N_22945);
xor UO_310 (O_310,N_19111,N_23312);
and UO_311 (O_311,N_20276,N_20185);
nor UO_312 (O_312,N_24877,N_24510);
xnor UO_313 (O_313,N_22597,N_19945);
nor UO_314 (O_314,N_23830,N_18911);
nor UO_315 (O_315,N_21341,N_19698);
xor UO_316 (O_316,N_23481,N_22877);
xnor UO_317 (O_317,N_22741,N_22983);
or UO_318 (O_318,N_20260,N_21530);
or UO_319 (O_319,N_18758,N_20403);
nor UO_320 (O_320,N_21496,N_18883);
nor UO_321 (O_321,N_21844,N_20644);
xnor UO_322 (O_322,N_19674,N_22196);
or UO_323 (O_323,N_24006,N_22653);
nor UO_324 (O_324,N_24672,N_20940);
nor UO_325 (O_325,N_23258,N_21648);
or UO_326 (O_326,N_20542,N_24740);
nand UO_327 (O_327,N_23584,N_24615);
nand UO_328 (O_328,N_23799,N_23752);
nand UO_329 (O_329,N_22323,N_19951);
or UO_330 (O_330,N_23293,N_22381);
and UO_331 (O_331,N_21545,N_21778);
nand UO_332 (O_332,N_19796,N_22659);
and UO_333 (O_333,N_23975,N_19581);
and UO_334 (O_334,N_23125,N_24739);
nand UO_335 (O_335,N_23967,N_19438);
nor UO_336 (O_336,N_21470,N_19209);
xor UO_337 (O_337,N_19218,N_22098);
nand UO_338 (O_338,N_21429,N_22433);
or UO_339 (O_339,N_21641,N_24822);
nand UO_340 (O_340,N_21293,N_23816);
nor UO_341 (O_341,N_24688,N_22186);
or UO_342 (O_342,N_24780,N_24089);
nand UO_343 (O_343,N_23035,N_23706);
or UO_344 (O_344,N_22955,N_23239);
nand UO_345 (O_345,N_20290,N_21123);
and UO_346 (O_346,N_22225,N_22612);
nor UO_347 (O_347,N_22825,N_23857);
and UO_348 (O_348,N_19475,N_23715);
xnor UO_349 (O_349,N_23971,N_21682);
and UO_350 (O_350,N_22744,N_23209);
or UO_351 (O_351,N_21918,N_19700);
nand UO_352 (O_352,N_22260,N_20763);
and UO_353 (O_353,N_23004,N_23190);
and UO_354 (O_354,N_20450,N_20054);
and UO_355 (O_355,N_22999,N_24130);
nor UO_356 (O_356,N_20643,N_19819);
nor UO_357 (O_357,N_21206,N_21610);
xnor UO_358 (O_358,N_24829,N_20928);
and UO_359 (O_359,N_24668,N_21435);
nor UO_360 (O_360,N_24571,N_21044);
nor UO_361 (O_361,N_21232,N_24805);
nor UO_362 (O_362,N_23412,N_22298);
or UO_363 (O_363,N_24288,N_21220);
xnor UO_364 (O_364,N_24357,N_24137);
xor UO_365 (O_365,N_21997,N_21780);
and UO_366 (O_366,N_20688,N_22509);
or UO_367 (O_367,N_20963,N_22317);
nand UO_368 (O_368,N_20480,N_21846);
and UO_369 (O_369,N_20492,N_18909);
or UO_370 (O_370,N_24174,N_23264);
xor UO_371 (O_371,N_22554,N_20031);
or UO_372 (O_372,N_19760,N_19069);
or UO_373 (O_373,N_22971,N_24770);
nor UO_374 (O_374,N_19801,N_20055);
xor UO_375 (O_375,N_24960,N_24738);
and UO_376 (O_376,N_20993,N_19381);
and UO_377 (O_377,N_23592,N_23052);
and UO_378 (O_378,N_22593,N_20647);
and UO_379 (O_379,N_21387,N_22085);
nor UO_380 (O_380,N_18871,N_23392);
xor UO_381 (O_381,N_22458,N_19068);
nand UO_382 (O_382,N_18991,N_21415);
or UO_383 (O_383,N_23375,N_20540);
nor UO_384 (O_384,N_18868,N_20543);
and UO_385 (O_385,N_23997,N_23489);
and UO_386 (O_386,N_20151,N_19765);
nor UO_387 (O_387,N_19203,N_23718);
xor UO_388 (O_388,N_22532,N_19467);
and UO_389 (O_389,N_22778,N_22375);
or UO_390 (O_390,N_19860,N_20957);
nor UO_391 (O_391,N_22162,N_24514);
nor UO_392 (O_392,N_21977,N_23774);
or UO_393 (O_393,N_19990,N_19343);
xor UO_394 (O_394,N_22682,N_22053);
xnor UO_395 (O_395,N_21799,N_23428);
xnor UO_396 (O_396,N_23679,N_24538);
or UO_397 (O_397,N_24690,N_21427);
nand UO_398 (O_398,N_23623,N_22412);
xnor UO_399 (O_399,N_19547,N_23999);
or UO_400 (O_400,N_21369,N_19348);
nor UO_401 (O_401,N_24745,N_22271);
nand UO_402 (O_402,N_19220,N_21898);
nor UO_403 (O_403,N_19992,N_21214);
or UO_404 (O_404,N_18837,N_24649);
or UO_405 (O_405,N_18881,N_24661);
xor UO_406 (O_406,N_22378,N_24747);
nor UO_407 (O_407,N_22560,N_23001);
xnor UO_408 (O_408,N_19261,N_20383);
nand UO_409 (O_409,N_21830,N_24078);
nor UO_410 (O_410,N_18822,N_20964);
xor UO_411 (O_411,N_22048,N_21061);
nor UO_412 (O_412,N_19202,N_24129);
and UO_413 (O_413,N_24529,N_20057);
and UO_414 (O_414,N_20223,N_18967);
nand UO_415 (O_415,N_22719,N_22428);
nand UO_416 (O_416,N_19827,N_18957);
nand UO_417 (O_417,N_20224,N_20726);
xnor UO_418 (O_418,N_22350,N_24417);
or UO_419 (O_419,N_24683,N_21309);
or UO_420 (O_420,N_24684,N_21731);
xnor UO_421 (O_421,N_22689,N_18974);
xor UO_422 (O_422,N_20715,N_21109);
xor UO_423 (O_423,N_19952,N_22197);
xor UO_424 (O_424,N_23502,N_19707);
or UO_425 (O_425,N_22524,N_21948);
nand UO_426 (O_426,N_24127,N_20070);
or UO_427 (O_427,N_24657,N_21086);
nand UO_428 (O_428,N_23123,N_19247);
nor UO_429 (O_429,N_24754,N_24970);
nand UO_430 (O_430,N_19717,N_24472);
xor UO_431 (O_431,N_23579,N_24343);
and UO_432 (O_432,N_22725,N_18770);
nor UO_433 (O_433,N_19925,N_21351);
nor UO_434 (O_434,N_22872,N_22034);
xnor UO_435 (O_435,N_21636,N_18947);
nor UO_436 (O_436,N_20409,N_20100);
or UO_437 (O_437,N_21485,N_20736);
xnor UO_438 (O_438,N_19942,N_24001);
or UO_439 (O_439,N_19073,N_23569);
nand UO_440 (O_440,N_19917,N_22734);
or UO_441 (O_441,N_22103,N_21069);
nand UO_442 (O_442,N_20317,N_21916);
xor UO_443 (O_443,N_20517,N_20210);
xnor UO_444 (O_444,N_24125,N_24534);
nand UO_445 (O_445,N_22864,N_23030);
or UO_446 (O_446,N_22054,N_20278);
xnor UO_447 (O_447,N_23089,N_19693);
xor UO_448 (O_448,N_24769,N_23536);
nor UO_449 (O_449,N_19848,N_19034);
nand UO_450 (O_450,N_23363,N_21983);
nand UO_451 (O_451,N_21654,N_20011);
xor UO_452 (O_452,N_23839,N_19533);
and UO_453 (O_453,N_22576,N_19464);
and UO_454 (O_454,N_22747,N_23912);
and UO_455 (O_455,N_23572,N_22483);
nand UO_456 (O_456,N_24517,N_20404);
nor UO_457 (O_457,N_20323,N_18783);
nor UO_458 (O_458,N_19048,N_19732);
xor UO_459 (O_459,N_19177,N_20227);
or UO_460 (O_460,N_24415,N_24911);
nor UO_461 (O_461,N_21030,N_20738);
or UO_462 (O_462,N_20427,N_24445);
and UO_463 (O_463,N_20949,N_22070);
and UO_464 (O_464,N_21152,N_23259);
or UO_465 (O_465,N_21114,N_19451);
nand UO_466 (O_466,N_19514,N_23959);
and UO_467 (O_467,N_24626,N_19971);
nor UO_468 (O_468,N_22564,N_20789);
and UO_469 (O_469,N_20881,N_23506);
or UO_470 (O_470,N_24782,N_21149);
xnor UO_471 (O_471,N_20922,N_24126);
xnor UO_472 (O_472,N_20371,N_21907);
or UO_473 (O_473,N_22807,N_23464);
xnor UO_474 (O_474,N_22168,N_24477);
nand UO_475 (O_475,N_23908,N_24968);
xor UO_476 (O_476,N_21273,N_20334);
nand UO_477 (O_477,N_24181,N_20889);
nand UO_478 (O_478,N_20080,N_22123);
and UO_479 (O_479,N_20640,N_21839);
or UO_480 (O_480,N_21856,N_24723);
xor UO_481 (O_481,N_22464,N_20439);
and UO_482 (O_482,N_19854,N_20233);
nand UO_483 (O_483,N_24864,N_19767);
nand UO_484 (O_484,N_23457,N_20663);
nor UO_485 (O_485,N_19067,N_19121);
and UO_486 (O_486,N_22880,N_23953);
or UO_487 (O_487,N_23302,N_20823);
nand UO_488 (O_488,N_19211,N_22132);
xor UO_489 (O_489,N_21606,N_22209);
or UO_490 (O_490,N_19712,N_21444);
and UO_491 (O_491,N_22528,N_21468);
or UO_492 (O_492,N_21200,N_20402);
nand UO_493 (O_493,N_24178,N_20350);
and UO_494 (O_494,N_19652,N_20422);
xnor UO_495 (O_495,N_24643,N_18841);
nand UO_496 (O_496,N_24362,N_20564);
or UO_497 (O_497,N_21411,N_19655);
or UO_498 (O_498,N_23073,N_24188);
xor UO_499 (O_499,N_24474,N_19637);
or UO_500 (O_500,N_19544,N_22023);
nor UO_501 (O_501,N_22875,N_21593);
nor UO_502 (O_502,N_19377,N_23172);
and UO_503 (O_503,N_24180,N_23000);
nand UO_504 (O_504,N_24906,N_21405);
or UO_505 (O_505,N_18971,N_22926);
and UO_506 (O_506,N_20857,N_23458);
or UO_507 (O_507,N_21313,N_20206);
xnor UO_508 (O_508,N_20984,N_24214);
nor UO_509 (O_509,N_20134,N_19216);
xnor UO_510 (O_510,N_18862,N_24594);
nor UO_511 (O_511,N_24090,N_24601);
or UO_512 (O_512,N_22865,N_23148);
nand UO_513 (O_513,N_22881,N_21226);
nor UO_514 (O_514,N_18919,N_19826);
or UO_515 (O_515,N_19295,N_23545);
xnor UO_516 (O_516,N_24256,N_22961);
or UO_517 (O_517,N_24329,N_20589);
xor UO_518 (O_518,N_23903,N_21937);
xnor UO_519 (O_519,N_23532,N_23982);
xnor UO_520 (O_520,N_19422,N_21513);
and UO_521 (O_521,N_20629,N_23698);
nand UO_522 (O_522,N_19131,N_21517);
or UO_523 (O_523,N_19791,N_23225);
and UO_524 (O_524,N_21522,N_24201);
and UO_525 (O_525,N_24818,N_23187);
or UO_526 (O_526,N_20706,N_21205);
nand UO_527 (O_527,N_24358,N_21346);
or UO_528 (O_528,N_22771,N_20132);
and UO_529 (O_529,N_24900,N_23809);
nand UO_530 (O_530,N_19256,N_24369);
xnor UO_531 (O_531,N_19191,N_19568);
nand UO_532 (O_532,N_20622,N_19424);
nand UO_533 (O_533,N_18951,N_22649);
nand UO_534 (O_534,N_22752,N_23909);
nor UO_535 (O_535,N_19850,N_23968);
nor UO_536 (O_536,N_18779,N_21979);
xnor UO_537 (O_537,N_24625,N_22500);
nand UO_538 (O_538,N_21960,N_22710);
nand UO_539 (O_539,N_24192,N_23132);
and UO_540 (O_540,N_20796,N_22257);
and UO_541 (O_541,N_19682,N_24106);
nor UO_542 (O_542,N_23845,N_21027);
and UO_543 (O_543,N_19148,N_21422);
xnor UO_544 (O_544,N_22787,N_23749);
xnor UO_545 (O_545,N_23241,N_19164);
xnor UO_546 (O_546,N_19174,N_23992);
nor UO_547 (O_547,N_20938,N_22730);
and UO_548 (O_548,N_20546,N_24166);
and UO_549 (O_549,N_21473,N_24637);
nand UO_550 (O_550,N_21573,N_24212);
nand UO_551 (O_551,N_20397,N_21139);
and UO_552 (O_552,N_21873,N_20844);
and UO_553 (O_553,N_20781,N_23196);
nor UO_554 (O_554,N_22346,N_19649);
nor UO_555 (O_555,N_19878,N_24393);
and UO_556 (O_556,N_21418,N_22480);
xnor UO_557 (O_557,N_21569,N_21614);
xor UO_558 (O_558,N_23948,N_23775);
nor UO_559 (O_559,N_22749,N_24604);
nor UO_560 (O_560,N_21456,N_23639);
nand UO_561 (O_561,N_23208,N_24627);
or UO_562 (O_562,N_22282,N_22127);
nor UO_563 (O_563,N_19718,N_20202);
or UO_564 (O_564,N_24297,N_24086);
nor UO_565 (O_565,N_19623,N_19858);
and UO_566 (O_566,N_23580,N_21741);
or UO_567 (O_567,N_24294,N_19207);
nand UO_568 (O_568,N_22842,N_24899);
or UO_569 (O_569,N_24271,N_19095);
and UO_570 (O_570,N_23410,N_20155);
and UO_571 (O_571,N_21835,N_23888);
nand UO_572 (O_572,N_24389,N_24691);
xor UO_573 (O_573,N_23273,N_21721);
or UO_574 (O_574,N_22046,N_18843);
nor UO_575 (O_575,N_24453,N_19772);
nand UO_576 (O_576,N_20926,N_23918);
nor UO_577 (O_577,N_22051,N_22658);
nor UO_578 (O_578,N_24564,N_20318);
or UO_579 (O_579,N_18952,N_21328);
and UO_580 (O_580,N_24645,N_19890);
and UO_581 (O_581,N_19645,N_19189);
nor UO_582 (O_582,N_20526,N_23694);
and UO_583 (O_583,N_21426,N_22767);
and UO_584 (O_584,N_18993,N_20391);
nor UO_585 (O_585,N_24113,N_22818);
or UO_586 (O_586,N_19124,N_21239);
or UO_587 (O_587,N_22477,N_18961);
nand UO_588 (O_588,N_20078,N_21911);
and UO_589 (O_589,N_24976,N_24863);
or UO_590 (O_590,N_23759,N_19534);
nand UO_591 (O_591,N_20216,N_19226);
nor UO_592 (O_592,N_24183,N_21345);
or UO_593 (O_593,N_22363,N_24431);
nand UO_594 (O_594,N_22972,N_21253);
or UO_595 (O_595,N_22967,N_20873);
nand UO_596 (O_596,N_21638,N_23029);
xor UO_597 (O_597,N_20454,N_24055);
nand UO_598 (O_598,N_20800,N_22430);
or UO_599 (O_599,N_21199,N_23068);
nand UO_600 (O_600,N_20660,N_24315);
or UO_601 (O_601,N_23709,N_20005);
nor UO_602 (O_602,N_20558,N_23608);
nor UO_603 (O_603,N_21793,N_24375);
nor UO_604 (O_604,N_24576,N_24017);
nor UO_605 (O_605,N_23868,N_24384);
nor UO_606 (O_606,N_20032,N_20535);
or UO_607 (O_607,N_24365,N_21259);
and UO_608 (O_608,N_23082,N_21978);
xor UO_609 (O_609,N_21582,N_24326);
nand UO_610 (O_610,N_19240,N_22634);
nand UO_611 (O_611,N_24794,N_23553);
nor UO_612 (O_612,N_22213,N_21157);
nor UO_613 (O_613,N_21382,N_22269);
nand UO_614 (O_614,N_18755,N_18937);
and UO_615 (O_615,N_21715,N_22648);
xnor UO_616 (O_616,N_22377,N_24617);
or UO_617 (O_617,N_20508,N_19151);
nor UO_618 (O_618,N_24374,N_22773);
xor UO_619 (O_619,N_23452,N_19483);
and UO_620 (O_620,N_21951,N_19839);
nor UO_621 (O_621,N_21129,N_24088);
and UO_622 (O_622,N_23825,N_18753);
xnor UO_623 (O_623,N_20297,N_23065);
nor UO_624 (O_624,N_22287,N_24687);
and UO_625 (O_625,N_20567,N_19004);
xnor UO_626 (O_626,N_20244,N_22846);
or UO_627 (O_627,N_20639,N_24224);
nand UO_628 (O_628,N_24603,N_20955);
and UO_629 (O_629,N_20161,N_22929);
nand UO_630 (O_630,N_19662,N_23115);
nand UO_631 (O_631,N_18977,N_18966);
and UO_632 (O_632,N_19969,N_24578);
xor UO_633 (O_633,N_19455,N_23031);
nand UO_634 (O_634,N_22329,N_19813);
and UO_635 (O_635,N_23386,N_18789);
nand UO_636 (O_636,N_22095,N_22608);
nand UO_637 (O_637,N_20041,N_24784);
and UO_638 (O_638,N_20826,N_22463);
nor UO_639 (O_639,N_24994,N_22692);
nor UO_640 (O_640,N_21811,N_20425);
and UO_641 (O_641,N_19330,N_20326);
nor UO_642 (O_642,N_19653,N_18893);
nor UO_643 (O_643,N_20252,N_19239);
nand UO_644 (O_644,N_19874,N_22146);
or UO_645 (O_645,N_24029,N_19539);
or UO_646 (O_646,N_21359,N_24807);
xor UO_647 (O_647,N_19374,N_23858);
xor UO_648 (O_648,N_23915,N_21605);
and UO_649 (O_649,N_23886,N_22998);
xor UO_650 (O_650,N_20693,N_23595);
nor UO_651 (O_651,N_19953,N_20264);
and UO_652 (O_652,N_23782,N_22988);
nor UO_653 (O_653,N_23519,N_24437);
xnor UO_654 (O_654,N_23263,N_18912);
nand UO_655 (O_655,N_21450,N_23813);
nor UO_656 (O_656,N_24023,N_22166);
or UO_657 (O_657,N_24925,N_20846);
nor UO_658 (O_658,N_20787,N_18917);
nand UO_659 (O_659,N_21102,N_21002);
nor UO_660 (O_660,N_19577,N_22928);
and UO_661 (O_661,N_22187,N_21807);
nor UO_662 (O_662,N_21763,N_23603);
and UO_663 (O_663,N_20109,N_19643);
xnor UO_664 (O_664,N_21305,N_20962);
xor UO_665 (O_665,N_21843,N_21525);
and UO_666 (O_666,N_21765,N_21008);
or UO_667 (O_667,N_21613,N_21448);
and UO_668 (O_668,N_24609,N_19336);
and UO_669 (O_669,N_23795,N_19979);
xor UO_670 (O_670,N_23057,N_22379);
xor UO_671 (O_671,N_22756,N_21402);
xor UO_672 (O_672,N_20678,N_23070);
nand UO_673 (O_673,N_22656,N_18776);
nor UO_674 (O_674,N_21975,N_22102);
nand UO_675 (O_675,N_21698,N_22713);
xnor UO_676 (O_676,N_23966,N_21540);
or UO_677 (O_677,N_23855,N_22026);
and UO_678 (O_678,N_18925,N_20628);
nor UO_679 (O_679,N_20583,N_23510);
nor UO_680 (O_680,N_21675,N_19055);
nand UO_681 (O_681,N_21461,N_19127);
nor UO_682 (O_682,N_20462,N_24447);
and UO_683 (O_683,N_21383,N_21662);
or UO_684 (O_684,N_24432,N_21025);
xor UO_685 (O_685,N_22019,N_23854);
xnor UO_686 (O_686,N_23741,N_22913);
nand UO_687 (O_687,N_23655,N_24917);
or UO_688 (O_688,N_20933,N_22450);
and UO_689 (O_689,N_22772,N_23778);
xor UO_690 (O_690,N_20827,N_19708);
or UO_691 (O_691,N_24671,N_23153);
xnor UO_692 (O_692,N_18972,N_18978);
or UO_693 (O_693,N_21609,N_24346);
nand UO_694 (O_694,N_23352,N_19407);
xnor UO_695 (O_695,N_24630,N_20891);
nand UO_696 (O_696,N_23009,N_24573);
nor UO_697 (O_697,N_23880,N_22376);
and UO_698 (O_698,N_20956,N_18985);
and UO_699 (O_699,N_21718,N_20060);
nand UO_700 (O_700,N_22976,N_23379);
xor UO_701 (O_701,N_21127,N_21914);
or UO_702 (O_702,N_23473,N_21816);
xor UO_703 (O_703,N_24080,N_23345);
xor UO_704 (O_704,N_24774,N_20092);
and UO_705 (O_705,N_24002,N_24102);
and UO_706 (O_706,N_24299,N_21228);
xnor UO_707 (O_707,N_23049,N_22037);
or UO_708 (O_708,N_18870,N_21574);
and UO_709 (O_709,N_20851,N_22279);
and UO_710 (O_710,N_21808,N_22720);
and UO_711 (O_711,N_22432,N_24039);
or UO_712 (O_712,N_18852,N_24659);
xnor UO_713 (O_713,N_21625,N_23803);
nor UO_714 (O_714,N_24208,N_24164);
nor UO_715 (O_715,N_20885,N_20098);
and UO_716 (O_716,N_21775,N_19340);
or UO_717 (O_717,N_22650,N_22069);
xnor UO_718 (O_718,N_21692,N_20200);
or UO_719 (O_719,N_24442,N_19820);
xnor UO_720 (O_720,N_23893,N_22444);
xor UO_721 (O_721,N_19861,N_24199);
and UO_722 (O_722,N_20308,N_23744);
and UO_723 (O_723,N_24713,N_20443);
nor UO_724 (O_724,N_21348,N_22614);
xnor UO_725 (O_725,N_21452,N_23383);
xnor UO_726 (O_726,N_19178,N_19477);
nor UO_727 (O_727,N_21179,N_24053);
or UO_728 (O_728,N_21249,N_19001);
xnor UO_729 (O_729,N_23496,N_20447);
nor UO_730 (O_730,N_21037,N_19587);
or UO_731 (O_731,N_18794,N_19186);
nor UO_732 (O_732,N_24111,N_23620);
and UO_733 (O_733,N_22632,N_23708);
or UO_734 (O_734,N_24562,N_18790);
or UO_735 (O_735,N_19527,N_20865);
xnor UO_736 (O_736,N_19926,N_18799);
xnor UO_737 (O_737,N_19353,N_23254);
or UO_738 (O_738,N_24073,N_24232);
nand UO_739 (O_739,N_19571,N_19790);
nand UO_740 (O_740,N_22631,N_19166);
nand UO_741 (O_741,N_23353,N_23929);
or UO_742 (O_742,N_24396,N_21929);
nor UO_743 (O_743,N_21284,N_23409);
or UO_744 (O_744,N_23007,N_19409);
and UO_745 (O_745,N_18774,N_19532);
and UO_746 (O_746,N_22558,N_21178);
or UO_747 (O_747,N_23734,N_23083);
and UO_748 (O_748,N_20421,N_20650);
nand UO_749 (O_749,N_20428,N_21110);
xor UO_750 (O_750,N_24895,N_22488);
nand UO_751 (O_751,N_19162,N_21766);
or UO_752 (O_752,N_23794,N_21868);
xor UO_753 (O_753,N_23523,N_24908);
or UO_754 (O_754,N_21566,N_21925);
xnor UO_755 (O_755,N_23890,N_22735);
nor UO_756 (O_756,N_24595,N_19258);
nor UO_757 (O_757,N_21004,N_19689);
or UO_758 (O_758,N_24508,N_19559);
nor UO_759 (O_759,N_19835,N_22422);
nand UO_760 (O_760,N_19642,N_24340);
or UO_761 (O_761,N_19497,N_20909);
xnor UO_762 (O_762,N_19460,N_23735);
nand UO_763 (O_763,N_22154,N_24743);
and UO_764 (O_764,N_19305,N_19919);
xor UO_765 (O_765,N_22522,N_22190);
and UO_766 (O_766,N_19022,N_19713);
or UO_767 (O_767,N_24715,N_23420);
xor UO_768 (O_768,N_23384,N_22418);
nand UO_769 (O_769,N_22621,N_22997);
or UO_770 (O_770,N_24173,N_21536);
or UO_771 (O_771,N_22003,N_19242);
nand UO_772 (O_772,N_20602,N_19175);
xor UO_773 (O_773,N_22547,N_24610);
nor UO_774 (O_774,N_23726,N_19701);
xor UO_775 (O_775,N_22056,N_24797);
nor UO_776 (O_776,N_20160,N_22615);
xnor UO_777 (O_777,N_24741,N_23441);
xor UO_778 (O_778,N_20665,N_24236);
xnor UO_779 (O_779,N_19397,N_19208);
xor UO_780 (O_780,N_23633,N_22121);
nor UO_781 (O_781,N_20483,N_18905);
and UO_782 (O_782,N_21758,N_20053);
xnor UO_783 (O_783,N_23682,N_19783);
nand UO_784 (O_784,N_24706,N_21436);
xnor UO_785 (O_785,N_22076,N_19506);
or UO_786 (O_786,N_23634,N_23404);
and UO_787 (O_787,N_23662,N_23013);
or UO_788 (O_788,N_22740,N_24655);
nand UO_789 (O_789,N_19695,N_22768);
xnor UO_790 (O_790,N_19968,N_19927);
nand UO_791 (O_791,N_20003,N_20584);
and UO_792 (O_792,N_20561,N_24660);
and UO_793 (O_793,N_22466,N_24099);
nand UO_794 (O_794,N_20052,N_22262);
xor UO_795 (O_795,N_18778,N_18829);
nor UO_796 (O_796,N_22549,N_24128);
or UO_797 (O_797,N_20870,N_19872);
nand UO_798 (O_798,N_22673,N_19074);
nand UO_799 (O_799,N_19098,N_18784);
xnor UO_800 (O_800,N_24874,N_21733);
nor UO_801 (O_801,N_22338,N_21704);
nand UO_802 (O_802,N_23728,N_24451);
xnor UO_803 (O_803,N_20258,N_24244);
and UO_804 (O_804,N_24753,N_21794);
and UO_805 (O_805,N_21552,N_21292);
and UO_806 (O_806,N_22726,N_23071);
and UO_807 (O_807,N_24098,N_24422);
and UO_808 (O_808,N_20380,N_20574);
or UO_809 (O_809,N_22038,N_23842);
and UO_810 (O_810,N_21391,N_21311);
xor UO_811 (O_811,N_23896,N_23116);
nand UO_812 (O_812,N_22072,N_20177);
nor UO_813 (O_813,N_19720,N_22387);
nor UO_814 (O_814,N_22434,N_20791);
and UO_815 (O_815,N_20897,N_22559);
nand UO_816 (O_816,N_19428,N_23466);
and UO_817 (O_817,N_18767,N_23402);
xnor UO_818 (O_818,N_23852,N_24669);
and UO_819 (O_819,N_21020,N_23637);
nor UO_820 (O_820,N_23131,N_21730);
or UO_821 (O_821,N_22133,N_20982);
xnor UO_822 (O_822,N_20248,N_20721);
or UO_823 (O_823,N_20293,N_23137);
nand UO_824 (O_824,N_22936,N_22891);
and UO_825 (O_825,N_21589,N_20338);
nor UO_826 (O_826,N_23859,N_22663);
nor UO_827 (O_827,N_23349,N_22964);
nor UO_828 (O_828,N_22078,N_19507);
or UO_829 (O_829,N_20815,N_20205);
and UO_830 (O_830,N_23670,N_22405);
or UO_831 (O_831,N_21981,N_20525);
nor UO_832 (O_832,N_20804,N_19035);
or UO_833 (O_833,N_21621,N_20710);
nand UO_834 (O_834,N_24479,N_21707);
nor UO_835 (O_835,N_24709,N_23150);
or UO_836 (O_836,N_20550,N_21159);
or UO_837 (O_837,N_19318,N_22370);
and UO_838 (O_838,N_22010,N_22007);
nand UO_839 (O_839,N_24901,N_18754);
nor UO_840 (O_840,N_21409,N_24061);
or UO_841 (O_841,N_22039,N_24842);
xor UO_842 (O_842,N_22061,N_23162);
nor UO_843 (O_843,N_18788,N_22987);
xor UO_844 (O_844,N_20904,N_19445);
or UO_845 (O_845,N_19978,N_22966);
nand UO_846 (O_846,N_24231,N_23361);
nand UO_847 (O_847,N_19276,N_23010);
xnor UO_848 (O_848,N_21045,N_19398);
nand UO_849 (O_849,N_24209,N_22042);
or UO_850 (O_850,N_22530,N_19354);
and UO_851 (O_851,N_19052,N_23962);
nand UO_852 (O_852,N_23804,N_23197);
nor UO_853 (O_853,N_21584,N_24558);
nor UO_854 (O_854,N_22591,N_23556);
or UO_855 (O_855,N_18827,N_22636);
nand UO_856 (O_856,N_19465,N_20807);
nand UO_857 (O_857,N_23102,N_22447);
nor UO_858 (O_858,N_20819,N_19550);
xnor UO_859 (O_859,N_23060,N_22288);
and UO_860 (O_860,N_22199,N_23200);
xnor UO_861 (O_861,N_19009,N_23022);
nor UO_862 (O_862,N_19597,N_23660);
xor UO_863 (O_863,N_23028,N_20434);
and UO_864 (O_864,N_18785,N_23819);
xor UO_865 (O_865,N_21655,N_19491);
nand UO_866 (O_866,N_22306,N_19510);
or UO_867 (O_867,N_24091,N_24685);
and UO_868 (O_868,N_19182,N_23507);
xnor UO_869 (O_869,N_21208,N_24497);
nor UO_870 (O_870,N_20310,N_24904);
nor UO_871 (O_871,N_21130,N_19110);
nor UO_872 (O_872,N_23503,N_23856);
nand UO_873 (O_873,N_19543,N_21795);
xor UO_874 (O_874,N_24349,N_19250);
or UO_875 (O_875,N_24872,N_22281);
and UO_876 (O_876,N_24964,N_20510);
nor UO_877 (O_877,N_22167,N_19521);
nor UO_878 (O_878,N_21708,N_20110);
and UO_879 (O_879,N_19082,N_23828);
xor UO_880 (O_880,N_22668,N_19738);
nand UO_881 (O_881,N_23431,N_19913);
nand UO_882 (O_882,N_23588,N_19730);
or UO_883 (O_883,N_21318,N_23612);
xnor UO_884 (O_884,N_22094,N_22241);
xnor UO_885 (O_885,N_24996,N_23945);
nand UO_886 (O_886,N_21591,N_24544);
xnor UO_887 (O_887,N_22089,N_18819);
xor UO_888 (O_888,N_21442,N_23296);
nand UO_889 (O_889,N_20331,N_19320);
nand UO_890 (O_890,N_21377,N_19291);
and UO_891 (O_891,N_18820,N_19462);
nand UO_892 (O_892,N_22600,N_24140);
and UO_893 (O_893,N_22284,N_19946);
or UO_894 (O_894,N_22871,N_21524);
xor UO_895 (O_895,N_24791,N_22439);
nand UO_896 (O_896,N_24153,N_20679);
nor UO_897 (O_897,N_22189,N_24156);
and UO_898 (O_898,N_20168,N_23415);
nand UO_899 (O_899,N_22651,N_24300);
nand UO_900 (O_900,N_24339,N_19725);
and UO_901 (O_901,N_23900,N_20894);
or UO_902 (O_902,N_19386,N_18878);
nor UO_903 (O_903,N_22340,N_23826);
and UO_904 (O_904,N_20816,N_21923);
xor UO_905 (O_905,N_23399,N_22900);
nor UO_906 (O_906,N_24759,N_22494);
and UO_907 (O_907,N_20978,N_19188);
nand UO_908 (O_908,N_23832,N_21712);
xor UO_909 (O_909,N_20803,N_20339);
nand UO_910 (O_910,N_21047,N_22321);
nand UO_911 (O_911,N_24308,N_24333);
or UO_912 (O_912,N_18930,N_22515);
and UO_913 (O_913,N_24919,N_19185);
nand UO_914 (O_914,N_24697,N_24575);
nand UO_915 (O_915,N_24819,N_21144);
nor UO_916 (O_916,N_20913,N_21938);
xor UO_917 (O_917,N_21646,N_23299);
nand UO_918 (O_918,N_23181,N_19516);
xor UO_919 (O_919,N_24221,N_18836);
xnor UO_920 (O_920,N_19756,N_22908);
nand UO_921 (O_921,N_19235,N_22174);
nor UO_922 (O_922,N_22137,N_22517);
or UO_923 (O_923,N_24134,N_19699);
nand UO_924 (O_924,N_22043,N_23791);
nor UO_925 (O_925,N_20424,N_20166);
nor UO_926 (O_926,N_19877,N_18975);
nand UO_927 (O_927,N_20971,N_19852);
nor UO_928 (O_928,N_21245,N_20009);
xnor UO_929 (O_929,N_20732,N_21571);
and UO_930 (O_930,N_24580,N_23434);
or UO_931 (O_931,N_20728,N_20022);
nand UO_932 (O_932,N_24285,N_21073);
xnor UO_933 (O_933,N_22060,N_20062);
nand UO_934 (O_934,N_19196,N_20752);
nor UO_935 (O_935,N_24830,N_24677);
and UO_936 (O_936,N_24413,N_20120);
nor UO_937 (O_937,N_24798,N_21446);
nor UO_938 (O_938,N_23848,N_20833);
and UO_939 (O_939,N_18918,N_20049);
xor UO_940 (O_940,N_23050,N_22993);
and UO_941 (O_941,N_22981,N_21054);
xor UO_942 (O_942,N_20315,N_22620);
xor UO_943 (O_943,N_23808,N_21096);
xnor UO_944 (O_944,N_20652,N_24019);
or UO_945 (O_945,N_21392,N_22203);
xor UO_946 (O_946,N_24949,N_18884);
and UO_947 (O_947,N_20808,N_21529);
xor UO_948 (O_948,N_21822,N_20991);
nor UO_949 (O_949,N_19598,N_19096);
and UO_950 (O_950,N_21121,N_19575);
or UO_951 (O_951,N_19636,N_19837);
xnor UO_952 (O_952,N_23463,N_19206);
or UO_953 (O_953,N_18929,N_21033);
or UO_954 (O_954,N_19078,N_22695);
nand UO_955 (O_955,N_19705,N_20271);
xnor UO_956 (O_956,N_21104,N_22206);
xor UO_957 (O_957,N_23081,N_23129);
or UO_958 (O_958,N_23849,N_20748);
or UO_959 (O_959,N_21572,N_20294);
and UO_960 (O_960,N_21828,N_23985);
xor UO_961 (O_961,N_19679,N_20615);
and UO_962 (O_962,N_20432,N_19564);
nand UO_963 (O_963,N_20319,N_19651);
nand UO_964 (O_964,N_24947,N_23783);
xor UO_965 (O_965,N_21512,N_19248);
nand UO_966 (O_966,N_19831,N_21695);
and UO_967 (O_967,N_22774,N_20313);
or UO_968 (O_968,N_23587,N_20536);
nand UO_969 (O_969,N_19167,N_23382);
nand UO_970 (O_970,N_22107,N_19442);
or UO_971 (O_971,N_21592,N_20772);
nor UO_972 (O_972,N_20541,N_20704);
nor UO_973 (O_973,N_21017,N_21278);
xnor UO_974 (O_974,N_22922,N_24487);
nor UO_975 (O_975,N_21410,N_23223);
and UO_976 (O_976,N_19284,N_20681);
or UO_977 (O_977,N_23938,N_19125);
and UO_978 (O_978,N_21538,N_19232);
xnor UO_979 (O_979,N_19026,N_21076);
nand UO_980 (O_980,N_24496,N_24674);
nor UO_981 (O_981,N_21855,N_20144);
or UO_982 (O_982,N_23678,N_19362);
nor UO_983 (O_983,N_24663,N_23630);
and UO_984 (O_984,N_20146,N_18844);
nand UO_985 (O_985,N_24158,N_22931);
xnor UO_986 (O_986,N_22783,N_20677);
nand UO_987 (O_987,N_20162,N_21833);
nor UO_988 (O_988,N_20912,N_24775);
nor UO_989 (O_989,N_23003,N_20332);
nand UO_990 (O_990,N_19828,N_19747);
or UO_991 (O_991,N_20755,N_24831);
nor UO_992 (O_992,N_21268,N_22581);
nand UO_993 (O_993,N_21155,N_19308);
nand UO_994 (O_994,N_23385,N_21336);
xnor UO_995 (O_995,N_21241,N_20394);
nor UO_996 (O_996,N_21643,N_20435);
and UO_997 (O_997,N_19051,N_22332);
nor UO_998 (O_998,N_24891,N_24119);
nor UO_999 (O_999,N_20038,N_24656);
or UO_1000 (O_1000,N_19139,N_23822);
nor UO_1001 (O_1001,N_19932,N_19459);
and UO_1002 (O_1002,N_21480,N_22696);
and UO_1003 (O_1003,N_20010,N_22192);
nor UO_1004 (O_1004,N_19286,N_21904);
and UO_1005 (O_1005,N_21454,N_21219);
and UO_1006 (O_1006,N_21840,N_23658);
and UO_1007 (O_1007,N_23554,N_18859);
and UO_1008 (O_1008,N_20201,N_20340);
xor UO_1009 (O_1009,N_23437,N_22543);
nor UO_1010 (O_1010,N_22170,N_20379);
nor UO_1011 (O_1011,N_22135,N_21063);
nor UO_1012 (O_1012,N_18916,N_22942);
xnor UO_1013 (O_1013,N_21842,N_20754);
or UO_1014 (O_1014,N_19147,N_20852);
nor UO_1015 (O_1015,N_21687,N_24391);
and UO_1016 (O_1016,N_23521,N_23417);
xor UO_1017 (O_1017,N_21779,N_19076);
nand UO_1018 (O_1018,N_24532,N_22124);
nand UO_1019 (O_1019,N_19498,N_23654);
or UO_1020 (O_1020,N_21999,N_24632);
nor UO_1021 (O_1021,N_19163,N_23365);
xnor UO_1022 (O_1022,N_20855,N_21058);
or UO_1023 (O_1023,N_21751,N_20725);
nor UO_1024 (O_1024,N_18933,N_18955);
xor UO_1025 (O_1025,N_21853,N_24486);
nand UO_1026 (O_1026,N_21222,N_21031);
nand UO_1027 (O_1027,N_20983,N_20874);
xnor UO_1028 (O_1028,N_19028,N_21699);
nor UO_1029 (O_1029,N_24952,N_24421);
and UO_1030 (O_1030,N_24159,N_22088);
and UO_1031 (O_1031,N_19201,N_19617);
nor UO_1032 (O_1032,N_19370,N_21817);
and UO_1033 (O_1033,N_20945,N_23571);
and UO_1034 (O_1034,N_20004,N_20335);
xnor UO_1035 (O_1035,N_22333,N_21244);
nand UO_1036 (O_1036,N_21304,N_22850);
or UO_1037 (O_1037,N_22215,N_23812);
and UO_1038 (O_1038,N_21652,N_23433);
nand UO_1039 (O_1039,N_24941,N_20351);
xnor UO_1040 (O_1040,N_23252,N_24992);
xnor UO_1041 (O_1041,N_24698,N_24281);
nor UO_1042 (O_1042,N_22421,N_22782);
xor UO_1043 (O_1043,N_19822,N_19729);
or UO_1044 (O_1044,N_24507,N_24284);
or UO_1045 (O_1045,N_20683,N_24865);
xnor UO_1046 (O_1046,N_20077,N_23939);
and UO_1047 (O_1047,N_21240,N_22086);
and UO_1048 (O_1048,N_23733,N_19031);
nand UO_1049 (O_1049,N_18924,N_22229);
nand UO_1050 (O_1050,N_19105,N_19780);
or UO_1051 (O_1051,N_20623,N_22706);
nor UO_1052 (O_1052,N_22845,N_20433);
or UO_1053 (O_1053,N_20300,N_18938);
nand UO_1054 (O_1054,N_24062,N_20883);
xnor UO_1055 (O_1055,N_20316,N_24347);
and UO_1056 (O_1056,N_21635,N_21300);
and UO_1057 (O_1057,N_19692,N_24013);
xor UO_1058 (O_1058,N_23558,N_24939);
and UO_1059 (O_1059,N_24696,N_21441);
and UO_1060 (O_1060,N_24440,N_21936);
or UO_1061 (O_1061,N_22812,N_22588);
xor UO_1062 (O_1062,N_21307,N_24586);
or UO_1063 (O_1063,N_20029,N_19224);
or UO_1064 (O_1064,N_24883,N_22687);
xor UO_1065 (O_1065,N_24270,N_22064);
xnor UO_1066 (O_1066,N_22397,N_21935);
nand UO_1067 (O_1067,N_18857,N_20785);
xnor UO_1068 (O_1068,N_21347,N_19093);
nand UO_1069 (O_1069,N_23641,N_20555);
nand UO_1070 (O_1070,N_24133,N_19383);
and UO_1071 (O_1071,N_24954,N_22736);
or UO_1072 (O_1072,N_19245,N_21942);
and UO_1073 (O_1073,N_21657,N_20179);
nand UO_1074 (O_1074,N_21827,N_21585);
xor UO_1075 (O_1075,N_24545,N_22420);
and UO_1076 (O_1076,N_21122,N_19998);
or UO_1077 (O_1077,N_22527,N_19050);
or UO_1078 (O_1078,N_19132,N_23002);
and UO_1079 (O_1079,N_21286,N_24548);
nand UO_1080 (O_1080,N_20064,N_19156);
nand UO_1081 (O_1081,N_20591,N_23924);
nor UO_1082 (O_1082,N_19231,N_20330);
nand UO_1083 (O_1083,N_23245,N_19171);
and UO_1084 (O_1084,N_23677,N_19959);
or UO_1085 (O_1085,N_19815,N_21495);
and UO_1086 (O_1086,N_22491,N_19976);
nand UO_1087 (O_1087,N_19757,N_19625);
nor UO_1088 (O_1088,N_19103,N_19228);
and UO_1089 (O_1089,N_22195,N_20761);
nand UO_1090 (O_1090,N_21289,N_21697);
or UO_1091 (O_1091,N_21554,N_19524);
and UO_1092 (O_1092,N_19591,N_23505);
or UO_1093 (O_1093,N_19351,N_24386);
xor UO_1094 (O_1094,N_20895,N_23462);
nor UO_1095 (O_1095,N_21234,N_21317);
and UO_1096 (O_1096,N_24000,N_22468);
and UO_1097 (O_1097,N_23005,N_22847);
or UO_1098 (O_1098,N_24854,N_21967);
nor UO_1099 (O_1099,N_20191,N_20580);
xor UO_1100 (O_1100,N_23023,N_22507);
nand UO_1101 (O_1101,N_21143,N_18874);
or UO_1102 (O_1102,N_21184,N_20159);
xnor UO_1103 (O_1103,N_22242,N_22893);
xnor UO_1104 (O_1104,N_24518,N_18812);
nand UO_1105 (O_1105,N_22451,N_23565);
and UO_1106 (O_1106,N_22178,N_19473);
and UO_1107 (O_1107,N_23756,N_24878);
nor UO_1108 (O_1108,N_24930,N_19980);
or UO_1109 (O_1109,N_21877,N_20176);
or UO_1110 (O_1110,N_20352,N_18759);
or UO_1111 (O_1111,N_19668,N_20782);
and UO_1112 (O_1112,N_18987,N_19255);
xor UO_1113 (O_1113,N_20042,N_23371);
and UO_1114 (O_1114,N_19800,N_24095);
and UO_1115 (O_1115,N_24169,N_23389);
nand UO_1116 (O_1116,N_19380,N_20914);
or UO_1117 (O_1117,N_24566,N_23747);
and UO_1118 (O_1118,N_22278,N_24011);
and UO_1119 (O_1119,N_23605,N_22096);
nor UO_1120 (O_1120,N_21022,N_23161);
nor UO_1121 (O_1121,N_22392,N_24694);
nand UO_1122 (O_1122,N_21215,N_23098);
and UO_1123 (O_1123,N_21787,N_22808);
nor UO_1124 (O_1124,N_20420,N_22290);
xor UO_1125 (O_1125,N_23817,N_21953);
nor UO_1126 (O_1126,N_19638,N_22230);
or UO_1127 (O_1127,N_24277,N_24666);
and UO_1128 (O_1128,N_24373,N_19396);
xor UO_1129 (O_1129,N_24806,N_20739);
nor UO_1130 (O_1130,N_21301,N_20165);
xor UO_1131 (O_1131,N_20214,N_19950);
xnor UO_1132 (O_1132,N_23234,N_21282);
nor UO_1133 (O_1133,N_22980,N_21472);
nor UO_1134 (O_1134,N_21332,N_19898);
nor UO_1135 (O_1135,N_23619,N_19137);
xnor UO_1136 (O_1136,N_19338,N_20469);
or UO_1137 (O_1137,N_20226,N_18798);
xnor UO_1138 (O_1138,N_19840,N_19683);
nor UO_1139 (O_1139,N_18867,N_20821);
nand UO_1140 (O_1140,N_20232,N_20412);
or UO_1141 (O_1141,N_24956,N_23862);
nand UO_1142 (O_1142,N_20130,N_22646);
and UO_1143 (O_1143,N_19635,N_22339);
and UO_1144 (O_1144,N_23305,N_19436);
nand UO_1145 (O_1145,N_22489,N_19761);
nor UO_1146 (O_1146,N_19272,N_22866);
xor UO_1147 (O_1147,N_21570,N_20641);
and UO_1148 (O_1148,N_20291,N_19606);
xnor UO_1149 (O_1149,N_24705,N_19294);
xor UO_1150 (O_1150,N_22431,N_20104);
or UO_1151 (O_1151,N_20929,N_21754);
and UO_1152 (O_1152,N_19676,N_19614);
nand UO_1153 (O_1153,N_21954,N_23540);
xor UO_1154 (O_1154,N_21294,N_20384);
nand UO_1155 (O_1155,N_19545,N_24915);
xor UO_1156 (O_1156,N_19149,N_19488);
nand UO_1157 (O_1157,N_21598,N_19654);
and UO_1158 (O_1158,N_20484,N_21260);
and UO_1159 (O_1159,N_21006,N_23631);
nand UO_1160 (O_1160,N_21195,N_20153);
nand UO_1161 (O_1161,N_21117,N_22536);
or UO_1162 (O_1162,N_21619,N_20257);
nor UO_1163 (O_1163,N_19014,N_18979);
or UO_1164 (O_1164,N_21388,N_24054);
and UO_1165 (O_1165,N_22834,N_23821);
xor UO_1166 (O_1166,N_24702,N_20947);
nand UO_1167 (O_1167,N_24342,N_21075);
nor UO_1168 (O_1168,N_20192,N_19991);
xor UO_1169 (O_1169,N_22841,N_19719);
or UO_1170 (O_1170,N_23340,N_22709);
and UO_1171 (O_1171,N_23127,N_24356);
xor UO_1172 (O_1172,N_20398,N_24522);
or UO_1173 (O_1173,N_22440,N_19414);
xor UO_1174 (O_1174,N_20127,N_23979);
and UO_1175 (O_1175,N_21693,N_20700);
xnor UO_1176 (O_1176,N_19714,N_21684);
xor UO_1177 (O_1177,N_21269,N_24974);
or UO_1178 (O_1178,N_19560,N_21390);
and UO_1179 (O_1179,N_23261,N_24746);
or UO_1180 (O_1180,N_24304,N_21478);
or UO_1181 (O_1181,N_24261,N_20618);
and UO_1182 (O_1182,N_19199,N_20878);
nor UO_1183 (O_1183,N_22765,N_22956);
nor UO_1184 (O_1184,N_23954,N_21026);
and UO_1185 (O_1185,N_24060,N_19472);
nand UO_1186 (O_1186,N_24275,N_24707);
or UO_1187 (O_1187,N_19933,N_20998);
nand UO_1188 (O_1188,N_19114,N_23006);
and UO_1189 (O_1189,N_19776,N_22294);
xor UO_1190 (O_1190,N_24438,N_18839);
xnor UO_1191 (O_1191,N_23914,N_24751);
and UO_1192 (O_1192,N_20825,N_20105);
or UO_1193 (O_1193,N_20582,N_24387);
and UO_1194 (O_1194,N_19611,N_23873);
nor UO_1195 (O_1195,N_18760,N_24044);
or UO_1196 (O_1196,N_22250,N_20178);
xnor UO_1197 (O_1197,N_23785,N_21202);
xor UO_1198 (O_1198,N_22844,N_23653);
nor UO_1199 (O_1199,N_22904,N_23575);
nand UO_1200 (O_1200,N_23320,N_21453);
xor UO_1201 (O_1201,N_24468,N_24292);
xor UO_1202 (O_1202,N_20879,N_24764);
or UO_1203 (O_1203,N_19895,N_19357);
and UO_1204 (O_1204,N_20596,N_19270);
xor UO_1205 (O_1205,N_24825,N_20703);
or UO_1206 (O_1206,N_21229,N_20664);
and UO_1207 (O_1207,N_24026,N_19519);
nor UO_1208 (O_1208,N_20245,N_20980);
nand UO_1209 (O_1209,N_24436,N_24980);
and UO_1210 (O_1210,N_22935,N_23872);
or UO_1211 (O_1211,N_20073,N_22685);
xnor UO_1212 (O_1212,N_20518,N_20362);
xnor UO_1213 (O_1213,N_19593,N_24733);
or UO_1214 (O_1214,N_23700,N_23221);
or UO_1215 (O_1215,N_20576,N_21847);
nand UO_1216 (O_1216,N_18751,N_24852);
or UO_1217 (O_1217,N_21557,N_21396);
nand UO_1218 (O_1218,N_22529,N_24072);
xor UO_1219 (O_1219,N_22589,N_21588);
xor UO_1220 (O_1220,N_23027,N_19733);
nor UO_1221 (O_1221,N_20353,N_23671);
and UO_1222 (O_1222,N_21417,N_20932);
nand UO_1223 (O_1223,N_24951,N_21103);
or UO_1224 (O_1224,N_24004,N_24903);
nor UO_1225 (O_1225,N_21380,N_22238);
and UO_1226 (O_1226,N_23366,N_23243);
nor UO_1227 (O_1227,N_22382,N_21177);
nor UO_1228 (O_1228,N_24771,N_24989);
nor UO_1229 (O_1229,N_21078,N_19891);
or UO_1230 (O_1230,N_19678,N_20944);
nand UO_1231 (O_1231,N_21138,N_21755);
nor UO_1232 (O_1232,N_19019,N_20875);
and UO_1233 (O_1233,N_23657,N_23475);
xor UO_1234 (O_1234,N_22514,N_24892);
nand UO_1235 (O_1235,N_21056,N_21932);
and UO_1236 (O_1236,N_19480,N_21998);
xnor UO_1237 (O_1237,N_22539,N_22342);
nor UO_1238 (O_1238,N_24732,N_23974);
or UO_1239 (O_1239,N_21258,N_18943);
and UO_1240 (O_1240,N_19903,N_21055);
nand UO_1241 (O_1241,N_20438,N_20958);
or UO_1242 (O_1242,N_20336,N_20012);
nand UO_1243 (O_1243,N_23219,N_20654);
xor UO_1244 (O_1244,N_23090,N_21642);
nor UO_1245 (O_1245,N_20707,N_21974);
and UO_1246 (O_1246,N_19358,N_22131);
and UO_1247 (O_1247,N_22890,N_24898);
or UO_1248 (O_1248,N_22327,N_22911);
xnor UO_1249 (O_1249,N_23251,N_22185);
nand UO_1250 (O_1250,N_24070,N_23450);
or UO_1251 (O_1251,N_22073,N_24849);
and UO_1252 (O_1252,N_21361,N_22035);
and UO_1253 (O_1253,N_19476,N_22590);
xnor UO_1254 (O_1254,N_20813,N_23950);
and UO_1255 (O_1255,N_24803,N_19432);
xnor UO_1256 (O_1256,N_21906,N_22183);
xnor UO_1257 (O_1257,N_19920,N_21716);
nor UO_1258 (O_1258,N_22181,N_20547);
and UO_1259 (O_1259,N_24085,N_19159);
xnor UO_1260 (O_1260,N_23043,N_24839);
or UO_1261 (O_1261,N_24441,N_21761);
xor UO_1262 (O_1262,N_24176,N_18873);
and UO_1263 (O_1263,N_22804,N_23229);
nand UO_1264 (O_1264,N_20637,N_18899);
nor UO_1265 (O_1265,N_20814,N_22315);
xor UO_1266 (O_1266,N_22180,N_19345);
or UO_1267 (O_1267,N_20281,N_20632);
or UO_1268 (O_1268,N_20033,N_21190);
or UO_1269 (O_1269,N_23322,N_20382);
nand UO_1270 (O_1270,N_21447,N_24537);
and UO_1271 (O_1271,N_24418,N_20613);
or UO_1272 (O_1272,N_19214,N_18973);
or UO_1273 (O_1273,N_22996,N_24667);
nand UO_1274 (O_1274,N_24003,N_18970);
nor UO_1275 (O_1275,N_22478,N_19770);
nor UO_1276 (O_1276,N_22211,N_20674);
xnor UO_1277 (O_1277,N_23577,N_23666);
xnor UO_1278 (O_1278,N_22492,N_24455);
and UO_1279 (O_1279,N_19194,N_21326);
and UO_1280 (O_1280,N_21084,N_21854);
and UO_1281 (O_1281,N_22326,N_19955);
xor UO_1282 (O_1282,N_21407,N_21800);
or UO_1283 (O_1283,N_23061,N_22110);
and UO_1284 (O_1284,N_22711,N_24165);
nor UO_1285 (O_1285,N_19337,N_20626);
nor UO_1286 (O_1286,N_22384,N_22401);
nand UO_1287 (O_1287,N_19869,N_23100);
xor UO_1288 (O_1288,N_19097,N_19894);
or UO_1289 (O_1289,N_20496,N_23743);
nor UO_1290 (O_1290,N_24307,N_23542);
and UO_1291 (O_1291,N_22508,N_20777);
or UO_1292 (O_1292,N_19158,N_20994);
nor UO_1293 (O_1293,N_24633,N_20071);
and UO_1294 (O_1294,N_20083,N_20820);
or UO_1295 (O_1295,N_21542,N_21246);
nand UO_1296 (O_1296,N_20118,N_20578);
xor UO_1297 (O_1297,N_20036,N_20699);
nor UO_1298 (O_1298,N_20051,N_22545);
xor UO_1299 (O_1299,N_23773,N_19789);
xnor UO_1300 (O_1300,N_24205,N_23451);
or UO_1301 (O_1301,N_22903,N_20666);
and UO_1302 (O_1302,N_19400,N_20740);
or UO_1303 (O_1303,N_19489,N_19716);
xor UO_1304 (O_1304,N_22679,N_22079);
nor UO_1305 (O_1305,N_23274,N_20269);
or UO_1306 (O_1306,N_23611,N_19426);
nand UO_1307 (O_1307,N_24234,N_21660);
xor UO_1308 (O_1308,N_24726,N_20174);
or UO_1309 (O_1309,N_24048,N_20590);
and UO_1310 (O_1310,N_19528,N_22253);
nand UO_1311 (O_1311,N_22619,N_22062);
nor UO_1312 (O_1312,N_24729,N_21349);
or UO_1313 (O_1313,N_22435,N_19470);
xor UO_1314 (O_1314,N_23012,N_22443);
nor UO_1315 (O_1315,N_24423,N_19349);
or UO_1316 (O_1316,N_21000,N_21262);
xor UO_1317 (O_1317,N_22388,N_21443);
and UO_1318 (O_1318,N_21381,N_18786);
or UO_1319 (O_1319,N_21577,N_21634);
and UO_1320 (O_1320,N_20723,N_24100);
xor UO_1321 (O_1321,N_23490,N_22635);
xnor UO_1322 (O_1322,N_19931,N_22789);
xor UO_1323 (O_1323,N_19871,N_22822);
or UO_1324 (O_1324,N_21996,N_24840);
nand UO_1325 (O_1325,N_24291,N_20393);
nand UO_1326 (O_1326,N_19122,N_18761);
and UO_1327 (O_1327,N_23731,N_23037);
nand UO_1328 (O_1328,N_22065,N_21128);
and UO_1329 (O_1329,N_24020,N_21628);
and UO_1330 (O_1330,N_21213,N_23032);
or UO_1331 (O_1331,N_19118,N_19970);
xnor UO_1332 (O_1332,N_19372,N_23600);
and UO_1333 (O_1333,N_24016,N_23622);
or UO_1334 (O_1334,N_21342,N_22905);
nand UO_1335 (O_1335,N_20301,N_18823);
nand UO_1336 (O_1336,N_20458,N_22623);
xor UO_1337 (O_1337,N_19275,N_22777);
xnor UO_1338 (O_1338,N_19886,N_22201);
nand UO_1339 (O_1339,N_24331,N_21263);
xor UO_1340 (O_1340,N_20465,N_19711);
xnor UO_1341 (O_1341,N_24034,N_22754);
or UO_1342 (O_1342,N_19556,N_21989);
nand UO_1343 (O_1343,N_21661,N_24485);
xnor UO_1344 (O_1344,N_23978,N_18984);
and UO_1345 (O_1345,N_21801,N_21949);
or UO_1346 (O_1346,N_23847,N_20597);
nor UO_1347 (O_1347,N_22349,N_20198);
xor UO_1348 (O_1348,N_21072,N_22748);
and UO_1349 (O_1349,N_23368,N_23777);
nand UO_1350 (O_1350,N_19257,N_24439);
and UO_1351 (O_1351,N_21374,N_20774);
and UO_1352 (O_1352,N_20303,N_20734);
nor UO_1353 (O_1353,N_23645,N_22283);
or UO_1354 (O_1354,N_19999,N_22264);
nor UO_1355 (O_1355,N_22002,N_23455);
nor UO_1356 (O_1356,N_19387,N_22571);
nand UO_1357 (O_1357,N_20992,N_24320);
nand UO_1358 (O_1358,N_23943,N_22407);
xnor UO_1359 (O_1359,N_21338,N_19005);
nand UO_1360 (O_1360,N_22633,N_21824);
and UO_1361 (O_1361,N_20250,N_19486);
nor UO_1362 (O_1362,N_19064,N_21231);
and UO_1363 (O_1363,N_23511,N_23044);
xnor UO_1364 (O_1364,N_23277,N_19077);
nand UO_1365 (O_1365,N_22032,N_20988);
nor UO_1366 (O_1366,N_23140,N_19283);
nand UO_1367 (O_1367,N_20445,N_23333);
or UO_1368 (O_1368,N_21225,N_23632);
or UO_1369 (O_1369,N_23801,N_19296);
or UO_1370 (O_1370,N_20150,N_21858);
nand UO_1371 (O_1371,N_21691,N_22305);
or UO_1372 (O_1372,N_21792,N_19157);
or UO_1373 (O_1373,N_20139,N_22851);
and UO_1374 (O_1374,N_20069,N_22858);
nor UO_1375 (O_1375,N_22481,N_19830);
xnor UO_1376 (O_1376,N_20592,N_21163);
and UO_1377 (O_1377,N_22759,N_19285);
or UO_1378 (O_1378,N_21940,N_24306);
nor UO_1379 (O_1379,N_21537,N_22563);
nor UO_1380 (O_1380,N_18906,N_20222);
or UO_1381 (O_1381,N_21036,N_23236);
nand UO_1382 (O_1382,N_24886,N_19726);
xor UO_1383 (O_1383,N_20621,N_19325);
and UO_1384 (O_1384,N_18880,N_24922);
or UO_1385 (O_1385,N_24405,N_22204);
nand UO_1386 (O_1386,N_23403,N_22882);
nand UO_1387 (O_1387,N_23762,N_23769);
xnor UO_1388 (O_1388,N_20346,N_18996);
nand UO_1389 (O_1389,N_20024,N_20920);
xnor UO_1390 (O_1390,N_20718,N_22912);
and UO_1391 (O_1391,N_19347,N_19660);
nor UO_1392 (O_1392,N_20670,N_21040);
xor UO_1393 (O_1393,N_21702,N_23529);
nand UO_1394 (O_1394,N_21686,N_23697);
nand UO_1395 (O_1395,N_23078,N_21962);
or UO_1396 (O_1396,N_19605,N_19576);
or UO_1397 (O_1397,N_19628,N_19680);
nor UO_1398 (O_1398,N_24652,N_23313);
nor UO_1399 (O_1399,N_23695,N_21271);
nand UO_1400 (O_1400,N_23738,N_24600);
nand UO_1401 (O_1401,N_19454,N_21802);
xnor UO_1402 (O_1402,N_21713,N_20143);
and UO_1403 (O_1403,N_22246,N_24341);
xnor UO_1404 (O_1404,N_20369,N_22212);
or UO_1405 (O_1405,N_19977,N_20129);
xor UO_1406 (O_1406,N_20461,N_23837);
xor UO_1407 (O_1407,N_20695,N_19236);
and UO_1408 (O_1408,N_19855,N_22797);
or UO_1409 (O_1409,N_22580,N_20671);
or UO_1410 (O_1410,N_20631,N_23516);
and UO_1411 (O_1411,N_19018,N_21945);
or UO_1412 (O_1412,N_24946,N_19751);
xor UO_1413 (O_1413,N_22833,N_21165);
and UO_1414 (O_1414,N_21624,N_19728);
nor UO_1415 (O_1415,N_20934,N_19779);
xnor UO_1416 (O_1416,N_22296,N_20959);
and UO_1417 (O_1417,N_24800,N_23664);
xor UO_1418 (O_1418,N_19344,N_21653);
and UO_1419 (O_1419,N_23977,N_22361);
or UO_1420 (O_1420,N_24533,N_19376);
nand UO_1421 (O_1421,N_18828,N_20600);
xor UO_1422 (O_1422,N_23213,N_19823);
nand UO_1423 (O_1423,N_23811,N_21829);
and UO_1424 (O_1424,N_20343,N_23248);
and UO_1425 (O_1425,N_20968,N_23624);
nand UO_1426 (O_1426,N_21965,N_20520);
nor UO_1427 (O_1427,N_21362,N_18989);
and UO_1428 (O_1428,N_22254,N_21310);
nor UO_1429 (O_1429,N_21007,N_23499);
or UO_1430 (O_1430,N_23910,N_19269);
or UO_1431 (O_1431,N_21576,N_22813);
or UO_1432 (O_1432,N_21750,N_20831);
and UO_1433 (O_1433,N_19145,N_21492);
or UO_1434 (O_1434,N_21672,N_18908);
and UO_1435 (O_1435,N_23494,N_19948);
and UO_1436 (O_1436,N_19784,N_19072);
and UO_1437 (O_1437,N_21663,N_22585);
nand UO_1438 (O_1438,N_24503,N_24216);
nor UO_1439 (O_1439,N_19736,N_22968);
nor UO_1440 (O_1440,N_24902,N_19142);
nand UO_1441 (O_1441,N_19864,N_22737);
nor UO_1442 (O_1442,N_24488,N_18953);
nor UO_1443 (O_1443,N_23732,N_19434);
nand UO_1444 (O_1444,N_19085,N_19450);
and UO_1445 (O_1445,N_23509,N_22302);
nand UO_1446 (O_1446,N_24354,N_19341);
and UO_1447 (O_1447,N_20838,N_20537);
nor UO_1448 (O_1448,N_24037,N_19315);
nand UO_1449 (O_1449,N_20727,N_21516);
nand UO_1450 (O_1450,N_19596,N_22551);
nor UO_1451 (O_1451,N_23445,N_21564);
and UO_1452 (O_1452,N_22899,N_20937);
xnor UO_1453 (O_1453,N_21203,N_18811);
nor UO_1454 (O_1454,N_19463,N_18765);
xnor UO_1455 (O_1455,N_21395,N_24646);
and UO_1456 (O_1456,N_22609,N_21863);
or UO_1457 (O_1457,N_18926,N_19493);
nor UO_1458 (O_1458,N_21189,N_23613);
nor UO_1459 (O_1459,N_22786,N_23550);
nand UO_1460 (O_1460,N_23625,N_19658);
xnor UO_1461 (O_1461,N_20877,N_18923);
nand UO_1462 (O_1462,N_22962,N_23470);
nor UO_1463 (O_1463,N_22453,N_19406);
and UO_1464 (O_1464,N_19217,N_23405);
xor UO_1465 (O_1465,N_21376,N_19586);
or UO_1466 (O_1466,N_24525,N_23278);
xnor UO_1467 (O_1467,N_24265,N_23356);
nand UO_1468 (O_1468,N_23206,N_18824);
xnor UO_1469 (O_1469,N_22486,N_19212);
xor UO_1470 (O_1470,N_20533,N_21790);
and UO_1471 (O_1471,N_21705,N_18945);
or UO_1472 (O_1472,N_19943,N_21608);
or UO_1473 (O_1473,N_22208,N_22733);
and UO_1474 (O_1474,N_20479,N_20531);
and UO_1475 (O_1475,N_20850,N_19403);
nor UO_1476 (O_1476,N_21815,N_22511);
nor UO_1477 (O_1477,N_20298,N_22602);
nand UO_1478 (O_1478,N_21913,N_22944);
or UO_1479 (O_1479,N_22232,N_23291);
nor UO_1480 (O_1480,N_24311,N_23761);
nor UO_1481 (O_1481,N_21857,N_23926);
nor UO_1482 (O_1482,N_23205,N_20365);
xnor UO_1483 (O_1483,N_23956,N_22669);
and UO_1484 (O_1484,N_23114,N_20203);
nor UO_1485 (O_1485,N_24394,N_19900);
or UO_1486 (O_1486,N_21814,N_24047);
nand UO_1487 (O_1487,N_23723,N_23539);
and UO_1488 (O_1488,N_22516,N_21905);
nor UO_1489 (O_1489,N_19769,N_22838);
nor UO_1490 (O_1490,N_23203,N_22556);
and UO_1491 (O_1491,N_21881,N_22892);
or UO_1492 (O_1492,N_24096,N_19496);
or UO_1493 (O_1493,N_22091,N_22111);
or UO_1494 (O_1494,N_21323,N_23413);
nand UO_1495 (O_1495,N_20385,N_24460);
nor UO_1496 (O_1496,N_18897,N_23838);
nor UO_1497 (O_1497,N_22112,N_21982);
nor UO_1498 (O_1498,N_20733,N_20884);
nand UO_1499 (O_1499,N_19530,N_23286);
or UO_1500 (O_1500,N_24966,N_19508);
or UO_1501 (O_1501,N_19000,N_19845);
nand UO_1502 (O_1502,N_24040,N_24912);
and UO_1503 (O_1503,N_20890,N_23301);
xor UO_1504 (O_1504,N_22757,N_19128);
nand UO_1505 (O_1505,N_19429,N_24206);
xor UO_1506 (O_1506,N_20091,N_21927);
xnor UO_1507 (O_1507,N_23578,N_19619);
xor UO_1508 (O_1508,N_21809,N_24998);
nor UO_1509 (O_1509,N_21723,N_19116);
xor UO_1510 (O_1510,N_19032,N_23789);
nor UO_1511 (O_1511,N_21647,N_18805);
nand UO_1512 (O_1512,N_19100,N_19901);
and UO_1513 (O_1513,N_19882,N_23497);
nand UO_1514 (O_1514,N_21559,N_23139);
and UO_1515 (O_1515,N_24241,N_19546);
nor UO_1516 (O_1516,N_21340,N_22120);
xor UO_1517 (O_1517,N_22474,N_20145);
nor UO_1518 (O_1518,N_19838,N_19401);
or UO_1519 (O_1519,N_21357,N_19071);
nor UO_1520 (O_1520,N_24945,N_19238);
and UO_1521 (O_1521,N_19618,N_19456);
and UO_1522 (O_1522,N_18763,N_23017);
nor UO_1523 (O_1523,N_20020,N_19204);
xor UO_1524 (O_1524,N_20229,N_19183);
nor UO_1525 (O_1525,N_21217,N_21988);
and UO_1526 (O_1526,N_21583,N_19007);
nor UO_1527 (O_1527,N_23517,N_18766);
nor UO_1528 (O_1528,N_24430,N_22601);
or UO_1529 (O_1529,N_23861,N_21658);
nor UO_1530 (O_1530,N_21601,N_19888);
and UO_1531 (O_1531,N_23884,N_23110);
nand UO_1532 (O_1532,N_20950,N_19902);
or UO_1533 (O_1533,N_21711,N_23594);
nor UO_1534 (O_1534,N_23429,N_24756);
nand UO_1535 (O_1535,N_19663,N_23538);
nor UO_1536 (O_1536,N_24230,N_22325);
nor UO_1537 (O_1537,N_21438,N_23720);
nor UO_1538 (O_1538,N_22016,N_19492);
xnor UO_1539 (O_1539,N_20231,N_21888);
or UO_1540 (O_1540,N_19924,N_20569);
and UO_1541 (O_1541,N_19333,N_22746);
or UO_1542 (O_1542,N_24101,N_22724);
and UO_1543 (O_1543,N_19444,N_23549);
xnor UO_1544 (O_1544,N_23960,N_23136);
nand UO_1545 (O_1545,N_24647,N_20722);
and UO_1546 (O_1546,N_24410,N_24620);
xor UO_1547 (O_1547,N_24790,N_22047);
or UO_1548 (O_1548,N_23336,N_20830);
nor UO_1549 (O_1549,N_23486,N_19313);
nand UO_1550 (O_1550,N_22156,N_23827);
nor UO_1551 (O_1551,N_18791,N_22731);
nand UO_1552 (O_1552,N_20368,N_21560);
or UO_1553 (O_1553,N_18863,N_24139);
nand UO_1554 (O_1554,N_22691,N_22228);
xor UO_1555 (O_1555,N_19282,N_22832);
nand UO_1556 (O_1556,N_22902,N_22568);
xnor UO_1557 (O_1557,N_18968,N_20995);
or UO_1558 (O_1558,N_21543,N_24480);
nand UO_1559 (O_1559,N_18768,N_20263);
or UO_1560 (O_1560,N_24380,N_24021);
nor UO_1561 (O_1561,N_20485,N_21423);
or UO_1562 (O_1562,N_24490,N_21742);
nor UO_1563 (O_1563,N_23784,N_24662);
or UO_1564 (O_1564,N_22082,N_24570);
xnor UO_1565 (O_1565,N_22336,N_21893);
and UO_1566 (O_1566,N_23069,N_20548);
and UO_1567 (O_1567,N_19604,N_20114);
nor UO_1568 (O_1568,N_19280,N_21645);
xnor UO_1569 (O_1569,N_22226,N_19752);
and UO_1570 (O_1570,N_21316,N_23753);
and UO_1571 (O_1571,N_22629,N_20730);
and UO_1572 (O_1572,N_19038,N_23300);
or UO_1573 (O_1573,N_19956,N_24990);
nand UO_1574 (O_1574,N_21595,N_21637);
nor UO_1575 (O_1575,N_23987,N_24985);
or UO_1576 (O_1576,N_20358,N_19439);
nand UO_1577 (O_1577,N_20169,N_23332);
or UO_1578 (O_1578,N_21759,N_22499);
or UO_1579 (O_1579,N_21462,N_19704);
xnor UO_1580 (O_1580,N_21694,N_21142);
nand UO_1581 (O_1581,N_24619,N_22345);
or UO_1582 (O_1582,N_21079,N_19853);
nor UO_1583 (O_1583,N_22785,N_19399);
and UO_1584 (O_1584,N_19123,N_19870);
xor UO_1585 (O_1585,N_22068,N_19419);
and UO_1586 (O_1586,N_24569,N_20417);
nand UO_1587 (O_1587,N_24443,N_18856);
xor UO_1588 (O_1588,N_20251,N_22105);
xor UO_1589 (O_1589,N_21798,N_19954);
or UO_1590 (O_1590,N_24193,N_19319);
xor UO_1591 (O_1591,N_21373,N_24464);
nand UO_1592 (O_1592,N_21251,N_24714);
or UO_1593 (O_1593,N_20701,N_21622);
and UO_1594 (O_1594,N_20375,N_23237);
or UO_1595 (O_1595,N_24876,N_22723);
and UO_1596 (O_1596,N_21420,N_23020);
nand UO_1597 (O_1597,N_24092,N_20858);
and UO_1598 (O_1598,N_20503,N_21261);
xnor UO_1599 (O_1599,N_20943,N_20312);
xnor UO_1600 (O_1600,N_23359,N_19579);
or UO_1601 (O_1601,N_22550,N_20282);
xnor UO_1602 (O_1602,N_19522,N_19589);
nor UO_1603 (O_1603,N_21216,N_21867);
and UO_1604 (O_1604,N_19515,N_24837);
nor UO_1605 (O_1605,N_24847,N_20919);
and UO_1606 (O_1606,N_20512,N_20900);
xnor UO_1607 (O_1607,N_23551,N_23360);
nor UO_1608 (O_1608,N_23851,N_22191);
and UO_1609 (O_1609,N_24109,N_21600);
xnor UO_1610 (O_1610,N_21832,N_20519);
nand UO_1611 (O_1611,N_20429,N_22565);
or UO_1612 (O_1612,N_24074,N_19834);
nor UO_1613 (O_1613,N_21627,N_24727);
nand UO_1614 (O_1614,N_19303,N_21964);
nor UO_1615 (O_1615,N_24736,N_20014);
xor UO_1616 (O_1616,N_23427,N_21549);
or UO_1617 (O_1617,N_22261,N_23552);
or UO_1618 (O_1618,N_21920,N_20568);
nand UO_1619 (O_1619,N_23262,N_21620);
nand UO_1620 (O_1620,N_24608,N_20771);
nand UO_1621 (O_1621,N_20135,N_21180);
nor UO_1622 (O_1622,N_21012,N_21247);
xor UO_1623 (O_1623,N_20812,N_23642);
nand UO_1624 (O_1624,N_24175,N_21980);
nand UO_1625 (O_1625,N_22184,N_19549);
nor UO_1626 (O_1626,N_24416,N_23688);
nand UO_1627 (O_1627,N_23547,N_24093);
xnor UO_1628 (O_1628,N_19554,N_24520);
xor UO_1629 (O_1629,N_22788,N_21514);
or UO_1630 (O_1630,N_18998,N_24360);
or UO_1631 (O_1631,N_23046,N_20302);
and UO_1632 (O_1632,N_19879,N_22173);
or UO_1633 (O_1633,N_20586,N_24493);
and UO_1634 (O_1634,N_18941,N_19440);
nor UO_1635 (O_1635,N_20673,N_21449);
or UO_1636 (O_1636,N_18800,N_20341);
nand UO_1637 (O_1637,N_21264,N_23614);
or UO_1638 (O_1638,N_18853,N_22081);
nor UO_1639 (O_1639,N_23390,N_23815);
and UO_1640 (O_1640,N_21014,N_22835);
nor UO_1641 (O_1641,N_21728,N_20923);
or UO_1642 (O_1642,N_21043,N_22448);
nand UO_1643 (O_1643,N_22626,N_23831);
xnor UO_1644 (O_1644,N_23443,N_24454);
nor UO_1645 (O_1645,N_23537,N_23758);
nand UO_1646 (O_1646,N_19379,N_21295);
or UO_1647 (O_1647,N_24772,N_22661);
nand UO_1648 (O_1648,N_18851,N_19873);
and UO_1649 (O_1649,N_21211,N_20538);
or UO_1650 (O_1650,N_20296,N_23311);
xor UO_1651 (O_1651,N_19762,N_20446);
nor UO_1652 (O_1652,N_21837,N_22704);
xnor UO_1653 (O_1653,N_19155,N_22099);
xnor UO_1654 (O_1654,N_24752,N_22941);
nor UO_1655 (O_1655,N_24038,N_23372);
or UO_1656 (O_1656,N_23991,N_23941);
nand UO_1657 (O_1657,N_24809,N_20400);
and UO_1658 (O_1658,N_22320,N_24742);
or UO_1659 (O_1659,N_22829,N_22055);
nand UO_1660 (O_1660,N_23944,N_23883);
xnor UO_1661 (O_1661,N_19062,N_22402);
nor UO_1662 (O_1662,N_19474,N_18849);
and UO_1663 (O_1663,N_20016,N_24881);
and UO_1664 (O_1664,N_22273,N_23106);
nor UO_1665 (O_1665,N_24258,N_21299);
nor UO_1666 (O_1666,N_20019,N_24539);
and UO_1667 (O_1667,N_24587,N_18804);
or UO_1668 (O_1668,N_23923,N_23797);
nor UO_1669 (O_1669,N_21547,N_19346);
and UO_1670 (O_1670,N_18866,N_19251);
nor UO_1671 (O_1671,N_19552,N_24512);
xnor UO_1672 (O_1672,N_24145,N_23211);
xor UO_1673 (O_1673,N_20387,N_20306);
xnor UO_1674 (O_1674,N_20745,N_19246);
xnor UO_1675 (O_1675,N_20411,N_24542);
or UO_1676 (O_1676,N_19334,N_18808);
and UO_1677 (O_1677,N_19410,N_24971);
nand UO_1678 (O_1678,N_24718,N_23216);
nor UO_1679 (O_1679,N_23699,N_21891);
or UO_1680 (O_1680,N_24722,N_24154);
and UO_1681 (O_1681,N_19469,N_23934);
nand UO_1682 (O_1682,N_19412,N_24115);
xor UO_1683 (O_1683,N_22126,N_20116);
nand UO_1684 (O_1684,N_24433,N_23370);
nor UO_1685 (O_1685,N_19017,N_24254);
and UO_1686 (O_1686,N_23246,N_20267);
and UO_1687 (O_1687,N_23396,N_21312);
and UO_1688 (O_1688,N_20786,N_20783);
and UO_1689 (O_1689,N_21736,N_20194);
and UO_1690 (O_1690,N_23188,N_23224);
xor UO_1691 (O_1691,N_20680,N_20440);
nand UO_1692 (O_1692,N_24228,N_20388);
or UO_1693 (O_1693,N_22006,N_23727);
xor UO_1694 (O_1694,N_19583,N_20948);
and UO_1695 (O_1695,N_24152,N_20690);
nand UO_1696 (O_1696,N_21201,N_22839);
or UO_1697 (O_1697,N_20901,N_23596);
or UO_1698 (O_1698,N_19487,N_22823);
or UO_1699 (O_1699,N_20355,N_24296);
nor UO_1700 (O_1700,N_21993,N_21520);
and UO_1701 (O_1701,N_22125,N_20067);
nor UO_1702 (O_1702,N_19501,N_21275);
nand UO_1703 (O_1703,N_19221,N_19385);
nand UO_1704 (O_1704,N_24717,N_22937);
nand UO_1705 (O_1705,N_19630,N_22769);
nor UO_1706 (O_1706,N_20505,N_19648);
xnor UO_1707 (O_1707,N_21562,N_19378);
nor UO_1708 (O_1708,N_20357,N_20324);
nand UO_1709 (O_1709,N_22013,N_20742);
or UO_1710 (O_1710,N_21431,N_24266);
or UO_1711 (O_1711,N_21013,N_20620);
and UO_1712 (O_1712,N_22144,N_22427);
nand UO_1713 (O_1713,N_22188,N_23796);
nor UO_1714 (O_1714,N_21329,N_21135);
nand UO_1715 (O_1715,N_24235,N_22583);
nand UO_1716 (O_1716,N_23649,N_24259);
xor UO_1717 (O_1717,N_22821,N_22939);
and UO_1718 (O_1718,N_20635,N_20088);
xnor UO_1719 (O_1719,N_18793,N_23790);
xor UO_1720 (O_1720,N_24924,N_20930);
nand UO_1721 (O_1721,N_21133,N_19909);
nor UO_1722 (O_1722,N_23334,N_22671);
nand UO_1723 (O_1723,N_20523,N_18887);
nor UO_1724 (O_1724,N_20952,N_21257);
xor UO_1725 (O_1725,N_23879,N_21283);
nand UO_1726 (O_1726,N_21690,N_22352);
and UO_1727 (O_1727,N_22889,N_20906);
nor UO_1728 (O_1728,N_19104,N_24588);
xor UO_1729 (O_1729,N_19448,N_23492);
and UO_1730 (O_1730,N_23887,N_22160);
and UO_1731 (O_1731,N_18782,N_18949);
nor UO_1732 (O_1732,N_23981,N_24147);
xor UO_1733 (O_1733,N_19811,N_23141);
and UO_1734 (O_1734,N_23317,N_21947);
or UO_1735 (O_1735,N_23546,N_22625);
and UO_1736 (O_1736,N_20649,N_21673);
and UO_1737 (O_1737,N_22728,N_20847);
nor UO_1738 (O_1738,N_21334,N_24317);
or UO_1739 (O_1739,N_23901,N_21963);
nor UO_1740 (O_1740,N_20180,N_24491);
or UO_1741 (O_1741,N_24851,N_21255);
xnor UO_1742 (O_1742,N_21327,N_20076);
and UO_1743 (O_1743,N_22268,N_19690);
or UO_1744 (O_1744,N_24848,N_20973);
nor UO_1745 (O_1745,N_21089,N_21164);
or UO_1746 (O_1746,N_23996,N_23230);
nor UO_1747 (O_1747,N_24893,N_24461);
nor UO_1748 (O_1748,N_22220,N_22059);
nor UO_1749 (O_1749,N_24596,N_23288);
xnor UO_1750 (O_1750,N_19613,N_24802);
xnor UO_1751 (O_1751,N_20946,N_21518);
and UO_1752 (O_1752,N_23284,N_22473);
xnor UO_1753 (O_1753,N_24427,N_18803);
or UO_1754 (O_1754,N_21080,N_23843);
nor UO_1755 (O_1755,N_23388,N_21667);
and UO_1756 (O_1756,N_22140,N_23062);
xnor UO_1757 (O_1757,N_19798,N_24838);
or UO_1758 (O_1758,N_23019,N_21298);
and UO_1759 (O_1759,N_20039,N_18845);
nand UO_1760 (O_1760,N_22837,N_21024);
and UO_1761 (O_1761,N_19993,N_21777);
xor UO_1762 (O_1762,N_21871,N_19037);
nor UO_1763 (O_1763,N_21958,N_23927);
or UO_1764 (O_1764,N_23563,N_24940);
xor UO_1765 (O_1765,N_21147,N_21424);
and UO_1766 (O_1766,N_19542,N_24110);
nand UO_1767 (O_1767,N_24182,N_23103);
nor UO_1768 (O_1768,N_23447,N_21136);
nor UO_1769 (O_1769,N_23599,N_24597);
xor UO_1770 (O_1770,N_21976,N_22664);
xnor UO_1771 (O_1771,N_20285,N_23609);
xor UO_1772 (O_1772,N_22157,N_22573);
or UO_1773 (O_1773,N_22643,N_23561);
nand UO_1774 (O_1774,N_23086,N_23319);
nand UO_1775 (O_1775,N_19940,N_24777);
nand UO_1776 (O_1776,N_18928,N_21230);
nand UO_1777 (O_1777,N_23112,N_19856);
and UO_1778 (O_1778,N_24552,N_19988);
nor UO_1779 (O_1779,N_22256,N_19863);
nand UO_1780 (O_1780,N_20476,N_23998);
nor UO_1781 (O_1781,N_24276,N_21368);
nand UO_1782 (O_1782,N_23541,N_22505);
nand UO_1783 (O_1783,N_20491,N_24622);
nor UO_1784 (O_1784,N_19054,N_23568);
nor UO_1785 (O_1785,N_21489,N_22090);
xnor UO_1786 (O_1786,N_24249,N_21869);
nor UO_1787 (O_1787,N_23802,N_20188);
xnor UO_1788 (O_1788,N_24198,N_20345);
nor UO_1789 (O_1789,N_19866,N_22360);
or UO_1790 (O_1790,N_22924,N_24884);
and UO_1791 (O_1791,N_22561,N_24866);
and UO_1792 (O_1792,N_21335,N_24725);
nor UO_1793 (O_1793,N_24210,N_19814);
or UO_1794 (O_1794,N_19669,N_19290);
nor UO_1795 (O_1795,N_20818,N_21649);
xor UO_1796 (O_1796,N_23287,N_21924);
and UO_1797 (O_1797,N_19293,N_20381);
or UO_1798 (O_1798,N_18771,N_19722);
nor UO_1799 (O_1799,N_22214,N_21483);
and UO_1800 (O_1800,N_23807,N_22040);
nand UO_1801 (O_1801,N_23693,N_20075);
nor UO_1802 (O_1802,N_21578,N_20685);
and UO_1803 (O_1803,N_22083,N_22351);
nor UO_1804 (O_1804,N_20514,N_24132);
xnor UO_1805 (O_1805,N_20246,N_23227);
and UO_1806 (O_1806,N_21851,N_24469);
or UO_1807 (O_1807,N_23176,N_19230);
nand UO_1808 (O_1808,N_24185,N_24720);
nand UO_1809 (O_1809,N_22408,N_24267);
xor UO_1810 (O_1810,N_21944,N_19200);
xor UO_1811 (O_1811,N_19020,N_19807);
or UO_1812 (O_1812,N_20243,N_20824);
nand UO_1813 (O_1813,N_24888,N_21091);
or UO_1814 (O_1814,N_20103,N_22469);
nor UO_1815 (O_1815,N_23869,N_22639);
or UO_1816 (O_1816,N_20487,N_24162);
or UO_1817 (O_1817,N_23681,N_24077);
and UO_1818 (O_1818,N_20138,N_22738);
xor UO_1819 (O_1819,N_22210,N_21360);
xnor UO_1820 (O_1820,N_23474,N_21678);
xor UO_1821 (O_1821,N_22784,N_20187);
nand UO_1822 (O_1822,N_24282,N_19574);
nor UO_1823 (O_1823,N_24719,N_20573);
nor UO_1824 (O_1824,N_23917,N_20131);
or UO_1825 (O_1825,N_22586,N_19039);
nand UO_1826 (O_1826,N_20097,N_19395);
nor UO_1827 (O_1827,N_19889,N_22484);
nor UO_1828 (O_1828,N_24398,N_24799);
xor UO_1829 (O_1829,N_20669,N_21580);
or UO_1830 (O_1830,N_22077,N_24972);
nor UO_1831 (O_1831,N_24724,N_20377);
nor UO_1832 (O_1832,N_24870,N_20442);
and UO_1833 (O_1833,N_21596,N_22106);
xor UO_1834 (O_1834,N_24982,N_23369);
xnor UO_1835 (O_1835,N_19915,N_21154);
nor UO_1836 (O_1836,N_21876,N_23395);
nand UO_1837 (O_1837,N_23350,N_24058);
nor UO_1838 (O_1838,N_24933,N_22915);
nand UO_1839 (O_1839,N_20941,N_23407);
nand UO_1840 (O_1840,N_20581,N_18750);
nor UO_1841 (O_1841,N_18787,N_24383);
xor UO_1842 (O_1842,N_23526,N_20773);
and UO_1843 (O_1843,N_21726,N_24009);
or UO_1844 (O_1844,N_23617,N_23155);
and UO_1845 (O_1845,N_24278,N_23107);
xor UO_1846 (O_1846,N_24942,N_19350);
and UO_1847 (O_1847,N_21440,N_20516);
and UO_1848 (O_1848,N_21188,N_21227);
or UO_1849 (O_1849,N_21494,N_21049);
nor UO_1850 (O_1850,N_20195,N_19706);
nor UO_1851 (O_1851,N_23736,N_20587);
and UO_1852 (O_1852,N_21768,N_24826);
nand UO_1853 (O_1853,N_24257,N_24094);
nor UO_1854 (O_1854,N_24397,N_20534);
nor UO_1855 (O_1855,N_18891,N_19003);
nand UO_1856 (O_1856,N_22952,N_24064);
nand UO_1857 (O_1857,N_19253,N_21599);
and UO_1858 (O_1858,N_21003,N_21237);
nand UO_1859 (O_1859,N_22328,N_23472);
xor UO_1860 (O_1860,N_24834,N_22237);
or UO_1861 (O_1861,N_22959,N_18896);
or UO_1862 (O_1862,N_24700,N_24084);
nand UO_1863 (O_1863,N_23269,N_20034);
or UO_1864 (O_1864,N_24289,N_21021);
xnor UO_1865 (O_1865,N_19670,N_24332);
xor UO_1866 (O_1866,N_20295,N_23298);
nor UO_1867 (O_1867,N_23672,N_20322);
and UO_1868 (O_1868,N_18756,N_19513);
or UO_1869 (O_1869,N_24328,N_19053);
nand UO_1870 (O_1870,N_20171,N_18752);
nand UO_1871 (O_1871,N_22364,N_22857);
nor UO_1872 (O_1872,N_22989,N_20544);
or UO_1873 (O_1873,N_22914,N_24935);
nand UO_1874 (O_1874,N_23729,N_18910);
xnor UO_1875 (O_1875,N_22594,N_21901);
nand UO_1876 (O_1876,N_21774,N_23895);
or UO_1877 (O_1877,N_20563,N_20835);
xor UO_1878 (O_1878,N_23416,N_21527);
or UO_1879 (O_1879,N_24022,N_19740);
xor UO_1880 (O_1880,N_23567,N_20241);
or UO_1881 (O_1881,N_24385,N_24814);
xnor UO_1882 (O_1882,N_18997,N_20235);
or UO_1883 (O_1883,N_23074,N_21192);
xor UO_1884 (O_1884,N_23099,N_21094);
or UO_1885 (O_1885,N_20283,N_23875);
nor UO_1886 (O_1886,N_20498,N_21688);
nand UO_1887 (O_1887,N_18999,N_24561);
xnor UO_1888 (O_1888,N_21398,N_20528);
xor UO_1889 (O_1889,N_23329,N_19402);
nand UO_1890 (O_1890,N_24484,N_21413);
nor UO_1891 (O_1891,N_19369,N_24821);
and UO_1892 (O_1892,N_22806,N_24918);
nand UO_1893 (O_1893,N_22618,N_20158);
xor UO_1894 (O_1894,N_22627,N_22224);
nor UO_1895 (O_1895,N_22957,N_19836);
or UO_1896 (O_1896,N_22700,N_18810);
and UO_1897 (O_1897,N_23573,N_24243);
nand UO_1898 (O_1898,N_24492,N_23075);
xnor UO_1899 (O_1899,N_19033,N_18907);
nor UO_1900 (O_1900,N_22853,N_24255);
and UO_1901 (O_1901,N_18773,N_24984);
and UO_1902 (O_1902,N_21330,N_20770);
nor UO_1903 (O_1903,N_24467,N_21745);
and UO_1904 (O_1904,N_20598,N_20747);
and UO_1905 (O_1905,N_24555,N_24873);
and UO_1906 (O_1906,N_20604,N_21083);
nand UO_1907 (O_1907,N_21223,N_20975);
and UO_1908 (O_1908,N_18807,N_24177);
nand UO_1909 (O_1909,N_20902,N_24395);
nor UO_1910 (O_1910,N_19584,N_23256);
xor UO_1911 (O_1911,N_22592,N_21151);
and UO_1912 (O_1912,N_22604,N_20363);
or UO_1913 (O_1913,N_20712,N_20694);
and UO_1914 (O_1914,N_20840,N_22359);
and UO_1915 (O_1915,N_20493,N_19266);
xor UO_1916 (O_1916,N_22542,N_22429);
xnor UO_1917 (O_1917,N_20616,N_18831);
xor UO_1918 (O_1918,N_23754,N_20405);
or UO_1919 (O_1919,N_21886,N_23198);
nor UO_1920 (O_1920,N_19143,N_23629);
xnor UO_1921 (O_1921,N_22334,N_20996);
nand UO_1922 (O_1922,N_22024,N_20378);
or UO_1923 (O_1923,N_24991,N_20482);
xnor UO_1924 (O_1924,N_23341,N_22973);
nand UO_1925 (O_1925,N_19675,N_21469);
and UO_1926 (O_1926,N_21358,N_21541);
xor UO_1927 (O_1927,N_22800,N_19192);
nand UO_1928 (O_1928,N_24710,N_20702);
xor UO_1929 (O_1929,N_23337,N_22218);
xor UO_1930 (O_1930,N_22414,N_21504);
or UO_1931 (O_1931,N_21703,N_20170);
nor UO_1932 (O_1932,N_22849,N_20452);
and UO_1933 (O_1933,N_23418,N_19983);
and UO_1934 (O_1934,N_19471,N_19365);
or UO_1935 (O_1935,N_24583,N_19621);
xnor UO_1936 (O_1936,N_24670,N_22555);
or UO_1937 (O_1937,N_24519,N_23342);
nor UO_1938 (O_1938,N_19322,N_24179);
xor UO_1939 (O_1939,N_22567,N_24412);
xor UO_1940 (O_1940,N_24168,N_22391);
nand UO_1941 (O_1941,N_20321,N_20645);
nand UO_1942 (O_1942,N_23304,N_24755);
xor UO_1943 (O_1943,N_24896,N_20154);
nand UO_1944 (O_1944,N_20199,N_22526);
or UO_1945 (O_1945,N_19608,N_20778);
or UO_1946 (O_1946,N_20273,N_22309);
xnor UO_1947 (O_1947,N_20986,N_23094);
nor UO_1948 (O_1948,N_20967,N_19963);
nor UO_1949 (O_1949,N_20063,N_22128);
and UO_1950 (O_1950,N_20636,N_23696);
xnor UO_1951 (O_1951,N_20553,N_24462);
nand UO_1952 (O_1952,N_19570,N_24200);
nand UO_1953 (O_1953,N_23072,N_21615);
xnor UO_1954 (O_1954,N_23663,N_19558);
nor UO_1955 (O_1955,N_23710,N_20888);
nor UO_1956 (O_1956,N_18858,N_23635);
nor UO_1957 (O_1957,N_20237,N_22301);
nor UO_1958 (O_1958,N_19041,N_18818);
nor UO_1959 (O_1959,N_24014,N_24024);
and UO_1960 (O_1960,N_19563,N_19225);
or UO_1961 (O_1961,N_20656,N_24678);
and UO_1962 (O_1962,N_20841,N_24402);
nor UO_1963 (O_1963,N_22071,N_23792);
nor UO_1964 (O_1964,N_18825,N_21910);
or UO_1965 (O_1965,N_19744,N_21186);
nor UO_1966 (O_1966,N_21303,N_22795);
or UO_1967 (O_1967,N_23518,N_20753);
nor UO_1968 (O_1968,N_22780,N_24031);
or UO_1969 (O_1969,N_21523,N_20667);
nor UO_1970 (O_1970,N_19388,N_22415);
nor UO_1971 (O_1971,N_20486,N_20471);
xor UO_1972 (O_1972,N_20836,N_19443);
xor UO_1973 (O_1973,N_24028,N_19664);
and UO_1974 (O_1974,N_19816,N_20050);
or UO_1975 (O_1975,N_22898,N_22410);
and UO_1976 (O_1976,N_18877,N_23835);
nor UO_1977 (O_1977,N_22816,N_23513);
and UO_1978 (O_1978,N_20489,N_24889);
xnor UO_1979 (O_1979,N_24593,N_19960);
and UO_1980 (O_1980,N_22307,N_19941);
or UO_1981 (O_1981,N_24909,N_24066);
xnor UO_1982 (O_1982,N_24711,N_23355);
xnor UO_1983 (O_1983,N_21016,N_19273);
nand UO_1984 (O_1984,N_21254,N_22805);
xor UO_1985 (O_1985,N_21957,N_24471);
xor UO_1986 (O_1986,N_24910,N_22122);
and UO_1987 (O_1987,N_23564,N_20464);
or UO_1988 (O_1988,N_18775,N_20364);
or UO_1989 (O_1989,N_24987,N_18806);
and UO_1990 (O_1990,N_20606,N_20577);
nand UO_1991 (O_1991,N_20416,N_24327);
and UO_1992 (O_1992,N_21337,N_23684);
nand UO_1993 (O_1993,N_19314,N_22108);
nor UO_1994 (O_1994,N_21445,N_20797);
or UO_1995 (O_1995,N_24184,N_22118);
xor UO_1996 (O_1996,N_22297,N_19195);
and UO_1997 (O_1997,N_19205,N_20186);
and UO_1998 (O_1998,N_20970,N_22574);
and UO_1999 (O_1999,N_21019,N_20472);
nor UO_2000 (O_2000,N_23436,N_24827);
nor UO_2001 (O_2001,N_19686,N_19923);
xor UO_2002 (O_2002,N_22236,N_24163);
nand UO_2003 (O_2003,N_19084,N_24207);
xor UO_2004 (O_2004,N_20676,N_21922);
and UO_2005 (O_2005,N_24644,N_21848);
xor UO_2006 (O_2006,N_22888,N_19352);
or UO_2007 (O_2007,N_24334,N_23750);
xnor UO_2008 (O_2008,N_19404,N_19944);
and UO_2009 (O_2009,N_23182,N_22923);
xor UO_2010 (O_2010,N_21831,N_23495);
and UO_2011 (O_2011,N_19634,N_24559);
nor UO_2012 (O_2012,N_24131,N_23548);
nor UO_2013 (O_2013,N_20072,N_19907);
or UO_2014 (O_2014,N_22467,N_20802);
nand UO_2015 (O_2015,N_24465,N_22652);
and UO_2016 (O_2016,N_18795,N_20953);
nor UO_2017 (O_2017,N_21956,N_20288);
and UO_2018 (O_2018,N_21385,N_24378);
nand UO_2019 (O_2019,N_20453,N_24796);
nor UO_2020 (O_2020,N_20376,N_21556);
nor UO_2021 (O_2021,N_20107,N_24370);
nor UO_2022 (O_2022,N_23643,N_21511);
xor UO_2023 (O_2023,N_19536,N_20494);
nor UO_2024 (O_2024,N_18895,N_20625);
nor UO_2025 (O_2025,N_21823,N_22234);
xnor UO_2026 (O_2026,N_22313,N_23133);
nor UO_2027 (O_2027,N_22701,N_22852);
xnor UO_2028 (O_2028,N_24953,N_18838);
xnor UO_2029 (O_2029,N_21162,N_20570);
nand UO_2030 (O_2030,N_20280,N_24426);
or UO_2031 (O_2031,N_18813,N_22919);
and UO_2032 (O_2032,N_20190,N_22920);
and UO_2033 (O_2033,N_21508,N_21486);
nand UO_2034 (O_2034,N_19511,N_23810);
xnor UO_2035 (O_2035,N_19324,N_24605);
and UO_2036 (O_2036,N_24781,N_19384);
or UO_2037 (O_2037,N_21836,N_23321);
xor UO_2038 (O_2038,N_20979,N_23180);
nand UO_2039 (O_2039,N_22498,N_19989);
nand UO_2040 (O_2040,N_22150,N_22482);
nand UO_2041 (O_2041,N_22277,N_18965);
and UO_2042 (O_2042,N_24734,N_23866);
xor UO_2043 (O_2043,N_20172,N_20002);
xor UO_2044 (O_2044,N_20735,N_23877);
or UO_2045 (O_2045,N_20981,N_24171);
xnor UO_2046 (O_2046,N_21302,N_20719);
xnor UO_2047 (O_2047,N_21066,N_21743);
nor UO_2048 (O_2048,N_21548,N_24018);
or UO_2049 (O_2049,N_19766,N_21256);
and UO_2050 (O_2050,N_23628,N_24628);
nand UO_2051 (O_2051,N_21365,N_19117);
nand UO_2052 (O_2052,N_23574,N_23925);
and UO_2053 (O_2053,N_20068,N_22308);
or UO_2054 (O_2054,N_18801,N_19538);
and UO_2055 (O_2055,N_21819,N_20843);
xor UO_2056 (O_2056,N_20768,N_19222);
nand UO_2057 (O_2057,N_24502,N_19010);
xnor UO_2058 (O_2058,N_20795,N_19304);
nand UO_2059 (O_2059,N_22874,N_20262);
and UO_2060 (O_2060,N_22803,N_18892);
xnor UO_2061 (O_2061,N_19086,N_23157);
nor UO_2062 (O_2062,N_24457,N_21280);
or UO_2063 (O_2063,N_22285,N_23467);
and UO_2064 (O_2064,N_24783,N_23240);
xor UO_2065 (O_2065,N_24824,N_18764);
or UO_2066 (O_2066,N_24639,N_23378);
or UO_2067 (O_2067,N_24995,N_21032);
xnor UO_2068 (O_2068,N_24624,N_21539);
nand UO_2069 (O_2069,N_23491,N_19021);
or UO_2070 (O_2070,N_19047,N_24483);
or UO_2071 (O_2071,N_19227,N_20459);
nor UO_2072 (O_2072,N_24563,N_21757);
or UO_2073 (O_2073,N_22537,N_24868);
or UO_2074 (O_2074,N_23674,N_24658);
or UO_2075 (O_2075,N_20234,N_24591);
or UO_2076 (O_2076,N_20040,N_22227);
or UO_2077 (O_2077,N_23717,N_21375);
xor UO_2078 (O_2078,N_23199,N_23152);
xor UO_2079 (O_2079,N_20515,N_21028);
or UO_2080 (O_2080,N_19223,N_19092);
nor UO_2081 (O_2081,N_24638,N_22293);
or UO_2082 (O_2082,N_22992,N_19753);
nand UO_2083 (O_2083,N_24116,N_23590);
xnor UO_2084 (O_2084,N_22824,N_22883);
nand UO_2085 (O_2085,N_21433,N_24735);
xor UO_2086 (O_2086,N_24680,N_19375);
nor UO_2087 (O_2087,N_19764,N_20880);
nor UO_2088 (O_2088,N_22843,N_20207);
or UO_2089 (O_2089,N_22779,N_20437);
nor UO_2090 (O_2090,N_24429,N_21674);
xnor UO_2091 (O_2091,N_20359,N_24689);
nor UO_2092 (O_2092,N_21946,N_23725);
nand UO_2093 (O_2093,N_24815,N_23339);
or UO_2094 (O_2094,N_23120,N_21288);
and UO_2095 (O_2095,N_24521,N_21493);
xnor UO_2096 (O_2096,N_20392,N_18956);
nand UO_2097 (O_2097,N_20749,N_24832);
and UO_2098 (O_2098,N_22647,N_19478);
xor UO_2099 (O_2099,N_23204,N_24635);
nand UO_2100 (O_2100,N_22751,N_20611);
or UO_2101 (O_2101,N_23257,N_19694);
nand UO_2102 (O_2102,N_22840,N_22182);
nor UO_2103 (O_2103,N_19974,N_20794);
xnor UO_2104 (O_2104,N_21394,N_22770);
xor UO_2105 (O_2105,N_24290,N_24403);
nor UO_2106 (O_2106,N_23247,N_20506);
xnor UO_2107 (O_2107,N_23308,N_21558);
and UO_2108 (O_2108,N_19847,N_21389);
and UO_2109 (O_2109,N_19996,N_19639);
nor UO_2110 (O_2110,N_20225,N_23846);
xnor UO_2111 (O_2111,N_19042,N_22579);
nand UO_2112 (O_2112,N_22916,N_21865);
xnor UO_2113 (O_2113,N_24607,N_18821);
or UO_2114 (O_2114,N_24452,N_21046);
or UO_2115 (O_2115,N_24273,N_18894);
or UO_2116 (O_2116,N_20684,N_19301);
nor UO_2117 (O_2117,N_20646,N_21344);
and UO_2118 (O_2118,N_23297,N_22548);
or UO_2119 (O_2119,N_22799,N_20942);
or UO_2120 (O_2120,N_20314,N_21782);
nand UO_2121 (O_2121,N_20788,N_20286);
or UO_2122 (O_2122,N_22383,N_23560);
and UO_2123 (O_2123,N_24379,N_22424);
or UO_2124 (O_2124,N_20798,N_24793);
xor UO_2125 (O_2125,N_24194,N_22863);
and UO_2126 (O_2126,N_19746,N_23059);
or UO_2127 (O_2127,N_18988,N_20399);
xor UO_2128 (O_2128,N_24141,N_23993);
nand UO_2129 (O_2129,N_19785,N_23374);
nor UO_2130 (O_2130,N_24219,N_19112);
nand UO_2131 (O_2131,N_19632,N_22544);
xnor UO_2132 (O_2132,N_22177,N_18792);
nor UO_2133 (O_2133,N_19449,N_24664);
xor UO_2134 (O_2134,N_18833,N_22930);
or UO_2135 (O_2135,N_21105,N_23080);
or UO_2136 (O_2136,N_21994,N_18932);
xnor UO_2137 (O_2137,N_18872,N_22005);
and UO_2138 (O_2138,N_21594,N_24779);
or UO_2139 (O_2139,N_24812,N_21866);
xor UO_2140 (O_2140,N_24260,N_19154);
nand UO_2141 (O_2141,N_22938,N_22151);
nor UO_2142 (O_2142,N_20872,N_24245);
or UO_2143 (O_2143,N_23508,N_22572);
xnor UO_2144 (O_2144,N_23973,N_24103);
nor UO_2145 (O_2145,N_24081,N_20149);
xnor UO_2146 (O_2146,N_23806,N_24083);
nand UO_2147 (O_2147,N_24527,N_19696);
nor UO_2148 (O_2148,N_20714,N_22485);
and UO_2149 (O_2149,N_20605,N_18865);
xor UO_2150 (O_2150,N_23220,N_20751);
xnor UO_2151 (O_2151,N_24765,N_21804);
nor UO_2152 (O_2152,N_21567,N_24679);
or UO_2153 (O_2153,N_22152,N_20085);
nor UO_2154 (O_2154,N_21709,N_19106);
nand UO_2155 (O_2155,N_23130,N_23576);
or UO_2156 (O_2156,N_22974,N_22217);
nand UO_2157 (O_2157,N_24030,N_24773);
xor UO_2158 (O_2158,N_20249,N_23468);
nand UO_2159 (O_2159,N_19832,N_24458);
nor UO_2160 (O_2160,N_21052,N_24218);
xor UO_2161 (O_2161,N_22932,N_24932);
nor UO_2162 (O_2162,N_21862,N_21010);
xnor UO_2163 (O_2163,N_23424,N_19499);
xor UO_2164 (O_2164,N_23408,N_20215);
or UO_2165 (O_2165,N_24050,N_24841);
or UO_2166 (O_2166,N_19146,N_20853);
nand UO_2167 (O_2167,N_22165,N_21515);
or UO_2168 (O_2168,N_19415,N_23905);
or UO_2169 (O_2169,N_22008,N_21669);
xor UO_2170 (O_2170,N_22462,N_23952);
nand UO_2171 (O_2171,N_20829,N_19582);
nor UO_2172 (O_2172,N_21035,N_22163);
or UO_2173 (O_2173,N_22798,N_19935);
and UO_2174 (O_2174,N_19457,N_23310);
nand UO_2175 (O_2175,N_21221,N_20691);
nor UO_2176 (O_2176,N_19773,N_20000);
or UO_2177 (O_2177,N_24478,N_21771);
or UO_2178 (O_2178,N_20037,N_23306);
or UO_2179 (O_2179,N_21057,N_23618);
nand UO_2180 (O_2180,N_24355,N_24869);
and UO_2181 (O_2181,N_19317,N_23244);
xor UO_2182 (O_2182,N_20366,N_24950);
nand UO_2183 (O_2183,N_22628,N_19809);
nor UO_2184 (O_2184,N_22856,N_23160);
nand UO_2185 (O_2185,N_21632,N_23484);
nor UO_2186 (O_2186,N_23442,N_24042);
or UO_2187 (O_2187,N_20675,N_22141);
nand UO_2188 (O_2188,N_22456,N_24712);
and UO_2189 (O_2189,N_23338,N_19793);
nand UO_2190 (O_2190,N_23177,N_23894);
nor UO_2191 (O_2191,N_19089,N_22501);
and UO_2192 (O_2192,N_23164,N_19452);
nand UO_2193 (O_2193,N_24978,N_22244);
xor UO_2194 (O_2194,N_24959,N_23117);
and UO_2195 (O_2195,N_19115,N_19278);
nand UO_2196 (O_2196,N_20951,N_19081);
nor UO_2197 (O_2197,N_19842,N_22001);
nor UO_2198 (O_2198,N_23669,N_19502);
and UO_2199 (O_2199,N_20638,N_23936);
nor UO_2200 (O_2200,N_19710,N_20954);
nand UO_2201 (O_2201,N_20522,N_18914);
nor UO_2202 (O_2202,N_21860,N_20834);
nor UO_2203 (O_2203,N_20045,N_22138);
or UO_2204 (O_2204,N_24143,N_24371);
or UO_2205 (O_2205,N_20687,N_23036);
nor UO_2206 (O_2206,N_21158,N_24778);
nand UO_2207 (O_2207,N_21140,N_23881);
nand UO_2208 (O_2208,N_24748,N_22521);
and UO_2209 (O_2209,N_21607,N_19490);
nand UO_2210 (O_2210,N_23995,N_22533);
xor UO_2211 (O_2211,N_20087,N_24411);
nand UO_2212 (O_2212,N_18850,N_22690);
or UO_2213 (O_2213,N_22022,N_23818);
or UO_2214 (O_2214,N_21265,N_23652);
or UO_2215 (O_2215,N_22300,N_19929);
nor UO_2216 (O_2216,N_21272,N_20466);
or UO_2217 (O_2217,N_23067,N_18915);
xor UO_2218 (O_2218,N_20765,N_21233);
nor UO_2219 (O_2219,N_19735,N_20408);
or UO_2220 (O_2220,N_23651,N_23779);
and UO_2221 (O_2221,N_20457,N_19849);
nand UO_2222 (O_2222,N_19531,N_23335);
nor UO_2223 (O_2223,N_21403,N_20255);
nor UO_2224 (O_2224,N_24238,N_23686);
nor UO_2225 (O_2225,N_24314,N_21510);
or UO_2226 (O_2226,N_23095,N_22036);
or UO_2227 (O_2227,N_22358,N_22790);
xor UO_2228 (O_2228,N_20662,N_20842);
and UO_2229 (O_2229,N_24404,N_23303);
xnor UO_2230 (O_2230,N_19887,N_22513);
nor UO_2231 (O_2231,N_18864,N_22423);
nand UO_2232 (O_2232,N_19724,N_20882);
nor UO_2233 (O_2233,N_20460,N_22272);
nand UO_2234 (O_2234,N_19997,N_19013);
and UO_2235 (O_2235,N_21193,N_23166);
and UO_2236 (O_2236,N_19063,N_24348);
nand UO_2237 (O_2237,N_23626,N_21343);
nand UO_2238 (O_2238,N_19083,N_21568);
xor UO_2239 (O_2239,N_19108,N_19681);
nand UO_2240 (O_2240,N_20776,N_20758);
nor UO_2241 (O_2241,N_23920,N_24293);
or UO_2242 (O_2242,N_19321,N_19525);
or UO_2243 (O_2243,N_19833,N_22641);
and UO_2244 (O_2244,N_23327,N_23836);
xor UO_2245 (O_2245,N_19537,N_23586);
nor UO_2246 (O_2246,N_19750,N_20513);
xnor UO_2247 (O_2247,N_19922,N_22142);
or UO_2248 (O_2248,N_21631,N_20867);
xnor UO_2249 (O_2249,N_24268,N_24005);
nor UO_2250 (O_2250,N_19181,N_19994);
and UO_2251 (O_2251,N_24012,N_21266);
nand UO_2252 (O_2252,N_23268,N_24082);
and UO_2253 (O_2253,N_22512,N_23544);
xor UO_2254 (O_2254,N_19962,N_21739);
and UO_2255 (O_2255,N_24075,N_24885);
or UO_2256 (O_2256,N_24654,N_22495);
and UO_2257 (O_2257,N_23522,N_21320);
and UO_2258 (O_2258,N_23400,N_23712);
and UO_2259 (O_2259,N_23823,N_23724);
and UO_2260 (O_2260,N_24250,N_23422);
nor UO_2261 (O_2261,N_20059,N_23940);
xor UO_2262 (O_2262,N_21587,N_20579);
and UO_2263 (O_2263,N_20289,N_19731);
nand UO_2264 (O_2264,N_22665,N_21696);
nor UO_2265 (O_2265,N_24247,N_23942);
and UO_2266 (O_2266,N_18942,N_20551);
nand UO_2267 (O_2267,N_21331,N_19446);
xnor UO_2268 (O_2268,N_24069,N_19609);
nor UO_2269 (O_2269,N_22067,N_23478);
nor UO_2270 (O_2270,N_24916,N_23593);
xnor UO_2271 (O_2271,N_23154,N_22781);
nor UO_2272 (O_2272,N_24811,N_19794);
and UO_2273 (O_2273,N_22610,N_21378);
or UO_2274 (O_2274,N_21500,N_22221);
nor UO_2275 (O_2275,N_23085,N_19569);
and UO_2276 (O_2276,N_23922,N_19949);
nor UO_2277 (O_2277,N_22946,N_20274);
or UO_2278 (O_2278,N_20211,N_20907);
nand UO_2279 (O_2279,N_22179,N_19631);
and UO_2280 (O_2280,N_19616,N_19417);
and UO_2281 (O_2281,N_22276,N_19787);
and UO_2282 (O_2282,N_24287,N_21350);
nor UO_2283 (O_2283,N_22520,N_24046);
nor UO_2284 (O_2284,N_22357,N_22965);
xor UO_2285 (O_2285,N_22139,N_23646);
nand UO_2286 (O_2286,N_20189,N_19862);
xor UO_2287 (O_2287,N_20966,N_24123);
nand UO_2288 (O_2288,N_20279,N_24170);
and UO_2289 (O_2289,N_24135,N_23039);
and UO_2290 (O_2290,N_24318,N_20630);
or UO_2291 (O_2291,N_22470,N_19423);
and UO_2292 (O_2292,N_19518,N_19512);
or UO_2293 (O_2293,N_20893,N_19557);
and UO_2294 (O_2294,N_23294,N_24890);
and UO_2295 (O_2295,N_21629,N_21506);
and UO_2296 (O_2296,N_22490,N_20093);
nand UO_2297 (O_2297,N_19307,N_23212);
and UO_2298 (O_2298,N_20532,N_23583);
or UO_2299 (O_2299,N_23128,N_19102);
nand UO_2300 (O_2300,N_24948,N_22606);
or UO_2301 (O_2301,N_24695,N_22341);
nor UO_2302 (O_2302,N_19759,N_20594);
nand UO_2303 (O_2303,N_24027,N_21120);
or UO_2304 (O_2304,N_19161,N_20356);
and UO_2305 (O_2305,N_22605,N_21626);
xnor UO_2306 (O_2306,N_20862,N_24616);
or UO_2307 (O_2307,N_21681,N_22136);
or UO_2308 (O_2308,N_24223,N_20708);
and UO_2309 (O_2309,N_18948,N_20724);
xnor UO_2310 (O_2310,N_24196,N_24071);
and UO_2311 (O_2311,N_20475,N_24237);
xnor UO_2312 (O_2312,N_23159,N_24816);
nor UO_2313 (O_2313,N_19985,N_22732);
nand UO_2314 (O_2314,N_21894,N_23373);
and UO_2315 (O_2315,N_21071,N_19287);
nor UO_2316 (O_2316,N_23640,N_22917);
nor UO_2317 (O_2317,N_21106,N_20839);
or UO_2318 (O_2318,N_19987,N_21107);
nor UO_2319 (O_2319,N_23994,N_20268);
and UO_2320 (O_2320,N_19044,N_24121);
nor UO_2321 (O_2321,N_24045,N_21972);
nor UO_2322 (O_2322,N_21725,N_22027);
or UO_2323 (O_2323,N_18814,N_23683);
xor UO_2324 (O_2324,N_20559,N_18832);
xor UO_2325 (O_2325,N_22519,N_19529);
and UO_2326 (O_2326,N_21903,N_23093);
and UO_2327 (O_2327,N_18840,N_23928);
nor UO_2328 (O_2328,N_22198,N_20043);
xor UO_2329 (O_2329,N_20259,N_23279);
and UO_2330 (O_2330,N_19795,N_19306);
xnor UO_2331 (O_2331,N_23770,N_21579);
nand UO_2332 (O_2332,N_23891,N_22599);
nand UO_2333 (O_2333,N_21134,N_19363);
and UO_2334 (O_2334,N_24229,N_19259);
or UO_2335 (O_2335,N_21285,N_24509);
nor UO_2336 (O_2336,N_24526,N_23685);
nor UO_2337 (O_2337,N_22050,N_21281);
and UO_2338 (O_2338,N_24144,N_23101);
nor UO_2339 (O_2339,N_20253,N_23850);
nand UO_2340 (O_2340,N_22403,N_24225);
xnor UO_2341 (O_2341,N_19036,N_23704);
and UO_2342 (O_2342,N_19709,N_24148);
and UO_2343 (O_2343,N_23958,N_19727);
or UO_2344 (O_2344,N_21810,N_18802);
nor UO_2345 (O_2345,N_22886,N_22506);
nand UO_2346 (O_2346,N_22240,N_20609);
and UO_2347 (O_2347,N_22977,N_20585);
and UO_2348 (O_2348,N_19986,N_22365);
xnor UO_2349 (O_2349,N_24967,N_23990);
nand UO_2350 (O_2350,N_21296,N_21092);
xnor UO_2351 (O_2351,N_24969,N_22775);
nand UO_2352 (O_2352,N_18936,N_22145);
nand UO_2353 (O_2353,N_21884,N_24572);
xor UO_2354 (O_2354,N_20860,N_24117);
or UO_2355 (O_2355,N_20572,N_22712);
or UO_2356 (O_2356,N_24079,N_24204);
nor UO_2357 (O_2357,N_19169,N_18902);
xnor UO_2358 (O_2358,N_22504,N_20648);
xnor UO_2359 (O_2359,N_24693,N_19332);
or UO_2360 (O_2360,N_23874,N_23648);
nand UO_2361 (O_2361,N_22380,N_22044);
and UO_2362 (O_2362,N_21528,N_20419);
nor UO_2363 (O_2363,N_24390,N_23766);
and UO_2364 (O_2364,N_19281,N_24157);
xnor UO_2365 (O_2365,N_22114,N_18888);
nand UO_2366 (O_2366,N_21826,N_19087);
nor UO_2367 (O_2367,N_22045,N_24274);
nand UO_2368 (O_2368,N_23748,N_23045);
and UO_2369 (O_2369,N_22963,N_24977);
xnor UO_2370 (O_2370,N_22502,N_23582);
nor UO_2371 (O_2371,N_24937,N_19390);
and UO_2372 (O_2372,N_23719,N_19938);
or UO_2373 (O_2373,N_21476,N_19804);
nand UO_2374 (O_2374,N_20448,N_23183);
and UO_2375 (O_2375,N_22479,N_24025);
nand UO_2376 (O_2376,N_23555,N_21065);
and UO_2377 (O_2377,N_22873,N_20240);
or UO_2378 (O_2378,N_22820,N_22353);
xor UO_2379 (O_2379,N_22762,N_24435);
or UO_2380 (O_2380,N_24921,N_18921);
or UO_2381 (O_2381,N_22074,N_22115);
nand UO_2382 (O_2382,N_23171,N_23331);
or UO_2383 (O_2383,N_23668,N_20488);
nand UO_2384 (O_2384,N_22176,N_24760);
or UO_2385 (O_2385,N_22686,N_20099);
nand UO_2386 (O_2386,N_23647,N_22802);
or UO_2387 (O_2387,N_19912,N_24651);
or UO_2388 (O_2388,N_19326,N_19316);
nand UO_2389 (O_2389,N_21969,N_20810);
nand UO_2390 (O_2390,N_24353,N_23191);
nand UO_2391 (O_2391,N_23460,N_24523);
or UO_2392 (O_2392,N_23946,N_24407);
and UO_2393 (O_2393,N_23493,N_23535);
xnor UO_2394 (O_2394,N_22640,N_22243);
and UO_2395 (O_2395,N_20575,N_22487);
and UO_2396 (O_2396,N_21464,N_21093);
nor UO_2397 (O_2397,N_22534,N_19012);
nor UO_2398 (O_2398,N_24599,N_24312);
and UO_2399 (O_2399,N_22459,N_23440);
nor UO_2400 (O_2400,N_23504,N_24516);
nor UO_2401 (O_2401,N_24579,N_24582);
or UO_2402 (O_2402,N_18976,N_19626);
nand UO_2403 (O_2403,N_22876,N_19580);
nand UO_2404 (O_2404,N_22471,N_20775);
nor UO_2405 (O_2405,N_22343,N_22012);
and UO_2406 (O_2406,N_19973,N_21187);
xnor UO_2407 (O_2407,N_20987,N_24701);
and UO_2408 (O_2408,N_20074,N_21834);
and UO_2409 (O_2409,N_24189,N_21460);
or UO_2410 (O_2410,N_23534,N_22084);
or UO_2411 (O_2411,N_20082,N_19671);
or UO_2412 (O_2412,N_19364,N_24263);
and UO_2413 (O_2413,N_18931,N_24913);
nand UO_2414 (O_2414,N_23562,N_19421);
nand UO_2415 (O_2415,N_21039,N_19288);
and UO_2416 (O_2416,N_21077,N_21861);
nand UO_2417 (O_2417,N_24758,N_21224);
nor UO_2418 (O_2418,N_19846,N_19984);
nand UO_2419 (O_2419,N_21099,N_22366);
and UO_2420 (O_2420,N_23346,N_19934);
and UO_2421 (O_2421,N_19249,N_20762);
nand UO_2422 (O_2422,N_24810,N_24036);
and UO_2423 (O_2423,N_22538,N_22155);
nand UO_2424 (O_2424,N_19774,N_19624);
nand UO_2425 (O_2425,N_24553,N_20527);
nand UO_2426 (O_2426,N_23955,N_23079);
or UO_2427 (O_2427,N_23055,N_21919);
xnor UO_2428 (O_2428,N_19590,N_20935);
nand UO_2429 (O_2429,N_20413,N_24540);
nor UO_2430 (O_2430,N_21928,N_22354);
xnor UO_2431 (O_2431,N_23713,N_23899);
and UO_2432 (O_2432,N_24499,N_24309);
and UO_2433 (O_2433,N_24057,N_23118);
xnor UO_2434 (O_2434,N_19030,N_24150);
and UO_2435 (O_2435,N_20254,N_23421);
and UO_2436 (O_2436,N_21892,N_19011);
and UO_2437 (O_2437,N_21680,N_24730);
and UO_2438 (O_2438,N_19080,N_22041);
nand UO_2439 (O_2439,N_20624,N_22009);
or UO_2440 (O_2440,N_20686,N_21277);
and UO_2441 (O_2441,N_22223,N_20090);
or UO_2442 (O_2442,N_21820,N_24844);
nand UO_2443 (O_2443,N_24981,N_24979);
xnor UO_2444 (O_2444,N_22011,N_24151);
nand UO_2445 (O_2445,N_23690,N_20196);
xnor UO_2446 (O_2446,N_24120,N_23465);
nor UO_2447 (O_2447,N_20661,N_19865);
and UO_2448 (O_2448,N_22867,N_24007);
nand UO_2449 (O_2449,N_20917,N_20456);
xor UO_2450 (O_2450,N_19749,N_22969);
nor UO_2451 (O_2451,N_19715,N_20348);
or UO_2452 (O_2452,N_21575,N_23289);
and UO_2453 (O_2453,N_21841,N_20044);
and UO_2454 (O_2454,N_19180,N_21481);
xnor UO_2455 (O_2455,N_20848,N_22698);
or UO_2456 (O_2456,N_22705,N_24215);
nand UO_2457 (O_2457,N_23292,N_21274);
nor UO_2458 (O_2458,N_19677,N_23426);
nand UO_2459 (O_2459,N_22324,N_22355);
nor UO_2460 (O_2460,N_20571,N_22097);
and UO_2461 (O_2461,N_23897,N_23076);
and UO_2462 (O_2462,N_21034,N_18796);
or UO_2463 (O_2463,N_22815,N_22219);
nand UO_2464 (O_2464,N_24795,N_24629);
nor UO_2465 (O_2465,N_24313,N_20653);
xnor UO_2466 (O_2466,N_19578,N_19277);
nor UO_2467 (O_2467,N_22057,N_18901);
and UO_2468 (O_2468,N_19758,N_22231);
or UO_2469 (O_2469,N_19176,N_19829);
and UO_2470 (O_2470,N_22814,N_19868);
xor UO_2471 (O_2471,N_22753,N_19413);
xnor UO_2472 (O_2472,N_21812,N_22493);
and UO_2473 (O_2473,N_24368,N_21535);
and UO_2474 (O_2474,N_20936,N_21917);
and UO_2475 (O_2475,N_23916,N_19430);
and UO_2476 (O_2476,N_20817,N_19045);
nor UO_2477 (O_2477,N_24359,N_23175);
and UO_2478 (O_2478,N_19517,N_23871);
or UO_2479 (O_2479,N_23391,N_20910);
nor UO_2480 (O_2480,N_19775,N_24269);
nand UO_2481 (O_2481,N_24195,N_23276);
nand UO_2482 (O_2482,N_24489,N_18797);
nand UO_2483 (O_2483,N_22531,N_19595);
nand UO_2484 (O_2484,N_18995,N_20184);
nand UO_2485 (O_2485,N_19972,N_22727);
or UO_2486 (O_2486,N_19408,N_21764);
xnor UO_2487 (O_2487,N_22681,N_23195);
nor UO_2488 (O_2488,N_20784,N_21603);
nor UO_2489 (O_2489,N_23469,N_24482);
xor UO_2490 (O_2490,N_21785,N_22817);
xor UO_2491 (O_2491,N_21889,N_20668);
xor UO_2492 (O_2492,N_21781,N_20275);
or UO_2493 (O_2493,N_19572,N_21825);
nor UO_2494 (O_2494,N_23627,N_20617);
xor UO_2495 (O_2495,N_19585,N_21544);
nor UO_2496 (O_2496,N_22445,N_22394);
and UO_2497 (O_2497,N_22248,N_21145);
nand UO_2498 (O_2498,N_20128,N_18842);
and UO_2499 (O_2499,N_19394,N_21604);
nand UO_2500 (O_2500,N_24504,N_24613);
nand UO_2501 (O_2501,N_22374,N_20868);
nand UO_2502 (O_2502,N_20985,N_20696);
nor UO_2503 (O_2503,N_22147,N_24692);
nor UO_2504 (O_2504,N_23324,N_19802);
nand UO_2505 (O_2505,N_20599,N_24059);
nand UO_2506 (O_2506,N_24749,N_23330);
nor UO_2507 (O_2507,N_24961,N_19484);
or UO_2508 (O_2508,N_22879,N_20746);
nand UO_2509 (O_2509,N_22598,N_22104);
nor UO_2510 (O_2510,N_21683,N_24879);
nor UO_2511 (O_2511,N_23210,N_19688);
and UO_2512 (O_2512,N_24104,N_19008);
nand UO_2513 (O_2513,N_23772,N_19359);
or UO_2514 (O_2514,N_22540,N_21617);
xnor UO_2515 (O_2515,N_24010,N_19101);
nand UO_2516 (O_2516,N_19113,N_20136);
and UO_2517 (O_2517,N_19172,N_23500);
xor UO_2518 (O_2518,N_22080,N_23026);
or UO_2519 (O_2519,N_21875,N_20960);
xnor UO_2520 (O_2520,N_22793,N_19136);
nor UO_2521 (O_2521,N_23040,N_22385);
and UO_2522 (O_2522,N_19070,N_19672);
and UO_2523 (O_2523,N_21896,N_20759);
or UO_2524 (O_2524,N_22990,N_18960);
and UO_2525 (O_2525,N_24621,N_23607);
xnor UO_2526 (O_2526,N_21762,N_23722);
or UO_2527 (O_2527,N_23167,N_19418);
xor UO_2528 (O_2528,N_19803,N_24338);
xnor UO_2529 (O_2529,N_19821,N_21236);
xnor UO_2530 (O_2530,N_22252,N_22596);
nor UO_2531 (O_2531,N_19666,N_21191);
nand UO_2532 (O_2532,N_24636,N_20557);
nor UO_2533 (O_2533,N_23419,N_22644);
nand UO_2534 (O_2534,N_21339,N_20220);
or UO_2535 (O_2535,N_20478,N_20999);
xor UO_2536 (O_2536,N_24515,N_19565);
xor UO_2537 (O_2537,N_23930,N_22025);
or UO_2538 (O_2538,N_19881,N_21852);
nor UO_2539 (O_2539,N_23097,N_20892);
nor UO_2540 (O_2540,N_19548,N_20349);
nand UO_2541 (O_2541,N_21772,N_22109);
and UO_2542 (O_2542,N_21909,N_24428);
and UO_2543 (O_2543,N_21788,N_23111);
xnor UO_2544 (O_2544,N_23824,N_19904);
nand UO_2545 (O_2545,N_22809,N_20221);
nor UO_2546 (O_2546,N_19311,N_20720);
xnor UO_2547 (O_2547,N_19219,N_22831);
or UO_2548 (O_2548,N_21477,N_24446);
and UO_2549 (O_2549,N_21784,N_24211);
xnor UO_2550 (O_2550,N_24388,N_24197);
xnor UO_2551 (O_2551,N_23354,N_20374);
nand UO_2552 (O_2552,N_23314,N_23602);
xor UO_2553 (O_2553,N_22172,N_18854);
nor UO_2554 (O_2554,N_21915,N_22921);
xor UO_2555 (O_2555,N_24556,N_23644);
xor UO_2556 (O_2556,N_23963,N_23739);
nor UO_2557 (O_2557,N_20741,N_24792);
nor UO_2558 (O_2558,N_20047,N_23692);
nand UO_2559 (O_2559,N_22660,N_23215);
nand UO_2560 (O_2560,N_23394,N_19975);
or UO_2561 (O_2561,N_21432,N_23531);
or UO_2562 (O_2562,N_23438,N_24409);
xnor UO_2563 (O_2563,N_19302,N_23969);
nor UO_2564 (O_2564,N_20672,N_20112);
xnor UO_2565 (O_2565,N_23024,N_18830);
nor UO_2566 (O_2566,N_19520,N_22416);
or UO_2567 (O_2567,N_21550,N_22411);
nand UO_2568 (O_2568,N_20058,N_22776);
xor UO_2569 (O_2569,N_21082,N_24155);
or UO_2570 (O_2570,N_24957,N_23659);
and UO_2571 (O_2571,N_18969,N_23104);
xor UO_2572 (O_2572,N_20634,N_23656);
and UO_2573 (O_2573,N_23751,N_19914);
and UO_2574 (O_2574,N_21995,N_18757);
and UO_2575 (O_2575,N_20025,N_21011);
nor UO_2576 (O_2576,N_22688,N_21252);
or UO_2577 (O_2577,N_22859,N_24861);
nor UO_2578 (O_2578,N_23343,N_21490);
and UO_2579 (O_2579,N_23282,N_23755);
nor UO_2580 (O_2580,N_24217,N_20799);
nand UO_2581 (O_2581,N_21685,N_20265);
nor UO_2582 (O_2582,N_20659,N_22654);
or UO_2583 (O_2583,N_20125,N_24681);
and UO_2584 (O_2584,N_19966,N_19107);
or UO_2585 (O_2585,N_19741,N_24323);
xor UO_2586 (O_2586,N_22991,N_21101);
nor UO_2587 (O_2587,N_19526,N_21111);
or UO_2588 (O_2588,N_21561,N_20272);
nand UO_2589 (O_2589,N_23041,N_20436);
or UO_2590 (O_2590,N_22425,N_21644);
nor UO_2591 (O_2591,N_19505,N_21183);
nand UO_2592 (O_2592,N_19567,N_19198);
nor UO_2593 (O_2593,N_24035,N_23053);
and UO_2594 (O_2594,N_22677,N_21563);
or UO_2595 (O_2595,N_24301,N_21532);
or UO_2596 (O_2596,N_20147,N_24087);
xor UO_2597 (O_2597,N_19391,N_19734);
nor UO_2598 (O_2598,N_22113,N_22566);
or UO_2599 (O_2599,N_21197,N_22535);
or UO_2600 (O_2600,N_20156,N_21670);
nor UO_2601 (O_2601,N_22552,N_24068);
and UO_2602 (O_2602,N_21941,N_19271);
or UO_2603 (O_2603,N_24076,N_18762);
and UO_2604 (O_2604,N_20406,N_19685);
nand UO_2605 (O_2605,N_21404,N_24253);
nand UO_2606 (O_2606,N_20903,N_19667);
xor UO_2607 (O_2607,N_21618,N_21400);
nand UO_2608 (O_2608,N_20163,N_20327);
or UO_2609 (O_2609,N_21503,N_23135);
xor UO_2610 (O_2610,N_24721,N_24303);
or UO_2611 (O_2611,N_21887,N_23008);
nand UO_2612 (O_2612,N_20119,N_21051);
xor UO_2613 (O_2613,N_21769,N_19964);
nand UO_2614 (O_2614,N_21356,N_24623);
xor UO_2615 (O_2615,N_23184,N_22978);
xnor UO_2616 (O_2616,N_20023,N_23814);
nand UO_2617 (O_2617,N_23559,N_24227);
nor UO_2618 (O_2618,N_19782,N_23066);
or UO_2619 (O_2619,N_24202,N_22830);
nor UO_2620 (O_2620,N_23280,N_20711);
nor UO_2621 (O_2621,N_20861,N_23989);
and UO_2622 (O_2622,N_20780,N_19768);
xor UO_2623 (O_2623,N_24246,N_21023);
and UO_2624 (O_2624,N_22836,N_22718);
nor UO_2625 (O_2625,N_22616,N_22828);
xnor UO_2626 (O_2626,N_20126,N_19897);
nand UO_2627 (O_2627,N_21465,N_23124);
xor UO_2628 (O_2628,N_20197,N_20822);
nand UO_2629 (O_2629,N_23480,N_21060);
nor UO_2630 (O_2630,N_19661,N_21738);
nand UO_2631 (O_2631,N_24557,N_24476);
nand UO_2632 (O_2632,N_20242,N_19911);
nor UO_2633 (O_2633,N_24737,N_19153);
xnor UO_2634 (O_2634,N_23471,N_23864);
xor UO_2635 (O_2635,N_24324,N_24804);
or UO_2636 (O_2636,N_19244,N_22207);
xor UO_2637 (O_2637,N_23745,N_23488);
xor UO_2638 (O_2638,N_23347,N_24280);
or UO_2639 (O_2639,N_24762,N_24481);
xnor UO_2640 (O_2640,N_22994,N_22438);
xnor UO_2641 (O_2641,N_21182,N_21125);
or UO_2642 (O_2642,N_19928,N_22100);
nor UO_2643 (O_2643,N_24382,N_20593);
and UO_2644 (O_2644,N_19965,N_24634);
xor UO_2645 (O_2645,N_23853,N_19371);
nand UO_2646 (O_2646,N_22553,N_19015);
and UO_2647 (O_2647,N_22216,N_24242);
and UO_2648 (O_2648,N_20837,N_20347);
xor UO_2649 (O_2649,N_23192,N_22670);
or UO_2650 (O_2650,N_20805,N_18980);
nand UO_2651 (O_2651,N_20193,N_23064);
xor UO_2652 (O_2652,N_21198,N_23876);
or UO_2653 (O_2653,N_23527,N_20247);
nor UO_2654 (O_2654,N_19781,N_23740);
or UO_2655 (O_2655,N_20939,N_23272);
and UO_2656 (O_2656,N_21166,N_22318);
nor UO_2657 (O_2657,N_24788,N_24631);
nor UO_2658 (O_2658,N_20299,N_24015);
nand UO_2659 (O_2659,N_22310,N_22101);
nor UO_2660 (O_2660,N_24524,N_23834);
nor UO_2661 (O_2661,N_22694,N_20266);
xnor UO_2662 (O_2662,N_22239,N_22299);
xor UO_2663 (O_2663,N_21458,N_20990);
or UO_2664 (O_2664,N_24248,N_23768);
xor UO_2665 (O_2665,N_21353,N_18847);
and UO_2666 (O_2666,N_24789,N_22758);
nand UO_2667 (O_2667,N_21930,N_23348);
xor UO_2668 (O_2668,N_21735,N_23449);
xnor UO_2669 (O_2669,N_21169,N_24406);
nor UO_2670 (O_2670,N_22134,N_24352);
and UO_2671 (O_2671,N_20495,N_24731);
nor UO_2672 (O_2672,N_24744,N_19179);
nor UO_2673 (O_2673,N_21250,N_19958);
nand UO_2674 (O_2674,N_21116,N_19173);
xor UO_2675 (O_2675,N_22703,N_19435);
xnor UO_2676 (O_2676,N_21248,N_19573);
or UO_2677 (O_2677,N_23805,N_20389);
and UO_2678 (O_2678,N_22721,N_22158);
or UO_2679 (O_2679,N_21710,N_23063);
or UO_2680 (O_2680,N_24122,N_21161);
nor UO_2681 (O_2681,N_21467,N_19896);
xor UO_2682 (O_2682,N_22406,N_20238);
nand UO_2683 (O_2683,N_24993,N_20270);
nor UO_2684 (O_2684,N_23249,N_18835);
or UO_2685 (O_2685,N_22292,N_20407);
nand UO_2686 (O_2686,N_22630,N_21551);
nand UO_2687 (O_2687,N_19141,N_19937);
nor UO_2688 (O_2688,N_22258,N_21062);
xor UO_2689 (O_2689,N_18815,N_19743);
and UO_2690 (O_2690,N_19190,N_23189);
and UO_2691 (O_2691,N_23377,N_22092);
nor UO_2692 (O_2692,N_21306,N_23841);
xnor UO_2693 (O_2693,N_21845,N_21354);
and UO_2694 (O_2694,N_20141,N_19691);
nor UO_2695 (O_2695,N_24105,N_23238);
or UO_2696 (O_2696,N_21612,N_20361);
xor UO_2697 (O_2697,N_23351,N_20767);
nor UO_2698 (O_2698,N_23798,N_20750);
nand UO_2699 (O_2699,N_21973,N_23109);
nor UO_2700 (O_2700,N_20856,N_24560);
xnor UO_2701 (O_2701,N_18990,N_19058);
xnor UO_2702 (O_2702,N_22465,N_21399);
and UO_2703 (O_2703,N_20560,N_20757);
or UO_2704 (O_2704,N_24286,N_22417);
nand UO_2705 (O_2705,N_24043,N_19237);
nand UO_2706 (O_2706,N_21488,N_23638);
nor UO_2707 (O_2707,N_21783,N_22367);
nand UO_2708 (O_2708,N_20095,N_22249);
nand UO_2709 (O_2709,N_19555,N_23771);
nand UO_2710 (O_2710,N_22861,N_24262);
xnor UO_2711 (O_2711,N_24648,N_20612);
and UO_2712 (O_2712,N_21773,N_22275);
and UO_2713 (O_2713,N_19094,N_19279);
nor UO_2714 (O_2714,N_22460,N_23512);
and UO_2715 (O_2715,N_20021,N_19356);
and UO_2716 (O_2716,N_19592,N_24673);
nor UO_2717 (O_2717,N_22541,N_19298);
and UO_2718 (O_2718,N_19057,N_22371);
and UO_2719 (O_2719,N_24682,N_22235);
or UO_2720 (O_2720,N_24653,N_21950);
or UO_2721 (O_2721,N_24108,N_20441);
xnor UO_2722 (O_2722,N_24161,N_20896);
xor UO_2723 (O_2723,N_23011,N_23840);
nor UO_2724 (O_2724,N_23179,N_19824);
nor UO_2725 (O_2725,N_22982,N_22655);
nand UO_2726 (O_2726,N_21970,N_21276);
and UO_2727 (O_2727,N_20916,N_20698);
or UO_2728 (O_2728,N_21421,N_23757);
or UO_2729 (O_2729,N_22578,N_24251);
or UO_2730 (O_2730,N_18946,N_19633);
and UO_2731 (O_2731,N_20370,N_19697);
nand UO_2732 (O_2732,N_20121,N_19059);
or UO_2733 (O_2733,N_22715,N_21717);
nand UO_2734 (O_2734,N_19327,N_21124);
or UO_2735 (O_2735,N_23570,N_19297);
nand UO_2736 (O_2736,N_20426,N_24032);
xnor UO_2737 (O_2737,N_21018,N_21633);
or UO_2738 (O_2738,N_22951,N_22794);
and UO_2739 (O_2739,N_20769,N_21207);
and UO_2740 (O_2740,N_21119,N_19197);
and UO_2741 (O_2741,N_24699,N_21813);
xor UO_2742 (O_2742,N_18855,N_22667);
nand UO_2743 (O_2743,N_21818,N_19657);
nor UO_2744 (O_2744,N_20182,N_21212);
xnor UO_2745 (O_2745,N_19778,N_24336);
nor UO_2746 (O_2746,N_24926,N_24381);
xor UO_2747 (O_2747,N_24934,N_20705);
xor UO_2748 (O_2748,N_19921,N_22954);
or UO_2749 (O_2749,N_22819,N_19748);
and UO_2750 (O_2750,N_24590,N_21991);
and UO_2751 (O_2751,N_23459,N_22761);
or UO_2752 (O_2752,N_20401,N_21519);
and UO_2753 (O_2753,N_23165,N_20756);
xnor UO_2754 (O_2754,N_23016,N_21459);
or UO_2755 (O_2755,N_20977,N_19485);
and UO_2756 (O_2756,N_22947,N_21796);
and UO_2757 (O_2757,N_22940,N_23844);
xnor UO_2758 (O_2758,N_24938,N_20102);
nand UO_2759 (O_2759,N_23919,N_19957);
nor UO_2760 (O_2760,N_23446,N_24213);
or UO_2761 (O_2761,N_20549,N_19503);
and UO_2762 (O_2762,N_21005,N_23326);
or UO_2763 (O_2763,N_18900,N_21805);
nor UO_2764 (O_2764,N_23233,N_24894);
and UO_2765 (O_2765,N_22093,N_20367);
nor UO_2766 (O_2766,N_19274,N_23898);
and UO_2767 (O_2767,N_23362,N_23406);
nand UO_2768 (O_2768,N_22895,N_23025);
and UO_2769 (O_2769,N_23255,N_19427);
nand UO_2770 (O_2770,N_23787,N_19160);
xor UO_2771 (O_2771,N_24716,N_24149);
xor UO_2772 (O_2772,N_22161,N_22657);
and UO_2773 (O_2773,N_22854,N_22437);
or UO_2774 (O_2774,N_19420,N_23376);
xnor UO_2775 (O_2775,N_21502,N_21015);
and UO_2776 (O_2776,N_22461,N_24962);
or UO_2777 (O_2777,N_21677,N_24568);
nand UO_2778 (O_2778,N_24530,N_20157);
xnor UO_2779 (O_2779,N_24920,N_20287);
or UO_2780 (O_2780,N_23533,N_20595);
nor UO_2781 (O_2781,N_19405,N_18834);
xor UO_2782 (O_2782,N_19481,N_19841);
and UO_2783 (O_2783,N_19859,N_22319);
or UO_2784 (O_2784,N_18962,N_22194);
nor UO_2785 (O_2785,N_23226,N_22457);
nor UO_2786 (O_2786,N_24850,N_19523);
or UO_2787 (O_2787,N_21146,N_22441);
and UO_2788 (O_2788,N_22148,N_23581);
or UO_2789 (O_2789,N_24240,N_20444);
nand UO_2790 (O_2790,N_23034,N_20545);
nand UO_2791 (O_2791,N_18922,N_19602);
nand UO_2792 (O_2792,N_21439,N_23780);
nor UO_2793 (O_2793,N_18848,N_23650);
nor UO_2794 (O_2794,N_23911,N_23800);
nand UO_2795 (O_2795,N_24867,N_24463);
xor UO_2796 (O_2796,N_22622,N_18994);
and UO_2797 (O_2797,N_24546,N_21679);
nor UO_2798 (O_2798,N_19540,N_20828);
nor UO_2799 (O_2799,N_23601,N_23483);
and UO_2800 (O_2800,N_19857,N_21746);
and UO_2801 (O_2801,N_22476,N_22021);
xnor UO_2802 (O_2802,N_23228,N_24345);
nand UO_2803 (O_2803,N_21048,N_23961);
xnor UO_2804 (O_2804,N_23448,N_20731);
nand UO_2805 (O_2805,N_21242,N_21968);
or UO_2806 (O_2806,N_23776,N_19024);
and UO_2807 (O_2807,N_21955,N_18780);
nor UO_2808 (O_2808,N_24470,N_23270);
xor UO_2809 (O_2809,N_23860,N_21238);
xnor UO_2810 (O_2810,N_22557,N_23514);
xor UO_2811 (O_2811,N_23381,N_21586);
xnor UO_2812 (O_2812,N_23158,N_19687);
nor UO_2813 (O_2813,N_24049,N_20614);
nand UO_2814 (O_2814,N_23557,N_24565);
or UO_2815 (O_2815,N_22251,N_23833);
nor UO_2816 (O_2816,N_19612,N_21471);
nor UO_2817 (O_2817,N_22678,N_18816);
or UO_2818 (O_2818,N_19360,N_24305);
or UO_2819 (O_2819,N_21386,N_21719);
xor UO_2820 (O_2820,N_24459,N_21611);
nor UO_2821 (O_2821,N_19805,N_19109);
and UO_2822 (O_2822,N_18944,N_19300);
nand UO_2823 (O_2823,N_19918,N_24400);
nand UO_2824 (O_2824,N_22033,N_24444);
and UO_2825 (O_2825,N_20089,N_20305);
xnor UO_2826 (O_2826,N_20395,N_19884);
or UO_2827 (O_2827,N_19588,N_18982);
or UO_2828 (O_2828,N_19561,N_19126);
and UO_2829 (O_2829,N_21880,N_23201);
xnor UO_2830 (O_2830,N_18963,N_21210);
nor UO_2831 (O_2831,N_22868,N_20521);
xor UO_2832 (O_2832,N_19187,N_19425);
nand UO_2833 (O_2833,N_22289,N_24097);
nand UO_2834 (O_2834,N_21428,N_22684);
and UO_2835 (O_2835,N_23984,N_19066);
or UO_2836 (O_2836,N_19947,N_23411);
nand UO_2837 (O_2837,N_21287,N_23423);
xor UO_2838 (O_2838,N_22714,N_22510);
nand UO_2839 (O_2839,N_24008,N_21590);
xnor UO_2840 (O_2840,N_19910,N_23530);
and UO_2841 (O_2841,N_22587,N_20218);
and UO_2842 (O_2842,N_23788,N_19170);
xor UO_2843 (O_2843,N_19673,N_24138);
and UO_2844 (O_2844,N_21850,N_19328);
xor UO_2845 (O_2845,N_23703,N_20455);
nand UO_2846 (O_2846,N_24887,N_21555);
and UO_2847 (O_2847,N_21171,N_23665);
nand UO_2848 (O_2848,N_20006,N_19600);
or UO_2849 (O_2849,N_24943,N_19040);
and UO_2850 (O_2850,N_20449,N_19665);
nand UO_2851 (O_2851,N_23156,N_20845);
nor UO_2852 (O_2852,N_23134,N_21959);
and UO_2853 (O_2853,N_24279,N_20122);
nor UO_2854 (O_2854,N_23054,N_21090);
nor UO_2855 (O_2855,N_24366,N_21009);
nor UO_2856 (O_2856,N_22722,N_22164);
nor UO_2857 (O_2857,N_24107,N_20908);
and UO_2858 (O_2858,N_22575,N_24686);
and UO_2859 (O_2859,N_21097,N_23882);
xnor UO_2860 (O_2860,N_21324,N_22570);
or UO_2861 (O_2861,N_24295,N_23716);
xor UO_2862 (O_2862,N_21553,N_21067);
xnor UO_2863 (O_2863,N_21196,N_24905);
xor UO_2864 (O_2864,N_20017,N_23096);
nand UO_2865 (O_2865,N_22049,N_21482);
and UO_2866 (O_2866,N_22909,N_21085);
or UO_2867 (O_2867,N_21895,N_20497);
nor UO_2868 (O_2868,N_24856,N_20470);
or UO_2869 (O_2869,N_19234,N_19875);
xnor UO_2870 (O_2870,N_22708,N_20423);
and UO_2871 (O_2871,N_24642,N_24928);
and UO_2872 (O_2872,N_22910,N_22525);
nand UO_2873 (O_2873,N_24845,N_22750);
xor UO_2874 (O_2874,N_24414,N_22020);
xnor UO_2875 (O_2875,N_20915,N_24528);
or UO_2876 (O_2876,N_23174,N_23721);
xor UO_2877 (O_2877,N_22562,N_23170);
or UO_2878 (O_2878,N_24728,N_20307);
xor UO_2879 (O_2879,N_23147,N_23680);
nand UO_2880 (O_2880,N_22316,N_20529);
nor UO_2881 (O_2881,N_19893,N_18920);
nand UO_2882 (O_2882,N_24408,N_21533);
nor UO_2883 (O_2883,N_20320,N_20849);
or UO_2884 (O_2884,N_20056,N_20137);
nand UO_2885 (O_2885,N_24882,N_23217);
and UO_2886 (O_2886,N_19260,N_22202);
xnor UO_2887 (O_2887,N_19541,N_24536);
xnor UO_2888 (O_2888,N_21108,N_23271);
nor UO_2889 (O_2889,N_22611,N_19366);
nand UO_2890 (O_2890,N_21308,N_19025);
or UO_2891 (O_2891,N_21899,N_22702);
nand UO_2892 (O_2892,N_24541,N_22523);
xnor UO_2893 (O_2893,N_19389,N_24052);
xnor UO_2894 (O_2894,N_19808,N_21565);
or UO_2895 (O_2895,N_21770,N_19065);
nor UO_2896 (O_2896,N_19393,N_22742);
or UO_2897 (O_2897,N_21041,N_24337);
or UO_2898 (O_2898,N_20208,N_22948);
xor UO_2899 (O_2899,N_22896,N_24283);
nand UO_2900 (O_2900,N_21885,N_22368);
nor UO_2901 (O_2901,N_19851,N_20261);
nor UO_2902 (O_2902,N_23498,N_24361);
and UO_2903 (O_2903,N_21534,N_19641);
nand UO_2904 (O_2904,N_23453,N_23142);
nand UO_2905 (O_2905,N_18882,N_19535);
nand UO_2906 (O_2906,N_22263,N_19594);
or UO_2907 (O_2907,N_19210,N_23021);
nor UO_2908 (O_2908,N_24316,N_21115);
or UO_2909 (O_2909,N_19892,N_19373);
nor UO_2910 (O_2910,N_20304,N_23242);
or UO_2911 (O_2911,N_23933,N_18876);
or UO_2912 (O_2912,N_23186,N_19152);
nor UO_2913 (O_2913,N_21322,N_23309);
nor UO_2914 (O_2914,N_24973,N_23702);
and UO_2915 (O_2915,N_20565,N_18954);
or UO_2916 (O_2916,N_24364,N_21902);
nand UO_2917 (O_2917,N_24975,N_20793);
nand UO_2918 (O_2918,N_21068,N_19184);
and UO_2919 (O_2919,N_24828,N_21650);
xor UO_2920 (O_2920,N_20811,N_19091);
nand UO_2921 (O_2921,N_24350,N_21430);
nand UO_2922 (O_2922,N_23214,N_22087);
xor UO_2923 (O_2923,N_24585,N_21160);
nand UO_2924 (O_2924,N_22335,N_24450);
nand UO_2925 (O_2925,N_20481,N_22455);
nor UO_2926 (O_2926,N_21581,N_20026);
xnor UO_2927 (O_2927,N_22796,N_21934);
and UO_2928 (O_2928,N_20737,N_23604);
nor UO_2929 (O_2929,N_20965,N_23524);
xnor UO_2930 (O_2930,N_21786,N_23501);
nand UO_2931 (O_2931,N_22907,N_20743);
xor UO_2932 (O_2932,N_19755,N_22255);
xnor UO_2933 (O_2933,N_24363,N_20530);
nand UO_2934 (O_2934,N_21167,N_21156);
xnor UO_2935 (O_2935,N_23904,N_18777);
or UO_2936 (O_2936,N_23307,N_18986);
or UO_2937 (O_2937,N_20230,N_21100);
nand UO_2938 (O_2938,N_23038,N_19133);
nor UO_2939 (O_2939,N_19229,N_19088);
nand UO_2940 (O_2940,N_20015,N_22743);
and UO_2941 (O_2941,N_19610,N_21270);
and UO_2942 (O_2942,N_18940,N_21185);
nand UO_2943 (O_2943,N_20792,N_23222);
nor UO_2944 (O_2944,N_20164,N_22801);
xnor UO_2945 (O_2945,N_23786,N_20976);
or UO_2946 (O_2946,N_23315,N_20801);
xor UO_2947 (O_2947,N_24136,N_20046);
xor UO_2948 (O_2948,N_24233,N_19771);
xnor UO_2949 (O_2949,N_18958,N_22058);
nor UO_2950 (O_2950,N_24124,N_24592);
xor UO_2951 (O_2951,N_20065,N_19930);
nor UO_2952 (O_2952,N_19495,N_23048);
xnor UO_2953 (O_2953,N_21463,N_21870);
nand UO_2954 (O_2954,N_20887,N_20048);
or UO_2955 (O_2955,N_20501,N_22699);
nor UO_2956 (O_2956,N_21297,N_22400);
nor UO_2957 (O_2957,N_23691,N_21882);
and UO_2958 (O_2958,N_22222,N_24500);
nor UO_2959 (O_2959,N_24853,N_19006);
nor UO_2960 (O_2960,N_23344,N_19844);
or UO_2961 (O_2961,N_22884,N_23323);
xnor UO_2962 (O_2962,N_20219,N_23088);
nand UO_2963 (O_2963,N_21434,N_20689);
xnor UO_2964 (O_2964,N_19099,N_18890);
or UO_2965 (O_2965,N_21521,N_19329);
nand UO_2966 (O_2966,N_22870,N_19562);
nand UO_2967 (O_2967,N_19323,N_24434);
nor UO_2968 (O_2968,N_23763,N_22638);
nand UO_2969 (O_2969,N_20790,N_23615);
nand UO_2970 (O_2970,N_21926,N_21112);
and UO_2971 (O_2971,N_23318,N_22348);
xnor UO_2972 (O_2972,N_22894,N_19292);
xor UO_2973 (O_2973,N_24456,N_24602);
nor UO_2974 (O_2974,N_22897,N_21325);
or UO_2975 (O_2975,N_24813,N_21393);
xnor UO_2976 (O_2976,N_23746,N_24419);
and UO_2977 (O_2977,N_22390,N_20142);
and UO_2978 (O_2978,N_23367,N_20927);
xor UO_2979 (O_2979,N_20152,N_19482);
or UO_2980 (O_2980,N_24606,N_24252);
or UO_2981 (O_2981,N_19447,N_22143);
xnor UO_2982 (O_2982,N_21753,N_20228);
or UO_2983 (O_2983,N_20342,N_19431);
nand UO_2984 (O_2984,N_23168,N_20028);
nor UO_2985 (O_2985,N_19500,N_21070);
or UO_2986 (O_2986,N_24823,N_22449);
nand UO_2987 (O_2987,N_22314,N_20013);
and UO_2988 (O_2988,N_21176,N_18886);
and UO_2989 (O_2989,N_19981,N_19967);
or UO_2990 (O_2990,N_23957,N_21602);
and UO_2991 (O_2991,N_23281,N_23711);
or UO_2992 (O_2992,N_19043,N_23606);
or UO_2993 (O_2993,N_24914,N_24787);
nand UO_2994 (O_2994,N_22280,N_20931);
or UO_2995 (O_2995,N_22031,N_22766);
or UO_2996 (O_2996,N_21148,N_20899);
nand UO_2997 (O_2997,N_21416,N_21668);
and UO_2998 (O_2998,N_20386,N_21372);
xnor UO_2999 (O_2999,N_24377,N_20989);
endmodule