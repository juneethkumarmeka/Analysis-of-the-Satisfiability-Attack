module basic_1500_15000_2000_10_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_78,In_122);
xor U1 (N_1,In_1108,In_896);
nor U2 (N_2,In_1342,In_377);
or U3 (N_3,In_554,In_1404);
nor U4 (N_4,In_713,In_1492);
or U5 (N_5,In_340,In_822);
or U6 (N_6,In_1271,In_1105);
nand U7 (N_7,In_1018,In_685);
or U8 (N_8,In_1038,In_1229);
nor U9 (N_9,In_150,In_166);
nand U10 (N_10,In_625,In_1071);
and U11 (N_11,In_101,In_755);
and U12 (N_12,In_341,In_427);
and U13 (N_13,In_407,In_1310);
and U14 (N_14,In_1383,In_1489);
or U15 (N_15,In_485,In_1259);
and U16 (N_16,In_663,In_1056);
nand U17 (N_17,In_1099,In_947);
nand U18 (N_18,In_1266,In_84);
nand U19 (N_19,In_849,In_571);
and U20 (N_20,In_786,In_677);
nor U21 (N_21,In_1374,In_59);
nor U22 (N_22,In_1043,In_610);
nor U23 (N_23,In_293,In_1185);
nor U24 (N_24,In_739,In_1488);
or U25 (N_25,In_172,In_98);
nand U26 (N_26,In_1371,In_1390);
nor U27 (N_27,In_632,In_1093);
nor U28 (N_28,In_1382,In_66);
and U29 (N_29,In_388,In_1397);
nand U30 (N_30,In_288,In_906);
or U31 (N_31,In_575,In_477);
and U32 (N_32,In_420,In_451);
xor U33 (N_33,In_1336,In_164);
or U34 (N_34,In_593,In_1021);
xor U35 (N_35,In_842,In_363);
and U36 (N_36,In_1211,In_301);
and U37 (N_37,In_633,In_576);
or U38 (N_38,In_463,In_144);
and U39 (N_39,In_133,In_179);
or U40 (N_40,In_985,In_1347);
nor U41 (N_41,In_740,In_1244);
and U42 (N_42,In_467,In_320);
nor U43 (N_43,In_80,In_1332);
nor U44 (N_44,In_1328,In_81);
and U45 (N_45,In_1017,In_989);
or U46 (N_46,In_729,In_1373);
nand U47 (N_47,In_1364,In_520);
or U48 (N_48,In_20,In_603);
nor U49 (N_49,In_843,In_1308);
and U50 (N_50,In_319,In_531);
or U51 (N_51,In_1098,In_631);
and U52 (N_52,In_519,In_234);
or U53 (N_53,In_1034,In_55);
nand U54 (N_54,In_549,In_1317);
nor U55 (N_55,In_1475,In_154);
nand U56 (N_56,In_1073,In_1370);
nand U57 (N_57,In_656,In_1321);
and U58 (N_58,In_850,In_698);
nand U59 (N_59,In_371,In_717);
nand U60 (N_60,In_572,In_4);
or U61 (N_61,In_830,In_801);
nand U62 (N_62,In_362,In_1050);
nor U63 (N_63,In_27,In_917);
nand U64 (N_64,In_408,In_403);
or U65 (N_65,In_457,In_646);
nand U66 (N_66,In_500,In_967);
nor U67 (N_67,In_969,In_148);
nand U68 (N_68,In_1316,In_758);
and U69 (N_69,In_282,In_74);
xnor U70 (N_70,In_1025,In_1035);
nand U71 (N_71,In_957,In_1394);
and U72 (N_72,In_1412,In_1353);
nor U73 (N_73,In_1134,In_1222);
xnor U74 (N_74,In_903,In_796);
nand U75 (N_75,In_670,In_644);
or U76 (N_76,In_1172,In_1441);
nor U77 (N_77,In_1274,In_980);
and U78 (N_78,In_870,In_60);
nor U79 (N_79,In_863,In_955);
and U80 (N_80,In_691,In_752);
nor U81 (N_81,In_1204,In_1241);
or U82 (N_82,In_1365,In_475);
nand U83 (N_83,In_323,In_1423);
nand U84 (N_84,In_1341,In_1294);
and U85 (N_85,In_276,In_1337);
and U86 (N_86,In_318,In_1232);
and U87 (N_87,In_1398,In_415);
and U88 (N_88,In_834,In_744);
or U89 (N_89,In_1486,In_515);
and U90 (N_90,In_11,In_426);
and U91 (N_91,In_538,In_33);
or U92 (N_92,In_902,In_1000);
and U93 (N_93,In_298,In_1131);
nor U94 (N_94,In_687,In_558);
or U95 (N_95,In_1401,In_961);
and U96 (N_96,In_52,In_1260);
xnor U97 (N_97,In_839,In_1490);
nor U98 (N_98,In_1453,In_1142);
xnor U99 (N_99,In_1302,In_569);
nand U100 (N_100,In_750,In_1235);
and U101 (N_101,In_361,In_1225);
or U102 (N_102,In_99,In_794);
or U103 (N_103,In_1262,In_1165);
or U104 (N_104,In_1206,In_88);
or U105 (N_105,In_1305,In_806);
nand U106 (N_106,In_846,In_1377);
nor U107 (N_107,In_1372,In_85);
nor U108 (N_108,In_394,In_452);
nor U109 (N_109,In_704,In_913);
and U110 (N_110,In_329,In_1496);
or U111 (N_111,In_1419,In_991);
nand U112 (N_112,In_769,In_127);
and U113 (N_113,In_1233,In_285);
and U114 (N_114,In_1261,In_277);
nand U115 (N_115,In_437,In_1173);
xor U116 (N_116,In_608,In_1003);
and U117 (N_117,In_997,In_322);
or U118 (N_118,In_1022,In_959);
or U119 (N_119,In_1216,In_220);
and U120 (N_120,In_354,In_1436);
xnor U121 (N_121,In_1163,In_266);
xnor U122 (N_122,In_208,In_1209);
or U123 (N_123,In_871,In_481);
or U124 (N_124,In_1445,In_389);
nor U125 (N_125,In_130,In_1298);
or U126 (N_126,In_391,In_881);
nand U127 (N_127,In_159,In_49);
and U128 (N_128,In_552,In_775);
nand U129 (N_129,In_129,In_584);
or U130 (N_130,In_296,In_1471);
nand U131 (N_131,In_792,In_286);
nand U132 (N_132,In_1236,In_737);
or U133 (N_133,In_165,In_516);
nand U134 (N_134,In_197,In_507);
nand U135 (N_135,In_1491,In_594);
nor U136 (N_136,In_675,In_1053);
or U137 (N_137,In_879,In_171);
xnor U138 (N_138,In_347,In_667);
and U139 (N_139,In_652,In_890);
xnor U140 (N_140,In_1177,In_158);
nor U141 (N_141,In_905,In_766);
xnor U142 (N_142,In_1121,In_1118);
nand U143 (N_143,In_506,In_1051);
nor U144 (N_144,In_1167,In_615);
or U145 (N_145,In_604,In_1077);
nor U146 (N_146,In_77,In_1095);
or U147 (N_147,In_264,In_1117);
or U148 (N_148,In_1484,In_18);
nor U149 (N_149,In_69,In_272);
nor U150 (N_150,In_970,In_707);
or U151 (N_151,In_1013,In_909);
xor U152 (N_152,In_1387,In_385);
and U153 (N_153,In_920,In_1092);
nor U154 (N_154,In_599,In_180);
or U155 (N_155,In_1460,In_173);
nor U156 (N_156,In_421,In_1433);
or U157 (N_157,In_819,In_458);
and U158 (N_158,In_824,In_1499);
xnor U159 (N_159,In_1350,In_901);
nand U160 (N_160,In_797,In_735);
and U161 (N_161,In_848,In_1447);
or U162 (N_162,In_1313,In_702);
or U163 (N_163,In_629,In_1146);
and U164 (N_164,In_254,In_372);
or U165 (N_165,In_390,In_46);
or U166 (N_166,In_1381,In_86);
or U167 (N_167,In_351,In_1089);
or U168 (N_168,In_944,In_462);
or U169 (N_169,In_683,In_1415);
or U170 (N_170,In_1465,In_606);
nand U171 (N_171,In_13,In_732);
or U172 (N_172,In_1187,In_492);
or U173 (N_173,In_338,In_1155);
nor U174 (N_174,In_812,In_1180);
and U175 (N_175,In_1307,In_756);
nor U176 (N_176,In_627,In_1088);
and U177 (N_177,In_104,In_776);
or U178 (N_178,In_994,In_126);
and U179 (N_179,In_641,In_513);
nand U180 (N_180,In_1368,In_1032);
or U181 (N_181,In_268,In_512);
nor U182 (N_182,In_308,In_253);
nand U183 (N_183,In_1468,In_249);
nor U184 (N_184,In_125,In_423);
and U185 (N_185,In_79,In_337);
nor U186 (N_186,In_899,In_754);
or U187 (N_187,In_1223,In_940);
xor U188 (N_188,In_470,In_1144);
and U189 (N_189,In_1124,In_1422);
and U190 (N_190,In_30,In_676);
and U191 (N_191,In_202,In_517);
and U192 (N_192,In_218,In_1255);
nor U193 (N_193,In_1091,In_161);
or U194 (N_194,In_1132,In_194);
nand U195 (N_195,In_1215,In_1231);
and U196 (N_196,In_724,In_482);
and U197 (N_197,In_726,In_696);
nand U198 (N_198,In_541,In_1399);
and U199 (N_199,In_473,In_487);
nor U200 (N_200,In_406,In_216);
nand U201 (N_201,In_356,In_1199);
and U202 (N_202,In_145,In_1202);
nand U203 (N_203,In_1060,In_260);
xor U204 (N_204,In_1076,In_954);
or U205 (N_205,In_605,In_1312);
or U206 (N_206,In_1213,In_914);
or U207 (N_207,In_1319,In_278);
nor U208 (N_208,In_1362,In_859);
and U209 (N_209,In_1301,In_1147);
nand U210 (N_210,In_853,In_722);
or U211 (N_211,In_450,In_201);
nand U212 (N_212,In_1116,In_1041);
xor U213 (N_213,In_416,In_39);
xor U214 (N_214,In_175,In_804);
nor U215 (N_215,In_1192,In_353);
xnor U216 (N_216,In_1281,In_1046);
xor U217 (N_217,In_1174,In_1400);
and U218 (N_218,In_841,In_837);
nand U219 (N_219,In_1031,In_418);
or U220 (N_220,In_1435,In_828);
or U221 (N_221,In_461,In_771);
nand U222 (N_222,In_731,In_818);
nor U223 (N_223,In_92,In_1424);
or U224 (N_224,In_73,In_1380);
and U225 (N_225,In_1268,In_851);
or U226 (N_226,In_706,In_336);
xor U227 (N_227,In_1348,In_1094);
nor U228 (N_228,In_762,In_67);
and U229 (N_229,In_586,In_9);
or U230 (N_230,In_432,In_366);
nand U231 (N_231,In_188,In_833);
nor U232 (N_232,In_118,In_2);
nor U233 (N_233,In_258,In_561);
nor U234 (N_234,In_128,In_207);
nand U235 (N_235,In_952,In_497);
nor U236 (N_236,In_1285,In_190);
nor U237 (N_237,In_24,In_813);
xor U238 (N_238,In_357,In_883);
nor U239 (N_239,In_1361,In_121);
nor U240 (N_240,In_456,In_1254);
nor U241 (N_241,In_559,In_343);
and U242 (N_242,In_236,In_267);
nor U243 (N_243,In_768,In_435);
nor U244 (N_244,In_1396,In_365);
and U245 (N_245,In_680,In_1195);
nand U246 (N_246,In_623,In_5);
or U247 (N_247,In_205,In_177);
or U248 (N_248,In_412,In_1123);
or U249 (N_249,In_1277,In_1487);
nand U250 (N_250,In_928,In_537);
and U251 (N_251,In_1210,In_619);
or U252 (N_252,In_1482,In_54);
nand U253 (N_253,In_251,In_484);
nor U254 (N_254,In_304,In_1090);
and U255 (N_255,In_352,In_369);
nor U256 (N_256,In_783,In_1459);
nor U257 (N_257,In_607,In_898);
xnor U258 (N_258,In_1275,In_132);
and U259 (N_259,In_810,In_654);
and U260 (N_260,In_476,In_1284);
xnor U261 (N_261,In_772,In_678);
nor U262 (N_262,In_324,In_934);
nor U263 (N_263,In_1110,In_163);
nand U264 (N_264,In_431,In_359);
or U265 (N_265,In_1085,In_397);
and U266 (N_266,In_892,In_156);
and U267 (N_267,In_413,In_72);
and U268 (N_268,In_314,In_109);
nor U269 (N_269,In_686,In_1066);
or U270 (N_270,In_1219,In_139);
or U271 (N_271,In_243,In_1061);
xnor U272 (N_272,In_1251,In_743);
and U273 (N_273,In_616,In_660);
xnor U274 (N_274,In_47,In_1005);
nor U275 (N_275,In_1367,In_921);
and U276 (N_276,In_630,In_1303);
and U277 (N_277,In_1161,In_1087);
or U278 (N_278,In_1019,In_1080);
nand U279 (N_279,In_521,In_113);
xnor U280 (N_280,In_233,In_581);
or U281 (N_281,In_455,In_1265);
xnor U282 (N_282,In_727,In_310);
and U283 (N_283,In_560,In_1104);
nor U284 (N_284,In_595,In_1291);
nand U285 (N_285,In_788,In_1193);
nand U286 (N_286,In_1253,In_543);
nand U287 (N_287,In_930,In_488);
nand U288 (N_288,In_1340,In_893);
nor U289 (N_289,In_326,In_1137);
and U290 (N_290,In_332,In_142);
nor U291 (N_291,In_45,In_291);
or U292 (N_292,In_1280,In_742);
and U293 (N_293,In_1024,In_378);
nor U294 (N_294,In_1333,In_998);
and U295 (N_295,In_1318,In_247);
or U296 (N_296,In_1205,In_1249);
nor U297 (N_297,In_741,In_1326);
nor U298 (N_298,In_760,In_651);
nand U299 (N_299,In_1227,In_618);
or U300 (N_300,In_7,In_137);
and U301 (N_301,In_1448,In_811);
nor U302 (N_302,In_831,In_454);
nand U303 (N_303,In_719,In_429);
and U304 (N_304,In_669,In_219);
or U305 (N_305,In_1048,In_1068);
and U306 (N_306,In_1217,In_1191);
nand U307 (N_307,In_414,In_907);
and U308 (N_308,In_425,In_916);
or U309 (N_309,In_1114,In_376);
xor U310 (N_310,In_975,In_335);
nor U311 (N_311,In_1036,In_405);
nand U312 (N_312,In_1242,In_131);
and U313 (N_313,In_478,In_635);
and U314 (N_314,In_986,In_662);
or U315 (N_315,In_17,In_638);
nor U316 (N_316,In_770,In_505);
and U317 (N_317,In_620,In_1355);
or U318 (N_318,In_299,In_1343);
nand U319 (N_319,In_82,In_87);
nand U320 (N_320,In_1464,In_8);
or U321 (N_321,In_590,In_189);
and U322 (N_322,In_1411,In_1074);
nor U323 (N_323,In_915,In_200);
or U324 (N_324,In_439,In_275);
nand U325 (N_325,In_518,In_1228);
xnor U326 (N_326,In_246,In_1410);
nand U327 (N_327,In_1430,In_1052);
and U328 (N_328,In_370,In_259);
and U329 (N_329,In_826,In_628);
and U330 (N_330,In_1140,In_53);
nor U331 (N_331,In_241,In_1200);
or U332 (N_332,In_57,In_1029);
nand U333 (N_333,In_682,In_483);
and U334 (N_334,In_995,In_1290);
nand U335 (N_335,In_401,In_1357);
and U336 (N_336,In_230,In_910);
and U337 (N_337,In_1111,In_1197);
or U338 (N_338,In_589,In_637);
or U339 (N_339,In_1010,In_551);
nor U340 (N_340,In_26,In_874);
and U341 (N_341,In_965,In_1378);
or U342 (N_342,In_624,In_501);
or U343 (N_343,In_261,In_1349);
or U344 (N_344,In_1276,In_578);
nand U345 (N_345,In_221,In_872);
and U346 (N_346,In_274,In_545);
nand U347 (N_347,In_1449,In_938);
and U348 (N_348,In_582,In_300);
or U349 (N_349,In_281,In_976);
nor U350 (N_350,In_1292,In_1469);
xor U351 (N_351,In_474,In_529);
or U352 (N_352,In_239,In_417);
nand U353 (N_353,In_950,In_346);
and U354 (N_354,In_393,In_1102);
and U355 (N_355,In_865,In_399);
nor U356 (N_356,In_35,In_438);
nand U357 (N_357,In_773,In_527);
nor U358 (N_358,In_658,In_953);
and U359 (N_359,In_1327,In_212);
nor U360 (N_360,In_184,In_613);
and U361 (N_361,In_41,In_511);
or U362 (N_362,In_927,In_321);
nor U363 (N_363,In_522,In_809);
nand U364 (N_364,In_1175,In_1008);
and U365 (N_365,In_925,In_494);
and U366 (N_366,In_867,In_1156);
or U367 (N_367,In_912,In_655);
nand U368 (N_368,In_1126,In_964);
nand U369 (N_369,In_866,In_1282);
xnor U370 (N_370,In_671,In_1462);
nor U371 (N_371,In_96,In_1369);
nor U372 (N_372,In_147,In_718);
nor U373 (N_373,In_1039,In_238);
nor U374 (N_374,In_857,In_793);
or U375 (N_375,In_224,In_1478);
xnor U376 (N_376,In_1078,In_248);
nor U377 (N_377,In_926,In_140);
or U378 (N_378,In_1176,In_1356);
and U379 (N_379,In_922,In_21);
nand U380 (N_380,In_697,In_56);
nand U381 (N_381,In_1446,In_779);
nand U382 (N_382,In_1030,In_700);
xor U383 (N_383,In_273,In_1403);
nor U384 (N_384,In_703,In_1086);
and U385 (N_385,In_860,In_222);
or U386 (N_386,In_192,In_753);
or U387 (N_387,In_315,In_1477);
or U388 (N_388,In_1256,In_245);
nor U389 (N_389,In_1346,In_1162);
or U390 (N_390,In_384,In_1179);
nand U391 (N_391,In_526,In_751);
and U392 (N_392,In_213,In_579);
nor U393 (N_393,In_1442,In_1335);
xor U394 (N_394,In_1004,In_856);
nor U395 (N_395,In_1315,In_789);
or U396 (N_396,In_854,In_1221);
or U397 (N_397,In_577,In_168);
or U398 (N_398,In_585,In_210);
or U399 (N_399,In_1166,In_31);
and U400 (N_400,In_1037,In_728);
nor U401 (N_401,In_990,In_782);
and U402 (N_402,In_374,In_368);
and U403 (N_403,In_306,In_499);
nor U404 (N_404,In_889,In_436);
and U405 (N_405,In_1324,In_565);
xor U406 (N_406,In_673,In_102);
nand U407 (N_407,In_1323,In_1141);
xor U408 (N_408,In_1494,In_864);
nand U409 (N_409,In_858,In_1109);
and U410 (N_410,In_510,In_193);
nor U411 (N_411,In_1426,In_948);
nor U412 (N_412,In_689,In_1263);
or U413 (N_413,In_1427,In_958);
or U414 (N_414,In_107,In_891);
or U415 (N_415,In_714,In_1354);
nand U416 (N_416,In_1322,In_761);
nand U417 (N_417,In_402,In_609);
nand U418 (N_418,In_580,In_1047);
nor U419 (N_419,In_262,In_963);
nand U420 (N_420,In_548,In_328);
nand U421 (N_421,In_570,In_790);
nand U422 (N_422,In_1239,In_183);
nand U423 (N_423,In_977,In_532);
nor U424 (N_424,In_1020,In_1264);
nand U425 (N_425,In_1212,In_636);
nand U426 (N_426,In_781,In_38);
and U427 (N_427,In_97,In_12);
and U428 (N_428,In_844,In_1157);
or U429 (N_429,In_1084,In_540);
or U430 (N_430,In_480,In_279);
and U431 (N_431,In_75,In_100);
or U432 (N_432,In_895,In_530);
nand U433 (N_433,In_486,In_1352);
nand U434 (N_434,In_877,In_19);
or U435 (N_435,In_1287,In_240);
nand U436 (N_436,In_1112,In_434);
nor U437 (N_437,In_1011,In_411);
or U438 (N_438,In_1295,In_94);
nor U439 (N_439,In_647,In_446);
and U440 (N_440,In_225,In_982);
or U441 (N_441,In_535,In_367);
or U442 (N_442,In_592,In_1473);
or U443 (N_443,In_290,In_330);
or U444 (N_444,In_1325,In_1395);
xor U445 (N_445,In_1338,In_1304);
and U446 (N_446,In_124,In_1392);
nor U447 (N_447,In_777,In_382);
or U448 (N_448,In_1306,In_992);
nor U449 (N_449,In_1456,In_1149);
nor U450 (N_450,In_136,In_862);
xnor U451 (N_451,In_387,In_723);
xnor U452 (N_452,In_1138,In_1042);
nand U453 (N_453,In_114,In_869);
and U454 (N_454,In_380,In_23);
nor U455 (N_455,In_1472,In_404);
or U456 (N_456,In_1145,In_533);
or U457 (N_457,In_978,In_829);
or U458 (N_458,In_1181,In_765);
xnor U459 (N_459,In_993,In_1168);
or U460 (N_460,In_400,In_588);
or U461 (N_461,In_1289,In_550);
or U462 (N_462,In_1238,In_747);
or U463 (N_463,In_648,In_1186);
nor U464 (N_464,In_14,In_265);
nor U465 (N_465,In_885,In_110);
or U466 (N_466,In_297,In_1001);
or U467 (N_467,In_1330,In_504);
nor U468 (N_468,In_36,In_123);
or U469 (N_469,In_795,In_601);
nand U470 (N_470,In_1384,In_509);
or U471 (N_471,In_746,In_1044);
or U472 (N_472,In_191,In_1040);
and U473 (N_473,In_821,In_381);
or U474 (N_474,In_311,In_815);
nor U475 (N_475,In_448,In_1479);
or U476 (N_476,In_1386,In_199);
xor U477 (N_477,In_115,In_937);
xor U478 (N_478,In_206,In_116);
and U479 (N_479,In_942,In_1064);
and U480 (N_480,In_302,In_1079);
and U481 (N_481,In_784,In_1407);
nor U482 (N_482,In_981,In_1360);
or U483 (N_483,In_256,In_469);
or U484 (N_484,In_1075,In_1016);
or U485 (N_485,In_1439,In_386);
or U486 (N_486,In_1409,In_919);
or U487 (N_487,In_489,In_269);
xnor U488 (N_488,In_1497,In_665);
nor U489 (N_489,In_650,In_1451);
nor U490 (N_490,In_1220,In_802);
or U491 (N_491,In_640,In_226);
and U492 (N_492,In_232,In_987);
nand U493 (N_493,In_16,In_162);
or U494 (N_494,In_886,In_546);
and U495 (N_495,In_373,In_466);
or U496 (N_496,In_1115,In_316);
and U497 (N_497,In_514,In_419);
xor U498 (N_498,In_1476,In_502);
nor U499 (N_499,In_534,In_563);
or U500 (N_500,In_1059,In_555);
or U501 (N_501,In_1130,In_1391);
nand U502 (N_502,In_430,In_433);
nor U503 (N_503,In_1178,In_410);
and U504 (N_504,In_642,In_1148);
xnor U505 (N_505,In_176,In_138);
or U506 (N_506,In_42,In_943);
nor U507 (N_507,In_1429,In_1431);
and U508 (N_508,In_1272,In_904);
or U509 (N_509,In_568,In_1120);
nand U510 (N_510,In_61,In_1358);
nand U511 (N_511,In_1258,In_1158);
nor U512 (N_512,In_460,In_157);
xor U513 (N_513,In_229,In_873);
or U514 (N_514,In_465,In_688);
nand U515 (N_515,In_1113,In_539);
nor U516 (N_516,In_1379,In_1495);
or U517 (N_517,In_270,In_339);
and U518 (N_518,In_1127,In_945);
nor U519 (N_519,In_32,In_612);
and U520 (N_520,In_182,In_204);
nand U521 (N_521,In_1237,In_152);
xor U522 (N_522,In_1257,In_375);
nor U523 (N_523,In_536,In_1443);
nand U524 (N_524,In_827,In_1028);
nor U525 (N_525,In_287,In_542);
or U526 (N_526,In_64,In_263);
or U527 (N_527,In_887,In_996);
and U528 (N_528,In_120,In_449);
or U529 (N_529,In_344,In_699);
nand U530 (N_530,In_106,In_1062);
or U531 (N_531,In_911,In_880);
nand U532 (N_532,In_1345,In_1006);
xor U533 (N_533,In_1485,In_1065);
and U534 (N_534,In_1466,In_918);
nor U535 (N_535,In_360,In_44);
nor U536 (N_536,In_358,In_1483);
or U537 (N_537,In_1026,In_228);
and U538 (N_538,In_1097,In_1329);
nor U539 (N_539,In_1432,In_1293);
or U540 (N_540,In_591,In_573);
nand U541 (N_541,In_491,In_111);
or U542 (N_542,In_445,In_1214);
and U543 (N_543,In_933,In_949);
or U544 (N_544,In_383,In_701);
nor U545 (N_545,In_600,In_721);
and U546 (N_546,In_51,In_187);
xor U547 (N_547,In_1009,In_1153);
xnor U548 (N_548,In_845,In_453);
nand U549 (N_549,In_151,In_1245);
nor U550 (N_550,In_1393,In_468);
and U551 (N_551,In_90,In_694);
nand U552 (N_552,In_71,In_1082);
nand U553 (N_553,In_1070,In_1139);
and U554 (N_554,In_237,In_1190);
or U555 (N_555,In_807,In_712);
or U556 (N_556,In_639,In_649);
and U557 (N_557,In_908,In_155);
nor U558 (N_558,In_250,In_141);
nor U559 (N_559,In_745,In_882);
nand U560 (N_560,In_1182,In_1402);
and U561 (N_561,In_271,In_1063);
nand U562 (N_562,In_1438,In_720);
or U563 (N_563,In_235,In_1055);
or U564 (N_564,In_1270,In_1184);
and U565 (N_565,In_495,In_350);
and U566 (N_566,In_923,In_1170);
nor U567 (N_567,In_1481,In_602);
nand U568 (N_568,In_1188,In_498);
or U569 (N_569,In_170,In_1033);
nand U570 (N_570,In_146,In_659);
nand U571 (N_571,In_1416,In_672);
nor U572 (N_572,In_661,In_1027);
and U573 (N_573,In_999,In_40);
or U574 (N_574,In_342,In_223);
and U575 (N_575,In_447,In_444);
and U576 (N_576,In_823,In_1457);
nand U577 (N_577,In_1100,In_305);
and U578 (N_578,In_58,In_799);
or U579 (N_579,In_710,In_617);
nor U580 (N_580,In_596,In_748);
or U581 (N_581,In_974,In_1418);
or U582 (N_582,In_91,In_544);
xnor U583 (N_583,In_1359,In_1122);
or U584 (N_584,In_1351,In_15);
nand U585 (N_585,In_664,In_1119);
or U586 (N_586,In_257,In_1234);
and U587 (N_587,In_876,In_621);
nand U588 (N_588,In_1331,In_875);
xor U589 (N_589,In_855,In_215);
xor U590 (N_590,In_634,In_763);
or U591 (N_591,In_178,In_1311);
and U592 (N_592,In_1425,In_626);
nand U593 (N_593,In_1363,In_1101);
nor U594 (N_594,In_1269,In_1297);
xnor U595 (N_595,In_557,In_1414);
nand U596 (N_596,In_1151,In_89);
or U597 (N_597,In_774,In_1183);
or U598 (N_598,In_459,In_653);
and U599 (N_599,In_1283,In_1081);
or U600 (N_600,In_692,In_800);
nor U601 (N_601,In_135,In_1096);
nor U602 (N_602,In_1454,In_832);
xor U603 (N_603,In_1171,In_894);
nand U604 (N_604,In_428,In_62);
and U605 (N_605,In_160,In_674);
nor U606 (N_606,In_838,In_1150);
or U607 (N_607,In_708,In_1434);
and U608 (N_608,In_1420,In_490);
nor U609 (N_609,In_935,In_666);
nor U610 (N_610,In_946,In_1169);
and U611 (N_611,In_1198,In_968);
nand U612 (N_612,In_803,In_1388);
or U613 (N_613,In_931,In_105);
and U614 (N_614,In_76,In_255);
or U615 (N_615,In_1203,In_331);
nor U616 (N_616,In_112,In_1240);
xnor U617 (N_617,In_979,In_1461);
and U618 (N_618,In_1,In_292);
or U619 (N_619,In_1154,In_852);
or U620 (N_620,In_1133,In_3);
or U621 (N_621,In_614,In_1467);
nand U622 (N_622,In_169,In_1455);
and U623 (N_623,In_611,In_1014);
nand U624 (N_624,In_303,In_1207);
nand U625 (N_625,In_1299,In_1196);
or U626 (N_626,In_1470,In_787);
and U627 (N_627,In_294,In_587);
nand U628 (N_628,In_1375,In_1230);
nor U629 (N_629,In_556,In_553);
and U630 (N_630,In_167,In_333);
nand U631 (N_631,In_730,In_1248);
nand U632 (N_632,In_244,In_814);
and U633 (N_633,In_681,In_1023);
nand U634 (N_634,In_1246,In_817);
or U635 (N_635,In_1135,In_395);
nand U636 (N_636,In_242,In_734);
nor U637 (N_637,In_503,In_547);
and U638 (N_638,In_214,In_1273);
nand U639 (N_639,In_312,In_43);
xnor U640 (N_640,In_349,In_508);
xor U641 (N_641,In_816,In_791);
or U642 (N_642,In_1057,In_757);
nand U643 (N_643,In_861,In_440);
nand U644 (N_644,In_37,In_929);
nand U645 (N_645,In_645,In_442);
or U646 (N_646,In_1458,In_203);
xor U647 (N_647,In_868,In_392);
and U648 (N_648,In_1224,In_1279);
nand U649 (N_649,In_186,In_1069);
and U650 (N_650,In_888,In_984);
nand U651 (N_651,In_1189,In_1437);
and U652 (N_652,In_29,In_643);
nand U653 (N_653,In_134,In_778);
or U654 (N_654,In_196,In_693);
nor U655 (N_655,In_1480,In_1125);
and U656 (N_656,In_884,In_780);
nand U657 (N_657,In_897,In_1286);
nand U658 (N_658,In_443,In_396);
nor U659 (N_659,In_983,In_1278);
nor U660 (N_660,In_690,In_1498);
or U661 (N_661,In_68,In_348);
nand U662 (N_662,In_1413,In_725);
xor U663 (N_663,In_528,In_1344);
or U664 (N_664,In_1136,In_657);
nand U665 (N_665,In_70,In_562);
or U666 (N_666,In_1152,In_524);
or U667 (N_667,In_209,In_0);
and U668 (N_668,In_956,In_280);
or U669 (N_669,In_1440,In_317);
nand U670 (N_670,In_960,In_759);
or U671 (N_671,In_1252,In_1194);
and U672 (N_672,In_1128,In_878);
nor U673 (N_673,In_1160,In_1243);
or U674 (N_674,In_1129,In_1007);
nand U675 (N_675,In_334,In_1159);
and U676 (N_676,In_1107,In_1417);
nor U677 (N_677,In_1045,In_932);
and U678 (N_678,In_327,In_805);
xnor U679 (N_679,In_785,In_988);
nand U680 (N_680,In_1300,In_1067);
and U681 (N_681,In_1002,In_622);
nor U682 (N_682,In_1218,In_198);
and U683 (N_683,In_149,In_409);
nor U684 (N_684,In_195,In_1428);
nand U685 (N_685,In_1208,In_597);
xnor U686 (N_686,In_181,In_95);
nor U687 (N_687,In_295,In_313);
nand U688 (N_688,In_325,In_103);
xor U689 (N_689,In_836,In_227);
xnor U690 (N_690,In_1072,In_1226);
nand U691 (N_691,In_1444,In_379);
nand U692 (N_692,In_1267,In_525);
or U693 (N_693,In_289,In_1406);
nor U694 (N_694,In_1058,In_34);
or U695 (N_695,In_1452,In_355);
xor U696 (N_696,In_840,In_749);
or U697 (N_697,In_598,In_1366);
xnor U698 (N_698,In_962,In_566);
nand U699 (N_699,In_10,In_464);
nor U700 (N_700,In_48,In_564);
or U701 (N_701,In_119,In_174);
xnor U702 (N_702,In_951,In_1015);
and U703 (N_703,In_939,In_143);
or U704 (N_704,In_1334,In_825);
and U705 (N_705,In_1339,In_808);
and U706 (N_706,In_6,In_28);
nor U707 (N_707,In_1405,In_231);
xnor U708 (N_708,In_252,In_583);
nand U709 (N_709,In_211,In_217);
nor U710 (N_710,In_668,In_767);
nand U711 (N_711,In_83,In_1385);
and U712 (N_712,In_567,In_1389);
xnor U713 (N_713,In_733,In_1103);
and U714 (N_714,In_1421,In_185);
xnor U715 (N_715,In_93,In_65);
and U716 (N_716,In_1054,In_709);
or U717 (N_717,In_1296,In_764);
nor U718 (N_718,In_472,In_1474);
nor U719 (N_719,In_1049,In_798);
nand U720 (N_720,In_1376,In_364);
nor U721 (N_721,In_283,In_1164);
nor U722 (N_722,In_738,In_1309);
and U723 (N_723,In_736,In_715);
nand U724 (N_724,In_309,In_496);
or U725 (N_725,In_345,In_936);
nand U726 (N_726,In_479,In_1247);
nand U727 (N_727,In_711,In_1012);
nor U728 (N_728,In_441,In_1450);
nor U729 (N_729,In_523,In_705);
nor U730 (N_730,In_1493,In_22);
and U731 (N_731,In_574,In_1320);
and U732 (N_732,In_972,In_900);
and U733 (N_733,In_284,In_684);
nor U734 (N_734,In_971,In_1106);
or U735 (N_735,In_716,In_820);
nand U736 (N_736,In_398,In_63);
nand U737 (N_737,In_471,In_941);
nand U738 (N_738,In_153,In_835);
xor U739 (N_739,In_1408,In_679);
or U740 (N_740,In_307,In_424);
or U741 (N_741,In_1083,In_422);
or U742 (N_742,In_117,In_847);
or U743 (N_743,In_493,In_1250);
nand U744 (N_744,In_1201,In_25);
or U745 (N_745,In_1143,In_966);
and U746 (N_746,In_973,In_50);
nand U747 (N_747,In_1463,In_1288);
or U748 (N_748,In_1314,In_695);
nand U749 (N_749,In_924,In_108);
or U750 (N_750,In_581,In_472);
nor U751 (N_751,In_567,In_1164);
nor U752 (N_752,In_76,In_1321);
or U753 (N_753,In_930,In_1349);
nand U754 (N_754,In_1368,In_371);
xor U755 (N_755,In_1442,In_481);
nor U756 (N_756,In_1266,In_306);
and U757 (N_757,In_431,In_735);
xor U758 (N_758,In_1169,In_568);
or U759 (N_759,In_1494,In_1046);
and U760 (N_760,In_825,In_458);
nand U761 (N_761,In_208,In_844);
nand U762 (N_762,In_1307,In_394);
and U763 (N_763,In_934,In_1443);
xnor U764 (N_764,In_1443,In_909);
and U765 (N_765,In_1307,In_535);
or U766 (N_766,In_933,In_410);
or U767 (N_767,In_357,In_661);
and U768 (N_768,In_738,In_1316);
nand U769 (N_769,In_1394,In_50);
or U770 (N_770,In_354,In_155);
nor U771 (N_771,In_236,In_992);
and U772 (N_772,In_1123,In_1350);
or U773 (N_773,In_1222,In_549);
and U774 (N_774,In_700,In_1157);
or U775 (N_775,In_772,In_1150);
and U776 (N_776,In_124,In_622);
nor U777 (N_777,In_1168,In_1460);
nand U778 (N_778,In_1461,In_273);
nor U779 (N_779,In_564,In_1473);
or U780 (N_780,In_50,In_705);
and U781 (N_781,In_836,In_45);
and U782 (N_782,In_1469,In_1163);
nor U783 (N_783,In_500,In_876);
and U784 (N_784,In_1250,In_1040);
or U785 (N_785,In_301,In_116);
nor U786 (N_786,In_773,In_757);
and U787 (N_787,In_1165,In_908);
nand U788 (N_788,In_142,In_945);
and U789 (N_789,In_414,In_1244);
or U790 (N_790,In_173,In_1072);
or U791 (N_791,In_1406,In_498);
nor U792 (N_792,In_441,In_801);
nand U793 (N_793,In_224,In_1492);
and U794 (N_794,In_714,In_772);
and U795 (N_795,In_682,In_922);
or U796 (N_796,In_709,In_783);
or U797 (N_797,In_386,In_860);
and U798 (N_798,In_610,In_402);
and U799 (N_799,In_1035,In_1165);
nor U800 (N_800,In_146,In_1447);
nor U801 (N_801,In_797,In_418);
nand U802 (N_802,In_547,In_765);
xnor U803 (N_803,In_95,In_1435);
or U804 (N_804,In_1367,In_993);
nor U805 (N_805,In_141,In_998);
and U806 (N_806,In_114,In_134);
xor U807 (N_807,In_1176,In_1242);
and U808 (N_808,In_151,In_184);
and U809 (N_809,In_316,In_494);
or U810 (N_810,In_708,In_180);
xnor U811 (N_811,In_346,In_14);
or U812 (N_812,In_601,In_1104);
nand U813 (N_813,In_460,In_411);
xor U814 (N_814,In_654,In_1416);
nor U815 (N_815,In_1271,In_1208);
and U816 (N_816,In_900,In_1017);
or U817 (N_817,In_542,In_918);
nor U818 (N_818,In_937,In_1101);
xor U819 (N_819,In_238,In_186);
and U820 (N_820,In_1233,In_123);
and U821 (N_821,In_879,In_1345);
nor U822 (N_822,In_1224,In_302);
nor U823 (N_823,In_997,In_206);
nor U824 (N_824,In_184,In_378);
and U825 (N_825,In_1007,In_1016);
or U826 (N_826,In_1456,In_688);
or U827 (N_827,In_361,In_442);
or U828 (N_828,In_1260,In_1451);
nand U829 (N_829,In_1478,In_607);
nand U830 (N_830,In_543,In_784);
nor U831 (N_831,In_633,In_606);
nor U832 (N_832,In_194,In_19);
nor U833 (N_833,In_574,In_1047);
nand U834 (N_834,In_235,In_1089);
nand U835 (N_835,In_12,In_28);
nand U836 (N_836,In_567,In_167);
nor U837 (N_837,In_107,In_1246);
nand U838 (N_838,In_768,In_1350);
nor U839 (N_839,In_593,In_1482);
or U840 (N_840,In_426,In_669);
nand U841 (N_841,In_36,In_1421);
xnor U842 (N_842,In_623,In_1440);
or U843 (N_843,In_1156,In_19);
nor U844 (N_844,In_435,In_884);
nor U845 (N_845,In_147,In_1248);
or U846 (N_846,In_1354,In_1035);
nor U847 (N_847,In_1184,In_1354);
nand U848 (N_848,In_1427,In_290);
xnor U849 (N_849,In_100,In_443);
nor U850 (N_850,In_33,In_1334);
or U851 (N_851,In_1244,In_8);
nor U852 (N_852,In_286,In_1085);
or U853 (N_853,In_248,In_392);
nor U854 (N_854,In_552,In_480);
nand U855 (N_855,In_1002,In_565);
nand U856 (N_856,In_21,In_1125);
xnor U857 (N_857,In_666,In_441);
or U858 (N_858,In_1361,In_481);
nand U859 (N_859,In_1024,In_964);
nand U860 (N_860,In_1085,In_544);
nor U861 (N_861,In_1341,In_1199);
nor U862 (N_862,In_146,In_286);
nand U863 (N_863,In_117,In_1058);
nor U864 (N_864,In_885,In_571);
nor U865 (N_865,In_745,In_1013);
and U866 (N_866,In_188,In_1041);
and U867 (N_867,In_1498,In_733);
nor U868 (N_868,In_543,In_1172);
nand U869 (N_869,In_242,In_452);
and U870 (N_870,In_196,In_513);
and U871 (N_871,In_283,In_1113);
nor U872 (N_872,In_327,In_516);
nor U873 (N_873,In_1232,In_32);
nand U874 (N_874,In_90,In_531);
or U875 (N_875,In_518,In_63);
nor U876 (N_876,In_427,In_78);
nor U877 (N_877,In_122,In_419);
nor U878 (N_878,In_277,In_1394);
or U879 (N_879,In_737,In_1240);
nand U880 (N_880,In_616,In_833);
and U881 (N_881,In_938,In_1300);
nor U882 (N_882,In_706,In_747);
nand U883 (N_883,In_445,In_574);
nand U884 (N_884,In_155,In_1278);
or U885 (N_885,In_142,In_257);
or U886 (N_886,In_1392,In_1251);
nand U887 (N_887,In_1029,In_146);
and U888 (N_888,In_474,In_737);
nor U889 (N_889,In_966,In_1102);
xor U890 (N_890,In_395,In_299);
and U891 (N_891,In_1266,In_504);
xnor U892 (N_892,In_152,In_134);
xnor U893 (N_893,In_277,In_998);
nand U894 (N_894,In_1313,In_474);
and U895 (N_895,In_74,In_473);
or U896 (N_896,In_586,In_1255);
nand U897 (N_897,In_243,In_1152);
nor U898 (N_898,In_640,In_666);
nand U899 (N_899,In_114,In_495);
xor U900 (N_900,In_985,In_1247);
nand U901 (N_901,In_1284,In_175);
and U902 (N_902,In_612,In_16);
nor U903 (N_903,In_1445,In_1073);
nand U904 (N_904,In_394,In_11);
or U905 (N_905,In_1149,In_1345);
or U906 (N_906,In_95,In_292);
or U907 (N_907,In_777,In_756);
or U908 (N_908,In_50,In_900);
or U909 (N_909,In_189,In_285);
nand U910 (N_910,In_1071,In_1251);
or U911 (N_911,In_936,In_629);
and U912 (N_912,In_976,In_1342);
nor U913 (N_913,In_1179,In_757);
nand U914 (N_914,In_1008,In_707);
nor U915 (N_915,In_295,In_376);
or U916 (N_916,In_464,In_1483);
and U917 (N_917,In_739,In_635);
or U918 (N_918,In_163,In_233);
nor U919 (N_919,In_1390,In_501);
nor U920 (N_920,In_1113,In_579);
nand U921 (N_921,In_340,In_503);
nor U922 (N_922,In_1061,In_297);
or U923 (N_923,In_1493,In_149);
nor U924 (N_924,In_228,In_1406);
nand U925 (N_925,In_985,In_1040);
nand U926 (N_926,In_330,In_708);
xnor U927 (N_927,In_993,In_1322);
nand U928 (N_928,In_1496,In_1203);
or U929 (N_929,In_586,In_958);
nand U930 (N_930,In_839,In_1165);
nand U931 (N_931,In_197,In_234);
nor U932 (N_932,In_310,In_972);
xnor U933 (N_933,In_106,In_751);
or U934 (N_934,In_143,In_750);
xnor U935 (N_935,In_652,In_315);
nand U936 (N_936,In_1426,In_1012);
xnor U937 (N_937,In_983,In_617);
nor U938 (N_938,In_1057,In_253);
or U939 (N_939,In_400,In_1142);
or U940 (N_940,In_477,In_596);
nand U941 (N_941,In_612,In_665);
or U942 (N_942,In_1117,In_779);
and U943 (N_943,In_253,In_1170);
and U944 (N_944,In_1390,In_431);
nand U945 (N_945,In_226,In_618);
nand U946 (N_946,In_654,In_896);
or U947 (N_947,In_763,In_641);
xor U948 (N_948,In_1437,In_1407);
nor U949 (N_949,In_583,In_1414);
nand U950 (N_950,In_1103,In_1458);
and U951 (N_951,In_657,In_4);
nand U952 (N_952,In_141,In_940);
nor U953 (N_953,In_1199,In_449);
or U954 (N_954,In_163,In_1271);
nand U955 (N_955,In_832,In_1124);
or U956 (N_956,In_241,In_1375);
and U957 (N_957,In_1051,In_491);
nand U958 (N_958,In_1302,In_271);
and U959 (N_959,In_718,In_1329);
nor U960 (N_960,In_818,In_734);
nor U961 (N_961,In_864,In_694);
and U962 (N_962,In_23,In_565);
and U963 (N_963,In_189,In_360);
nand U964 (N_964,In_1227,In_849);
nor U965 (N_965,In_931,In_58);
or U966 (N_966,In_142,In_1135);
nand U967 (N_967,In_703,In_697);
and U968 (N_968,In_403,In_621);
and U969 (N_969,In_1439,In_536);
or U970 (N_970,In_524,In_1233);
nor U971 (N_971,In_1093,In_1235);
and U972 (N_972,In_422,In_631);
and U973 (N_973,In_71,In_912);
and U974 (N_974,In_934,In_57);
and U975 (N_975,In_98,In_1199);
nand U976 (N_976,In_412,In_920);
and U977 (N_977,In_763,In_1036);
and U978 (N_978,In_653,In_338);
or U979 (N_979,In_1257,In_639);
nand U980 (N_980,In_1268,In_1017);
and U981 (N_981,In_988,In_1016);
xnor U982 (N_982,In_88,In_1016);
xnor U983 (N_983,In_1,In_734);
xnor U984 (N_984,In_716,In_1068);
and U985 (N_985,In_1183,In_571);
or U986 (N_986,In_670,In_332);
or U987 (N_987,In_702,In_624);
nor U988 (N_988,In_953,In_952);
nand U989 (N_989,In_761,In_1275);
and U990 (N_990,In_1391,In_311);
and U991 (N_991,In_252,In_1409);
nand U992 (N_992,In_506,In_1377);
and U993 (N_993,In_1066,In_355);
or U994 (N_994,In_1152,In_1361);
nor U995 (N_995,In_770,In_1265);
nand U996 (N_996,In_1103,In_293);
or U997 (N_997,In_683,In_524);
nor U998 (N_998,In_858,In_677);
or U999 (N_999,In_402,In_1482);
or U1000 (N_1000,In_492,In_1417);
and U1001 (N_1001,In_1253,In_901);
or U1002 (N_1002,In_607,In_1121);
xnor U1003 (N_1003,In_1258,In_1242);
or U1004 (N_1004,In_685,In_945);
nor U1005 (N_1005,In_719,In_97);
nand U1006 (N_1006,In_697,In_897);
nand U1007 (N_1007,In_648,In_54);
xnor U1008 (N_1008,In_121,In_1050);
nand U1009 (N_1009,In_423,In_1106);
nor U1010 (N_1010,In_1379,In_73);
nor U1011 (N_1011,In_790,In_340);
nor U1012 (N_1012,In_1340,In_931);
nor U1013 (N_1013,In_1495,In_633);
nor U1014 (N_1014,In_686,In_909);
nand U1015 (N_1015,In_259,In_1395);
xor U1016 (N_1016,In_41,In_980);
xnor U1017 (N_1017,In_726,In_1373);
or U1018 (N_1018,In_61,In_682);
nor U1019 (N_1019,In_261,In_838);
nor U1020 (N_1020,In_567,In_579);
nand U1021 (N_1021,In_141,In_1396);
and U1022 (N_1022,In_129,In_690);
nor U1023 (N_1023,In_39,In_383);
nand U1024 (N_1024,In_605,In_119);
xor U1025 (N_1025,In_222,In_773);
nor U1026 (N_1026,In_257,In_651);
or U1027 (N_1027,In_81,In_630);
or U1028 (N_1028,In_752,In_965);
or U1029 (N_1029,In_497,In_991);
xor U1030 (N_1030,In_1222,In_1440);
or U1031 (N_1031,In_680,In_30);
nor U1032 (N_1032,In_185,In_649);
xnor U1033 (N_1033,In_1192,In_360);
and U1034 (N_1034,In_1309,In_401);
nand U1035 (N_1035,In_1324,In_430);
and U1036 (N_1036,In_809,In_1165);
nand U1037 (N_1037,In_1470,In_1184);
and U1038 (N_1038,In_1499,In_189);
and U1039 (N_1039,In_551,In_1115);
and U1040 (N_1040,In_1483,In_1359);
and U1041 (N_1041,In_287,In_1249);
nor U1042 (N_1042,In_376,In_974);
nor U1043 (N_1043,In_234,In_957);
or U1044 (N_1044,In_553,In_544);
nor U1045 (N_1045,In_77,In_358);
nand U1046 (N_1046,In_822,In_259);
nand U1047 (N_1047,In_1314,In_1202);
xnor U1048 (N_1048,In_54,In_896);
or U1049 (N_1049,In_460,In_345);
xor U1050 (N_1050,In_484,In_758);
and U1051 (N_1051,In_64,In_1474);
or U1052 (N_1052,In_814,In_752);
nand U1053 (N_1053,In_566,In_1470);
or U1054 (N_1054,In_293,In_1114);
or U1055 (N_1055,In_1291,In_1105);
and U1056 (N_1056,In_1162,In_303);
nand U1057 (N_1057,In_1482,In_1269);
nor U1058 (N_1058,In_1069,In_817);
or U1059 (N_1059,In_972,In_1192);
nand U1060 (N_1060,In_1020,In_1383);
xnor U1061 (N_1061,In_1299,In_757);
and U1062 (N_1062,In_910,In_247);
nand U1063 (N_1063,In_1381,In_461);
and U1064 (N_1064,In_1284,In_533);
or U1065 (N_1065,In_274,In_1439);
or U1066 (N_1066,In_662,In_702);
or U1067 (N_1067,In_298,In_90);
and U1068 (N_1068,In_443,In_877);
nor U1069 (N_1069,In_637,In_1243);
nand U1070 (N_1070,In_240,In_1208);
nor U1071 (N_1071,In_1286,In_499);
or U1072 (N_1072,In_1307,In_1420);
and U1073 (N_1073,In_909,In_857);
or U1074 (N_1074,In_1200,In_457);
nand U1075 (N_1075,In_1444,In_398);
or U1076 (N_1076,In_164,In_399);
nand U1077 (N_1077,In_1366,In_766);
nand U1078 (N_1078,In_367,In_583);
or U1079 (N_1079,In_405,In_209);
or U1080 (N_1080,In_676,In_243);
nor U1081 (N_1081,In_1056,In_1487);
nand U1082 (N_1082,In_98,In_547);
nand U1083 (N_1083,In_765,In_270);
xor U1084 (N_1084,In_621,In_295);
nor U1085 (N_1085,In_1256,In_1095);
and U1086 (N_1086,In_411,In_1144);
or U1087 (N_1087,In_555,In_194);
nor U1088 (N_1088,In_1040,In_1039);
nand U1089 (N_1089,In_490,In_1282);
and U1090 (N_1090,In_84,In_325);
nand U1091 (N_1091,In_482,In_1185);
and U1092 (N_1092,In_1404,In_31);
nand U1093 (N_1093,In_478,In_717);
and U1094 (N_1094,In_407,In_1093);
or U1095 (N_1095,In_500,In_353);
nor U1096 (N_1096,In_615,In_1426);
xor U1097 (N_1097,In_641,In_1130);
or U1098 (N_1098,In_812,In_144);
nor U1099 (N_1099,In_316,In_732);
and U1100 (N_1100,In_1253,In_1473);
and U1101 (N_1101,In_32,In_191);
nor U1102 (N_1102,In_972,In_1048);
nor U1103 (N_1103,In_1186,In_794);
nor U1104 (N_1104,In_898,In_661);
and U1105 (N_1105,In_1074,In_813);
and U1106 (N_1106,In_779,In_96);
nand U1107 (N_1107,In_1144,In_929);
nand U1108 (N_1108,In_556,In_1338);
or U1109 (N_1109,In_890,In_707);
nor U1110 (N_1110,In_520,In_388);
nand U1111 (N_1111,In_1322,In_471);
nor U1112 (N_1112,In_1029,In_435);
nor U1113 (N_1113,In_703,In_1461);
nor U1114 (N_1114,In_1380,In_24);
nand U1115 (N_1115,In_1192,In_1020);
xnor U1116 (N_1116,In_365,In_907);
or U1117 (N_1117,In_857,In_1426);
or U1118 (N_1118,In_1219,In_1384);
or U1119 (N_1119,In_1458,In_1420);
xor U1120 (N_1120,In_212,In_1078);
nand U1121 (N_1121,In_639,In_869);
nor U1122 (N_1122,In_1272,In_1345);
or U1123 (N_1123,In_586,In_625);
nor U1124 (N_1124,In_873,In_1412);
and U1125 (N_1125,In_212,In_1290);
nor U1126 (N_1126,In_797,In_1330);
nand U1127 (N_1127,In_1239,In_173);
xor U1128 (N_1128,In_1393,In_1128);
nand U1129 (N_1129,In_228,In_1155);
nor U1130 (N_1130,In_1383,In_152);
or U1131 (N_1131,In_1296,In_964);
xnor U1132 (N_1132,In_101,In_1235);
and U1133 (N_1133,In_552,In_1083);
and U1134 (N_1134,In_93,In_668);
nor U1135 (N_1135,In_233,In_1063);
or U1136 (N_1136,In_608,In_1030);
nand U1137 (N_1137,In_1020,In_254);
nor U1138 (N_1138,In_1298,In_603);
nand U1139 (N_1139,In_7,In_681);
and U1140 (N_1140,In_470,In_533);
nand U1141 (N_1141,In_755,In_1300);
or U1142 (N_1142,In_1125,In_29);
or U1143 (N_1143,In_1210,In_1212);
xnor U1144 (N_1144,In_608,In_72);
or U1145 (N_1145,In_880,In_971);
or U1146 (N_1146,In_449,In_329);
nand U1147 (N_1147,In_655,In_211);
xnor U1148 (N_1148,In_1353,In_1203);
and U1149 (N_1149,In_1067,In_1107);
xnor U1150 (N_1150,In_874,In_1132);
nand U1151 (N_1151,In_1258,In_1121);
nand U1152 (N_1152,In_840,In_1323);
or U1153 (N_1153,In_197,In_213);
and U1154 (N_1154,In_862,In_184);
nor U1155 (N_1155,In_323,In_275);
xor U1156 (N_1156,In_1346,In_1304);
or U1157 (N_1157,In_71,In_209);
xor U1158 (N_1158,In_692,In_1264);
nand U1159 (N_1159,In_1035,In_262);
nand U1160 (N_1160,In_758,In_1411);
or U1161 (N_1161,In_621,In_263);
nor U1162 (N_1162,In_75,In_682);
nor U1163 (N_1163,In_517,In_1171);
or U1164 (N_1164,In_1455,In_610);
and U1165 (N_1165,In_1147,In_1285);
nor U1166 (N_1166,In_1128,In_1469);
and U1167 (N_1167,In_179,In_1377);
xnor U1168 (N_1168,In_1440,In_1178);
nor U1169 (N_1169,In_457,In_519);
and U1170 (N_1170,In_388,In_307);
or U1171 (N_1171,In_426,In_559);
or U1172 (N_1172,In_1144,In_739);
and U1173 (N_1173,In_144,In_366);
nor U1174 (N_1174,In_971,In_630);
nor U1175 (N_1175,In_347,In_884);
nor U1176 (N_1176,In_43,In_125);
nor U1177 (N_1177,In_1177,In_125);
or U1178 (N_1178,In_1255,In_136);
nand U1179 (N_1179,In_1379,In_506);
nor U1180 (N_1180,In_1140,In_841);
or U1181 (N_1181,In_1009,In_1059);
nor U1182 (N_1182,In_1410,In_1312);
nand U1183 (N_1183,In_1293,In_1116);
xnor U1184 (N_1184,In_721,In_1062);
nand U1185 (N_1185,In_535,In_344);
or U1186 (N_1186,In_625,In_853);
or U1187 (N_1187,In_630,In_809);
nor U1188 (N_1188,In_1139,In_1078);
or U1189 (N_1189,In_332,In_1440);
nor U1190 (N_1190,In_928,In_587);
and U1191 (N_1191,In_258,In_660);
nor U1192 (N_1192,In_836,In_369);
nand U1193 (N_1193,In_1392,In_74);
or U1194 (N_1194,In_181,In_676);
nor U1195 (N_1195,In_468,In_843);
and U1196 (N_1196,In_219,In_1148);
or U1197 (N_1197,In_947,In_692);
and U1198 (N_1198,In_448,In_191);
and U1199 (N_1199,In_611,In_1118);
xnor U1200 (N_1200,In_158,In_1358);
nand U1201 (N_1201,In_1035,In_692);
xor U1202 (N_1202,In_572,In_1134);
and U1203 (N_1203,In_142,In_1294);
or U1204 (N_1204,In_799,In_118);
or U1205 (N_1205,In_1293,In_931);
xor U1206 (N_1206,In_1333,In_641);
nor U1207 (N_1207,In_591,In_815);
and U1208 (N_1208,In_1190,In_276);
or U1209 (N_1209,In_272,In_178);
nand U1210 (N_1210,In_625,In_152);
or U1211 (N_1211,In_1198,In_622);
nor U1212 (N_1212,In_51,In_246);
nand U1213 (N_1213,In_1181,In_730);
nor U1214 (N_1214,In_1236,In_1034);
and U1215 (N_1215,In_931,In_1419);
or U1216 (N_1216,In_1290,In_1013);
and U1217 (N_1217,In_122,In_466);
or U1218 (N_1218,In_272,In_104);
nand U1219 (N_1219,In_199,In_236);
nand U1220 (N_1220,In_1028,In_133);
and U1221 (N_1221,In_1133,In_1395);
and U1222 (N_1222,In_1006,In_613);
and U1223 (N_1223,In_1445,In_1218);
or U1224 (N_1224,In_778,In_220);
nand U1225 (N_1225,In_487,In_945);
nand U1226 (N_1226,In_856,In_902);
or U1227 (N_1227,In_73,In_1045);
and U1228 (N_1228,In_187,In_1451);
nor U1229 (N_1229,In_229,In_1128);
nor U1230 (N_1230,In_980,In_910);
nor U1231 (N_1231,In_86,In_1244);
nor U1232 (N_1232,In_190,In_759);
or U1233 (N_1233,In_719,In_1471);
nand U1234 (N_1234,In_1485,In_204);
nor U1235 (N_1235,In_487,In_885);
and U1236 (N_1236,In_632,In_366);
nor U1237 (N_1237,In_324,In_594);
nor U1238 (N_1238,In_685,In_1070);
and U1239 (N_1239,In_318,In_444);
nor U1240 (N_1240,In_819,In_1113);
nor U1241 (N_1241,In_995,In_1358);
nor U1242 (N_1242,In_1307,In_1461);
nand U1243 (N_1243,In_929,In_1145);
nor U1244 (N_1244,In_610,In_457);
and U1245 (N_1245,In_25,In_717);
nand U1246 (N_1246,In_634,In_764);
nand U1247 (N_1247,In_890,In_634);
nand U1248 (N_1248,In_448,In_377);
xnor U1249 (N_1249,In_698,In_521);
or U1250 (N_1250,In_5,In_1061);
nor U1251 (N_1251,In_89,In_565);
nand U1252 (N_1252,In_420,In_652);
or U1253 (N_1253,In_340,In_560);
nand U1254 (N_1254,In_1250,In_899);
xnor U1255 (N_1255,In_1165,In_1047);
and U1256 (N_1256,In_1025,In_1083);
or U1257 (N_1257,In_110,In_822);
or U1258 (N_1258,In_495,In_1354);
and U1259 (N_1259,In_367,In_406);
nand U1260 (N_1260,In_28,In_1231);
or U1261 (N_1261,In_22,In_1293);
and U1262 (N_1262,In_1149,In_587);
and U1263 (N_1263,In_720,In_1411);
nand U1264 (N_1264,In_124,In_1087);
nand U1265 (N_1265,In_1211,In_1309);
and U1266 (N_1266,In_1167,In_186);
or U1267 (N_1267,In_583,In_631);
or U1268 (N_1268,In_757,In_114);
or U1269 (N_1269,In_1462,In_400);
or U1270 (N_1270,In_1072,In_1166);
nor U1271 (N_1271,In_412,In_1193);
or U1272 (N_1272,In_13,In_558);
nor U1273 (N_1273,In_527,In_65);
or U1274 (N_1274,In_469,In_1285);
and U1275 (N_1275,In_475,In_316);
nor U1276 (N_1276,In_443,In_1306);
nand U1277 (N_1277,In_183,In_94);
nand U1278 (N_1278,In_1090,In_1294);
nor U1279 (N_1279,In_409,In_1062);
or U1280 (N_1280,In_1171,In_1470);
and U1281 (N_1281,In_1015,In_83);
and U1282 (N_1282,In_1331,In_1274);
nand U1283 (N_1283,In_821,In_590);
and U1284 (N_1284,In_1380,In_507);
or U1285 (N_1285,In_1390,In_585);
xnor U1286 (N_1286,In_622,In_280);
nand U1287 (N_1287,In_1146,In_783);
nor U1288 (N_1288,In_1337,In_24);
nor U1289 (N_1289,In_517,In_685);
nand U1290 (N_1290,In_1022,In_558);
xnor U1291 (N_1291,In_1337,In_1262);
or U1292 (N_1292,In_1176,In_1106);
or U1293 (N_1293,In_219,In_1165);
nand U1294 (N_1294,In_891,In_946);
xor U1295 (N_1295,In_936,In_976);
nand U1296 (N_1296,In_1364,In_507);
nor U1297 (N_1297,In_531,In_579);
nand U1298 (N_1298,In_53,In_949);
xnor U1299 (N_1299,In_1483,In_773);
nand U1300 (N_1300,In_473,In_730);
nand U1301 (N_1301,In_1449,In_814);
or U1302 (N_1302,In_966,In_771);
or U1303 (N_1303,In_575,In_979);
nor U1304 (N_1304,In_405,In_728);
and U1305 (N_1305,In_420,In_107);
or U1306 (N_1306,In_355,In_1040);
nand U1307 (N_1307,In_1120,In_1041);
or U1308 (N_1308,In_1442,In_977);
and U1309 (N_1309,In_30,In_374);
nand U1310 (N_1310,In_105,In_1389);
nor U1311 (N_1311,In_1245,In_179);
nand U1312 (N_1312,In_986,In_212);
nor U1313 (N_1313,In_1416,In_1172);
nand U1314 (N_1314,In_1471,In_326);
or U1315 (N_1315,In_358,In_625);
or U1316 (N_1316,In_1495,In_1020);
nor U1317 (N_1317,In_1206,In_596);
nand U1318 (N_1318,In_41,In_973);
nand U1319 (N_1319,In_631,In_1314);
and U1320 (N_1320,In_478,In_1408);
nand U1321 (N_1321,In_449,In_966);
or U1322 (N_1322,In_1358,In_1266);
nand U1323 (N_1323,In_630,In_844);
or U1324 (N_1324,In_432,In_697);
nor U1325 (N_1325,In_111,In_284);
or U1326 (N_1326,In_360,In_167);
or U1327 (N_1327,In_284,In_270);
xor U1328 (N_1328,In_351,In_561);
or U1329 (N_1329,In_1474,In_135);
nand U1330 (N_1330,In_1176,In_578);
nand U1331 (N_1331,In_785,In_200);
nor U1332 (N_1332,In_126,In_497);
nand U1333 (N_1333,In_645,In_502);
and U1334 (N_1334,In_551,In_69);
and U1335 (N_1335,In_475,In_448);
nand U1336 (N_1336,In_715,In_721);
or U1337 (N_1337,In_688,In_435);
or U1338 (N_1338,In_826,In_1211);
or U1339 (N_1339,In_619,In_607);
or U1340 (N_1340,In_208,In_941);
nor U1341 (N_1341,In_435,In_560);
or U1342 (N_1342,In_844,In_467);
nand U1343 (N_1343,In_125,In_1138);
xor U1344 (N_1344,In_362,In_925);
nand U1345 (N_1345,In_59,In_176);
nand U1346 (N_1346,In_1443,In_125);
and U1347 (N_1347,In_417,In_385);
xor U1348 (N_1348,In_800,In_23);
xor U1349 (N_1349,In_282,In_77);
nor U1350 (N_1350,In_359,In_1325);
nor U1351 (N_1351,In_1084,In_1093);
and U1352 (N_1352,In_1010,In_540);
or U1353 (N_1353,In_1003,In_276);
nand U1354 (N_1354,In_1108,In_818);
nand U1355 (N_1355,In_284,In_709);
and U1356 (N_1356,In_741,In_606);
nand U1357 (N_1357,In_532,In_587);
xor U1358 (N_1358,In_398,In_116);
nor U1359 (N_1359,In_896,In_381);
nor U1360 (N_1360,In_1102,In_1053);
nor U1361 (N_1361,In_1335,In_1215);
nand U1362 (N_1362,In_609,In_134);
nand U1363 (N_1363,In_651,In_16);
or U1364 (N_1364,In_1252,In_67);
nor U1365 (N_1365,In_436,In_803);
and U1366 (N_1366,In_583,In_703);
or U1367 (N_1367,In_860,In_1331);
nor U1368 (N_1368,In_748,In_1386);
nand U1369 (N_1369,In_550,In_150);
nand U1370 (N_1370,In_180,In_1158);
nor U1371 (N_1371,In_1112,In_1443);
and U1372 (N_1372,In_109,In_916);
nand U1373 (N_1373,In_961,In_214);
or U1374 (N_1374,In_1471,In_1330);
nor U1375 (N_1375,In_779,In_1067);
nor U1376 (N_1376,In_482,In_1390);
and U1377 (N_1377,In_248,In_1382);
nor U1378 (N_1378,In_413,In_1277);
or U1379 (N_1379,In_1318,In_952);
nand U1380 (N_1380,In_878,In_100);
or U1381 (N_1381,In_1394,In_1162);
nor U1382 (N_1382,In_52,In_1075);
or U1383 (N_1383,In_742,In_41);
or U1384 (N_1384,In_443,In_1101);
or U1385 (N_1385,In_1443,In_305);
nor U1386 (N_1386,In_1186,In_472);
xor U1387 (N_1387,In_1000,In_871);
or U1388 (N_1388,In_904,In_1351);
and U1389 (N_1389,In_63,In_1272);
nand U1390 (N_1390,In_655,In_617);
and U1391 (N_1391,In_967,In_1099);
and U1392 (N_1392,In_359,In_417);
or U1393 (N_1393,In_1099,In_1112);
or U1394 (N_1394,In_962,In_1013);
nor U1395 (N_1395,In_869,In_906);
or U1396 (N_1396,In_1018,In_583);
nand U1397 (N_1397,In_809,In_683);
or U1398 (N_1398,In_1202,In_744);
xnor U1399 (N_1399,In_259,In_718);
nand U1400 (N_1400,In_310,In_990);
nor U1401 (N_1401,In_775,In_1362);
xor U1402 (N_1402,In_103,In_49);
or U1403 (N_1403,In_634,In_1059);
nor U1404 (N_1404,In_646,In_541);
xnor U1405 (N_1405,In_50,In_1254);
or U1406 (N_1406,In_644,In_1410);
nand U1407 (N_1407,In_195,In_1450);
nand U1408 (N_1408,In_563,In_1213);
or U1409 (N_1409,In_165,In_546);
and U1410 (N_1410,In_977,In_353);
and U1411 (N_1411,In_333,In_144);
and U1412 (N_1412,In_1403,In_93);
and U1413 (N_1413,In_67,In_1241);
nor U1414 (N_1414,In_1460,In_857);
or U1415 (N_1415,In_1236,In_643);
nor U1416 (N_1416,In_819,In_1149);
nor U1417 (N_1417,In_752,In_817);
or U1418 (N_1418,In_298,In_643);
and U1419 (N_1419,In_492,In_651);
or U1420 (N_1420,In_866,In_913);
nor U1421 (N_1421,In_70,In_342);
or U1422 (N_1422,In_130,In_1482);
nand U1423 (N_1423,In_345,In_1368);
or U1424 (N_1424,In_1138,In_347);
and U1425 (N_1425,In_645,In_328);
and U1426 (N_1426,In_297,In_365);
and U1427 (N_1427,In_712,In_1426);
and U1428 (N_1428,In_415,In_411);
and U1429 (N_1429,In_803,In_1260);
nor U1430 (N_1430,In_307,In_678);
or U1431 (N_1431,In_1399,In_347);
xor U1432 (N_1432,In_423,In_292);
and U1433 (N_1433,In_255,In_648);
or U1434 (N_1434,In_19,In_130);
or U1435 (N_1435,In_139,In_795);
or U1436 (N_1436,In_1425,In_962);
xnor U1437 (N_1437,In_891,In_196);
nor U1438 (N_1438,In_167,In_417);
and U1439 (N_1439,In_432,In_22);
or U1440 (N_1440,In_1170,In_1267);
nor U1441 (N_1441,In_701,In_404);
or U1442 (N_1442,In_1385,In_515);
nor U1443 (N_1443,In_138,In_786);
nor U1444 (N_1444,In_1478,In_455);
or U1445 (N_1445,In_585,In_1389);
nand U1446 (N_1446,In_951,In_238);
and U1447 (N_1447,In_1461,In_288);
and U1448 (N_1448,In_412,In_948);
or U1449 (N_1449,In_238,In_982);
nand U1450 (N_1450,In_709,In_883);
xnor U1451 (N_1451,In_69,In_159);
or U1452 (N_1452,In_726,In_1173);
nor U1453 (N_1453,In_948,In_855);
xnor U1454 (N_1454,In_172,In_277);
and U1455 (N_1455,In_1049,In_916);
nor U1456 (N_1456,In_187,In_200);
nor U1457 (N_1457,In_1018,In_621);
or U1458 (N_1458,In_862,In_1112);
xnor U1459 (N_1459,In_1499,In_1373);
nor U1460 (N_1460,In_1237,In_1478);
nand U1461 (N_1461,In_1331,In_1132);
nand U1462 (N_1462,In_1278,In_1178);
or U1463 (N_1463,In_421,In_473);
nand U1464 (N_1464,In_1118,In_450);
and U1465 (N_1465,In_67,In_308);
nand U1466 (N_1466,In_1376,In_1315);
nand U1467 (N_1467,In_229,In_1394);
nor U1468 (N_1468,In_1379,In_627);
or U1469 (N_1469,In_306,In_585);
nor U1470 (N_1470,In_1451,In_189);
and U1471 (N_1471,In_1189,In_790);
nand U1472 (N_1472,In_87,In_301);
xnor U1473 (N_1473,In_1224,In_144);
and U1474 (N_1474,In_435,In_1265);
nand U1475 (N_1475,In_147,In_1099);
or U1476 (N_1476,In_251,In_1070);
nand U1477 (N_1477,In_369,In_480);
or U1478 (N_1478,In_1248,In_254);
nor U1479 (N_1479,In_600,In_656);
and U1480 (N_1480,In_736,In_1259);
or U1481 (N_1481,In_1321,In_526);
or U1482 (N_1482,In_14,In_996);
and U1483 (N_1483,In_129,In_1381);
or U1484 (N_1484,In_658,In_87);
and U1485 (N_1485,In_491,In_676);
or U1486 (N_1486,In_921,In_1263);
nand U1487 (N_1487,In_784,In_1397);
nand U1488 (N_1488,In_719,In_1370);
nor U1489 (N_1489,In_1087,In_1200);
nor U1490 (N_1490,In_1272,In_1236);
nor U1491 (N_1491,In_1080,In_115);
nand U1492 (N_1492,In_456,In_1246);
nor U1493 (N_1493,In_362,In_784);
nand U1494 (N_1494,In_602,In_1235);
nand U1495 (N_1495,In_762,In_950);
and U1496 (N_1496,In_1373,In_1126);
nand U1497 (N_1497,In_314,In_1208);
xnor U1498 (N_1498,In_548,In_1330);
nor U1499 (N_1499,In_953,In_1188);
nor U1500 (N_1500,N_1393,N_842);
or U1501 (N_1501,N_393,N_131);
xor U1502 (N_1502,N_594,N_338);
nand U1503 (N_1503,N_616,N_283);
nand U1504 (N_1504,N_529,N_1201);
nor U1505 (N_1505,N_662,N_1056);
or U1506 (N_1506,N_1466,N_812);
nand U1507 (N_1507,N_1002,N_996);
nor U1508 (N_1508,N_1165,N_1348);
or U1509 (N_1509,N_1055,N_1275);
nand U1510 (N_1510,N_598,N_526);
or U1511 (N_1511,N_916,N_319);
nand U1512 (N_1512,N_1232,N_637);
and U1513 (N_1513,N_344,N_314);
nand U1514 (N_1514,N_1279,N_560);
or U1515 (N_1515,N_824,N_122);
and U1516 (N_1516,N_337,N_72);
nor U1517 (N_1517,N_321,N_511);
nor U1518 (N_1518,N_373,N_818);
or U1519 (N_1519,N_1140,N_660);
xnor U1520 (N_1520,N_1099,N_172);
nor U1521 (N_1521,N_721,N_801);
nor U1522 (N_1522,N_472,N_1262);
or U1523 (N_1523,N_686,N_1346);
or U1524 (N_1524,N_775,N_836);
nand U1525 (N_1525,N_1032,N_254);
nand U1526 (N_1526,N_556,N_290);
xnor U1527 (N_1527,N_835,N_901);
nand U1528 (N_1528,N_1322,N_1085);
nand U1529 (N_1529,N_942,N_42);
or U1530 (N_1530,N_1033,N_1060);
xnor U1531 (N_1531,N_833,N_1254);
and U1532 (N_1532,N_800,N_1186);
and U1533 (N_1533,N_700,N_1481);
and U1534 (N_1534,N_706,N_96);
nand U1535 (N_1535,N_950,N_218);
or U1536 (N_1536,N_565,N_647);
or U1537 (N_1537,N_1013,N_555);
nor U1538 (N_1538,N_742,N_713);
xor U1539 (N_1539,N_1432,N_729);
and U1540 (N_1540,N_1461,N_878);
and U1541 (N_1541,N_1310,N_705);
and U1542 (N_1542,N_855,N_212);
and U1543 (N_1543,N_1106,N_1065);
or U1544 (N_1544,N_1390,N_1258);
and U1545 (N_1545,N_476,N_286);
nand U1546 (N_1546,N_1394,N_694);
and U1547 (N_1547,N_1082,N_368);
or U1548 (N_1548,N_315,N_217);
xor U1549 (N_1549,N_214,N_640);
and U1550 (N_1550,N_355,N_967);
xor U1551 (N_1551,N_1204,N_1272);
or U1552 (N_1552,N_57,N_1485);
and U1553 (N_1553,N_1286,N_1281);
nand U1554 (N_1554,N_264,N_175);
or U1555 (N_1555,N_304,N_443);
nand U1556 (N_1556,N_1453,N_1471);
nand U1557 (N_1557,N_843,N_573);
xor U1558 (N_1558,N_1087,N_1486);
xnor U1559 (N_1559,N_1494,N_965);
or U1560 (N_1560,N_612,N_1226);
or U1561 (N_1561,N_1045,N_890);
xor U1562 (N_1562,N_1396,N_200);
xor U1563 (N_1563,N_75,N_948);
and U1564 (N_1564,N_245,N_1230);
and U1565 (N_1565,N_743,N_1206);
xnor U1566 (N_1566,N_894,N_495);
or U1567 (N_1567,N_78,N_410);
xnor U1568 (N_1568,N_1323,N_572);
and U1569 (N_1569,N_1111,N_1324);
nand U1570 (N_1570,N_678,N_1264);
and U1571 (N_1571,N_649,N_1020);
nand U1572 (N_1572,N_617,N_1001);
or U1573 (N_1573,N_177,N_752);
or U1574 (N_1574,N_430,N_825);
nand U1575 (N_1575,N_1263,N_546);
nand U1576 (N_1576,N_575,N_188);
xnor U1577 (N_1577,N_1383,N_796);
or U1578 (N_1578,N_604,N_797);
nand U1579 (N_1579,N_334,N_385);
nor U1580 (N_1580,N_467,N_358);
nor U1581 (N_1581,N_263,N_990);
and U1582 (N_1582,N_514,N_1141);
nor U1583 (N_1583,N_167,N_1079);
xnor U1584 (N_1584,N_1340,N_416);
and U1585 (N_1585,N_317,N_105);
nand U1586 (N_1586,N_772,N_726);
and U1587 (N_1587,N_754,N_1381);
and U1588 (N_1588,N_858,N_777);
and U1589 (N_1589,N_943,N_1268);
xnor U1590 (N_1590,N_1078,N_95);
or U1591 (N_1591,N_829,N_359);
nand U1592 (N_1592,N_408,N_280);
nor U1593 (N_1593,N_932,N_866);
nor U1594 (N_1594,N_306,N_130);
and U1595 (N_1595,N_1156,N_310);
and U1596 (N_1596,N_930,N_251);
nand U1597 (N_1597,N_81,N_893);
xnor U1598 (N_1598,N_146,N_1473);
nor U1599 (N_1599,N_642,N_266);
nand U1600 (N_1600,N_515,N_82);
or U1601 (N_1601,N_924,N_1303);
and U1602 (N_1602,N_490,N_681);
or U1603 (N_1603,N_1255,N_684);
nand U1604 (N_1604,N_730,N_1212);
or U1605 (N_1605,N_1395,N_449);
nor U1606 (N_1606,N_1318,N_904);
nand U1607 (N_1607,N_345,N_1152);
nor U1608 (N_1608,N_1195,N_771);
nor U1609 (N_1609,N_891,N_453);
and U1610 (N_1610,N_428,N_540);
or U1611 (N_1611,N_494,N_623);
nor U1612 (N_1612,N_155,N_423);
nand U1613 (N_1613,N_1034,N_1122);
and U1614 (N_1614,N_44,N_1489);
or U1615 (N_1615,N_1153,N_1081);
nor U1616 (N_1616,N_570,N_1488);
or U1617 (N_1617,N_242,N_1339);
and U1618 (N_1618,N_614,N_21);
or U1619 (N_1619,N_504,N_823);
or U1620 (N_1620,N_1170,N_216);
nor U1621 (N_1621,N_1454,N_1313);
nor U1622 (N_1622,N_939,N_1353);
nor U1623 (N_1623,N_848,N_402);
and U1624 (N_1624,N_267,N_1220);
or U1625 (N_1625,N_1372,N_1108);
xnor U1626 (N_1626,N_790,N_320);
nor U1627 (N_1627,N_275,N_1282);
or U1628 (N_1628,N_1160,N_298);
nor U1629 (N_1629,N_277,N_1316);
and U1630 (N_1630,N_1084,N_946);
and U1631 (N_1631,N_1387,N_922);
nand U1632 (N_1632,N_1445,N_295);
and U1633 (N_1633,N_139,N_362);
nor U1634 (N_1634,N_941,N_1197);
nor U1635 (N_1635,N_676,N_1465);
and U1636 (N_1636,N_659,N_211);
and U1637 (N_1637,N_19,N_170);
nor U1638 (N_1638,N_725,N_1245);
nor U1639 (N_1639,N_438,N_346);
nand U1640 (N_1640,N_508,N_350);
nor U1641 (N_1641,N_774,N_1223);
or U1642 (N_1642,N_884,N_783);
nor U1643 (N_1643,N_1051,N_349);
nor U1644 (N_1644,N_1405,N_963);
or U1645 (N_1645,N_1467,N_1115);
and U1646 (N_1646,N_339,N_651);
nor U1647 (N_1647,N_849,N_1437);
nor U1648 (N_1648,N_1351,N_231);
and U1649 (N_1649,N_925,N_497);
nand U1650 (N_1650,N_528,N_577);
nand U1651 (N_1651,N_693,N_195);
and U1652 (N_1652,N_1447,N_1196);
or U1653 (N_1653,N_1419,N_1208);
or U1654 (N_1654,N_1180,N_1274);
xnor U1655 (N_1655,N_1040,N_284);
nand U1656 (N_1656,N_867,N_1298);
xor U1657 (N_1657,N_74,N_1378);
and U1658 (N_1658,N_962,N_837);
nor U1659 (N_1659,N_1007,N_786);
nor U1660 (N_1660,N_1219,N_1278);
nand U1661 (N_1661,N_988,N_1128);
and U1662 (N_1662,N_697,N_782);
and U1663 (N_1663,N_805,N_767);
or U1664 (N_1664,N_670,N_1482);
nor U1665 (N_1665,N_192,N_955);
nor U1666 (N_1666,N_677,N_199);
and U1667 (N_1667,N_50,N_535);
nor U1668 (N_1668,N_150,N_76);
xor U1669 (N_1669,N_1433,N_1028);
and U1670 (N_1670,N_287,N_137);
nand U1671 (N_1671,N_45,N_952);
and U1672 (N_1672,N_183,N_1308);
or U1673 (N_1673,N_1116,N_673);
and U1674 (N_1674,N_959,N_491);
nand U1675 (N_1675,N_1253,N_247);
nor U1676 (N_1676,N_1217,N_1431);
nor U1677 (N_1677,N_1071,N_1413);
and U1678 (N_1678,N_583,N_1290);
or U1679 (N_1679,N_225,N_525);
or U1680 (N_1680,N_854,N_1006);
nand U1681 (N_1681,N_1301,N_845);
nor U1682 (N_1682,N_1090,N_638);
or U1683 (N_1683,N_709,N_722);
nand U1684 (N_1684,N_166,N_731);
and U1685 (N_1685,N_973,N_1487);
and U1686 (N_1686,N_1236,N_778);
and U1687 (N_1687,N_1450,N_120);
or U1688 (N_1688,N_872,N_109);
or U1689 (N_1689,N_784,N_118);
and U1690 (N_1690,N_201,N_1434);
nand U1691 (N_1691,N_2,N_204);
or U1692 (N_1692,N_426,N_324);
nor U1693 (N_1693,N_701,N_1293);
or U1694 (N_1694,N_607,N_375);
and U1695 (N_1695,N_79,N_844);
and U1696 (N_1696,N_509,N_1270);
nor U1697 (N_1697,N_444,N_483);
nor U1698 (N_1698,N_559,N_1100);
or U1699 (N_1699,N_1297,N_1259);
xor U1700 (N_1700,N_853,N_1261);
or U1701 (N_1701,N_910,N_422);
or U1702 (N_1702,N_834,N_36);
xor U1703 (N_1703,N_1004,N_1070);
nand U1704 (N_1704,N_873,N_597);
or U1705 (N_1705,N_223,N_564);
and U1706 (N_1706,N_458,N_1092);
nand U1707 (N_1707,N_31,N_1172);
and U1708 (N_1708,N_586,N_1185);
and U1709 (N_1709,N_117,N_1247);
and U1710 (N_1710,N_751,N_1047);
or U1711 (N_1711,N_1101,N_1412);
or U1712 (N_1712,N_1144,N_921);
or U1713 (N_1713,N_152,N_568);
or U1714 (N_1714,N_1161,N_919);
nand U1715 (N_1715,N_505,N_1408);
nor U1716 (N_1716,N_1414,N_808);
nor U1717 (N_1717,N_271,N_209);
nor U1718 (N_1718,N_1222,N_1011);
nor U1719 (N_1719,N_1302,N_758);
nor U1720 (N_1720,N_1191,N_579);
xnor U1721 (N_1721,N_1399,N_482);
and U1722 (N_1722,N_1072,N_1010);
or U1723 (N_1723,N_1138,N_156);
or U1724 (N_1724,N_1363,N_456);
nand U1725 (N_1725,N_1416,N_196);
or U1726 (N_1726,N_1448,N_62);
xor U1727 (N_1727,N_915,N_64);
nand U1728 (N_1728,N_1117,N_895);
nand U1729 (N_1729,N_1231,N_104);
and U1730 (N_1730,N_813,N_562);
and U1731 (N_1731,N_1252,N_715);
nand U1732 (N_1732,N_633,N_87);
nor U1733 (N_1733,N_857,N_518);
or U1734 (N_1734,N_7,N_738);
nand U1735 (N_1735,N_803,N_70);
or U1736 (N_1736,N_432,N_99);
nor U1737 (N_1737,N_1088,N_1131);
xnor U1738 (N_1738,N_143,N_427);
nand U1739 (N_1739,N_1151,N_1015);
or U1740 (N_1740,N_322,N_182);
and U1741 (N_1741,N_1333,N_1306);
or U1742 (N_1742,N_61,N_1075);
nor U1743 (N_1743,N_1480,N_1407);
nor U1744 (N_1744,N_1440,N_762);
xor U1745 (N_1745,N_740,N_1022);
or U1746 (N_1746,N_881,N_1130);
or U1747 (N_1747,N_1364,N_328);
or U1748 (N_1748,N_58,N_8);
or U1749 (N_1749,N_148,N_365);
or U1750 (N_1750,N_142,N_420);
xor U1751 (N_1751,N_896,N_439);
and U1752 (N_1752,N_1190,N_871);
nor U1753 (N_1753,N_789,N_107);
nand U1754 (N_1754,N_958,N_934);
and U1755 (N_1755,N_114,N_794);
or U1756 (N_1756,N_1441,N_613);
or U1757 (N_1757,N_73,N_682);
and U1758 (N_1758,N_821,N_144);
nor U1759 (N_1759,N_374,N_12);
nand U1760 (N_1760,N_892,N_976);
or U1761 (N_1761,N_553,N_161);
or U1762 (N_1762,N_1164,N_1112);
nand U1763 (N_1763,N_499,N_29);
or U1764 (N_1764,N_1429,N_542);
xnor U1765 (N_1765,N_944,N_862);
or U1766 (N_1766,N_369,N_780);
nand U1767 (N_1767,N_138,N_773);
or U1768 (N_1768,N_691,N_634);
nand U1769 (N_1769,N_303,N_657);
and U1770 (N_1770,N_451,N_1127);
nor U1771 (N_1771,N_1183,N_1325);
xnor U1772 (N_1772,N_1398,N_352);
and U1773 (N_1773,N_1367,N_1273);
nor U1774 (N_1774,N_289,N_1402);
and U1775 (N_1775,N_814,N_1370);
nand U1776 (N_1776,N_1053,N_668);
nor U1777 (N_1777,N_331,N_1426);
or U1778 (N_1778,N_1406,N_437);
nor U1779 (N_1779,N_1446,N_918);
and U1780 (N_1780,N_1037,N_851);
and U1781 (N_1781,N_816,N_995);
nand U1782 (N_1782,N_1352,N_679);
and U1783 (N_1783,N_886,N_1228);
nand U1784 (N_1784,N_1076,N_127);
or U1785 (N_1785,N_533,N_645);
and U1786 (N_1786,N_1491,N_1299);
nor U1787 (N_1787,N_238,N_933);
or U1788 (N_1788,N_1241,N_1200);
and U1789 (N_1789,N_15,N_488);
or U1790 (N_1790,N_340,N_37);
or U1791 (N_1791,N_766,N_411);
and U1792 (N_1792,N_753,N_1);
and U1793 (N_1793,N_876,N_404);
nand U1794 (N_1794,N_1355,N_86);
and U1795 (N_1795,N_71,N_1000);
and U1796 (N_1796,N_1411,N_474);
nor U1797 (N_1797,N_1493,N_1309);
and U1798 (N_1798,N_1018,N_342);
xor U1799 (N_1799,N_1120,N_938);
and U1800 (N_1800,N_608,N_442);
nor U1801 (N_1801,N_228,N_1158);
and U1802 (N_1802,N_1058,N_785);
nor U1803 (N_1803,N_471,N_710);
and U1804 (N_1804,N_1104,N_388);
nand U1805 (N_1805,N_403,N_101);
nand U1806 (N_1806,N_123,N_975);
and U1807 (N_1807,N_1119,N_69);
nand U1808 (N_1808,N_1063,N_171);
nor U1809 (N_1809,N_448,N_235);
and U1810 (N_1810,N_477,N_220);
or U1811 (N_1811,N_1427,N_966);
nor U1812 (N_1812,N_1234,N_91);
and U1813 (N_1813,N_675,N_989);
and U1814 (N_1814,N_1029,N_190);
and U1815 (N_1815,N_549,N_256);
nor U1816 (N_1816,N_629,N_174);
and U1817 (N_1817,N_1187,N_436);
or U1818 (N_1818,N_1499,N_1495);
or U1819 (N_1819,N_1175,N_193);
and U1820 (N_1820,N_1118,N_1036);
and U1821 (N_1821,N_1094,N_191);
and U1822 (N_1822,N_548,N_1269);
nand U1823 (N_1823,N_595,N_305);
xnor U1824 (N_1824,N_378,N_103);
nand U1825 (N_1825,N_18,N_1404);
and U1826 (N_1826,N_689,N_429);
or U1827 (N_1827,N_1146,N_1061);
nand U1828 (N_1828,N_249,N_1443);
nor U1829 (N_1829,N_1062,N_1350);
or U1830 (N_1830,N_665,N_750);
or U1831 (N_1831,N_1041,N_1424);
or U1832 (N_1832,N_1439,N_899);
or U1833 (N_1833,N_819,N_563);
nor U1834 (N_1834,N_282,N_1246);
and U1835 (N_1835,N_1296,N_698);
and U1836 (N_1836,N_111,N_405);
or U1837 (N_1837,N_1113,N_11);
or U1838 (N_1838,N_759,N_291);
and U1839 (N_1839,N_1114,N_643);
nand U1840 (N_1840,N_1124,N_1421);
nand U1841 (N_1841,N_1218,N_23);
or U1842 (N_1842,N_961,N_68);
or U1843 (N_1843,N_1251,N_43);
nor U1844 (N_1844,N_396,N_52);
nand U1845 (N_1845,N_1295,N_671);
nand U1846 (N_1846,N_492,N_386);
nor U1847 (N_1847,N_53,N_512);
xnor U1848 (N_1848,N_360,N_661);
nand U1849 (N_1849,N_401,N_6);
and U1850 (N_1850,N_792,N_547);
or U1851 (N_1851,N_1143,N_1451);
nand U1852 (N_1852,N_557,N_397);
nand U1853 (N_1853,N_1288,N_720);
and U1854 (N_1854,N_116,N_981);
nor U1855 (N_1855,N_464,N_1096);
nand U1856 (N_1856,N_1256,N_917);
or U1857 (N_1857,N_89,N_1182);
and U1858 (N_1858,N_185,N_817);
or U1859 (N_1859,N_1225,N_567);
nand U1860 (N_1860,N_839,N_1319);
and U1861 (N_1861,N_911,N_566);
nor U1862 (N_1862,N_1052,N_316);
nand U1863 (N_1863,N_503,N_1046);
and U1864 (N_1864,N_1452,N_1360);
or U1865 (N_1865,N_389,N_311);
xor U1866 (N_1866,N_473,N_905);
and U1867 (N_1867,N_520,N_498);
and U1868 (N_1868,N_978,N_259);
and U1869 (N_1869,N_115,N_92);
and U1870 (N_1870,N_791,N_581);
nor U1871 (N_1871,N_452,N_1189);
and U1872 (N_1872,N_273,N_1386);
and U1873 (N_1873,N_584,N_1227);
and U1874 (N_1874,N_732,N_639);
nor U1875 (N_1875,N_1362,N_887);
nor U1876 (N_1876,N_1326,N_606);
nand U1877 (N_1877,N_1455,N_164);
nand U1878 (N_1878,N_846,N_827);
and U1879 (N_1879,N_1460,N_1205);
xor U1880 (N_1880,N_500,N_1089);
and U1881 (N_1881,N_409,N_860);
nor U1882 (N_1882,N_733,N_804);
nand U1883 (N_1883,N_487,N_244);
xnor U1884 (N_1884,N_151,N_1312);
nand U1885 (N_1885,N_433,N_840);
nand U1886 (N_1886,N_1043,N_1265);
nand U1887 (N_1887,N_224,N_688);
or U1888 (N_1888,N_1458,N_243);
nor U1889 (N_1889,N_1147,N_1250);
xnor U1890 (N_1890,N_173,N_920);
and U1891 (N_1891,N_672,N_1385);
or U1892 (N_1892,N_864,N_1202);
nand U1893 (N_1893,N_269,N_1024);
xnor U1894 (N_1894,N_1345,N_696);
and U1895 (N_1895,N_744,N_763);
nor U1896 (N_1896,N_1162,N_644);
nor U1897 (N_1897,N_1401,N_593);
nand U1898 (N_1898,N_1289,N_1430);
and U1899 (N_1899,N_234,N_1005);
or U1900 (N_1900,N_431,N_1472);
nor U1901 (N_1901,N_1462,N_147);
and U1902 (N_1902,N_382,N_1159);
and U1903 (N_1903,N_268,N_624);
or U1904 (N_1904,N_1347,N_1484);
or U1905 (N_1905,N_582,N_1442);
nand U1906 (N_1906,N_1285,N_1335);
or U1907 (N_1907,N_1016,N_1283);
nor U1908 (N_1908,N_717,N_213);
and U1909 (N_1909,N_983,N_711);
nand U1910 (N_1910,N_974,N_468);
or U1911 (N_1911,N_312,N_850);
or U1912 (N_1912,N_313,N_968);
or U1913 (N_1913,N_93,N_1490);
nor U1914 (N_1914,N_699,N_591);
xnor U1915 (N_1915,N_1026,N_538);
xor U1916 (N_1916,N_108,N_141);
nand U1917 (N_1917,N_366,N_658);
and U1918 (N_1918,N_596,N_882);
or U1919 (N_1919,N_718,N_727);
nor U1920 (N_1920,N_1169,N_66);
or U1921 (N_1921,N_907,N_463);
and U1922 (N_1922,N_361,N_372);
or U1923 (N_1923,N_145,N_793);
nor U1924 (N_1924,N_38,N_507);
or U1925 (N_1925,N_10,N_250);
and U1926 (N_1926,N_776,N_457);
or U1927 (N_1927,N_685,N_626);
nand U1928 (N_1928,N_1224,N_1209);
nand U1929 (N_1929,N_1136,N_735);
nand U1930 (N_1930,N_49,N_1049);
nand U1931 (N_1931,N_666,N_537);
or U1932 (N_1932,N_809,N_1365);
xnor U1933 (N_1933,N_460,N_765);
or U1934 (N_1934,N_993,N_466);
nor U1935 (N_1935,N_383,N_1388);
nor U1936 (N_1936,N_134,N_1199);
nand U1937 (N_1937,N_1376,N_252);
and U1938 (N_1938,N_294,N_325);
xnor U1939 (N_1939,N_1179,N_605);
and U1940 (N_1940,N_625,N_908);
and U1941 (N_1941,N_1157,N_59);
nand U1942 (N_1942,N_601,N_847);
nor U1943 (N_1943,N_859,N_736);
nor U1944 (N_1944,N_739,N_600);
nor U1945 (N_1945,N_187,N_986);
or U1946 (N_1946,N_326,N_832);
and U1947 (N_1947,N_1012,N_580);
or U1948 (N_1948,N_157,N_257);
and U1949 (N_1949,N_1330,N_335);
nand U1950 (N_1950,N_648,N_1331);
nor U1951 (N_1951,N_768,N_395);
nand U1952 (N_1952,N_926,N_1054);
nor U1953 (N_1953,N_1456,N_179);
nor U1954 (N_1954,N_723,N_205);
nor U1955 (N_1955,N_1139,N_802);
or U1956 (N_1956,N_1039,N_1329);
nand U1957 (N_1957,N_1221,N_1133);
nor U1958 (N_1958,N_336,N_88);
nor U1959 (N_1959,N_1057,N_1300);
or U1960 (N_1960,N_1328,N_1242);
and U1961 (N_1961,N_1135,N_189);
and U1962 (N_1962,N_576,N_1359);
and U1963 (N_1963,N_197,N_1248);
nor U1964 (N_1964,N_1358,N_879);
nor U1965 (N_1965,N_747,N_991);
or U1966 (N_1966,N_1377,N_332);
and U1967 (N_1967,N_712,N_496);
or U1968 (N_1968,N_830,N_16);
and U1969 (N_1969,N_100,N_1249);
nor U1970 (N_1970,N_128,N_1304);
and U1971 (N_1971,N_80,N_27);
nand U1972 (N_1972,N_384,N_714);
xnor U1973 (N_1973,N_516,N_25);
xor U1974 (N_1974,N_347,N_329);
nand U1975 (N_1975,N_1174,N_1468);
nand U1976 (N_1976,N_441,N_541);
nand U1977 (N_1977,N_1110,N_24);
nor U1978 (N_1978,N_1149,N_1371);
nor U1979 (N_1979,N_9,N_1163);
nor U1980 (N_1980,N_532,N_1192);
xnor U1981 (N_1981,N_501,N_1380);
nor U1982 (N_1982,N_30,N_154);
nand U1983 (N_1983,N_1497,N_883);
nor U1984 (N_1984,N_861,N_880);
and U1985 (N_1985,N_354,N_716);
or U1986 (N_1986,N_987,N_126);
and U1987 (N_1987,N_928,N_272);
nand U1988 (N_1988,N_279,N_1176);
and U1989 (N_1989,N_465,N_695);
and U1990 (N_1990,N_106,N_176);
nand U1991 (N_1991,N_877,N_1074);
or U1992 (N_1992,N_357,N_1344);
nor U1993 (N_1993,N_323,N_1315);
and U1994 (N_1994,N_206,N_455);
and U1995 (N_1995,N_274,N_1470);
xor U1996 (N_1996,N_947,N_574);
and U1997 (N_1997,N_348,N_125);
nor U1998 (N_1998,N_28,N_781);
nor U1999 (N_1999,N_1167,N_446);
nand U2000 (N_2000,N_353,N_940);
xnor U2001 (N_2001,N_534,N_1280);
or U2002 (N_2002,N_1420,N_419);
nor U2003 (N_2003,N_615,N_215);
or U2004 (N_2004,N_1321,N_390);
and U2005 (N_2005,N_129,N_1392);
or U2006 (N_2006,N_770,N_680);
and U2007 (N_2007,N_953,N_1103);
xor U2008 (N_2008,N_1177,N_470);
xnor U2009 (N_2009,N_1031,N_1211);
nand U2010 (N_2010,N_255,N_1477);
nand U2011 (N_2011,N_1444,N_168);
xor U2012 (N_2012,N_119,N_539);
or U2013 (N_2013,N_3,N_302);
or U2014 (N_2014,N_363,N_1354);
or U2015 (N_2015,N_1469,N_755);
nand U2016 (N_2016,N_379,N_960);
and U2017 (N_2017,N_262,N_764);
and U2018 (N_2018,N_459,N_392);
nor U2019 (N_2019,N_90,N_1498);
nand U2020 (N_2020,N_703,N_1327);
or U2021 (N_2021,N_798,N_391);
and U2022 (N_2022,N_517,N_788);
xor U2023 (N_2023,N_1240,N_1207);
nor U2024 (N_2024,N_1154,N_631);
and U2025 (N_2025,N_1203,N_519);
or U2026 (N_2026,N_531,N_728);
nand U2027 (N_2027,N_1093,N_870);
nand U2028 (N_2028,N_169,N_544);
nor U2029 (N_2029,N_1069,N_203);
or U2030 (N_2030,N_622,N_1171);
nand U2031 (N_2031,N_994,N_652);
and U2032 (N_2032,N_708,N_40);
nor U2033 (N_2033,N_110,N_1068);
nand U2034 (N_2034,N_863,N_377);
or U2035 (N_2035,N_1073,N_856);
nand U2036 (N_2036,N_779,N_1320);
nand U2037 (N_2037,N_674,N_121);
nor U2038 (N_2038,N_1107,N_653);
nand U2039 (N_2039,N_248,N_1042);
or U2040 (N_2040,N_1260,N_424);
and U2041 (N_2041,N_669,N_979);
xor U2042 (N_2042,N_707,N_1244);
or U2043 (N_2043,N_239,N_654);
xor U2044 (N_2044,N_875,N_84);
nor U2045 (N_2045,N_56,N_1166);
nor U2046 (N_2046,N_510,N_1391);
nand U2047 (N_2047,N_656,N_1243);
or U2048 (N_2048,N_413,N_258);
nor U2049 (N_2049,N_667,N_5);
and U2050 (N_2050,N_1409,N_999);
nor U2051 (N_2051,N_1287,N_435);
and U2052 (N_2052,N_39,N_636);
nor U2053 (N_2053,N_1438,N_936);
or U2054 (N_2054,N_461,N_55);
xnor U2055 (N_2055,N_1237,N_1317);
and U2056 (N_2056,N_184,N_646);
nor U2057 (N_2057,N_1483,N_4);
and U2058 (N_2058,N_14,N_132);
or U2059 (N_2059,N_1479,N_1213);
and U2060 (N_2060,N_34,N_977);
nand U2061 (N_2061,N_1428,N_888);
nand U2062 (N_2062,N_97,N_1334);
or U2063 (N_2063,N_1457,N_480);
and U2064 (N_2064,N_971,N_1129);
nor U2065 (N_2065,N_489,N_1435);
nand U2066 (N_2066,N_20,N_1474);
and U2067 (N_2067,N_1023,N_587);
and U2068 (N_2068,N_561,N_984);
xnor U2069 (N_2069,N_1038,N_48);
nand U2070 (N_2070,N_807,N_1083);
or U2071 (N_2071,N_1035,N_425);
or U2072 (N_2072,N_1266,N_588);
nor U2073 (N_2073,N_434,N_370);
nand U2074 (N_2074,N_202,N_909);
xnor U2075 (N_2075,N_1403,N_1375);
and U2076 (N_2076,N_297,N_1009);
and U2077 (N_2077,N_620,N_1305);
nand U2078 (N_2078,N_0,N_970);
or U2079 (N_2079,N_94,N_702);
or U2080 (N_2080,N_140,N_440);
nor U2081 (N_2081,N_1137,N_1233);
nand U2082 (N_2082,N_178,N_1337);
nor U2083 (N_2083,N_1008,N_136);
nor U2084 (N_2084,N_951,N_1193);
nand U2085 (N_2085,N_1475,N_506);
nor U2086 (N_2086,N_293,N_219);
nand U2087 (N_2087,N_618,N_153);
and U2088 (N_2088,N_1423,N_51);
nor U2089 (N_2089,N_1369,N_913);
nor U2090 (N_2090,N_609,N_1239);
and U2091 (N_2091,N_1019,N_318);
nand U2092 (N_2092,N_207,N_635);
nand U2093 (N_2093,N_1188,N_1086);
nor U2094 (N_2094,N_400,N_690);
xnor U2095 (N_2095,N_589,N_479);
xnor U2096 (N_2096,N_113,N_1336);
and U2097 (N_2097,N_931,N_1374);
and U2098 (N_2098,N_54,N_485);
or U2099 (N_2099,N_112,N_1194);
and U2100 (N_2100,N_769,N_1050);
and U2101 (N_2101,N_356,N_719);
nor U2102 (N_2102,N_929,N_462);
nand U2103 (N_2103,N_1235,N_683);
and U2104 (N_2104,N_945,N_927);
or U2105 (N_2105,N_22,N_826);
and U2106 (N_2106,N_554,N_1098);
or U2107 (N_2107,N_956,N_1397);
nand U2108 (N_2108,N_610,N_1292);
nor U2109 (N_2109,N_17,N_787);
and U2110 (N_2110,N_745,N_1030);
and U2111 (N_2111,N_1257,N_26);
or U2112 (N_2112,N_949,N_1021);
or U2113 (N_2113,N_527,N_276);
nand U2114 (N_2114,N_380,N_475);
or U2115 (N_2115,N_229,N_222);
and U2116 (N_2116,N_889,N_165);
and U2117 (N_2117,N_902,N_181);
nor U2118 (N_2118,N_417,N_445);
nor U2119 (N_2119,N_1436,N_1181);
and U2120 (N_2120,N_906,N_367);
xor U2121 (N_2121,N_757,N_1389);
nor U2122 (N_2122,N_1095,N_992);
and U2123 (N_2123,N_63,N_221);
or U2124 (N_2124,N_398,N_868);
and U2125 (N_2125,N_296,N_885);
nand U2126 (N_2126,N_32,N_1342);
nand U2127 (N_2127,N_550,N_964);
and U2128 (N_2128,N_603,N_1307);
or U2129 (N_2129,N_865,N_664);
nand U2130 (N_2130,N_13,N_233);
and U2131 (N_2131,N_545,N_1215);
and U2132 (N_2132,N_133,N_1121);
nand U2133 (N_2133,N_569,N_822);
nand U2134 (N_2134,N_1361,N_1459);
nand U2135 (N_2135,N_261,N_237);
or U2136 (N_2136,N_741,N_687);
nand U2137 (N_2137,N_102,N_486);
xor U2138 (N_2138,N_1417,N_874);
nor U2139 (N_2139,N_1425,N_611);
and U2140 (N_2140,N_1238,N_415);
nand U2141 (N_2141,N_543,N_281);
nand U2142 (N_2142,N_1368,N_1415);
or U2143 (N_2143,N_815,N_208);
or U2144 (N_2144,N_418,N_65);
nand U2145 (N_2145,N_1464,N_1148);
or U2146 (N_2146,N_799,N_1145);
and U2147 (N_2147,N_226,N_1332);
nor U2148 (N_2148,N_746,N_236);
and U2149 (N_2149,N_160,N_998);
and U2150 (N_2150,N_869,N_513);
or U2151 (N_2151,N_578,N_969);
and U2152 (N_2152,N_641,N_1059);
and U2153 (N_2153,N_1066,N_180);
or U2154 (N_2154,N_47,N_571);
nand U2155 (N_2155,N_1357,N_1003);
nor U2156 (N_2156,N_903,N_1294);
xnor U2157 (N_2157,N_1382,N_230);
or U2158 (N_2158,N_343,N_820);
or U2159 (N_2159,N_1343,N_241);
nor U2160 (N_2160,N_914,N_1027);
nand U2161 (N_2161,N_831,N_1184);
nor U2162 (N_2162,N_1410,N_1338);
xnor U2163 (N_2163,N_186,N_599);
nor U2164 (N_2164,N_1025,N_1476);
xor U2165 (N_2165,N_761,N_270);
or U2166 (N_2166,N_1102,N_1198);
nand U2167 (N_2167,N_1216,N_523);
xor U2168 (N_2168,N_1064,N_810);
xor U2169 (N_2169,N_1373,N_621);
nor U2170 (N_2170,N_997,N_1311);
xnor U2171 (N_2171,N_1048,N_811);
nor U2172 (N_2172,N_85,N_1356);
and U2173 (N_2173,N_590,N_67);
nand U2174 (N_2174,N_900,N_937);
and U2175 (N_2175,N_734,N_1091);
nand U2176 (N_2176,N_227,N_619);
or U2177 (N_2177,N_912,N_1463);
or U2178 (N_2178,N_806,N_655);
nor U2179 (N_2179,N_1276,N_524);
or U2180 (N_2180,N_285,N_83);
xnor U2181 (N_2181,N_1168,N_330);
or U2182 (N_2182,N_795,N_841);
nor U2183 (N_2183,N_162,N_954);
nand U2184 (N_2184,N_1379,N_1214);
nor U2185 (N_2185,N_935,N_159);
nand U2186 (N_2186,N_35,N_387);
or U2187 (N_2187,N_46,N_828);
and U2188 (N_2188,N_447,N_450);
nor U2189 (N_2189,N_1155,N_957);
or U2190 (N_2190,N_972,N_163);
nor U2191 (N_2191,N_756,N_898);
or U2192 (N_2192,N_1271,N_530);
nor U2193 (N_2193,N_265,N_246);
or U2194 (N_2194,N_1126,N_1349);
nand U2195 (N_2195,N_381,N_1067);
nor U2196 (N_2196,N_838,N_1422);
xor U2197 (N_2197,N_737,N_478);
and U2198 (N_2198,N_484,N_1277);
and U2199 (N_2199,N_33,N_982);
nand U2200 (N_2200,N_985,N_469);
and U2201 (N_2201,N_1284,N_632);
xor U2202 (N_2202,N_124,N_1173);
nor U2203 (N_2203,N_394,N_481);
nand U2204 (N_2204,N_1109,N_1492);
nor U2205 (N_2205,N_650,N_253);
or U2206 (N_2206,N_1142,N_60);
and U2207 (N_2207,N_502,N_292);
nor U2208 (N_2208,N_376,N_558);
xnor U2209 (N_2209,N_1314,N_1105);
or U2210 (N_2210,N_407,N_1341);
nor U2211 (N_2211,N_149,N_307);
and U2212 (N_2212,N_663,N_628);
and U2213 (N_2213,N_748,N_692);
and U2214 (N_2214,N_1123,N_1014);
nor U2215 (N_2215,N_897,N_585);
nand U2216 (N_2216,N_412,N_210);
nor U2217 (N_2217,N_602,N_1150);
nand U2218 (N_2218,N_1077,N_630);
and U2219 (N_2219,N_521,N_301);
nor U2220 (N_2220,N_98,N_198);
and U2221 (N_2221,N_1134,N_1210);
nand U2222 (N_2222,N_592,N_327);
nand U2223 (N_2223,N_1496,N_923);
xor U2224 (N_2224,N_1132,N_454);
and U2225 (N_2225,N_749,N_493);
or U2226 (N_2226,N_77,N_1291);
xor U2227 (N_2227,N_980,N_399);
and U2228 (N_2228,N_1017,N_364);
and U2229 (N_2229,N_1080,N_724);
nand U2230 (N_2230,N_522,N_552);
or U2231 (N_2231,N_299,N_1366);
nor U2232 (N_2232,N_308,N_135);
and U2233 (N_2233,N_1097,N_341);
and U2234 (N_2234,N_627,N_158);
and U2235 (N_2235,N_421,N_1449);
nor U2236 (N_2236,N_1267,N_1178);
or U2237 (N_2237,N_309,N_278);
or U2238 (N_2238,N_414,N_300);
and U2239 (N_2239,N_406,N_240);
nand U2240 (N_2240,N_536,N_1418);
and U2241 (N_2241,N_333,N_288);
nand U2242 (N_2242,N_1229,N_194);
and U2243 (N_2243,N_760,N_371);
or U2244 (N_2244,N_1478,N_852);
xnor U2245 (N_2245,N_260,N_1125);
nand U2246 (N_2246,N_551,N_41);
and U2247 (N_2247,N_1044,N_1384);
and U2248 (N_2248,N_351,N_232);
nand U2249 (N_2249,N_704,N_1400);
or U2250 (N_2250,N_1119,N_655);
nand U2251 (N_2251,N_386,N_61);
xnor U2252 (N_2252,N_623,N_205);
nor U2253 (N_2253,N_531,N_650);
nor U2254 (N_2254,N_27,N_763);
and U2255 (N_2255,N_98,N_329);
and U2256 (N_2256,N_244,N_1213);
xnor U2257 (N_2257,N_182,N_143);
nor U2258 (N_2258,N_447,N_656);
nor U2259 (N_2259,N_1425,N_131);
and U2260 (N_2260,N_686,N_1345);
xnor U2261 (N_2261,N_1190,N_544);
and U2262 (N_2262,N_481,N_889);
nor U2263 (N_2263,N_584,N_1237);
xnor U2264 (N_2264,N_923,N_1305);
nand U2265 (N_2265,N_20,N_209);
or U2266 (N_2266,N_1109,N_772);
and U2267 (N_2267,N_338,N_1090);
and U2268 (N_2268,N_83,N_161);
nor U2269 (N_2269,N_400,N_1421);
and U2270 (N_2270,N_829,N_577);
nand U2271 (N_2271,N_393,N_899);
and U2272 (N_2272,N_301,N_641);
nand U2273 (N_2273,N_1123,N_907);
or U2274 (N_2274,N_1499,N_550);
and U2275 (N_2275,N_1092,N_65);
or U2276 (N_2276,N_785,N_1310);
or U2277 (N_2277,N_425,N_325);
or U2278 (N_2278,N_521,N_386);
nor U2279 (N_2279,N_561,N_30);
and U2280 (N_2280,N_782,N_662);
and U2281 (N_2281,N_906,N_1364);
nand U2282 (N_2282,N_1341,N_186);
nand U2283 (N_2283,N_1439,N_475);
or U2284 (N_2284,N_1246,N_666);
nor U2285 (N_2285,N_858,N_456);
nor U2286 (N_2286,N_1478,N_213);
and U2287 (N_2287,N_290,N_115);
or U2288 (N_2288,N_809,N_397);
nor U2289 (N_2289,N_64,N_344);
nand U2290 (N_2290,N_50,N_1032);
nor U2291 (N_2291,N_62,N_200);
nand U2292 (N_2292,N_216,N_903);
and U2293 (N_2293,N_492,N_764);
nor U2294 (N_2294,N_1367,N_386);
and U2295 (N_2295,N_696,N_1143);
nand U2296 (N_2296,N_492,N_1235);
and U2297 (N_2297,N_667,N_1298);
nand U2298 (N_2298,N_520,N_64);
nor U2299 (N_2299,N_437,N_794);
and U2300 (N_2300,N_457,N_315);
nor U2301 (N_2301,N_311,N_11);
nand U2302 (N_2302,N_465,N_8);
and U2303 (N_2303,N_110,N_581);
nand U2304 (N_2304,N_428,N_594);
or U2305 (N_2305,N_745,N_290);
nor U2306 (N_2306,N_716,N_527);
xnor U2307 (N_2307,N_964,N_250);
nor U2308 (N_2308,N_1397,N_1427);
or U2309 (N_2309,N_418,N_1464);
nor U2310 (N_2310,N_303,N_1274);
nand U2311 (N_2311,N_716,N_38);
and U2312 (N_2312,N_126,N_366);
or U2313 (N_2313,N_1448,N_662);
or U2314 (N_2314,N_8,N_112);
and U2315 (N_2315,N_7,N_1406);
nand U2316 (N_2316,N_756,N_873);
and U2317 (N_2317,N_559,N_999);
and U2318 (N_2318,N_1235,N_599);
and U2319 (N_2319,N_1283,N_724);
nor U2320 (N_2320,N_687,N_1133);
nor U2321 (N_2321,N_286,N_1162);
xor U2322 (N_2322,N_40,N_918);
nand U2323 (N_2323,N_16,N_159);
and U2324 (N_2324,N_1474,N_1106);
or U2325 (N_2325,N_1001,N_1360);
nor U2326 (N_2326,N_1455,N_907);
nand U2327 (N_2327,N_935,N_1114);
xor U2328 (N_2328,N_328,N_312);
and U2329 (N_2329,N_67,N_766);
xor U2330 (N_2330,N_1085,N_186);
or U2331 (N_2331,N_951,N_813);
nor U2332 (N_2332,N_1021,N_338);
or U2333 (N_2333,N_1241,N_1289);
nand U2334 (N_2334,N_1458,N_1482);
nand U2335 (N_2335,N_1219,N_44);
or U2336 (N_2336,N_972,N_1070);
or U2337 (N_2337,N_1080,N_745);
and U2338 (N_2338,N_1348,N_679);
and U2339 (N_2339,N_1013,N_840);
xnor U2340 (N_2340,N_550,N_611);
or U2341 (N_2341,N_1041,N_273);
nor U2342 (N_2342,N_867,N_1248);
nor U2343 (N_2343,N_1153,N_746);
or U2344 (N_2344,N_1488,N_417);
nor U2345 (N_2345,N_1126,N_925);
and U2346 (N_2346,N_724,N_1378);
and U2347 (N_2347,N_996,N_686);
or U2348 (N_2348,N_361,N_251);
nor U2349 (N_2349,N_1425,N_1163);
nand U2350 (N_2350,N_404,N_1154);
nand U2351 (N_2351,N_623,N_550);
nor U2352 (N_2352,N_534,N_65);
and U2353 (N_2353,N_101,N_620);
nor U2354 (N_2354,N_643,N_1198);
and U2355 (N_2355,N_106,N_1360);
xnor U2356 (N_2356,N_377,N_90);
or U2357 (N_2357,N_454,N_772);
xnor U2358 (N_2358,N_742,N_1319);
and U2359 (N_2359,N_895,N_133);
or U2360 (N_2360,N_76,N_642);
or U2361 (N_2361,N_1097,N_944);
nor U2362 (N_2362,N_531,N_1431);
or U2363 (N_2363,N_35,N_1215);
nand U2364 (N_2364,N_258,N_1438);
nand U2365 (N_2365,N_947,N_897);
or U2366 (N_2366,N_236,N_459);
nand U2367 (N_2367,N_380,N_626);
xor U2368 (N_2368,N_694,N_53);
and U2369 (N_2369,N_739,N_1034);
or U2370 (N_2370,N_1106,N_287);
xnor U2371 (N_2371,N_1303,N_809);
nor U2372 (N_2372,N_1332,N_1197);
xor U2373 (N_2373,N_330,N_436);
and U2374 (N_2374,N_171,N_300);
nand U2375 (N_2375,N_57,N_444);
and U2376 (N_2376,N_672,N_1417);
nand U2377 (N_2377,N_526,N_852);
nor U2378 (N_2378,N_1489,N_329);
and U2379 (N_2379,N_1072,N_49);
nor U2380 (N_2380,N_1457,N_704);
and U2381 (N_2381,N_138,N_1231);
nand U2382 (N_2382,N_873,N_647);
and U2383 (N_2383,N_404,N_0);
or U2384 (N_2384,N_1207,N_1461);
nor U2385 (N_2385,N_675,N_1272);
and U2386 (N_2386,N_648,N_409);
nand U2387 (N_2387,N_546,N_652);
nor U2388 (N_2388,N_1478,N_1254);
nand U2389 (N_2389,N_382,N_541);
or U2390 (N_2390,N_1247,N_373);
and U2391 (N_2391,N_561,N_1028);
or U2392 (N_2392,N_24,N_1133);
nor U2393 (N_2393,N_1127,N_1085);
xor U2394 (N_2394,N_266,N_684);
xor U2395 (N_2395,N_854,N_601);
nor U2396 (N_2396,N_825,N_1391);
xor U2397 (N_2397,N_1215,N_732);
xor U2398 (N_2398,N_529,N_646);
and U2399 (N_2399,N_64,N_614);
nand U2400 (N_2400,N_932,N_728);
nand U2401 (N_2401,N_1142,N_609);
or U2402 (N_2402,N_279,N_725);
or U2403 (N_2403,N_64,N_397);
nand U2404 (N_2404,N_705,N_587);
nand U2405 (N_2405,N_679,N_85);
or U2406 (N_2406,N_705,N_1351);
nor U2407 (N_2407,N_515,N_1220);
nor U2408 (N_2408,N_1408,N_536);
or U2409 (N_2409,N_415,N_253);
and U2410 (N_2410,N_612,N_816);
nor U2411 (N_2411,N_783,N_1202);
nand U2412 (N_2412,N_595,N_434);
nor U2413 (N_2413,N_3,N_1047);
xor U2414 (N_2414,N_511,N_938);
or U2415 (N_2415,N_155,N_307);
nor U2416 (N_2416,N_1076,N_935);
xnor U2417 (N_2417,N_760,N_946);
and U2418 (N_2418,N_1286,N_647);
nand U2419 (N_2419,N_147,N_1075);
or U2420 (N_2420,N_1114,N_1453);
and U2421 (N_2421,N_884,N_270);
or U2422 (N_2422,N_1120,N_1339);
and U2423 (N_2423,N_420,N_90);
or U2424 (N_2424,N_568,N_594);
and U2425 (N_2425,N_573,N_295);
and U2426 (N_2426,N_314,N_368);
nand U2427 (N_2427,N_328,N_1126);
or U2428 (N_2428,N_1062,N_792);
nor U2429 (N_2429,N_809,N_1346);
nor U2430 (N_2430,N_761,N_755);
and U2431 (N_2431,N_339,N_76);
nor U2432 (N_2432,N_9,N_462);
nand U2433 (N_2433,N_379,N_956);
xor U2434 (N_2434,N_345,N_1158);
nand U2435 (N_2435,N_1102,N_50);
or U2436 (N_2436,N_684,N_118);
xnor U2437 (N_2437,N_522,N_344);
nor U2438 (N_2438,N_1287,N_749);
xor U2439 (N_2439,N_358,N_233);
and U2440 (N_2440,N_1012,N_1095);
nor U2441 (N_2441,N_844,N_1270);
or U2442 (N_2442,N_716,N_701);
or U2443 (N_2443,N_1073,N_1097);
and U2444 (N_2444,N_1062,N_1336);
or U2445 (N_2445,N_125,N_1183);
xnor U2446 (N_2446,N_968,N_431);
and U2447 (N_2447,N_367,N_165);
or U2448 (N_2448,N_469,N_1375);
or U2449 (N_2449,N_834,N_399);
nand U2450 (N_2450,N_751,N_80);
and U2451 (N_2451,N_1289,N_579);
nor U2452 (N_2452,N_94,N_1350);
and U2453 (N_2453,N_1373,N_1331);
nand U2454 (N_2454,N_992,N_203);
nand U2455 (N_2455,N_1311,N_1293);
nand U2456 (N_2456,N_1398,N_1244);
nor U2457 (N_2457,N_1250,N_897);
or U2458 (N_2458,N_698,N_1135);
nor U2459 (N_2459,N_589,N_570);
and U2460 (N_2460,N_664,N_1275);
nor U2461 (N_2461,N_889,N_1098);
nor U2462 (N_2462,N_470,N_1331);
nand U2463 (N_2463,N_1171,N_461);
nor U2464 (N_2464,N_485,N_923);
xnor U2465 (N_2465,N_821,N_644);
nor U2466 (N_2466,N_205,N_1310);
or U2467 (N_2467,N_885,N_693);
nand U2468 (N_2468,N_162,N_166);
or U2469 (N_2469,N_159,N_1401);
xnor U2470 (N_2470,N_42,N_872);
nand U2471 (N_2471,N_464,N_169);
nor U2472 (N_2472,N_582,N_376);
nand U2473 (N_2473,N_654,N_1165);
and U2474 (N_2474,N_8,N_912);
xor U2475 (N_2475,N_833,N_702);
or U2476 (N_2476,N_955,N_1012);
or U2477 (N_2477,N_1204,N_1179);
nand U2478 (N_2478,N_282,N_1327);
or U2479 (N_2479,N_1120,N_379);
nor U2480 (N_2480,N_35,N_1318);
nand U2481 (N_2481,N_855,N_89);
and U2482 (N_2482,N_1087,N_1315);
and U2483 (N_2483,N_1208,N_866);
and U2484 (N_2484,N_323,N_569);
and U2485 (N_2485,N_419,N_1030);
or U2486 (N_2486,N_540,N_162);
nand U2487 (N_2487,N_1337,N_1);
or U2488 (N_2488,N_1078,N_359);
xnor U2489 (N_2489,N_491,N_791);
nand U2490 (N_2490,N_815,N_590);
and U2491 (N_2491,N_69,N_1274);
nor U2492 (N_2492,N_867,N_1374);
nor U2493 (N_2493,N_1111,N_366);
nor U2494 (N_2494,N_1038,N_186);
or U2495 (N_2495,N_475,N_1288);
xor U2496 (N_2496,N_999,N_983);
xnor U2497 (N_2497,N_1145,N_470);
and U2498 (N_2498,N_291,N_301);
nand U2499 (N_2499,N_775,N_335);
and U2500 (N_2500,N_1321,N_222);
and U2501 (N_2501,N_1494,N_1050);
or U2502 (N_2502,N_562,N_524);
or U2503 (N_2503,N_113,N_589);
xnor U2504 (N_2504,N_1479,N_545);
nand U2505 (N_2505,N_1436,N_1455);
xnor U2506 (N_2506,N_1278,N_221);
nor U2507 (N_2507,N_175,N_253);
and U2508 (N_2508,N_592,N_728);
nor U2509 (N_2509,N_651,N_152);
or U2510 (N_2510,N_225,N_142);
or U2511 (N_2511,N_16,N_173);
nor U2512 (N_2512,N_1349,N_278);
nand U2513 (N_2513,N_1350,N_377);
and U2514 (N_2514,N_883,N_1471);
nand U2515 (N_2515,N_242,N_393);
and U2516 (N_2516,N_798,N_856);
nand U2517 (N_2517,N_1245,N_520);
nand U2518 (N_2518,N_1460,N_1350);
nor U2519 (N_2519,N_838,N_1475);
xor U2520 (N_2520,N_1133,N_526);
or U2521 (N_2521,N_12,N_1308);
and U2522 (N_2522,N_877,N_575);
nor U2523 (N_2523,N_833,N_1107);
and U2524 (N_2524,N_1223,N_733);
nand U2525 (N_2525,N_296,N_1);
and U2526 (N_2526,N_1457,N_304);
xor U2527 (N_2527,N_789,N_708);
nand U2528 (N_2528,N_851,N_1340);
and U2529 (N_2529,N_1326,N_1096);
or U2530 (N_2530,N_804,N_1479);
nand U2531 (N_2531,N_745,N_1461);
nor U2532 (N_2532,N_907,N_404);
nand U2533 (N_2533,N_312,N_1227);
and U2534 (N_2534,N_1407,N_1374);
nor U2535 (N_2535,N_1059,N_931);
nor U2536 (N_2536,N_347,N_1491);
xnor U2537 (N_2537,N_865,N_1006);
nor U2538 (N_2538,N_1197,N_46);
nor U2539 (N_2539,N_788,N_728);
nand U2540 (N_2540,N_1468,N_552);
and U2541 (N_2541,N_154,N_346);
and U2542 (N_2542,N_1241,N_398);
or U2543 (N_2543,N_118,N_61);
xor U2544 (N_2544,N_766,N_578);
nand U2545 (N_2545,N_1156,N_974);
and U2546 (N_2546,N_840,N_96);
or U2547 (N_2547,N_305,N_377);
xor U2548 (N_2548,N_180,N_426);
nor U2549 (N_2549,N_929,N_1061);
nor U2550 (N_2550,N_978,N_447);
nor U2551 (N_2551,N_1254,N_579);
and U2552 (N_2552,N_1326,N_1194);
nor U2553 (N_2553,N_155,N_762);
nor U2554 (N_2554,N_830,N_772);
nor U2555 (N_2555,N_792,N_793);
nor U2556 (N_2556,N_1148,N_813);
nand U2557 (N_2557,N_1218,N_321);
or U2558 (N_2558,N_620,N_994);
and U2559 (N_2559,N_990,N_1152);
nand U2560 (N_2560,N_375,N_1389);
nand U2561 (N_2561,N_1072,N_791);
nor U2562 (N_2562,N_600,N_1315);
nor U2563 (N_2563,N_900,N_1097);
or U2564 (N_2564,N_873,N_417);
or U2565 (N_2565,N_1476,N_1231);
nand U2566 (N_2566,N_548,N_688);
xor U2567 (N_2567,N_1330,N_767);
nor U2568 (N_2568,N_927,N_366);
or U2569 (N_2569,N_1105,N_986);
or U2570 (N_2570,N_1310,N_294);
or U2571 (N_2571,N_587,N_252);
and U2572 (N_2572,N_1459,N_846);
and U2573 (N_2573,N_523,N_238);
or U2574 (N_2574,N_1287,N_397);
or U2575 (N_2575,N_80,N_448);
or U2576 (N_2576,N_1285,N_1089);
or U2577 (N_2577,N_485,N_705);
or U2578 (N_2578,N_1108,N_389);
or U2579 (N_2579,N_775,N_1339);
and U2580 (N_2580,N_1144,N_139);
nor U2581 (N_2581,N_947,N_1126);
xor U2582 (N_2582,N_887,N_64);
nor U2583 (N_2583,N_1212,N_37);
or U2584 (N_2584,N_521,N_204);
nor U2585 (N_2585,N_1264,N_388);
and U2586 (N_2586,N_681,N_501);
nand U2587 (N_2587,N_737,N_1084);
or U2588 (N_2588,N_311,N_1336);
nand U2589 (N_2589,N_1450,N_798);
or U2590 (N_2590,N_125,N_655);
nand U2591 (N_2591,N_1352,N_245);
or U2592 (N_2592,N_481,N_53);
nor U2593 (N_2593,N_1224,N_119);
nand U2594 (N_2594,N_808,N_384);
or U2595 (N_2595,N_447,N_356);
nor U2596 (N_2596,N_346,N_750);
or U2597 (N_2597,N_349,N_136);
or U2598 (N_2598,N_959,N_427);
nand U2599 (N_2599,N_607,N_503);
nor U2600 (N_2600,N_335,N_62);
or U2601 (N_2601,N_1172,N_616);
nor U2602 (N_2602,N_938,N_311);
nand U2603 (N_2603,N_1441,N_1125);
nor U2604 (N_2604,N_546,N_231);
nor U2605 (N_2605,N_1309,N_545);
or U2606 (N_2606,N_405,N_789);
nor U2607 (N_2607,N_1157,N_802);
and U2608 (N_2608,N_114,N_629);
xor U2609 (N_2609,N_1315,N_114);
nand U2610 (N_2610,N_144,N_195);
nor U2611 (N_2611,N_1026,N_469);
or U2612 (N_2612,N_888,N_400);
xnor U2613 (N_2613,N_1439,N_469);
xnor U2614 (N_2614,N_873,N_750);
nand U2615 (N_2615,N_329,N_614);
nor U2616 (N_2616,N_542,N_793);
nor U2617 (N_2617,N_1158,N_668);
nor U2618 (N_2618,N_630,N_607);
nor U2619 (N_2619,N_1005,N_804);
xor U2620 (N_2620,N_1306,N_418);
nand U2621 (N_2621,N_1340,N_1436);
nand U2622 (N_2622,N_542,N_1364);
nor U2623 (N_2623,N_102,N_580);
nand U2624 (N_2624,N_1489,N_1093);
xnor U2625 (N_2625,N_7,N_1192);
and U2626 (N_2626,N_846,N_504);
or U2627 (N_2627,N_573,N_983);
nand U2628 (N_2628,N_1404,N_595);
and U2629 (N_2629,N_1307,N_558);
nand U2630 (N_2630,N_1089,N_159);
or U2631 (N_2631,N_358,N_45);
xnor U2632 (N_2632,N_234,N_735);
nand U2633 (N_2633,N_98,N_989);
nand U2634 (N_2634,N_615,N_1478);
nand U2635 (N_2635,N_667,N_905);
nor U2636 (N_2636,N_1267,N_364);
nand U2637 (N_2637,N_22,N_1413);
nand U2638 (N_2638,N_144,N_445);
nand U2639 (N_2639,N_423,N_232);
nand U2640 (N_2640,N_457,N_851);
nor U2641 (N_2641,N_1406,N_1090);
and U2642 (N_2642,N_1305,N_1061);
nand U2643 (N_2643,N_27,N_985);
nand U2644 (N_2644,N_1467,N_1163);
nand U2645 (N_2645,N_329,N_513);
nand U2646 (N_2646,N_1110,N_85);
nand U2647 (N_2647,N_923,N_551);
and U2648 (N_2648,N_256,N_1307);
nand U2649 (N_2649,N_404,N_1247);
or U2650 (N_2650,N_722,N_158);
nand U2651 (N_2651,N_517,N_64);
or U2652 (N_2652,N_1030,N_1476);
or U2653 (N_2653,N_696,N_1193);
nor U2654 (N_2654,N_1339,N_963);
or U2655 (N_2655,N_1410,N_0);
and U2656 (N_2656,N_696,N_1402);
nor U2657 (N_2657,N_305,N_782);
and U2658 (N_2658,N_1456,N_1435);
nand U2659 (N_2659,N_40,N_464);
or U2660 (N_2660,N_602,N_1249);
nand U2661 (N_2661,N_1082,N_1073);
nand U2662 (N_2662,N_410,N_1141);
xor U2663 (N_2663,N_1226,N_328);
nor U2664 (N_2664,N_491,N_1186);
nand U2665 (N_2665,N_1394,N_723);
or U2666 (N_2666,N_1144,N_1066);
and U2667 (N_2667,N_1323,N_21);
nand U2668 (N_2668,N_829,N_1330);
and U2669 (N_2669,N_198,N_732);
nor U2670 (N_2670,N_620,N_739);
nor U2671 (N_2671,N_336,N_1101);
nand U2672 (N_2672,N_358,N_780);
nand U2673 (N_2673,N_551,N_27);
or U2674 (N_2674,N_962,N_683);
or U2675 (N_2675,N_687,N_1371);
nand U2676 (N_2676,N_619,N_959);
nand U2677 (N_2677,N_1126,N_522);
or U2678 (N_2678,N_682,N_698);
nor U2679 (N_2679,N_573,N_1490);
or U2680 (N_2680,N_881,N_837);
and U2681 (N_2681,N_284,N_662);
nand U2682 (N_2682,N_1285,N_4);
and U2683 (N_2683,N_758,N_737);
and U2684 (N_2684,N_287,N_1109);
nand U2685 (N_2685,N_1494,N_1432);
or U2686 (N_2686,N_382,N_55);
xor U2687 (N_2687,N_1332,N_501);
nand U2688 (N_2688,N_1193,N_677);
nand U2689 (N_2689,N_1088,N_499);
nor U2690 (N_2690,N_851,N_683);
nand U2691 (N_2691,N_303,N_146);
or U2692 (N_2692,N_1180,N_500);
nor U2693 (N_2693,N_811,N_429);
or U2694 (N_2694,N_616,N_473);
xnor U2695 (N_2695,N_892,N_575);
nor U2696 (N_2696,N_1132,N_226);
or U2697 (N_2697,N_488,N_842);
or U2698 (N_2698,N_569,N_26);
or U2699 (N_2699,N_1217,N_5);
nor U2700 (N_2700,N_1335,N_1385);
or U2701 (N_2701,N_1403,N_334);
nand U2702 (N_2702,N_360,N_254);
nor U2703 (N_2703,N_43,N_485);
nand U2704 (N_2704,N_1413,N_525);
nand U2705 (N_2705,N_1036,N_462);
nand U2706 (N_2706,N_966,N_741);
nor U2707 (N_2707,N_364,N_1201);
nor U2708 (N_2708,N_1009,N_963);
and U2709 (N_2709,N_994,N_43);
xor U2710 (N_2710,N_309,N_419);
or U2711 (N_2711,N_1451,N_614);
nor U2712 (N_2712,N_368,N_864);
xor U2713 (N_2713,N_881,N_1437);
nor U2714 (N_2714,N_103,N_1126);
nor U2715 (N_2715,N_1318,N_394);
xnor U2716 (N_2716,N_1078,N_1219);
nor U2717 (N_2717,N_145,N_827);
nor U2718 (N_2718,N_453,N_12);
nor U2719 (N_2719,N_1168,N_99);
nand U2720 (N_2720,N_1268,N_273);
nor U2721 (N_2721,N_297,N_650);
and U2722 (N_2722,N_1056,N_359);
and U2723 (N_2723,N_312,N_1152);
nand U2724 (N_2724,N_1319,N_1196);
nor U2725 (N_2725,N_65,N_325);
xnor U2726 (N_2726,N_871,N_135);
nand U2727 (N_2727,N_452,N_1107);
or U2728 (N_2728,N_235,N_111);
nand U2729 (N_2729,N_624,N_1053);
and U2730 (N_2730,N_462,N_311);
xor U2731 (N_2731,N_48,N_245);
or U2732 (N_2732,N_1063,N_300);
nor U2733 (N_2733,N_713,N_50);
nand U2734 (N_2734,N_93,N_516);
xor U2735 (N_2735,N_65,N_1190);
and U2736 (N_2736,N_8,N_1097);
and U2737 (N_2737,N_808,N_662);
and U2738 (N_2738,N_613,N_1400);
and U2739 (N_2739,N_1036,N_553);
or U2740 (N_2740,N_493,N_1437);
nor U2741 (N_2741,N_944,N_840);
nand U2742 (N_2742,N_380,N_59);
or U2743 (N_2743,N_1121,N_45);
xor U2744 (N_2744,N_235,N_1322);
and U2745 (N_2745,N_914,N_855);
nor U2746 (N_2746,N_299,N_1058);
nor U2747 (N_2747,N_957,N_326);
nor U2748 (N_2748,N_235,N_600);
nand U2749 (N_2749,N_1172,N_1422);
nand U2750 (N_2750,N_760,N_1222);
or U2751 (N_2751,N_1406,N_882);
and U2752 (N_2752,N_86,N_966);
nand U2753 (N_2753,N_508,N_674);
and U2754 (N_2754,N_237,N_1441);
xnor U2755 (N_2755,N_1109,N_220);
xnor U2756 (N_2756,N_509,N_16);
nor U2757 (N_2757,N_42,N_578);
and U2758 (N_2758,N_1382,N_1153);
or U2759 (N_2759,N_348,N_615);
or U2760 (N_2760,N_20,N_405);
or U2761 (N_2761,N_885,N_954);
and U2762 (N_2762,N_219,N_730);
xnor U2763 (N_2763,N_1343,N_1203);
and U2764 (N_2764,N_821,N_755);
nand U2765 (N_2765,N_651,N_369);
xor U2766 (N_2766,N_594,N_1257);
xor U2767 (N_2767,N_1107,N_1091);
and U2768 (N_2768,N_1451,N_1134);
and U2769 (N_2769,N_1143,N_1198);
or U2770 (N_2770,N_1282,N_1356);
nor U2771 (N_2771,N_431,N_776);
or U2772 (N_2772,N_11,N_1148);
and U2773 (N_2773,N_688,N_545);
or U2774 (N_2774,N_861,N_562);
or U2775 (N_2775,N_902,N_1289);
nand U2776 (N_2776,N_281,N_493);
or U2777 (N_2777,N_994,N_93);
nand U2778 (N_2778,N_799,N_938);
nand U2779 (N_2779,N_768,N_495);
nor U2780 (N_2780,N_897,N_494);
nor U2781 (N_2781,N_598,N_961);
nor U2782 (N_2782,N_1171,N_818);
xnor U2783 (N_2783,N_337,N_244);
nand U2784 (N_2784,N_657,N_392);
and U2785 (N_2785,N_1301,N_487);
or U2786 (N_2786,N_403,N_259);
xor U2787 (N_2787,N_1348,N_1099);
and U2788 (N_2788,N_1390,N_1017);
nand U2789 (N_2789,N_14,N_930);
nor U2790 (N_2790,N_929,N_1376);
nor U2791 (N_2791,N_1117,N_333);
nand U2792 (N_2792,N_34,N_989);
or U2793 (N_2793,N_850,N_432);
nand U2794 (N_2794,N_1194,N_739);
nand U2795 (N_2795,N_595,N_636);
nor U2796 (N_2796,N_50,N_968);
nor U2797 (N_2797,N_1085,N_464);
or U2798 (N_2798,N_1411,N_856);
or U2799 (N_2799,N_842,N_1225);
xor U2800 (N_2800,N_671,N_203);
nor U2801 (N_2801,N_308,N_1394);
nor U2802 (N_2802,N_380,N_429);
xor U2803 (N_2803,N_920,N_169);
and U2804 (N_2804,N_406,N_1305);
nor U2805 (N_2805,N_1277,N_375);
nor U2806 (N_2806,N_349,N_119);
xor U2807 (N_2807,N_1420,N_153);
nand U2808 (N_2808,N_649,N_942);
or U2809 (N_2809,N_339,N_1292);
nor U2810 (N_2810,N_499,N_1142);
or U2811 (N_2811,N_1250,N_612);
nor U2812 (N_2812,N_361,N_544);
nand U2813 (N_2813,N_563,N_1028);
nor U2814 (N_2814,N_1197,N_82);
nor U2815 (N_2815,N_1080,N_49);
nand U2816 (N_2816,N_859,N_637);
nor U2817 (N_2817,N_1044,N_61);
nand U2818 (N_2818,N_1270,N_1445);
and U2819 (N_2819,N_1420,N_1453);
nor U2820 (N_2820,N_805,N_317);
nand U2821 (N_2821,N_1087,N_900);
nand U2822 (N_2822,N_818,N_38);
or U2823 (N_2823,N_564,N_298);
or U2824 (N_2824,N_598,N_1307);
nor U2825 (N_2825,N_937,N_1485);
nor U2826 (N_2826,N_954,N_773);
nand U2827 (N_2827,N_140,N_1210);
and U2828 (N_2828,N_216,N_1175);
nand U2829 (N_2829,N_289,N_590);
nor U2830 (N_2830,N_1264,N_645);
or U2831 (N_2831,N_1114,N_1350);
nor U2832 (N_2832,N_781,N_213);
nand U2833 (N_2833,N_196,N_582);
or U2834 (N_2834,N_1175,N_72);
or U2835 (N_2835,N_486,N_1464);
nand U2836 (N_2836,N_107,N_21);
nor U2837 (N_2837,N_1212,N_158);
or U2838 (N_2838,N_1212,N_905);
and U2839 (N_2839,N_251,N_741);
xor U2840 (N_2840,N_1494,N_275);
nand U2841 (N_2841,N_1338,N_62);
or U2842 (N_2842,N_575,N_1353);
or U2843 (N_2843,N_563,N_725);
xor U2844 (N_2844,N_103,N_600);
nand U2845 (N_2845,N_214,N_194);
or U2846 (N_2846,N_1084,N_226);
nand U2847 (N_2847,N_1420,N_1012);
and U2848 (N_2848,N_412,N_637);
or U2849 (N_2849,N_1281,N_1276);
or U2850 (N_2850,N_1128,N_533);
or U2851 (N_2851,N_411,N_1247);
and U2852 (N_2852,N_1168,N_949);
nor U2853 (N_2853,N_1399,N_298);
nor U2854 (N_2854,N_1425,N_319);
and U2855 (N_2855,N_462,N_745);
or U2856 (N_2856,N_1176,N_1399);
and U2857 (N_2857,N_701,N_1382);
and U2858 (N_2858,N_1114,N_300);
or U2859 (N_2859,N_753,N_451);
and U2860 (N_2860,N_1356,N_709);
nand U2861 (N_2861,N_311,N_587);
nor U2862 (N_2862,N_995,N_1298);
and U2863 (N_2863,N_926,N_1417);
xnor U2864 (N_2864,N_279,N_829);
nand U2865 (N_2865,N_534,N_912);
xor U2866 (N_2866,N_1497,N_972);
nor U2867 (N_2867,N_1037,N_16);
or U2868 (N_2868,N_1464,N_322);
or U2869 (N_2869,N_361,N_893);
and U2870 (N_2870,N_123,N_360);
xor U2871 (N_2871,N_1121,N_357);
or U2872 (N_2872,N_933,N_593);
nand U2873 (N_2873,N_748,N_178);
and U2874 (N_2874,N_1087,N_447);
nand U2875 (N_2875,N_1494,N_1164);
nand U2876 (N_2876,N_800,N_21);
and U2877 (N_2877,N_379,N_496);
nand U2878 (N_2878,N_128,N_1227);
and U2879 (N_2879,N_1346,N_1150);
nand U2880 (N_2880,N_666,N_332);
nand U2881 (N_2881,N_1397,N_831);
xor U2882 (N_2882,N_87,N_191);
nand U2883 (N_2883,N_1478,N_1095);
xor U2884 (N_2884,N_128,N_1412);
nand U2885 (N_2885,N_969,N_246);
or U2886 (N_2886,N_136,N_203);
nand U2887 (N_2887,N_1304,N_132);
nand U2888 (N_2888,N_1019,N_1063);
nand U2889 (N_2889,N_1292,N_361);
and U2890 (N_2890,N_315,N_833);
nor U2891 (N_2891,N_836,N_595);
nor U2892 (N_2892,N_828,N_1451);
xnor U2893 (N_2893,N_559,N_75);
nor U2894 (N_2894,N_1438,N_1446);
or U2895 (N_2895,N_772,N_1259);
or U2896 (N_2896,N_1288,N_327);
nor U2897 (N_2897,N_979,N_248);
and U2898 (N_2898,N_298,N_693);
nand U2899 (N_2899,N_1468,N_440);
and U2900 (N_2900,N_184,N_295);
nor U2901 (N_2901,N_293,N_413);
nor U2902 (N_2902,N_966,N_421);
xor U2903 (N_2903,N_601,N_1400);
and U2904 (N_2904,N_419,N_54);
nor U2905 (N_2905,N_401,N_1312);
nand U2906 (N_2906,N_1333,N_636);
xor U2907 (N_2907,N_497,N_402);
nor U2908 (N_2908,N_352,N_490);
xnor U2909 (N_2909,N_942,N_139);
xnor U2910 (N_2910,N_1257,N_1228);
nand U2911 (N_2911,N_1406,N_999);
nor U2912 (N_2912,N_1128,N_437);
nor U2913 (N_2913,N_1440,N_317);
nand U2914 (N_2914,N_548,N_106);
and U2915 (N_2915,N_669,N_1278);
and U2916 (N_2916,N_1423,N_569);
or U2917 (N_2917,N_1183,N_459);
nand U2918 (N_2918,N_1310,N_1008);
xor U2919 (N_2919,N_984,N_491);
nand U2920 (N_2920,N_190,N_1055);
or U2921 (N_2921,N_294,N_1455);
or U2922 (N_2922,N_1251,N_788);
or U2923 (N_2923,N_1305,N_1446);
nand U2924 (N_2924,N_1115,N_1438);
and U2925 (N_2925,N_669,N_814);
nand U2926 (N_2926,N_184,N_1064);
nor U2927 (N_2927,N_407,N_372);
nor U2928 (N_2928,N_262,N_253);
or U2929 (N_2929,N_535,N_980);
nor U2930 (N_2930,N_413,N_1441);
nand U2931 (N_2931,N_450,N_1469);
and U2932 (N_2932,N_1085,N_1363);
nor U2933 (N_2933,N_339,N_1104);
nor U2934 (N_2934,N_462,N_106);
nor U2935 (N_2935,N_278,N_39);
and U2936 (N_2936,N_658,N_1073);
or U2937 (N_2937,N_683,N_1098);
and U2938 (N_2938,N_1398,N_597);
nor U2939 (N_2939,N_1226,N_1342);
xnor U2940 (N_2940,N_648,N_816);
or U2941 (N_2941,N_1002,N_1215);
or U2942 (N_2942,N_1159,N_125);
or U2943 (N_2943,N_1398,N_1103);
xor U2944 (N_2944,N_1449,N_1099);
and U2945 (N_2945,N_677,N_246);
xnor U2946 (N_2946,N_1279,N_1164);
and U2947 (N_2947,N_593,N_665);
nand U2948 (N_2948,N_1004,N_511);
and U2949 (N_2949,N_1242,N_821);
or U2950 (N_2950,N_1467,N_1308);
and U2951 (N_2951,N_369,N_837);
and U2952 (N_2952,N_48,N_876);
nor U2953 (N_2953,N_1396,N_795);
nand U2954 (N_2954,N_1071,N_167);
or U2955 (N_2955,N_1427,N_315);
nor U2956 (N_2956,N_1089,N_390);
nand U2957 (N_2957,N_55,N_473);
xnor U2958 (N_2958,N_1372,N_321);
nand U2959 (N_2959,N_1054,N_938);
or U2960 (N_2960,N_1325,N_847);
or U2961 (N_2961,N_712,N_653);
nor U2962 (N_2962,N_733,N_307);
and U2963 (N_2963,N_1129,N_249);
nor U2964 (N_2964,N_971,N_783);
nand U2965 (N_2965,N_691,N_1489);
and U2966 (N_2966,N_574,N_1069);
or U2967 (N_2967,N_458,N_978);
nor U2968 (N_2968,N_118,N_503);
xnor U2969 (N_2969,N_682,N_225);
and U2970 (N_2970,N_446,N_480);
or U2971 (N_2971,N_162,N_360);
nand U2972 (N_2972,N_447,N_1288);
and U2973 (N_2973,N_202,N_265);
or U2974 (N_2974,N_1389,N_1288);
and U2975 (N_2975,N_1283,N_1360);
and U2976 (N_2976,N_161,N_1246);
and U2977 (N_2977,N_978,N_1114);
nor U2978 (N_2978,N_459,N_275);
or U2979 (N_2979,N_244,N_506);
or U2980 (N_2980,N_335,N_378);
nand U2981 (N_2981,N_260,N_276);
nand U2982 (N_2982,N_863,N_480);
nand U2983 (N_2983,N_1383,N_404);
and U2984 (N_2984,N_545,N_1024);
nor U2985 (N_2985,N_169,N_268);
nor U2986 (N_2986,N_519,N_763);
and U2987 (N_2987,N_149,N_679);
xnor U2988 (N_2988,N_453,N_1395);
nor U2989 (N_2989,N_1294,N_720);
or U2990 (N_2990,N_1196,N_1400);
or U2991 (N_2991,N_914,N_532);
and U2992 (N_2992,N_690,N_804);
or U2993 (N_2993,N_1111,N_1301);
and U2994 (N_2994,N_383,N_1062);
and U2995 (N_2995,N_1153,N_356);
and U2996 (N_2996,N_414,N_977);
nand U2997 (N_2997,N_895,N_236);
or U2998 (N_2998,N_922,N_455);
and U2999 (N_2999,N_767,N_217);
nand U3000 (N_3000,N_2066,N_2377);
nor U3001 (N_3001,N_1733,N_2045);
and U3002 (N_3002,N_2807,N_2405);
and U3003 (N_3003,N_2206,N_2239);
and U3004 (N_3004,N_2642,N_2976);
or U3005 (N_3005,N_1897,N_2559);
nor U3006 (N_3006,N_2743,N_2628);
or U3007 (N_3007,N_2654,N_1589);
nor U3008 (N_3008,N_2235,N_2151);
and U3009 (N_3009,N_2364,N_2091);
nand U3010 (N_3010,N_2831,N_2866);
nor U3011 (N_3011,N_2798,N_2689);
nand U3012 (N_3012,N_1618,N_2898);
and U3013 (N_3013,N_2508,N_1506);
nor U3014 (N_3014,N_1602,N_2453);
and U3015 (N_3015,N_2070,N_2375);
and U3016 (N_3016,N_1824,N_2115);
xnor U3017 (N_3017,N_1683,N_2777);
and U3018 (N_3018,N_2047,N_1871);
nand U3019 (N_3019,N_2495,N_2008);
nand U3020 (N_3020,N_1641,N_1832);
and U3021 (N_3021,N_2611,N_2282);
nand U3022 (N_3022,N_1638,N_2789);
or U3023 (N_3023,N_1890,N_1521);
nand U3024 (N_3024,N_2240,N_2549);
or U3025 (N_3025,N_2053,N_2722);
or U3026 (N_3026,N_1502,N_2744);
nor U3027 (N_3027,N_1561,N_2470);
nor U3028 (N_3028,N_2020,N_1863);
xnor U3029 (N_3029,N_1645,N_1840);
and U3030 (N_3030,N_2287,N_1825);
or U3031 (N_3031,N_1941,N_2466);
or U3032 (N_3032,N_1912,N_2249);
and U3033 (N_3033,N_2938,N_2809);
xnor U3034 (N_3034,N_2414,N_2254);
or U3035 (N_3035,N_2225,N_1792);
and U3036 (N_3036,N_1877,N_1859);
nor U3037 (N_3037,N_2877,N_1887);
and U3038 (N_3038,N_1766,N_1543);
nor U3039 (N_3039,N_1757,N_1965);
nand U3040 (N_3040,N_2551,N_2896);
nor U3041 (N_3041,N_2185,N_1553);
nor U3042 (N_3042,N_1624,N_2538);
nand U3043 (N_3043,N_2221,N_2431);
xnor U3044 (N_3044,N_2701,N_1868);
or U3045 (N_3045,N_1791,N_2144);
nand U3046 (N_3046,N_1558,N_2526);
nor U3047 (N_3047,N_2463,N_1844);
xor U3048 (N_3048,N_2016,N_2709);
and U3049 (N_3049,N_2887,N_1729);
nor U3050 (N_3050,N_2696,N_1940);
or U3051 (N_3051,N_2698,N_2399);
and U3052 (N_3052,N_2803,N_1956);
nor U3053 (N_3053,N_1904,N_2623);
xor U3054 (N_3054,N_1915,N_2356);
or U3055 (N_3055,N_2906,N_2686);
and U3056 (N_3056,N_2272,N_2592);
or U3057 (N_3057,N_2425,N_1636);
nor U3058 (N_3058,N_2557,N_2624);
nor U3059 (N_3059,N_2941,N_1793);
or U3060 (N_3060,N_2268,N_2299);
nand U3061 (N_3061,N_1749,N_2665);
nand U3062 (N_3062,N_2552,N_2649);
and U3063 (N_3063,N_2251,N_2378);
nand U3064 (N_3064,N_2710,N_1613);
nor U3065 (N_3065,N_2847,N_2093);
and U3066 (N_3066,N_1552,N_1807);
nand U3067 (N_3067,N_2325,N_2021);
nor U3068 (N_3068,N_2682,N_1660);
nor U3069 (N_3069,N_2633,N_2022);
nand U3070 (N_3070,N_1582,N_2494);
nand U3071 (N_3071,N_1635,N_1559);
nor U3072 (N_3072,N_1984,N_1934);
or U3073 (N_3073,N_2591,N_2864);
or U3074 (N_3074,N_1676,N_2339);
and U3075 (N_3075,N_1978,N_2781);
nor U3076 (N_3076,N_2818,N_2681);
or U3077 (N_3077,N_1574,N_2492);
nand U3078 (N_3078,N_1736,N_1668);
nor U3079 (N_3079,N_2622,N_2488);
nor U3080 (N_3080,N_1856,N_2291);
nor U3081 (N_3081,N_2835,N_2977);
or U3082 (N_3082,N_2715,N_2416);
and U3083 (N_3083,N_2933,N_1981);
nand U3084 (N_3084,N_2227,N_1776);
xor U3085 (N_3085,N_2300,N_2891);
or U3086 (N_3086,N_2385,N_1894);
and U3087 (N_3087,N_2674,N_2676);
xor U3088 (N_3088,N_2276,N_2188);
or U3089 (N_3089,N_1942,N_2612);
or U3090 (N_3090,N_2255,N_1741);
nor U3091 (N_3091,N_1661,N_2775);
nand U3092 (N_3092,N_2130,N_2918);
xor U3093 (N_3093,N_2027,N_2195);
nor U3094 (N_3094,N_2924,N_1518);
nand U3095 (N_3095,N_2156,N_2305);
nor U3096 (N_3096,N_2072,N_2384);
or U3097 (N_3097,N_1747,N_1560);
and U3098 (N_3098,N_1616,N_2764);
xor U3099 (N_3099,N_2514,N_1798);
nand U3100 (N_3100,N_2838,N_2018);
nor U3101 (N_3101,N_1900,N_2815);
nand U3102 (N_3102,N_1803,N_2229);
xnor U3103 (N_3103,N_1761,N_2830);
or U3104 (N_3104,N_2051,N_1533);
nand U3105 (N_3105,N_2015,N_2387);
or U3106 (N_3106,N_2161,N_2304);
or U3107 (N_3107,N_2913,N_2565);
or U3108 (N_3108,N_2921,N_1802);
nand U3109 (N_3109,N_2140,N_1622);
nand U3110 (N_3110,N_2245,N_2116);
xnor U3111 (N_3111,N_2410,N_2865);
nand U3112 (N_3112,N_1760,N_2162);
or U3113 (N_3113,N_2758,N_2226);
nor U3114 (N_3114,N_2203,N_2576);
or U3115 (N_3115,N_2736,N_1691);
nor U3116 (N_3116,N_2505,N_1516);
and U3117 (N_3117,N_2573,N_2491);
or U3118 (N_3118,N_2780,N_2089);
xor U3119 (N_3119,N_1918,N_1673);
and U3120 (N_3120,N_1637,N_1875);
and U3121 (N_3121,N_2895,N_1801);
nor U3122 (N_3122,N_2143,N_2450);
and U3123 (N_3123,N_2026,N_2944);
nand U3124 (N_3124,N_2121,N_2571);
xnor U3125 (N_3125,N_2783,N_1655);
or U3126 (N_3126,N_1563,N_2699);
nor U3127 (N_3127,N_2168,N_2312);
and U3128 (N_3128,N_1666,N_2587);
and U3129 (N_3129,N_2480,N_1753);
nor U3130 (N_3130,N_2473,N_2432);
and U3131 (N_3131,N_2281,N_1575);
nor U3132 (N_3132,N_2355,N_2313);
nor U3133 (N_3133,N_2760,N_2620);
xor U3134 (N_3134,N_2248,N_1706);
nand U3135 (N_3135,N_1961,N_1579);
nor U3136 (N_3136,N_2999,N_2678);
or U3137 (N_3137,N_2196,N_2128);
nor U3138 (N_3138,N_2001,N_2421);
and U3139 (N_3139,N_2094,N_2037);
nand U3140 (N_3140,N_2853,N_2347);
nor U3141 (N_3141,N_2522,N_2606);
nand U3142 (N_3142,N_2126,N_2497);
nand U3143 (N_3143,N_1500,N_2289);
and U3144 (N_3144,N_2985,N_1649);
and U3145 (N_3145,N_2036,N_1765);
nor U3146 (N_3146,N_1948,N_2409);
nand U3147 (N_3147,N_2258,N_2728);
or U3148 (N_3148,N_2321,N_1855);
and U3149 (N_3149,N_2261,N_2619);
and U3150 (N_3150,N_2250,N_2989);
nand U3151 (N_3151,N_2669,N_2537);
or U3152 (N_3152,N_2486,N_2543);
nand U3153 (N_3153,N_1848,N_1779);
nand U3154 (N_3154,N_2518,N_1669);
xor U3155 (N_3155,N_2039,N_2886);
nor U3156 (N_3156,N_2220,N_2031);
nor U3157 (N_3157,N_2296,N_2916);
or U3158 (N_3158,N_2101,N_2376);
xor U3159 (N_3159,N_2959,N_2626);
or U3160 (N_3160,N_1611,N_2230);
nand U3161 (N_3161,N_2407,N_2012);
and U3162 (N_3162,N_2829,N_1962);
nand U3163 (N_3163,N_2969,N_2653);
xor U3164 (N_3164,N_1991,N_1966);
nand U3165 (N_3165,N_2169,N_2788);
and U3166 (N_3166,N_1963,N_1999);
nand U3167 (N_3167,N_1805,N_2867);
nand U3168 (N_3168,N_1505,N_2228);
and U3169 (N_3169,N_1684,N_1708);
nand U3170 (N_3170,N_2640,N_2588);
nand U3171 (N_3171,N_1800,N_1540);
and U3172 (N_3172,N_1623,N_2883);
nor U3173 (N_3173,N_2216,N_1590);
or U3174 (N_3174,N_2186,N_2420);
nand U3175 (N_3175,N_1958,N_1536);
and U3176 (N_3176,N_2833,N_1763);
nor U3177 (N_3177,N_2310,N_1852);
or U3178 (N_3178,N_2350,N_2721);
nor U3179 (N_3179,N_2187,N_2753);
or U3180 (N_3180,N_2150,N_2825);
xor U3181 (N_3181,N_2232,N_2382);
nor U3182 (N_3182,N_1930,N_2610);
nand U3183 (N_3183,N_2604,N_2935);
and U3184 (N_3184,N_2981,N_2961);
nand U3185 (N_3185,N_2210,N_2550);
nand U3186 (N_3186,N_1921,N_2890);
or U3187 (N_3187,N_2556,N_2373);
nand U3188 (N_3188,N_2123,N_1599);
nand U3189 (N_3189,N_2801,N_2994);
nand U3190 (N_3190,N_1644,N_2205);
or U3191 (N_3191,N_1899,N_2451);
nand U3192 (N_3192,N_1833,N_1857);
nor U3193 (N_3193,N_1569,N_1537);
or U3194 (N_3194,N_2279,N_2629);
xor U3195 (N_3195,N_2814,N_1738);
or U3196 (N_3196,N_2060,N_2802);
and U3197 (N_3197,N_2554,N_2766);
or U3198 (N_3198,N_2396,N_1804);
and U3199 (N_3199,N_2761,N_1694);
nor U3200 (N_3200,N_1931,N_1898);
nand U3201 (N_3201,N_1994,N_1851);
or U3202 (N_3202,N_2157,N_2112);
nand U3203 (N_3203,N_2481,N_2395);
or U3204 (N_3204,N_2343,N_1628);
and U3205 (N_3205,N_2237,N_2908);
or U3206 (N_3206,N_1550,N_2437);
and U3207 (N_3207,N_2170,N_1843);
and U3208 (N_3208,N_1861,N_2820);
nand U3209 (N_3209,N_1858,N_2851);
xor U3210 (N_3210,N_2105,N_2411);
or U3211 (N_3211,N_2583,N_2530);
nor U3212 (N_3212,N_1593,N_1703);
xor U3213 (N_3213,N_1768,N_1634);
nor U3214 (N_3214,N_1773,N_2293);
and U3215 (N_3215,N_2794,N_2850);
and U3216 (N_3216,N_2134,N_2363);
nand U3217 (N_3217,N_1722,N_2749);
nand U3218 (N_3218,N_2233,N_2708);
nor U3219 (N_3219,N_2618,N_1514);
and U3220 (N_3220,N_2752,N_2878);
nand U3221 (N_3221,N_2058,N_2799);
or U3222 (N_3222,N_2177,N_2362);
and U3223 (N_3223,N_2462,N_2863);
xor U3224 (N_3224,N_1985,N_2418);
nand U3225 (N_3225,N_2962,N_2404);
nor U3226 (N_3226,N_1678,N_1554);
or U3227 (N_3227,N_2625,N_1874);
nand U3228 (N_3228,N_2762,N_2002);
nor U3229 (N_3229,N_2352,N_1925);
or U3230 (N_3230,N_2754,N_2381);
and U3231 (N_3231,N_1911,N_2246);
nor U3232 (N_3232,N_2900,N_2737);
and U3233 (N_3233,N_2991,N_1810);
xor U3234 (N_3234,N_2057,N_1996);
nand U3235 (N_3235,N_1546,N_1762);
and U3236 (N_3236,N_2957,N_2322);
nand U3237 (N_3237,N_1515,N_2950);
and U3238 (N_3238,N_1696,N_2525);
and U3239 (N_3239,N_1625,N_2178);
or U3240 (N_3240,N_2566,N_1631);
or U3241 (N_3241,N_1817,N_2848);
and U3242 (N_3242,N_1919,N_1547);
and U3243 (N_3243,N_2876,N_2067);
xor U3244 (N_3244,N_1971,N_2812);
nand U3245 (N_3245,N_2380,N_2262);
and U3246 (N_3246,N_2646,N_2298);
and U3247 (N_3247,N_1545,N_1995);
nor U3248 (N_3248,N_1924,N_2517);
or U3249 (N_3249,N_1835,N_1717);
nand U3250 (N_3250,N_2614,N_2454);
and U3251 (N_3251,N_2483,N_1781);
nor U3252 (N_3252,N_1656,N_2111);
nand U3253 (N_3253,N_2397,N_1821);
nor U3254 (N_3254,N_1876,N_1663);
nand U3255 (N_3255,N_2294,N_2617);
or U3256 (N_3256,N_2672,N_2953);
nor U3257 (N_3257,N_2796,N_1648);
or U3258 (N_3258,N_2076,N_2202);
and U3259 (N_3259,N_2541,N_2946);
and U3260 (N_3260,N_1734,N_2025);
or U3261 (N_3261,N_1621,N_2585);
nand U3262 (N_3262,N_2578,N_2309);
and U3263 (N_3263,N_2406,N_2048);
or U3264 (N_3264,N_1866,N_1604);
xnor U3265 (N_3265,N_2854,N_2207);
or U3266 (N_3266,N_2859,N_2997);
and U3267 (N_3267,N_1675,N_2603);
or U3268 (N_3268,N_1718,N_2844);
and U3269 (N_3269,N_1690,N_2855);
or U3270 (N_3270,N_2951,N_2677);
xor U3271 (N_3271,N_2934,N_2639);
nand U3272 (N_3272,N_2003,N_1846);
nor U3273 (N_3273,N_2042,N_2960);
or U3274 (N_3274,N_2930,N_2209);
nor U3275 (N_3275,N_2839,N_2723);
nand U3276 (N_3276,N_1724,N_1783);
or U3277 (N_3277,N_1600,N_2090);
nand U3278 (N_3278,N_2529,N_2063);
nand U3279 (N_3279,N_2073,N_1633);
nand U3280 (N_3280,N_2468,N_2137);
and U3281 (N_3281,N_1727,N_1939);
and U3282 (N_3282,N_1700,N_2106);
nand U3283 (N_3283,N_2443,N_1568);
nor U3284 (N_3284,N_2391,N_2852);
xor U3285 (N_3285,N_2160,N_1822);
nand U3286 (N_3286,N_2159,N_2065);
nand U3287 (N_3287,N_2357,N_2907);
and U3288 (N_3288,N_2504,N_2885);
or U3289 (N_3289,N_2903,N_2631);
or U3290 (N_3290,N_1680,N_2327);
and U3291 (N_3291,N_2474,N_2236);
nand U3292 (N_3292,N_2153,N_1620);
nand U3293 (N_3293,N_1617,N_1728);
or U3294 (N_3294,N_2475,N_2331);
or U3295 (N_3295,N_2388,N_2740);
nor U3296 (N_3296,N_2594,N_1752);
nor U3297 (N_3297,N_2398,N_2511);
nand U3298 (N_3298,N_2359,N_2318);
or U3299 (N_3299,N_2998,N_1555);
nand U3300 (N_3300,N_2992,N_2922);
nand U3301 (N_3301,N_2224,N_2011);
nand U3302 (N_3302,N_2755,N_2593);
xnor U3303 (N_3303,N_2061,N_2817);
nor U3304 (N_3304,N_2862,N_2806);
nor U3305 (N_3305,N_1658,N_2765);
nor U3306 (N_3306,N_2098,N_1571);
or U3307 (N_3307,N_1652,N_1959);
nor U3308 (N_3308,N_2064,N_2931);
nor U3309 (N_3309,N_1818,N_1699);
and U3310 (N_3310,N_2823,N_2727);
xnor U3311 (N_3311,N_2456,N_2487);
and U3312 (N_3312,N_2490,N_1748);
nand U3313 (N_3313,N_1881,N_2149);
nand U3314 (N_3314,N_1596,N_1585);
nor U3315 (N_3315,N_2006,N_1929);
xnor U3316 (N_3316,N_1686,N_1828);
or U3317 (N_3317,N_1778,N_2717);
and U3318 (N_3318,N_2129,N_2198);
and U3319 (N_3319,N_1601,N_2658);
nand U3320 (N_3320,N_1812,N_2241);
nand U3321 (N_3321,N_2660,N_2000);
nand U3322 (N_3322,N_2441,N_1964);
nor U3323 (N_3323,N_2104,N_1969);
and U3324 (N_3324,N_2974,N_1721);
nor U3325 (N_3325,N_2176,N_1998);
or U3326 (N_3326,N_2007,N_2670);
xor U3327 (N_3327,N_2182,N_2485);
nor U3328 (N_3328,N_2540,N_1665);
and U3329 (N_3329,N_2971,N_2125);
nand U3330 (N_3330,N_2029,N_2329);
or U3331 (N_3331,N_1549,N_2949);
and U3332 (N_3332,N_2663,N_1697);
and U3333 (N_3333,N_1970,N_2426);
or U3334 (N_3334,N_1667,N_1503);
or U3335 (N_3335,N_1777,N_2702);
and U3336 (N_3336,N_1993,N_2158);
and U3337 (N_3337,N_1643,N_2033);
and U3338 (N_3338,N_2257,N_2712);
nand U3339 (N_3339,N_2899,N_1716);
nand U3340 (N_3340,N_1759,N_2635);
nand U3341 (N_3341,N_1820,N_2284);
nor U3342 (N_3342,N_2657,N_1834);
nor U3343 (N_3343,N_2872,N_1854);
or U3344 (N_3344,N_2085,N_2983);
and U3345 (N_3345,N_2277,N_1770);
nor U3346 (N_3346,N_2086,N_2119);
or U3347 (N_3347,N_2668,N_2306);
nand U3348 (N_3348,N_1726,N_2030);
nor U3349 (N_3349,N_2449,N_1983);
xor U3350 (N_3350,N_2661,N_2138);
nand U3351 (N_3351,N_2703,N_2652);
nor U3352 (N_3352,N_2664,N_2135);
or U3353 (N_3353,N_1730,N_1764);
nor U3354 (N_3354,N_2122,N_2004);
nand U3355 (N_3355,N_2349,N_1879);
nor U3356 (N_3356,N_1735,N_1672);
or U3357 (N_3357,N_1862,N_2532);
nor U3358 (N_3358,N_1989,N_1682);
and U3359 (N_3359,N_2711,N_2786);
nand U3360 (N_3360,N_2856,N_1968);
or U3361 (N_3361,N_1509,N_1806);
or U3362 (N_3362,N_2328,N_1671);
nor U3363 (N_3363,N_1739,N_2726);
and U3364 (N_3364,N_2643,N_2184);
or U3365 (N_3365,N_2163,N_2013);
and U3366 (N_3366,N_2193,N_1938);
or U3367 (N_3367,N_1944,N_1860);
or U3368 (N_3368,N_1581,N_2621);
nand U3369 (N_3369,N_2731,N_2244);
nor U3370 (N_3370,N_1933,N_2730);
nand U3371 (N_3371,N_2679,N_2902);
nand U3372 (N_3372,N_2131,N_2127);
nor U3373 (N_3373,N_2601,N_2445);
nor U3374 (N_3374,N_2337,N_2354);
and U3375 (N_3375,N_2954,N_1586);
nor U3376 (N_3376,N_1814,N_2581);
or U3377 (N_3377,N_2613,N_2616);
and U3378 (N_3378,N_1827,N_2077);
nor U3379 (N_3379,N_1688,N_2572);
nand U3380 (N_3380,N_2145,N_2392);
nor U3381 (N_3381,N_2341,N_2231);
nand U3382 (N_3382,N_2014,N_2513);
and U3383 (N_3383,N_2995,N_2596);
or U3384 (N_3384,N_1997,N_1504);
xnor U3385 (N_3385,N_2857,N_2574);
or U3386 (N_3386,N_2133,N_2446);
nor U3387 (N_3387,N_2253,N_2502);
nor U3388 (N_3388,N_2422,N_2586);
or U3389 (N_3389,N_1744,N_2656);
and U3390 (N_3390,N_2455,N_2659);
and U3391 (N_3391,N_2560,N_1754);
or U3392 (N_3392,N_2174,N_2945);
or U3393 (N_3393,N_2769,N_1693);
or U3394 (N_3394,N_2440,N_2430);
nor U3395 (N_3395,N_1769,N_1932);
nand U3396 (N_3396,N_2461,N_2320);
nor U3397 (N_3397,N_2675,N_1654);
nand U3398 (N_3398,N_2211,N_2097);
and U3399 (N_3399,N_2925,N_2684);
nor U3400 (N_3400,N_2826,N_2988);
and U3401 (N_3401,N_2419,N_2993);
or U3402 (N_3402,N_2897,N_2412);
and U3403 (N_3403,N_2201,N_1960);
nor U3404 (N_3404,N_2632,N_1709);
nor U3405 (N_3405,N_2813,N_2084);
nand U3406 (N_3406,N_2627,N_2346);
nand U3407 (N_3407,N_2705,N_2793);
and U3408 (N_3408,N_2370,N_1903);
or U3409 (N_3409,N_1542,N_1723);
nand U3410 (N_3410,N_1507,N_2634);
nor U3411 (N_3411,N_2869,N_2519);
and U3412 (N_3412,N_2733,N_2259);
nand U3413 (N_3413,N_1979,N_1816);
and U3414 (N_3414,N_2165,N_2278);
or U3415 (N_3415,N_2283,N_2043);
or U3416 (N_3416,N_1784,N_2523);
and U3417 (N_3417,N_2314,N_2301);
and U3418 (N_3418,N_2046,N_1908);
nor U3419 (N_3419,N_1880,N_2353);
nor U3420 (N_3420,N_1975,N_1746);
xnor U3421 (N_3421,N_2963,N_2285);
or U3422 (N_3422,N_2570,N_2824);
nor U3423 (N_3423,N_2371,N_2503);
or U3424 (N_3424,N_2901,N_2846);
or U3425 (N_3425,N_2534,N_1914);
and U3426 (N_3426,N_1955,N_2630);
nand U3427 (N_3427,N_2732,N_1882);
or U3428 (N_3428,N_2875,N_2561);
nand U3429 (N_3429,N_1567,N_2427);
and U3430 (N_3430,N_1990,N_2054);
nand U3431 (N_3431,N_2081,N_1790);
and U3432 (N_3432,N_2303,N_1872);
nand U3433 (N_3433,N_2673,N_2536);
nor U3434 (N_3434,N_2790,N_2553);
and U3435 (N_3435,N_2360,N_2776);
nand U3436 (N_3436,N_1587,N_2548);
xor U3437 (N_3437,N_1570,N_1564);
or U3438 (N_3438,N_1954,N_2648);
or U3439 (N_3439,N_1603,N_2471);
and U3440 (N_3440,N_2947,N_2797);
and U3441 (N_3441,N_2800,N_2340);
or U3442 (N_3442,N_1529,N_2146);
nand U3443 (N_3443,N_2956,N_1949);
or U3444 (N_3444,N_2154,N_2372);
and U3445 (N_3445,N_2212,N_2142);
or U3446 (N_3446,N_2943,N_2920);
or U3447 (N_3447,N_1865,N_2939);
or U3448 (N_3448,N_1847,N_2290);
nor U3449 (N_3449,N_2386,N_2768);
or U3450 (N_3450,N_1640,N_1785);
nand U3451 (N_3451,N_1687,N_2942);
nor U3452 (N_3452,N_1850,N_1928);
nor U3453 (N_3453,N_1588,N_2269);
or U3454 (N_3454,N_1936,N_1523);
and U3455 (N_3455,N_1522,N_2926);
or U3456 (N_3456,N_2607,N_1685);
xnor U3457 (N_3457,N_2750,N_1953);
nor U3458 (N_3458,N_2336,N_2092);
nor U3459 (N_3459,N_1813,N_2512);
nor U3460 (N_3460,N_1520,N_2531);
nor U3461 (N_3461,N_2087,N_1945);
nand U3462 (N_3462,N_2720,N_2555);
nand U3463 (N_3463,N_1642,N_2102);
nand U3464 (N_3464,N_2265,N_2267);
or U3465 (N_3465,N_2344,N_1910);
nand U3466 (N_3466,N_2987,N_2271);
xor U3467 (N_3467,N_2476,N_2113);
or U3468 (N_3468,N_1614,N_2688);
nor U3469 (N_3469,N_2191,N_1646);
nand U3470 (N_3470,N_1526,N_1573);
nand U3471 (N_3471,N_2215,N_2024);
and U3472 (N_3472,N_2683,N_2990);
or U3473 (N_3473,N_2095,N_2457);
or U3474 (N_3474,N_2175,N_1973);
or U3475 (N_3475,N_2423,N_1532);
or U3476 (N_3476,N_2079,N_2501);
and U3477 (N_3477,N_2772,N_2589);
and U3478 (N_3478,N_2075,N_1565);
and U3479 (N_3479,N_2438,N_1630);
and U3480 (N_3480,N_2845,N_2521);
or U3481 (N_3481,N_2980,N_2773);
and U3482 (N_3482,N_1841,N_2197);
nor U3483 (N_3483,N_2904,N_1950);
or U3484 (N_3484,N_2996,N_2693);
xor U3485 (N_3485,N_2204,N_2275);
and U3486 (N_3486,N_2792,N_2316);
xnor U3487 (N_3487,N_1627,N_2034);
and U3488 (N_3488,N_2274,N_2568);
nor U3489 (N_3489,N_2107,N_2260);
nand U3490 (N_3490,N_2496,N_1775);
nor U3491 (N_3491,N_2986,N_1609);
and U3492 (N_3492,N_2400,N_1619);
and U3493 (N_3493,N_1838,N_1794);
nand U3494 (N_3494,N_2334,N_2893);
nor U3495 (N_3495,N_2811,N_1711);
or U3496 (N_3496,N_2784,N_1957);
or U3497 (N_3497,N_1750,N_2602);
nor U3498 (N_3498,N_2972,N_1819);
xor U3499 (N_3499,N_1982,N_2751);
or U3500 (N_3500,N_2484,N_1756);
and U3501 (N_3501,N_2879,N_2842);
nor U3502 (N_3502,N_1692,N_1809);
nand U3503 (N_3503,N_2725,N_1771);
nand U3504 (N_3504,N_2429,N_2167);
or U3505 (N_3505,N_2644,N_1888);
nand U3506 (N_3506,N_2685,N_2152);
and U3507 (N_3507,N_1527,N_2348);
and U3508 (N_3508,N_1951,N_1577);
nand U3509 (N_3509,N_2978,N_2071);
xor U3510 (N_3510,N_2108,N_2952);
nor U3511 (N_3511,N_2005,N_2888);
and U3512 (N_3512,N_2729,N_1829);
or U3513 (N_3513,N_2690,N_2936);
and U3514 (N_3514,N_2687,N_2597);
nand U3515 (N_3515,N_2464,N_1845);
or U3516 (N_3516,N_2940,N_2984);
and U3517 (N_3517,N_2074,N_2478);
and U3518 (N_3518,N_1943,N_2345);
nor U3519 (N_3519,N_2433,N_1831);
and U3520 (N_3520,N_2932,N_1556);
xor U3521 (N_3521,N_2637,N_2821);
and U3522 (N_3522,N_2771,N_2068);
nand U3523 (N_3523,N_2428,N_2691);
or U3524 (N_3524,N_1576,N_1710);
xnor U3525 (N_3525,N_2052,N_2038);
xnor U3526 (N_3526,N_2028,N_1952);
nor U3527 (N_3527,N_1704,N_1714);
or U3528 (N_3528,N_1701,N_2056);
and U3529 (N_3529,N_1650,N_2319);
xor U3530 (N_3530,N_2040,N_2124);
nand U3531 (N_3531,N_2332,N_1780);
or U3532 (N_3532,N_2242,N_2666);
xor U3533 (N_3533,N_2292,N_2270);
nor U3534 (N_3534,N_2724,N_2871);
xnor U3535 (N_3535,N_2841,N_2199);
or U3536 (N_3536,N_2390,N_2746);
and U3537 (N_3537,N_1713,N_2009);
or U3538 (N_3538,N_2444,N_2100);
nor U3539 (N_3539,N_1737,N_1799);
nand U3540 (N_3540,N_2834,N_2563);
nand U3541 (N_3541,N_1884,N_2194);
and U3542 (N_3542,N_2741,N_1541);
nor U3543 (N_3543,N_2335,N_2080);
or U3544 (N_3544,N_1517,N_2424);
nor U3545 (N_3545,N_2609,N_1886);
nor U3546 (N_3546,N_1705,N_1538);
and U3547 (N_3547,N_2498,N_2403);
nand U3548 (N_3548,N_2567,N_1572);
nor U3549 (N_3549,N_2655,N_1774);
xnor U3550 (N_3550,N_2582,N_1758);
or U3551 (N_3551,N_2062,N_1607);
nand U3552 (N_3552,N_2520,N_2408);
nor U3553 (N_3553,N_2117,N_1731);
or U3554 (N_3554,N_2791,N_2118);
or U3555 (N_3555,N_2533,N_1922);
xor U3556 (N_3556,N_2539,N_2819);
nand U3557 (N_3557,N_1980,N_1597);
or U3558 (N_3558,N_1895,N_2849);
nand U3559 (N_3559,N_2173,N_2605);
nand U3560 (N_3560,N_2966,N_2351);
and U3561 (N_3561,N_2767,N_1679);
xor U3562 (N_3562,N_2302,N_2266);
nand U3563 (N_3563,N_2049,N_1892);
and U3564 (N_3564,N_2584,N_1976);
nand U3565 (N_3565,N_1592,N_2223);
nor U3566 (N_3566,N_2078,N_1853);
and U3567 (N_3567,N_2779,N_2171);
nor U3568 (N_3568,N_2369,N_2238);
or U3569 (N_3569,N_1967,N_1519);
xor U3570 (N_3570,N_1539,N_2547);
xor U3571 (N_3571,N_2164,N_1767);
and U3572 (N_3572,N_2756,N_2546);
and U3573 (N_3573,N_2787,N_2874);
and U3574 (N_3574,N_2837,N_2172);
xnor U3575 (N_3575,N_2288,N_1839);
xor U3576 (N_3576,N_2970,N_2286);
nor U3577 (N_3577,N_2472,N_2413);
nor U3578 (N_3578,N_2645,N_1927);
and U3579 (N_3579,N_2096,N_1702);
nand U3580 (N_3580,N_2738,N_2840);
or U3581 (N_3581,N_2366,N_1902);
and U3582 (N_3582,N_1530,N_2650);
or U3583 (N_3583,N_2507,N_1836);
or U3584 (N_3584,N_2217,N_2114);
and U3585 (N_3585,N_1916,N_2600);
and U3586 (N_3586,N_2745,N_2082);
or U3587 (N_3587,N_2695,N_2694);
or U3588 (N_3588,N_2467,N_1751);
nand U3589 (N_3589,N_2330,N_2317);
nand U3590 (N_3590,N_2214,N_2843);
nand U3591 (N_3591,N_2367,N_2915);
and U3592 (N_3592,N_2208,N_2256);
nand U3593 (N_3593,N_1772,N_2032);
nor U3594 (N_3594,N_1524,N_1795);
or U3595 (N_3595,N_1732,N_1907);
and U3596 (N_3596,N_2035,N_1664);
or U3597 (N_3597,N_1878,N_2590);
and U3598 (N_3598,N_1528,N_2912);
or U3599 (N_3599,N_2782,N_2524);
nand U3600 (N_3600,N_2580,N_1849);
nand U3601 (N_3601,N_2379,N_2774);
nor U3602 (N_3602,N_2315,N_2911);
xor U3603 (N_3603,N_2010,N_2937);
nor U3604 (N_3604,N_1987,N_2132);
nor U3605 (N_3605,N_2295,N_1512);
nor U3606 (N_3606,N_2718,N_2393);
nand U3607 (N_3607,N_1913,N_2243);
or U3608 (N_3608,N_2110,N_2919);
nand U3609 (N_3609,N_2489,N_2465);
nor U3610 (N_3610,N_1869,N_2638);
nand U3611 (N_3611,N_2598,N_1786);
nand U3612 (N_3612,N_2770,N_1677);
or U3613 (N_3613,N_2234,N_1789);
and U3614 (N_3614,N_2023,N_2880);
and U3615 (N_3615,N_2434,N_2882);
nor U3616 (N_3616,N_1883,N_1653);
and U3617 (N_3617,N_2558,N_2383);
xor U3618 (N_3618,N_1889,N_2667);
nand U3619 (N_3619,N_2222,N_2822);
nand U3620 (N_3620,N_2759,N_2889);
nand U3621 (N_3621,N_2247,N_1901);
and U3622 (N_3622,N_2647,N_2479);
nor U3623 (N_3623,N_2059,N_2929);
nand U3624 (N_3624,N_2297,N_2482);
or U3625 (N_3625,N_2252,N_2735);
nor U3626 (N_3626,N_1787,N_2808);
nor U3627 (N_3627,N_2692,N_1632);
nor U3628 (N_3628,N_2280,N_2734);
nand U3629 (N_3629,N_2213,N_1674);
nand U3630 (N_3630,N_1594,N_2189);
nor U3631 (N_3631,N_1639,N_1808);
nand U3632 (N_3632,N_1974,N_1698);
and U3633 (N_3633,N_2183,N_1986);
and U3634 (N_3634,N_1811,N_2713);
and U3635 (N_3635,N_2019,N_2389);
and U3636 (N_3636,N_1651,N_2459);
and U3637 (N_3637,N_1867,N_2599);
nand U3638 (N_3638,N_2577,N_2704);
nand U3639 (N_3639,N_1662,N_2700);
nand U3640 (N_3640,N_1826,N_2477);
or U3641 (N_3641,N_2166,N_2055);
nand U3642 (N_3642,N_1906,N_2747);
and U3643 (N_3643,N_1584,N_2326);
xnor U3644 (N_3644,N_2447,N_1608);
nand U3645 (N_3645,N_2569,N_2615);
and U3646 (N_3646,N_1745,N_2575);
nor U3647 (N_3647,N_1501,N_2181);
and U3648 (N_3648,N_2982,N_2120);
and U3649 (N_3649,N_2263,N_1905);
or U3650 (N_3650,N_1891,N_1830);
nand U3651 (N_3651,N_1610,N_1525);
and U3652 (N_3652,N_2439,N_2545);
or U3653 (N_3653,N_2394,N_1815);
or U3654 (N_3654,N_1935,N_2069);
and U3655 (N_3655,N_2697,N_2192);
xnor U3656 (N_3656,N_2778,N_2562);
nand U3657 (N_3657,N_2968,N_1926);
nand U3658 (N_3658,N_2493,N_1917);
or U3659 (N_3659,N_1885,N_2499);
nand U3660 (N_3660,N_2083,N_1531);
xor U3661 (N_3661,N_2651,N_2636);
and U3662 (N_3662,N_1659,N_1715);
nor U3663 (N_3663,N_2763,N_1557);
nor U3664 (N_3664,N_2017,N_2923);
nor U3665 (N_3665,N_1920,N_2264);
nor U3666 (N_3666,N_1562,N_1896);
or U3667 (N_3667,N_1842,N_2516);
and U3668 (N_3668,N_1755,N_2311);
nor U3669 (N_3669,N_2358,N_1580);
xnor U3670 (N_3670,N_1544,N_1937);
nand U3671 (N_3671,N_1725,N_2979);
or U3672 (N_3672,N_2608,N_1551);
and U3673 (N_3673,N_2965,N_1591);
nor U3674 (N_3674,N_2827,N_1796);
and U3675 (N_3675,N_2884,N_2795);
nand U3676 (N_3676,N_1707,N_2958);
and U3677 (N_3677,N_2909,N_2155);
or U3678 (N_3678,N_1612,N_2948);
and U3679 (N_3679,N_2515,N_2506);
nand U3680 (N_3680,N_2324,N_2719);
and U3681 (N_3681,N_2103,N_1534);
or U3682 (N_3682,N_2180,N_2816);
nand U3683 (N_3683,N_1992,N_1873);
nand U3684 (N_3684,N_1510,N_2528);
nand U3685 (N_3685,N_2914,N_2870);
xor U3686 (N_3686,N_2535,N_1712);
nand U3687 (N_3687,N_2873,N_2050);
xnor U3688 (N_3688,N_1719,N_1864);
and U3689 (N_3689,N_2955,N_2109);
nor U3690 (N_3690,N_2307,N_1511);
or U3691 (N_3691,N_2739,N_1947);
nor U3692 (N_3692,N_1977,N_1988);
and U3693 (N_3693,N_2219,N_2860);
nand U3694 (N_3694,N_2148,N_1578);
nand U3695 (N_3695,N_2308,N_2402);
or U3696 (N_3696,N_1740,N_1615);
or U3697 (N_3697,N_1629,N_1946);
or U3698 (N_3698,N_1535,N_2323);
or U3699 (N_3699,N_2417,N_1893);
or U3700 (N_3700,N_2868,N_1837);
and U3701 (N_3701,N_2964,N_2810);
nand U3702 (N_3702,N_2706,N_2680);
xor U3703 (N_3703,N_1606,N_1788);
and U3704 (N_3704,N_2858,N_2141);
nor U3705 (N_3705,N_2975,N_1681);
nand U3706 (N_3706,N_1605,N_2448);
or U3707 (N_3707,N_2928,N_2044);
or U3708 (N_3708,N_2190,N_1670);
nand U3709 (N_3709,N_2200,N_1566);
nor U3710 (N_3710,N_2544,N_2716);
and U3711 (N_3711,N_2973,N_1647);
nor U3712 (N_3712,N_2342,N_1548);
nand U3713 (N_3713,N_2136,N_2714);
and U3714 (N_3714,N_2218,N_1695);
and U3715 (N_3715,N_2804,N_2564);
nor U3716 (N_3716,N_2401,N_2828);
nor U3717 (N_3717,N_2595,N_2442);
nand U3718 (N_3718,N_2579,N_1797);
nand U3719 (N_3719,N_2510,N_1583);
nand U3720 (N_3720,N_2707,N_2671);
nand U3721 (N_3721,N_2917,N_2905);
nand U3722 (N_3722,N_2805,N_1743);
nor U3723 (N_3723,N_2147,N_2368);
nor U3724 (N_3724,N_2361,N_1823);
or U3725 (N_3725,N_2748,N_2452);
nor U3726 (N_3726,N_1742,N_1909);
nor U3727 (N_3727,N_1626,N_2500);
nand U3728 (N_3728,N_2836,N_2861);
xor U3729 (N_3729,N_2469,N_2881);
xnor U3730 (N_3730,N_1720,N_2333);
nand U3731 (N_3731,N_1657,N_2435);
or U3732 (N_3732,N_2527,N_1972);
or U3733 (N_3733,N_2832,N_2509);
xor U3734 (N_3734,N_2641,N_1595);
nor U3735 (N_3735,N_2927,N_2742);
nand U3736 (N_3736,N_2542,N_2785);
xor U3737 (N_3737,N_2273,N_2910);
or U3738 (N_3738,N_2458,N_2041);
nor U3739 (N_3739,N_1870,N_2967);
nand U3740 (N_3740,N_2365,N_1923);
nor U3741 (N_3741,N_2338,N_2892);
nand U3742 (N_3742,N_2460,N_1689);
and U3743 (N_3743,N_2179,N_2757);
nor U3744 (N_3744,N_2099,N_2894);
xor U3745 (N_3745,N_2374,N_2088);
nand U3746 (N_3746,N_2662,N_1598);
and U3747 (N_3747,N_2415,N_1782);
and U3748 (N_3748,N_1513,N_2436);
nor U3749 (N_3749,N_1508,N_2139);
and U3750 (N_3750,N_2518,N_2982);
nor U3751 (N_3751,N_1604,N_2569);
nor U3752 (N_3752,N_2442,N_1829);
and U3753 (N_3753,N_2069,N_2461);
nor U3754 (N_3754,N_2370,N_2129);
xor U3755 (N_3755,N_2784,N_2849);
nand U3756 (N_3756,N_2982,N_2467);
and U3757 (N_3757,N_1550,N_1589);
and U3758 (N_3758,N_2025,N_2960);
xor U3759 (N_3759,N_2261,N_2050);
nand U3760 (N_3760,N_1673,N_2439);
or U3761 (N_3761,N_2739,N_1709);
and U3762 (N_3762,N_1634,N_2089);
nor U3763 (N_3763,N_2268,N_2407);
or U3764 (N_3764,N_1899,N_2258);
or U3765 (N_3765,N_1758,N_2648);
nand U3766 (N_3766,N_2866,N_1683);
nand U3767 (N_3767,N_2062,N_1987);
nand U3768 (N_3768,N_2138,N_2890);
nand U3769 (N_3769,N_2980,N_2765);
or U3770 (N_3770,N_2474,N_1702);
or U3771 (N_3771,N_2266,N_1746);
and U3772 (N_3772,N_2662,N_2058);
xor U3773 (N_3773,N_2110,N_1594);
nand U3774 (N_3774,N_1960,N_1882);
or U3775 (N_3775,N_1929,N_2395);
and U3776 (N_3776,N_1888,N_2412);
nand U3777 (N_3777,N_2962,N_2383);
or U3778 (N_3778,N_2888,N_2651);
nand U3779 (N_3779,N_1977,N_2646);
nor U3780 (N_3780,N_1533,N_2994);
or U3781 (N_3781,N_2748,N_2639);
or U3782 (N_3782,N_2736,N_1943);
and U3783 (N_3783,N_2686,N_1710);
or U3784 (N_3784,N_2711,N_2488);
and U3785 (N_3785,N_2500,N_2812);
xor U3786 (N_3786,N_2364,N_2831);
and U3787 (N_3787,N_1549,N_2891);
and U3788 (N_3788,N_1772,N_1546);
and U3789 (N_3789,N_2513,N_2522);
nor U3790 (N_3790,N_2320,N_2965);
or U3791 (N_3791,N_2491,N_2389);
nand U3792 (N_3792,N_2144,N_2671);
or U3793 (N_3793,N_1981,N_1607);
nor U3794 (N_3794,N_1541,N_1920);
nor U3795 (N_3795,N_2129,N_2288);
nor U3796 (N_3796,N_2974,N_1749);
xnor U3797 (N_3797,N_2696,N_2614);
nand U3798 (N_3798,N_2039,N_2120);
nand U3799 (N_3799,N_2038,N_1778);
and U3800 (N_3800,N_1614,N_2559);
nor U3801 (N_3801,N_1663,N_2070);
or U3802 (N_3802,N_2684,N_2780);
nand U3803 (N_3803,N_2214,N_2690);
or U3804 (N_3804,N_1962,N_2552);
nand U3805 (N_3805,N_2128,N_2276);
and U3806 (N_3806,N_2585,N_1775);
nand U3807 (N_3807,N_2963,N_2083);
and U3808 (N_3808,N_1716,N_2284);
or U3809 (N_3809,N_1858,N_1629);
or U3810 (N_3810,N_2226,N_2152);
nor U3811 (N_3811,N_1768,N_2893);
and U3812 (N_3812,N_1916,N_2757);
nand U3813 (N_3813,N_2431,N_2777);
or U3814 (N_3814,N_2923,N_2110);
or U3815 (N_3815,N_2681,N_1973);
nand U3816 (N_3816,N_1838,N_1996);
xnor U3817 (N_3817,N_2008,N_2537);
nor U3818 (N_3818,N_2181,N_2115);
xor U3819 (N_3819,N_2312,N_2210);
nand U3820 (N_3820,N_1984,N_2305);
xor U3821 (N_3821,N_1501,N_2145);
nor U3822 (N_3822,N_1894,N_2831);
nor U3823 (N_3823,N_1804,N_2352);
nand U3824 (N_3824,N_2039,N_2568);
or U3825 (N_3825,N_2393,N_2429);
nand U3826 (N_3826,N_1996,N_1752);
nor U3827 (N_3827,N_1614,N_2393);
and U3828 (N_3828,N_1511,N_2638);
nand U3829 (N_3829,N_1524,N_2717);
and U3830 (N_3830,N_1813,N_1885);
and U3831 (N_3831,N_1549,N_1710);
nor U3832 (N_3832,N_2614,N_2305);
nand U3833 (N_3833,N_2376,N_2303);
or U3834 (N_3834,N_2094,N_2690);
or U3835 (N_3835,N_1848,N_2273);
and U3836 (N_3836,N_2083,N_2329);
or U3837 (N_3837,N_2113,N_1643);
or U3838 (N_3838,N_2350,N_2662);
or U3839 (N_3839,N_2529,N_2815);
nor U3840 (N_3840,N_2246,N_2186);
nand U3841 (N_3841,N_2058,N_1665);
or U3842 (N_3842,N_2781,N_2504);
nand U3843 (N_3843,N_1812,N_2286);
xor U3844 (N_3844,N_2995,N_1875);
or U3845 (N_3845,N_1749,N_2011);
or U3846 (N_3846,N_1717,N_2502);
nand U3847 (N_3847,N_2659,N_2069);
and U3848 (N_3848,N_1690,N_2791);
and U3849 (N_3849,N_2911,N_2542);
and U3850 (N_3850,N_2513,N_2241);
nor U3851 (N_3851,N_1564,N_1806);
or U3852 (N_3852,N_2551,N_1708);
nor U3853 (N_3853,N_1691,N_2802);
nand U3854 (N_3854,N_2867,N_2950);
nor U3855 (N_3855,N_2926,N_2599);
nand U3856 (N_3856,N_2418,N_2688);
and U3857 (N_3857,N_2865,N_1793);
xor U3858 (N_3858,N_1900,N_1522);
and U3859 (N_3859,N_2725,N_2344);
nand U3860 (N_3860,N_1547,N_2026);
nand U3861 (N_3861,N_2175,N_2318);
nand U3862 (N_3862,N_1605,N_2357);
and U3863 (N_3863,N_1544,N_2849);
or U3864 (N_3864,N_1773,N_2060);
or U3865 (N_3865,N_2306,N_2385);
and U3866 (N_3866,N_2073,N_2484);
or U3867 (N_3867,N_1936,N_2987);
nand U3868 (N_3868,N_1746,N_1792);
nor U3869 (N_3869,N_1936,N_2902);
and U3870 (N_3870,N_2656,N_1508);
or U3871 (N_3871,N_2199,N_1728);
and U3872 (N_3872,N_1780,N_1870);
nand U3873 (N_3873,N_2014,N_1660);
or U3874 (N_3874,N_1924,N_1856);
xnor U3875 (N_3875,N_2050,N_2591);
and U3876 (N_3876,N_2140,N_2016);
nand U3877 (N_3877,N_1782,N_2336);
xor U3878 (N_3878,N_1883,N_2591);
nor U3879 (N_3879,N_2138,N_2583);
and U3880 (N_3880,N_2979,N_2293);
nand U3881 (N_3881,N_2827,N_1555);
nand U3882 (N_3882,N_1503,N_2810);
nor U3883 (N_3883,N_2746,N_2963);
nor U3884 (N_3884,N_1880,N_2412);
and U3885 (N_3885,N_2182,N_2930);
nor U3886 (N_3886,N_1683,N_2492);
xnor U3887 (N_3887,N_2099,N_1810);
xor U3888 (N_3888,N_2435,N_2326);
xor U3889 (N_3889,N_2827,N_2152);
or U3890 (N_3890,N_2580,N_1759);
nand U3891 (N_3891,N_1881,N_2912);
or U3892 (N_3892,N_2669,N_2601);
xor U3893 (N_3893,N_1979,N_1975);
or U3894 (N_3894,N_2042,N_2629);
xnor U3895 (N_3895,N_1891,N_1695);
nor U3896 (N_3896,N_2485,N_2737);
nand U3897 (N_3897,N_2870,N_2734);
nor U3898 (N_3898,N_1840,N_2330);
nand U3899 (N_3899,N_2102,N_2504);
nand U3900 (N_3900,N_2855,N_1927);
xnor U3901 (N_3901,N_1625,N_1553);
and U3902 (N_3902,N_1643,N_2056);
and U3903 (N_3903,N_1737,N_2953);
and U3904 (N_3904,N_2628,N_2727);
nand U3905 (N_3905,N_2322,N_2426);
and U3906 (N_3906,N_1834,N_2559);
nand U3907 (N_3907,N_2686,N_2439);
nand U3908 (N_3908,N_2790,N_2992);
nor U3909 (N_3909,N_1651,N_2013);
or U3910 (N_3910,N_2692,N_1728);
nor U3911 (N_3911,N_2943,N_2267);
nand U3912 (N_3912,N_2836,N_2152);
and U3913 (N_3913,N_1720,N_2215);
xnor U3914 (N_3914,N_1602,N_2592);
or U3915 (N_3915,N_2019,N_2591);
xor U3916 (N_3916,N_1502,N_2089);
nand U3917 (N_3917,N_2391,N_2053);
nor U3918 (N_3918,N_2234,N_1904);
and U3919 (N_3919,N_2156,N_2210);
xor U3920 (N_3920,N_2493,N_2467);
nor U3921 (N_3921,N_1526,N_2774);
xnor U3922 (N_3922,N_2252,N_2003);
nand U3923 (N_3923,N_1652,N_1607);
or U3924 (N_3924,N_2168,N_2858);
and U3925 (N_3925,N_1661,N_1709);
and U3926 (N_3926,N_2593,N_1706);
and U3927 (N_3927,N_2349,N_2264);
or U3928 (N_3928,N_2793,N_2569);
nor U3929 (N_3929,N_1968,N_2356);
xnor U3930 (N_3930,N_2053,N_1785);
and U3931 (N_3931,N_2781,N_2540);
nor U3932 (N_3932,N_2764,N_2789);
nor U3933 (N_3933,N_2165,N_2985);
nand U3934 (N_3934,N_1843,N_1786);
nand U3935 (N_3935,N_2776,N_2890);
nor U3936 (N_3936,N_1595,N_2943);
and U3937 (N_3937,N_2337,N_2822);
nor U3938 (N_3938,N_1877,N_2238);
nor U3939 (N_3939,N_2676,N_2352);
xor U3940 (N_3940,N_2566,N_1935);
nor U3941 (N_3941,N_1774,N_2858);
nor U3942 (N_3942,N_1818,N_2959);
nand U3943 (N_3943,N_2394,N_1809);
and U3944 (N_3944,N_1575,N_2858);
nand U3945 (N_3945,N_2615,N_2544);
nor U3946 (N_3946,N_1572,N_1664);
or U3947 (N_3947,N_1692,N_2796);
nand U3948 (N_3948,N_1939,N_1839);
and U3949 (N_3949,N_2085,N_1698);
nand U3950 (N_3950,N_1593,N_2215);
and U3951 (N_3951,N_2998,N_2796);
xor U3952 (N_3952,N_2996,N_1915);
and U3953 (N_3953,N_2359,N_2254);
and U3954 (N_3954,N_2584,N_1815);
nand U3955 (N_3955,N_1517,N_2999);
xor U3956 (N_3956,N_1557,N_2698);
nand U3957 (N_3957,N_2526,N_1960);
and U3958 (N_3958,N_2512,N_2331);
nand U3959 (N_3959,N_1915,N_2083);
and U3960 (N_3960,N_2971,N_2826);
xnor U3961 (N_3961,N_2403,N_2043);
or U3962 (N_3962,N_1615,N_2885);
and U3963 (N_3963,N_2397,N_2670);
nand U3964 (N_3964,N_2109,N_2852);
nand U3965 (N_3965,N_2892,N_2461);
or U3966 (N_3966,N_1676,N_1825);
xor U3967 (N_3967,N_1577,N_1735);
xnor U3968 (N_3968,N_2069,N_2201);
nor U3969 (N_3969,N_2937,N_2282);
or U3970 (N_3970,N_1748,N_2277);
or U3971 (N_3971,N_2967,N_2165);
or U3972 (N_3972,N_2116,N_1864);
or U3973 (N_3973,N_2437,N_2971);
or U3974 (N_3974,N_2957,N_1892);
nor U3975 (N_3975,N_1559,N_2459);
and U3976 (N_3976,N_2163,N_2499);
nand U3977 (N_3977,N_2945,N_1501);
nand U3978 (N_3978,N_2703,N_2540);
nor U3979 (N_3979,N_1500,N_2069);
and U3980 (N_3980,N_1907,N_2830);
or U3981 (N_3981,N_2248,N_1759);
nand U3982 (N_3982,N_1984,N_1826);
nand U3983 (N_3983,N_2049,N_2281);
xor U3984 (N_3984,N_2716,N_2637);
nor U3985 (N_3985,N_2651,N_2510);
and U3986 (N_3986,N_2483,N_1724);
and U3987 (N_3987,N_1892,N_1931);
xnor U3988 (N_3988,N_2835,N_1516);
nand U3989 (N_3989,N_1596,N_1823);
or U3990 (N_3990,N_1534,N_2296);
nor U3991 (N_3991,N_2906,N_2710);
nand U3992 (N_3992,N_2605,N_1931);
nand U3993 (N_3993,N_2486,N_2181);
nand U3994 (N_3994,N_1558,N_1838);
nor U3995 (N_3995,N_1630,N_2071);
nor U3996 (N_3996,N_1533,N_2845);
nor U3997 (N_3997,N_2415,N_1659);
nand U3998 (N_3998,N_2731,N_2927);
or U3999 (N_3999,N_1721,N_1791);
xor U4000 (N_4000,N_1958,N_2581);
or U4001 (N_4001,N_2968,N_2787);
nor U4002 (N_4002,N_2110,N_2557);
and U4003 (N_4003,N_1982,N_2365);
nor U4004 (N_4004,N_2694,N_1971);
xor U4005 (N_4005,N_2772,N_1994);
xor U4006 (N_4006,N_2392,N_2521);
nor U4007 (N_4007,N_2601,N_2844);
nor U4008 (N_4008,N_2636,N_2384);
or U4009 (N_4009,N_1813,N_1709);
or U4010 (N_4010,N_2455,N_2400);
and U4011 (N_4011,N_2151,N_1841);
nor U4012 (N_4012,N_2451,N_1691);
nand U4013 (N_4013,N_1532,N_2199);
nand U4014 (N_4014,N_2540,N_1671);
or U4015 (N_4015,N_1655,N_2209);
and U4016 (N_4016,N_1564,N_1782);
or U4017 (N_4017,N_2477,N_2077);
or U4018 (N_4018,N_1675,N_2329);
or U4019 (N_4019,N_2567,N_2688);
and U4020 (N_4020,N_2060,N_1636);
nor U4021 (N_4021,N_2068,N_1798);
or U4022 (N_4022,N_2158,N_1622);
nand U4023 (N_4023,N_2586,N_1992);
and U4024 (N_4024,N_1743,N_2602);
nand U4025 (N_4025,N_2860,N_2408);
and U4026 (N_4026,N_2247,N_2214);
and U4027 (N_4027,N_2624,N_2757);
nor U4028 (N_4028,N_2262,N_2192);
nand U4029 (N_4029,N_1664,N_1595);
or U4030 (N_4030,N_1861,N_1956);
or U4031 (N_4031,N_2598,N_1861);
and U4032 (N_4032,N_2922,N_2108);
nor U4033 (N_4033,N_2883,N_1517);
nand U4034 (N_4034,N_1994,N_1563);
nor U4035 (N_4035,N_2867,N_2334);
and U4036 (N_4036,N_2244,N_2309);
nand U4037 (N_4037,N_1613,N_1825);
nor U4038 (N_4038,N_2425,N_2011);
xor U4039 (N_4039,N_2057,N_2806);
or U4040 (N_4040,N_1875,N_2283);
and U4041 (N_4041,N_2742,N_2998);
and U4042 (N_4042,N_2759,N_1763);
nand U4043 (N_4043,N_2395,N_2203);
nand U4044 (N_4044,N_2590,N_2428);
nand U4045 (N_4045,N_1660,N_1554);
nor U4046 (N_4046,N_2669,N_2448);
xor U4047 (N_4047,N_1874,N_1519);
and U4048 (N_4048,N_2319,N_2180);
and U4049 (N_4049,N_2458,N_2733);
and U4050 (N_4050,N_2376,N_1964);
or U4051 (N_4051,N_2760,N_2277);
xor U4052 (N_4052,N_1652,N_1974);
or U4053 (N_4053,N_2287,N_1818);
nand U4054 (N_4054,N_1635,N_2644);
nand U4055 (N_4055,N_2140,N_2500);
and U4056 (N_4056,N_2136,N_2447);
and U4057 (N_4057,N_2822,N_2955);
or U4058 (N_4058,N_2138,N_2839);
nand U4059 (N_4059,N_2060,N_2115);
xnor U4060 (N_4060,N_2013,N_2274);
nand U4061 (N_4061,N_2369,N_2239);
or U4062 (N_4062,N_1877,N_2175);
nor U4063 (N_4063,N_1980,N_2609);
nand U4064 (N_4064,N_2276,N_2815);
or U4065 (N_4065,N_2974,N_1888);
nor U4066 (N_4066,N_1602,N_1728);
nor U4067 (N_4067,N_2004,N_2793);
nor U4068 (N_4068,N_2477,N_2276);
nor U4069 (N_4069,N_1610,N_2761);
nand U4070 (N_4070,N_1884,N_2905);
nand U4071 (N_4071,N_2740,N_2205);
nor U4072 (N_4072,N_2651,N_1711);
and U4073 (N_4073,N_2767,N_1622);
nand U4074 (N_4074,N_2710,N_1853);
nor U4075 (N_4075,N_2532,N_1821);
xor U4076 (N_4076,N_2718,N_2682);
xnor U4077 (N_4077,N_2206,N_2494);
or U4078 (N_4078,N_1997,N_1723);
xnor U4079 (N_4079,N_2843,N_2659);
xor U4080 (N_4080,N_1743,N_2762);
xor U4081 (N_4081,N_2445,N_2511);
nor U4082 (N_4082,N_2167,N_1641);
xnor U4083 (N_4083,N_1631,N_2002);
and U4084 (N_4084,N_1506,N_1756);
and U4085 (N_4085,N_1920,N_2534);
nor U4086 (N_4086,N_2592,N_2801);
nand U4087 (N_4087,N_2973,N_1949);
or U4088 (N_4088,N_2425,N_2362);
and U4089 (N_4089,N_2138,N_1814);
nand U4090 (N_4090,N_1859,N_2841);
nand U4091 (N_4091,N_1927,N_2393);
xor U4092 (N_4092,N_2829,N_2032);
nand U4093 (N_4093,N_2745,N_2497);
nand U4094 (N_4094,N_1556,N_1979);
and U4095 (N_4095,N_1544,N_2251);
or U4096 (N_4096,N_1598,N_1866);
and U4097 (N_4097,N_2024,N_2025);
or U4098 (N_4098,N_1745,N_2462);
nand U4099 (N_4099,N_2265,N_1725);
and U4100 (N_4100,N_1859,N_2895);
nor U4101 (N_4101,N_1743,N_2268);
nand U4102 (N_4102,N_1865,N_2754);
nor U4103 (N_4103,N_2322,N_1659);
xnor U4104 (N_4104,N_2211,N_2769);
or U4105 (N_4105,N_2339,N_2974);
nor U4106 (N_4106,N_2075,N_2036);
nor U4107 (N_4107,N_1626,N_2830);
nor U4108 (N_4108,N_2352,N_1812);
and U4109 (N_4109,N_2899,N_1786);
nor U4110 (N_4110,N_1663,N_1729);
and U4111 (N_4111,N_2279,N_2829);
or U4112 (N_4112,N_1897,N_2803);
and U4113 (N_4113,N_2378,N_2102);
nor U4114 (N_4114,N_2208,N_2664);
nor U4115 (N_4115,N_1849,N_1921);
nor U4116 (N_4116,N_1860,N_1967);
and U4117 (N_4117,N_2855,N_2428);
nand U4118 (N_4118,N_1999,N_1944);
or U4119 (N_4119,N_1927,N_2134);
nand U4120 (N_4120,N_2963,N_2088);
nor U4121 (N_4121,N_2105,N_1787);
xnor U4122 (N_4122,N_2044,N_2060);
or U4123 (N_4123,N_2752,N_1661);
or U4124 (N_4124,N_2023,N_2372);
nand U4125 (N_4125,N_2866,N_1560);
nand U4126 (N_4126,N_1787,N_2352);
nor U4127 (N_4127,N_2027,N_1866);
or U4128 (N_4128,N_1832,N_2151);
or U4129 (N_4129,N_1830,N_1509);
or U4130 (N_4130,N_2442,N_1532);
nor U4131 (N_4131,N_1933,N_2143);
nor U4132 (N_4132,N_1979,N_2972);
xor U4133 (N_4133,N_2335,N_1994);
nor U4134 (N_4134,N_2337,N_2675);
nand U4135 (N_4135,N_2525,N_2762);
xor U4136 (N_4136,N_1964,N_2757);
nor U4137 (N_4137,N_2667,N_1947);
or U4138 (N_4138,N_2058,N_1929);
and U4139 (N_4139,N_1529,N_1609);
and U4140 (N_4140,N_2934,N_2187);
or U4141 (N_4141,N_1850,N_1955);
nor U4142 (N_4142,N_2353,N_1743);
nor U4143 (N_4143,N_2353,N_2427);
nand U4144 (N_4144,N_2467,N_2037);
nor U4145 (N_4145,N_2981,N_1741);
nand U4146 (N_4146,N_2456,N_2139);
nor U4147 (N_4147,N_2091,N_2738);
and U4148 (N_4148,N_1976,N_1825);
or U4149 (N_4149,N_2092,N_1629);
nand U4150 (N_4150,N_2963,N_2160);
and U4151 (N_4151,N_2387,N_1679);
nand U4152 (N_4152,N_2813,N_2679);
or U4153 (N_4153,N_2608,N_2580);
nor U4154 (N_4154,N_2452,N_2671);
nor U4155 (N_4155,N_1871,N_1752);
xor U4156 (N_4156,N_1586,N_1526);
xor U4157 (N_4157,N_2686,N_2924);
or U4158 (N_4158,N_1973,N_2740);
or U4159 (N_4159,N_2791,N_2923);
or U4160 (N_4160,N_1898,N_1770);
nor U4161 (N_4161,N_1538,N_1758);
or U4162 (N_4162,N_1631,N_2856);
nand U4163 (N_4163,N_2157,N_2493);
nor U4164 (N_4164,N_2350,N_1916);
or U4165 (N_4165,N_2852,N_2938);
xnor U4166 (N_4166,N_1906,N_2082);
nor U4167 (N_4167,N_2758,N_2953);
xnor U4168 (N_4168,N_2293,N_2666);
or U4169 (N_4169,N_2522,N_2287);
nor U4170 (N_4170,N_1886,N_2042);
and U4171 (N_4171,N_2306,N_1539);
and U4172 (N_4172,N_2986,N_2177);
nand U4173 (N_4173,N_2816,N_2987);
nand U4174 (N_4174,N_2687,N_2602);
nor U4175 (N_4175,N_2668,N_2953);
nand U4176 (N_4176,N_1780,N_2488);
nor U4177 (N_4177,N_2143,N_2487);
xnor U4178 (N_4178,N_2122,N_2249);
and U4179 (N_4179,N_1565,N_1761);
nor U4180 (N_4180,N_2556,N_1737);
and U4181 (N_4181,N_2349,N_2190);
nand U4182 (N_4182,N_2036,N_1891);
nor U4183 (N_4183,N_2153,N_2764);
and U4184 (N_4184,N_2668,N_1789);
or U4185 (N_4185,N_2706,N_2414);
nand U4186 (N_4186,N_2356,N_2418);
nand U4187 (N_4187,N_1703,N_1796);
nor U4188 (N_4188,N_1779,N_2378);
or U4189 (N_4189,N_2401,N_2335);
xor U4190 (N_4190,N_2447,N_2690);
and U4191 (N_4191,N_1933,N_1844);
nand U4192 (N_4192,N_2830,N_2453);
and U4193 (N_4193,N_2618,N_1681);
and U4194 (N_4194,N_1566,N_2854);
or U4195 (N_4195,N_2882,N_2464);
nand U4196 (N_4196,N_1995,N_1655);
nand U4197 (N_4197,N_2656,N_1995);
xnor U4198 (N_4198,N_1595,N_1765);
nor U4199 (N_4199,N_1732,N_2677);
nand U4200 (N_4200,N_2923,N_1882);
or U4201 (N_4201,N_2102,N_2627);
or U4202 (N_4202,N_2154,N_2266);
and U4203 (N_4203,N_2262,N_1627);
nor U4204 (N_4204,N_1710,N_2963);
and U4205 (N_4205,N_2678,N_2289);
nor U4206 (N_4206,N_2838,N_1741);
or U4207 (N_4207,N_2104,N_1673);
xnor U4208 (N_4208,N_1764,N_1766);
nand U4209 (N_4209,N_1746,N_2491);
nor U4210 (N_4210,N_2945,N_2104);
and U4211 (N_4211,N_2971,N_1708);
and U4212 (N_4212,N_2966,N_2515);
or U4213 (N_4213,N_1650,N_2881);
or U4214 (N_4214,N_2592,N_2007);
nor U4215 (N_4215,N_2569,N_1508);
nand U4216 (N_4216,N_2804,N_1524);
nand U4217 (N_4217,N_1970,N_2701);
and U4218 (N_4218,N_1872,N_2249);
and U4219 (N_4219,N_2848,N_1780);
and U4220 (N_4220,N_2697,N_2961);
nand U4221 (N_4221,N_2779,N_2708);
nor U4222 (N_4222,N_2520,N_2794);
nand U4223 (N_4223,N_2012,N_1693);
nand U4224 (N_4224,N_2356,N_1619);
nor U4225 (N_4225,N_2528,N_1993);
xor U4226 (N_4226,N_2025,N_2443);
or U4227 (N_4227,N_2608,N_2437);
xnor U4228 (N_4228,N_2959,N_2791);
xnor U4229 (N_4229,N_1629,N_1791);
nand U4230 (N_4230,N_1719,N_2474);
and U4231 (N_4231,N_2109,N_2933);
nor U4232 (N_4232,N_2350,N_1910);
nand U4233 (N_4233,N_2415,N_2507);
nand U4234 (N_4234,N_1694,N_2915);
nor U4235 (N_4235,N_2256,N_2670);
and U4236 (N_4236,N_2917,N_2644);
and U4237 (N_4237,N_2614,N_2811);
nand U4238 (N_4238,N_2962,N_2218);
nor U4239 (N_4239,N_2546,N_2651);
or U4240 (N_4240,N_2892,N_1921);
or U4241 (N_4241,N_1970,N_1827);
or U4242 (N_4242,N_2950,N_2142);
and U4243 (N_4243,N_1646,N_1628);
nor U4244 (N_4244,N_2901,N_1505);
nor U4245 (N_4245,N_2146,N_2641);
and U4246 (N_4246,N_2589,N_2093);
nand U4247 (N_4247,N_2126,N_2687);
nor U4248 (N_4248,N_1854,N_2674);
and U4249 (N_4249,N_2965,N_1578);
nand U4250 (N_4250,N_2055,N_2057);
xor U4251 (N_4251,N_2625,N_2278);
and U4252 (N_4252,N_2329,N_1656);
nand U4253 (N_4253,N_2983,N_1672);
or U4254 (N_4254,N_1964,N_1737);
nand U4255 (N_4255,N_2974,N_2840);
nor U4256 (N_4256,N_2554,N_2178);
nor U4257 (N_4257,N_2949,N_2634);
nor U4258 (N_4258,N_1968,N_1656);
nor U4259 (N_4259,N_1628,N_2442);
and U4260 (N_4260,N_2701,N_2778);
or U4261 (N_4261,N_2491,N_2021);
xor U4262 (N_4262,N_2944,N_2749);
and U4263 (N_4263,N_1723,N_1591);
nand U4264 (N_4264,N_2506,N_2158);
or U4265 (N_4265,N_2738,N_2140);
nor U4266 (N_4266,N_2939,N_1605);
nor U4267 (N_4267,N_2827,N_1931);
nor U4268 (N_4268,N_2727,N_2268);
nand U4269 (N_4269,N_2730,N_1791);
or U4270 (N_4270,N_2694,N_1976);
and U4271 (N_4271,N_2779,N_2746);
xor U4272 (N_4272,N_1952,N_2795);
and U4273 (N_4273,N_2205,N_1657);
xnor U4274 (N_4274,N_2140,N_1580);
and U4275 (N_4275,N_2180,N_1762);
nor U4276 (N_4276,N_1908,N_2556);
nor U4277 (N_4277,N_1907,N_2260);
and U4278 (N_4278,N_2193,N_2827);
xnor U4279 (N_4279,N_2590,N_2831);
nor U4280 (N_4280,N_2172,N_2014);
xor U4281 (N_4281,N_2406,N_2949);
and U4282 (N_4282,N_2300,N_1975);
and U4283 (N_4283,N_1733,N_2889);
and U4284 (N_4284,N_2622,N_2410);
nor U4285 (N_4285,N_1758,N_1654);
nor U4286 (N_4286,N_1608,N_2104);
nand U4287 (N_4287,N_2146,N_2951);
or U4288 (N_4288,N_2153,N_1641);
xnor U4289 (N_4289,N_2892,N_2911);
nand U4290 (N_4290,N_1847,N_2249);
nand U4291 (N_4291,N_1852,N_2752);
or U4292 (N_4292,N_2378,N_1847);
nor U4293 (N_4293,N_2166,N_1797);
nor U4294 (N_4294,N_2375,N_1526);
nor U4295 (N_4295,N_2955,N_1994);
nor U4296 (N_4296,N_2006,N_1581);
or U4297 (N_4297,N_2936,N_2903);
and U4298 (N_4298,N_1583,N_2172);
and U4299 (N_4299,N_2093,N_1891);
nor U4300 (N_4300,N_1582,N_2639);
or U4301 (N_4301,N_1635,N_2228);
or U4302 (N_4302,N_2495,N_2568);
xor U4303 (N_4303,N_2664,N_2074);
nor U4304 (N_4304,N_2119,N_1657);
nor U4305 (N_4305,N_2427,N_1584);
and U4306 (N_4306,N_2926,N_2121);
nand U4307 (N_4307,N_1968,N_2276);
nand U4308 (N_4308,N_2257,N_2019);
nor U4309 (N_4309,N_2824,N_1643);
or U4310 (N_4310,N_1791,N_2617);
xnor U4311 (N_4311,N_1874,N_1673);
nand U4312 (N_4312,N_1542,N_1678);
nand U4313 (N_4313,N_2580,N_2059);
and U4314 (N_4314,N_1608,N_2935);
xnor U4315 (N_4315,N_1704,N_1619);
or U4316 (N_4316,N_1541,N_2195);
and U4317 (N_4317,N_2140,N_2497);
or U4318 (N_4318,N_2824,N_2591);
nand U4319 (N_4319,N_2794,N_2239);
or U4320 (N_4320,N_2808,N_2761);
and U4321 (N_4321,N_1512,N_1919);
nor U4322 (N_4322,N_2193,N_1667);
xor U4323 (N_4323,N_2101,N_1770);
or U4324 (N_4324,N_2118,N_2340);
nor U4325 (N_4325,N_2505,N_1534);
and U4326 (N_4326,N_2493,N_2002);
xnor U4327 (N_4327,N_2045,N_2338);
or U4328 (N_4328,N_2895,N_2070);
or U4329 (N_4329,N_2700,N_2480);
xnor U4330 (N_4330,N_1891,N_2787);
and U4331 (N_4331,N_2754,N_2713);
nand U4332 (N_4332,N_1944,N_2592);
and U4333 (N_4333,N_2534,N_1551);
nor U4334 (N_4334,N_1729,N_2252);
or U4335 (N_4335,N_2410,N_1887);
nand U4336 (N_4336,N_2965,N_1508);
nor U4337 (N_4337,N_2674,N_1546);
nand U4338 (N_4338,N_1520,N_1828);
nand U4339 (N_4339,N_1516,N_2555);
nor U4340 (N_4340,N_2458,N_2198);
nor U4341 (N_4341,N_2516,N_2128);
nand U4342 (N_4342,N_2224,N_2827);
xor U4343 (N_4343,N_2039,N_1653);
or U4344 (N_4344,N_2012,N_2181);
and U4345 (N_4345,N_2591,N_1763);
nor U4346 (N_4346,N_2016,N_1917);
nand U4347 (N_4347,N_2454,N_2832);
or U4348 (N_4348,N_2851,N_1669);
or U4349 (N_4349,N_2727,N_1733);
or U4350 (N_4350,N_2351,N_2579);
and U4351 (N_4351,N_2846,N_1817);
and U4352 (N_4352,N_1692,N_2746);
nand U4353 (N_4353,N_2091,N_1952);
nor U4354 (N_4354,N_2170,N_1576);
nand U4355 (N_4355,N_2890,N_1952);
xnor U4356 (N_4356,N_2732,N_2609);
xor U4357 (N_4357,N_1972,N_2855);
or U4358 (N_4358,N_2464,N_2229);
nor U4359 (N_4359,N_2479,N_1632);
nand U4360 (N_4360,N_1983,N_2966);
and U4361 (N_4361,N_1911,N_2402);
nor U4362 (N_4362,N_2500,N_2997);
and U4363 (N_4363,N_2871,N_2665);
or U4364 (N_4364,N_2206,N_2337);
or U4365 (N_4365,N_1671,N_2154);
nor U4366 (N_4366,N_2099,N_1901);
or U4367 (N_4367,N_2414,N_2441);
and U4368 (N_4368,N_2802,N_1733);
or U4369 (N_4369,N_2108,N_2162);
nor U4370 (N_4370,N_1507,N_1633);
and U4371 (N_4371,N_2192,N_2630);
nand U4372 (N_4372,N_2796,N_2253);
nor U4373 (N_4373,N_2655,N_2259);
nor U4374 (N_4374,N_2988,N_2714);
nand U4375 (N_4375,N_2285,N_1555);
nand U4376 (N_4376,N_2323,N_2737);
and U4377 (N_4377,N_2261,N_1731);
nand U4378 (N_4378,N_2317,N_2833);
and U4379 (N_4379,N_2842,N_2835);
or U4380 (N_4380,N_1755,N_2374);
and U4381 (N_4381,N_2039,N_2893);
nand U4382 (N_4382,N_1979,N_1874);
or U4383 (N_4383,N_1704,N_2802);
and U4384 (N_4384,N_1985,N_1516);
nand U4385 (N_4385,N_2785,N_2900);
and U4386 (N_4386,N_1969,N_2996);
and U4387 (N_4387,N_1823,N_2107);
xor U4388 (N_4388,N_2508,N_2931);
and U4389 (N_4389,N_2342,N_1642);
xnor U4390 (N_4390,N_1926,N_2637);
nand U4391 (N_4391,N_2365,N_1508);
nand U4392 (N_4392,N_1514,N_2351);
and U4393 (N_4393,N_2077,N_1674);
and U4394 (N_4394,N_1574,N_1824);
nand U4395 (N_4395,N_2210,N_2757);
or U4396 (N_4396,N_2060,N_2067);
or U4397 (N_4397,N_2435,N_2685);
or U4398 (N_4398,N_1804,N_1948);
or U4399 (N_4399,N_2205,N_2395);
or U4400 (N_4400,N_1969,N_1585);
xnor U4401 (N_4401,N_2144,N_2484);
nor U4402 (N_4402,N_2106,N_2952);
nand U4403 (N_4403,N_1648,N_2954);
and U4404 (N_4404,N_1872,N_2171);
or U4405 (N_4405,N_2459,N_2785);
nand U4406 (N_4406,N_1540,N_2549);
nor U4407 (N_4407,N_2678,N_2770);
nand U4408 (N_4408,N_1828,N_1628);
and U4409 (N_4409,N_2602,N_2508);
nand U4410 (N_4410,N_1543,N_2362);
or U4411 (N_4411,N_1871,N_2108);
or U4412 (N_4412,N_2803,N_2129);
xor U4413 (N_4413,N_2712,N_1536);
and U4414 (N_4414,N_1683,N_2365);
nand U4415 (N_4415,N_2605,N_2875);
and U4416 (N_4416,N_1798,N_2680);
or U4417 (N_4417,N_2264,N_1622);
nand U4418 (N_4418,N_2977,N_2404);
nor U4419 (N_4419,N_2006,N_1843);
nand U4420 (N_4420,N_1940,N_2698);
nand U4421 (N_4421,N_2634,N_1588);
nor U4422 (N_4422,N_2767,N_2152);
and U4423 (N_4423,N_1848,N_2801);
or U4424 (N_4424,N_1755,N_1748);
nand U4425 (N_4425,N_2782,N_2037);
nand U4426 (N_4426,N_2798,N_1834);
or U4427 (N_4427,N_2831,N_2756);
and U4428 (N_4428,N_2476,N_2535);
xor U4429 (N_4429,N_2440,N_2843);
xor U4430 (N_4430,N_2990,N_2922);
and U4431 (N_4431,N_2743,N_2415);
nor U4432 (N_4432,N_1814,N_1811);
or U4433 (N_4433,N_2556,N_2466);
nor U4434 (N_4434,N_1837,N_1774);
nand U4435 (N_4435,N_1970,N_2548);
nand U4436 (N_4436,N_2140,N_2194);
or U4437 (N_4437,N_2237,N_1605);
nor U4438 (N_4438,N_2777,N_1565);
xnor U4439 (N_4439,N_1714,N_2269);
nor U4440 (N_4440,N_2416,N_2571);
and U4441 (N_4441,N_2013,N_1738);
nand U4442 (N_4442,N_1862,N_1972);
or U4443 (N_4443,N_2344,N_2097);
nor U4444 (N_4444,N_2534,N_2649);
nand U4445 (N_4445,N_1577,N_2198);
nand U4446 (N_4446,N_1569,N_2986);
xor U4447 (N_4447,N_2893,N_2331);
or U4448 (N_4448,N_2459,N_1803);
xor U4449 (N_4449,N_1992,N_1833);
nor U4450 (N_4450,N_2933,N_1780);
and U4451 (N_4451,N_2480,N_1946);
xnor U4452 (N_4452,N_2112,N_2979);
nor U4453 (N_4453,N_2531,N_2332);
and U4454 (N_4454,N_2789,N_2306);
and U4455 (N_4455,N_2686,N_1618);
nor U4456 (N_4456,N_2728,N_1623);
or U4457 (N_4457,N_1756,N_1524);
and U4458 (N_4458,N_2169,N_2350);
nand U4459 (N_4459,N_2030,N_2193);
or U4460 (N_4460,N_1516,N_2625);
nand U4461 (N_4461,N_2096,N_2916);
and U4462 (N_4462,N_2505,N_2619);
nor U4463 (N_4463,N_2700,N_1747);
xor U4464 (N_4464,N_1950,N_1710);
and U4465 (N_4465,N_2852,N_2549);
nand U4466 (N_4466,N_2889,N_1921);
nand U4467 (N_4467,N_2141,N_2280);
nor U4468 (N_4468,N_2020,N_2835);
nand U4469 (N_4469,N_2244,N_2934);
and U4470 (N_4470,N_2326,N_2718);
or U4471 (N_4471,N_2844,N_2044);
nor U4472 (N_4472,N_2330,N_1695);
nor U4473 (N_4473,N_2985,N_2689);
nor U4474 (N_4474,N_2587,N_2515);
or U4475 (N_4475,N_2217,N_1988);
xor U4476 (N_4476,N_2211,N_2278);
xnor U4477 (N_4477,N_2447,N_2967);
or U4478 (N_4478,N_2210,N_1508);
or U4479 (N_4479,N_2280,N_2966);
nand U4480 (N_4480,N_2350,N_2134);
nor U4481 (N_4481,N_2483,N_2649);
xnor U4482 (N_4482,N_2672,N_2759);
or U4483 (N_4483,N_2773,N_2635);
and U4484 (N_4484,N_2914,N_1674);
nand U4485 (N_4485,N_2827,N_2644);
or U4486 (N_4486,N_2633,N_1905);
nand U4487 (N_4487,N_1975,N_1848);
nor U4488 (N_4488,N_2496,N_1558);
and U4489 (N_4489,N_1554,N_2555);
nand U4490 (N_4490,N_2803,N_2598);
nor U4491 (N_4491,N_2026,N_1681);
and U4492 (N_4492,N_2115,N_2795);
or U4493 (N_4493,N_1566,N_2128);
and U4494 (N_4494,N_1502,N_2170);
or U4495 (N_4495,N_2882,N_2784);
or U4496 (N_4496,N_1582,N_2421);
or U4497 (N_4497,N_2829,N_2709);
nand U4498 (N_4498,N_2373,N_1972);
and U4499 (N_4499,N_2610,N_2190);
nor U4500 (N_4500,N_3877,N_3725);
nand U4501 (N_4501,N_4241,N_3665);
and U4502 (N_4502,N_3497,N_3970);
or U4503 (N_4503,N_3105,N_3135);
nand U4504 (N_4504,N_3142,N_3998);
nor U4505 (N_4505,N_3741,N_4437);
and U4506 (N_4506,N_3512,N_3723);
nor U4507 (N_4507,N_3358,N_3492);
or U4508 (N_4508,N_3412,N_3250);
nor U4509 (N_4509,N_3165,N_4433);
or U4510 (N_4510,N_4285,N_4348);
xor U4511 (N_4511,N_3567,N_3447);
nand U4512 (N_4512,N_3040,N_4386);
or U4513 (N_4513,N_3559,N_3697);
or U4514 (N_4514,N_4216,N_3526);
and U4515 (N_4515,N_3022,N_3989);
and U4516 (N_4516,N_3574,N_4017);
nand U4517 (N_4517,N_3798,N_3228);
nor U4518 (N_4518,N_4217,N_3516);
nand U4519 (N_4519,N_4377,N_3538);
and U4520 (N_4520,N_4031,N_3416);
nand U4521 (N_4521,N_3427,N_3924);
nand U4522 (N_4522,N_4033,N_3084);
nor U4523 (N_4523,N_3552,N_4035);
or U4524 (N_4524,N_4109,N_3299);
nor U4525 (N_4525,N_3896,N_4292);
or U4526 (N_4526,N_3783,N_3733);
or U4527 (N_4527,N_3764,N_3077);
and U4528 (N_4528,N_3611,N_3980);
xnor U4529 (N_4529,N_3223,N_3923);
nand U4530 (N_4530,N_3939,N_3781);
and U4531 (N_4531,N_3953,N_3279);
nor U4532 (N_4532,N_3351,N_4221);
nor U4533 (N_4533,N_3820,N_4062);
and U4534 (N_4534,N_3500,N_3450);
nand U4535 (N_4535,N_3442,N_3964);
nand U4536 (N_4536,N_3999,N_3187);
or U4537 (N_4537,N_3286,N_3336);
nor U4538 (N_4538,N_3128,N_3839);
nor U4539 (N_4539,N_3395,N_3817);
or U4540 (N_4540,N_3340,N_3487);
or U4541 (N_4541,N_3703,N_3828);
nand U4542 (N_4542,N_3504,N_3963);
xor U4543 (N_4543,N_3701,N_3151);
nor U4544 (N_4544,N_3090,N_4481);
nand U4545 (N_4545,N_3911,N_3280);
nand U4546 (N_4546,N_4007,N_3672);
or U4547 (N_4547,N_4191,N_3052);
nand U4548 (N_4548,N_3739,N_4462);
nand U4549 (N_4549,N_3962,N_3950);
and U4550 (N_4550,N_3735,N_4232);
or U4551 (N_4551,N_4209,N_3523);
nand U4552 (N_4552,N_4101,N_3276);
nand U4553 (N_4553,N_3385,N_3848);
xor U4554 (N_4554,N_3401,N_3372);
nor U4555 (N_4555,N_3083,N_4372);
nand U4556 (N_4556,N_4336,N_4270);
nand U4557 (N_4557,N_3232,N_4340);
or U4558 (N_4558,N_4063,N_3146);
nor U4559 (N_4559,N_3321,N_3251);
or U4560 (N_4560,N_3932,N_3186);
and U4561 (N_4561,N_3485,N_3916);
nor U4562 (N_4562,N_3136,N_4163);
nand U4563 (N_4563,N_4029,N_3503);
and U4564 (N_4564,N_4065,N_3490);
xnor U4565 (N_4565,N_3753,N_4376);
and U4566 (N_4566,N_3515,N_3059);
or U4567 (N_4567,N_4180,N_4395);
nor U4568 (N_4568,N_3803,N_3646);
and U4569 (N_4569,N_3566,N_3638);
nor U4570 (N_4570,N_4161,N_3884);
nand U4571 (N_4571,N_3293,N_3027);
nor U4572 (N_4572,N_3092,N_3683);
nor U4573 (N_4573,N_3102,N_3029);
nand U4574 (N_4574,N_4457,N_3061);
and U4575 (N_4575,N_4173,N_3007);
and U4576 (N_4576,N_4020,N_3235);
nor U4577 (N_4577,N_3690,N_3806);
nor U4578 (N_4578,N_3586,N_3630);
nand U4579 (N_4579,N_3288,N_3231);
nor U4580 (N_4580,N_3938,N_3431);
nor U4581 (N_4581,N_3020,N_4042);
nor U4582 (N_4582,N_3705,N_4260);
nor U4583 (N_4583,N_3317,N_4126);
nand U4584 (N_4584,N_3238,N_4305);
nand U4585 (N_4585,N_3951,N_3847);
or U4586 (N_4586,N_3054,N_4047);
nand U4587 (N_4587,N_3969,N_3650);
or U4588 (N_4588,N_3555,N_3324);
nand U4589 (N_4589,N_4154,N_3031);
nor U4590 (N_4590,N_4067,N_3551);
or U4591 (N_4591,N_4186,N_3343);
nor U4592 (N_4592,N_4210,N_3775);
nand U4593 (N_4593,N_3906,N_3687);
xnor U4594 (N_4594,N_3987,N_3444);
or U4595 (N_4595,N_3995,N_4150);
nor U4596 (N_4596,N_3443,N_3382);
and U4597 (N_4597,N_3898,N_4284);
or U4598 (N_4598,N_3274,N_3118);
nor U4599 (N_4599,N_4080,N_3393);
nor U4600 (N_4600,N_4034,N_3320);
and U4601 (N_4601,N_3166,N_3901);
or U4602 (N_4602,N_3270,N_4324);
xnor U4603 (N_4603,N_4152,N_4118);
nor U4604 (N_4604,N_3239,N_3009);
xnor U4605 (N_4605,N_3263,N_3153);
nor U4606 (N_4606,N_3921,N_3300);
nand U4607 (N_4607,N_3058,N_3063);
xor U4608 (N_4608,N_3873,N_3233);
nor U4609 (N_4609,N_3508,N_4106);
nand U4610 (N_4610,N_3008,N_3653);
nor U4611 (N_4611,N_4235,N_3615);
and U4612 (N_4612,N_4002,N_4061);
and U4613 (N_4613,N_3282,N_4429);
and U4614 (N_4614,N_3434,N_3837);
nor U4615 (N_4615,N_3868,N_3674);
or U4616 (N_4616,N_3547,N_3047);
nor U4617 (N_4617,N_4351,N_3180);
or U4618 (N_4618,N_3907,N_3678);
and U4619 (N_4619,N_4281,N_3339);
nor U4620 (N_4620,N_3377,N_3821);
xnor U4621 (N_4621,N_3120,N_3517);
and U4622 (N_4622,N_3928,N_4265);
or U4623 (N_4623,N_3660,N_3578);
or U4624 (N_4624,N_3730,N_3316);
nand U4625 (N_4625,N_3082,N_3438);
nand U4626 (N_4626,N_4022,N_3230);
and U4627 (N_4627,N_4129,N_3307);
or U4628 (N_4628,N_3600,N_4276);
and U4629 (N_4629,N_3761,N_3494);
and U4630 (N_4630,N_4011,N_3297);
xor U4631 (N_4631,N_3954,N_4293);
nand U4632 (N_4632,N_4024,N_4330);
and U4633 (N_4633,N_4289,N_3154);
nand U4634 (N_4634,N_3131,N_3161);
nand U4635 (N_4635,N_4113,N_3979);
or U4636 (N_4636,N_3298,N_3356);
and U4637 (N_4637,N_4309,N_3724);
or U4638 (N_4638,N_3430,N_3426);
nor U4639 (N_4639,N_3091,N_3460);
nor U4640 (N_4640,N_3941,N_3693);
nand U4641 (N_4641,N_3897,N_3489);
nand U4642 (N_4642,N_3342,N_3220);
or U4643 (N_4643,N_3456,N_4468);
nand U4644 (N_4644,N_4399,N_4127);
nor U4645 (N_4645,N_3062,N_3642);
nor U4646 (N_4646,N_3287,N_4038);
nor U4647 (N_4647,N_4425,N_4411);
or U4648 (N_4648,N_3234,N_4082);
nor U4649 (N_4649,N_4428,N_4475);
nor U4650 (N_4650,N_4103,N_3134);
nor U4651 (N_4651,N_4280,N_4383);
nand U4652 (N_4652,N_4205,N_3719);
xnor U4653 (N_4653,N_3432,N_4440);
and U4654 (N_4654,N_3915,N_3992);
nand U4655 (N_4655,N_3772,N_4257);
nand U4656 (N_4656,N_3689,N_3913);
or U4657 (N_4657,N_4350,N_3874);
nand U4658 (N_4658,N_3405,N_4146);
xnor U4659 (N_4659,N_3588,N_4486);
nor U4660 (N_4660,N_3985,N_3418);
and U4661 (N_4661,N_3943,N_3776);
and U4662 (N_4662,N_3005,N_4489);
nand U4663 (N_4663,N_3086,N_3127);
xnor U4664 (N_4664,N_4215,N_4242);
and U4665 (N_4665,N_3347,N_4357);
nand U4666 (N_4666,N_3577,N_4325);
nor U4667 (N_4667,N_3527,N_3840);
xor U4668 (N_4668,N_4201,N_4159);
and U4669 (N_4669,N_3625,N_3173);
or U4670 (N_4670,N_3277,N_3056);
nand U4671 (N_4671,N_3016,N_3591);
nor U4672 (N_4672,N_4111,N_3870);
or U4673 (N_4673,N_3064,N_4054);
and U4674 (N_4674,N_3666,N_3309);
nor U4675 (N_4675,N_4479,N_3685);
or U4676 (N_4676,N_3659,N_3836);
and U4677 (N_4677,N_4250,N_3830);
and U4678 (N_4678,N_4439,N_4172);
xor U4679 (N_4679,N_3268,N_4246);
nor U4680 (N_4680,N_3914,N_3209);
xor U4681 (N_4681,N_3773,N_3010);
and U4682 (N_4682,N_3875,N_3306);
nor U4683 (N_4683,N_3422,N_3344);
nor U4684 (N_4684,N_3483,N_3604);
nor U4685 (N_4685,N_4368,N_3856);
nand U4686 (N_4686,N_3721,N_3408);
and U4687 (N_4687,N_3057,N_3449);
and U4688 (N_4688,N_4361,N_3179);
or U4689 (N_4689,N_3150,N_3766);
nand U4690 (N_4690,N_3986,N_4308);
and U4691 (N_4691,N_3070,N_3688);
nand U4692 (N_4692,N_4473,N_4435);
nor U4693 (N_4693,N_4236,N_4389);
and U4694 (N_4694,N_4119,N_4043);
nor U4695 (N_4695,N_3885,N_3505);
nand U4696 (N_4696,N_3144,N_3758);
nor U4697 (N_4697,N_3114,N_3194);
and U4698 (N_4698,N_3853,N_4066);
nand U4699 (N_4699,N_4313,N_3881);
and U4700 (N_4700,N_3493,N_3810);
nor U4701 (N_4701,N_4014,N_3423);
or U4702 (N_4702,N_3147,N_4140);
or U4703 (N_4703,N_4358,N_4298);
xor U4704 (N_4704,N_3132,N_3794);
nand U4705 (N_4705,N_3681,N_3258);
or U4706 (N_4706,N_4245,N_3190);
or U4707 (N_4707,N_3355,N_3854);
nand U4708 (N_4708,N_3167,N_3381);
or U4709 (N_4709,N_3119,N_4401);
and U4710 (N_4710,N_3218,N_4070);
nor U4711 (N_4711,N_3759,N_4114);
nand U4712 (N_4712,N_3049,N_4446);
nand U4713 (N_4713,N_3155,N_3272);
or U4714 (N_4714,N_3708,N_3479);
and U4715 (N_4715,N_3349,N_3918);
nor U4716 (N_4716,N_3371,N_3583);
and U4717 (N_4717,N_3731,N_3971);
and U4718 (N_4718,N_3636,N_4177);
xor U4719 (N_4719,N_4064,N_3651);
nand U4720 (N_4720,N_3922,N_3389);
or U4721 (N_4721,N_3905,N_4384);
and U4722 (N_4722,N_4072,N_3858);
xnor U4723 (N_4723,N_4342,N_3774);
nor U4724 (N_4724,N_4090,N_4073);
and U4725 (N_4725,N_3936,N_4477);
nand U4726 (N_4726,N_4162,N_3544);
nor U4727 (N_4727,N_3826,N_3476);
or U4728 (N_4728,N_3023,N_3619);
xor U4729 (N_4729,N_3663,N_3601);
xor U4730 (N_4730,N_3707,N_3871);
nand U4731 (N_4731,N_3370,N_4431);
nand U4732 (N_4732,N_3825,N_4105);
nor U4733 (N_4733,N_4028,N_3894);
xor U4734 (N_4734,N_3213,N_3097);
nor U4735 (N_4735,N_3303,N_4121);
and U4736 (N_4736,N_4458,N_4332);
nand U4737 (N_4737,N_3872,N_3641);
and U4738 (N_4738,N_3704,N_4053);
nand U4739 (N_4739,N_4412,N_3260);
nor U4740 (N_4740,N_4418,N_3139);
and U4741 (N_4741,N_3602,N_3219);
or U4742 (N_4742,N_4199,N_4497);
nand U4743 (N_4743,N_3815,N_3661);
and U4744 (N_4744,N_3664,N_3934);
nand U4745 (N_4745,N_3787,N_3368);
nor U4746 (N_4746,N_3445,N_3181);
or U4747 (N_4747,N_3278,N_4030);
nand U4748 (N_4748,N_4198,N_3603);
nand U4749 (N_4749,N_4192,N_4083);
or U4750 (N_4750,N_3495,N_3419);
xnor U4751 (N_4751,N_4123,N_4353);
and U4752 (N_4752,N_4006,N_3961);
and U4753 (N_4753,N_3107,N_3554);
or U4754 (N_4754,N_4465,N_3327);
nand U4755 (N_4755,N_4422,N_4436);
nand U4756 (N_4756,N_4003,N_4086);
and U4757 (N_4757,N_4365,N_3657);
or U4758 (N_4758,N_4300,N_3745);
or U4759 (N_4759,N_3050,N_4442);
and U4760 (N_4760,N_3085,N_3305);
nand U4761 (N_4761,N_4144,N_3096);
and U4762 (N_4762,N_3388,N_4315);
xor U4763 (N_4763,N_3246,N_3126);
or U4764 (N_4764,N_3365,N_3518);
nand U4765 (N_4765,N_3413,N_3514);
nand U4766 (N_4766,N_3562,N_3015);
xor U4767 (N_4767,N_4012,N_4491);
or U4768 (N_4768,N_3789,N_3751);
or U4769 (N_4769,N_3121,N_3930);
or U4770 (N_4770,N_3784,N_3750);
and U4771 (N_4771,N_3677,N_3754);
nand U4772 (N_4772,N_3882,N_4183);
or U4773 (N_4773,N_3100,N_3507);
xor U4774 (N_4774,N_3537,N_3545);
nand U4775 (N_4775,N_3396,N_4312);
nand U4776 (N_4776,N_3631,N_3076);
and U4777 (N_4777,N_3786,N_4098);
nand U4778 (N_4778,N_3205,N_3192);
and U4779 (N_4779,N_3557,N_4166);
or U4780 (N_4780,N_3628,N_3752);
and U4781 (N_4781,N_3065,N_4455);
or U4782 (N_4782,N_4295,N_4249);
and U4783 (N_4783,N_3698,N_3536);
and U4784 (N_4784,N_3458,N_3225);
or U4785 (N_4785,N_3940,N_3041);
xnor U4786 (N_4786,N_3446,N_3594);
or U4787 (N_4787,N_4356,N_4147);
and U4788 (N_4788,N_3499,N_4075);
nand U4789 (N_4789,N_3302,N_4165);
nor U4790 (N_4790,N_3346,N_3204);
or U4791 (N_4791,N_4269,N_3221);
and U4792 (N_4792,N_3908,N_3269);
xnor U4793 (N_4793,N_4032,N_3193);
nand U4794 (N_4794,N_3384,N_3807);
or U4795 (N_4795,N_3414,N_4445);
nand U4796 (N_4796,N_3296,N_4419);
nand U4797 (N_4797,N_3101,N_3795);
or U4798 (N_4798,N_3402,N_4362);
and U4799 (N_4799,N_3360,N_4008);
nor U4800 (N_4800,N_4096,N_3867);
and U4801 (N_4801,N_3257,N_3273);
nand U4802 (N_4802,N_3823,N_4282);
nor U4803 (N_4803,N_3177,N_4149);
nor U4804 (N_4804,N_3624,N_3087);
and U4805 (N_4805,N_3767,N_3822);
or U4806 (N_4806,N_3138,N_3778);
and U4807 (N_4807,N_4088,N_3094);
or U4808 (N_4808,N_4181,N_3634);
nand U4809 (N_4809,N_3977,N_3684);
and U4810 (N_4810,N_3560,N_3457);
nand U4811 (N_4811,N_3799,N_3379);
and U4812 (N_4812,N_3202,N_4447);
nor U4813 (N_4813,N_3715,N_4333);
nand U4814 (N_4814,N_3982,N_3312);
or U4815 (N_4815,N_3919,N_3433);
nand U4816 (N_4816,N_4402,N_4262);
and U4817 (N_4817,N_3838,N_3929);
and U4818 (N_4818,N_4396,N_3044);
nand U4819 (N_4819,N_4370,N_3331);
nor U4820 (N_4820,N_3319,N_4174);
and U4821 (N_4821,N_3033,N_4005);
and U4822 (N_4822,N_3670,N_3909);
nor U4823 (N_4823,N_3859,N_4297);
or U4824 (N_4824,N_3359,N_3981);
and U4825 (N_4825,N_3744,N_3627);
nand U4826 (N_4826,N_3073,N_3944);
and U4827 (N_4827,N_4296,N_3648);
or U4828 (N_4828,N_4077,N_3960);
xor U4829 (N_4829,N_4335,N_3264);
nand U4830 (N_4830,N_3742,N_4321);
xor U4831 (N_4831,N_4423,N_3472);
or U4832 (N_4832,N_3722,N_3649);
nand U4833 (N_4833,N_4499,N_4448);
nand U4834 (N_4834,N_4317,N_4404);
nor U4835 (N_4835,N_3013,N_3647);
nand U4836 (N_4836,N_4466,N_4229);
xor U4837 (N_4837,N_4452,N_3927);
nor U4838 (N_4838,N_3511,N_4339);
or U4839 (N_4839,N_3607,N_3169);
or U4840 (N_4840,N_3183,N_3081);
nor U4841 (N_4841,N_4001,N_4320);
and U4842 (N_4842,N_4287,N_3680);
or U4843 (N_4843,N_3548,N_3301);
or U4844 (N_4844,N_3691,N_3437);
or U4845 (N_4845,N_3069,N_4311);
nor U4846 (N_4846,N_3935,N_4449);
nor U4847 (N_4847,N_3018,N_4274);
and U4848 (N_4848,N_4048,N_3322);
nand U4849 (N_4849,N_3095,N_4102);
nand U4850 (N_4850,N_3407,N_3606);
nor U4851 (N_4851,N_3878,N_3428);
or U4852 (N_4852,N_3522,N_3640);
or U4853 (N_4853,N_4375,N_4454);
nand U4854 (N_4854,N_3417,N_3525);
nor U4855 (N_4855,N_4403,N_4444);
nand U4856 (N_4856,N_3055,N_3243);
nor U4857 (N_4857,N_3410,N_3596);
xnor U4858 (N_4858,N_4156,N_3348);
and U4859 (N_4859,N_3869,N_4139);
xor U4860 (N_4860,N_3189,N_4044);
or U4861 (N_4861,N_3866,N_3644);
or U4862 (N_4862,N_3006,N_4329);
nand U4863 (N_4863,N_3903,N_4107);
or U4864 (N_4864,N_4112,N_3968);
or U4865 (N_4865,N_3686,N_4220);
and U4866 (N_4866,N_3785,N_3597);
nor U4867 (N_4867,N_4286,N_4299);
xor U4868 (N_4868,N_4234,N_3335);
nor U4869 (N_4869,N_3409,N_4239);
or U4870 (N_4870,N_4304,N_3176);
nor U4871 (N_4871,N_3592,N_3156);
nor U4872 (N_4872,N_3149,N_4359);
xor U4873 (N_4873,N_4104,N_4438);
or U4874 (N_4874,N_3354,N_3639);
xor U4875 (N_4875,N_4087,N_4469);
nand U4876 (N_4876,N_3550,N_4223);
and U4877 (N_4877,N_3206,N_4273);
and U4878 (N_4878,N_4266,N_3652);
nand U4879 (N_4879,N_4204,N_4097);
or U4880 (N_4880,N_4197,N_3088);
and U4881 (N_4881,N_4218,N_4405);
xor U4882 (N_4882,N_4347,N_3802);
nor U4883 (N_4883,N_4427,N_3956);
nor U4884 (N_4884,N_4247,N_3112);
and U4885 (N_4885,N_3845,N_3482);
or U4886 (N_4886,N_3108,N_4164);
nand U4887 (N_4887,N_3030,N_3695);
and U4888 (N_4888,N_4158,N_4195);
nor U4889 (N_4889,N_3865,N_3829);
xnor U4890 (N_4890,N_4476,N_4202);
nor U4891 (N_4891,N_4142,N_4049);
nor U4892 (N_4892,N_3561,N_3310);
and U4893 (N_4893,N_3337,N_4040);
xnor U4894 (N_4894,N_3814,N_4301);
and U4895 (N_4895,N_3966,N_4327);
or U4896 (N_4896,N_3496,N_4196);
or U4897 (N_4897,N_3612,N_4243);
and U4898 (N_4898,N_3621,N_3974);
nand U4899 (N_4899,N_4443,N_4125);
nor U4900 (N_4900,N_3290,N_3478);
nand U4901 (N_4901,N_3195,N_4175);
or U4902 (N_4902,N_3109,N_4135);
and U4903 (N_4903,N_3208,N_3833);
nor U4904 (N_4904,N_3256,N_3171);
and U4905 (N_4905,N_4290,N_4254);
or U4906 (N_4906,N_4398,N_3311);
and U4907 (N_4907,N_3972,N_3984);
nand U4908 (N_4908,N_3148,N_4294);
nor U4909 (N_4909,N_3104,N_4382);
or U4910 (N_4910,N_3726,N_3771);
nor U4911 (N_4911,N_3051,N_4379);
xor U4912 (N_4912,N_4354,N_3308);
nand U4913 (N_4913,N_3967,N_4413);
nor U4914 (N_4914,N_3217,N_3610);
nand U4915 (N_4915,N_4264,N_3860);
nor U4916 (N_4916,N_3667,N_3952);
and U4917 (N_4917,N_3528,N_3747);
or U4918 (N_4918,N_3618,N_4390);
nor U4919 (N_4919,N_3990,N_4226);
nand U4920 (N_4920,N_3598,N_4136);
nor U4921 (N_4921,N_4148,N_4143);
nor U4922 (N_4922,N_3480,N_4345);
xor U4923 (N_4923,N_3808,N_4071);
or U4924 (N_4924,N_4338,N_4076);
nand U4925 (N_4925,N_3117,N_3613);
and U4926 (N_4926,N_3740,N_3780);
or U4927 (N_4927,N_3014,N_4021);
nor U4928 (N_4928,N_3262,N_3352);
or U4929 (N_4929,N_4453,N_3463);
nor U4930 (N_4930,N_3702,N_3593);
nor U4931 (N_4931,N_3790,N_3888);
nand U4932 (N_4932,N_3762,N_4424);
or U4933 (N_4933,N_3454,N_3556);
or U4934 (N_4934,N_3345,N_3743);
nor U4935 (N_4935,N_3484,N_3247);
nand U4936 (N_4936,N_3633,N_3032);
and U4937 (N_4937,N_4492,N_4349);
and U4938 (N_4938,N_3068,N_4170);
nor U4939 (N_4939,N_3330,N_3415);
and U4940 (N_4940,N_3425,N_3214);
and U4941 (N_4941,N_4208,N_4261);
or U4942 (N_4942,N_3696,N_3453);
and U4943 (N_4943,N_3849,N_3043);
or U4944 (N_4944,N_3501,N_3011);
nand U4945 (N_4945,N_3519,N_3113);
nand U4946 (N_4946,N_4441,N_3241);
and U4947 (N_4947,N_3668,N_3760);
nand U4948 (N_4948,N_4407,N_3284);
nor U4949 (N_4949,N_3720,N_4000);
xor U4950 (N_4950,N_4434,N_3471);
and U4951 (N_4951,N_3948,N_3899);
and U4952 (N_4952,N_4224,N_3585);
or U4953 (N_4953,N_3012,N_4256);
nand U4954 (N_4954,N_4228,N_3152);
or U4955 (N_4955,N_3175,N_3542);
and U4956 (N_4956,N_3185,N_3216);
and U4957 (N_4957,N_4253,N_3852);
or U4958 (N_4958,N_4275,N_3851);
nor U4959 (N_4959,N_3568,N_4117);
nor U4960 (N_4960,N_3832,N_4472);
and U4961 (N_4961,N_4364,N_3635);
xor U4962 (N_4962,N_4027,N_3332);
xor U4963 (N_4963,N_3746,N_4120);
xor U4964 (N_4964,N_4025,N_3699);
nand U4965 (N_4965,N_3571,N_3540);
or U4966 (N_4966,N_3991,N_4341);
xnor U4967 (N_4967,N_4023,N_3124);
nand U4968 (N_4968,N_3271,N_4037);
xnor U4969 (N_4969,N_3622,N_4267);
and U4970 (N_4970,N_3283,N_4093);
xnor U4971 (N_4971,N_4495,N_3563);
xnor U4972 (N_4972,N_3338,N_3617);
nand U4973 (N_4973,N_4346,N_4084);
and U4974 (N_4974,N_3048,N_4231);
xor U4975 (N_4975,N_3580,N_4095);
and U4976 (N_4976,N_3711,N_3253);
nand U4977 (N_4977,N_4493,N_3364);
nand U4978 (N_4978,N_4463,N_3157);
nor U4979 (N_4979,N_4133,N_4369);
or U4980 (N_4980,N_4451,N_3163);
or U4981 (N_4981,N_4426,N_4450);
nand U4982 (N_4982,N_3679,N_3245);
and U4983 (N_4983,N_3474,N_3749);
xor U4984 (N_4984,N_3110,N_3658);
nand U4985 (N_4985,N_3455,N_4214);
or U4986 (N_4986,N_3768,N_4310);
nand U4987 (N_4987,N_4406,N_3714);
nand U4988 (N_4988,N_3748,N_4355);
nand U4989 (N_4989,N_3796,N_3025);
nor U4990 (N_4990,N_3988,N_3390);
xnor U4991 (N_4991,N_3266,N_4171);
nor U4992 (N_4992,N_3066,N_4206);
or U4993 (N_4993,N_4291,N_4288);
and U4994 (N_4994,N_3757,N_3367);
and U4995 (N_4995,N_4374,N_4050);
or U4996 (N_4996,N_3394,N_4116);
nor U4997 (N_4997,N_4233,N_3524);
and U4998 (N_4998,N_3530,N_4019);
xnor U4999 (N_4999,N_3019,N_4485);
nand U5000 (N_5000,N_3350,N_3811);
and U5001 (N_5001,N_3261,N_3846);
and U5002 (N_5002,N_3682,N_4193);
or U5003 (N_5003,N_3130,N_3797);
and U5004 (N_5004,N_4130,N_3188);
nand U5005 (N_5005,N_3576,N_4091);
nand U5006 (N_5006,N_3958,N_3021);
nor U5007 (N_5007,N_3392,N_3957);
nor U5008 (N_5008,N_3326,N_3565);
nand U5009 (N_5009,N_4138,N_3123);
nor U5010 (N_5010,N_3197,N_4013);
and U5011 (N_5011,N_3067,N_3439);
nor U5012 (N_5012,N_3357,N_3673);
nand U5013 (N_5013,N_3855,N_4055);
or U5014 (N_5014,N_3391,N_4074);
and U5015 (N_5015,N_3626,N_4387);
nand U5016 (N_5016,N_4251,N_3397);
or U5017 (N_5017,N_3994,N_4343);
nand U5018 (N_5018,N_3804,N_3996);
or U5019 (N_5019,N_3361,N_3373);
or U5020 (N_5020,N_3159,N_3451);
or U5021 (N_5021,N_4051,N_3737);
nor U5022 (N_5022,N_3770,N_3464);
or U5023 (N_5023,N_4259,N_4371);
nor U5024 (N_5024,N_4459,N_3226);
nand U5025 (N_5025,N_4268,N_4316);
nor U5026 (N_5026,N_3582,N_3089);
and U5027 (N_5027,N_4494,N_4385);
or U5028 (N_5028,N_3281,N_3595);
nand U5029 (N_5029,N_3184,N_3890);
nor U5030 (N_5030,N_3782,N_4211);
or U5031 (N_5031,N_3178,N_4252);
and U5032 (N_5032,N_3045,N_3671);
nor U5033 (N_5033,N_3529,N_3801);
or U5034 (N_5034,N_4360,N_4212);
xnor U5035 (N_5035,N_3053,N_4081);
and U5036 (N_5036,N_3718,N_3831);
nor U5037 (N_5037,N_4456,N_3003);
and U5038 (N_5038,N_4169,N_3942);
or U5039 (N_5039,N_4160,N_3717);
xnor U5040 (N_5040,N_3543,N_4155);
or U5041 (N_5041,N_3325,N_3421);
nor U5042 (N_5042,N_4039,N_3889);
nor U5043 (N_5043,N_3656,N_3229);
nand U5044 (N_5044,N_4004,N_3933);
nand U5045 (N_5045,N_3313,N_4238);
nand U5046 (N_5046,N_4487,N_3949);
nand U5047 (N_5047,N_3765,N_4225);
nand U5048 (N_5048,N_4393,N_3265);
nor U5049 (N_5049,N_4244,N_3459);
nor U5050 (N_5050,N_3605,N_3369);
nor U5051 (N_5051,N_4460,N_3819);
and U5052 (N_5052,N_3289,N_3549);
or U5053 (N_5053,N_3534,N_3486);
nand U5054 (N_5054,N_3535,N_3920);
and U5055 (N_5055,N_4068,N_4482);
or U5056 (N_5056,N_3026,N_4132);
and U5057 (N_5057,N_3440,N_3805);
and U5058 (N_5058,N_3676,N_3513);
nand U5059 (N_5059,N_4421,N_3792);
nand U5060 (N_5060,N_3608,N_3675);
nor U5061 (N_5061,N_4367,N_3240);
and U5062 (N_5062,N_4094,N_3842);
or U5063 (N_5063,N_3328,N_3201);
xnor U5064 (N_5064,N_3692,N_3376);
xor U5065 (N_5065,N_3141,N_4222);
nand U5066 (N_5066,N_3755,N_3912);
nand U5067 (N_5067,N_3706,N_3506);
nor U5068 (N_5068,N_3098,N_4137);
nor U5069 (N_5069,N_3039,N_4314);
and U5070 (N_5070,N_3902,N_3353);
nand U5071 (N_5071,N_4392,N_4373);
or U5072 (N_5072,N_3387,N_4153);
nand U5073 (N_5073,N_4248,N_3294);
and U5074 (N_5074,N_3420,N_4178);
and U5075 (N_5075,N_3042,N_3267);
and U5076 (N_5076,N_4478,N_3643);
xnor U5077 (N_5077,N_3469,N_3531);
nand U5078 (N_5078,N_3491,N_3237);
nor U5079 (N_5079,N_3818,N_3099);
or U5080 (N_5080,N_4272,N_4179);
nor U5081 (N_5081,N_4484,N_4018);
xor U5082 (N_5082,N_4157,N_3200);
nor U5083 (N_5083,N_4240,N_3669);
or U5084 (N_5084,N_3891,N_3017);
nand U5085 (N_5085,N_3236,N_3000);
or U5086 (N_5086,N_3122,N_3366);
and U5087 (N_5087,N_3375,N_3162);
and U5088 (N_5088,N_3700,N_3170);
and U5089 (N_5089,N_3462,N_3071);
and U5090 (N_5090,N_4134,N_3024);
or U5091 (N_5091,N_3570,N_3581);
nand U5092 (N_5092,N_3254,N_4203);
nand U5093 (N_5093,N_3255,N_3709);
and U5094 (N_5094,N_3843,N_4141);
nor U5095 (N_5095,N_4200,N_3072);
or U5096 (N_5096,N_4058,N_4471);
nor U5097 (N_5097,N_3481,N_3710);
nand U5098 (N_5098,N_3203,N_3386);
or U5099 (N_5099,N_3861,N_3959);
nand U5100 (N_5100,N_3196,N_3424);
nor U5101 (N_5101,N_3572,N_3103);
nand U5102 (N_5102,N_4219,N_4036);
and U5103 (N_5103,N_3973,N_3738);
and U5104 (N_5104,N_3242,N_3111);
nand U5105 (N_5105,N_3931,N_4124);
and U5106 (N_5106,N_3028,N_4318);
or U5107 (N_5107,N_4488,N_4344);
and U5108 (N_5108,N_3864,N_3965);
xnor U5109 (N_5109,N_3400,N_3917);
nand U5110 (N_5110,N_3564,N_4009);
or U5111 (N_5111,N_3140,N_4323);
and U5112 (N_5112,N_3632,N_3106);
nor U5113 (N_5113,N_3546,N_4237);
nor U5114 (N_5114,N_3448,N_4303);
nor U5115 (N_5115,N_3587,N_3769);
or U5116 (N_5116,N_3079,N_3654);
nand U5117 (N_5117,N_3191,N_4131);
xnor U5118 (N_5118,N_3521,N_4430);
or U5119 (N_5119,N_3716,N_3655);
or U5120 (N_5120,N_4115,N_3475);
nand U5121 (N_5121,N_3403,N_4496);
xor U5122 (N_5122,N_3441,N_3133);
nand U5123 (N_5123,N_4408,N_4227);
nor U5124 (N_5124,N_3212,N_3925);
nor U5125 (N_5125,N_3498,N_3468);
and U5126 (N_5126,N_3404,N_3841);
or U5127 (N_5127,N_4122,N_4328);
or U5128 (N_5128,N_3895,N_4417);
and U5129 (N_5129,N_4194,N_4184);
nor U5130 (N_5130,N_3900,N_4056);
or U5131 (N_5131,N_3558,N_3292);
xor U5132 (N_5132,N_3978,N_4331);
xor U5133 (N_5133,N_3116,N_3883);
nor U5134 (N_5134,N_3168,N_4026);
and U5135 (N_5135,N_3034,N_4283);
nor U5136 (N_5136,N_3174,N_3502);
nor U5137 (N_5137,N_3158,N_3729);
nor U5138 (N_5138,N_3318,N_3252);
or U5139 (N_5139,N_4089,N_3645);
xnor U5140 (N_5140,N_4322,N_3093);
and U5141 (N_5141,N_4016,N_3182);
nand U5142 (N_5142,N_3827,N_3363);
nor U5143 (N_5143,N_4366,N_3452);
nand U5144 (N_5144,N_3662,N_3809);
xnor U5145 (N_5145,N_3734,N_3926);
nor U5146 (N_5146,N_3259,N_3910);
or U5147 (N_5147,N_3470,N_3609);
nand U5148 (N_5148,N_3210,N_4416);
nand U5149 (N_5149,N_3616,N_3520);
and U5150 (N_5150,N_3732,N_3466);
or U5151 (N_5151,N_3590,N_3275);
nand U5152 (N_5152,N_4059,N_3694);
or U5153 (N_5153,N_3850,N_3465);
nor U5154 (N_5154,N_3145,N_3863);
xnor U5155 (N_5155,N_4474,N_3004);
and U5156 (N_5156,N_4263,N_3380);
nand U5157 (N_5157,N_3892,N_4464);
nor U5158 (N_5158,N_4079,N_4483);
nor U5159 (N_5159,N_4278,N_3993);
nand U5160 (N_5160,N_4420,N_3314);
or U5161 (N_5161,N_3813,N_4167);
nand U5162 (N_5162,N_4319,N_3078);
or U5163 (N_5163,N_3137,N_4052);
and U5164 (N_5164,N_4381,N_4394);
and U5165 (N_5165,N_3411,N_3291);
nor U5166 (N_5166,N_3036,N_3477);
or U5167 (N_5167,N_3997,N_3857);
and U5168 (N_5168,N_4397,N_3763);
and U5169 (N_5169,N_3955,N_3406);
and U5170 (N_5170,N_3244,N_3333);
nor U5171 (N_5171,N_3510,N_3461);
and U5172 (N_5172,N_4189,N_4352);
nand U5173 (N_5173,N_3541,N_4168);
or U5174 (N_5174,N_3637,N_3887);
nand U5175 (N_5175,N_3046,N_3579);
nand U5176 (N_5176,N_3876,N_4078);
and U5177 (N_5177,N_4060,N_3211);
or U5178 (N_5178,N_3788,N_3791);
and U5179 (N_5179,N_4057,N_3374);
xor U5180 (N_5180,N_4190,N_3975);
or U5181 (N_5181,N_3488,N_3834);
and U5182 (N_5182,N_3589,N_4302);
and U5183 (N_5183,N_4176,N_4069);
nor U5184 (N_5184,N_3224,N_3378);
or U5185 (N_5185,N_3074,N_3947);
nor U5186 (N_5186,N_3383,N_4409);
and U5187 (N_5187,N_3728,N_3777);
or U5188 (N_5188,N_4461,N_3756);
nand U5189 (N_5189,N_3575,N_4015);
and U5190 (N_5190,N_3323,N_4277);
and U5191 (N_5191,N_3249,N_3080);
nor U5192 (N_5192,N_4010,N_3115);
or U5193 (N_5193,N_3584,N_4188);
xor U5194 (N_5194,N_4378,N_3800);
or U5195 (N_5195,N_4041,N_4480);
and U5196 (N_5196,N_3599,N_3125);
or U5197 (N_5197,N_4306,N_4414);
nor U5198 (N_5198,N_3334,N_4187);
nor U5199 (N_5199,N_4145,N_3946);
or U5200 (N_5200,N_4388,N_3160);
nand U5201 (N_5201,N_3060,N_3295);
xnor U5202 (N_5202,N_3429,N_3614);
or U5203 (N_5203,N_4182,N_3509);
xnor U5204 (N_5204,N_3248,N_3937);
and U5205 (N_5205,N_3793,N_4432);
and U5206 (N_5206,N_3727,N_3129);
or U5207 (N_5207,N_3983,N_3533);
nor U5208 (N_5208,N_4337,N_3222);
and U5209 (N_5209,N_4258,N_3399);
nand U5210 (N_5210,N_4415,N_4380);
nor U5211 (N_5211,N_3207,N_4085);
nand U5212 (N_5212,N_3143,N_3285);
nand U5213 (N_5213,N_4467,N_4498);
and U5214 (N_5214,N_3341,N_4363);
xor U5215 (N_5215,N_3835,N_4307);
nor U5216 (N_5216,N_4400,N_3227);
nand U5217 (N_5217,N_3569,N_3215);
nor U5218 (N_5218,N_3329,N_3002);
nor U5219 (N_5219,N_3573,N_4271);
nand U5220 (N_5220,N_4326,N_3198);
nand U5221 (N_5221,N_4046,N_4099);
and U5222 (N_5222,N_4045,N_4230);
and U5223 (N_5223,N_3976,N_4100);
nor U5224 (N_5224,N_3880,N_3862);
nand U5225 (N_5225,N_3879,N_4092);
nor U5226 (N_5226,N_3945,N_4110);
or U5227 (N_5227,N_3620,N_3362);
or U5228 (N_5228,N_3816,N_3893);
nor U5229 (N_5229,N_3001,N_3315);
nor U5230 (N_5230,N_4128,N_4490);
nor U5231 (N_5231,N_3553,N_3886);
nand U5232 (N_5232,N_3037,N_3172);
nor U5233 (N_5233,N_4391,N_3736);
nor U5234 (N_5234,N_3844,N_4410);
or U5235 (N_5235,N_3164,N_3812);
and U5236 (N_5236,N_3435,N_3473);
and U5237 (N_5237,N_3038,N_3467);
and U5238 (N_5238,N_3304,N_3398);
or U5239 (N_5239,N_4108,N_3539);
or U5240 (N_5240,N_4151,N_3623);
nand U5241 (N_5241,N_3904,N_3436);
nand U5242 (N_5242,N_4213,N_3629);
or U5243 (N_5243,N_3532,N_4470);
and U5244 (N_5244,N_3199,N_4334);
xor U5245 (N_5245,N_4185,N_4279);
xnor U5246 (N_5246,N_3824,N_4255);
nand U5247 (N_5247,N_3035,N_3779);
and U5248 (N_5248,N_3712,N_3713);
nand U5249 (N_5249,N_4207,N_3075);
nand U5250 (N_5250,N_4274,N_3841);
xnor U5251 (N_5251,N_3455,N_4181);
or U5252 (N_5252,N_3199,N_4185);
nand U5253 (N_5253,N_3190,N_4094);
and U5254 (N_5254,N_4426,N_3617);
nand U5255 (N_5255,N_3217,N_3177);
nand U5256 (N_5256,N_4362,N_3306);
nor U5257 (N_5257,N_4324,N_4443);
xnor U5258 (N_5258,N_3671,N_4185);
or U5259 (N_5259,N_3819,N_3625);
nor U5260 (N_5260,N_3697,N_4223);
xnor U5261 (N_5261,N_4007,N_3216);
nand U5262 (N_5262,N_3674,N_4402);
xnor U5263 (N_5263,N_3997,N_3592);
nand U5264 (N_5264,N_4106,N_3826);
or U5265 (N_5265,N_3391,N_3615);
nand U5266 (N_5266,N_4029,N_3090);
or U5267 (N_5267,N_3076,N_4222);
nor U5268 (N_5268,N_3807,N_3367);
nand U5269 (N_5269,N_3256,N_3515);
nor U5270 (N_5270,N_3870,N_3109);
nand U5271 (N_5271,N_3514,N_4302);
nor U5272 (N_5272,N_3444,N_3485);
or U5273 (N_5273,N_4015,N_3401);
nor U5274 (N_5274,N_4296,N_3976);
and U5275 (N_5275,N_3409,N_4401);
and U5276 (N_5276,N_3844,N_3587);
and U5277 (N_5277,N_4435,N_3893);
or U5278 (N_5278,N_4138,N_3116);
or U5279 (N_5279,N_3520,N_4272);
nand U5280 (N_5280,N_3274,N_4376);
or U5281 (N_5281,N_3275,N_3982);
nor U5282 (N_5282,N_4183,N_3142);
or U5283 (N_5283,N_3804,N_3148);
and U5284 (N_5284,N_3133,N_3693);
or U5285 (N_5285,N_4080,N_4127);
and U5286 (N_5286,N_3012,N_4125);
and U5287 (N_5287,N_3753,N_3025);
and U5288 (N_5288,N_3140,N_3740);
nor U5289 (N_5289,N_3554,N_3377);
nand U5290 (N_5290,N_3195,N_4477);
nor U5291 (N_5291,N_3276,N_3560);
nor U5292 (N_5292,N_3119,N_3063);
nand U5293 (N_5293,N_4272,N_3062);
nand U5294 (N_5294,N_3528,N_3672);
or U5295 (N_5295,N_3924,N_3858);
or U5296 (N_5296,N_3302,N_3602);
and U5297 (N_5297,N_4435,N_4032);
nor U5298 (N_5298,N_4272,N_3456);
nor U5299 (N_5299,N_3535,N_4000);
and U5300 (N_5300,N_4238,N_3317);
and U5301 (N_5301,N_3392,N_4394);
nand U5302 (N_5302,N_3164,N_3263);
or U5303 (N_5303,N_4085,N_4009);
and U5304 (N_5304,N_3217,N_4316);
xnor U5305 (N_5305,N_4125,N_4005);
and U5306 (N_5306,N_4338,N_4216);
nor U5307 (N_5307,N_3530,N_3590);
and U5308 (N_5308,N_4246,N_3807);
nor U5309 (N_5309,N_3244,N_3330);
nand U5310 (N_5310,N_4206,N_3145);
or U5311 (N_5311,N_3109,N_3657);
nand U5312 (N_5312,N_3863,N_3016);
nand U5313 (N_5313,N_3721,N_4068);
nand U5314 (N_5314,N_3434,N_3311);
and U5315 (N_5315,N_3711,N_4057);
xor U5316 (N_5316,N_4434,N_3705);
and U5317 (N_5317,N_3347,N_4174);
and U5318 (N_5318,N_3509,N_3206);
nand U5319 (N_5319,N_3395,N_3254);
or U5320 (N_5320,N_4249,N_3081);
nand U5321 (N_5321,N_4402,N_4043);
and U5322 (N_5322,N_4219,N_3769);
nand U5323 (N_5323,N_3125,N_3462);
nand U5324 (N_5324,N_4013,N_3915);
and U5325 (N_5325,N_4208,N_4014);
and U5326 (N_5326,N_3237,N_3980);
xnor U5327 (N_5327,N_3836,N_3075);
nand U5328 (N_5328,N_4153,N_4215);
nand U5329 (N_5329,N_4268,N_3943);
nand U5330 (N_5330,N_3959,N_3167);
and U5331 (N_5331,N_3334,N_3981);
nor U5332 (N_5332,N_4465,N_3632);
nor U5333 (N_5333,N_3957,N_3027);
nand U5334 (N_5334,N_4295,N_3463);
nand U5335 (N_5335,N_3654,N_3314);
and U5336 (N_5336,N_4344,N_4092);
and U5337 (N_5337,N_3396,N_3766);
nor U5338 (N_5338,N_4453,N_3413);
and U5339 (N_5339,N_3486,N_3474);
nand U5340 (N_5340,N_3523,N_4105);
xor U5341 (N_5341,N_3074,N_3753);
and U5342 (N_5342,N_3467,N_3324);
or U5343 (N_5343,N_3632,N_3228);
or U5344 (N_5344,N_4382,N_4221);
xnor U5345 (N_5345,N_3558,N_3283);
and U5346 (N_5346,N_3512,N_3851);
xor U5347 (N_5347,N_3525,N_3549);
nand U5348 (N_5348,N_3569,N_3680);
nor U5349 (N_5349,N_3686,N_3547);
nor U5350 (N_5350,N_3727,N_3246);
xor U5351 (N_5351,N_3947,N_3000);
nor U5352 (N_5352,N_4494,N_4357);
or U5353 (N_5353,N_3058,N_4400);
nand U5354 (N_5354,N_3416,N_4452);
nand U5355 (N_5355,N_4261,N_4383);
or U5356 (N_5356,N_3074,N_3770);
xnor U5357 (N_5357,N_3255,N_3254);
nor U5358 (N_5358,N_3861,N_3462);
or U5359 (N_5359,N_4323,N_4152);
or U5360 (N_5360,N_3247,N_3173);
nand U5361 (N_5361,N_4189,N_3383);
nand U5362 (N_5362,N_3044,N_3432);
or U5363 (N_5363,N_3638,N_3725);
xor U5364 (N_5364,N_3021,N_3990);
and U5365 (N_5365,N_3445,N_4234);
nand U5366 (N_5366,N_3370,N_3736);
nand U5367 (N_5367,N_4131,N_3006);
and U5368 (N_5368,N_4053,N_3864);
and U5369 (N_5369,N_4055,N_3191);
xor U5370 (N_5370,N_3641,N_3274);
nor U5371 (N_5371,N_3836,N_3323);
xor U5372 (N_5372,N_4411,N_3164);
and U5373 (N_5373,N_3709,N_3654);
nor U5374 (N_5374,N_3037,N_4017);
nand U5375 (N_5375,N_3343,N_3041);
nand U5376 (N_5376,N_4341,N_3559);
nand U5377 (N_5377,N_4151,N_4321);
nor U5378 (N_5378,N_3127,N_4465);
nor U5379 (N_5379,N_3927,N_4169);
nor U5380 (N_5380,N_4193,N_3746);
and U5381 (N_5381,N_3691,N_4112);
or U5382 (N_5382,N_4078,N_4430);
xor U5383 (N_5383,N_4110,N_4416);
nand U5384 (N_5384,N_3751,N_4018);
nor U5385 (N_5385,N_4149,N_3306);
or U5386 (N_5386,N_3556,N_4075);
nor U5387 (N_5387,N_3221,N_3824);
nand U5388 (N_5388,N_3979,N_3997);
nor U5389 (N_5389,N_3643,N_4129);
and U5390 (N_5390,N_3465,N_4167);
nor U5391 (N_5391,N_3543,N_3145);
xnor U5392 (N_5392,N_3424,N_3400);
or U5393 (N_5393,N_3255,N_3100);
xnor U5394 (N_5394,N_4337,N_3697);
or U5395 (N_5395,N_3720,N_3257);
or U5396 (N_5396,N_3506,N_4427);
and U5397 (N_5397,N_3812,N_3624);
or U5398 (N_5398,N_3335,N_4446);
and U5399 (N_5399,N_4049,N_3302);
and U5400 (N_5400,N_4232,N_4245);
or U5401 (N_5401,N_3037,N_3539);
nand U5402 (N_5402,N_3917,N_4460);
and U5403 (N_5403,N_4434,N_3291);
nor U5404 (N_5404,N_4291,N_3726);
nor U5405 (N_5405,N_3016,N_3054);
nor U5406 (N_5406,N_4248,N_3464);
or U5407 (N_5407,N_3502,N_3625);
nor U5408 (N_5408,N_4085,N_3834);
or U5409 (N_5409,N_3680,N_4374);
or U5410 (N_5410,N_3359,N_4056);
nand U5411 (N_5411,N_3081,N_4367);
nand U5412 (N_5412,N_4182,N_3483);
nand U5413 (N_5413,N_3366,N_3541);
nor U5414 (N_5414,N_3753,N_3003);
or U5415 (N_5415,N_3961,N_3262);
nor U5416 (N_5416,N_4151,N_3063);
xnor U5417 (N_5417,N_3680,N_4052);
xor U5418 (N_5418,N_4382,N_4202);
and U5419 (N_5419,N_4402,N_4498);
nand U5420 (N_5420,N_3957,N_4424);
nand U5421 (N_5421,N_4124,N_3620);
or U5422 (N_5422,N_3939,N_4250);
or U5423 (N_5423,N_3376,N_3837);
xnor U5424 (N_5424,N_4201,N_3670);
or U5425 (N_5425,N_4446,N_3537);
xnor U5426 (N_5426,N_4348,N_4471);
or U5427 (N_5427,N_3303,N_4257);
and U5428 (N_5428,N_3543,N_4219);
nand U5429 (N_5429,N_3412,N_3255);
nand U5430 (N_5430,N_3356,N_3359);
nor U5431 (N_5431,N_3035,N_3750);
or U5432 (N_5432,N_4432,N_3903);
nand U5433 (N_5433,N_3605,N_3830);
nor U5434 (N_5434,N_3457,N_4394);
xor U5435 (N_5435,N_4079,N_3939);
nor U5436 (N_5436,N_4049,N_3691);
nand U5437 (N_5437,N_4242,N_4278);
nor U5438 (N_5438,N_4265,N_3408);
nor U5439 (N_5439,N_4488,N_3859);
and U5440 (N_5440,N_3482,N_3747);
or U5441 (N_5441,N_3107,N_3749);
or U5442 (N_5442,N_3781,N_3147);
or U5443 (N_5443,N_3117,N_3691);
nor U5444 (N_5444,N_4045,N_3409);
nand U5445 (N_5445,N_4109,N_3062);
xnor U5446 (N_5446,N_3549,N_4369);
and U5447 (N_5447,N_4490,N_3287);
nand U5448 (N_5448,N_3931,N_4346);
nor U5449 (N_5449,N_3545,N_3734);
and U5450 (N_5450,N_4273,N_3329);
and U5451 (N_5451,N_3547,N_3928);
or U5452 (N_5452,N_3741,N_3284);
or U5453 (N_5453,N_4409,N_3046);
and U5454 (N_5454,N_3926,N_4442);
or U5455 (N_5455,N_3377,N_3096);
and U5456 (N_5456,N_3993,N_3533);
nor U5457 (N_5457,N_3923,N_3603);
xor U5458 (N_5458,N_3415,N_4290);
or U5459 (N_5459,N_3263,N_3332);
or U5460 (N_5460,N_3560,N_3833);
nor U5461 (N_5461,N_3019,N_3044);
xor U5462 (N_5462,N_4370,N_4008);
or U5463 (N_5463,N_4075,N_3906);
nor U5464 (N_5464,N_4163,N_4378);
nor U5465 (N_5465,N_4038,N_3952);
xor U5466 (N_5466,N_3507,N_4039);
nand U5467 (N_5467,N_3163,N_3912);
nand U5468 (N_5468,N_3076,N_3491);
and U5469 (N_5469,N_3905,N_3281);
nor U5470 (N_5470,N_4265,N_3546);
or U5471 (N_5471,N_3603,N_3326);
nand U5472 (N_5472,N_3491,N_3015);
and U5473 (N_5473,N_3719,N_4480);
nand U5474 (N_5474,N_3116,N_3177);
xor U5475 (N_5475,N_3236,N_4388);
nand U5476 (N_5476,N_3281,N_3400);
or U5477 (N_5477,N_4423,N_4433);
nand U5478 (N_5478,N_3613,N_3796);
nand U5479 (N_5479,N_4426,N_4222);
nor U5480 (N_5480,N_3128,N_3052);
nand U5481 (N_5481,N_3380,N_4439);
and U5482 (N_5482,N_4446,N_3865);
or U5483 (N_5483,N_4155,N_3353);
nand U5484 (N_5484,N_3911,N_4311);
nor U5485 (N_5485,N_3491,N_4127);
nor U5486 (N_5486,N_4301,N_3705);
and U5487 (N_5487,N_3750,N_3730);
nor U5488 (N_5488,N_3847,N_4334);
or U5489 (N_5489,N_4450,N_4400);
and U5490 (N_5490,N_3174,N_3913);
nor U5491 (N_5491,N_4483,N_3246);
or U5492 (N_5492,N_3583,N_4397);
and U5493 (N_5493,N_3434,N_3849);
or U5494 (N_5494,N_4051,N_4443);
xor U5495 (N_5495,N_4059,N_3573);
or U5496 (N_5496,N_3965,N_4420);
nand U5497 (N_5497,N_3720,N_3775);
nand U5498 (N_5498,N_3776,N_4137);
or U5499 (N_5499,N_3843,N_3761);
or U5500 (N_5500,N_3136,N_3578);
and U5501 (N_5501,N_4294,N_3950);
and U5502 (N_5502,N_3912,N_3292);
and U5503 (N_5503,N_4115,N_4284);
nor U5504 (N_5504,N_4189,N_4172);
and U5505 (N_5505,N_3561,N_4079);
nor U5506 (N_5506,N_4276,N_4016);
and U5507 (N_5507,N_3019,N_4242);
and U5508 (N_5508,N_3161,N_3954);
or U5509 (N_5509,N_4457,N_4347);
xor U5510 (N_5510,N_4430,N_3749);
nor U5511 (N_5511,N_3733,N_3010);
or U5512 (N_5512,N_3341,N_3814);
or U5513 (N_5513,N_4491,N_3574);
or U5514 (N_5514,N_3584,N_4106);
or U5515 (N_5515,N_3142,N_4188);
or U5516 (N_5516,N_3662,N_3648);
nor U5517 (N_5517,N_3546,N_3948);
nand U5518 (N_5518,N_3176,N_3791);
nand U5519 (N_5519,N_3861,N_4319);
nor U5520 (N_5520,N_3732,N_3233);
and U5521 (N_5521,N_3540,N_3229);
nor U5522 (N_5522,N_3438,N_4043);
or U5523 (N_5523,N_4216,N_3606);
and U5524 (N_5524,N_3383,N_4494);
and U5525 (N_5525,N_3676,N_4322);
nand U5526 (N_5526,N_3655,N_3758);
and U5527 (N_5527,N_4210,N_4013);
nor U5528 (N_5528,N_3381,N_4226);
and U5529 (N_5529,N_3220,N_3267);
or U5530 (N_5530,N_3669,N_3794);
and U5531 (N_5531,N_4178,N_4003);
and U5532 (N_5532,N_3413,N_3538);
nor U5533 (N_5533,N_3392,N_4477);
or U5534 (N_5534,N_3075,N_4472);
xnor U5535 (N_5535,N_3819,N_3905);
and U5536 (N_5536,N_3244,N_3969);
nor U5537 (N_5537,N_3953,N_3614);
nor U5538 (N_5538,N_4026,N_3209);
nand U5539 (N_5539,N_4169,N_3569);
xor U5540 (N_5540,N_4433,N_3239);
nand U5541 (N_5541,N_4084,N_3354);
nand U5542 (N_5542,N_3739,N_4315);
or U5543 (N_5543,N_3038,N_3175);
or U5544 (N_5544,N_3700,N_4460);
or U5545 (N_5545,N_4108,N_3784);
or U5546 (N_5546,N_4230,N_4315);
and U5547 (N_5547,N_4422,N_4093);
nand U5548 (N_5548,N_4147,N_4292);
and U5549 (N_5549,N_3674,N_3026);
and U5550 (N_5550,N_4316,N_3074);
nand U5551 (N_5551,N_3917,N_3122);
and U5552 (N_5552,N_4398,N_4121);
or U5553 (N_5553,N_4175,N_4102);
or U5554 (N_5554,N_3909,N_3078);
xor U5555 (N_5555,N_3738,N_3200);
and U5556 (N_5556,N_3738,N_4429);
or U5557 (N_5557,N_3016,N_4066);
nor U5558 (N_5558,N_3627,N_3651);
xor U5559 (N_5559,N_3970,N_3789);
and U5560 (N_5560,N_3176,N_4384);
nand U5561 (N_5561,N_4068,N_3728);
xnor U5562 (N_5562,N_3720,N_3165);
nand U5563 (N_5563,N_3792,N_3880);
nor U5564 (N_5564,N_3776,N_4037);
nor U5565 (N_5565,N_4361,N_3528);
xor U5566 (N_5566,N_3407,N_3619);
nor U5567 (N_5567,N_3645,N_3932);
nor U5568 (N_5568,N_3586,N_3789);
and U5569 (N_5569,N_3224,N_3177);
or U5570 (N_5570,N_3778,N_3444);
or U5571 (N_5571,N_3980,N_3249);
nor U5572 (N_5572,N_4029,N_4073);
nor U5573 (N_5573,N_3334,N_3661);
xnor U5574 (N_5574,N_3753,N_4329);
and U5575 (N_5575,N_4413,N_3156);
xor U5576 (N_5576,N_3322,N_3064);
or U5577 (N_5577,N_3366,N_3261);
nand U5578 (N_5578,N_4155,N_3984);
xnor U5579 (N_5579,N_3975,N_3377);
or U5580 (N_5580,N_3406,N_3054);
nand U5581 (N_5581,N_4079,N_3332);
and U5582 (N_5582,N_3563,N_4082);
or U5583 (N_5583,N_3461,N_3932);
and U5584 (N_5584,N_4404,N_3856);
nand U5585 (N_5585,N_3759,N_4093);
nor U5586 (N_5586,N_3047,N_3437);
and U5587 (N_5587,N_4380,N_3409);
and U5588 (N_5588,N_3636,N_4389);
nand U5589 (N_5589,N_3373,N_4352);
nand U5590 (N_5590,N_3048,N_4125);
or U5591 (N_5591,N_3415,N_4124);
xor U5592 (N_5592,N_3139,N_3955);
nor U5593 (N_5593,N_3788,N_3312);
nor U5594 (N_5594,N_3475,N_4436);
nand U5595 (N_5595,N_3074,N_4038);
nor U5596 (N_5596,N_3349,N_3161);
or U5597 (N_5597,N_4468,N_4045);
nor U5598 (N_5598,N_3537,N_4066);
and U5599 (N_5599,N_3823,N_3668);
nor U5600 (N_5600,N_3162,N_3157);
nor U5601 (N_5601,N_3624,N_3607);
or U5602 (N_5602,N_3561,N_3528);
or U5603 (N_5603,N_4066,N_3684);
nand U5604 (N_5604,N_4097,N_3921);
nand U5605 (N_5605,N_3171,N_3973);
nand U5606 (N_5606,N_3410,N_3066);
and U5607 (N_5607,N_3363,N_3164);
xor U5608 (N_5608,N_3140,N_4456);
and U5609 (N_5609,N_3015,N_3131);
nand U5610 (N_5610,N_3028,N_3250);
and U5611 (N_5611,N_3020,N_3973);
and U5612 (N_5612,N_4364,N_3863);
nor U5613 (N_5613,N_4177,N_4386);
and U5614 (N_5614,N_3966,N_3355);
nor U5615 (N_5615,N_3952,N_3424);
and U5616 (N_5616,N_3454,N_3690);
or U5617 (N_5617,N_3889,N_4282);
and U5618 (N_5618,N_4248,N_4356);
nand U5619 (N_5619,N_3735,N_3759);
nand U5620 (N_5620,N_3591,N_3917);
and U5621 (N_5621,N_3350,N_3650);
nand U5622 (N_5622,N_3910,N_3563);
xor U5623 (N_5623,N_4030,N_3945);
and U5624 (N_5624,N_3909,N_4012);
xnor U5625 (N_5625,N_4201,N_3464);
xor U5626 (N_5626,N_3899,N_3148);
or U5627 (N_5627,N_4462,N_4275);
nand U5628 (N_5628,N_3217,N_4246);
nand U5629 (N_5629,N_3219,N_4387);
and U5630 (N_5630,N_4421,N_4437);
and U5631 (N_5631,N_3700,N_3025);
nand U5632 (N_5632,N_3348,N_4419);
and U5633 (N_5633,N_3668,N_4178);
and U5634 (N_5634,N_3191,N_3282);
or U5635 (N_5635,N_3382,N_4447);
xnor U5636 (N_5636,N_3405,N_3288);
nand U5637 (N_5637,N_3473,N_4274);
nand U5638 (N_5638,N_4021,N_4280);
and U5639 (N_5639,N_4072,N_3278);
and U5640 (N_5640,N_4380,N_3096);
or U5641 (N_5641,N_3512,N_3813);
xnor U5642 (N_5642,N_4164,N_3508);
nor U5643 (N_5643,N_3070,N_3382);
and U5644 (N_5644,N_3327,N_3921);
or U5645 (N_5645,N_3602,N_4172);
and U5646 (N_5646,N_3251,N_3839);
nand U5647 (N_5647,N_3213,N_3719);
xnor U5648 (N_5648,N_3600,N_3381);
or U5649 (N_5649,N_3744,N_3602);
and U5650 (N_5650,N_4036,N_3455);
nor U5651 (N_5651,N_3536,N_3086);
nand U5652 (N_5652,N_4206,N_3360);
or U5653 (N_5653,N_3268,N_3625);
nand U5654 (N_5654,N_4059,N_4353);
or U5655 (N_5655,N_3243,N_3477);
nor U5656 (N_5656,N_4174,N_3160);
and U5657 (N_5657,N_3374,N_3266);
xor U5658 (N_5658,N_3099,N_3289);
and U5659 (N_5659,N_3635,N_3143);
or U5660 (N_5660,N_4385,N_3026);
xor U5661 (N_5661,N_4329,N_3465);
or U5662 (N_5662,N_3673,N_3869);
nor U5663 (N_5663,N_4238,N_3435);
or U5664 (N_5664,N_4003,N_4222);
nand U5665 (N_5665,N_3480,N_4425);
and U5666 (N_5666,N_3728,N_3274);
nand U5667 (N_5667,N_3397,N_3611);
or U5668 (N_5668,N_4370,N_3123);
and U5669 (N_5669,N_4201,N_3058);
and U5670 (N_5670,N_4434,N_3569);
and U5671 (N_5671,N_4196,N_3297);
nor U5672 (N_5672,N_3667,N_3060);
nor U5673 (N_5673,N_3864,N_4323);
xnor U5674 (N_5674,N_4253,N_3346);
nand U5675 (N_5675,N_3231,N_3586);
nor U5676 (N_5676,N_4172,N_4141);
and U5677 (N_5677,N_3638,N_3203);
and U5678 (N_5678,N_3256,N_3374);
nor U5679 (N_5679,N_4012,N_4258);
nand U5680 (N_5680,N_3858,N_3972);
or U5681 (N_5681,N_3981,N_4210);
and U5682 (N_5682,N_4366,N_3491);
nor U5683 (N_5683,N_3889,N_3304);
nor U5684 (N_5684,N_3682,N_3640);
xnor U5685 (N_5685,N_3430,N_4247);
or U5686 (N_5686,N_3820,N_4176);
and U5687 (N_5687,N_3373,N_3503);
and U5688 (N_5688,N_4260,N_3866);
and U5689 (N_5689,N_4330,N_4263);
nor U5690 (N_5690,N_4017,N_3521);
xnor U5691 (N_5691,N_4368,N_4190);
nand U5692 (N_5692,N_4461,N_3657);
nand U5693 (N_5693,N_4339,N_3399);
or U5694 (N_5694,N_4263,N_3860);
xor U5695 (N_5695,N_3153,N_4484);
and U5696 (N_5696,N_3082,N_3325);
or U5697 (N_5697,N_3396,N_4139);
and U5698 (N_5698,N_3598,N_4445);
or U5699 (N_5699,N_3663,N_3588);
nor U5700 (N_5700,N_3598,N_3009);
nor U5701 (N_5701,N_3841,N_3115);
nand U5702 (N_5702,N_3268,N_3859);
nand U5703 (N_5703,N_4151,N_3465);
nor U5704 (N_5704,N_3802,N_4355);
nand U5705 (N_5705,N_3211,N_3506);
or U5706 (N_5706,N_4349,N_3114);
nand U5707 (N_5707,N_3240,N_3386);
nor U5708 (N_5708,N_3017,N_4127);
nor U5709 (N_5709,N_3838,N_4180);
nand U5710 (N_5710,N_4186,N_3240);
and U5711 (N_5711,N_3333,N_3425);
nor U5712 (N_5712,N_4295,N_4435);
nand U5713 (N_5713,N_4006,N_3763);
nand U5714 (N_5714,N_4288,N_3198);
nand U5715 (N_5715,N_3626,N_3441);
and U5716 (N_5716,N_4358,N_4010);
nand U5717 (N_5717,N_3419,N_3564);
and U5718 (N_5718,N_3811,N_3846);
nand U5719 (N_5719,N_3427,N_3153);
or U5720 (N_5720,N_3264,N_3569);
or U5721 (N_5721,N_3676,N_3152);
nor U5722 (N_5722,N_3087,N_3571);
nor U5723 (N_5723,N_3091,N_3736);
xor U5724 (N_5724,N_3155,N_3227);
nor U5725 (N_5725,N_3182,N_4169);
nor U5726 (N_5726,N_4173,N_3831);
xor U5727 (N_5727,N_3485,N_3260);
and U5728 (N_5728,N_4387,N_4263);
and U5729 (N_5729,N_4166,N_3664);
nand U5730 (N_5730,N_3969,N_3653);
nand U5731 (N_5731,N_4021,N_3226);
and U5732 (N_5732,N_4367,N_3477);
nor U5733 (N_5733,N_3268,N_3237);
xnor U5734 (N_5734,N_3606,N_4308);
or U5735 (N_5735,N_4186,N_3264);
and U5736 (N_5736,N_3025,N_3612);
and U5737 (N_5737,N_4059,N_3145);
or U5738 (N_5738,N_4108,N_4071);
or U5739 (N_5739,N_3456,N_4226);
nor U5740 (N_5740,N_3776,N_3099);
xnor U5741 (N_5741,N_3076,N_3901);
nor U5742 (N_5742,N_3988,N_3731);
nor U5743 (N_5743,N_3248,N_3726);
nand U5744 (N_5744,N_3135,N_4188);
nand U5745 (N_5745,N_3814,N_4338);
nor U5746 (N_5746,N_3259,N_3575);
nand U5747 (N_5747,N_4180,N_4315);
and U5748 (N_5748,N_4276,N_3075);
nor U5749 (N_5749,N_4037,N_3654);
nand U5750 (N_5750,N_4025,N_3264);
nor U5751 (N_5751,N_3726,N_3799);
nor U5752 (N_5752,N_4490,N_4347);
xnor U5753 (N_5753,N_3816,N_4492);
and U5754 (N_5754,N_3201,N_3719);
and U5755 (N_5755,N_3501,N_3232);
or U5756 (N_5756,N_3434,N_4205);
and U5757 (N_5757,N_3075,N_3032);
nor U5758 (N_5758,N_3091,N_3887);
xor U5759 (N_5759,N_4041,N_3602);
and U5760 (N_5760,N_3491,N_3347);
or U5761 (N_5761,N_3360,N_4105);
nand U5762 (N_5762,N_4219,N_3674);
or U5763 (N_5763,N_4268,N_4113);
nand U5764 (N_5764,N_4011,N_3597);
nor U5765 (N_5765,N_3678,N_4452);
nor U5766 (N_5766,N_3379,N_4261);
and U5767 (N_5767,N_4086,N_3781);
or U5768 (N_5768,N_4015,N_4102);
and U5769 (N_5769,N_4273,N_3516);
and U5770 (N_5770,N_3834,N_4021);
nor U5771 (N_5771,N_4179,N_3964);
nor U5772 (N_5772,N_3350,N_3638);
nand U5773 (N_5773,N_3609,N_3524);
nor U5774 (N_5774,N_3986,N_3682);
nand U5775 (N_5775,N_3941,N_3322);
nand U5776 (N_5776,N_3922,N_3378);
and U5777 (N_5777,N_4016,N_3402);
nand U5778 (N_5778,N_4172,N_3246);
nand U5779 (N_5779,N_3845,N_3019);
or U5780 (N_5780,N_4437,N_3657);
or U5781 (N_5781,N_3646,N_4020);
or U5782 (N_5782,N_3946,N_3539);
and U5783 (N_5783,N_4144,N_3700);
nor U5784 (N_5784,N_4248,N_3254);
nand U5785 (N_5785,N_4286,N_3458);
and U5786 (N_5786,N_3167,N_4020);
and U5787 (N_5787,N_3546,N_3488);
and U5788 (N_5788,N_4342,N_3234);
nor U5789 (N_5789,N_3324,N_3335);
nand U5790 (N_5790,N_4456,N_4153);
and U5791 (N_5791,N_3751,N_4075);
and U5792 (N_5792,N_3550,N_3785);
or U5793 (N_5793,N_3854,N_4319);
or U5794 (N_5794,N_3381,N_3879);
nand U5795 (N_5795,N_4059,N_3191);
nor U5796 (N_5796,N_4427,N_4138);
and U5797 (N_5797,N_3679,N_3042);
and U5798 (N_5798,N_4011,N_3991);
or U5799 (N_5799,N_3291,N_3382);
nor U5800 (N_5800,N_3706,N_3159);
nor U5801 (N_5801,N_3889,N_4011);
xor U5802 (N_5802,N_4220,N_3329);
nand U5803 (N_5803,N_3053,N_3668);
and U5804 (N_5804,N_4417,N_3226);
nor U5805 (N_5805,N_3216,N_3618);
nand U5806 (N_5806,N_3993,N_3794);
xnor U5807 (N_5807,N_3383,N_3125);
nand U5808 (N_5808,N_4190,N_3727);
and U5809 (N_5809,N_4386,N_3174);
nor U5810 (N_5810,N_3576,N_4051);
nor U5811 (N_5811,N_3470,N_3356);
nand U5812 (N_5812,N_3501,N_4097);
nand U5813 (N_5813,N_3611,N_4107);
and U5814 (N_5814,N_3484,N_3064);
and U5815 (N_5815,N_3947,N_4136);
or U5816 (N_5816,N_3837,N_4192);
nand U5817 (N_5817,N_3973,N_3528);
or U5818 (N_5818,N_4410,N_4274);
or U5819 (N_5819,N_3310,N_3872);
xnor U5820 (N_5820,N_3801,N_4045);
nor U5821 (N_5821,N_4492,N_4036);
nand U5822 (N_5822,N_3907,N_3701);
xnor U5823 (N_5823,N_3092,N_3967);
or U5824 (N_5824,N_3337,N_3445);
or U5825 (N_5825,N_3822,N_4249);
or U5826 (N_5826,N_4119,N_4271);
nand U5827 (N_5827,N_4143,N_4117);
or U5828 (N_5828,N_3641,N_4214);
nor U5829 (N_5829,N_4419,N_3364);
nor U5830 (N_5830,N_3231,N_3374);
nand U5831 (N_5831,N_3543,N_4415);
and U5832 (N_5832,N_3907,N_3236);
or U5833 (N_5833,N_3337,N_3960);
nor U5834 (N_5834,N_3237,N_3714);
or U5835 (N_5835,N_3550,N_3238);
or U5836 (N_5836,N_3608,N_4019);
nand U5837 (N_5837,N_3534,N_4139);
or U5838 (N_5838,N_4325,N_3637);
or U5839 (N_5839,N_3920,N_3213);
or U5840 (N_5840,N_3228,N_4415);
nand U5841 (N_5841,N_4436,N_4382);
or U5842 (N_5842,N_3516,N_3071);
xor U5843 (N_5843,N_3800,N_4370);
or U5844 (N_5844,N_3334,N_3173);
or U5845 (N_5845,N_4424,N_4147);
nand U5846 (N_5846,N_4011,N_3599);
or U5847 (N_5847,N_4480,N_3218);
and U5848 (N_5848,N_3420,N_4222);
nor U5849 (N_5849,N_3182,N_4470);
nand U5850 (N_5850,N_4287,N_4212);
nand U5851 (N_5851,N_3929,N_3258);
nor U5852 (N_5852,N_3663,N_4416);
nand U5853 (N_5853,N_3854,N_3653);
xnor U5854 (N_5854,N_3487,N_3253);
nor U5855 (N_5855,N_4098,N_3093);
or U5856 (N_5856,N_3311,N_3532);
xnor U5857 (N_5857,N_3262,N_3041);
nor U5858 (N_5858,N_4074,N_3332);
and U5859 (N_5859,N_3551,N_3418);
nor U5860 (N_5860,N_3565,N_4348);
or U5861 (N_5861,N_3695,N_3563);
xor U5862 (N_5862,N_3740,N_4221);
nor U5863 (N_5863,N_3077,N_3625);
and U5864 (N_5864,N_4082,N_3336);
and U5865 (N_5865,N_3064,N_3024);
or U5866 (N_5866,N_3588,N_3021);
or U5867 (N_5867,N_3327,N_4203);
or U5868 (N_5868,N_3697,N_4455);
or U5869 (N_5869,N_4361,N_3442);
nand U5870 (N_5870,N_4143,N_4446);
nor U5871 (N_5871,N_4481,N_4112);
and U5872 (N_5872,N_4417,N_3430);
nand U5873 (N_5873,N_4269,N_4111);
nand U5874 (N_5874,N_3624,N_4207);
nor U5875 (N_5875,N_4021,N_3554);
nor U5876 (N_5876,N_3958,N_4376);
or U5877 (N_5877,N_4080,N_3226);
nor U5878 (N_5878,N_3043,N_3449);
nor U5879 (N_5879,N_3942,N_3576);
nor U5880 (N_5880,N_4002,N_3429);
nor U5881 (N_5881,N_3321,N_3842);
nor U5882 (N_5882,N_3212,N_3924);
and U5883 (N_5883,N_4396,N_4286);
nand U5884 (N_5884,N_3546,N_3790);
nor U5885 (N_5885,N_4453,N_3280);
nand U5886 (N_5886,N_4436,N_3943);
nand U5887 (N_5887,N_4407,N_4401);
and U5888 (N_5888,N_3241,N_3326);
nand U5889 (N_5889,N_4445,N_4003);
nand U5890 (N_5890,N_3635,N_4310);
and U5891 (N_5891,N_3365,N_3799);
nor U5892 (N_5892,N_3825,N_4237);
or U5893 (N_5893,N_3050,N_4431);
nor U5894 (N_5894,N_4179,N_4248);
and U5895 (N_5895,N_3202,N_3072);
xnor U5896 (N_5896,N_4245,N_4329);
nand U5897 (N_5897,N_3263,N_3896);
xnor U5898 (N_5898,N_3005,N_3807);
and U5899 (N_5899,N_3136,N_3927);
nand U5900 (N_5900,N_3116,N_4169);
nor U5901 (N_5901,N_3264,N_3223);
nor U5902 (N_5902,N_4341,N_4449);
nand U5903 (N_5903,N_3659,N_3345);
nor U5904 (N_5904,N_3665,N_3977);
xor U5905 (N_5905,N_4068,N_3921);
or U5906 (N_5906,N_4445,N_3659);
nor U5907 (N_5907,N_3856,N_4177);
and U5908 (N_5908,N_3102,N_3770);
and U5909 (N_5909,N_3044,N_4478);
or U5910 (N_5910,N_3438,N_4351);
xor U5911 (N_5911,N_3134,N_4458);
nor U5912 (N_5912,N_4443,N_3399);
nand U5913 (N_5913,N_3655,N_4391);
or U5914 (N_5914,N_3401,N_4396);
nand U5915 (N_5915,N_3510,N_3765);
nor U5916 (N_5916,N_3132,N_3536);
xnor U5917 (N_5917,N_4441,N_4412);
or U5918 (N_5918,N_4134,N_3670);
nor U5919 (N_5919,N_3867,N_3268);
or U5920 (N_5920,N_3312,N_3476);
nor U5921 (N_5921,N_3818,N_3526);
nand U5922 (N_5922,N_4008,N_4248);
nor U5923 (N_5923,N_4036,N_3162);
or U5924 (N_5924,N_4056,N_4003);
and U5925 (N_5925,N_3111,N_3309);
nor U5926 (N_5926,N_4314,N_3111);
nor U5927 (N_5927,N_3480,N_4213);
nand U5928 (N_5928,N_4484,N_3938);
and U5929 (N_5929,N_3060,N_3364);
or U5930 (N_5930,N_4064,N_4075);
or U5931 (N_5931,N_3876,N_3215);
or U5932 (N_5932,N_3653,N_4417);
nor U5933 (N_5933,N_3151,N_4005);
nand U5934 (N_5934,N_4448,N_3225);
nor U5935 (N_5935,N_3065,N_3134);
nand U5936 (N_5936,N_3554,N_4490);
and U5937 (N_5937,N_4149,N_3088);
nand U5938 (N_5938,N_4156,N_3351);
nand U5939 (N_5939,N_3247,N_4482);
or U5940 (N_5940,N_3215,N_3754);
nand U5941 (N_5941,N_4085,N_4249);
and U5942 (N_5942,N_4412,N_4464);
xor U5943 (N_5943,N_4120,N_3864);
nor U5944 (N_5944,N_4287,N_3060);
and U5945 (N_5945,N_4085,N_3599);
or U5946 (N_5946,N_3863,N_3827);
or U5947 (N_5947,N_3661,N_4060);
nor U5948 (N_5948,N_3887,N_3078);
nand U5949 (N_5949,N_3021,N_4356);
or U5950 (N_5950,N_3227,N_4228);
nor U5951 (N_5951,N_4115,N_4192);
or U5952 (N_5952,N_3189,N_3871);
and U5953 (N_5953,N_4448,N_4382);
and U5954 (N_5954,N_4347,N_3626);
xnor U5955 (N_5955,N_3644,N_3436);
or U5956 (N_5956,N_3396,N_3281);
and U5957 (N_5957,N_4386,N_4420);
nand U5958 (N_5958,N_4265,N_3678);
xnor U5959 (N_5959,N_3285,N_3824);
xor U5960 (N_5960,N_3340,N_4122);
or U5961 (N_5961,N_3858,N_4166);
nor U5962 (N_5962,N_3592,N_3977);
or U5963 (N_5963,N_4078,N_3054);
nor U5964 (N_5964,N_3067,N_4345);
nand U5965 (N_5965,N_3825,N_3337);
nand U5966 (N_5966,N_3338,N_4203);
nand U5967 (N_5967,N_3952,N_3557);
or U5968 (N_5968,N_3030,N_3614);
and U5969 (N_5969,N_3110,N_3852);
nand U5970 (N_5970,N_4369,N_4370);
nand U5971 (N_5971,N_4378,N_3062);
xor U5972 (N_5972,N_3021,N_3071);
and U5973 (N_5973,N_4226,N_4233);
or U5974 (N_5974,N_3557,N_3793);
nor U5975 (N_5975,N_3431,N_3488);
xnor U5976 (N_5976,N_3798,N_4281);
xnor U5977 (N_5977,N_3707,N_3169);
or U5978 (N_5978,N_3765,N_4146);
nand U5979 (N_5979,N_4150,N_4308);
nand U5980 (N_5980,N_4051,N_3111);
and U5981 (N_5981,N_4270,N_3834);
nand U5982 (N_5982,N_3508,N_3205);
nand U5983 (N_5983,N_3066,N_4128);
and U5984 (N_5984,N_4004,N_3430);
xor U5985 (N_5985,N_3793,N_4051);
nor U5986 (N_5986,N_3225,N_4429);
and U5987 (N_5987,N_4234,N_3172);
nor U5988 (N_5988,N_3776,N_3617);
nand U5989 (N_5989,N_3985,N_3285);
nor U5990 (N_5990,N_3765,N_4069);
nand U5991 (N_5991,N_3828,N_3684);
or U5992 (N_5992,N_4479,N_3339);
nand U5993 (N_5993,N_4135,N_3044);
or U5994 (N_5994,N_3151,N_4184);
or U5995 (N_5995,N_3169,N_3105);
nand U5996 (N_5996,N_3733,N_3922);
xnor U5997 (N_5997,N_3056,N_3647);
or U5998 (N_5998,N_3144,N_3290);
xnor U5999 (N_5999,N_4226,N_3710);
and U6000 (N_6000,N_4855,N_4862);
or U6001 (N_6001,N_5938,N_4845);
nor U6002 (N_6002,N_5120,N_5882);
or U6003 (N_6003,N_4658,N_5198);
nor U6004 (N_6004,N_5878,N_4939);
or U6005 (N_6005,N_5418,N_4560);
xnor U6006 (N_6006,N_5399,N_5038);
nand U6007 (N_6007,N_4955,N_5027);
and U6008 (N_6008,N_4577,N_5694);
and U6009 (N_6009,N_4891,N_5477);
and U6010 (N_6010,N_4950,N_4598);
and U6011 (N_6011,N_5787,N_5087);
xor U6012 (N_6012,N_5309,N_4595);
nor U6013 (N_6013,N_4974,N_5398);
and U6014 (N_6014,N_5638,N_5282);
xor U6015 (N_6015,N_4832,N_4758);
nor U6016 (N_6016,N_4791,N_4659);
nand U6017 (N_6017,N_5154,N_4611);
or U6018 (N_6018,N_5011,N_4669);
nand U6019 (N_6019,N_5425,N_5849);
nand U6020 (N_6020,N_4581,N_4857);
nor U6021 (N_6021,N_4667,N_5046);
or U6022 (N_6022,N_4701,N_4705);
nand U6023 (N_6023,N_4930,N_5953);
or U6024 (N_6024,N_4784,N_5085);
nor U6025 (N_6025,N_4524,N_5862);
nor U6026 (N_6026,N_5419,N_4601);
or U6027 (N_6027,N_4990,N_5677);
nor U6028 (N_6028,N_4580,N_5002);
xnor U6029 (N_6029,N_5243,N_5816);
and U6030 (N_6030,N_4660,N_4689);
nand U6031 (N_6031,N_5393,N_4633);
nor U6032 (N_6032,N_5003,N_5904);
and U6033 (N_6033,N_4706,N_4536);
nor U6034 (N_6034,N_5396,N_4762);
xor U6035 (N_6035,N_4926,N_5760);
and U6036 (N_6036,N_5640,N_5054);
nor U6037 (N_6037,N_4795,N_5505);
or U6038 (N_6038,N_4743,N_4788);
nand U6039 (N_6039,N_5860,N_4715);
or U6040 (N_6040,N_5701,N_4892);
xor U6041 (N_6041,N_5102,N_4613);
nand U6042 (N_6042,N_5471,N_5684);
and U6043 (N_6043,N_5139,N_4878);
nand U6044 (N_6044,N_4693,N_5337);
nor U6045 (N_6045,N_4526,N_5680);
or U6046 (N_6046,N_4945,N_4516);
and U6047 (N_6047,N_4702,N_5806);
nor U6048 (N_6048,N_5109,N_5014);
or U6049 (N_6049,N_5976,N_5526);
xor U6050 (N_6050,N_5698,N_5813);
or U6051 (N_6051,N_5015,N_4805);
nor U6052 (N_6052,N_5788,N_5898);
nand U6053 (N_6053,N_5868,N_5746);
nor U6054 (N_6054,N_4563,N_5415);
xor U6055 (N_6055,N_5402,N_4834);
nor U6056 (N_6056,N_5847,N_4948);
nand U6057 (N_6057,N_5101,N_5263);
or U6058 (N_6058,N_4671,N_4681);
nor U6059 (N_6059,N_5594,N_4804);
or U6060 (N_6060,N_5836,N_4809);
nand U6061 (N_6061,N_5707,N_5215);
or U6062 (N_6062,N_5678,N_4638);
nand U6063 (N_6063,N_5919,N_5785);
or U6064 (N_6064,N_5357,N_5962);
nand U6065 (N_6065,N_5855,N_4906);
xnor U6066 (N_6066,N_5628,N_4854);
nand U6067 (N_6067,N_4873,N_5850);
or U6068 (N_6068,N_5254,N_5292);
nor U6069 (N_6069,N_5016,N_5531);
or U6070 (N_6070,N_5539,N_5278);
nand U6071 (N_6071,N_5079,N_5876);
nor U6072 (N_6072,N_5358,N_4925);
and U6073 (N_6073,N_5774,N_5761);
nand U6074 (N_6074,N_5590,N_5567);
or U6075 (N_6075,N_4707,N_5366);
or U6076 (N_6076,N_5853,N_5889);
nand U6077 (N_6077,N_5173,N_5652);
nand U6078 (N_6078,N_5975,N_5161);
nor U6079 (N_6079,N_4952,N_5744);
and U6080 (N_6080,N_5752,N_5374);
or U6081 (N_6081,N_4896,N_5729);
or U6082 (N_6082,N_4986,N_5851);
nor U6083 (N_6083,N_5627,N_5621);
nor U6084 (N_6084,N_5513,N_5560);
nand U6085 (N_6085,N_4650,N_4898);
nand U6086 (N_6086,N_5148,N_5696);
and U6087 (N_6087,N_5410,N_5714);
and U6088 (N_6088,N_5424,N_5227);
nor U6089 (N_6089,N_5685,N_4709);
nand U6090 (N_6090,N_5940,N_5755);
or U6091 (N_6091,N_4760,N_4517);
or U6092 (N_6092,N_5636,N_5769);
nor U6093 (N_6093,N_4901,N_5069);
or U6094 (N_6094,N_4724,N_5792);
nand U6095 (N_6095,N_5327,N_5197);
nand U6096 (N_6096,N_5965,N_5454);
nand U6097 (N_6097,N_5821,N_5075);
nand U6098 (N_6098,N_5153,N_5713);
nor U6099 (N_6099,N_5405,N_5974);
and U6100 (N_6100,N_5112,N_5029);
nand U6101 (N_6101,N_5558,N_5190);
xor U6102 (N_6102,N_5020,N_4818);
nor U6103 (N_6103,N_4992,N_5325);
nand U6104 (N_6104,N_5599,N_5146);
nor U6105 (N_6105,N_5651,N_4645);
nor U6106 (N_6106,N_5500,N_5004);
or U6107 (N_6107,N_5935,N_5013);
nand U6108 (N_6108,N_5482,N_5320);
and U6109 (N_6109,N_4867,N_4769);
nand U6110 (N_6110,N_5926,N_4940);
nor U6111 (N_6111,N_4782,N_4923);
and U6112 (N_6112,N_5529,N_4808);
and U6113 (N_6113,N_5068,N_5213);
nand U6114 (N_6114,N_5209,N_4648);
nor U6115 (N_6115,N_5059,N_5747);
nand U6116 (N_6116,N_5416,N_5492);
nor U6117 (N_6117,N_5629,N_4604);
or U6118 (N_6118,N_4876,N_5283);
nor U6119 (N_6119,N_5447,N_5715);
or U6120 (N_6120,N_4778,N_4897);
or U6121 (N_6121,N_5194,N_5000);
and U6122 (N_6122,N_5913,N_5247);
or U6123 (N_6123,N_4872,N_5439);
nand U6124 (N_6124,N_4972,N_5909);
nor U6125 (N_6125,N_5830,N_4583);
nor U6126 (N_6126,N_5995,N_5165);
nor U6127 (N_6127,N_5386,N_5201);
nor U6128 (N_6128,N_5668,N_4713);
xor U6129 (N_6129,N_5519,N_5767);
nor U6130 (N_6130,N_4614,N_4728);
nor U6131 (N_6131,N_5289,N_4554);
and U6132 (N_6132,N_5892,N_5181);
and U6133 (N_6133,N_5056,N_5506);
nand U6134 (N_6134,N_5080,N_5572);
nor U6135 (N_6135,N_5062,N_5196);
and U6136 (N_6136,N_5954,N_5097);
nand U6137 (N_6137,N_5809,N_5508);
nor U6138 (N_6138,N_5899,N_4840);
nor U6139 (N_6139,N_5566,N_4970);
nor U6140 (N_6140,N_5268,N_4550);
or U6141 (N_6141,N_4936,N_4523);
and U6142 (N_6142,N_5269,N_5286);
nand U6143 (N_6143,N_5642,N_4775);
nor U6144 (N_6144,N_4703,N_4932);
and U6145 (N_6145,N_5711,N_5001);
nor U6146 (N_6146,N_5193,N_4785);
nor U6147 (N_6147,N_5491,N_4924);
nand U6148 (N_6148,N_5695,N_4719);
or U6149 (N_6149,N_5923,N_4666);
nand U6150 (N_6150,N_5228,N_5671);
nand U6151 (N_6151,N_4831,N_4911);
nand U6152 (N_6152,N_4734,N_4989);
xor U6153 (N_6153,N_5277,N_4838);
nor U6154 (N_6154,N_4649,N_4875);
nand U6155 (N_6155,N_5478,N_4879);
and U6156 (N_6156,N_4670,N_5351);
nand U6157 (N_6157,N_4531,N_5987);
or U6158 (N_6158,N_5406,N_5992);
nand U6159 (N_6159,N_5687,N_5972);
and U6160 (N_6160,N_5635,N_5782);
xnor U6161 (N_6161,N_5431,N_5328);
xor U6162 (N_6162,N_4973,N_5552);
nand U6163 (N_6163,N_5933,N_4912);
xnor U6164 (N_6164,N_4625,N_4616);
xnor U6165 (N_6165,N_5622,N_5149);
nor U6166 (N_6166,N_5615,N_4542);
or U6167 (N_6167,N_5261,N_5632);
xor U6168 (N_6168,N_5208,N_5455);
nand U6169 (N_6169,N_4700,N_5699);
nor U6170 (N_6170,N_5423,N_4889);
or U6171 (N_6171,N_5249,N_5412);
nor U6172 (N_6172,N_4870,N_4815);
xor U6173 (N_6173,N_5749,N_5129);
and U6174 (N_6174,N_5742,N_5185);
and U6175 (N_6175,N_5570,N_4914);
and U6176 (N_6176,N_4535,N_4573);
nor U6177 (N_6177,N_4880,N_5989);
nor U6178 (N_6178,N_4806,N_5260);
xnor U6179 (N_6179,N_4732,N_4800);
nor U6180 (N_6180,N_5061,N_5817);
nand U6181 (N_6181,N_5661,N_5693);
or U6182 (N_6182,N_5872,N_4835);
and U6183 (N_6183,N_5676,N_4518);
and U6184 (N_6184,N_4929,N_5446);
nor U6185 (N_6185,N_5319,N_5907);
nand U6186 (N_6186,N_5221,N_5238);
or U6187 (N_6187,N_5559,N_4773);
nor U6188 (N_6188,N_4755,N_5473);
nor U6189 (N_6189,N_5229,N_5818);
or U6190 (N_6190,N_4810,N_5956);
nor U6191 (N_6191,N_5379,N_5512);
or U6192 (N_6192,N_4506,N_5541);
nor U6193 (N_6193,N_5662,N_5440);
nor U6194 (N_6194,N_5470,N_4890);
nand U6195 (N_6195,N_4748,N_5771);
nor U6196 (N_6196,N_5138,N_5382);
or U6197 (N_6197,N_4764,N_4586);
nor U6198 (N_6198,N_4844,N_5515);
nand U6199 (N_6199,N_4640,N_5784);
nor U6200 (N_6200,N_5397,N_4786);
nand U6201 (N_6201,N_5312,N_4623);
nand U6202 (N_6202,N_5563,N_5609);
or U6203 (N_6203,N_5799,N_5834);
nor U6204 (N_6204,N_5308,N_4942);
nand U6205 (N_6205,N_5066,N_5646);
and U6206 (N_6206,N_4672,N_4678);
nor U6207 (N_6207,N_5144,N_5712);
nor U6208 (N_6208,N_5468,N_5321);
nand U6209 (N_6209,N_4673,N_4803);
or U6210 (N_6210,N_5955,N_5465);
nand U6211 (N_6211,N_4657,N_4979);
xnor U6212 (N_6212,N_5795,N_4982);
and U6213 (N_6213,N_5996,N_4736);
or U6214 (N_6214,N_4731,N_4829);
xnor U6215 (N_6215,N_5305,N_4602);
and U6216 (N_6216,N_4621,N_5307);
or U6217 (N_6217,N_5039,N_5207);
nor U6218 (N_6218,N_4908,N_4720);
nand U6219 (N_6219,N_5272,N_4918);
nand U6220 (N_6220,N_5350,N_5338);
and U6221 (N_6221,N_5751,N_4859);
nor U6222 (N_6222,N_4874,N_4722);
xnor U6223 (N_6223,N_5302,N_5259);
nand U6224 (N_6224,N_5130,N_4994);
and U6225 (N_6225,N_4528,N_5532);
nand U6226 (N_6226,N_5579,N_4742);
and U6227 (N_6227,N_5819,N_5918);
or U6228 (N_6228,N_5377,N_5951);
nor U6229 (N_6229,N_5533,N_5610);
and U6230 (N_6230,N_4676,N_5511);
nor U6231 (N_6231,N_5562,N_5945);
nor U6232 (N_6232,N_5331,N_4564);
or U6233 (N_6233,N_5043,N_5219);
nor U6234 (N_6234,N_5591,N_4863);
nand U6235 (N_6235,N_5256,N_5490);
nand U6236 (N_6236,N_5091,N_5762);
or U6237 (N_6237,N_5902,N_5815);
and U6238 (N_6238,N_4916,N_5537);
nor U6239 (N_6239,N_4981,N_5811);
or U6240 (N_6240,N_5116,N_4813);
and U6241 (N_6241,N_5222,N_4587);
nand U6242 (N_6242,N_5401,N_4954);
and U6243 (N_6243,N_5450,N_5518);
nor U6244 (N_6244,N_4735,N_5527);
and U6245 (N_6245,N_5077,N_4740);
nand U6246 (N_6246,N_5589,N_5502);
nand U6247 (N_6247,N_4774,N_4591);
and U6248 (N_6248,N_4675,N_5369);
nand U6249 (N_6249,N_5287,N_5117);
nand U6250 (N_6250,N_5791,N_4860);
nand U6251 (N_6251,N_5820,N_5607);
xnor U6252 (N_6252,N_5352,N_5666);
and U6253 (N_6253,N_5187,N_5800);
or U6254 (N_6254,N_5757,N_5373);
or U6255 (N_6255,N_5253,N_5794);
or U6256 (N_6256,N_5070,N_5167);
and U6257 (N_6257,N_4971,N_4605);
or U6258 (N_6258,N_4522,N_5394);
nand U6259 (N_6259,N_4861,N_5550);
nand U6260 (N_6260,N_5275,N_5252);
xnor U6261 (N_6261,N_5353,N_5499);
nand U6262 (N_6262,N_5279,N_5223);
nand U6263 (N_6263,N_4894,N_5875);
nor U6264 (N_6264,N_5006,N_4883);
and U6265 (N_6265,N_5643,N_5304);
or U6266 (N_6266,N_4593,N_4600);
nor U6267 (N_6267,N_5485,N_5999);
or U6268 (N_6268,N_5801,N_4824);
xnor U6269 (N_6269,N_4776,N_5530);
and U6270 (N_6270,N_5990,N_4631);
nor U6271 (N_6271,N_5957,N_5549);
xnor U6272 (N_6272,N_4946,N_5498);
xnor U6273 (N_6273,N_5143,N_5157);
or U6274 (N_6274,N_4569,N_5180);
or U6275 (N_6275,N_5895,N_5597);
or U6276 (N_6276,N_5191,N_5125);
xor U6277 (N_6277,N_5690,N_5780);
nor U6278 (N_6278,N_5947,N_5561);
nor U6279 (N_6279,N_5808,N_4744);
or U6280 (N_6280,N_4910,N_5964);
nor U6281 (N_6281,N_4796,N_5072);
nand U6282 (N_6282,N_4960,N_4754);
nor U6283 (N_6283,N_4933,N_5152);
nor U6284 (N_6284,N_5585,N_5348);
or U6285 (N_6285,N_5950,N_4884);
and U6286 (N_6286,N_5035,N_5104);
xnor U6287 (N_6287,N_4823,N_5534);
nand U6288 (N_6288,N_4641,N_5683);
or U6289 (N_6289,N_5248,N_5958);
or U6290 (N_6290,N_5928,N_5578);
nand U6291 (N_6291,N_5576,N_5472);
nor U6292 (N_6292,N_4541,N_5970);
nor U6293 (N_6293,N_5121,N_5119);
nor U6294 (N_6294,N_5639,N_4661);
nor U6295 (N_6295,N_5914,N_4651);
or U6296 (N_6296,N_5298,N_5391);
nand U6297 (N_6297,N_5442,N_4966);
or U6298 (N_6298,N_5865,N_5370);
and U6299 (N_6299,N_5433,N_5335);
xor U6300 (N_6300,N_5720,N_5825);
and U6301 (N_6301,N_5390,N_5984);
nand U6302 (N_6302,N_4726,N_5625);
nand U6303 (N_6303,N_5368,N_5520);
or U6304 (N_6304,N_5235,N_4557);
and U6305 (N_6305,N_5839,N_4699);
nor U6306 (N_6306,N_4751,N_5569);
nor U6307 (N_6307,N_5702,N_5978);
nor U6308 (N_6308,N_5703,N_4548);
xnor U6309 (N_6309,N_5007,N_4729);
nor U6310 (N_6310,N_5900,N_5326);
nor U6311 (N_6311,N_4770,N_5600);
nand U6312 (N_6312,N_5837,N_4698);
and U6313 (N_6313,N_5034,N_4768);
or U6314 (N_6314,N_4747,N_5944);
and U6315 (N_6315,N_5967,N_5294);
or U6316 (N_6316,N_4652,N_4919);
xor U6317 (N_6317,N_5092,N_5731);
or U6318 (N_6318,N_4852,N_4525);
nor U6319 (N_6319,N_4686,N_4576);
nor U6320 (N_6320,N_5008,N_5267);
xor U6321 (N_6321,N_5665,N_4882);
xor U6322 (N_6322,N_5961,N_5067);
nor U6323 (N_6323,N_5859,N_4963);
and U6324 (N_6324,N_5555,N_4642);
xnor U6325 (N_6325,N_5057,N_5115);
nand U6326 (N_6326,N_4841,N_5732);
nand U6327 (N_6327,N_4688,N_5886);
nand U6328 (N_6328,N_5280,N_4997);
xor U6329 (N_6329,N_4630,N_5789);
or U6330 (N_6330,N_5748,N_5186);
nand U6331 (N_6331,N_5841,N_5273);
and U6332 (N_6332,N_5224,N_4510);
and U6333 (N_6333,N_5735,N_5218);
nand U6334 (N_6334,N_5573,N_4848);
nand U6335 (N_6335,N_4802,N_5188);
or U6336 (N_6336,N_5618,N_5340);
nor U6337 (N_6337,N_4561,N_5740);
nor U6338 (N_6338,N_4811,N_5291);
or U6339 (N_6339,N_5064,N_4655);
and U6340 (N_6340,N_5400,N_5910);
nand U6341 (N_6341,N_5613,N_4512);
or U6342 (N_6342,N_5241,N_5611);
or U6343 (N_6343,N_5546,N_5420);
nor U6344 (N_6344,N_5796,N_4664);
and U6345 (N_6345,N_5237,N_5088);
and U6346 (N_6346,N_5941,N_5032);
or U6347 (N_6347,N_5018,N_5495);
nand U6348 (N_6348,N_5060,N_5045);
or U6349 (N_6349,N_5606,N_5971);
nor U6350 (N_6350,N_5959,N_5612);
xnor U6351 (N_6351,N_5347,N_4567);
and U6352 (N_6352,N_5790,N_4738);
nand U6353 (N_6353,N_4509,N_4812);
nand U6354 (N_6354,N_4837,N_4527);
and U6355 (N_6355,N_5988,N_5462);
and U6356 (N_6356,N_5336,N_5486);
or U6357 (N_6357,N_5575,N_4961);
or U6358 (N_6358,N_4606,N_4827);
nand U6359 (N_6359,N_5783,N_5881);
nor U6360 (N_6360,N_4777,N_4987);
nor U6361 (N_6361,N_5041,N_5344);
nor U6362 (N_6362,N_5009,N_5436);
nand U6363 (N_6363,N_5290,N_5487);
nand U6364 (N_6364,N_4714,N_5040);
nor U6365 (N_6365,N_5132,N_5604);
or U6366 (N_6366,N_5324,N_5083);
xnor U6367 (N_6367,N_5966,N_4568);
nand U6368 (N_6368,N_4749,N_5301);
and U6369 (N_6369,N_4644,N_5276);
or U6370 (N_6370,N_5176,N_4781);
and U6371 (N_6371,N_5538,N_4597);
nand U6372 (N_6372,N_5557,N_4656);
nand U6373 (N_6373,N_5897,N_5133);
nor U6374 (N_6374,N_4502,N_5262);
or U6375 (N_6375,N_5548,N_5633);
and U6376 (N_6376,N_4530,N_5584);
and U6377 (N_6377,N_5669,N_5595);
nor U6378 (N_6378,N_4763,N_5588);
xnor U6379 (N_6379,N_4765,N_5673);
xor U6380 (N_6380,N_4575,N_5392);
and U6381 (N_6381,N_4725,N_4902);
and U6382 (N_6382,N_4552,N_4716);
nor U6383 (N_6383,N_4967,N_5395);
nand U6384 (N_6384,N_5051,N_4787);
nor U6385 (N_6385,N_5883,N_4622);
and U6386 (N_6386,N_5688,N_5058);
and U6387 (N_6387,N_5773,N_5619);
nor U6388 (N_6388,N_4615,N_5764);
nor U6389 (N_6389,N_5217,N_4682);
nor U6390 (N_6390,N_4962,N_5587);
or U6391 (N_6391,N_5159,N_5106);
or U6392 (N_6392,N_4501,N_4694);
and U6393 (N_6393,N_5124,N_5998);
nor U6394 (N_6394,N_5509,N_5355);
nand U6395 (N_6395,N_5689,N_4637);
xnor U6396 (N_6396,N_5758,N_5725);
or U6397 (N_6397,N_4904,N_4964);
nand U6398 (N_6398,N_5936,N_5494);
or U6399 (N_6399,N_5310,N_5441);
or U6400 (N_6400,N_5210,N_5281);
and U6401 (N_6401,N_4627,N_4584);
or U6402 (N_6402,N_4980,N_5778);
nand U6403 (N_6403,N_5943,N_5905);
xor U6404 (N_6404,N_5536,N_5543);
and U6405 (N_6405,N_5963,N_5380);
nor U6406 (N_6406,N_5523,N_4590);
and U6407 (N_6407,N_4572,N_5111);
nand U6408 (N_6408,N_4558,N_5997);
and U6409 (N_6409,N_5048,N_4909);
or U6410 (N_6410,N_5503,N_4723);
nand U6411 (N_6411,N_4692,N_5723);
and U6412 (N_6412,N_5031,N_5081);
and U6413 (N_6413,N_5036,N_5522);
nand U6414 (N_6414,N_4935,N_5983);
and U6415 (N_6415,N_4985,N_4816);
and U6416 (N_6416,N_5750,N_5717);
and U6417 (N_6417,N_5623,N_5657);
or U6418 (N_6418,N_5314,N_4999);
nand U6419 (N_6419,N_5202,N_5843);
and U6420 (N_6420,N_5738,N_5903);
or U6421 (N_6421,N_5094,N_5655);
nor U6422 (N_6422,N_5867,N_5356);
or U6423 (N_6423,N_4520,N_4500);
nor U6424 (N_6424,N_4543,N_4968);
and U6425 (N_6425,N_5183,N_5244);
nor U6426 (N_6426,N_5074,N_5797);
nand U6427 (N_6427,N_5164,N_5147);
and U6428 (N_6428,N_5318,N_5675);
or U6429 (N_6429,N_5343,N_5220);
or U6430 (N_6430,N_5274,N_4565);
nand U6431 (N_6431,N_4913,N_5387);
nand U6432 (N_6432,N_4757,N_5814);
and U6433 (N_6433,N_4790,N_5718);
and U6434 (N_6434,N_5616,N_4507);
xnor U6435 (N_6435,N_5832,N_4534);
xnor U6436 (N_6436,N_4938,N_4846);
and U6437 (N_6437,N_5672,N_5826);
or U6438 (N_6438,N_4739,N_4975);
nand U6439 (N_6439,N_5551,N_5017);
or U6440 (N_6440,N_5894,N_5982);
nand U6441 (N_6441,N_5427,N_5199);
and U6442 (N_6442,N_4574,N_4941);
or U6443 (N_6443,N_4881,N_4976);
nand U6444 (N_6444,N_5756,N_5448);
xnor U6445 (N_6445,N_5245,N_5359);
nor U6446 (N_6446,N_5545,N_5216);
xor U6447 (N_6447,N_5367,N_5103);
nand U6448 (N_6448,N_4792,N_4922);
nand U6449 (N_6449,N_5136,N_5802);
nand U6450 (N_6450,N_5838,N_5175);
and U6451 (N_6451,N_5047,N_4856);
nor U6452 (N_6452,N_5901,N_4599);
nor U6453 (N_6453,N_4610,N_5844);
or U6454 (N_6454,N_5554,N_5630);
nand U6455 (N_6455,N_4514,N_5388);
nand U6456 (N_6456,N_4920,N_4704);
or U6457 (N_6457,N_5107,N_4690);
or U6458 (N_6458,N_5288,N_4585);
nand U6459 (N_6459,N_4907,N_5805);
nor U6460 (N_6460,N_5601,N_5948);
and U6461 (N_6461,N_5848,N_5428);
nor U6462 (N_6462,N_5863,N_5650);
nor U6463 (N_6463,N_5052,N_5484);
and U6464 (N_6464,N_5179,N_4545);
nand U6465 (N_6465,N_5925,N_5877);
nand U6466 (N_6466,N_5389,N_5251);
or U6467 (N_6467,N_4727,N_5409);
nand U6468 (N_6468,N_4903,N_4866);
nor U6469 (N_6469,N_4825,N_5917);
and U6470 (N_6470,N_5127,N_4915);
or U6471 (N_6471,N_5524,N_4503);
or U6472 (N_6472,N_4836,N_4579);
or U6473 (N_6473,N_5177,N_5915);
nand U6474 (N_6474,N_5890,N_4839);
or U6475 (N_6475,N_4708,N_5775);
and U6476 (N_6476,N_5211,N_5323);
and U6477 (N_6477,N_4820,N_5417);
nor U6478 (N_6478,N_4830,N_5765);
nand U6479 (N_6479,N_4959,N_5602);
nand U6480 (N_6480,N_5023,N_5645);
nand U6481 (N_6481,N_5189,N_5766);
nand U6482 (N_6482,N_5170,N_5076);
or U6483 (N_6483,N_5030,N_4793);
or U6484 (N_6484,N_4944,N_4588);
and U6485 (N_6485,N_4737,N_5535);
and U6486 (N_6486,N_4592,N_4877);
xnor U6487 (N_6487,N_4869,N_5354);
nand U6488 (N_6488,N_5908,N_5073);
nand U6489 (N_6489,N_4871,N_4799);
or U6490 (N_6490,N_5285,N_5239);
nand U6491 (N_6491,N_5481,N_5710);
or U6492 (N_6492,N_5376,N_5322);
nor U6493 (N_6493,N_4521,N_5654);
nor U6494 (N_6494,N_5828,N_5293);
nor U6495 (N_6495,N_5582,N_4556);
and U6496 (N_6496,N_5303,N_4993);
and U6497 (N_6497,N_4928,N_4680);
nand U6498 (N_6498,N_5497,N_5295);
nand U6499 (N_6499,N_5994,N_5706);
nor U6500 (N_6500,N_5174,N_5206);
nor U6501 (N_6501,N_5037,N_5663);
nor U6502 (N_6502,N_5822,N_4629);
or U6503 (N_6503,N_5460,N_5184);
or U6504 (N_6504,N_4547,N_5553);
nor U6505 (N_6505,N_4780,N_5577);
nor U6506 (N_6506,N_4632,N_4783);
nor U6507 (N_6507,N_5242,N_4998);
nand U6508 (N_6508,N_4772,N_4977);
nor U6509 (N_6509,N_5580,N_5300);
or U6510 (N_6510,N_5445,N_4582);
nand U6511 (N_6511,N_5949,N_4771);
and U6512 (N_6512,N_5985,N_5960);
or U6513 (N_6513,N_5339,N_5649);
and U6514 (N_6514,N_4549,N_5055);
nor U6515 (N_6515,N_5150,N_4538);
or U6516 (N_6516,N_5719,N_4895);
nor U6517 (N_6517,N_4504,N_4662);
nand U6518 (N_6518,N_5574,N_4899);
or U6519 (N_6519,N_5044,N_5873);
nor U6520 (N_6520,N_5459,N_5306);
nand U6521 (N_6521,N_5979,N_5807);
and U6522 (N_6522,N_5686,N_4596);
or U6523 (N_6523,N_5861,N_4821);
nand U6524 (N_6524,N_5086,N_5476);
or U6525 (N_6525,N_4798,N_5605);
nand U6526 (N_6526,N_5258,N_5246);
and U6527 (N_6527,N_5099,N_5010);
and U6528 (N_6528,N_5362,N_5082);
or U6529 (N_6529,N_5458,N_5980);
nand U6530 (N_6530,N_5065,N_4733);
nor U6531 (N_6531,N_5469,N_5641);
xnor U6532 (N_6532,N_5781,N_5846);
or U6533 (N_6533,N_5722,N_4620);
or U6534 (N_6534,N_5516,N_5842);
and U6535 (N_6535,N_4628,N_4851);
and U6536 (N_6536,N_5297,N_5528);
nor U6537 (N_6537,N_5346,N_5544);
xnor U6538 (N_6538,N_4607,N_5042);
nand U6539 (N_6539,N_5608,N_4779);
xor U6540 (N_6540,N_5168,N_4537);
and U6541 (N_6541,N_4544,N_4794);
nand U6542 (N_6542,N_5525,N_5946);
xor U6543 (N_6543,N_4943,N_4636);
or U6544 (N_6544,N_4647,N_4646);
nor U6545 (N_6545,N_5429,N_5345);
or U6546 (N_6546,N_5110,N_5810);
or U6547 (N_6547,N_4814,N_4745);
or U6548 (N_6548,N_5916,N_5697);
nand U6549 (N_6549,N_5866,N_4654);
or U6550 (N_6550,N_4965,N_4949);
and U6551 (N_6551,N_5835,N_4893);
and U6552 (N_6552,N_5063,N_5571);
and U6553 (N_6553,N_5141,N_4511);
or U6554 (N_6554,N_5178,N_4712);
or U6555 (N_6555,N_5583,N_4589);
or U6556 (N_6556,N_4957,N_4842);
and U6557 (N_6557,N_5664,N_4515);
nand U6558 (N_6558,N_5005,N_5736);
xor U6559 (N_6559,N_5977,N_5426);
or U6560 (N_6560,N_4562,N_4766);
nor U6561 (N_6561,N_5874,N_5421);
nor U6562 (N_6562,N_5973,N_4519);
nand U6563 (N_6563,N_5856,N_4753);
xnor U6564 (N_6564,N_5026,N_4691);
and U6565 (N_6565,N_5365,N_5586);
nor U6566 (N_6566,N_4991,N_5670);
nor U6567 (N_6567,N_5430,N_4619);
and U6568 (N_6568,N_4505,N_5659);
and U6569 (N_6569,N_5050,N_5078);
and U6570 (N_6570,N_5404,N_4931);
and U6571 (N_6571,N_5869,N_5403);
or U6572 (N_6572,N_4789,N_4746);
nand U6573 (N_6573,N_4847,N_5644);
nand U6574 (N_6574,N_5793,N_5432);
xor U6575 (N_6575,N_4653,N_5656);
xnor U6576 (N_6576,N_5829,N_5371);
nor U6577 (N_6577,N_5931,N_4626);
xnor U6578 (N_6578,N_5169,N_4665);
nor U6579 (N_6579,N_4730,N_5614);
or U6580 (N_6580,N_5479,N_5200);
or U6581 (N_6581,N_4634,N_5496);
nand U6582 (N_6582,N_4969,N_4546);
and U6583 (N_6583,N_5240,N_5071);
nor U6584 (N_6584,N_5547,N_5438);
nand U6585 (N_6585,N_5381,N_5777);
nand U6586 (N_6586,N_5924,N_5932);
or U6587 (N_6587,N_5507,N_4674);
xor U6588 (N_6588,N_5332,N_5705);
nand U6589 (N_6589,N_5726,N_5451);
and U6590 (N_6590,N_5233,N_5691);
or U6591 (N_6591,N_4684,N_5679);
nor U6592 (N_6592,N_4677,N_5313);
or U6593 (N_6593,N_4868,N_5823);
or U6594 (N_6594,N_5375,N_4983);
nand U6595 (N_6595,N_5779,N_4687);
and U6596 (N_6596,N_5135,N_5271);
and U6597 (N_6597,N_5753,N_5893);
nor U6598 (N_6598,N_4513,N_5739);
nor U6599 (N_6599,N_5768,N_5192);
or U6600 (N_6600,N_5708,N_5212);
xnor U6601 (N_6601,N_5372,N_5596);
or U6602 (N_6602,N_4921,N_5880);
and U6603 (N_6603,N_4752,N_4609);
nor U6604 (N_6604,N_5896,N_5033);
nand U6605 (N_6605,N_5105,N_4721);
and U6606 (N_6606,N_5151,N_5879);
or U6607 (N_6607,N_5284,N_5226);
or U6608 (N_6608,N_5108,N_5021);
and U6609 (N_6609,N_4819,N_4508);
xor U6610 (N_6610,N_4618,N_5857);
or U6611 (N_6611,N_4612,N_4885);
nand U6612 (N_6612,N_5126,N_5493);
and U6613 (N_6613,N_5854,N_5232);
nand U6614 (N_6614,N_5122,N_5234);
nand U6615 (N_6615,N_5884,N_4988);
xnor U6616 (N_6616,N_5329,N_4635);
or U6617 (N_6617,N_5840,N_4807);
or U6618 (N_6618,N_5598,N_4683);
xor U6619 (N_6619,N_5763,N_5142);
nor U6620 (N_6620,N_5422,N_5700);
and U6621 (N_6621,N_4828,N_5028);
and U6622 (N_6622,N_5911,N_5437);
nand U6623 (N_6623,N_5991,N_5203);
nor U6624 (N_6624,N_5123,N_5333);
or U6625 (N_6625,N_4533,N_5658);
nand U6626 (N_6626,N_5255,N_5467);
nor U6627 (N_6627,N_5118,N_5349);
and U6628 (N_6628,N_5128,N_5934);
nand U6629 (N_6629,N_5134,N_5231);
or U6630 (N_6630,N_5025,N_4958);
nand U6631 (N_6631,N_4937,N_5114);
nand U6632 (N_6632,N_5089,N_5137);
nor U6633 (N_6633,N_5734,N_4858);
nor U6634 (N_6634,N_5162,N_5759);
or U6635 (N_6635,N_5682,N_5824);
nor U6636 (N_6636,N_4559,N_5969);
or U6637 (N_6637,N_5986,N_5317);
nand U6638 (N_6638,N_4643,N_5592);
nor U6639 (N_6639,N_5564,N_4532);
nor U6640 (N_6640,N_5937,N_5411);
nor U6641 (N_6641,N_4826,N_5160);
and U6642 (N_6642,N_5885,N_5163);
or U6643 (N_6643,N_5444,N_5870);
and U6644 (N_6644,N_4617,N_5704);
or U6645 (N_6645,N_5648,N_4953);
or U6646 (N_6646,N_5634,N_4797);
nand U6647 (N_6647,N_4540,N_5090);
nand U6648 (N_6648,N_4529,N_5993);
nand U6649 (N_6649,N_5456,N_5012);
nand U6650 (N_6650,N_4553,N_4603);
or U6651 (N_6651,N_5334,N_5770);
xor U6652 (N_6652,N_4718,N_4956);
nand U6653 (N_6653,N_4822,N_5929);
nor U6654 (N_6654,N_5754,N_5360);
nand U6655 (N_6655,N_5724,N_5236);
or U6656 (N_6656,N_5413,N_5158);
nand U6657 (N_6657,N_5653,N_5435);
nand U6658 (N_6658,N_5205,N_5449);
nand U6659 (N_6659,N_5385,N_5912);
or U6660 (N_6660,N_5145,N_5831);
nand U6661 (N_6661,N_5716,N_5674);
or U6662 (N_6662,N_5786,N_5316);
or U6663 (N_6663,N_4539,N_4696);
nand U6664 (N_6664,N_5845,N_5593);
xor U6665 (N_6665,N_5019,N_5510);
nand U6666 (N_6666,N_5521,N_4767);
nor U6667 (N_6667,N_5084,N_5833);
nand U6668 (N_6668,N_4984,N_4668);
nor U6669 (N_6669,N_5155,N_5093);
nor U6670 (N_6670,N_4947,N_5342);
or U6671 (N_6671,N_5637,N_5501);
or U6672 (N_6672,N_4717,N_5647);
nor U6673 (N_6673,N_5930,N_5457);
nand U6674 (N_6674,N_4817,N_5542);
nand U6675 (N_6675,N_5384,N_5743);
or U6676 (N_6676,N_4570,N_4849);
and U6677 (N_6677,N_5888,N_5182);
or U6678 (N_6678,N_5053,N_5266);
xnor U6679 (N_6679,N_5741,N_5363);
nand U6680 (N_6680,N_5812,N_5581);
or U6681 (N_6681,N_5730,N_5968);
and U6682 (N_6682,N_5172,N_4917);
nor U6683 (N_6683,N_5772,N_5939);
nor U6684 (N_6684,N_5852,N_5667);
and U6685 (N_6685,N_5981,N_5452);
nor U6686 (N_6686,N_5483,N_5942);
nand U6687 (N_6687,N_5434,N_4951);
nand U6688 (N_6688,N_4888,N_5858);
or U6689 (N_6689,N_5315,N_5631);
xnor U6690 (N_6690,N_5568,N_5250);
nand U6691 (N_6691,N_4663,N_5727);
nor U6692 (N_6692,N_5098,N_5096);
and U6693 (N_6693,N_5095,N_4996);
nor U6694 (N_6694,N_4850,N_5341);
and U6695 (N_6695,N_4865,N_4741);
nand U6696 (N_6696,N_4759,N_4639);
xnor U6697 (N_6697,N_5383,N_5517);
or U6698 (N_6698,N_4710,N_5049);
nand U6699 (N_6699,N_5166,N_5709);
or U6700 (N_6700,N_4756,N_4695);
nor U6701 (N_6701,N_5364,N_5776);
nand U6702 (N_6702,N_4551,N_5504);
and U6703 (N_6703,N_5265,N_5171);
or U6704 (N_6704,N_4571,N_4685);
nor U6705 (N_6705,N_5296,N_5556);
xor U6706 (N_6706,N_4578,N_5264);
and U6707 (N_6707,N_5681,N_5480);
nand U6708 (N_6708,N_5952,N_5407);
nor U6709 (N_6709,N_5692,N_4843);
nand U6710 (N_6710,N_4853,N_5721);
nand U6711 (N_6711,N_5921,N_4801);
nor U6712 (N_6712,N_5156,N_5378);
xor U6713 (N_6713,N_5617,N_5022);
nor U6714 (N_6714,N_5540,N_4555);
or U6715 (N_6715,N_4905,N_4566);
or U6716 (N_6716,N_5443,N_5140);
nor U6717 (N_6717,N_5453,N_5733);
or U6718 (N_6718,N_5906,N_4978);
nor U6719 (N_6719,N_5474,N_5922);
xor U6720 (N_6720,N_5864,N_4697);
and U6721 (N_6721,N_5414,N_5871);
nor U6722 (N_6722,N_5624,N_4608);
or U6723 (N_6723,N_5311,N_5475);
and U6724 (N_6724,N_5803,N_4679);
nand U6725 (N_6725,N_5603,N_5920);
and U6726 (N_6726,N_4711,N_5361);
nand U6727 (N_6727,N_5100,N_5464);
and U6728 (N_6728,N_5927,N_5626);
nand U6729 (N_6729,N_5024,N_4833);
nand U6730 (N_6730,N_4927,N_5270);
or U6731 (N_6731,N_5214,N_4761);
or U6732 (N_6732,N_4594,N_4900);
or U6733 (N_6733,N_4886,N_5620);
and U6734 (N_6734,N_4995,N_5489);
nand U6735 (N_6735,N_4864,N_5113);
xnor U6736 (N_6736,N_5745,N_5257);
nand U6737 (N_6737,N_5466,N_5230);
nand U6738 (N_6738,N_5195,N_5565);
nor U6739 (N_6739,N_4887,N_5887);
or U6740 (N_6740,N_5330,N_5660);
nor U6741 (N_6741,N_5299,N_5408);
nand U6742 (N_6742,N_5798,N_4750);
and U6743 (N_6743,N_4624,N_5225);
nand U6744 (N_6744,N_5461,N_5488);
or U6745 (N_6745,N_5204,N_5728);
nor U6746 (N_6746,N_5463,N_5804);
and U6747 (N_6747,N_4934,N_5131);
or U6748 (N_6748,N_5514,N_5827);
and U6749 (N_6749,N_5737,N_5891);
or U6750 (N_6750,N_5834,N_5741);
nor U6751 (N_6751,N_4608,N_4514);
xor U6752 (N_6752,N_5501,N_5478);
nand U6753 (N_6753,N_4576,N_4805);
nor U6754 (N_6754,N_5739,N_5280);
nor U6755 (N_6755,N_4889,N_5241);
or U6756 (N_6756,N_4683,N_5150);
and U6757 (N_6757,N_5059,N_5480);
and U6758 (N_6758,N_5603,N_5815);
or U6759 (N_6759,N_5254,N_5520);
nand U6760 (N_6760,N_5670,N_5819);
and U6761 (N_6761,N_5189,N_5570);
or U6762 (N_6762,N_4522,N_5200);
or U6763 (N_6763,N_5591,N_5497);
and U6764 (N_6764,N_5862,N_4762);
or U6765 (N_6765,N_5916,N_4504);
or U6766 (N_6766,N_5656,N_5107);
or U6767 (N_6767,N_5315,N_5665);
and U6768 (N_6768,N_5560,N_5176);
and U6769 (N_6769,N_5421,N_4835);
or U6770 (N_6770,N_4528,N_4603);
nor U6771 (N_6771,N_5155,N_5366);
nand U6772 (N_6772,N_5703,N_4910);
or U6773 (N_6773,N_5999,N_5941);
or U6774 (N_6774,N_4836,N_4684);
and U6775 (N_6775,N_5601,N_4707);
nand U6776 (N_6776,N_5654,N_5692);
and U6777 (N_6777,N_5317,N_5571);
xor U6778 (N_6778,N_4647,N_5474);
nand U6779 (N_6779,N_4722,N_5236);
or U6780 (N_6780,N_4505,N_5044);
or U6781 (N_6781,N_5136,N_5708);
and U6782 (N_6782,N_5494,N_4590);
xnor U6783 (N_6783,N_5618,N_5969);
and U6784 (N_6784,N_5518,N_4973);
or U6785 (N_6785,N_5744,N_4973);
nand U6786 (N_6786,N_5320,N_5291);
and U6787 (N_6787,N_5113,N_5811);
and U6788 (N_6788,N_4824,N_4884);
or U6789 (N_6789,N_5147,N_5291);
and U6790 (N_6790,N_5786,N_4788);
and U6791 (N_6791,N_5331,N_4916);
xor U6792 (N_6792,N_5745,N_5068);
and U6793 (N_6793,N_5941,N_5031);
and U6794 (N_6794,N_5228,N_4558);
or U6795 (N_6795,N_4934,N_5740);
or U6796 (N_6796,N_5906,N_5879);
nand U6797 (N_6797,N_4622,N_4530);
and U6798 (N_6798,N_5717,N_5827);
xnor U6799 (N_6799,N_4619,N_5984);
nand U6800 (N_6800,N_5641,N_4737);
nand U6801 (N_6801,N_4539,N_5942);
nor U6802 (N_6802,N_4835,N_5728);
or U6803 (N_6803,N_5220,N_5589);
nor U6804 (N_6804,N_5745,N_5752);
and U6805 (N_6805,N_5129,N_5001);
or U6806 (N_6806,N_5027,N_5617);
or U6807 (N_6807,N_4597,N_5945);
or U6808 (N_6808,N_5614,N_5087);
or U6809 (N_6809,N_5425,N_5963);
nand U6810 (N_6810,N_5330,N_5915);
or U6811 (N_6811,N_5763,N_4723);
nand U6812 (N_6812,N_5908,N_5505);
nor U6813 (N_6813,N_5375,N_4866);
or U6814 (N_6814,N_5009,N_4739);
nor U6815 (N_6815,N_5131,N_5285);
nor U6816 (N_6816,N_5653,N_5634);
nor U6817 (N_6817,N_5007,N_5476);
and U6818 (N_6818,N_5343,N_5357);
nor U6819 (N_6819,N_4798,N_5852);
nor U6820 (N_6820,N_5257,N_5404);
nand U6821 (N_6821,N_5341,N_4716);
and U6822 (N_6822,N_5630,N_4777);
nand U6823 (N_6823,N_5536,N_5898);
xor U6824 (N_6824,N_5714,N_5473);
nand U6825 (N_6825,N_5123,N_5962);
and U6826 (N_6826,N_5831,N_5726);
or U6827 (N_6827,N_5416,N_4560);
xor U6828 (N_6828,N_5058,N_4989);
or U6829 (N_6829,N_5673,N_4756);
nor U6830 (N_6830,N_5776,N_5275);
and U6831 (N_6831,N_5160,N_5107);
and U6832 (N_6832,N_5086,N_5447);
xnor U6833 (N_6833,N_5572,N_5971);
nor U6834 (N_6834,N_5844,N_5469);
nand U6835 (N_6835,N_4502,N_5520);
and U6836 (N_6836,N_5095,N_5173);
xnor U6837 (N_6837,N_5436,N_5471);
nor U6838 (N_6838,N_5166,N_4612);
and U6839 (N_6839,N_5566,N_5044);
xnor U6840 (N_6840,N_5573,N_4746);
and U6841 (N_6841,N_5516,N_5896);
or U6842 (N_6842,N_5512,N_5492);
nand U6843 (N_6843,N_4841,N_5738);
and U6844 (N_6844,N_5086,N_5239);
or U6845 (N_6845,N_5734,N_5866);
nand U6846 (N_6846,N_5855,N_4513);
or U6847 (N_6847,N_5662,N_5485);
nor U6848 (N_6848,N_5241,N_4595);
nor U6849 (N_6849,N_5468,N_4704);
and U6850 (N_6850,N_5990,N_4623);
or U6851 (N_6851,N_4866,N_5053);
nor U6852 (N_6852,N_5262,N_4635);
and U6853 (N_6853,N_5350,N_4628);
nor U6854 (N_6854,N_5927,N_5076);
or U6855 (N_6855,N_4907,N_5649);
or U6856 (N_6856,N_5465,N_5043);
or U6857 (N_6857,N_4502,N_5358);
xnor U6858 (N_6858,N_4618,N_5746);
nand U6859 (N_6859,N_5824,N_5812);
or U6860 (N_6860,N_5088,N_5910);
or U6861 (N_6861,N_4972,N_4767);
or U6862 (N_6862,N_5544,N_4962);
nand U6863 (N_6863,N_5918,N_5669);
nand U6864 (N_6864,N_5625,N_4846);
nand U6865 (N_6865,N_4915,N_4812);
nor U6866 (N_6866,N_5976,N_4640);
nand U6867 (N_6867,N_5032,N_5546);
nand U6868 (N_6868,N_5556,N_4909);
xor U6869 (N_6869,N_5655,N_5027);
nand U6870 (N_6870,N_5623,N_5729);
nand U6871 (N_6871,N_4586,N_5999);
xor U6872 (N_6872,N_5846,N_5400);
and U6873 (N_6873,N_4699,N_4502);
nand U6874 (N_6874,N_5865,N_5029);
nor U6875 (N_6875,N_5652,N_5455);
xor U6876 (N_6876,N_5486,N_5417);
or U6877 (N_6877,N_4754,N_5159);
or U6878 (N_6878,N_5826,N_4532);
or U6879 (N_6879,N_4966,N_5207);
or U6880 (N_6880,N_5016,N_4693);
nor U6881 (N_6881,N_5557,N_5061);
nand U6882 (N_6882,N_4850,N_4679);
nand U6883 (N_6883,N_5252,N_5512);
nor U6884 (N_6884,N_5660,N_5431);
nor U6885 (N_6885,N_5381,N_5901);
nor U6886 (N_6886,N_5586,N_4961);
xnor U6887 (N_6887,N_4878,N_5150);
or U6888 (N_6888,N_4948,N_4953);
nand U6889 (N_6889,N_5554,N_5892);
or U6890 (N_6890,N_5417,N_5808);
nand U6891 (N_6891,N_4751,N_5346);
nand U6892 (N_6892,N_4679,N_5018);
nor U6893 (N_6893,N_4976,N_5787);
and U6894 (N_6894,N_5734,N_4782);
nand U6895 (N_6895,N_5927,N_4775);
or U6896 (N_6896,N_5227,N_4775);
and U6897 (N_6897,N_4957,N_4757);
nor U6898 (N_6898,N_5532,N_5027);
or U6899 (N_6899,N_5382,N_5567);
and U6900 (N_6900,N_4641,N_4715);
nand U6901 (N_6901,N_5237,N_4840);
and U6902 (N_6902,N_4798,N_4568);
or U6903 (N_6903,N_5844,N_4795);
nor U6904 (N_6904,N_5751,N_5230);
or U6905 (N_6905,N_4785,N_4668);
and U6906 (N_6906,N_5323,N_5244);
and U6907 (N_6907,N_5097,N_5535);
nand U6908 (N_6908,N_5790,N_4698);
nand U6909 (N_6909,N_5869,N_4842);
xnor U6910 (N_6910,N_4765,N_5451);
or U6911 (N_6911,N_5883,N_5862);
nor U6912 (N_6912,N_5736,N_5780);
nor U6913 (N_6913,N_5344,N_5428);
nor U6914 (N_6914,N_5436,N_5492);
and U6915 (N_6915,N_5293,N_5478);
and U6916 (N_6916,N_4631,N_5391);
or U6917 (N_6917,N_5579,N_4998);
nand U6918 (N_6918,N_5762,N_4525);
xor U6919 (N_6919,N_5235,N_4892);
or U6920 (N_6920,N_4579,N_4989);
nor U6921 (N_6921,N_5807,N_4875);
or U6922 (N_6922,N_5438,N_5918);
and U6923 (N_6923,N_4634,N_4564);
nor U6924 (N_6924,N_5494,N_4888);
nand U6925 (N_6925,N_4961,N_5992);
xor U6926 (N_6926,N_5385,N_4570);
or U6927 (N_6927,N_5793,N_4621);
or U6928 (N_6928,N_4927,N_5682);
nor U6929 (N_6929,N_4821,N_4675);
and U6930 (N_6930,N_5666,N_5939);
and U6931 (N_6931,N_4966,N_5627);
and U6932 (N_6932,N_5059,N_5030);
nand U6933 (N_6933,N_5935,N_5696);
or U6934 (N_6934,N_4927,N_5669);
or U6935 (N_6935,N_5960,N_5705);
nor U6936 (N_6936,N_5518,N_5700);
and U6937 (N_6937,N_4875,N_4743);
or U6938 (N_6938,N_5987,N_4960);
nand U6939 (N_6939,N_5706,N_5140);
and U6940 (N_6940,N_5893,N_5273);
and U6941 (N_6941,N_5211,N_4771);
xor U6942 (N_6942,N_5223,N_5724);
nand U6943 (N_6943,N_5067,N_4825);
and U6944 (N_6944,N_5935,N_4557);
or U6945 (N_6945,N_5379,N_4747);
nand U6946 (N_6946,N_5489,N_4998);
nor U6947 (N_6947,N_5310,N_4876);
nand U6948 (N_6948,N_5569,N_4792);
and U6949 (N_6949,N_4907,N_5066);
xor U6950 (N_6950,N_5043,N_5319);
nand U6951 (N_6951,N_5885,N_5301);
xor U6952 (N_6952,N_5009,N_5754);
nand U6953 (N_6953,N_5725,N_5172);
and U6954 (N_6954,N_5865,N_5336);
and U6955 (N_6955,N_4792,N_4629);
or U6956 (N_6956,N_5844,N_5261);
or U6957 (N_6957,N_4961,N_5990);
nand U6958 (N_6958,N_5787,N_5913);
nor U6959 (N_6959,N_5220,N_5794);
xnor U6960 (N_6960,N_5336,N_4830);
xnor U6961 (N_6961,N_5630,N_5446);
nor U6962 (N_6962,N_4682,N_4971);
and U6963 (N_6963,N_4618,N_5480);
or U6964 (N_6964,N_4957,N_5771);
and U6965 (N_6965,N_5313,N_5454);
and U6966 (N_6966,N_4633,N_5384);
and U6967 (N_6967,N_5059,N_4795);
or U6968 (N_6968,N_5726,N_5982);
nand U6969 (N_6969,N_5098,N_4573);
nor U6970 (N_6970,N_5723,N_4558);
or U6971 (N_6971,N_5095,N_5915);
nor U6972 (N_6972,N_5046,N_5191);
nand U6973 (N_6973,N_4858,N_4727);
nor U6974 (N_6974,N_5370,N_5828);
nor U6975 (N_6975,N_4676,N_5058);
or U6976 (N_6976,N_5928,N_4724);
and U6977 (N_6977,N_4555,N_5239);
or U6978 (N_6978,N_5488,N_5911);
nand U6979 (N_6979,N_5753,N_5713);
nand U6980 (N_6980,N_5172,N_5057);
and U6981 (N_6981,N_5717,N_5193);
nor U6982 (N_6982,N_5924,N_4862);
and U6983 (N_6983,N_4532,N_4740);
nand U6984 (N_6984,N_5639,N_5514);
or U6985 (N_6985,N_5258,N_5139);
nand U6986 (N_6986,N_4853,N_4829);
nor U6987 (N_6987,N_5835,N_5196);
and U6988 (N_6988,N_5775,N_5107);
or U6989 (N_6989,N_5729,N_5402);
nand U6990 (N_6990,N_5755,N_5177);
or U6991 (N_6991,N_5804,N_5123);
nor U6992 (N_6992,N_5551,N_5578);
and U6993 (N_6993,N_5383,N_4976);
xnor U6994 (N_6994,N_5386,N_5226);
xnor U6995 (N_6995,N_5009,N_5274);
nand U6996 (N_6996,N_5275,N_5121);
nor U6997 (N_6997,N_5982,N_4785);
nand U6998 (N_6998,N_4991,N_4579);
nand U6999 (N_6999,N_4981,N_5097);
nand U7000 (N_7000,N_5413,N_5878);
or U7001 (N_7001,N_5408,N_5443);
nor U7002 (N_7002,N_4953,N_5184);
nor U7003 (N_7003,N_5818,N_4515);
or U7004 (N_7004,N_5214,N_4576);
nand U7005 (N_7005,N_5628,N_5990);
xor U7006 (N_7006,N_5244,N_5534);
nand U7007 (N_7007,N_5983,N_4719);
or U7008 (N_7008,N_5414,N_4973);
nand U7009 (N_7009,N_5988,N_5742);
or U7010 (N_7010,N_5562,N_5671);
or U7011 (N_7011,N_5624,N_5323);
nand U7012 (N_7012,N_5135,N_5104);
nand U7013 (N_7013,N_4818,N_4914);
and U7014 (N_7014,N_4792,N_4909);
nand U7015 (N_7015,N_5348,N_4782);
nor U7016 (N_7016,N_5065,N_5416);
or U7017 (N_7017,N_5345,N_5061);
and U7018 (N_7018,N_5542,N_5814);
xor U7019 (N_7019,N_5511,N_5207);
nor U7020 (N_7020,N_4587,N_4549);
nand U7021 (N_7021,N_5373,N_5791);
nand U7022 (N_7022,N_4942,N_4660);
xor U7023 (N_7023,N_5360,N_5554);
nor U7024 (N_7024,N_5836,N_5430);
or U7025 (N_7025,N_4982,N_5069);
nand U7026 (N_7026,N_4658,N_5471);
and U7027 (N_7027,N_5435,N_5448);
and U7028 (N_7028,N_5872,N_4761);
nand U7029 (N_7029,N_4871,N_5153);
or U7030 (N_7030,N_5271,N_5430);
nor U7031 (N_7031,N_4609,N_5790);
or U7032 (N_7032,N_4835,N_5197);
or U7033 (N_7033,N_4695,N_5391);
nand U7034 (N_7034,N_5731,N_4660);
nand U7035 (N_7035,N_5128,N_4586);
nand U7036 (N_7036,N_5926,N_5766);
nor U7037 (N_7037,N_5105,N_5073);
nand U7038 (N_7038,N_5402,N_4673);
nand U7039 (N_7039,N_4723,N_5518);
or U7040 (N_7040,N_4900,N_5022);
nor U7041 (N_7041,N_5378,N_4810);
or U7042 (N_7042,N_5526,N_5277);
nor U7043 (N_7043,N_5845,N_5906);
nor U7044 (N_7044,N_5254,N_4869);
xor U7045 (N_7045,N_4995,N_5457);
xor U7046 (N_7046,N_4772,N_4788);
and U7047 (N_7047,N_5221,N_4516);
nor U7048 (N_7048,N_5308,N_4859);
and U7049 (N_7049,N_5427,N_4756);
nand U7050 (N_7050,N_5074,N_4648);
xor U7051 (N_7051,N_5918,N_4903);
or U7052 (N_7052,N_5818,N_5154);
and U7053 (N_7053,N_5324,N_5412);
nand U7054 (N_7054,N_5006,N_5328);
or U7055 (N_7055,N_5442,N_4692);
or U7056 (N_7056,N_5032,N_5840);
nor U7057 (N_7057,N_5692,N_4730);
xnor U7058 (N_7058,N_4846,N_4807);
or U7059 (N_7059,N_5673,N_5513);
or U7060 (N_7060,N_4912,N_5602);
nand U7061 (N_7061,N_5581,N_5680);
nand U7062 (N_7062,N_5446,N_5958);
or U7063 (N_7063,N_4515,N_5231);
nor U7064 (N_7064,N_5702,N_5408);
nand U7065 (N_7065,N_4740,N_5841);
or U7066 (N_7066,N_5157,N_5691);
xor U7067 (N_7067,N_4811,N_4873);
xor U7068 (N_7068,N_5783,N_5276);
nor U7069 (N_7069,N_5951,N_5792);
and U7070 (N_7070,N_5946,N_5599);
nor U7071 (N_7071,N_4581,N_5480);
nand U7072 (N_7072,N_5073,N_4639);
nor U7073 (N_7073,N_5073,N_5257);
nor U7074 (N_7074,N_5238,N_4793);
xor U7075 (N_7075,N_5951,N_4946);
nand U7076 (N_7076,N_4886,N_5829);
nor U7077 (N_7077,N_4707,N_4870);
nor U7078 (N_7078,N_5752,N_4598);
nor U7079 (N_7079,N_5257,N_5674);
nor U7080 (N_7080,N_5814,N_5197);
nand U7081 (N_7081,N_5748,N_5439);
and U7082 (N_7082,N_5007,N_5929);
and U7083 (N_7083,N_5785,N_4920);
and U7084 (N_7084,N_5935,N_5805);
and U7085 (N_7085,N_4820,N_4577);
and U7086 (N_7086,N_5611,N_5504);
and U7087 (N_7087,N_4541,N_4617);
nor U7088 (N_7088,N_5038,N_5837);
nand U7089 (N_7089,N_5276,N_5540);
or U7090 (N_7090,N_5919,N_5162);
xor U7091 (N_7091,N_5466,N_5546);
and U7092 (N_7092,N_5592,N_5161);
nor U7093 (N_7093,N_5771,N_5422);
nand U7094 (N_7094,N_4557,N_5696);
nand U7095 (N_7095,N_4888,N_5561);
or U7096 (N_7096,N_5867,N_5815);
nor U7097 (N_7097,N_4694,N_5299);
and U7098 (N_7098,N_4694,N_5311);
nor U7099 (N_7099,N_5684,N_5303);
or U7100 (N_7100,N_4580,N_5731);
nand U7101 (N_7101,N_5467,N_5099);
and U7102 (N_7102,N_5160,N_5088);
or U7103 (N_7103,N_4514,N_5817);
nor U7104 (N_7104,N_5093,N_4628);
or U7105 (N_7105,N_5888,N_5738);
and U7106 (N_7106,N_5125,N_5155);
nand U7107 (N_7107,N_4822,N_4945);
nor U7108 (N_7108,N_5832,N_5154);
nor U7109 (N_7109,N_5322,N_4792);
nor U7110 (N_7110,N_5997,N_4595);
nor U7111 (N_7111,N_4917,N_5727);
nor U7112 (N_7112,N_5633,N_5656);
and U7113 (N_7113,N_4734,N_4795);
and U7114 (N_7114,N_4798,N_5647);
nor U7115 (N_7115,N_4724,N_5559);
and U7116 (N_7116,N_5625,N_4697);
nand U7117 (N_7117,N_5977,N_5337);
xor U7118 (N_7118,N_4690,N_5924);
nor U7119 (N_7119,N_4830,N_5176);
and U7120 (N_7120,N_5889,N_5630);
or U7121 (N_7121,N_5604,N_4834);
or U7122 (N_7122,N_5338,N_5619);
or U7123 (N_7123,N_5225,N_4923);
nor U7124 (N_7124,N_5477,N_5392);
or U7125 (N_7125,N_4730,N_5936);
nand U7126 (N_7126,N_4521,N_5146);
nand U7127 (N_7127,N_5789,N_4969);
nor U7128 (N_7128,N_5228,N_5296);
nand U7129 (N_7129,N_4601,N_4747);
and U7130 (N_7130,N_4905,N_5999);
nor U7131 (N_7131,N_5377,N_5299);
nor U7132 (N_7132,N_4836,N_5762);
and U7133 (N_7133,N_5686,N_5206);
and U7134 (N_7134,N_5215,N_5832);
nor U7135 (N_7135,N_5149,N_4817);
xor U7136 (N_7136,N_5799,N_4991);
and U7137 (N_7137,N_4816,N_4521);
nor U7138 (N_7138,N_5370,N_4500);
or U7139 (N_7139,N_5092,N_4602);
and U7140 (N_7140,N_5455,N_4784);
or U7141 (N_7141,N_4540,N_5849);
nor U7142 (N_7142,N_4708,N_5810);
nor U7143 (N_7143,N_5314,N_5814);
nand U7144 (N_7144,N_5346,N_5612);
and U7145 (N_7145,N_5234,N_5242);
nand U7146 (N_7146,N_5562,N_5460);
or U7147 (N_7147,N_4605,N_5030);
and U7148 (N_7148,N_4931,N_4717);
and U7149 (N_7149,N_5991,N_4874);
or U7150 (N_7150,N_5354,N_4997);
nand U7151 (N_7151,N_5983,N_5266);
and U7152 (N_7152,N_5226,N_5762);
nor U7153 (N_7153,N_4517,N_4943);
and U7154 (N_7154,N_5643,N_4921);
nand U7155 (N_7155,N_5256,N_4673);
nand U7156 (N_7156,N_5755,N_5600);
and U7157 (N_7157,N_4764,N_5139);
nand U7158 (N_7158,N_5797,N_5234);
nand U7159 (N_7159,N_5637,N_5619);
or U7160 (N_7160,N_5915,N_5626);
nor U7161 (N_7161,N_4910,N_4994);
nor U7162 (N_7162,N_5827,N_5977);
nor U7163 (N_7163,N_5349,N_5345);
and U7164 (N_7164,N_4917,N_4514);
and U7165 (N_7165,N_5143,N_4903);
nor U7166 (N_7166,N_5281,N_5087);
nor U7167 (N_7167,N_4963,N_5957);
nand U7168 (N_7168,N_5339,N_4835);
nand U7169 (N_7169,N_5073,N_5909);
nand U7170 (N_7170,N_5003,N_5941);
or U7171 (N_7171,N_5452,N_5907);
nand U7172 (N_7172,N_4582,N_5033);
nand U7173 (N_7173,N_4626,N_5947);
nor U7174 (N_7174,N_4922,N_5143);
and U7175 (N_7175,N_4897,N_5950);
nor U7176 (N_7176,N_4665,N_4693);
nor U7177 (N_7177,N_4702,N_4528);
nor U7178 (N_7178,N_5119,N_4947);
nor U7179 (N_7179,N_5284,N_5213);
or U7180 (N_7180,N_5303,N_5661);
nand U7181 (N_7181,N_5954,N_5768);
nor U7182 (N_7182,N_4769,N_5418);
and U7183 (N_7183,N_5712,N_4816);
and U7184 (N_7184,N_4506,N_4555);
and U7185 (N_7185,N_5050,N_5949);
and U7186 (N_7186,N_4720,N_5074);
and U7187 (N_7187,N_4799,N_4603);
or U7188 (N_7188,N_5627,N_4780);
nand U7189 (N_7189,N_5892,N_5686);
nand U7190 (N_7190,N_4623,N_4826);
xor U7191 (N_7191,N_5394,N_5728);
and U7192 (N_7192,N_5168,N_5133);
nand U7193 (N_7193,N_5901,N_4561);
nor U7194 (N_7194,N_5560,N_5754);
nor U7195 (N_7195,N_5801,N_5061);
nand U7196 (N_7196,N_5255,N_5070);
or U7197 (N_7197,N_5860,N_5619);
xnor U7198 (N_7198,N_4839,N_4995);
xnor U7199 (N_7199,N_5524,N_5137);
or U7200 (N_7200,N_5452,N_5636);
xor U7201 (N_7201,N_5810,N_5870);
and U7202 (N_7202,N_5189,N_4867);
nand U7203 (N_7203,N_4879,N_5115);
and U7204 (N_7204,N_5657,N_4691);
nand U7205 (N_7205,N_5501,N_5778);
xor U7206 (N_7206,N_5000,N_5617);
or U7207 (N_7207,N_5532,N_5880);
and U7208 (N_7208,N_4704,N_4583);
and U7209 (N_7209,N_5617,N_5071);
nor U7210 (N_7210,N_5613,N_5625);
nor U7211 (N_7211,N_5365,N_5557);
or U7212 (N_7212,N_5704,N_4868);
and U7213 (N_7213,N_4638,N_5303);
nor U7214 (N_7214,N_5660,N_4792);
and U7215 (N_7215,N_5001,N_5510);
nand U7216 (N_7216,N_5439,N_5892);
nand U7217 (N_7217,N_5164,N_5932);
or U7218 (N_7218,N_5618,N_5815);
nand U7219 (N_7219,N_5549,N_5424);
nand U7220 (N_7220,N_5235,N_4844);
and U7221 (N_7221,N_5867,N_5624);
or U7222 (N_7222,N_5850,N_4746);
nor U7223 (N_7223,N_5486,N_5263);
and U7224 (N_7224,N_5057,N_5850);
and U7225 (N_7225,N_5704,N_4908);
and U7226 (N_7226,N_5403,N_5142);
nor U7227 (N_7227,N_5578,N_4879);
nand U7228 (N_7228,N_4807,N_4781);
xor U7229 (N_7229,N_5245,N_5300);
nor U7230 (N_7230,N_4813,N_5062);
nand U7231 (N_7231,N_5936,N_4864);
or U7232 (N_7232,N_5174,N_5883);
xnor U7233 (N_7233,N_5673,N_5525);
xor U7234 (N_7234,N_5720,N_4888);
or U7235 (N_7235,N_5094,N_4732);
and U7236 (N_7236,N_5969,N_5790);
nor U7237 (N_7237,N_5327,N_5587);
nor U7238 (N_7238,N_5738,N_5664);
nand U7239 (N_7239,N_5958,N_5651);
or U7240 (N_7240,N_5603,N_5954);
nor U7241 (N_7241,N_4558,N_5159);
and U7242 (N_7242,N_5335,N_5264);
nor U7243 (N_7243,N_5754,N_5341);
and U7244 (N_7244,N_5964,N_5886);
or U7245 (N_7245,N_5754,N_5301);
nand U7246 (N_7246,N_5992,N_4938);
and U7247 (N_7247,N_5821,N_4520);
and U7248 (N_7248,N_5629,N_5997);
nor U7249 (N_7249,N_5711,N_5877);
and U7250 (N_7250,N_4858,N_4768);
nor U7251 (N_7251,N_4979,N_5371);
and U7252 (N_7252,N_4628,N_4825);
nand U7253 (N_7253,N_5386,N_4570);
nand U7254 (N_7254,N_5938,N_5397);
or U7255 (N_7255,N_5102,N_5263);
xor U7256 (N_7256,N_5009,N_4880);
or U7257 (N_7257,N_4903,N_4859);
nor U7258 (N_7258,N_5890,N_5508);
nor U7259 (N_7259,N_4987,N_4940);
and U7260 (N_7260,N_4627,N_5767);
nand U7261 (N_7261,N_5596,N_5541);
nor U7262 (N_7262,N_5276,N_4846);
nor U7263 (N_7263,N_5506,N_4988);
and U7264 (N_7264,N_4719,N_5758);
xor U7265 (N_7265,N_4682,N_5350);
or U7266 (N_7266,N_4824,N_5891);
and U7267 (N_7267,N_5456,N_5137);
and U7268 (N_7268,N_4726,N_4509);
or U7269 (N_7269,N_4989,N_5781);
or U7270 (N_7270,N_5902,N_5718);
nand U7271 (N_7271,N_4716,N_4970);
nor U7272 (N_7272,N_4822,N_5620);
xor U7273 (N_7273,N_4678,N_5266);
or U7274 (N_7274,N_5056,N_4995);
nand U7275 (N_7275,N_5758,N_4952);
nand U7276 (N_7276,N_5186,N_5529);
nand U7277 (N_7277,N_5752,N_5416);
and U7278 (N_7278,N_5477,N_4625);
or U7279 (N_7279,N_5288,N_5402);
xnor U7280 (N_7280,N_4829,N_4990);
xnor U7281 (N_7281,N_4909,N_5213);
nand U7282 (N_7282,N_5413,N_5973);
and U7283 (N_7283,N_4819,N_5172);
and U7284 (N_7284,N_5527,N_5985);
or U7285 (N_7285,N_4662,N_5871);
and U7286 (N_7286,N_5268,N_4563);
nor U7287 (N_7287,N_4555,N_5778);
and U7288 (N_7288,N_5321,N_4554);
nand U7289 (N_7289,N_5676,N_5706);
and U7290 (N_7290,N_5683,N_5247);
xor U7291 (N_7291,N_5415,N_4890);
nor U7292 (N_7292,N_5742,N_4956);
xor U7293 (N_7293,N_4963,N_4713);
nand U7294 (N_7294,N_5043,N_5628);
and U7295 (N_7295,N_5848,N_4773);
and U7296 (N_7296,N_5552,N_4607);
nor U7297 (N_7297,N_4997,N_5704);
nor U7298 (N_7298,N_4782,N_5976);
and U7299 (N_7299,N_5945,N_5584);
or U7300 (N_7300,N_5060,N_5844);
and U7301 (N_7301,N_5970,N_5222);
nand U7302 (N_7302,N_5329,N_4606);
nand U7303 (N_7303,N_5764,N_4517);
nor U7304 (N_7304,N_5624,N_5239);
nand U7305 (N_7305,N_5947,N_5784);
nor U7306 (N_7306,N_5364,N_5782);
and U7307 (N_7307,N_4747,N_5283);
nand U7308 (N_7308,N_5410,N_5906);
and U7309 (N_7309,N_5929,N_5060);
or U7310 (N_7310,N_4570,N_5526);
and U7311 (N_7311,N_4766,N_5430);
nand U7312 (N_7312,N_5963,N_5304);
or U7313 (N_7313,N_5695,N_5852);
or U7314 (N_7314,N_5482,N_5671);
nor U7315 (N_7315,N_4500,N_4992);
xnor U7316 (N_7316,N_5532,N_5960);
nor U7317 (N_7317,N_4841,N_4700);
and U7318 (N_7318,N_4728,N_5914);
nand U7319 (N_7319,N_4925,N_5097);
nand U7320 (N_7320,N_5939,N_5137);
and U7321 (N_7321,N_5328,N_4955);
and U7322 (N_7322,N_5570,N_5652);
nand U7323 (N_7323,N_5613,N_5594);
and U7324 (N_7324,N_5743,N_4697);
or U7325 (N_7325,N_4973,N_4844);
and U7326 (N_7326,N_4763,N_5236);
and U7327 (N_7327,N_5451,N_5101);
nand U7328 (N_7328,N_4858,N_4807);
and U7329 (N_7329,N_5627,N_4507);
and U7330 (N_7330,N_5764,N_5792);
xnor U7331 (N_7331,N_4729,N_4892);
nand U7332 (N_7332,N_5214,N_5547);
nand U7333 (N_7333,N_5393,N_4551);
xor U7334 (N_7334,N_5350,N_5397);
nand U7335 (N_7335,N_5106,N_4687);
or U7336 (N_7336,N_5796,N_5121);
or U7337 (N_7337,N_5324,N_4725);
and U7338 (N_7338,N_5864,N_5917);
xnor U7339 (N_7339,N_5316,N_5185);
and U7340 (N_7340,N_5897,N_5512);
or U7341 (N_7341,N_4834,N_5371);
and U7342 (N_7342,N_5757,N_5987);
nand U7343 (N_7343,N_5408,N_5258);
nand U7344 (N_7344,N_5083,N_5657);
and U7345 (N_7345,N_5794,N_5833);
or U7346 (N_7346,N_4636,N_4730);
or U7347 (N_7347,N_5348,N_4711);
xnor U7348 (N_7348,N_4930,N_5624);
or U7349 (N_7349,N_5040,N_5469);
and U7350 (N_7350,N_5845,N_4632);
nor U7351 (N_7351,N_5945,N_4690);
nand U7352 (N_7352,N_5293,N_5862);
nor U7353 (N_7353,N_4817,N_4999);
and U7354 (N_7354,N_4759,N_5157);
and U7355 (N_7355,N_4820,N_5904);
and U7356 (N_7356,N_4682,N_4608);
and U7357 (N_7357,N_5782,N_5521);
nand U7358 (N_7358,N_5476,N_4820);
nor U7359 (N_7359,N_5853,N_4728);
nor U7360 (N_7360,N_5396,N_4786);
and U7361 (N_7361,N_5175,N_5454);
nor U7362 (N_7362,N_5159,N_4827);
or U7363 (N_7363,N_5161,N_4947);
nor U7364 (N_7364,N_5849,N_5633);
nor U7365 (N_7365,N_4798,N_5763);
nor U7366 (N_7366,N_5186,N_5575);
and U7367 (N_7367,N_4835,N_4571);
or U7368 (N_7368,N_5471,N_5738);
nor U7369 (N_7369,N_5208,N_5266);
xnor U7370 (N_7370,N_5694,N_4690);
nand U7371 (N_7371,N_5086,N_4927);
or U7372 (N_7372,N_5218,N_4828);
xnor U7373 (N_7373,N_5741,N_5610);
or U7374 (N_7374,N_5333,N_5429);
nor U7375 (N_7375,N_5925,N_5739);
nor U7376 (N_7376,N_4593,N_5566);
nand U7377 (N_7377,N_5979,N_5093);
nand U7378 (N_7378,N_5345,N_5311);
nand U7379 (N_7379,N_4925,N_5474);
nand U7380 (N_7380,N_5034,N_5250);
and U7381 (N_7381,N_5324,N_5257);
or U7382 (N_7382,N_4866,N_5274);
or U7383 (N_7383,N_5190,N_5410);
nand U7384 (N_7384,N_5319,N_5866);
or U7385 (N_7385,N_4505,N_5881);
and U7386 (N_7386,N_4968,N_4893);
or U7387 (N_7387,N_5570,N_5489);
nand U7388 (N_7388,N_5482,N_5053);
nand U7389 (N_7389,N_5684,N_5624);
and U7390 (N_7390,N_5521,N_5772);
nor U7391 (N_7391,N_4676,N_5851);
nand U7392 (N_7392,N_5674,N_5288);
or U7393 (N_7393,N_5031,N_5925);
or U7394 (N_7394,N_4596,N_5149);
and U7395 (N_7395,N_4826,N_5748);
nand U7396 (N_7396,N_4672,N_5993);
and U7397 (N_7397,N_4783,N_5835);
nor U7398 (N_7398,N_4803,N_4659);
or U7399 (N_7399,N_4980,N_4876);
nor U7400 (N_7400,N_5330,N_4981);
nor U7401 (N_7401,N_5467,N_5035);
or U7402 (N_7402,N_5774,N_5029);
xnor U7403 (N_7403,N_5276,N_5602);
and U7404 (N_7404,N_5248,N_5615);
nand U7405 (N_7405,N_5435,N_5176);
and U7406 (N_7406,N_5153,N_5964);
xnor U7407 (N_7407,N_5383,N_4793);
xor U7408 (N_7408,N_5378,N_5530);
and U7409 (N_7409,N_5078,N_4938);
and U7410 (N_7410,N_5613,N_5465);
or U7411 (N_7411,N_4564,N_5689);
nand U7412 (N_7412,N_4850,N_4634);
nand U7413 (N_7413,N_4725,N_4799);
xnor U7414 (N_7414,N_5150,N_5109);
nand U7415 (N_7415,N_5298,N_5072);
and U7416 (N_7416,N_5617,N_4515);
nor U7417 (N_7417,N_5960,N_5389);
nor U7418 (N_7418,N_5301,N_4691);
nand U7419 (N_7419,N_5322,N_5849);
and U7420 (N_7420,N_5922,N_4726);
and U7421 (N_7421,N_4841,N_5855);
and U7422 (N_7422,N_4638,N_5285);
nand U7423 (N_7423,N_4765,N_4509);
xor U7424 (N_7424,N_5733,N_5779);
and U7425 (N_7425,N_4818,N_5780);
nor U7426 (N_7426,N_5113,N_4625);
and U7427 (N_7427,N_5539,N_4732);
nor U7428 (N_7428,N_5400,N_5987);
nor U7429 (N_7429,N_5081,N_4614);
xnor U7430 (N_7430,N_4886,N_5952);
or U7431 (N_7431,N_5613,N_5748);
and U7432 (N_7432,N_5460,N_4990);
nor U7433 (N_7433,N_4632,N_4979);
nor U7434 (N_7434,N_4838,N_5009);
or U7435 (N_7435,N_5713,N_5736);
nand U7436 (N_7436,N_5754,N_4731);
nor U7437 (N_7437,N_5456,N_4575);
or U7438 (N_7438,N_5889,N_4614);
and U7439 (N_7439,N_4655,N_5513);
or U7440 (N_7440,N_4611,N_5058);
or U7441 (N_7441,N_5515,N_5593);
nor U7442 (N_7442,N_5178,N_4916);
xor U7443 (N_7443,N_4975,N_5258);
and U7444 (N_7444,N_4682,N_5490);
nand U7445 (N_7445,N_5916,N_5588);
nor U7446 (N_7446,N_5361,N_5041);
nor U7447 (N_7447,N_4624,N_5420);
xor U7448 (N_7448,N_5991,N_4574);
or U7449 (N_7449,N_5403,N_5635);
nor U7450 (N_7450,N_5586,N_4891);
nand U7451 (N_7451,N_5737,N_4772);
and U7452 (N_7452,N_5537,N_5391);
nor U7453 (N_7453,N_5366,N_4834);
nand U7454 (N_7454,N_4971,N_5660);
nor U7455 (N_7455,N_5218,N_4749);
nand U7456 (N_7456,N_5632,N_5628);
nand U7457 (N_7457,N_4885,N_5963);
nand U7458 (N_7458,N_5081,N_4576);
nand U7459 (N_7459,N_5408,N_5655);
or U7460 (N_7460,N_4954,N_5074);
xor U7461 (N_7461,N_4582,N_5376);
and U7462 (N_7462,N_5731,N_4670);
or U7463 (N_7463,N_5107,N_5453);
and U7464 (N_7464,N_5590,N_5240);
and U7465 (N_7465,N_5132,N_5191);
or U7466 (N_7466,N_5837,N_5431);
and U7467 (N_7467,N_4665,N_4918);
nand U7468 (N_7468,N_5380,N_5281);
or U7469 (N_7469,N_5174,N_4867);
nand U7470 (N_7470,N_5984,N_5220);
and U7471 (N_7471,N_4561,N_5407);
nor U7472 (N_7472,N_5403,N_5321);
or U7473 (N_7473,N_5369,N_5350);
nand U7474 (N_7474,N_4910,N_5728);
nor U7475 (N_7475,N_5623,N_5766);
and U7476 (N_7476,N_4762,N_5171);
xnor U7477 (N_7477,N_4813,N_5256);
or U7478 (N_7478,N_5819,N_5870);
nor U7479 (N_7479,N_4976,N_5089);
or U7480 (N_7480,N_5987,N_5539);
or U7481 (N_7481,N_4812,N_5574);
nor U7482 (N_7482,N_5283,N_4678);
xor U7483 (N_7483,N_5131,N_4890);
and U7484 (N_7484,N_5029,N_5002);
nand U7485 (N_7485,N_5799,N_5644);
xor U7486 (N_7486,N_4864,N_5102);
and U7487 (N_7487,N_5621,N_5448);
and U7488 (N_7488,N_4967,N_4832);
nand U7489 (N_7489,N_4629,N_4777);
nand U7490 (N_7490,N_5959,N_4621);
xor U7491 (N_7491,N_5535,N_4609);
nor U7492 (N_7492,N_5281,N_5517);
or U7493 (N_7493,N_5032,N_5989);
nand U7494 (N_7494,N_5738,N_4654);
nand U7495 (N_7495,N_5842,N_5024);
or U7496 (N_7496,N_5900,N_5651);
and U7497 (N_7497,N_5221,N_5336);
nand U7498 (N_7498,N_5369,N_5006);
nand U7499 (N_7499,N_5341,N_5464);
xor U7500 (N_7500,N_6878,N_6240);
and U7501 (N_7501,N_6162,N_6027);
nor U7502 (N_7502,N_7047,N_7171);
nand U7503 (N_7503,N_7105,N_7038);
and U7504 (N_7504,N_6875,N_6838);
and U7505 (N_7505,N_7003,N_7054);
and U7506 (N_7506,N_6450,N_7265);
or U7507 (N_7507,N_7396,N_6273);
or U7508 (N_7508,N_6228,N_7445);
nand U7509 (N_7509,N_6396,N_7410);
nor U7510 (N_7510,N_6511,N_6525);
nand U7511 (N_7511,N_7052,N_6800);
and U7512 (N_7512,N_6327,N_6121);
and U7513 (N_7513,N_6363,N_6248);
or U7514 (N_7514,N_7018,N_6245);
or U7515 (N_7515,N_7454,N_7013);
or U7516 (N_7516,N_7042,N_6891);
and U7517 (N_7517,N_6760,N_6215);
and U7518 (N_7518,N_6413,N_6792);
nand U7519 (N_7519,N_6138,N_6779);
nand U7520 (N_7520,N_6565,N_6866);
nand U7521 (N_7521,N_6671,N_6232);
nand U7522 (N_7522,N_6103,N_6177);
and U7523 (N_7523,N_6622,N_6345);
and U7524 (N_7524,N_6942,N_6764);
xor U7525 (N_7525,N_7148,N_7235);
xor U7526 (N_7526,N_7019,N_6064);
or U7527 (N_7527,N_6678,N_6881);
nand U7528 (N_7528,N_6674,N_6989);
or U7529 (N_7529,N_7205,N_7413);
xnor U7530 (N_7530,N_6262,N_6733);
nand U7531 (N_7531,N_6761,N_7168);
or U7532 (N_7532,N_7301,N_6333);
or U7533 (N_7533,N_6137,N_6068);
or U7534 (N_7534,N_6646,N_6855);
nand U7535 (N_7535,N_6583,N_6022);
or U7536 (N_7536,N_6863,N_7182);
and U7537 (N_7537,N_6729,N_6252);
nand U7538 (N_7538,N_6966,N_7362);
nor U7539 (N_7539,N_6578,N_7025);
nand U7540 (N_7540,N_6325,N_6210);
nand U7541 (N_7541,N_6642,N_7093);
and U7542 (N_7542,N_6604,N_6379);
nor U7543 (N_7543,N_7156,N_7474);
and U7544 (N_7544,N_7214,N_6939);
xnor U7545 (N_7545,N_6540,N_6432);
nand U7546 (N_7546,N_6174,N_6649);
and U7547 (N_7547,N_7473,N_7268);
nor U7548 (N_7548,N_6842,N_7333);
and U7549 (N_7549,N_6291,N_6999);
nand U7550 (N_7550,N_6282,N_6721);
nor U7551 (N_7551,N_6028,N_6380);
nand U7552 (N_7552,N_6487,N_6778);
and U7553 (N_7553,N_6735,N_7325);
nand U7554 (N_7554,N_6835,N_7437);
nor U7555 (N_7555,N_6915,N_6600);
and U7556 (N_7556,N_7056,N_6912);
or U7557 (N_7557,N_7067,N_6482);
nand U7558 (N_7558,N_7299,N_6148);
xor U7559 (N_7559,N_6935,N_7045);
or U7560 (N_7560,N_6048,N_7210);
xnor U7561 (N_7561,N_6595,N_7359);
nor U7562 (N_7562,N_6020,N_6627);
and U7563 (N_7563,N_6730,N_6417);
or U7564 (N_7564,N_7203,N_7024);
nor U7565 (N_7565,N_7406,N_6409);
and U7566 (N_7566,N_7337,N_6029);
and U7567 (N_7567,N_7472,N_6105);
xnor U7568 (N_7568,N_7139,N_6624);
and U7569 (N_7569,N_6362,N_6375);
xor U7570 (N_7570,N_6293,N_7364);
or U7571 (N_7571,N_6909,N_6127);
nor U7572 (N_7572,N_7141,N_6478);
nand U7573 (N_7573,N_6013,N_7146);
nand U7574 (N_7574,N_6200,N_6077);
nand U7575 (N_7575,N_6739,N_6752);
and U7576 (N_7576,N_6071,N_6968);
and U7577 (N_7577,N_7387,N_6904);
or U7578 (N_7578,N_6444,N_7342);
nand U7579 (N_7579,N_6474,N_6548);
or U7580 (N_7580,N_6611,N_7267);
xor U7581 (N_7581,N_7232,N_6637);
xor U7582 (N_7582,N_6285,N_7099);
or U7583 (N_7583,N_6633,N_6211);
or U7584 (N_7584,N_6250,N_6987);
nor U7585 (N_7585,N_6789,N_6193);
nor U7586 (N_7586,N_6795,N_6757);
nand U7587 (N_7587,N_7429,N_7159);
and U7588 (N_7588,N_7307,N_6157);
nand U7589 (N_7589,N_7190,N_6539);
or U7590 (N_7590,N_7069,N_7378);
or U7591 (N_7591,N_6256,N_6903);
or U7592 (N_7592,N_7303,N_6019);
nor U7593 (N_7593,N_7094,N_6315);
and U7594 (N_7594,N_6585,N_6360);
or U7595 (N_7595,N_6353,N_7494);
nand U7596 (N_7596,N_6581,N_7459);
nand U7597 (N_7597,N_6209,N_6230);
or U7598 (N_7598,N_6065,N_6534);
nor U7599 (N_7599,N_7471,N_6339);
or U7600 (N_7600,N_7255,N_6088);
nand U7601 (N_7601,N_7125,N_7485);
nand U7602 (N_7602,N_6806,N_6988);
nor U7603 (N_7603,N_6544,N_7444);
nand U7604 (N_7604,N_6166,N_7109);
and U7605 (N_7605,N_6686,N_7136);
and U7606 (N_7606,N_6069,N_7225);
and U7607 (N_7607,N_7347,N_6884);
nor U7608 (N_7608,N_6158,N_6199);
or U7609 (N_7609,N_6083,N_7394);
nand U7610 (N_7610,N_6475,N_7432);
nor U7611 (N_7611,N_6094,N_6893);
nand U7612 (N_7612,N_6859,N_6203);
nor U7613 (N_7613,N_6976,N_6269);
nand U7614 (N_7614,N_6823,N_7183);
and U7615 (N_7615,N_6507,N_6306);
nor U7616 (N_7616,N_6164,N_7341);
and U7617 (N_7617,N_6251,N_6247);
or U7618 (N_7618,N_6060,N_7240);
and U7619 (N_7619,N_7124,N_7468);
nor U7620 (N_7620,N_6612,N_7039);
nor U7621 (N_7621,N_6206,N_7016);
nor U7622 (N_7622,N_6395,N_6221);
or U7623 (N_7623,N_6223,N_6731);
or U7624 (N_7624,N_7311,N_6412);
nand U7625 (N_7625,N_7479,N_6798);
or U7626 (N_7626,N_7211,N_7011);
nor U7627 (N_7627,N_7319,N_7499);
nand U7628 (N_7628,N_6383,N_7077);
nor U7629 (N_7629,N_6407,N_6876);
nor U7630 (N_7630,N_6953,N_6602);
nor U7631 (N_7631,N_6990,N_6862);
nor U7632 (N_7632,N_7022,N_6769);
or U7633 (N_7633,N_6120,N_7356);
or U7634 (N_7634,N_7464,N_6411);
nor U7635 (N_7635,N_7244,N_6403);
nor U7636 (N_7636,N_6505,N_6224);
nand U7637 (N_7637,N_6389,N_6593);
nor U7638 (N_7638,N_6442,N_6851);
nand U7639 (N_7639,N_6179,N_6402);
nand U7640 (N_7640,N_7126,N_7493);
nor U7641 (N_7641,N_7300,N_6196);
and U7642 (N_7642,N_6194,N_7480);
xor U7643 (N_7643,N_6826,N_6919);
or U7644 (N_7644,N_7170,N_7172);
nor U7645 (N_7645,N_6342,N_6722);
nand U7646 (N_7646,N_6771,N_7089);
nor U7647 (N_7647,N_6770,N_6217);
nand U7648 (N_7648,N_7229,N_6697);
nor U7649 (N_7649,N_6931,N_7250);
nor U7650 (N_7650,N_6153,N_6322);
or U7651 (N_7651,N_7271,N_7491);
and U7652 (N_7652,N_7334,N_6767);
and U7653 (N_7653,N_6212,N_7030);
xor U7654 (N_7654,N_7379,N_7247);
or U7655 (N_7655,N_6374,N_6737);
nor U7656 (N_7656,N_6218,N_7061);
xnor U7657 (N_7657,N_6554,N_6335);
nand U7658 (N_7658,N_7135,N_6497);
and U7659 (N_7659,N_6744,N_7496);
nor U7660 (N_7660,N_7082,N_7407);
nor U7661 (N_7661,N_6689,N_6489);
nand U7662 (N_7662,N_6388,N_6473);
nor U7663 (N_7663,N_6580,N_6846);
and U7664 (N_7664,N_6009,N_7103);
nor U7665 (N_7665,N_6370,N_6108);
or U7666 (N_7666,N_6479,N_6055);
and U7667 (N_7667,N_6628,N_7425);
nor U7668 (N_7668,N_6645,N_7065);
or U7669 (N_7669,N_7184,N_6503);
and U7670 (N_7670,N_6040,N_6390);
nor U7671 (N_7671,N_6704,N_6541);
and U7672 (N_7672,N_6310,N_7145);
nor U7673 (N_7673,N_6061,N_6857);
and U7674 (N_7674,N_7157,N_7179);
and U7675 (N_7675,N_6254,N_7287);
or U7676 (N_7676,N_6829,N_7401);
or U7677 (N_7677,N_6720,N_6455);
or U7678 (N_7678,N_7147,N_6096);
and U7679 (N_7679,N_6922,N_6141);
and U7680 (N_7680,N_6590,N_6101);
nand U7681 (N_7681,N_6382,N_6132);
nor U7682 (N_7682,N_6261,N_6808);
and U7683 (N_7683,N_6399,N_6928);
or U7684 (N_7684,N_7367,N_6130);
or U7685 (N_7685,N_6449,N_6181);
or U7686 (N_7686,N_6941,N_6097);
xor U7687 (N_7687,N_6810,N_7257);
and U7688 (N_7688,N_6234,N_6677);
or U7689 (N_7689,N_7350,N_7374);
or U7690 (N_7690,N_7292,N_7308);
nor U7691 (N_7691,N_7409,N_6386);
and U7692 (N_7692,N_6352,N_7453);
nor U7693 (N_7693,N_6710,N_7162);
nand U7694 (N_7694,N_6422,N_6281);
and U7695 (N_7695,N_7073,N_6226);
nand U7696 (N_7696,N_7017,N_7115);
nor U7697 (N_7697,N_6465,N_6705);
nor U7698 (N_7698,N_6051,N_6125);
nand U7699 (N_7699,N_7218,N_6781);
or U7700 (N_7700,N_7296,N_6286);
nor U7701 (N_7701,N_7389,N_6186);
nor U7702 (N_7702,N_7284,N_7262);
or U7703 (N_7703,N_7175,N_7092);
xor U7704 (N_7704,N_7490,N_6517);
or U7705 (N_7705,N_6551,N_6197);
and U7706 (N_7706,N_7423,N_6378);
nor U7707 (N_7707,N_7012,N_6368);
and U7708 (N_7708,N_7239,N_6093);
nor U7709 (N_7709,N_6925,N_7302);
nand U7710 (N_7710,N_7353,N_6317);
or U7711 (N_7711,N_7314,N_7028);
or U7712 (N_7712,N_7066,N_7201);
nor U7713 (N_7713,N_7155,N_6266);
nand U7714 (N_7714,N_6324,N_6995);
nand U7715 (N_7715,N_6567,N_6787);
or U7716 (N_7716,N_7117,N_7368);
and U7717 (N_7717,N_6471,N_6530);
xor U7718 (N_7718,N_6434,N_6491);
nor U7719 (N_7719,N_7484,N_6484);
nand U7720 (N_7720,N_6280,N_7304);
or U7721 (N_7721,N_6618,N_6329);
nand U7722 (N_7722,N_6170,N_6560);
or U7723 (N_7723,N_7110,N_6472);
nor U7724 (N_7724,N_6005,N_6713);
xnor U7725 (N_7725,N_6632,N_7273);
nand U7726 (N_7726,N_6668,N_7336);
nor U7727 (N_7727,N_6140,N_6205);
nand U7728 (N_7728,N_7071,N_7053);
and U7729 (N_7729,N_6259,N_6133);
nor U7730 (N_7730,N_7352,N_6948);
or U7731 (N_7731,N_6086,N_6260);
or U7732 (N_7732,N_6579,N_6452);
nand U7733 (N_7733,N_6607,N_6997);
nand U7734 (N_7734,N_7181,N_6684);
and U7735 (N_7735,N_6986,N_7060);
nand U7736 (N_7736,N_6896,N_7046);
nand U7737 (N_7737,N_7116,N_6309);
nor U7738 (N_7738,N_6975,N_6518);
or U7739 (N_7739,N_6372,N_6959);
and U7740 (N_7740,N_6433,N_6850);
nand U7741 (N_7741,N_6592,N_6092);
nand U7742 (N_7742,N_6090,N_7402);
or U7743 (N_7743,N_7068,N_6746);
nand U7744 (N_7744,N_6406,N_6742);
nand U7745 (N_7745,N_7291,N_7264);
nor U7746 (N_7746,N_6337,N_6355);
or U7747 (N_7747,N_6204,N_7121);
nand U7748 (N_7748,N_7180,N_6718);
or U7749 (N_7749,N_6822,N_7037);
and U7750 (N_7750,N_6128,N_7006);
or U7751 (N_7751,N_6198,N_6113);
and U7752 (N_7752,N_7462,N_6707);
nor U7753 (N_7753,N_6082,N_6219);
or U7754 (N_7754,N_7329,N_6774);
and U7755 (N_7755,N_7414,N_6034);
nand U7756 (N_7756,N_6328,N_6877);
or U7757 (N_7757,N_6424,N_7279);
nand U7758 (N_7758,N_7059,N_6991);
nand U7759 (N_7759,N_6287,N_7080);
xnor U7760 (N_7760,N_6498,N_6364);
xnor U7761 (N_7761,N_7004,N_6682);
nor U7762 (N_7762,N_7294,N_6623);
nor U7763 (N_7763,N_6458,N_6715);
nor U7764 (N_7764,N_7400,N_6122);
or U7765 (N_7765,N_6075,N_6002);
nand U7766 (N_7766,N_6553,N_7062);
and U7767 (N_7767,N_6947,N_6110);
or U7768 (N_7768,N_7312,N_7275);
or U7769 (N_7769,N_6320,N_6311);
nand U7770 (N_7770,N_6845,N_7431);
nand U7771 (N_7771,N_6296,N_7152);
nor U7772 (N_7772,N_6070,N_6246);
or U7773 (N_7773,N_6830,N_7122);
or U7774 (N_7774,N_6883,N_6868);
or U7775 (N_7775,N_6818,N_6425);
nor U7776 (N_7776,N_7108,N_7165);
nand U7777 (N_7777,N_7249,N_6703);
nor U7778 (N_7778,N_6811,N_7123);
nand U7779 (N_7779,N_7107,N_6816);
or U7780 (N_7780,N_7370,N_6946);
nand U7781 (N_7781,N_6233,N_6298);
nor U7782 (N_7782,N_6726,N_7321);
and U7783 (N_7783,N_6369,N_7023);
and U7784 (N_7784,N_7160,N_7128);
and U7785 (N_7785,N_6949,N_6300);
or U7786 (N_7786,N_7243,N_7404);
nand U7787 (N_7787,N_6777,N_6817);
nand U7788 (N_7788,N_7150,N_7032);
and U7789 (N_7789,N_6741,N_7487);
nand U7790 (N_7790,N_6880,N_6546);
nand U7791 (N_7791,N_6867,N_7057);
and U7792 (N_7792,N_6938,N_7388);
nor U7793 (N_7793,N_6629,N_6923);
and U7794 (N_7794,N_7119,N_6522);
nand U7795 (N_7795,N_6634,N_7241);
nor U7796 (N_7796,N_6640,N_7095);
or U7797 (N_7797,N_6238,N_7140);
nor U7798 (N_7798,N_7021,N_6118);
nand U7799 (N_7799,N_6169,N_7408);
or U7800 (N_7800,N_7441,N_7392);
or U7801 (N_7801,N_6468,N_7083);
or U7802 (N_7802,N_7272,N_6410);
or U7803 (N_7803,N_6102,N_6314);
nor U7804 (N_7804,N_7452,N_6049);
or U7805 (N_7805,N_6954,N_7256);
or U7806 (N_7806,N_7274,N_6012);
or U7807 (N_7807,N_7443,N_6911);
and U7808 (N_7808,N_6676,N_6316);
or U7809 (N_7809,N_7498,N_6080);
xor U7810 (N_7810,N_6493,N_6937);
nand U7811 (N_7811,N_7209,N_6807);
nand U7812 (N_7812,N_6340,N_6227);
and U7813 (N_7813,N_6147,N_6992);
nand U7814 (N_7814,N_7365,N_6568);
nor U7815 (N_7815,N_6323,N_6920);
or U7816 (N_7816,N_7169,N_7290);
nand U7817 (N_7817,N_7034,N_6466);
nand U7818 (N_7818,N_7282,N_6043);
nor U7819 (N_7819,N_6371,N_6150);
or U7820 (N_7820,N_6932,N_6902);
xnor U7821 (N_7821,N_6780,N_7221);
nand U7822 (N_7822,N_6485,N_6036);
and U7823 (N_7823,N_7224,N_6755);
nor U7824 (N_7824,N_6330,N_6584);
or U7825 (N_7825,N_6439,N_6214);
xnor U7826 (N_7826,N_6708,N_6839);
and U7827 (N_7827,N_7091,N_6143);
and U7828 (N_7828,N_6732,N_6492);
or U7829 (N_7829,N_7127,N_6679);
or U7830 (N_7830,N_7219,N_6486);
nand U7831 (N_7831,N_6301,N_6848);
and U7832 (N_7832,N_6066,N_6004);
or U7833 (N_7833,N_6516,N_6814);
or U7834 (N_7834,N_7102,N_7488);
xor U7835 (N_7835,N_6619,N_7258);
or U7836 (N_7836,N_6343,N_6588);
nand U7837 (N_7837,N_6344,N_7164);
or U7838 (N_7838,N_6985,N_6973);
xnor U7839 (N_7839,N_7481,N_6702);
nand U7840 (N_7840,N_7316,N_6898);
nor U7841 (N_7841,N_6873,N_7455);
and U7842 (N_7842,N_6756,N_6574);
nor U7843 (N_7843,N_6258,N_6161);
nor U7844 (N_7844,N_6834,N_7202);
or U7845 (N_7845,N_7167,N_6562);
nor U7846 (N_7846,N_6794,N_6144);
nand U7847 (N_7847,N_7072,N_6762);
xor U7848 (N_7848,N_6044,N_6304);
or U7849 (N_7849,N_6586,N_6532);
nor U7850 (N_7850,N_6313,N_6667);
and U7851 (N_7851,N_7438,N_6786);
nand U7852 (N_7852,N_6295,N_6481);
nor U7853 (N_7853,N_6201,N_6297);
nor U7854 (N_7854,N_6361,N_6124);
nor U7855 (N_7855,N_6837,N_6496);
nor U7856 (N_7856,N_6334,N_7349);
and U7857 (N_7857,N_6114,N_6605);
nand U7858 (N_7858,N_7385,N_6126);
xor U7859 (N_7859,N_6289,N_6035);
nand U7860 (N_7860,N_6957,N_6979);
and U7861 (N_7861,N_6683,N_7014);
and U7862 (N_7862,N_7405,N_6016);
nand U7863 (N_7863,N_6426,N_7354);
nor U7864 (N_7864,N_6885,N_7440);
nor U7865 (N_7865,N_7058,N_6319);
nor U7866 (N_7866,N_6501,N_7376);
or U7867 (N_7867,N_6620,N_7463);
or U7868 (N_7868,N_6136,N_6006);
nand U7869 (N_7869,N_6681,N_7465);
and U7870 (N_7870,N_6725,N_6828);
nand U7871 (N_7871,N_6241,N_7433);
nor U7872 (N_7872,N_6067,N_6970);
xor U7873 (N_7873,N_7174,N_7231);
or U7874 (N_7874,N_7313,N_6052);
or U7875 (N_7875,N_6601,N_7278);
nand U7876 (N_7876,N_7087,N_6860);
and U7877 (N_7877,N_6457,N_6772);
xor U7878 (N_7878,N_6139,N_6026);
nand U7879 (N_7879,N_6358,N_7420);
or U7880 (N_7880,N_7040,N_6913);
or U7881 (N_7881,N_7000,N_7436);
nor U7882 (N_7882,N_6943,N_7154);
nand U7883 (N_7883,N_7434,N_6847);
nor U7884 (N_7884,N_6914,N_6994);
or U7885 (N_7885,N_6572,N_6950);
and U7886 (N_7886,N_6597,N_6576);
or U7887 (N_7887,N_6190,N_7447);
nand U7888 (N_7888,N_6341,N_6533);
and U7889 (N_7889,N_6087,N_6010);
or U7890 (N_7890,N_7216,N_6239);
and U7891 (N_7891,N_7358,N_6663);
and U7892 (N_7892,N_6504,N_7002);
nand U7893 (N_7893,N_6400,N_7277);
xor U7894 (N_7894,N_7204,N_6962);
nand U7895 (N_7895,N_6173,N_6793);
nor U7896 (N_7896,N_6175,N_7360);
and U7897 (N_7897,N_7086,N_6542);
xor U7898 (N_7898,N_6813,N_6115);
nor U7899 (N_7899,N_6709,N_6490);
nand U7900 (N_7900,N_6187,N_6603);
and U7901 (N_7901,N_6998,N_6796);
xor U7902 (N_7902,N_7085,N_6268);
nor U7903 (N_7903,N_6738,N_7330);
xor U7904 (N_7904,N_6745,N_6208);
nand U7905 (N_7905,N_6644,N_6299);
nor U7906 (N_7906,N_7192,N_6030);
nor U7907 (N_7907,N_7220,N_6294);
nand U7908 (N_7908,N_6236,N_6665);
or U7909 (N_7909,N_6336,N_6537);
or U7910 (N_7910,N_7373,N_6418);
and U7911 (N_7911,N_6930,N_7134);
nor U7912 (N_7912,N_6917,N_6000);
or U7913 (N_7913,N_7486,N_6167);
nor U7914 (N_7914,N_6747,N_6754);
and U7915 (N_7915,N_6753,N_6841);
or U7916 (N_7916,N_7270,N_6751);
or U7917 (N_7917,N_6955,N_6680);
xnor U7918 (N_7918,N_6523,N_7417);
and U7919 (N_7919,N_6833,N_6971);
or U7920 (N_7920,N_6480,N_7114);
nand U7921 (N_7921,N_6587,N_6515);
and U7922 (N_7922,N_6984,N_6111);
or U7923 (N_7923,N_6900,N_6940);
and U7924 (N_7924,N_6427,N_6307);
xnor U7925 (N_7925,N_6235,N_6748);
and U7926 (N_7926,N_7297,N_7029);
nand U7927 (N_7927,N_6561,N_6706);
nand U7928 (N_7928,N_6391,N_7390);
nand U7929 (N_7929,N_6081,N_7309);
nand U7930 (N_7930,N_6393,N_6782);
and U7931 (N_7931,N_7031,N_7327);
or U7932 (N_7932,N_6275,N_6454);
nor U7933 (N_7933,N_7415,N_6116);
nand U7934 (N_7934,N_7081,N_6695);
and U7935 (N_7935,N_6563,N_6448);
or U7936 (N_7936,N_6151,N_6536);
or U7937 (N_7937,N_7288,N_6556);
or U7938 (N_7938,N_6263,N_6356);
and U7939 (N_7939,N_6951,N_6895);
xor U7940 (N_7940,N_6963,N_7371);
nand U7941 (N_7941,N_6423,N_6785);
nor U7942 (N_7942,N_6073,N_6416);
and U7943 (N_7943,N_7158,N_6685);
xor U7944 (N_7944,N_6543,N_6119);
or U7945 (N_7945,N_6346,N_6146);
nand U7946 (N_7946,N_6499,N_7033);
nand U7947 (N_7947,N_7163,N_7186);
nor U7948 (N_7948,N_6625,N_7227);
nand U7949 (N_7949,N_7133,N_6662);
and U7950 (N_7950,N_6156,N_6797);
xnor U7951 (N_7951,N_6283,N_6621);
or U7952 (N_7952,N_7338,N_7144);
and U7953 (N_7953,N_6249,N_6445);
nand U7954 (N_7954,N_6723,N_7369);
nor U7955 (N_7955,N_7377,N_6609);
nand U7956 (N_7956,N_6017,N_6651);
nor U7957 (N_7957,N_6596,N_7252);
xor U7958 (N_7958,N_7153,N_7345);
nand U7959 (N_7959,N_6521,N_7084);
or U7960 (N_7960,N_6047,N_7188);
xnor U7961 (N_7961,N_6840,N_7478);
xnor U7962 (N_7962,N_7254,N_6104);
nand U7963 (N_7963,N_6582,N_6821);
or U7964 (N_7964,N_7010,N_6719);
and U7965 (N_7965,N_7467,N_7412);
or U7966 (N_7966,N_6265,N_7009);
and U7967 (N_7967,N_7280,N_7090);
nor U7968 (N_7968,N_6024,N_6229);
and U7969 (N_7969,N_6408,N_6892);
and U7970 (N_7970,N_6776,N_6469);
or U7971 (N_7971,N_7212,N_6519);
nor U7972 (N_7972,N_6791,N_7331);
nor U7973 (N_7973,N_6549,N_6025);
xor U7974 (N_7974,N_6699,N_7129);
xnor U7975 (N_7975,N_7149,N_6693);
nand U7976 (N_7976,N_6961,N_6129);
and U7977 (N_7977,N_6435,N_6354);
and U7978 (N_7978,N_6357,N_7366);
or U7979 (N_7979,N_6788,N_6244);
and U7980 (N_7980,N_7283,N_7355);
nand U7981 (N_7981,N_7098,N_7251);
nor U7982 (N_7982,N_6367,N_6267);
xnor U7983 (N_7983,N_6401,N_6509);
or U7984 (N_7984,N_6091,N_7096);
xor U7985 (N_7985,N_6936,N_7315);
nor U7986 (N_7986,N_6461,N_6216);
xnor U7987 (N_7987,N_6253,N_6655);
and U7988 (N_7988,N_6736,N_7375);
xnor U7989 (N_7989,N_6694,N_6773);
and U7990 (N_7990,N_7199,N_7048);
nand U7991 (N_7991,N_7266,N_6057);
xnor U7992 (N_7992,N_7005,N_7450);
nand U7993 (N_7993,N_6185,N_6222);
xnor U7994 (N_7994,N_6366,N_7469);
nand U7995 (N_7995,N_7489,N_6886);
or U7996 (N_7996,N_7185,N_6459);
and U7997 (N_7997,N_7222,N_7476);
and U7998 (N_7998,N_6392,N_6397);
nand U7999 (N_7999,N_7197,N_7448);
and U8000 (N_8000,N_6616,N_6441);
and U8001 (N_8001,N_7344,N_6566);
or U8002 (N_8002,N_6456,N_6500);
xor U8003 (N_8003,N_6058,N_6759);
nand U8004 (N_8004,N_6277,N_6790);
and U8005 (N_8005,N_7064,N_6802);
and U8006 (N_8006,N_6871,N_7120);
nor U8007 (N_8007,N_6008,N_6431);
or U8008 (N_8008,N_6617,N_6042);
or U8009 (N_8009,N_6451,N_6318);
xor U8010 (N_8010,N_6384,N_6347);
xnor U8011 (N_8011,N_6023,N_6727);
or U8012 (N_8012,N_6076,N_6189);
xor U8013 (N_8013,N_7020,N_7189);
or U8014 (N_8014,N_6557,N_7248);
nor U8015 (N_8015,N_6978,N_6123);
nor U8016 (N_8016,N_6656,N_6606);
and U8017 (N_8017,N_6373,N_7426);
or U8018 (N_8018,N_6278,N_7215);
nor U8019 (N_8019,N_7112,N_7466);
nor U8020 (N_8020,N_6714,N_7276);
or U8021 (N_8021,N_6112,N_7346);
and U8022 (N_8022,N_6809,N_6046);
nand U8023 (N_8023,N_6591,N_6326);
and U8024 (N_8024,N_6934,N_7442);
xor U8025 (N_8025,N_6749,N_7395);
nand U8026 (N_8026,N_6376,N_6856);
nand U8027 (N_8027,N_6916,N_6514);
nor U8028 (N_8028,N_7234,N_7446);
nor U8029 (N_8029,N_7026,N_6661);
or U8030 (N_8030,N_7317,N_6428);
nand U8031 (N_8031,N_6559,N_7260);
or U8032 (N_8032,N_7195,N_6470);
nand U8033 (N_8033,N_6415,N_6547);
or U8034 (N_8034,N_6700,N_7397);
xor U8035 (N_8035,N_6062,N_6865);
or U8036 (N_8036,N_6430,N_6910);
nor U8037 (N_8037,N_6599,N_7318);
or U8038 (N_8038,N_6279,N_6405);
nor U8039 (N_8039,N_6569,N_6870);
nor U8040 (N_8040,N_6899,N_6453);
nor U8041 (N_8041,N_6944,N_6958);
and U8042 (N_8042,N_7439,N_7079);
nand U8043 (N_8043,N_6972,N_6508);
and U8044 (N_8044,N_7391,N_6996);
nand U8045 (N_8045,N_6312,N_6476);
and U8046 (N_8046,N_7422,N_6163);
nor U8047 (N_8047,N_6882,N_7381);
and U8048 (N_8048,N_7497,N_6155);
or U8049 (N_8049,N_7137,N_6824);
nor U8050 (N_8050,N_6648,N_6168);
nor U8051 (N_8051,N_6184,N_7424);
nand U8052 (N_8052,N_6849,N_6220);
or U8053 (N_8053,N_6879,N_7173);
and U8054 (N_8054,N_6843,N_6929);
nand U8055 (N_8055,N_6615,N_6853);
or U8056 (N_8056,N_7332,N_6555);
nor U8057 (N_8057,N_6933,N_6274);
nor U8058 (N_8058,N_7130,N_7238);
or U8059 (N_8059,N_6564,N_6172);
nor U8060 (N_8060,N_6982,N_6825);
or U8061 (N_8061,N_6072,N_6037);
nand U8062 (N_8062,N_6084,N_7044);
nor U8063 (N_8063,N_6812,N_6510);
xor U8064 (N_8064,N_7118,N_6657);
and U8065 (N_8065,N_6135,N_7233);
and U8066 (N_8066,N_7306,N_7289);
or U8067 (N_8067,N_7335,N_6803);
and U8068 (N_8068,N_6359,N_7399);
nor U8069 (N_8069,N_6467,N_6039);
or U8070 (N_8070,N_7324,N_6890);
nor U8071 (N_8071,N_6763,N_6038);
nor U8072 (N_8072,N_6610,N_6460);
nor U8073 (N_8073,N_7482,N_7176);
xnor U8074 (N_8074,N_6117,N_6573);
xor U8075 (N_8075,N_7113,N_6387);
nor U8076 (N_8076,N_7097,N_6192);
nand U8077 (N_8077,N_6981,N_6815);
nand U8078 (N_8078,N_7036,N_6302);
nand U8079 (N_8079,N_6740,N_7326);
and U8080 (N_8080,N_6688,N_7380);
and U8081 (N_8081,N_6905,N_7228);
or U8082 (N_8082,N_7253,N_7049);
xor U8083 (N_8083,N_7298,N_6011);
and U8084 (N_8084,N_6176,N_6728);
nand U8085 (N_8085,N_7340,N_7131);
or U8086 (N_8086,N_6716,N_6183);
and U8087 (N_8087,N_6483,N_6419);
nand U8088 (N_8088,N_6272,N_6696);
nand U8089 (N_8089,N_6032,N_7269);
and U8090 (N_8090,N_6191,N_6014);
nor U8091 (N_8091,N_6854,N_6918);
and U8092 (N_8092,N_7207,N_6641);
nand U8093 (N_8093,N_6734,N_7470);
nand U8094 (N_8094,N_7348,N_7419);
nor U8095 (N_8095,N_6652,N_6784);
nor U8096 (N_8096,N_7206,N_6675);
or U8097 (N_8097,N_7461,N_6015);
xnor U8098 (N_8098,N_6820,N_7398);
nor U8099 (N_8099,N_6659,N_7078);
nand U8100 (N_8100,N_6290,N_6321);
and U8101 (N_8101,N_7435,N_7143);
nand U8102 (N_8102,N_6437,N_6207);
and U8103 (N_8103,N_6231,N_6160);
and U8104 (N_8104,N_6552,N_6965);
nand U8105 (N_8105,N_6255,N_6443);
nand U8106 (N_8106,N_6712,N_6074);
nand U8107 (N_8107,N_6613,N_6888);
and U8108 (N_8108,N_7001,N_6063);
or U8109 (N_8109,N_6570,N_7421);
or U8110 (N_8110,N_7245,N_7043);
nand U8111 (N_8111,N_6717,N_6897);
or U8112 (N_8112,N_7142,N_6213);
nor U8113 (N_8113,N_6131,N_6099);
or U8114 (N_8114,N_7343,N_6054);
nor U8115 (N_8115,N_6477,N_7427);
xor U8116 (N_8116,N_6513,N_6526);
and U8117 (N_8117,N_6658,N_6801);
and U8118 (N_8118,N_6171,N_7106);
or U8119 (N_8119,N_6142,N_7223);
and U8120 (N_8120,N_6438,N_6874);
or U8121 (N_8121,N_7194,N_6003);
or U8122 (N_8122,N_6257,N_7483);
nand U8123 (N_8123,N_6724,N_7035);
or U8124 (N_8124,N_6033,N_6506);
nor U8125 (N_8125,N_6805,N_7196);
or U8126 (N_8126,N_6538,N_6983);
or U8127 (N_8127,N_7416,N_6308);
or U8128 (N_8128,N_6098,N_7074);
nand U8129 (N_8129,N_6494,N_6145);
or U8130 (N_8130,N_6365,N_6558);
or U8131 (N_8131,N_7449,N_6832);
and U8132 (N_8132,N_6348,N_6377);
xor U8133 (N_8133,N_7177,N_6698);
nand U8134 (N_8134,N_6927,N_6974);
xor U8135 (N_8135,N_6237,N_7070);
or U8136 (N_8136,N_7383,N_6945);
or U8137 (N_8137,N_7295,N_6284);
or U8138 (N_8138,N_6385,N_6050);
or U8139 (N_8139,N_6664,N_7339);
xor U8140 (N_8140,N_7363,N_6872);
and U8141 (N_8141,N_6571,N_6993);
nor U8142 (N_8142,N_7208,N_6758);
or U8143 (N_8143,N_6350,N_7495);
or U8144 (N_8144,N_6673,N_6095);
and U8145 (N_8145,N_6969,N_7242);
nand U8146 (N_8146,N_7477,N_6404);
and U8147 (N_8147,N_7007,N_6398);
and U8148 (N_8148,N_7246,N_6089);
xor U8149 (N_8149,N_7008,N_6906);
xor U8150 (N_8150,N_6059,N_6420);
nand U8151 (N_8151,N_7178,N_6159);
or U8152 (N_8152,N_6512,N_6654);
nand U8153 (N_8153,N_7063,N_6440);
nand U8154 (N_8154,N_6670,N_6529);
and U8155 (N_8155,N_7310,N_6647);
and U8156 (N_8156,N_6638,N_6165);
nand U8157 (N_8157,N_7382,N_6018);
and U8158 (N_8158,N_6079,N_7475);
nand U8159 (N_8159,N_6669,N_6690);
xnor U8160 (N_8160,N_6852,N_6577);
nand U8161 (N_8161,N_6178,N_7351);
xnor U8162 (N_8162,N_6134,N_6907);
nor U8163 (N_8163,N_6188,N_7418);
and U8164 (N_8164,N_6535,N_6643);
nor U8165 (N_8165,N_7101,N_7286);
nor U8166 (N_8166,N_6804,N_7193);
nor U8167 (N_8167,N_6653,N_6414);
nor U8168 (N_8168,N_6031,N_6264);
nand U8169 (N_8169,N_7460,N_6550);
or U8170 (N_8170,N_6041,N_7015);
and U8171 (N_8171,N_6276,N_6351);
or U8172 (N_8172,N_6887,N_6531);
or U8173 (N_8173,N_6956,N_6100);
xor U8174 (N_8174,N_6660,N_7372);
or U8175 (N_8175,N_6429,N_6889);
and U8176 (N_8176,N_6598,N_7458);
and U8177 (N_8177,N_6594,N_7041);
nor U8178 (N_8178,N_7261,N_7213);
xor U8179 (N_8179,N_6225,N_6575);
xor U8180 (N_8180,N_7050,N_6908);
or U8181 (N_8181,N_7457,N_7132);
and U8182 (N_8182,N_7411,N_6149);
nor U8183 (N_8183,N_6980,N_6836);
or U8184 (N_8184,N_6446,N_6864);
nor U8185 (N_8185,N_6672,N_6524);
and U8186 (N_8186,N_7305,N_6766);
nand U8187 (N_8187,N_6614,N_6520);
or U8188 (N_8188,N_6305,N_6381);
or U8189 (N_8189,N_6332,N_6819);
nor U8190 (N_8190,N_6303,N_6349);
or U8191 (N_8191,N_7237,N_7230);
and U8192 (N_8192,N_6650,N_6894);
nor U8193 (N_8193,N_6783,N_6488);
and U8194 (N_8194,N_6589,N_6926);
or U8195 (N_8195,N_6921,N_6827);
or U8196 (N_8196,N_7451,N_7357);
xor U8197 (N_8197,N_7492,N_6858);
or U8198 (N_8198,N_6152,N_6463);
nor U8199 (N_8199,N_6608,N_7285);
or U8200 (N_8200,N_7263,N_6799);
nand U8201 (N_8201,N_6636,N_6775);
nand U8202 (N_8202,N_7320,N_7138);
and U8203 (N_8203,N_7191,N_6924);
nand U8204 (N_8204,N_6626,N_7198);
and U8205 (N_8205,N_7055,N_6631);
and U8206 (N_8206,N_7226,N_6666);
and U8207 (N_8207,N_7393,N_6687);
nor U8208 (N_8208,N_6270,N_6495);
nor U8209 (N_8209,N_6502,N_6045);
nor U8210 (N_8210,N_6701,N_6869);
nand U8211 (N_8211,N_6180,N_6195);
nand U8212 (N_8212,N_6964,N_6743);
and U8213 (N_8213,N_6154,N_7187);
or U8214 (N_8214,N_6394,N_7200);
nand U8215 (N_8215,N_7281,N_6338);
xor U8216 (N_8216,N_7384,N_6109);
and U8217 (N_8217,N_7430,N_6635);
nor U8218 (N_8218,N_6639,N_6462);
nor U8219 (N_8219,N_6085,N_6967);
or U8220 (N_8220,N_7076,N_6765);
or U8221 (N_8221,N_6692,N_7075);
nand U8222 (N_8222,N_6901,N_7217);
nor U8223 (N_8223,N_6447,N_7293);
nor U8224 (N_8224,N_7161,N_6243);
nor U8225 (N_8225,N_6271,N_7361);
nand U8226 (N_8226,N_6464,N_7151);
or U8227 (N_8227,N_6711,N_6528);
nand U8228 (N_8228,N_6768,N_6861);
and U8229 (N_8229,N_7403,N_6182);
nand U8230 (N_8230,N_7428,N_7088);
or U8231 (N_8231,N_7100,N_7322);
nor U8232 (N_8232,N_6202,N_6421);
or U8233 (N_8233,N_6545,N_6106);
nor U8234 (N_8234,N_6527,N_6107);
nor U8235 (N_8235,N_7051,N_6007);
nand U8236 (N_8236,N_6952,N_7104);
and U8237 (N_8237,N_6630,N_7456);
or U8238 (N_8238,N_6844,N_6750);
and U8239 (N_8239,N_6331,N_6292);
xor U8240 (N_8240,N_6056,N_6001);
and U8241 (N_8241,N_6288,N_7236);
or U8242 (N_8242,N_6436,N_7027);
nor U8243 (N_8243,N_7386,N_6977);
or U8244 (N_8244,N_6960,N_6021);
nor U8245 (N_8245,N_7166,N_6831);
nor U8246 (N_8246,N_6078,N_7111);
nand U8247 (N_8247,N_7328,N_6053);
nor U8248 (N_8248,N_6242,N_7323);
or U8249 (N_8249,N_6691,N_7259);
and U8250 (N_8250,N_7353,N_6974);
or U8251 (N_8251,N_6562,N_7338);
and U8252 (N_8252,N_6410,N_7428);
and U8253 (N_8253,N_6736,N_7268);
and U8254 (N_8254,N_7225,N_6065);
and U8255 (N_8255,N_6867,N_6259);
and U8256 (N_8256,N_6604,N_6710);
and U8257 (N_8257,N_7481,N_6272);
nor U8258 (N_8258,N_6344,N_6818);
nor U8259 (N_8259,N_6910,N_6275);
xnor U8260 (N_8260,N_7476,N_7352);
xor U8261 (N_8261,N_7449,N_6379);
or U8262 (N_8262,N_6643,N_7276);
or U8263 (N_8263,N_6367,N_7199);
nor U8264 (N_8264,N_6527,N_6748);
nor U8265 (N_8265,N_6327,N_6758);
nand U8266 (N_8266,N_6054,N_7403);
or U8267 (N_8267,N_7142,N_6845);
and U8268 (N_8268,N_6268,N_7347);
nor U8269 (N_8269,N_6196,N_7279);
xor U8270 (N_8270,N_6769,N_6909);
nand U8271 (N_8271,N_6532,N_6942);
and U8272 (N_8272,N_6960,N_6784);
nor U8273 (N_8273,N_6453,N_6411);
nand U8274 (N_8274,N_6130,N_6018);
and U8275 (N_8275,N_6312,N_7422);
nor U8276 (N_8276,N_6929,N_6986);
and U8277 (N_8277,N_6056,N_7096);
nor U8278 (N_8278,N_6565,N_6459);
nor U8279 (N_8279,N_6817,N_7438);
xnor U8280 (N_8280,N_6828,N_6635);
nand U8281 (N_8281,N_6841,N_6396);
nand U8282 (N_8282,N_6061,N_6178);
xnor U8283 (N_8283,N_6793,N_6854);
nor U8284 (N_8284,N_6226,N_6102);
nor U8285 (N_8285,N_6497,N_7219);
or U8286 (N_8286,N_6705,N_7172);
and U8287 (N_8287,N_6430,N_7431);
nand U8288 (N_8288,N_6497,N_6318);
or U8289 (N_8289,N_6712,N_6579);
or U8290 (N_8290,N_7127,N_6231);
xnor U8291 (N_8291,N_6905,N_7402);
nor U8292 (N_8292,N_6432,N_6522);
nand U8293 (N_8293,N_7016,N_6886);
nand U8294 (N_8294,N_6086,N_6189);
or U8295 (N_8295,N_6106,N_6945);
nand U8296 (N_8296,N_6345,N_7342);
or U8297 (N_8297,N_7193,N_7481);
or U8298 (N_8298,N_7364,N_6706);
nor U8299 (N_8299,N_6309,N_7041);
nand U8300 (N_8300,N_7060,N_7011);
nor U8301 (N_8301,N_6501,N_6649);
and U8302 (N_8302,N_6060,N_6654);
or U8303 (N_8303,N_7084,N_7454);
xnor U8304 (N_8304,N_6341,N_6680);
and U8305 (N_8305,N_6186,N_7253);
or U8306 (N_8306,N_6075,N_6115);
nand U8307 (N_8307,N_7337,N_6568);
nand U8308 (N_8308,N_6577,N_6824);
nor U8309 (N_8309,N_7120,N_7366);
and U8310 (N_8310,N_6945,N_7497);
nand U8311 (N_8311,N_6342,N_6404);
and U8312 (N_8312,N_6934,N_6521);
nand U8313 (N_8313,N_6213,N_6179);
and U8314 (N_8314,N_6618,N_6553);
nor U8315 (N_8315,N_6842,N_7283);
or U8316 (N_8316,N_7047,N_6470);
or U8317 (N_8317,N_6512,N_7024);
nor U8318 (N_8318,N_6597,N_6345);
or U8319 (N_8319,N_7112,N_7050);
or U8320 (N_8320,N_7482,N_6967);
or U8321 (N_8321,N_7063,N_6363);
and U8322 (N_8322,N_6414,N_6255);
nand U8323 (N_8323,N_7106,N_6872);
nor U8324 (N_8324,N_7221,N_6094);
nor U8325 (N_8325,N_6681,N_6346);
nand U8326 (N_8326,N_7170,N_7405);
or U8327 (N_8327,N_6324,N_6052);
nand U8328 (N_8328,N_6317,N_6928);
nor U8329 (N_8329,N_6097,N_6641);
nand U8330 (N_8330,N_7014,N_6695);
nor U8331 (N_8331,N_6825,N_6469);
nand U8332 (N_8332,N_7389,N_6916);
nand U8333 (N_8333,N_6800,N_6161);
nand U8334 (N_8334,N_6816,N_6581);
nor U8335 (N_8335,N_7243,N_6987);
nor U8336 (N_8336,N_6561,N_6660);
nor U8337 (N_8337,N_6324,N_7428);
or U8338 (N_8338,N_6064,N_6768);
nand U8339 (N_8339,N_6166,N_7097);
xor U8340 (N_8340,N_6748,N_7037);
or U8341 (N_8341,N_6368,N_7085);
or U8342 (N_8342,N_6593,N_7077);
or U8343 (N_8343,N_6558,N_7068);
nor U8344 (N_8344,N_6292,N_6655);
nand U8345 (N_8345,N_7444,N_6856);
nand U8346 (N_8346,N_6897,N_6507);
nand U8347 (N_8347,N_7200,N_6751);
nand U8348 (N_8348,N_6212,N_7227);
xor U8349 (N_8349,N_7316,N_6630);
nand U8350 (N_8350,N_7119,N_6632);
nor U8351 (N_8351,N_6305,N_6346);
nor U8352 (N_8352,N_6239,N_7198);
nor U8353 (N_8353,N_6134,N_7453);
and U8354 (N_8354,N_6844,N_6114);
nand U8355 (N_8355,N_7448,N_6093);
and U8356 (N_8356,N_6068,N_6541);
or U8357 (N_8357,N_7415,N_6809);
nand U8358 (N_8358,N_7032,N_6587);
nor U8359 (N_8359,N_7447,N_6360);
nor U8360 (N_8360,N_6661,N_6277);
nand U8361 (N_8361,N_6584,N_6431);
nor U8362 (N_8362,N_6864,N_7416);
nand U8363 (N_8363,N_6766,N_7465);
nand U8364 (N_8364,N_6424,N_6386);
xor U8365 (N_8365,N_7282,N_6315);
or U8366 (N_8366,N_6700,N_7289);
nor U8367 (N_8367,N_6231,N_6537);
xnor U8368 (N_8368,N_7439,N_7068);
or U8369 (N_8369,N_6816,N_6781);
and U8370 (N_8370,N_6998,N_7419);
nor U8371 (N_8371,N_7000,N_7339);
or U8372 (N_8372,N_6673,N_6713);
nor U8373 (N_8373,N_6349,N_6535);
xor U8374 (N_8374,N_7029,N_6592);
and U8375 (N_8375,N_6066,N_6851);
and U8376 (N_8376,N_7283,N_7301);
nor U8377 (N_8377,N_6784,N_6791);
nor U8378 (N_8378,N_6198,N_6279);
nand U8379 (N_8379,N_6087,N_7322);
nor U8380 (N_8380,N_7233,N_6375);
or U8381 (N_8381,N_6377,N_6762);
or U8382 (N_8382,N_6713,N_6083);
nand U8383 (N_8383,N_6557,N_7092);
or U8384 (N_8384,N_6512,N_7412);
nand U8385 (N_8385,N_6061,N_7458);
and U8386 (N_8386,N_7350,N_7064);
or U8387 (N_8387,N_7408,N_6306);
nor U8388 (N_8388,N_7037,N_6104);
nor U8389 (N_8389,N_6915,N_7073);
or U8390 (N_8390,N_6179,N_6286);
nor U8391 (N_8391,N_6354,N_6083);
or U8392 (N_8392,N_7455,N_7279);
and U8393 (N_8393,N_7303,N_6652);
xor U8394 (N_8394,N_6410,N_7435);
nor U8395 (N_8395,N_6900,N_7012);
nor U8396 (N_8396,N_6778,N_6635);
nand U8397 (N_8397,N_6284,N_6679);
nor U8398 (N_8398,N_6723,N_6940);
or U8399 (N_8399,N_6081,N_7477);
or U8400 (N_8400,N_6780,N_6449);
and U8401 (N_8401,N_7213,N_7220);
or U8402 (N_8402,N_6868,N_7272);
or U8403 (N_8403,N_7160,N_6200);
or U8404 (N_8404,N_6977,N_6941);
or U8405 (N_8405,N_6095,N_7406);
nand U8406 (N_8406,N_6066,N_6164);
or U8407 (N_8407,N_6441,N_6993);
nand U8408 (N_8408,N_7029,N_6395);
or U8409 (N_8409,N_6110,N_6786);
xor U8410 (N_8410,N_6818,N_6851);
or U8411 (N_8411,N_6452,N_6978);
nor U8412 (N_8412,N_6532,N_6736);
nor U8413 (N_8413,N_6678,N_6674);
or U8414 (N_8414,N_6871,N_7025);
nor U8415 (N_8415,N_7390,N_6662);
and U8416 (N_8416,N_7088,N_6023);
or U8417 (N_8417,N_7275,N_7149);
and U8418 (N_8418,N_6148,N_6756);
nor U8419 (N_8419,N_6824,N_6755);
or U8420 (N_8420,N_6916,N_6006);
or U8421 (N_8421,N_7349,N_7478);
xor U8422 (N_8422,N_7119,N_6800);
and U8423 (N_8423,N_6435,N_6494);
nor U8424 (N_8424,N_6765,N_7269);
or U8425 (N_8425,N_6807,N_6750);
or U8426 (N_8426,N_6082,N_6970);
and U8427 (N_8427,N_6010,N_7440);
nand U8428 (N_8428,N_7299,N_6244);
and U8429 (N_8429,N_7256,N_6036);
or U8430 (N_8430,N_6094,N_6187);
nand U8431 (N_8431,N_6976,N_6958);
nor U8432 (N_8432,N_7467,N_7146);
nor U8433 (N_8433,N_7268,N_6524);
and U8434 (N_8434,N_6459,N_6508);
xnor U8435 (N_8435,N_6125,N_6560);
xnor U8436 (N_8436,N_6492,N_6048);
and U8437 (N_8437,N_7013,N_6356);
nor U8438 (N_8438,N_6281,N_7112);
nor U8439 (N_8439,N_6533,N_6045);
or U8440 (N_8440,N_6869,N_6079);
or U8441 (N_8441,N_6473,N_6619);
nand U8442 (N_8442,N_6020,N_6894);
nand U8443 (N_8443,N_6555,N_6949);
nand U8444 (N_8444,N_7002,N_6261);
and U8445 (N_8445,N_6595,N_7023);
and U8446 (N_8446,N_7004,N_6277);
and U8447 (N_8447,N_7320,N_6932);
xnor U8448 (N_8448,N_7443,N_6704);
and U8449 (N_8449,N_6636,N_6602);
or U8450 (N_8450,N_7038,N_6900);
nor U8451 (N_8451,N_6102,N_7432);
nor U8452 (N_8452,N_6033,N_6835);
nand U8453 (N_8453,N_7443,N_7065);
nand U8454 (N_8454,N_6811,N_6665);
nand U8455 (N_8455,N_7225,N_6441);
nor U8456 (N_8456,N_6164,N_6505);
nor U8457 (N_8457,N_6459,N_7446);
nor U8458 (N_8458,N_7377,N_6076);
nor U8459 (N_8459,N_7206,N_6203);
nor U8460 (N_8460,N_7293,N_6850);
nor U8461 (N_8461,N_7015,N_6609);
or U8462 (N_8462,N_6274,N_6149);
nand U8463 (N_8463,N_6084,N_7118);
nand U8464 (N_8464,N_6636,N_6599);
or U8465 (N_8465,N_6016,N_7268);
nor U8466 (N_8466,N_6019,N_7236);
xor U8467 (N_8467,N_6538,N_6171);
nand U8468 (N_8468,N_6924,N_7174);
nand U8469 (N_8469,N_7202,N_6125);
or U8470 (N_8470,N_7497,N_6652);
or U8471 (N_8471,N_6104,N_6730);
nand U8472 (N_8472,N_7281,N_6252);
nor U8473 (N_8473,N_7378,N_6706);
nand U8474 (N_8474,N_7061,N_6331);
nor U8475 (N_8475,N_7039,N_6478);
nand U8476 (N_8476,N_6369,N_6785);
nand U8477 (N_8477,N_7447,N_7122);
xor U8478 (N_8478,N_7328,N_6314);
or U8479 (N_8479,N_7353,N_7245);
nand U8480 (N_8480,N_6229,N_7464);
nor U8481 (N_8481,N_6824,N_6175);
nand U8482 (N_8482,N_6442,N_7214);
or U8483 (N_8483,N_7210,N_7257);
nand U8484 (N_8484,N_6872,N_7310);
and U8485 (N_8485,N_6007,N_6720);
and U8486 (N_8486,N_7263,N_7392);
xnor U8487 (N_8487,N_7328,N_6255);
or U8488 (N_8488,N_6508,N_6793);
or U8489 (N_8489,N_7131,N_7497);
and U8490 (N_8490,N_7496,N_7129);
or U8491 (N_8491,N_6599,N_6745);
xor U8492 (N_8492,N_6977,N_7228);
nand U8493 (N_8493,N_6788,N_6955);
nand U8494 (N_8494,N_6193,N_6680);
nor U8495 (N_8495,N_6802,N_6957);
or U8496 (N_8496,N_6455,N_6875);
or U8497 (N_8497,N_6659,N_6145);
nand U8498 (N_8498,N_6452,N_7220);
nor U8499 (N_8499,N_6680,N_7061);
nor U8500 (N_8500,N_7045,N_6674);
xnor U8501 (N_8501,N_6241,N_7208);
nand U8502 (N_8502,N_6568,N_7456);
nand U8503 (N_8503,N_6344,N_7276);
nor U8504 (N_8504,N_6412,N_7121);
nand U8505 (N_8505,N_6467,N_6777);
or U8506 (N_8506,N_6163,N_6953);
or U8507 (N_8507,N_7163,N_7409);
nor U8508 (N_8508,N_6915,N_7428);
and U8509 (N_8509,N_6034,N_6791);
and U8510 (N_8510,N_6075,N_6230);
or U8511 (N_8511,N_7158,N_6411);
and U8512 (N_8512,N_6928,N_6907);
and U8513 (N_8513,N_6383,N_7486);
nor U8514 (N_8514,N_6167,N_6386);
and U8515 (N_8515,N_7212,N_7085);
nand U8516 (N_8516,N_7223,N_6954);
nor U8517 (N_8517,N_6428,N_6372);
or U8518 (N_8518,N_6172,N_6826);
nor U8519 (N_8519,N_6860,N_6974);
or U8520 (N_8520,N_7076,N_6278);
nor U8521 (N_8521,N_6652,N_6438);
xor U8522 (N_8522,N_6495,N_6650);
and U8523 (N_8523,N_6927,N_6670);
and U8524 (N_8524,N_6376,N_7155);
or U8525 (N_8525,N_6216,N_6252);
xor U8526 (N_8526,N_6818,N_7426);
and U8527 (N_8527,N_6173,N_6882);
nor U8528 (N_8528,N_6853,N_6450);
or U8529 (N_8529,N_6174,N_6056);
nand U8530 (N_8530,N_7118,N_7294);
and U8531 (N_8531,N_7441,N_6339);
and U8532 (N_8532,N_7375,N_7138);
nand U8533 (N_8533,N_7014,N_7176);
nor U8534 (N_8534,N_7277,N_6784);
nor U8535 (N_8535,N_6017,N_6136);
or U8536 (N_8536,N_6041,N_7429);
or U8537 (N_8537,N_7331,N_6916);
nand U8538 (N_8538,N_6035,N_6741);
xnor U8539 (N_8539,N_6674,N_7461);
and U8540 (N_8540,N_6366,N_7238);
and U8541 (N_8541,N_6097,N_7397);
nor U8542 (N_8542,N_6958,N_6576);
or U8543 (N_8543,N_6388,N_7055);
and U8544 (N_8544,N_6223,N_6421);
nor U8545 (N_8545,N_7075,N_7096);
nand U8546 (N_8546,N_7127,N_7295);
or U8547 (N_8547,N_7456,N_6380);
nor U8548 (N_8548,N_6910,N_6292);
and U8549 (N_8549,N_6686,N_6312);
xor U8550 (N_8550,N_7040,N_6175);
nand U8551 (N_8551,N_6716,N_7001);
nor U8552 (N_8552,N_7382,N_6452);
nand U8553 (N_8553,N_7037,N_7348);
or U8554 (N_8554,N_6404,N_7032);
or U8555 (N_8555,N_6768,N_6840);
or U8556 (N_8556,N_7478,N_6286);
or U8557 (N_8557,N_6688,N_6740);
or U8558 (N_8558,N_6909,N_7380);
nand U8559 (N_8559,N_7476,N_6532);
and U8560 (N_8560,N_7452,N_6092);
and U8561 (N_8561,N_7296,N_6506);
nor U8562 (N_8562,N_6723,N_7011);
or U8563 (N_8563,N_6166,N_6969);
and U8564 (N_8564,N_7278,N_7035);
nand U8565 (N_8565,N_7181,N_6624);
nand U8566 (N_8566,N_6432,N_6448);
or U8567 (N_8567,N_6327,N_7303);
nand U8568 (N_8568,N_7315,N_6042);
or U8569 (N_8569,N_6425,N_6418);
and U8570 (N_8570,N_6821,N_6563);
nor U8571 (N_8571,N_7147,N_6523);
nand U8572 (N_8572,N_7445,N_6710);
nand U8573 (N_8573,N_6880,N_7467);
or U8574 (N_8574,N_6196,N_6031);
or U8575 (N_8575,N_6223,N_6096);
or U8576 (N_8576,N_6568,N_6400);
nor U8577 (N_8577,N_6444,N_6261);
nand U8578 (N_8578,N_6595,N_6898);
nor U8579 (N_8579,N_6278,N_6313);
nor U8580 (N_8580,N_7025,N_6988);
or U8581 (N_8581,N_6694,N_6576);
nor U8582 (N_8582,N_6428,N_6228);
or U8583 (N_8583,N_7484,N_6400);
or U8584 (N_8584,N_7109,N_7202);
nor U8585 (N_8585,N_7169,N_6321);
and U8586 (N_8586,N_6170,N_7081);
nand U8587 (N_8587,N_7056,N_6110);
nand U8588 (N_8588,N_7421,N_7358);
xor U8589 (N_8589,N_6448,N_7032);
or U8590 (N_8590,N_6974,N_6165);
xor U8591 (N_8591,N_7134,N_6730);
xnor U8592 (N_8592,N_7449,N_6619);
nor U8593 (N_8593,N_6678,N_6627);
or U8594 (N_8594,N_6771,N_6268);
or U8595 (N_8595,N_6624,N_6198);
nor U8596 (N_8596,N_6347,N_6811);
xor U8597 (N_8597,N_6754,N_7461);
or U8598 (N_8598,N_7230,N_7343);
or U8599 (N_8599,N_6784,N_7204);
and U8600 (N_8600,N_7356,N_6600);
and U8601 (N_8601,N_6124,N_6297);
and U8602 (N_8602,N_6972,N_7315);
nand U8603 (N_8603,N_6489,N_6394);
and U8604 (N_8604,N_6054,N_6286);
or U8605 (N_8605,N_6105,N_7326);
and U8606 (N_8606,N_7496,N_6477);
nor U8607 (N_8607,N_6818,N_6068);
and U8608 (N_8608,N_6728,N_6195);
nand U8609 (N_8609,N_6200,N_6961);
and U8610 (N_8610,N_6724,N_6380);
or U8611 (N_8611,N_7410,N_6508);
or U8612 (N_8612,N_7095,N_7169);
or U8613 (N_8613,N_7151,N_6205);
nor U8614 (N_8614,N_7052,N_6530);
nand U8615 (N_8615,N_7276,N_6273);
nor U8616 (N_8616,N_6887,N_7313);
or U8617 (N_8617,N_6360,N_6224);
and U8618 (N_8618,N_6320,N_6661);
nor U8619 (N_8619,N_6704,N_7097);
xnor U8620 (N_8620,N_6525,N_6625);
nor U8621 (N_8621,N_6306,N_6624);
or U8622 (N_8622,N_6099,N_6423);
nor U8623 (N_8623,N_7416,N_6775);
nor U8624 (N_8624,N_7394,N_6660);
nand U8625 (N_8625,N_7422,N_7189);
and U8626 (N_8626,N_6907,N_6126);
nand U8627 (N_8627,N_7042,N_6860);
and U8628 (N_8628,N_7081,N_6491);
nand U8629 (N_8629,N_6622,N_6420);
and U8630 (N_8630,N_6636,N_6098);
nand U8631 (N_8631,N_6005,N_6374);
or U8632 (N_8632,N_6274,N_6751);
nor U8633 (N_8633,N_6170,N_7203);
nor U8634 (N_8634,N_6987,N_6376);
and U8635 (N_8635,N_6867,N_6184);
nor U8636 (N_8636,N_7307,N_6488);
and U8637 (N_8637,N_6247,N_6839);
and U8638 (N_8638,N_7231,N_6302);
and U8639 (N_8639,N_6551,N_7220);
and U8640 (N_8640,N_6729,N_7062);
nor U8641 (N_8641,N_7257,N_6317);
xnor U8642 (N_8642,N_7421,N_7322);
and U8643 (N_8643,N_6639,N_6343);
nor U8644 (N_8644,N_6280,N_7472);
xnor U8645 (N_8645,N_6078,N_6477);
and U8646 (N_8646,N_6371,N_6367);
nand U8647 (N_8647,N_6391,N_7225);
nand U8648 (N_8648,N_6362,N_6095);
or U8649 (N_8649,N_6514,N_7462);
nor U8650 (N_8650,N_7315,N_7030);
nand U8651 (N_8651,N_6215,N_7232);
nor U8652 (N_8652,N_7254,N_7301);
and U8653 (N_8653,N_6874,N_6500);
xnor U8654 (N_8654,N_6638,N_7023);
and U8655 (N_8655,N_6552,N_6657);
xor U8656 (N_8656,N_7128,N_6060);
xnor U8657 (N_8657,N_6939,N_6178);
nor U8658 (N_8658,N_7484,N_7132);
and U8659 (N_8659,N_6620,N_6627);
nor U8660 (N_8660,N_6004,N_6337);
or U8661 (N_8661,N_7307,N_6917);
or U8662 (N_8662,N_6603,N_6633);
xnor U8663 (N_8663,N_6764,N_6739);
xor U8664 (N_8664,N_7404,N_6956);
nor U8665 (N_8665,N_6661,N_6507);
nand U8666 (N_8666,N_6992,N_7453);
xnor U8667 (N_8667,N_7207,N_6120);
nor U8668 (N_8668,N_6028,N_6013);
xnor U8669 (N_8669,N_6609,N_6355);
xnor U8670 (N_8670,N_6460,N_6696);
and U8671 (N_8671,N_7332,N_6832);
xnor U8672 (N_8672,N_7181,N_6165);
and U8673 (N_8673,N_7101,N_6443);
or U8674 (N_8674,N_6636,N_6136);
and U8675 (N_8675,N_6454,N_7014);
and U8676 (N_8676,N_6008,N_6200);
nand U8677 (N_8677,N_6961,N_6046);
xor U8678 (N_8678,N_7431,N_6686);
nor U8679 (N_8679,N_6542,N_6953);
and U8680 (N_8680,N_6343,N_6861);
nand U8681 (N_8681,N_6341,N_6923);
and U8682 (N_8682,N_6914,N_6878);
or U8683 (N_8683,N_6347,N_6725);
nand U8684 (N_8684,N_6683,N_7255);
or U8685 (N_8685,N_6112,N_7178);
nand U8686 (N_8686,N_6567,N_7016);
nor U8687 (N_8687,N_7226,N_6033);
nor U8688 (N_8688,N_7482,N_6587);
xnor U8689 (N_8689,N_6283,N_6790);
nand U8690 (N_8690,N_6695,N_6427);
and U8691 (N_8691,N_6452,N_6859);
nand U8692 (N_8692,N_6654,N_6869);
nand U8693 (N_8693,N_6195,N_6246);
nor U8694 (N_8694,N_6057,N_7003);
nand U8695 (N_8695,N_7435,N_6337);
or U8696 (N_8696,N_6213,N_7481);
or U8697 (N_8697,N_6932,N_7415);
xor U8698 (N_8698,N_6791,N_6731);
or U8699 (N_8699,N_7226,N_6911);
nor U8700 (N_8700,N_7236,N_7311);
xor U8701 (N_8701,N_6926,N_7021);
and U8702 (N_8702,N_6251,N_6941);
nor U8703 (N_8703,N_6062,N_7167);
nand U8704 (N_8704,N_6579,N_7310);
nor U8705 (N_8705,N_7127,N_6731);
nor U8706 (N_8706,N_6268,N_6184);
and U8707 (N_8707,N_7292,N_6041);
xor U8708 (N_8708,N_6630,N_6636);
or U8709 (N_8709,N_6313,N_7062);
nor U8710 (N_8710,N_6208,N_7040);
nor U8711 (N_8711,N_6805,N_6405);
and U8712 (N_8712,N_7106,N_6964);
nor U8713 (N_8713,N_6331,N_6133);
xnor U8714 (N_8714,N_6737,N_6235);
nand U8715 (N_8715,N_7216,N_6486);
or U8716 (N_8716,N_6851,N_7448);
and U8717 (N_8717,N_6689,N_6574);
or U8718 (N_8718,N_6811,N_7298);
or U8719 (N_8719,N_6506,N_6030);
nand U8720 (N_8720,N_6862,N_6432);
nor U8721 (N_8721,N_6547,N_6546);
nor U8722 (N_8722,N_6644,N_7395);
nand U8723 (N_8723,N_6342,N_6085);
nand U8724 (N_8724,N_6781,N_6516);
nand U8725 (N_8725,N_6886,N_6924);
or U8726 (N_8726,N_6258,N_7417);
and U8727 (N_8727,N_7042,N_6424);
nor U8728 (N_8728,N_6605,N_6603);
nor U8729 (N_8729,N_7255,N_6121);
nor U8730 (N_8730,N_6502,N_6072);
or U8731 (N_8731,N_6338,N_7002);
or U8732 (N_8732,N_6713,N_7085);
and U8733 (N_8733,N_6219,N_6794);
and U8734 (N_8734,N_6087,N_6869);
or U8735 (N_8735,N_6764,N_6420);
xor U8736 (N_8736,N_6171,N_6211);
and U8737 (N_8737,N_6276,N_7243);
xnor U8738 (N_8738,N_7445,N_6346);
nand U8739 (N_8739,N_7219,N_7051);
and U8740 (N_8740,N_7488,N_7417);
and U8741 (N_8741,N_6772,N_6845);
and U8742 (N_8742,N_7160,N_6731);
nand U8743 (N_8743,N_7423,N_7487);
and U8744 (N_8744,N_7480,N_7238);
nor U8745 (N_8745,N_6998,N_7243);
nor U8746 (N_8746,N_7334,N_6979);
nand U8747 (N_8747,N_6600,N_6159);
and U8748 (N_8748,N_7230,N_7328);
nor U8749 (N_8749,N_7319,N_6494);
nand U8750 (N_8750,N_6597,N_7455);
nand U8751 (N_8751,N_6465,N_7263);
or U8752 (N_8752,N_6564,N_6028);
and U8753 (N_8753,N_6565,N_7077);
and U8754 (N_8754,N_6688,N_6405);
nor U8755 (N_8755,N_7182,N_7155);
nor U8756 (N_8756,N_6933,N_6313);
nand U8757 (N_8757,N_7240,N_6597);
nor U8758 (N_8758,N_6704,N_6561);
and U8759 (N_8759,N_6030,N_6625);
xnor U8760 (N_8760,N_6676,N_7125);
nand U8761 (N_8761,N_7419,N_6464);
nand U8762 (N_8762,N_6738,N_7115);
and U8763 (N_8763,N_6235,N_6987);
or U8764 (N_8764,N_6608,N_6135);
nand U8765 (N_8765,N_6900,N_6702);
xnor U8766 (N_8766,N_6958,N_7052);
nor U8767 (N_8767,N_6008,N_6982);
nor U8768 (N_8768,N_6352,N_7260);
nand U8769 (N_8769,N_7410,N_7188);
and U8770 (N_8770,N_7139,N_6239);
nor U8771 (N_8771,N_6953,N_7316);
nor U8772 (N_8772,N_6832,N_7047);
xnor U8773 (N_8773,N_7029,N_6690);
and U8774 (N_8774,N_6092,N_7142);
nor U8775 (N_8775,N_6888,N_7068);
or U8776 (N_8776,N_6933,N_6218);
and U8777 (N_8777,N_7197,N_6594);
nor U8778 (N_8778,N_6399,N_6696);
nand U8779 (N_8779,N_6773,N_7096);
or U8780 (N_8780,N_7407,N_7156);
or U8781 (N_8781,N_6308,N_6959);
nand U8782 (N_8782,N_6988,N_6710);
and U8783 (N_8783,N_7138,N_6127);
nor U8784 (N_8784,N_6519,N_6329);
nand U8785 (N_8785,N_6594,N_7029);
nand U8786 (N_8786,N_7114,N_6369);
or U8787 (N_8787,N_6372,N_6160);
nand U8788 (N_8788,N_6946,N_7063);
or U8789 (N_8789,N_6002,N_7367);
nor U8790 (N_8790,N_6716,N_6356);
nor U8791 (N_8791,N_7178,N_6423);
nand U8792 (N_8792,N_6414,N_6135);
nand U8793 (N_8793,N_6472,N_7045);
or U8794 (N_8794,N_6553,N_6026);
and U8795 (N_8795,N_6366,N_6807);
xnor U8796 (N_8796,N_6839,N_7343);
nor U8797 (N_8797,N_6737,N_6308);
nor U8798 (N_8798,N_7215,N_6358);
nand U8799 (N_8799,N_7265,N_6160);
and U8800 (N_8800,N_6584,N_6760);
nand U8801 (N_8801,N_6565,N_6009);
or U8802 (N_8802,N_6142,N_7042);
nand U8803 (N_8803,N_6092,N_7343);
nand U8804 (N_8804,N_7267,N_7459);
xnor U8805 (N_8805,N_6261,N_6366);
nand U8806 (N_8806,N_6957,N_6320);
nand U8807 (N_8807,N_6167,N_6610);
xnor U8808 (N_8808,N_7199,N_6415);
or U8809 (N_8809,N_6103,N_7088);
or U8810 (N_8810,N_6468,N_6486);
xor U8811 (N_8811,N_7123,N_6268);
or U8812 (N_8812,N_6104,N_7023);
nand U8813 (N_8813,N_6991,N_6142);
nor U8814 (N_8814,N_6445,N_7145);
or U8815 (N_8815,N_7381,N_6454);
and U8816 (N_8816,N_6286,N_7128);
nor U8817 (N_8817,N_6708,N_7485);
and U8818 (N_8818,N_6270,N_6268);
nand U8819 (N_8819,N_6330,N_6233);
and U8820 (N_8820,N_6417,N_6103);
nand U8821 (N_8821,N_6468,N_7176);
nor U8822 (N_8822,N_7229,N_6442);
nand U8823 (N_8823,N_6930,N_6698);
nor U8824 (N_8824,N_6988,N_7145);
and U8825 (N_8825,N_6511,N_7283);
or U8826 (N_8826,N_7031,N_6254);
and U8827 (N_8827,N_6135,N_7280);
xor U8828 (N_8828,N_7473,N_6356);
or U8829 (N_8829,N_7273,N_7134);
nand U8830 (N_8830,N_7010,N_6553);
nor U8831 (N_8831,N_6387,N_6258);
and U8832 (N_8832,N_6990,N_7119);
nor U8833 (N_8833,N_6051,N_6266);
and U8834 (N_8834,N_7027,N_6224);
nor U8835 (N_8835,N_6644,N_7186);
nor U8836 (N_8836,N_7389,N_6603);
or U8837 (N_8837,N_6402,N_7250);
and U8838 (N_8838,N_7380,N_6549);
or U8839 (N_8839,N_6301,N_6051);
nand U8840 (N_8840,N_7117,N_6429);
nand U8841 (N_8841,N_6792,N_7029);
nand U8842 (N_8842,N_6480,N_7157);
nor U8843 (N_8843,N_7259,N_7172);
and U8844 (N_8844,N_7167,N_6079);
or U8845 (N_8845,N_6245,N_6323);
nor U8846 (N_8846,N_7303,N_7164);
nor U8847 (N_8847,N_6934,N_6177);
nor U8848 (N_8848,N_6709,N_6924);
and U8849 (N_8849,N_7258,N_6273);
and U8850 (N_8850,N_6686,N_6170);
or U8851 (N_8851,N_6216,N_6037);
nand U8852 (N_8852,N_6242,N_7054);
nor U8853 (N_8853,N_6863,N_6793);
nand U8854 (N_8854,N_6807,N_6131);
nor U8855 (N_8855,N_6383,N_7347);
or U8856 (N_8856,N_6340,N_6147);
nand U8857 (N_8857,N_6354,N_7235);
and U8858 (N_8858,N_6894,N_6954);
and U8859 (N_8859,N_6331,N_6793);
or U8860 (N_8860,N_7429,N_6042);
or U8861 (N_8861,N_7146,N_6906);
and U8862 (N_8862,N_6183,N_7138);
and U8863 (N_8863,N_6918,N_6695);
xor U8864 (N_8864,N_6178,N_7033);
or U8865 (N_8865,N_7361,N_7255);
or U8866 (N_8866,N_7076,N_7014);
nand U8867 (N_8867,N_6722,N_7302);
and U8868 (N_8868,N_6170,N_6897);
nand U8869 (N_8869,N_6596,N_7097);
nand U8870 (N_8870,N_6456,N_7415);
nand U8871 (N_8871,N_7011,N_6088);
nand U8872 (N_8872,N_6973,N_7069);
nor U8873 (N_8873,N_6280,N_6690);
nand U8874 (N_8874,N_6933,N_6105);
nor U8875 (N_8875,N_6281,N_6665);
nor U8876 (N_8876,N_6259,N_6027);
and U8877 (N_8877,N_6330,N_7052);
xor U8878 (N_8878,N_7476,N_6153);
nor U8879 (N_8879,N_6979,N_6792);
and U8880 (N_8880,N_6327,N_6231);
nand U8881 (N_8881,N_7445,N_7172);
and U8882 (N_8882,N_7427,N_6067);
and U8883 (N_8883,N_6708,N_6563);
nor U8884 (N_8884,N_7494,N_6684);
nor U8885 (N_8885,N_6999,N_7123);
or U8886 (N_8886,N_6661,N_7042);
nor U8887 (N_8887,N_7194,N_6021);
nand U8888 (N_8888,N_6848,N_7461);
or U8889 (N_8889,N_6923,N_6104);
nand U8890 (N_8890,N_6585,N_6531);
nor U8891 (N_8891,N_6568,N_7062);
nand U8892 (N_8892,N_6230,N_7190);
or U8893 (N_8893,N_6646,N_6609);
nor U8894 (N_8894,N_7077,N_7289);
or U8895 (N_8895,N_6325,N_6179);
nand U8896 (N_8896,N_6073,N_7031);
xnor U8897 (N_8897,N_7253,N_7007);
and U8898 (N_8898,N_6988,N_6957);
xor U8899 (N_8899,N_6384,N_6359);
xor U8900 (N_8900,N_6262,N_6458);
nor U8901 (N_8901,N_6006,N_6819);
nor U8902 (N_8902,N_7381,N_6553);
and U8903 (N_8903,N_6854,N_7429);
and U8904 (N_8904,N_6964,N_6932);
and U8905 (N_8905,N_7346,N_7077);
nand U8906 (N_8906,N_6127,N_6670);
or U8907 (N_8907,N_6043,N_7379);
or U8908 (N_8908,N_6338,N_7381);
and U8909 (N_8909,N_6275,N_7010);
nor U8910 (N_8910,N_7456,N_6918);
and U8911 (N_8911,N_6357,N_7268);
nor U8912 (N_8912,N_7132,N_6145);
or U8913 (N_8913,N_6874,N_6510);
nand U8914 (N_8914,N_6470,N_6466);
or U8915 (N_8915,N_6051,N_7445);
xor U8916 (N_8916,N_7477,N_6416);
nor U8917 (N_8917,N_6774,N_6873);
nor U8918 (N_8918,N_7194,N_6998);
and U8919 (N_8919,N_6259,N_6733);
nor U8920 (N_8920,N_6612,N_6190);
or U8921 (N_8921,N_7264,N_7138);
and U8922 (N_8922,N_6884,N_6578);
or U8923 (N_8923,N_6129,N_7205);
or U8924 (N_8924,N_6318,N_6487);
nand U8925 (N_8925,N_6831,N_6912);
and U8926 (N_8926,N_7077,N_6660);
nand U8927 (N_8927,N_6678,N_6111);
nand U8928 (N_8928,N_6790,N_6631);
or U8929 (N_8929,N_7258,N_6390);
and U8930 (N_8930,N_6741,N_7004);
xnor U8931 (N_8931,N_6501,N_7251);
and U8932 (N_8932,N_6444,N_7479);
nand U8933 (N_8933,N_6745,N_7214);
and U8934 (N_8934,N_6574,N_6239);
or U8935 (N_8935,N_6711,N_6250);
nand U8936 (N_8936,N_7327,N_6007);
nor U8937 (N_8937,N_7315,N_6427);
nand U8938 (N_8938,N_6249,N_6605);
xor U8939 (N_8939,N_6109,N_6205);
or U8940 (N_8940,N_7227,N_7494);
nand U8941 (N_8941,N_6011,N_6075);
xor U8942 (N_8942,N_6734,N_6703);
nor U8943 (N_8943,N_6627,N_6110);
or U8944 (N_8944,N_7473,N_7372);
nand U8945 (N_8945,N_6345,N_7319);
nand U8946 (N_8946,N_7398,N_6733);
nand U8947 (N_8947,N_7272,N_6815);
or U8948 (N_8948,N_7428,N_7426);
nor U8949 (N_8949,N_7110,N_6278);
nor U8950 (N_8950,N_6397,N_7371);
nand U8951 (N_8951,N_7072,N_6592);
and U8952 (N_8952,N_6479,N_6462);
nor U8953 (N_8953,N_6004,N_6244);
and U8954 (N_8954,N_6680,N_6177);
nor U8955 (N_8955,N_6821,N_7150);
nand U8956 (N_8956,N_7472,N_6558);
nor U8957 (N_8957,N_6472,N_6309);
or U8958 (N_8958,N_6190,N_6127);
nand U8959 (N_8959,N_6891,N_6505);
and U8960 (N_8960,N_7416,N_6433);
nand U8961 (N_8961,N_6419,N_6937);
or U8962 (N_8962,N_6784,N_7417);
nor U8963 (N_8963,N_6530,N_6590);
or U8964 (N_8964,N_6220,N_7287);
and U8965 (N_8965,N_6136,N_6693);
nor U8966 (N_8966,N_6675,N_6158);
and U8967 (N_8967,N_7016,N_6383);
nand U8968 (N_8968,N_7097,N_7248);
and U8969 (N_8969,N_7386,N_7109);
or U8970 (N_8970,N_6117,N_6203);
or U8971 (N_8971,N_7201,N_6063);
xnor U8972 (N_8972,N_6828,N_6342);
nor U8973 (N_8973,N_7420,N_6571);
or U8974 (N_8974,N_6992,N_7156);
nand U8975 (N_8975,N_7289,N_6468);
or U8976 (N_8976,N_6346,N_6758);
or U8977 (N_8977,N_6932,N_6508);
and U8978 (N_8978,N_7219,N_6021);
and U8979 (N_8979,N_6782,N_6467);
nand U8980 (N_8980,N_6386,N_7117);
xor U8981 (N_8981,N_6926,N_6746);
or U8982 (N_8982,N_6025,N_6193);
nor U8983 (N_8983,N_7332,N_6423);
or U8984 (N_8984,N_6290,N_7256);
nand U8985 (N_8985,N_6652,N_7047);
and U8986 (N_8986,N_6921,N_6325);
nor U8987 (N_8987,N_6655,N_6270);
and U8988 (N_8988,N_6592,N_7094);
nand U8989 (N_8989,N_6872,N_7130);
and U8990 (N_8990,N_6065,N_6632);
and U8991 (N_8991,N_7496,N_6079);
xnor U8992 (N_8992,N_6656,N_6266);
and U8993 (N_8993,N_6691,N_6008);
and U8994 (N_8994,N_7375,N_7242);
nand U8995 (N_8995,N_6189,N_7024);
nor U8996 (N_8996,N_6573,N_7410);
nand U8997 (N_8997,N_7485,N_6427);
nor U8998 (N_8998,N_7006,N_6550);
or U8999 (N_8999,N_6544,N_6751);
nor U9000 (N_9000,N_8242,N_7531);
nand U9001 (N_9001,N_8469,N_8507);
xor U9002 (N_9002,N_8705,N_8014);
or U9003 (N_9003,N_8930,N_8569);
nand U9004 (N_9004,N_7891,N_8187);
nand U9005 (N_9005,N_8832,N_8167);
xnor U9006 (N_9006,N_7654,N_8642);
or U9007 (N_9007,N_8075,N_7853);
nand U9008 (N_9008,N_8621,N_8882);
or U9009 (N_9009,N_7994,N_7593);
and U9010 (N_9010,N_8160,N_7665);
nand U9011 (N_9011,N_8592,N_7591);
nor U9012 (N_9012,N_7752,N_7524);
nor U9013 (N_9013,N_8750,N_7921);
and U9014 (N_9014,N_7525,N_7913);
nand U9015 (N_9015,N_8227,N_7661);
nor U9016 (N_9016,N_8541,N_8009);
nor U9017 (N_9017,N_8808,N_7727);
nand U9018 (N_9018,N_8931,N_7729);
xnor U9019 (N_9019,N_7938,N_8021);
or U9020 (N_9020,N_7579,N_8577);
xor U9021 (N_9021,N_7588,N_7605);
xnor U9022 (N_9022,N_8258,N_8069);
and U9023 (N_9023,N_8056,N_8364);
and U9024 (N_9024,N_8863,N_8399);
and U9025 (N_9025,N_7587,N_7860);
or U9026 (N_9026,N_7718,N_8422);
and U9027 (N_9027,N_7970,N_7825);
nand U9028 (N_9028,N_8086,N_7968);
or U9029 (N_9029,N_8235,N_8264);
nand U9030 (N_9030,N_7804,N_8827);
nand U9031 (N_9031,N_7644,N_7864);
or U9032 (N_9032,N_8620,N_8505);
and U9033 (N_9033,N_8408,N_7540);
or U9034 (N_9034,N_8550,N_8736);
nor U9035 (N_9035,N_8945,N_8968);
nor U9036 (N_9036,N_8983,N_8270);
or U9037 (N_9037,N_8532,N_8654);
nand U9038 (N_9038,N_8022,N_8209);
or U9039 (N_9039,N_8825,N_8011);
or U9040 (N_9040,N_7966,N_8959);
nand U9041 (N_9041,N_7725,N_8820);
nand U9042 (N_9042,N_7926,N_8023);
and U9043 (N_9043,N_7716,N_8604);
or U9044 (N_9044,N_7851,N_8783);
nor U9045 (N_9045,N_8907,N_7557);
nor U9046 (N_9046,N_7739,N_8530);
nor U9047 (N_9047,N_7855,N_8026);
nor U9048 (N_9048,N_8984,N_7656);
or U9049 (N_9049,N_7694,N_8581);
nor U9050 (N_9050,N_8551,N_7614);
and U9051 (N_9051,N_8282,N_7563);
or U9052 (N_9052,N_7936,N_7880);
nand U9053 (N_9053,N_7801,N_8338);
and U9054 (N_9054,N_8899,N_8673);
nor U9055 (N_9055,N_8094,N_8400);
nor U9056 (N_9056,N_8320,N_7840);
nor U9057 (N_9057,N_8644,N_7923);
nand U9058 (N_9058,N_8806,N_8564);
or U9059 (N_9059,N_8097,N_8156);
nor U9060 (N_9060,N_8589,N_7998);
nand U9061 (N_9061,N_7874,N_7599);
and U9062 (N_9062,N_7683,N_8789);
nor U9063 (N_9063,N_7712,N_7693);
and U9064 (N_9064,N_8918,N_7787);
nand U9065 (N_9065,N_8043,N_7948);
or U9066 (N_9066,N_7818,N_8548);
and U9067 (N_9067,N_8451,N_8689);
or U9068 (N_9068,N_8535,N_7626);
nand U9069 (N_9069,N_8509,N_8200);
nor U9070 (N_9070,N_8842,N_8031);
and U9071 (N_9071,N_8328,N_8168);
nand U9072 (N_9072,N_8602,N_8652);
nand U9073 (N_9073,N_7771,N_7511);
and U9074 (N_9074,N_7692,N_7810);
nor U9075 (N_9075,N_7709,N_7543);
xor U9076 (N_9076,N_8790,N_7522);
and U9077 (N_9077,N_8138,N_7909);
xnor U9078 (N_9078,N_7786,N_8908);
and U9079 (N_9079,N_8275,N_8429);
nand U9080 (N_9080,N_8524,N_7581);
xor U9081 (N_9081,N_8609,N_8890);
and U9082 (N_9082,N_7737,N_7837);
nor U9083 (N_9083,N_8278,N_8543);
xor U9084 (N_9084,N_7941,N_7514);
and U9085 (N_9085,N_7987,N_7854);
nor U9086 (N_9086,N_8103,N_8397);
xnor U9087 (N_9087,N_8841,N_7770);
or U9088 (N_9088,N_8540,N_8512);
nor U9089 (N_9089,N_7884,N_7567);
and U9090 (N_9090,N_8109,N_8361);
or U9091 (N_9091,N_8089,N_7964);
nand U9092 (N_9092,N_8889,N_7623);
or U9093 (N_9093,N_8440,N_8517);
nand U9094 (N_9094,N_8865,N_8647);
nand U9095 (N_9095,N_8991,N_7643);
nand U9096 (N_9096,N_7832,N_8062);
or U9097 (N_9097,N_8926,N_8615);
nor U9098 (N_9098,N_8005,N_8566);
or U9099 (N_9099,N_8972,N_7714);
xor U9100 (N_9100,N_8101,N_8283);
nor U9101 (N_9101,N_7546,N_7549);
xor U9102 (N_9102,N_7753,N_8727);
xor U9103 (N_9103,N_8100,N_8775);
or U9104 (N_9104,N_8586,N_8289);
nand U9105 (N_9105,N_8963,N_8406);
nor U9106 (N_9106,N_7595,N_7889);
and U9107 (N_9107,N_8288,N_7611);
or U9108 (N_9108,N_7843,N_8178);
and U9109 (N_9109,N_8322,N_7877);
or U9110 (N_9110,N_8096,N_8631);
nand U9111 (N_9111,N_7664,N_8538);
and U9112 (N_9112,N_8302,N_8650);
xnor U9113 (N_9113,N_7585,N_7648);
and U9114 (N_9114,N_8117,N_7646);
nand U9115 (N_9115,N_7710,N_8247);
and U9116 (N_9116,N_8910,N_7780);
xnor U9117 (N_9117,N_7691,N_7961);
and U9118 (N_9118,N_8396,N_8822);
nor U9119 (N_9119,N_8697,N_8957);
or U9120 (N_9120,N_8425,N_8157);
or U9121 (N_9121,N_8664,N_8619);
xor U9122 (N_9122,N_8660,N_8271);
nor U9123 (N_9123,N_7735,N_8266);
nand U9124 (N_9124,N_8537,N_7507);
or U9125 (N_9125,N_8353,N_7930);
nor U9126 (N_9126,N_8737,N_8403);
and U9127 (N_9127,N_8110,N_8444);
nor U9128 (N_9128,N_7902,N_8210);
nor U9129 (N_9129,N_8600,N_8716);
nand U9130 (N_9130,N_8852,N_7527);
nand U9131 (N_9131,N_8587,N_8421);
or U9132 (N_9132,N_7895,N_8061);
nor U9133 (N_9133,N_7871,N_8107);
nand U9134 (N_9134,N_8277,N_8902);
nor U9135 (N_9135,N_8853,N_8259);
xor U9136 (N_9136,N_8297,N_8738);
nor U9137 (N_9137,N_8446,N_8035);
or U9138 (N_9138,N_8504,N_8758);
nor U9139 (N_9139,N_8601,N_7675);
and U9140 (N_9140,N_7845,N_8641);
nor U9141 (N_9141,N_8699,N_7820);
or U9142 (N_9142,N_8267,N_8241);
and U9143 (N_9143,N_8748,N_8950);
and U9144 (N_9144,N_7898,N_7669);
or U9145 (N_9145,N_8260,N_8552);
or U9146 (N_9146,N_7858,N_8745);
xor U9147 (N_9147,N_7751,N_8257);
nand U9148 (N_9148,N_8154,N_8503);
and U9149 (N_9149,N_8805,N_8800);
and U9150 (N_9150,N_7835,N_8340);
and U9151 (N_9151,N_8424,N_8730);
nor U9152 (N_9152,N_8268,N_8506);
nor U9153 (N_9153,N_8857,N_8966);
and U9154 (N_9154,N_7575,N_8747);
and U9155 (N_9155,N_7977,N_8939);
or U9156 (N_9156,N_8753,N_8152);
nor U9157 (N_9157,N_8012,N_8571);
and U9158 (N_9158,N_7668,N_7793);
or U9159 (N_9159,N_8801,N_8638);
and U9160 (N_9160,N_8193,N_8828);
and U9161 (N_9161,N_8740,N_8007);
nand U9162 (N_9162,N_8793,N_7848);
nand U9163 (N_9163,N_7897,N_8911);
nor U9164 (N_9164,N_7564,N_8561);
nor U9165 (N_9165,N_8462,N_8804);
and U9166 (N_9166,N_8778,N_8237);
xnor U9167 (N_9167,N_8625,N_8205);
and U9168 (N_9168,N_7574,N_8090);
xor U9169 (N_9169,N_7687,N_7682);
and U9170 (N_9170,N_8002,N_8649);
nor U9171 (N_9171,N_8690,N_8389);
nor U9172 (N_9172,N_8262,N_8667);
and U9173 (N_9173,N_7621,N_8946);
or U9174 (N_9174,N_8327,N_8643);
and U9175 (N_9175,N_8224,N_8719);
xnor U9176 (N_9176,N_7502,N_7911);
and U9177 (N_9177,N_8346,N_7728);
nor U9178 (N_9178,N_8752,N_8325);
or U9179 (N_9179,N_8197,N_7530);
or U9180 (N_9180,N_8384,N_7779);
or U9181 (N_9181,N_7500,N_8850);
nand U9182 (N_9182,N_7625,N_8420);
or U9183 (N_9183,N_8723,N_8663);
nand U9184 (N_9184,N_8722,N_8798);
nor U9185 (N_9185,N_8878,N_8046);
xnor U9186 (N_9186,N_8941,N_7636);
nor U9187 (N_9187,N_8682,N_8236);
nand U9188 (N_9188,N_7572,N_8081);
or U9189 (N_9189,N_8198,N_8411);
xor U9190 (N_9190,N_8996,N_7633);
nand U9191 (N_9191,N_8067,N_7767);
nand U9192 (N_9192,N_8711,N_8474);
or U9193 (N_9193,N_8671,N_7501);
or U9194 (N_9194,N_8216,N_7731);
or U9195 (N_9195,N_7758,N_8127);
nor U9196 (N_9196,N_7942,N_8557);
xor U9197 (N_9197,N_7560,N_8891);
and U9198 (N_9198,N_8943,N_8868);
and U9199 (N_9199,N_8376,N_7932);
or U9200 (N_9200,N_8226,N_7886);
nor U9201 (N_9201,N_8054,N_8767);
and U9202 (N_9202,N_8489,N_7537);
and U9203 (N_9203,N_8139,N_8993);
and U9204 (N_9204,N_8239,N_8659);
nor U9205 (N_9205,N_7974,N_8580);
nor U9206 (N_9206,N_7931,N_8093);
nand U9207 (N_9207,N_8618,N_8840);
nor U9208 (N_9208,N_8279,N_8779);
and U9209 (N_9209,N_7901,N_7736);
or U9210 (N_9210,N_7912,N_8675);
xnor U9211 (N_9211,N_8533,N_8632);
and U9212 (N_9212,N_8250,N_7515);
nand U9213 (N_9213,N_8534,N_8934);
or U9214 (N_9214,N_8265,N_8414);
and U9215 (N_9215,N_7756,N_8568);
or U9216 (N_9216,N_7551,N_8276);
or U9217 (N_9217,N_8839,N_7637);
nor U9218 (N_9218,N_8999,N_7673);
or U9219 (N_9219,N_8687,N_8718);
nand U9220 (N_9220,N_8284,N_7816);
xnor U9221 (N_9221,N_7565,N_7790);
nand U9222 (N_9222,N_7558,N_7918);
or U9223 (N_9223,N_8772,N_8831);
or U9224 (N_9224,N_7872,N_7797);
xor U9225 (N_9225,N_7956,N_7685);
nand U9226 (N_9226,N_8196,N_8102);
nand U9227 (N_9227,N_8499,N_7663);
or U9228 (N_9228,N_8872,N_7680);
xnor U9229 (N_9229,N_8544,N_8997);
nand U9230 (N_9230,N_8286,N_7606);
nand U9231 (N_9231,N_8465,N_8683);
nor U9232 (N_9232,N_8797,N_7952);
xnor U9233 (N_9233,N_8441,N_8252);
nand U9234 (N_9234,N_8662,N_8029);
or U9235 (N_9235,N_8788,N_8215);
nor U9236 (N_9236,N_7750,N_7700);
nor U9237 (N_9237,N_8217,N_7796);
or U9238 (N_9238,N_8933,N_7688);
nand U9239 (N_9239,N_7689,N_8150);
or U9240 (N_9240,N_8915,N_8634);
and U9241 (N_9241,N_8347,N_8811);
and U9242 (N_9242,N_7992,N_8481);
xnor U9243 (N_9243,N_8703,N_8058);
nor U9244 (N_9244,N_7686,N_8715);
nand U9245 (N_9245,N_8928,N_8920);
xor U9246 (N_9246,N_8686,N_8362);
nor U9247 (N_9247,N_8835,N_8803);
nor U9248 (N_9248,N_8763,N_7505);
or U9249 (N_9249,N_7681,N_8439);
xnor U9250 (N_9250,N_7713,N_8900);
nand U9251 (N_9251,N_8334,N_7844);
or U9252 (N_9252,N_7792,N_8480);
nor U9253 (N_9253,N_8377,N_8794);
xnor U9254 (N_9254,N_8243,N_7917);
nor U9255 (N_9255,N_8497,N_7984);
or U9256 (N_9256,N_7529,N_8815);
xor U9257 (N_9257,N_8856,N_8714);
or U9258 (N_9258,N_8897,N_8877);
nor U9259 (N_9259,N_8218,N_7960);
nor U9260 (N_9260,N_8375,N_8676);
nor U9261 (N_9261,N_8078,N_8597);
xnor U9262 (N_9262,N_8438,N_7678);
nand U9263 (N_9263,N_7925,N_8194);
or U9264 (N_9264,N_8245,N_8490);
xnor U9265 (N_9265,N_8706,N_7856);
nor U9266 (N_9266,N_8169,N_8762);
xnor U9267 (N_9267,N_8816,N_8887);
nand U9268 (N_9268,N_7747,N_8427);
nor U9269 (N_9269,N_7857,N_8940);
or U9270 (N_9270,N_7805,N_8073);
or U9271 (N_9271,N_7745,N_8554);
nand U9272 (N_9272,N_8881,N_8354);
or U9273 (N_9273,N_8818,N_8351);
nor U9274 (N_9274,N_8574,N_8436);
nand U9275 (N_9275,N_8536,N_8685);
nand U9276 (N_9276,N_7647,N_8492);
or U9277 (N_9277,N_8591,N_8653);
xor U9278 (N_9278,N_8136,N_8363);
nor U9279 (N_9279,N_7556,N_8498);
nor U9280 (N_9280,N_8185,N_7807);
and U9281 (N_9281,N_8859,N_7607);
nor U9282 (N_9282,N_7711,N_8883);
nor U9283 (N_9283,N_8024,N_7774);
nand U9284 (N_9284,N_7783,N_8929);
or U9285 (N_9285,N_8214,N_8336);
and U9286 (N_9286,N_7519,N_8263);
and U9287 (N_9287,N_8020,N_8843);
nand U9288 (N_9288,N_8823,N_8413);
nand U9289 (N_9289,N_8177,N_8721);
xnor U9290 (N_9290,N_7619,N_8953);
nand U9291 (N_9291,N_8596,N_7958);
nor U9292 (N_9292,N_8125,N_8371);
nand U9293 (N_9293,N_7981,N_7963);
xor U9294 (N_9294,N_8074,N_8948);
nor U9295 (N_9295,N_7809,N_7520);
nand U9296 (N_9296,N_7730,N_8385);
nor U9297 (N_9297,N_8314,N_8688);
and U9298 (N_9298,N_8759,N_7715);
nand U9299 (N_9299,N_8973,N_8179);
and U9300 (N_9300,N_7883,N_8372);
nand U9301 (N_9301,N_7562,N_8165);
or U9302 (N_9302,N_7781,N_7584);
nor U9303 (N_9303,N_7510,N_8526);
nor U9304 (N_9304,N_7831,N_8381);
and U9305 (N_9305,N_8546,N_8040);
or U9306 (N_9306,N_8848,N_7734);
nand U9307 (N_9307,N_7888,N_8851);
and U9308 (N_9308,N_8121,N_7841);
xor U9309 (N_9309,N_8341,N_8515);
nand U9310 (N_9310,N_8188,N_8287);
and U9311 (N_9311,N_8594,N_8112);
nor U9312 (N_9312,N_8545,N_8782);
nand U9313 (N_9313,N_8437,N_8922);
nor U9314 (N_9314,N_7724,N_8486);
or U9315 (N_9315,N_7914,N_8126);
or U9316 (N_9316,N_7592,N_8885);
or U9317 (N_9317,N_7629,N_8830);
nor U9318 (N_9318,N_7915,N_8605);
and U9319 (N_9319,N_8404,N_8207);
or U9320 (N_9320,N_8909,N_8016);
nor U9321 (N_9321,N_8518,N_8133);
nand U9322 (N_9322,N_8358,N_7638);
or U9323 (N_9323,N_8628,N_7996);
and U9324 (N_9324,N_8204,N_8261);
or U9325 (N_9325,N_8994,N_8180);
nor U9326 (N_9326,N_8635,N_8769);
or U9327 (N_9327,N_7568,N_7659);
nor U9328 (N_9328,N_8837,N_8978);
xor U9329 (N_9329,N_7823,N_7777);
nand U9330 (N_9330,N_7878,N_8388);
and U9331 (N_9331,N_8416,N_7632);
nor U9332 (N_9332,N_7658,N_8796);
nor U9333 (N_9333,N_8563,N_7953);
nand U9334 (N_9334,N_7577,N_8316);
and U9335 (N_9335,N_7554,N_8802);
and U9336 (N_9336,N_7763,N_8123);
nor U9337 (N_9337,N_8974,N_8124);
or U9338 (N_9338,N_7553,N_8064);
and U9339 (N_9339,N_7817,N_7699);
or U9340 (N_9340,N_8116,N_8709);
xnor U9341 (N_9341,N_8129,N_7965);
or U9342 (N_9342,N_7900,N_8454);
nor U9343 (N_9343,N_8291,N_8369);
nor U9344 (N_9344,N_7634,N_8785);
or U9345 (N_9345,N_8050,N_8076);
or U9346 (N_9346,N_7749,N_7922);
and U9347 (N_9347,N_7896,N_7892);
nand U9348 (N_9348,N_7703,N_8921);
nand U9349 (N_9349,N_8791,N_8459);
xnor U9350 (N_9350,N_7904,N_8880);
and U9351 (N_9351,N_7652,N_7865);
nor U9352 (N_9352,N_8888,N_8562);
and U9353 (N_9353,N_8624,N_8598);
xnor U9354 (N_9354,N_7822,N_8244);
nand U9355 (N_9355,N_7706,N_8448);
or U9356 (N_9356,N_8228,N_8255);
nor U9357 (N_9357,N_7516,N_8944);
nor U9358 (N_9358,N_8764,N_8903);
nor U9359 (N_9359,N_7861,N_7867);
nor U9360 (N_9360,N_7944,N_8896);
and U9361 (N_9361,N_7830,N_8549);
nor U9362 (N_9362,N_7821,N_7616);
or U9363 (N_9363,N_7833,N_8080);
nand U9364 (N_9364,N_8071,N_7766);
nand U9365 (N_9365,N_8335,N_8045);
nand U9366 (N_9366,N_7732,N_7535);
nor U9367 (N_9367,N_8114,N_7806);
and U9368 (N_9368,N_7907,N_8395);
and U9369 (N_9369,N_8761,N_8290);
nand U9370 (N_9370,N_8976,N_8980);
and U9371 (N_9371,N_8418,N_8195);
nor U9372 (N_9372,N_7755,N_8570);
or U9373 (N_9373,N_7622,N_7972);
or U9374 (N_9374,N_7513,N_7929);
or U9375 (N_9375,N_8623,N_8989);
nand U9376 (N_9376,N_8616,N_8412);
and U9377 (N_9377,N_8698,N_8161);
or U9378 (N_9378,N_8070,N_8923);
and U9379 (N_9379,N_7990,N_7708);
nand U9380 (N_9380,N_8186,N_8345);
nand U9381 (N_9381,N_7744,N_7834);
nor U9382 (N_9382,N_7959,N_8158);
xnor U9383 (N_9383,N_8443,N_8969);
and U9384 (N_9384,N_8824,N_8223);
xor U9385 (N_9385,N_8333,N_8442);
nand U9386 (N_9386,N_8331,N_7866);
and U9387 (N_9387,N_8231,N_8373);
or U9388 (N_9388,N_8661,N_8471);
and U9389 (N_9389,N_8352,N_8666);
and U9390 (N_9390,N_7982,N_7667);
xor U9391 (N_9391,N_7604,N_7875);
and U9392 (N_9392,N_8724,N_7951);
nand U9393 (N_9393,N_8329,N_7776);
and U9394 (N_9394,N_8240,N_7784);
nor U9395 (N_9395,N_8985,N_7868);
or U9396 (N_9396,N_8935,N_8047);
and U9397 (N_9397,N_8990,N_8527);
xor U9398 (N_9398,N_8799,N_8886);
nor U9399 (N_9399,N_8754,N_8182);
or U9400 (N_9400,N_8912,N_7993);
or U9401 (N_9401,N_8982,N_8428);
and U9402 (N_9402,N_8305,N_8303);
or U9403 (N_9403,N_8781,N_8479);
xor U9404 (N_9404,N_7962,N_7506);
nor U9405 (N_9405,N_7662,N_7795);
and U9406 (N_9406,N_8221,N_8144);
nand U9407 (N_9407,N_8068,N_8988);
and U9408 (N_9408,N_8203,N_8967);
nand U9409 (N_9409,N_8529,N_8051);
or U9410 (N_9410,N_8836,N_7772);
and U9411 (N_9411,N_8039,N_8206);
nor U9412 (N_9412,N_8720,N_8269);
and U9413 (N_9413,N_8300,N_8344);
xnor U9414 (N_9414,N_8584,N_8468);
nor U9415 (N_9415,N_8274,N_8163);
and U9416 (N_9416,N_8784,N_8710);
and U9417 (N_9417,N_8904,N_7639);
or U9418 (N_9418,N_8829,N_8234);
or U9419 (N_9419,N_7824,N_8674);
nor U9420 (N_9420,N_7782,N_7569);
nand U9421 (N_9421,N_8432,N_8099);
and U9422 (N_9422,N_8987,N_8726);
or U9423 (N_9423,N_7666,N_8360);
or U9424 (N_9424,N_8648,N_8118);
nand U9425 (N_9425,N_8213,N_8105);
and U9426 (N_9426,N_8522,N_7852);
or U9427 (N_9427,N_8220,N_8128);
nor U9428 (N_9428,N_8108,N_8960);
nand U9429 (N_9429,N_8066,N_7934);
nand U9430 (N_9430,N_7943,N_7802);
and U9431 (N_9431,N_7627,N_8183);
or U9432 (N_9432,N_8746,N_7679);
nor U9433 (N_9433,N_8640,N_8555);
nand U9434 (N_9434,N_8033,N_8694);
nand U9435 (N_9435,N_8603,N_7828);
and U9436 (N_9436,N_8478,N_7609);
or U9437 (N_9437,N_8159,N_8614);
nor U9438 (N_9438,N_7971,N_8513);
and U9439 (N_9439,N_8955,N_8704);
and U9440 (N_9440,N_7597,N_8938);
xnor U9441 (N_9441,N_8645,N_7539);
nor U9442 (N_9442,N_7578,N_8956);
nand U9443 (N_9443,N_8810,N_7827);
nand U9444 (N_9444,N_8001,N_8142);
xor U9445 (N_9445,N_8323,N_8181);
and U9446 (N_9446,N_8433,N_7999);
or U9447 (N_9447,N_8019,N_8707);
nand U9448 (N_9448,N_8057,N_7723);
and U9449 (N_9449,N_8326,N_8656);
nand U9450 (N_9450,N_8582,N_7975);
nor U9451 (N_9451,N_8387,N_8409);
or U9452 (N_9452,N_7814,N_8393);
nor U9453 (N_9453,N_7547,N_8677);
xor U9454 (N_9454,N_7976,N_8435);
and U9455 (N_9455,N_8575,N_8310);
nor U9456 (N_9456,N_7642,N_8787);
and U9457 (N_9457,N_7550,N_8053);
or U9458 (N_9458,N_8272,N_8495);
and U9459 (N_9459,N_7594,N_7521);
nor U9460 (N_9460,N_8470,N_8453);
nand U9461 (N_9461,N_7545,N_8668);
nand U9462 (N_9462,N_7863,N_8547);
nor U9463 (N_9463,N_8669,N_8304);
nand U9464 (N_9464,N_7617,N_8693);
and U9465 (N_9465,N_7989,N_7978);
nand U9466 (N_9466,N_7903,N_8971);
or U9467 (N_9467,N_7676,N_8906);
or U9468 (N_9468,N_8192,N_8398);
nor U9469 (N_9469,N_8042,N_8251);
nand U9470 (N_9470,N_7702,N_8655);
xor U9471 (N_9471,N_8256,N_8088);
nor U9472 (N_9472,N_8059,N_8475);
xor U9473 (N_9473,N_8010,N_7742);
or U9474 (N_9474,N_8249,N_8807);
or U9475 (N_9475,N_8041,N_8523);
and U9476 (N_9476,N_7649,N_8317);
and U9477 (N_9477,N_7985,N_8961);
nand U9478 (N_9478,N_8572,N_8739);
nor U9479 (N_9479,N_7719,N_8229);
or U9480 (N_9480,N_8731,N_8964);
xnor U9481 (N_9481,N_8771,N_8858);
and U9482 (N_9482,N_7697,N_8315);
and U9483 (N_9483,N_8032,N_8646);
nand U9484 (N_9484,N_7997,N_8083);
and U9485 (N_9485,N_7935,N_8981);
nor U9486 (N_9486,N_7819,N_8273);
nand U9487 (N_9487,N_8780,N_7769);
and U9488 (N_9488,N_8415,N_8500);
and U9489 (N_9489,N_8253,N_7846);
xnor U9490 (N_9490,N_8895,N_8044);
xor U9491 (N_9491,N_8391,N_7778);
nor U9492 (N_9492,N_8528,N_7566);
nand U9493 (N_9493,N_8927,N_7967);
and U9494 (N_9494,N_7768,N_7799);
xor U9495 (N_9495,N_8977,N_8149);
nand U9496 (N_9496,N_8488,N_8342);
or U9497 (N_9497,N_8456,N_7726);
and U9498 (N_9498,N_8348,N_7559);
nor U9499 (N_9499,N_8006,N_7544);
or U9500 (N_9500,N_8884,N_8670);
or U9501 (N_9501,N_7586,N_8084);
nand U9502 (N_9502,N_7876,N_7541);
nor U9503 (N_9503,N_7601,N_8082);
and U9504 (N_9504,N_7839,N_7655);
or U9505 (N_9505,N_7596,N_8862);
xor U9506 (N_9506,N_8542,N_8319);
nand U9507 (N_9507,N_7672,N_8622);
nand U9508 (N_9508,N_7570,N_8430);
nor U9509 (N_9509,N_8833,N_7800);
or U9510 (N_9510,N_8606,N_7785);
and U9511 (N_9511,N_8246,N_7641);
nor U9512 (N_9512,N_8749,N_7696);
and U9513 (N_9513,N_8508,N_8639);
and U9514 (N_9514,N_8355,N_8386);
nor U9515 (N_9515,N_8607,N_7881);
or U9516 (N_9516,N_7503,N_7677);
nor U9517 (N_9517,N_8208,N_8467);
nand U9518 (N_9518,N_8464,N_8864);
xnor U9519 (N_9519,N_7631,N_8611);
nor U9520 (N_9520,N_8636,N_7517);
xnor U9521 (N_9521,N_8485,N_7671);
nand U9522 (N_9522,N_8717,N_8849);
nand U9523 (N_9523,N_8212,N_8854);
xnor U9524 (N_9524,N_7610,N_8452);
and U9525 (N_9525,N_7536,N_8773);
nor U9526 (N_9526,N_7869,N_8175);
nor U9527 (N_9527,N_8725,N_8332);
nor U9528 (N_9528,N_8565,N_8392);
and U9529 (N_9529,N_8588,N_8349);
nor U9530 (N_9530,N_8700,N_7580);
and U9531 (N_9531,N_7630,N_8135);
or U9532 (N_9532,N_8861,N_7608);
nor U9533 (N_9533,N_8743,N_8153);
nand U9534 (N_9534,N_7789,N_8306);
and U9535 (N_9535,N_8519,N_8087);
nor U9536 (N_9536,N_8608,N_7945);
xor U9537 (N_9537,N_8410,N_8225);
and U9538 (N_9538,N_7534,N_8368);
nor U9539 (N_9539,N_8155,N_7620);
nor U9540 (N_9540,N_8106,N_8015);
nor U9541 (N_9541,N_8164,N_8482);
and U9542 (N_9542,N_8869,N_8484);
nand U9543 (N_9543,N_7969,N_8491);
or U9544 (N_9544,N_7933,N_8583);
or U9545 (N_9545,N_8576,N_8766);
nand U9546 (N_9546,N_7748,N_8817);
and U9547 (N_9547,N_8120,N_8146);
nor U9548 (N_9548,N_7741,N_7908);
or U9549 (N_9549,N_8343,N_7583);
nand U9550 (N_9550,N_8496,N_8612);
nor U9551 (N_9551,N_7940,N_8792);
nor U9552 (N_9552,N_7684,N_7873);
nor U9553 (N_9553,N_8115,N_8573);
nor U9554 (N_9554,N_8826,N_8521);
or U9555 (N_9555,N_7552,N_7651);
nand U9556 (N_9556,N_8367,N_7722);
xor U9557 (N_9557,N_8162,N_7894);
and U9558 (N_9558,N_8434,N_8735);
and U9559 (N_9559,N_8511,N_8423);
and U9560 (N_9560,N_8585,N_7920);
nand U9561 (N_9561,N_7615,N_8760);
nand U9562 (N_9562,N_8844,N_8190);
or U9563 (N_9563,N_7957,N_7598);
nor U9564 (N_9564,N_7657,N_7808);
and U9565 (N_9565,N_8510,N_8951);
or U9566 (N_9566,N_8457,N_8579);
and U9567 (N_9567,N_7508,N_7988);
or U9568 (N_9568,N_8151,N_7803);
nor U9569 (N_9569,N_7717,N_8558);
xnor U9570 (N_9570,N_7893,N_7635);
nand U9571 (N_9571,N_8233,N_8091);
nor U9572 (N_9572,N_7613,N_8713);
xnor U9573 (N_9573,N_8191,N_8184);
nor U9574 (N_9574,N_8917,N_8501);
and U9575 (N_9575,N_8299,N_8751);
and U9576 (N_9576,N_8085,N_7760);
or U9577 (N_9577,N_7850,N_7890);
or U9578 (N_9578,N_7859,N_8417);
nand U9579 (N_9579,N_8894,N_7532);
or U9580 (N_9580,N_8819,N_7542);
nor U9581 (N_9581,N_8756,N_7695);
or U9582 (N_9582,N_8295,N_7919);
xnor U9583 (N_9583,N_8487,N_8407);
nand U9584 (N_9584,N_8992,N_8166);
nand U9585 (N_9585,N_8855,N_7870);
nor U9586 (N_9586,N_8449,N_7813);
nand U9587 (N_9587,N_8063,N_8970);
nand U9588 (N_9588,N_8876,N_8008);
nand U9589 (N_9589,N_7523,N_8280);
or U9590 (N_9590,N_8460,N_8401);
and U9591 (N_9591,N_8131,N_8514);
or U9592 (N_9592,N_8795,N_8629);
nand U9593 (N_9593,N_8590,N_8390);
nand U9594 (N_9594,N_8357,N_8539);
and U9595 (N_9595,N_8916,N_8593);
and U9596 (N_9596,N_8060,N_7721);
or U9597 (N_9597,N_7937,N_8483);
or U9598 (N_9598,N_7528,N_8932);
xor U9599 (N_9599,N_8312,N_7576);
or U9600 (N_9600,N_7885,N_8048);
nor U9601 (N_9601,N_7899,N_7910);
or U9602 (N_9602,N_7950,N_7764);
and U9603 (N_9603,N_8025,N_8450);
or U9604 (N_9604,N_7955,N_7645);
nand U9605 (N_9605,N_8768,N_8958);
nor U9606 (N_9606,N_8170,N_7603);
nand U9607 (N_9607,N_7980,N_8017);
or U9608 (N_9608,N_8701,N_8294);
or U9609 (N_9609,N_8875,N_8952);
or U9610 (N_9610,N_7773,N_7618);
nor U9611 (N_9611,N_7571,N_8383);
nor U9612 (N_9612,N_8426,N_8702);
or U9613 (N_9613,N_8148,N_8405);
nand U9614 (N_9614,N_8898,N_8132);
nor U9615 (N_9615,N_8786,N_8776);
and U9616 (N_9616,N_8365,N_7704);
and U9617 (N_9617,N_8098,N_8757);
or U9618 (N_9618,N_8729,N_8962);
or U9619 (N_9619,N_8658,N_7939);
xor U9620 (N_9620,N_7862,N_7791);
or U9621 (N_9621,N_8913,N_7512);
and U9622 (N_9622,N_8419,N_7991);
or U9623 (N_9623,N_7650,N_8296);
nand U9624 (N_9624,N_8130,N_7879);
nand U9625 (N_9625,N_8691,N_7602);
nand U9626 (N_9626,N_7775,N_8378);
and U9627 (N_9627,N_8744,N_7954);
and U9628 (N_9628,N_8651,N_7924);
and U9629 (N_9629,N_8986,N_7947);
nand U9630 (N_9630,N_8866,N_7759);
and U9631 (N_9631,N_8493,N_8311);
nand U9632 (N_9632,N_8734,N_8366);
nand U9633 (N_9633,N_8741,N_8065);
or U9634 (N_9634,N_8285,N_8728);
nor U9635 (N_9635,N_7733,N_8141);
xor U9636 (N_9636,N_8814,N_8893);
xor U9637 (N_9637,N_8630,N_8111);
xnor U9638 (N_9638,N_8379,N_8140);
or U9639 (N_9639,N_8356,N_7690);
and U9640 (N_9640,N_8079,N_8145);
nor U9641 (N_9641,N_7788,N_7582);
and U9642 (N_9642,N_8254,N_7949);
or U9643 (N_9643,N_7628,N_8755);
and U9644 (N_9644,N_8293,N_8874);
and U9645 (N_9645,N_8339,N_7509);
and U9646 (N_9646,N_8695,N_8122);
and U9647 (N_9647,N_8679,N_8712);
nor U9648 (N_9648,N_7738,N_8777);
xnor U9649 (N_9649,N_8965,N_8995);
xnor U9650 (N_9650,N_8812,N_8219);
nand U9651 (N_9651,N_8202,N_8038);
nand U9652 (N_9652,N_7612,N_8937);
nor U9653 (N_9653,N_7533,N_8696);
nor U9654 (N_9654,N_8134,N_8301);
nor U9655 (N_9655,N_8979,N_8176);
nand U9656 (N_9656,N_8860,N_8998);
nand U9657 (N_9657,N_8402,N_7707);
nand U9658 (N_9658,N_8867,N_7829);
and U9659 (N_9659,N_8942,N_7986);
and U9660 (N_9660,N_8380,N_7761);
nor U9661 (N_9661,N_8461,N_7882);
or U9662 (N_9662,N_8947,N_7906);
and U9663 (N_9663,N_8004,N_8092);
xnor U9664 (N_9664,N_7811,N_8137);
nand U9665 (N_9665,N_8813,N_7548);
and U9666 (N_9666,N_8633,N_8447);
nand U9667 (N_9667,N_8560,N_7670);
xnor U9668 (N_9668,N_7740,N_7794);
nand U9669 (N_9669,N_8077,N_7927);
or U9670 (N_9670,N_8954,N_8879);
xor U9671 (N_9671,N_8637,N_8321);
or U9672 (N_9672,N_7887,N_7660);
xor U9673 (N_9673,N_7743,N_8692);
or U9674 (N_9674,N_7573,N_7757);
nand U9675 (N_9675,N_8770,N_8742);
nand U9676 (N_9676,N_8925,N_8281);
or U9677 (N_9677,N_8665,N_8613);
or U9678 (N_9678,N_8055,N_8525);
and U9679 (N_9679,N_8914,N_7842);
nand U9680 (N_9680,N_8313,N_8374);
or U9681 (N_9681,N_8578,N_8774);
or U9682 (N_9682,N_8027,N_8627);
nor U9683 (N_9683,N_8095,N_7815);
xnor U9684 (N_9684,N_8873,N_8143);
xnor U9685 (N_9685,N_8199,N_7946);
nand U9686 (N_9686,N_8298,N_8472);
nand U9687 (N_9687,N_7504,N_8901);
nand U9688 (N_9688,N_7836,N_8072);
nor U9689 (N_9689,N_8845,N_8473);
xnor U9690 (N_9690,N_8018,N_8104);
and U9691 (N_9691,N_8171,N_8049);
nor U9692 (N_9692,N_8476,N_7754);
and U9693 (N_9693,N_8455,N_7916);
nand U9694 (N_9694,N_8463,N_7838);
nand U9695 (N_9695,N_7826,N_8307);
and U9696 (N_9696,N_7812,N_7589);
nor U9697 (N_9697,N_8382,N_7555);
and U9698 (N_9698,N_8919,N_8765);
nor U9699 (N_9699,N_8000,N_8248);
nor U9700 (N_9700,N_7538,N_8337);
nor U9701 (N_9701,N_8230,N_8672);
nor U9702 (N_9702,N_7979,N_7674);
nand U9703 (N_9703,N_8949,N_8037);
nor U9704 (N_9704,N_8626,N_7849);
nor U9705 (N_9705,N_8892,N_8847);
nand U9706 (N_9706,N_8034,N_8147);
nor U9707 (N_9707,N_8477,N_8394);
nand U9708 (N_9708,N_8003,N_7765);
nand U9709 (N_9709,N_8821,N_8905);
and U9710 (N_9710,N_8028,N_7561);
and U9711 (N_9711,N_8350,N_7624);
nor U9712 (N_9712,N_8708,N_8466);
nand U9713 (N_9713,N_7995,N_8870);
nor U9714 (N_9714,N_7983,N_8445);
and U9715 (N_9715,N_8732,N_8595);
or U9716 (N_9716,N_8431,N_8309);
nand U9717 (N_9717,N_8324,N_8119);
nor U9718 (N_9718,N_7928,N_8553);
nor U9719 (N_9719,N_8680,N_8189);
or U9720 (N_9720,N_7746,N_8924);
xor U9721 (N_9721,N_7698,N_8678);
xor U9722 (N_9722,N_8871,N_7518);
nor U9723 (N_9723,N_8458,N_8052);
or U9724 (N_9724,N_7973,N_7600);
xor U9725 (N_9725,N_8494,N_8556);
and U9726 (N_9726,N_7640,N_8684);
nor U9727 (N_9727,N_8036,N_8174);
and U9728 (N_9728,N_8681,N_8370);
and U9729 (N_9729,N_7653,N_8232);
or U9730 (N_9730,N_8599,N_8173);
or U9731 (N_9731,N_8559,N_7705);
or U9732 (N_9732,N_7798,N_8809);
or U9733 (N_9733,N_8834,N_8222);
nor U9734 (N_9734,N_8308,N_8531);
or U9735 (N_9735,N_8838,N_8292);
nand U9736 (N_9736,N_8113,N_8359);
nor U9737 (N_9737,N_7526,N_8936);
or U9738 (N_9738,N_8030,N_8657);
or U9739 (N_9739,N_8617,N_8846);
and U9740 (N_9740,N_8502,N_7590);
nor U9741 (N_9741,N_8238,N_7905);
nor U9742 (N_9742,N_8975,N_8567);
nand U9743 (N_9743,N_8318,N_7847);
and U9744 (N_9744,N_7762,N_7701);
or U9745 (N_9745,N_8520,N_8211);
and U9746 (N_9746,N_8013,N_8201);
and U9747 (N_9747,N_8610,N_8516);
or U9748 (N_9748,N_7720,N_8330);
and U9749 (N_9749,N_8172,N_8733);
nor U9750 (N_9750,N_8147,N_8954);
nor U9751 (N_9751,N_8344,N_8625);
xor U9752 (N_9752,N_8554,N_8460);
nor U9753 (N_9753,N_8267,N_8982);
nand U9754 (N_9754,N_7946,N_8669);
and U9755 (N_9755,N_8431,N_7661);
nand U9756 (N_9756,N_7703,N_8488);
nand U9757 (N_9757,N_7820,N_8101);
nor U9758 (N_9758,N_7994,N_8038);
xor U9759 (N_9759,N_7923,N_8567);
nor U9760 (N_9760,N_7696,N_7621);
or U9761 (N_9761,N_8354,N_8477);
or U9762 (N_9762,N_7513,N_8100);
nor U9763 (N_9763,N_7902,N_7888);
and U9764 (N_9764,N_8698,N_8845);
nand U9765 (N_9765,N_7617,N_7641);
or U9766 (N_9766,N_7930,N_8449);
nand U9767 (N_9767,N_7542,N_8165);
or U9768 (N_9768,N_7674,N_7779);
xnor U9769 (N_9769,N_8305,N_8934);
or U9770 (N_9770,N_7962,N_8145);
and U9771 (N_9771,N_7939,N_7652);
nand U9772 (N_9772,N_7749,N_7807);
nand U9773 (N_9773,N_7862,N_7926);
xor U9774 (N_9774,N_7513,N_8156);
nor U9775 (N_9775,N_8678,N_8903);
or U9776 (N_9776,N_8106,N_7568);
nand U9777 (N_9777,N_8710,N_7752);
or U9778 (N_9778,N_8177,N_8868);
nand U9779 (N_9779,N_7642,N_8225);
and U9780 (N_9780,N_8341,N_8055);
or U9781 (N_9781,N_7848,N_7758);
nand U9782 (N_9782,N_8131,N_7723);
and U9783 (N_9783,N_8806,N_8413);
nor U9784 (N_9784,N_7848,N_8589);
xnor U9785 (N_9785,N_7781,N_8662);
nor U9786 (N_9786,N_8015,N_8156);
or U9787 (N_9787,N_7926,N_8234);
nand U9788 (N_9788,N_7783,N_8018);
and U9789 (N_9789,N_8538,N_8502);
and U9790 (N_9790,N_8570,N_8358);
and U9791 (N_9791,N_8200,N_8747);
or U9792 (N_9792,N_8056,N_8680);
xnor U9793 (N_9793,N_8256,N_8536);
nor U9794 (N_9794,N_8284,N_8356);
nand U9795 (N_9795,N_8346,N_7903);
nand U9796 (N_9796,N_8951,N_8180);
nand U9797 (N_9797,N_8410,N_8240);
xnor U9798 (N_9798,N_7741,N_8578);
or U9799 (N_9799,N_8772,N_8200);
nor U9800 (N_9800,N_7858,N_8329);
and U9801 (N_9801,N_8902,N_8995);
nor U9802 (N_9802,N_8902,N_8473);
nor U9803 (N_9803,N_8675,N_8788);
and U9804 (N_9804,N_8032,N_8457);
nand U9805 (N_9805,N_8486,N_7989);
xor U9806 (N_9806,N_8409,N_8499);
nand U9807 (N_9807,N_7707,N_8197);
or U9808 (N_9808,N_8075,N_8932);
or U9809 (N_9809,N_8867,N_8856);
nor U9810 (N_9810,N_8630,N_7941);
and U9811 (N_9811,N_8280,N_8391);
or U9812 (N_9812,N_8137,N_8124);
and U9813 (N_9813,N_7699,N_7508);
or U9814 (N_9814,N_8055,N_7803);
nand U9815 (N_9815,N_8169,N_8226);
xnor U9816 (N_9816,N_8571,N_8539);
nor U9817 (N_9817,N_8570,N_7552);
or U9818 (N_9818,N_7595,N_7836);
nand U9819 (N_9819,N_8360,N_8305);
nor U9820 (N_9820,N_7878,N_7543);
nand U9821 (N_9821,N_8101,N_7994);
or U9822 (N_9822,N_7969,N_7973);
and U9823 (N_9823,N_7544,N_8877);
or U9824 (N_9824,N_7592,N_8409);
xor U9825 (N_9825,N_8938,N_8155);
and U9826 (N_9826,N_8195,N_8257);
nor U9827 (N_9827,N_7502,N_8200);
or U9828 (N_9828,N_8134,N_8059);
nand U9829 (N_9829,N_8026,N_8879);
nand U9830 (N_9830,N_7577,N_8738);
and U9831 (N_9831,N_7719,N_8349);
nor U9832 (N_9832,N_7518,N_7814);
and U9833 (N_9833,N_7872,N_8365);
nor U9834 (N_9834,N_7550,N_8920);
nand U9835 (N_9835,N_7679,N_8305);
and U9836 (N_9836,N_7881,N_8967);
or U9837 (N_9837,N_7745,N_8772);
nor U9838 (N_9838,N_7634,N_7810);
xor U9839 (N_9839,N_8953,N_8198);
or U9840 (N_9840,N_7836,N_8453);
nand U9841 (N_9841,N_8735,N_8554);
and U9842 (N_9842,N_7836,N_8269);
nor U9843 (N_9843,N_8792,N_8504);
nand U9844 (N_9844,N_8020,N_8362);
nor U9845 (N_9845,N_8862,N_7932);
nor U9846 (N_9846,N_8316,N_7531);
nand U9847 (N_9847,N_8179,N_7987);
nand U9848 (N_9848,N_8091,N_8744);
nand U9849 (N_9849,N_7683,N_7547);
nand U9850 (N_9850,N_8778,N_8148);
or U9851 (N_9851,N_8815,N_7583);
or U9852 (N_9852,N_8201,N_8325);
nand U9853 (N_9853,N_8377,N_7558);
nor U9854 (N_9854,N_7588,N_8941);
xnor U9855 (N_9855,N_8701,N_8213);
or U9856 (N_9856,N_7694,N_7901);
nor U9857 (N_9857,N_7658,N_8293);
and U9858 (N_9858,N_8284,N_8403);
and U9859 (N_9859,N_8676,N_7762);
or U9860 (N_9860,N_7578,N_8090);
and U9861 (N_9861,N_7993,N_8575);
nor U9862 (N_9862,N_8800,N_8759);
and U9863 (N_9863,N_8587,N_8181);
nor U9864 (N_9864,N_8115,N_8228);
nor U9865 (N_9865,N_7902,N_8425);
xnor U9866 (N_9866,N_8916,N_8410);
nand U9867 (N_9867,N_7638,N_8409);
nand U9868 (N_9868,N_8020,N_7731);
or U9869 (N_9869,N_8319,N_8070);
and U9870 (N_9870,N_8418,N_8261);
or U9871 (N_9871,N_8589,N_8672);
nor U9872 (N_9872,N_8189,N_7662);
or U9873 (N_9873,N_7632,N_8473);
and U9874 (N_9874,N_8210,N_8995);
xnor U9875 (N_9875,N_8077,N_7603);
and U9876 (N_9876,N_7624,N_7956);
and U9877 (N_9877,N_8284,N_7717);
or U9878 (N_9878,N_7583,N_7732);
or U9879 (N_9879,N_7629,N_7878);
nand U9880 (N_9880,N_7958,N_7941);
and U9881 (N_9881,N_8218,N_8032);
nand U9882 (N_9882,N_7637,N_8454);
or U9883 (N_9883,N_8458,N_8639);
nand U9884 (N_9884,N_8483,N_7815);
or U9885 (N_9885,N_7543,N_8889);
nor U9886 (N_9886,N_7574,N_8150);
xor U9887 (N_9887,N_8677,N_8312);
nor U9888 (N_9888,N_8987,N_7586);
and U9889 (N_9889,N_7766,N_8203);
nor U9890 (N_9890,N_8666,N_7999);
nand U9891 (N_9891,N_8951,N_7518);
nand U9892 (N_9892,N_8144,N_8026);
nand U9893 (N_9893,N_8530,N_8222);
and U9894 (N_9894,N_8458,N_8335);
nor U9895 (N_9895,N_8076,N_8716);
nor U9896 (N_9896,N_8066,N_7546);
and U9897 (N_9897,N_8785,N_8754);
nor U9898 (N_9898,N_8512,N_7900);
and U9899 (N_9899,N_8951,N_8093);
and U9900 (N_9900,N_7684,N_7835);
or U9901 (N_9901,N_8702,N_8411);
or U9902 (N_9902,N_7549,N_8492);
nand U9903 (N_9903,N_8420,N_8316);
or U9904 (N_9904,N_8279,N_7516);
nand U9905 (N_9905,N_8523,N_7754);
xor U9906 (N_9906,N_7719,N_8514);
nand U9907 (N_9907,N_8042,N_8285);
and U9908 (N_9908,N_8344,N_7566);
xor U9909 (N_9909,N_7600,N_8587);
xor U9910 (N_9910,N_8417,N_8056);
nand U9911 (N_9911,N_7844,N_7839);
or U9912 (N_9912,N_8083,N_8637);
and U9913 (N_9913,N_8068,N_7524);
nand U9914 (N_9914,N_7840,N_7747);
or U9915 (N_9915,N_7925,N_8070);
or U9916 (N_9916,N_8895,N_7875);
nand U9917 (N_9917,N_8021,N_7897);
or U9918 (N_9918,N_8433,N_8235);
nor U9919 (N_9919,N_8640,N_8997);
and U9920 (N_9920,N_7614,N_7892);
and U9921 (N_9921,N_7565,N_8327);
nand U9922 (N_9922,N_8825,N_7690);
xor U9923 (N_9923,N_8768,N_7995);
nand U9924 (N_9924,N_8955,N_7748);
or U9925 (N_9925,N_8417,N_8000);
nor U9926 (N_9926,N_7608,N_8448);
xor U9927 (N_9927,N_8968,N_8123);
nand U9928 (N_9928,N_8857,N_8144);
nor U9929 (N_9929,N_8646,N_8114);
nand U9930 (N_9930,N_8953,N_7885);
and U9931 (N_9931,N_8894,N_7874);
nor U9932 (N_9932,N_8772,N_8321);
nand U9933 (N_9933,N_7990,N_8167);
xnor U9934 (N_9934,N_8131,N_8798);
and U9935 (N_9935,N_8347,N_8315);
nand U9936 (N_9936,N_8191,N_8666);
and U9937 (N_9937,N_8217,N_8884);
nand U9938 (N_9938,N_8321,N_7646);
nor U9939 (N_9939,N_8738,N_8077);
and U9940 (N_9940,N_7743,N_8502);
and U9941 (N_9941,N_8278,N_8118);
nor U9942 (N_9942,N_8203,N_8348);
or U9943 (N_9943,N_8969,N_8048);
and U9944 (N_9944,N_7774,N_8430);
nor U9945 (N_9945,N_7541,N_7597);
and U9946 (N_9946,N_8741,N_8865);
nor U9947 (N_9947,N_8682,N_8180);
nand U9948 (N_9948,N_8016,N_8408);
nand U9949 (N_9949,N_8234,N_8037);
and U9950 (N_9950,N_8986,N_7905);
nor U9951 (N_9951,N_7735,N_8001);
nor U9952 (N_9952,N_8653,N_8392);
and U9953 (N_9953,N_8927,N_8390);
nor U9954 (N_9954,N_8144,N_8619);
and U9955 (N_9955,N_8198,N_8373);
nor U9956 (N_9956,N_7956,N_8578);
nor U9957 (N_9957,N_7891,N_8468);
or U9958 (N_9958,N_8562,N_7513);
xnor U9959 (N_9959,N_7969,N_7767);
nor U9960 (N_9960,N_8817,N_8634);
nor U9961 (N_9961,N_8668,N_8264);
nand U9962 (N_9962,N_8217,N_8603);
or U9963 (N_9963,N_8437,N_7683);
nor U9964 (N_9964,N_8243,N_7628);
and U9965 (N_9965,N_7540,N_7554);
and U9966 (N_9966,N_7945,N_8786);
and U9967 (N_9967,N_8882,N_8217);
and U9968 (N_9968,N_7916,N_7609);
xor U9969 (N_9969,N_8297,N_8625);
nand U9970 (N_9970,N_7784,N_7693);
xnor U9971 (N_9971,N_7991,N_8944);
nand U9972 (N_9972,N_7797,N_8208);
nor U9973 (N_9973,N_7972,N_8748);
xor U9974 (N_9974,N_8938,N_7604);
nand U9975 (N_9975,N_8696,N_8298);
nand U9976 (N_9976,N_7941,N_7597);
or U9977 (N_9977,N_8110,N_8349);
and U9978 (N_9978,N_8370,N_7894);
xor U9979 (N_9979,N_8229,N_8614);
and U9980 (N_9980,N_7630,N_8097);
xnor U9981 (N_9981,N_8346,N_7950);
nand U9982 (N_9982,N_8509,N_8052);
nor U9983 (N_9983,N_8080,N_8467);
nand U9984 (N_9984,N_8037,N_8963);
or U9985 (N_9985,N_8605,N_8813);
or U9986 (N_9986,N_7966,N_7815);
nand U9987 (N_9987,N_8972,N_7885);
xor U9988 (N_9988,N_7748,N_8626);
and U9989 (N_9989,N_7526,N_7599);
xor U9990 (N_9990,N_8403,N_7785);
or U9991 (N_9991,N_7585,N_8632);
or U9992 (N_9992,N_8589,N_8952);
nor U9993 (N_9993,N_7927,N_7665);
xor U9994 (N_9994,N_8719,N_7534);
nand U9995 (N_9995,N_8387,N_8328);
nor U9996 (N_9996,N_8953,N_8893);
nand U9997 (N_9997,N_7572,N_7714);
and U9998 (N_9998,N_7520,N_8663);
or U9999 (N_9999,N_8176,N_7696);
and U10000 (N_10000,N_8587,N_8004);
and U10001 (N_10001,N_8931,N_8216);
and U10002 (N_10002,N_8278,N_7829);
and U10003 (N_10003,N_8900,N_7810);
xnor U10004 (N_10004,N_8212,N_8118);
nor U10005 (N_10005,N_7742,N_8745);
nor U10006 (N_10006,N_8645,N_7843);
nor U10007 (N_10007,N_7802,N_8189);
nand U10008 (N_10008,N_8620,N_8530);
or U10009 (N_10009,N_7503,N_7622);
or U10010 (N_10010,N_8561,N_8122);
nor U10011 (N_10011,N_8769,N_7509);
nor U10012 (N_10012,N_8537,N_8729);
and U10013 (N_10013,N_8014,N_7801);
nor U10014 (N_10014,N_8557,N_8190);
nand U10015 (N_10015,N_7748,N_7653);
nand U10016 (N_10016,N_7635,N_7920);
xnor U10017 (N_10017,N_8914,N_7592);
xor U10018 (N_10018,N_8488,N_8430);
nand U10019 (N_10019,N_8381,N_8012);
or U10020 (N_10020,N_8960,N_8538);
or U10021 (N_10021,N_8792,N_7887);
nor U10022 (N_10022,N_8594,N_8379);
or U10023 (N_10023,N_8087,N_8131);
or U10024 (N_10024,N_8681,N_7650);
and U10025 (N_10025,N_7766,N_8207);
or U10026 (N_10026,N_7590,N_8960);
nor U10027 (N_10027,N_7983,N_8785);
nand U10028 (N_10028,N_8950,N_8472);
xor U10029 (N_10029,N_8623,N_7894);
and U10030 (N_10030,N_7523,N_8285);
nor U10031 (N_10031,N_7730,N_8965);
nor U10032 (N_10032,N_8040,N_8415);
xnor U10033 (N_10033,N_8503,N_8932);
nor U10034 (N_10034,N_8076,N_8203);
and U10035 (N_10035,N_7524,N_7607);
xor U10036 (N_10036,N_8752,N_7671);
and U10037 (N_10037,N_7850,N_8605);
and U10038 (N_10038,N_7973,N_8934);
and U10039 (N_10039,N_8476,N_7834);
nand U10040 (N_10040,N_7580,N_8979);
nor U10041 (N_10041,N_8491,N_7869);
or U10042 (N_10042,N_8783,N_7644);
nor U10043 (N_10043,N_8004,N_7956);
nand U10044 (N_10044,N_8123,N_7583);
nand U10045 (N_10045,N_8131,N_8588);
nand U10046 (N_10046,N_8390,N_7852);
nand U10047 (N_10047,N_8509,N_8316);
xnor U10048 (N_10048,N_8433,N_8808);
and U10049 (N_10049,N_8593,N_8308);
and U10050 (N_10050,N_8128,N_8021);
nand U10051 (N_10051,N_8110,N_7918);
nand U10052 (N_10052,N_8743,N_7669);
and U10053 (N_10053,N_7619,N_7856);
xor U10054 (N_10054,N_7527,N_8796);
and U10055 (N_10055,N_7540,N_7530);
or U10056 (N_10056,N_8488,N_8978);
or U10057 (N_10057,N_8785,N_8452);
nor U10058 (N_10058,N_8422,N_8939);
xor U10059 (N_10059,N_8502,N_8664);
or U10060 (N_10060,N_7868,N_8371);
xnor U10061 (N_10061,N_7582,N_8631);
nand U10062 (N_10062,N_8684,N_8087);
and U10063 (N_10063,N_8388,N_8825);
nor U10064 (N_10064,N_7912,N_7705);
or U10065 (N_10065,N_8898,N_8775);
and U10066 (N_10066,N_7567,N_7716);
nor U10067 (N_10067,N_8687,N_8377);
and U10068 (N_10068,N_7587,N_8207);
xnor U10069 (N_10069,N_8020,N_8082);
xnor U10070 (N_10070,N_8149,N_7614);
nand U10071 (N_10071,N_8031,N_7546);
nand U10072 (N_10072,N_7781,N_7938);
nand U10073 (N_10073,N_8371,N_8301);
and U10074 (N_10074,N_8100,N_8931);
or U10075 (N_10075,N_8477,N_8398);
or U10076 (N_10076,N_8464,N_8093);
and U10077 (N_10077,N_8489,N_8379);
nor U10078 (N_10078,N_8734,N_7612);
and U10079 (N_10079,N_8886,N_7545);
and U10080 (N_10080,N_7954,N_8789);
nor U10081 (N_10081,N_8241,N_8660);
nand U10082 (N_10082,N_8380,N_8236);
or U10083 (N_10083,N_7657,N_7627);
nor U10084 (N_10084,N_8605,N_8121);
nand U10085 (N_10085,N_8696,N_8428);
nand U10086 (N_10086,N_7731,N_8432);
nor U10087 (N_10087,N_7550,N_8612);
or U10088 (N_10088,N_7933,N_8897);
and U10089 (N_10089,N_8926,N_8802);
or U10090 (N_10090,N_8964,N_8990);
nand U10091 (N_10091,N_8785,N_8990);
nand U10092 (N_10092,N_8961,N_8198);
and U10093 (N_10093,N_8793,N_8925);
nand U10094 (N_10094,N_8756,N_8883);
nor U10095 (N_10095,N_7953,N_8617);
or U10096 (N_10096,N_8389,N_8285);
nor U10097 (N_10097,N_8857,N_8440);
xnor U10098 (N_10098,N_7803,N_8369);
and U10099 (N_10099,N_8249,N_7770);
nand U10100 (N_10100,N_7731,N_8810);
xnor U10101 (N_10101,N_8221,N_8532);
nor U10102 (N_10102,N_8950,N_8487);
or U10103 (N_10103,N_7614,N_8608);
nor U10104 (N_10104,N_8614,N_8781);
nor U10105 (N_10105,N_8432,N_8170);
nor U10106 (N_10106,N_8235,N_7893);
and U10107 (N_10107,N_8804,N_8299);
nor U10108 (N_10108,N_8512,N_8288);
and U10109 (N_10109,N_8616,N_8993);
nor U10110 (N_10110,N_8872,N_7558);
nand U10111 (N_10111,N_8136,N_8120);
xnor U10112 (N_10112,N_7765,N_8284);
nor U10113 (N_10113,N_8541,N_8843);
and U10114 (N_10114,N_8795,N_7584);
and U10115 (N_10115,N_8210,N_8757);
nor U10116 (N_10116,N_7937,N_8980);
xnor U10117 (N_10117,N_8010,N_8065);
nor U10118 (N_10118,N_7942,N_7893);
and U10119 (N_10119,N_7579,N_7922);
and U10120 (N_10120,N_8581,N_8003);
nor U10121 (N_10121,N_8330,N_8275);
or U10122 (N_10122,N_8960,N_8684);
nand U10123 (N_10123,N_8671,N_8644);
nand U10124 (N_10124,N_8550,N_8647);
and U10125 (N_10125,N_7581,N_7886);
or U10126 (N_10126,N_8200,N_8271);
nand U10127 (N_10127,N_8236,N_8233);
xnor U10128 (N_10128,N_8341,N_7691);
nand U10129 (N_10129,N_7681,N_8690);
and U10130 (N_10130,N_7952,N_7818);
nand U10131 (N_10131,N_8826,N_7872);
or U10132 (N_10132,N_7781,N_8100);
or U10133 (N_10133,N_7723,N_8970);
nor U10134 (N_10134,N_7906,N_8972);
nand U10135 (N_10135,N_8266,N_8082);
and U10136 (N_10136,N_8234,N_8435);
nand U10137 (N_10137,N_8007,N_8697);
nand U10138 (N_10138,N_8327,N_8043);
nor U10139 (N_10139,N_8415,N_8930);
nor U10140 (N_10140,N_8404,N_8624);
nor U10141 (N_10141,N_8474,N_8802);
or U10142 (N_10142,N_8725,N_8174);
nor U10143 (N_10143,N_8742,N_7706);
or U10144 (N_10144,N_8507,N_7976);
and U10145 (N_10145,N_8140,N_8637);
nand U10146 (N_10146,N_8886,N_8788);
nand U10147 (N_10147,N_8432,N_8795);
and U10148 (N_10148,N_8038,N_7609);
nand U10149 (N_10149,N_7836,N_7582);
nor U10150 (N_10150,N_8500,N_7932);
and U10151 (N_10151,N_8828,N_7753);
and U10152 (N_10152,N_7595,N_8637);
or U10153 (N_10153,N_7651,N_8284);
nand U10154 (N_10154,N_8113,N_7976);
and U10155 (N_10155,N_7782,N_8375);
xnor U10156 (N_10156,N_8099,N_8526);
or U10157 (N_10157,N_8095,N_7602);
nor U10158 (N_10158,N_8450,N_8993);
and U10159 (N_10159,N_7993,N_8236);
and U10160 (N_10160,N_8470,N_8360);
nor U10161 (N_10161,N_7825,N_8441);
nor U10162 (N_10162,N_8254,N_7718);
nand U10163 (N_10163,N_7818,N_8082);
or U10164 (N_10164,N_8198,N_8138);
nor U10165 (N_10165,N_8071,N_8944);
and U10166 (N_10166,N_8131,N_8856);
and U10167 (N_10167,N_7520,N_8038);
and U10168 (N_10168,N_7790,N_8832);
and U10169 (N_10169,N_7633,N_7745);
and U10170 (N_10170,N_7793,N_8878);
nor U10171 (N_10171,N_8237,N_8882);
nor U10172 (N_10172,N_8671,N_8557);
or U10173 (N_10173,N_8773,N_8350);
nor U10174 (N_10174,N_8351,N_8757);
and U10175 (N_10175,N_7912,N_7776);
nor U10176 (N_10176,N_8879,N_8046);
nand U10177 (N_10177,N_8132,N_7722);
nor U10178 (N_10178,N_8468,N_8330);
xor U10179 (N_10179,N_7922,N_8838);
and U10180 (N_10180,N_8979,N_8446);
nor U10181 (N_10181,N_7875,N_8392);
or U10182 (N_10182,N_8705,N_8609);
nand U10183 (N_10183,N_7972,N_8849);
xor U10184 (N_10184,N_8343,N_7990);
nand U10185 (N_10185,N_7570,N_8969);
nor U10186 (N_10186,N_7534,N_7875);
or U10187 (N_10187,N_7617,N_7866);
nor U10188 (N_10188,N_7686,N_8381);
or U10189 (N_10189,N_7628,N_7585);
or U10190 (N_10190,N_8172,N_8463);
or U10191 (N_10191,N_8979,N_7677);
nor U10192 (N_10192,N_7711,N_7714);
nor U10193 (N_10193,N_8053,N_8559);
xor U10194 (N_10194,N_7557,N_8170);
and U10195 (N_10195,N_8418,N_7676);
xnor U10196 (N_10196,N_7728,N_7956);
and U10197 (N_10197,N_8034,N_7863);
and U10198 (N_10198,N_8598,N_8521);
xnor U10199 (N_10199,N_8928,N_8250);
and U10200 (N_10200,N_8371,N_8772);
or U10201 (N_10201,N_7512,N_8610);
nor U10202 (N_10202,N_8791,N_7964);
nor U10203 (N_10203,N_8402,N_8974);
nor U10204 (N_10204,N_7732,N_7934);
nand U10205 (N_10205,N_8764,N_7842);
xor U10206 (N_10206,N_8464,N_8219);
and U10207 (N_10207,N_8537,N_8528);
or U10208 (N_10208,N_8139,N_8073);
nand U10209 (N_10209,N_8812,N_7721);
nor U10210 (N_10210,N_8886,N_7798);
nand U10211 (N_10211,N_8161,N_8193);
nor U10212 (N_10212,N_8009,N_8870);
nand U10213 (N_10213,N_7950,N_7520);
nand U10214 (N_10214,N_8550,N_8934);
nor U10215 (N_10215,N_7856,N_8798);
or U10216 (N_10216,N_8599,N_8774);
nor U10217 (N_10217,N_8904,N_8108);
or U10218 (N_10218,N_8656,N_7733);
nand U10219 (N_10219,N_7543,N_7873);
and U10220 (N_10220,N_7979,N_8861);
or U10221 (N_10221,N_7619,N_8386);
nand U10222 (N_10222,N_7907,N_7669);
nand U10223 (N_10223,N_8542,N_8954);
and U10224 (N_10224,N_8583,N_8738);
and U10225 (N_10225,N_7518,N_7757);
or U10226 (N_10226,N_8853,N_8144);
and U10227 (N_10227,N_8307,N_8282);
xor U10228 (N_10228,N_7619,N_8427);
nand U10229 (N_10229,N_7868,N_8432);
nand U10230 (N_10230,N_8680,N_7918);
xnor U10231 (N_10231,N_7502,N_8477);
xnor U10232 (N_10232,N_8074,N_7894);
xor U10233 (N_10233,N_8978,N_8045);
nor U10234 (N_10234,N_8246,N_8802);
nor U10235 (N_10235,N_7698,N_8779);
nor U10236 (N_10236,N_8169,N_7995);
and U10237 (N_10237,N_8673,N_8495);
nor U10238 (N_10238,N_8798,N_8489);
nand U10239 (N_10239,N_8722,N_8139);
and U10240 (N_10240,N_7698,N_8957);
or U10241 (N_10241,N_7637,N_8414);
or U10242 (N_10242,N_8873,N_8486);
or U10243 (N_10243,N_8041,N_8984);
nand U10244 (N_10244,N_8609,N_8075);
or U10245 (N_10245,N_8938,N_8520);
and U10246 (N_10246,N_8458,N_8711);
nand U10247 (N_10247,N_7843,N_7920);
nor U10248 (N_10248,N_8933,N_7777);
xnor U10249 (N_10249,N_8529,N_8850);
nand U10250 (N_10250,N_8550,N_8740);
nand U10251 (N_10251,N_8817,N_8022);
nand U10252 (N_10252,N_8833,N_8330);
or U10253 (N_10253,N_7867,N_8896);
nor U10254 (N_10254,N_7912,N_8629);
nor U10255 (N_10255,N_8433,N_8765);
or U10256 (N_10256,N_8774,N_8723);
nand U10257 (N_10257,N_8737,N_8527);
or U10258 (N_10258,N_7568,N_7676);
and U10259 (N_10259,N_8734,N_7506);
xnor U10260 (N_10260,N_8119,N_7532);
or U10261 (N_10261,N_8379,N_8897);
nand U10262 (N_10262,N_8982,N_8146);
or U10263 (N_10263,N_8879,N_8890);
or U10264 (N_10264,N_8508,N_7924);
or U10265 (N_10265,N_7652,N_8213);
or U10266 (N_10266,N_8208,N_8506);
nor U10267 (N_10267,N_7743,N_7656);
and U10268 (N_10268,N_8812,N_7921);
or U10269 (N_10269,N_8594,N_8039);
nand U10270 (N_10270,N_8028,N_8883);
nand U10271 (N_10271,N_8237,N_8746);
xor U10272 (N_10272,N_8801,N_8123);
or U10273 (N_10273,N_7506,N_8409);
xnor U10274 (N_10274,N_8806,N_7754);
and U10275 (N_10275,N_8300,N_7821);
and U10276 (N_10276,N_8569,N_8440);
nor U10277 (N_10277,N_7582,N_7715);
or U10278 (N_10278,N_8559,N_8554);
or U10279 (N_10279,N_7665,N_8699);
nand U10280 (N_10280,N_8804,N_8917);
and U10281 (N_10281,N_7981,N_7577);
nand U10282 (N_10282,N_7554,N_7701);
nor U10283 (N_10283,N_7547,N_7696);
and U10284 (N_10284,N_8139,N_8396);
and U10285 (N_10285,N_8427,N_8147);
nand U10286 (N_10286,N_8379,N_7874);
nor U10287 (N_10287,N_8325,N_8969);
nor U10288 (N_10288,N_8546,N_7504);
nand U10289 (N_10289,N_8683,N_8262);
and U10290 (N_10290,N_7613,N_8193);
xnor U10291 (N_10291,N_7570,N_8762);
nor U10292 (N_10292,N_7967,N_8590);
xor U10293 (N_10293,N_7814,N_8435);
or U10294 (N_10294,N_8830,N_8093);
nand U10295 (N_10295,N_8067,N_7703);
or U10296 (N_10296,N_8969,N_8259);
xnor U10297 (N_10297,N_8722,N_8581);
nor U10298 (N_10298,N_8107,N_8009);
or U10299 (N_10299,N_8116,N_7895);
nand U10300 (N_10300,N_7752,N_8254);
and U10301 (N_10301,N_8460,N_8436);
nor U10302 (N_10302,N_7716,N_8817);
or U10303 (N_10303,N_8325,N_8473);
nand U10304 (N_10304,N_8633,N_8312);
nor U10305 (N_10305,N_8246,N_8094);
or U10306 (N_10306,N_7510,N_7655);
nand U10307 (N_10307,N_8003,N_8297);
or U10308 (N_10308,N_7701,N_7680);
nand U10309 (N_10309,N_7912,N_8467);
and U10310 (N_10310,N_8909,N_8872);
nor U10311 (N_10311,N_8727,N_8009);
or U10312 (N_10312,N_8512,N_8982);
nor U10313 (N_10313,N_7790,N_8551);
or U10314 (N_10314,N_7720,N_8456);
nor U10315 (N_10315,N_8950,N_7714);
and U10316 (N_10316,N_7921,N_8070);
and U10317 (N_10317,N_7659,N_8110);
or U10318 (N_10318,N_8591,N_8529);
nand U10319 (N_10319,N_8902,N_8164);
nor U10320 (N_10320,N_8368,N_8167);
and U10321 (N_10321,N_8360,N_8235);
nand U10322 (N_10322,N_7897,N_7686);
and U10323 (N_10323,N_8492,N_8341);
nor U10324 (N_10324,N_8585,N_7747);
or U10325 (N_10325,N_8253,N_7867);
xor U10326 (N_10326,N_8553,N_8305);
or U10327 (N_10327,N_7889,N_8724);
and U10328 (N_10328,N_8083,N_7562);
or U10329 (N_10329,N_8123,N_8725);
nor U10330 (N_10330,N_8416,N_7980);
nor U10331 (N_10331,N_8075,N_7825);
nand U10332 (N_10332,N_8291,N_7754);
or U10333 (N_10333,N_7910,N_8495);
nand U10334 (N_10334,N_8678,N_7604);
nor U10335 (N_10335,N_8197,N_7511);
nand U10336 (N_10336,N_7652,N_7709);
nand U10337 (N_10337,N_8974,N_7629);
nor U10338 (N_10338,N_7805,N_8098);
and U10339 (N_10339,N_8520,N_8961);
nand U10340 (N_10340,N_8946,N_7923);
nand U10341 (N_10341,N_8996,N_7729);
or U10342 (N_10342,N_7641,N_8974);
or U10343 (N_10343,N_8368,N_8390);
nand U10344 (N_10344,N_8225,N_8347);
nor U10345 (N_10345,N_8351,N_7812);
or U10346 (N_10346,N_7705,N_7893);
or U10347 (N_10347,N_7922,N_8740);
or U10348 (N_10348,N_8296,N_8537);
nand U10349 (N_10349,N_8181,N_8971);
nor U10350 (N_10350,N_8150,N_8192);
and U10351 (N_10351,N_7752,N_7949);
and U10352 (N_10352,N_8767,N_7659);
xnor U10353 (N_10353,N_7924,N_7518);
nor U10354 (N_10354,N_8624,N_7682);
nand U10355 (N_10355,N_7977,N_8760);
or U10356 (N_10356,N_7644,N_7571);
and U10357 (N_10357,N_8605,N_7619);
xnor U10358 (N_10358,N_7901,N_8881);
and U10359 (N_10359,N_8433,N_8729);
and U10360 (N_10360,N_7700,N_7576);
nand U10361 (N_10361,N_8276,N_8416);
and U10362 (N_10362,N_8026,N_8264);
nor U10363 (N_10363,N_7674,N_8883);
xnor U10364 (N_10364,N_8743,N_8127);
nand U10365 (N_10365,N_8519,N_7556);
nand U10366 (N_10366,N_7749,N_8225);
nor U10367 (N_10367,N_8243,N_8861);
or U10368 (N_10368,N_8360,N_8481);
and U10369 (N_10369,N_8133,N_8662);
and U10370 (N_10370,N_8419,N_8209);
or U10371 (N_10371,N_8794,N_8531);
nor U10372 (N_10372,N_8024,N_8011);
or U10373 (N_10373,N_7528,N_8446);
nor U10374 (N_10374,N_8563,N_8002);
nor U10375 (N_10375,N_7667,N_8831);
or U10376 (N_10376,N_8422,N_8719);
nor U10377 (N_10377,N_8168,N_7543);
nand U10378 (N_10378,N_8723,N_8143);
nand U10379 (N_10379,N_8953,N_8039);
xor U10380 (N_10380,N_7803,N_7649);
nand U10381 (N_10381,N_8903,N_7532);
and U10382 (N_10382,N_8742,N_7659);
nand U10383 (N_10383,N_8548,N_8518);
nand U10384 (N_10384,N_8570,N_8634);
and U10385 (N_10385,N_8234,N_8540);
xnor U10386 (N_10386,N_8485,N_7742);
or U10387 (N_10387,N_8351,N_8847);
and U10388 (N_10388,N_8565,N_8945);
nand U10389 (N_10389,N_8812,N_8757);
and U10390 (N_10390,N_8387,N_8497);
and U10391 (N_10391,N_7666,N_8701);
nor U10392 (N_10392,N_8538,N_8173);
nor U10393 (N_10393,N_8674,N_7601);
xor U10394 (N_10394,N_7856,N_8865);
nand U10395 (N_10395,N_7537,N_7764);
nor U10396 (N_10396,N_8157,N_7633);
nand U10397 (N_10397,N_8792,N_8370);
or U10398 (N_10398,N_8325,N_8671);
nand U10399 (N_10399,N_7669,N_8537);
nand U10400 (N_10400,N_8624,N_7815);
or U10401 (N_10401,N_8316,N_8116);
and U10402 (N_10402,N_8126,N_7674);
or U10403 (N_10403,N_7947,N_7714);
nand U10404 (N_10404,N_7781,N_8583);
or U10405 (N_10405,N_8481,N_7859);
or U10406 (N_10406,N_8446,N_8039);
nand U10407 (N_10407,N_8297,N_8069);
nor U10408 (N_10408,N_7758,N_8670);
and U10409 (N_10409,N_8339,N_7525);
or U10410 (N_10410,N_8838,N_7975);
nand U10411 (N_10411,N_7882,N_7837);
or U10412 (N_10412,N_8679,N_8187);
and U10413 (N_10413,N_8264,N_8204);
nor U10414 (N_10414,N_8703,N_7963);
nor U10415 (N_10415,N_8253,N_8261);
nand U10416 (N_10416,N_8177,N_7629);
or U10417 (N_10417,N_8527,N_8497);
nand U10418 (N_10418,N_8725,N_7608);
nand U10419 (N_10419,N_8382,N_7763);
or U10420 (N_10420,N_8065,N_8907);
or U10421 (N_10421,N_8029,N_8454);
nand U10422 (N_10422,N_8763,N_7645);
xor U10423 (N_10423,N_8996,N_7724);
or U10424 (N_10424,N_7902,N_8046);
or U10425 (N_10425,N_8272,N_8171);
or U10426 (N_10426,N_8962,N_8558);
nor U10427 (N_10427,N_7975,N_8226);
xor U10428 (N_10428,N_8936,N_8142);
and U10429 (N_10429,N_8814,N_8993);
or U10430 (N_10430,N_8246,N_8886);
or U10431 (N_10431,N_8973,N_7777);
and U10432 (N_10432,N_8163,N_8892);
and U10433 (N_10433,N_8668,N_8401);
and U10434 (N_10434,N_8219,N_7675);
or U10435 (N_10435,N_8995,N_8153);
nor U10436 (N_10436,N_8156,N_7693);
or U10437 (N_10437,N_8142,N_8459);
xor U10438 (N_10438,N_8048,N_8615);
and U10439 (N_10439,N_8568,N_7793);
or U10440 (N_10440,N_8609,N_7698);
xnor U10441 (N_10441,N_8496,N_8004);
nor U10442 (N_10442,N_7940,N_8171);
nor U10443 (N_10443,N_8466,N_8707);
nand U10444 (N_10444,N_7539,N_8034);
and U10445 (N_10445,N_8808,N_8630);
or U10446 (N_10446,N_8907,N_7569);
and U10447 (N_10447,N_7860,N_8586);
and U10448 (N_10448,N_7769,N_7931);
nor U10449 (N_10449,N_8632,N_7936);
or U10450 (N_10450,N_7774,N_8836);
xnor U10451 (N_10451,N_8436,N_7500);
nand U10452 (N_10452,N_8630,N_8258);
or U10453 (N_10453,N_7993,N_8879);
or U10454 (N_10454,N_8935,N_7690);
xor U10455 (N_10455,N_8865,N_8546);
xnor U10456 (N_10456,N_7546,N_8667);
nand U10457 (N_10457,N_8411,N_8804);
and U10458 (N_10458,N_8938,N_7987);
nand U10459 (N_10459,N_8932,N_8140);
nand U10460 (N_10460,N_7686,N_8863);
nand U10461 (N_10461,N_7555,N_8116);
nor U10462 (N_10462,N_8438,N_7666);
nor U10463 (N_10463,N_8940,N_7678);
and U10464 (N_10464,N_8837,N_8625);
and U10465 (N_10465,N_8284,N_7603);
or U10466 (N_10466,N_7898,N_7955);
nand U10467 (N_10467,N_7864,N_8656);
or U10468 (N_10468,N_7617,N_7739);
and U10469 (N_10469,N_7571,N_8634);
and U10470 (N_10470,N_8176,N_8510);
or U10471 (N_10471,N_8914,N_8713);
nand U10472 (N_10472,N_8698,N_8641);
and U10473 (N_10473,N_8697,N_8875);
nand U10474 (N_10474,N_8464,N_8759);
xor U10475 (N_10475,N_7787,N_8282);
or U10476 (N_10476,N_8743,N_8732);
xor U10477 (N_10477,N_7934,N_8674);
or U10478 (N_10478,N_8478,N_7578);
nand U10479 (N_10479,N_8779,N_8110);
nand U10480 (N_10480,N_8916,N_7648);
nor U10481 (N_10481,N_7751,N_8393);
nand U10482 (N_10482,N_7824,N_7880);
or U10483 (N_10483,N_7923,N_8094);
nor U10484 (N_10484,N_8683,N_7586);
nand U10485 (N_10485,N_8034,N_8518);
nand U10486 (N_10486,N_8074,N_8638);
and U10487 (N_10487,N_7942,N_8311);
nand U10488 (N_10488,N_7596,N_7951);
nor U10489 (N_10489,N_8475,N_8303);
or U10490 (N_10490,N_7745,N_8896);
or U10491 (N_10491,N_8619,N_7678);
nor U10492 (N_10492,N_8667,N_7837);
nand U10493 (N_10493,N_8274,N_8820);
xor U10494 (N_10494,N_7657,N_8262);
and U10495 (N_10495,N_7766,N_8459);
nor U10496 (N_10496,N_8503,N_8881);
nand U10497 (N_10497,N_7694,N_7840);
or U10498 (N_10498,N_8973,N_8236);
xor U10499 (N_10499,N_7601,N_7540);
nand U10500 (N_10500,N_9761,N_9608);
and U10501 (N_10501,N_10348,N_10491);
or U10502 (N_10502,N_9749,N_9946);
and U10503 (N_10503,N_9852,N_10175);
and U10504 (N_10504,N_9320,N_9037);
xnor U10505 (N_10505,N_10404,N_9527);
and U10506 (N_10506,N_9895,N_9600);
nor U10507 (N_10507,N_9162,N_9211);
and U10508 (N_10508,N_10007,N_9491);
xnor U10509 (N_10509,N_9110,N_9854);
or U10510 (N_10510,N_9356,N_9941);
nand U10511 (N_10511,N_9016,N_10420);
nand U10512 (N_10512,N_10119,N_10020);
and U10513 (N_10513,N_10457,N_9744);
nand U10514 (N_10514,N_9509,N_9953);
or U10515 (N_10515,N_9061,N_9611);
and U10516 (N_10516,N_9569,N_9406);
or U10517 (N_10517,N_10084,N_9970);
and U10518 (N_10518,N_10039,N_9118);
nand U10519 (N_10519,N_10398,N_9397);
and U10520 (N_10520,N_10330,N_10471);
nand U10521 (N_10521,N_9214,N_9695);
or U10522 (N_10522,N_10373,N_9480);
nand U10523 (N_10523,N_9699,N_9124);
or U10524 (N_10524,N_10217,N_9777);
nand U10525 (N_10525,N_9404,N_10280);
nand U10526 (N_10526,N_9660,N_9903);
nand U10527 (N_10527,N_9217,N_9187);
and U10528 (N_10528,N_9936,N_9785);
nor U10529 (N_10529,N_10079,N_9753);
nand U10530 (N_10530,N_10319,N_9666);
and U10531 (N_10531,N_9328,N_9713);
or U10532 (N_10532,N_9866,N_10257);
and U10533 (N_10533,N_10019,N_9440);
and U10534 (N_10534,N_10252,N_10120);
and U10535 (N_10535,N_9261,N_9776);
nor U10536 (N_10536,N_10183,N_9708);
xor U10537 (N_10537,N_9568,N_9161);
and U10538 (N_10538,N_10388,N_10052);
nand U10539 (N_10539,N_9846,N_10136);
and U10540 (N_10540,N_9621,N_9478);
or U10541 (N_10541,N_10075,N_10249);
and U10542 (N_10542,N_9437,N_10444);
nand U10543 (N_10543,N_9519,N_10387);
nand U10544 (N_10544,N_9090,N_9296);
nor U10545 (N_10545,N_9703,N_10029);
xnor U10546 (N_10546,N_9825,N_9726);
nor U10547 (N_10547,N_9318,N_10392);
or U10548 (N_10548,N_9487,N_10071);
nor U10549 (N_10549,N_9150,N_9091);
nor U10550 (N_10550,N_9691,N_9538);
nor U10551 (N_10551,N_9439,N_9121);
or U10552 (N_10552,N_10361,N_9531);
nand U10553 (N_10553,N_9779,N_9160);
nand U10554 (N_10554,N_10100,N_9553);
and U10555 (N_10555,N_9496,N_10043);
or U10556 (N_10556,N_9040,N_10307);
nand U10557 (N_10557,N_10167,N_9559);
nand U10558 (N_10558,N_9125,N_10146);
nand U10559 (N_10559,N_9712,N_9722);
and U10560 (N_10560,N_10322,N_9354);
nand U10561 (N_10561,N_9917,N_10439);
nor U10562 (N_10562,N_10226,N_10211);
or U10563 (N_10563,N_9624,N_10297);
or U10564 (N_10564,N_9286,N_9752);
and U10565 (N_10565,N_9780,N_9270);
nor U10566 (N_10566,N_9826,N_10378);
nor U10567 (N_10567,N_10011,N_10156);
or U10568 (N_10568,N_9649,N_10062);
and U10569 (N_10569,N_10158,N_10204);
and U10570 (N_10570,N_9801,N_9949);
nand U10571 (N_10571,N_9813,N_10376);
or U10572 (N_10572,N_9443,N_9802);
and U10573 (N_10573,N_9488,N_9358);
nor U10574 (N_10574,N_10213,N_9832);
nor U10575 (N_10575,N_9881,N_9363);
and U10576 (N_10576,N_10060,N_10061);
xnor U10577 (N_10577,N_9355,N_10144);
nand U10578 (N_10578,N_9892,N_9224);
nor U10579 (N_10579,N_10405,N_9789);
nor U10580 (N_10580,N_10097,N_9717);
and U10581 (N_10581,N_10448,N_9468);
xnor U10582 (N_10582,N_9079,N_9021);
nor U10583 (N_10583,N_10428,N_10401);
nor U10584 (N_10584,N_10181,N_10415);
nor U10585 (N_10585,N_9141,N_9741);
xor U10586 (N_10586,N_9380,N_9838);
or U10587 (N_10587,N_9032,N_10272);
xor U10588 (N_10588,N_9095,N_9921);
or U10589 (N_10589,N_9038,N_10261);
or U10590 (N_10590,N_9909,N_10406);
nand U10591 (N_10591,N_9830,N_9853);
nor U10592 (N_10592,N_9815,N_9479);
and U10593 (N_10593,N_9366,N_9714);
nor U10594 (N_10594,N_9275,N_10067);
or U10595 (N_10595,N_9481,N_9243);
nand U10596 (N_10596,N_9837,N_9414);
xor U10597 (N_10597,N_9996,N_9191);
nand U10598 (N_10598,N_9989,N_9075);
nand U10599 (N_10599,N_9044,N_9295);
nor U10600 (N_10600,N_10228,N_10018);
or U10601 (N_10601,N_9030,N_9539);
nand U10602 (N_10602,N_9516,N_9111);
or U10603 (N_10603,N_10174,N_10196);
nand U10604 (N_10604,N_9847,N_10314);
or U10605 (N_10605,N_9576,N_10054);
nand U10606 (N_10606,N_9051,N_9492);
nor U10607 (N_10607,N_9848,N_9638);
or U10608 (N_10608,N_9513,N_9563);
nand U10609 (N_10609,N_9522,N_9011);
and U10610 (N_10610,N_10273,N_9652);
nor U10611 (N_10611,N_9850,N_9346);
nor U10612 (N_10612,N_9601,N_9065);
xor U10613 (N_10613,N_10059,N_9822);
nand U10614 (N_10614,N_9583,N_10370);
xor U10615 (N_10615,N_10169,N_10161);
nor U10616 (N_10616,N_9705,N_9985);
and U10617 (N_10617,N_9631,N_9504);
nor U10618 (N_10618,N_9880,N_10472);
xor U10619 (N_10619,N_9581,N_10038);
nor U10620 (N_10620,N_9334,N_9849);
and U10621 (N_10621,N_9294,N_10206);
and U10622 (N_10622,N_9535,N_9341);
or U10623 (N_10623,N_9743,N_9507);
nor U10624 (N_10624,N_9928,N_9043);
nor U10625 (N_10625,N_9639,N_9344);
nor U10626 (N_10626,N_9461,N_10292);
and U10627 (N_10627,N_10334,N_9132);
nor U10628 (N_10628,N_9940,N_10031);
or U10629 (N_10629,N_10456,N_10078);
and U10630 (N_10630,N_9787,N_10131);
nand U10631 (N_10631,N_10188,N_9466);
nor U10632 (N_10632,N_10197,N_10362);
and U10633 (N_10633,N_10001,N_10024);
or U10634 (N_10634,N_9050,N_9693);
or U10635 (N_10635,N_9092,N_9742);
and U10636 (N_10636,N_9871,N_9590);
nand U10637 (N_10637,N_10032,N_9457);
nand U10638 (N_10638,N_9681,N_10123);
nor U10639 (N_10639,N_10186,N_10336);
or U10640 (N_10640,N_9603,N_10419);
or U10641 (N_10641,N_9382,N_9931);
nor U10642 (N_10642,N_9186,N_10000);
nor U10643 (N_10643,N_9001,N_9840);
and U10644 (N_10644,N_9416,N_9786);
nor U10645 (N_10645,N_9302,N_9063);
and U10646 (N_10646,N_10058,N_9374);
or U10647 (N_10647,N_9879,N_10089);
nor U10648 (N_10648,N_10423,N_10281);
xnor U10649 (N_10649,N_10070,N_10263);
or U10650 (N_10650,N_9335,N_10497);
and U10651 (N_10651,N_9300,N_10094);
and U10652 (N_10652,N_9325,N_9987);
nand U10653 (N_10653,N_10092,N_9348);
or U10654 (N_10654,N_9431,N_9922);
or U10655 (N_10655,N_9672,N_10085);
nor U10656 (N_10656,N_10172,N_9756);
xor U10657 (N_10657,N_9399,N_9113);
nor U10658 (N_10658,N_10008,N_9035);
nand U10659 (N_10659,N_9657,N_9448);
or U10660 (N_10660,N_10363,N_9209);
or U10661 (N_10661,N_9793,N_9782);
and U10662 (N_10662,N_9100,N_9526);
and U10663 (N_10663,N_9905,N_10027);
nor U10664 (N_10664,N_9271,N_9916);
nor U10665 (N_10665,N_9446,N_10076);
and U10666 (N_10666,N_9973,N_9867);
xor U10667 (N_10667,N_10074,N_9556);
nand U10668 (N_10668,N_9316,N_9907);
nor U10669 (N_10669,N_9870,N_9278);
nor U10670 (N_10670,N_9924,N_9421);
or U10671 (N_10671,N_9758,N_10244);
xnor U10672 (N_10672,N_10461,N_9904);
or U10673 (N_10673,N_9661,N_9855);
or U10674 (N_10674,N_9763,N_9284);
nand U10675 (N_10675,N_10256,N_9472);
and U10676 (N_10676,N_9925,N_9873);
and U10677 (N_10677,N_10137,N_9643);
nand U10678 (N_10678,N_9455,N_10486);
nand U10679 (N_10679,N_9747,N_9000);
or U10680 (N_10680,N_10125,N_9984);
and U10681 (N_10681,N_9817,N_10360);
xor U10682 (N_10682,N_9543,N_10332);
and U10683 (N_10683,N_9735,N_9860);
nand U10684 (N_10684,N_10436,N_9013);
and U10685 (N_10685,N_10237,N_9349);
or U10686 (N_10686,N_9142,N_10275);
or U10687 (N_10687,N_9963,N_9518);
or U10688 (N_10688,N_9449,N_10176);
nor U10689 (N_10689,N_10016,N_10493);
or U10690 (N_10690,N_10099,N_9140);
nor U10691 (N_10691,N_10238,N_9236);
nand U10692 (N_10692,N_9506,N_9645);
or U10693 (N_10693,N_9410,N_10301);
or U10694 (N_10694,N_9131,N_9595);
or U10695 (N_10695,N_10350,N_9309);
or U10696 (N_10696,N_9857,N_10165);
nor U10697 (N_10697,N_9444,N_9107);
and U10698 (N_10698,N_9195,N_10434);
or U10699 (N_10699,N_9408,N_10110);
or U10700 (N_10700,N_10202,N_9222);
nand U10701 (N_10701,N_10342,N_9223);
or U10702 (N_10702,N_10313,N_10382);
nand U10703 (N_10703,N_9676,N_10320);
or U10704 (N_10704,N_9024,N_10247);
and U10705 (N_10705,N_10379,N_9586);
nand U10706 (N_10706,N_10296,N_9541);
nand U10707 (N_10707,N_10106,N_10021);
or U10708 (N_10708,N_10259,N_10412);
and U10709 (N_10709,N_10484,N_9002);
xnor U10710 (N_10710,N_10278,N_10364);
nand U10711 (N_10711,N_9684,N_9423);
nand U10712 (N_10712,N_9663,N_9280);
and U10713 (N_10713,N_10338,N_10240);
and U10714 (N_10714,N_10317,N_9177);
and U10715 (N_10715,N_10080,N_9775);
or U10716 (N_10716,N_9700,N_10427);
or U10717 (N_10717,N_9613,N_9551);
or U10718 (N_10718,N_10105,N_9352);
xor U10719 (N_10719,N_10316,N_10145);
nand U10720 (N_10720,N_10205,N_10270);
and U10721 (N_10721,N_9598,N_9105);
and U10722 (N_10722,N_10453,N_9723);
xor U10723 (N_10723,N_10195,N_10390);
and U10724 (N_10724,N_9605,N_9218);
xor U10725 (N_10725,N_10480,N_10132);
nor U10726 (N_10726,N_10128,N_10250);
or U10727 (N_10727,N_10182,N_10114);
and U10728 (N_10728,N_9912,N_10288);
or U10729 (N_10729,N_9256,N_9788);
and U10730 (N_10730,N_9567,N_10231);
and U10731 (N_10731,N_10393,N_10285);
and U10732 (N_10732,N_10417,N_9650);
nand U10733 (N_10733,N_9642,N_10009);
and U10734 (N_10734,N_9829,N_9773);
and U10735 (N_10735,N_10303,N_9463);
nand U10736 (N_10736,N_9233,N_9493);
or U10737 (N_10737,N_9266,N_10284);
and U10738 (N_10738,N_9134,N_9086);
or U10739 (N_10739,N_10383,N_9894);
or U10740 (N_10740,N_10180,N_9505);
nand U10741 (N_10741,N_9047,N_9755);
and U10742 (N_10742,N_9384,N_9008);
xor U10743 (N_10743,N_10343,N_9625);
and U10744 (N_10744,N_9136,N_9738);
and U10745 (N_10745,N_9721,N_10050);
nand U10746 (N_10746,N_9732,N_10395);
and U10747 (N_10747,N_10358,N_10331);
nand U10748 (N_10748,N_9915,N_9791);
nand U10749 (N_10749,N_9696,N_9248);
or U10750 (N_10750,N_10044,N_10005);
or U10751 (N_10751,N_9620,N_10037);
or U10752 (N_10752,N_9938,N_9333);
and U10753 (N_10753,N_9199,N_9863);
or U10754 (N_10754,N_9685,N_10198);
and U10755 (N_10755,N_9843,N_9943);
or U10756 (N_10756,N_9015,N_9972);
or U10757 (N_10757,N_10143,N_9053);
nand U10758 (N_10758,N_9552,N_9350);
nand U10759 (N_10759,N_10066,N_10242);
nor U10760 (N_10760,N_10308,N_9206);
nor U10761 (N_10761,N_9144,N_9204);
and U10762 (N_10762,N_10015,N_9804);
nand U10763 (N_10763,N_9971,N_9094);
nand U10764 (N_10764,N_9719,N_9580);
and U10765 (N_10765,N_9687,N_9281);
xnor U10766 (N_10766,N_10366,N_9778);
or U10767 (N_10767,N_9899,N_9658);
xor U10768 (N_10768,N_10177,N_10006);
and U10769 (N_10769,N_9405,N_9314);
nor U10770 (N_10770,N_9495,N_10246);
xor U10771 (N_10771,N_10433,N_9428);
and U10772 (N_10772,N_9010,N_9438);
nand U10773 (N_10773,N_9361,N_10315);
xnor U10774 (N_10774,N_9088,N_9819);
nor U10775 (N_10775,N_9103,N_10209);
and U10776 (N_10776,N_9896,N_9022);
nand U10777 (N_10777,N_10460,N_9220);
and U10778 (N_10778,N_9549,N_10470);
nand U10779 (N_10779,N_9555,N_10260);
and U10780 (N_10780,N_9227,N_10450);
nand U10781 (N_10781,N_9716,N_9373);
or U10782 (N_10782,N_9082,N_9636);
or U10783 (N_10783,N_9564,N_10243);
nand U10784 (N_10784,N_9071,N_9876);
nand U10785 (N_10785,N_9189,N_9181);
nand U10786 (N_10786,N_10036,N_10269);
nor U10787 (N_10787,N_9036,N_10391);
or U10788 (N_10788,N_9720,N_10056);
nor U10789 (N_10789,N_10113,N_9565);
nand U10790 (N_10790,N_10115,N_9059);
or U10791 (N_10791,N_9212,N_10191);
or U10792 (N_10792,N_10289,N_9288);
or U10793 (N_10793,N_10164,N_10463);
nand U10794 (N_10794,N_9596,N_9751);
or U10795 (N_10795,N_10200,N_9554);
and U10796 (N_10796,N_9106,N_9797);
nand U10797 (N_10797,N_9612,N_9273);
xnor U10798 (N_10798,N_9766,N_9532);
and U10799 (N_10799,N_9485,N_9258);
nand U10800 (N_10800,N_9375,N_9178);
nand U10801 (N_10801,N_10236,N_10063);
nand U10802 (N_10802,N_9740,N_9087);
nand U10803 (N_10803,N_9683,N_9321);
nor U10804 (N_10804,N_10277,N_9025);
nor U10805 (N_10805,N_9795,N_10013);
nor U10806 (N_10806,N_9644,N_9913);
nor U10807 (N_10807,N_9471,N_9180);
or U10808 (N_10808,N_10357,N_9339);
nor U10809 (N_10809,N_9974,N_9677);
and U10810 (N_10810,N_9659,N_9622);
nor U10811 (N_10811,N_10218,N_9298);
nand U10812 (N_10812,N_9229,N_9164);
nor U10813 (N_10813,N_9007,N_9640);
nand U10814 (N_10814,N_10251,N_10048);
or U10815 (N_10815,N_9986,N_9772);
nor U10816 (N_10816,N_9415,N_9247);
and U10817 (N_10817,N_10046,N_10150);
nor U10818 (N_10818,N_10306,N_10481);
nor U10819 (N_10819,N_9458,N_9566);
nand U10820 (N_10820,N_10160,N_10349);
nor U10821 (N_10821,N_9514,N_10081);
nor U10822 (N_10822,N_9833,N_9948);
nand U10823 (N_10823,N_9332,N_9179);
nand U10824 (N_10824,N_9097,N_9285);
and U10825 (N_10825,N_10418,N_9221);
nand U10826 (N_10826,N_9289,N_9297);
and U10827 (N_10827,N_9155,N_10411);
nand U10828 (N_10828,N_10445,N_10371);
nor U10829 (N_10829,N_9133,N_10309);
or U10830 (N_10830,N_9099,N_9653);
nor U10831 (N_10831,N_9319,N_9052);
nand U10832 (N_10832,N_9089,N_9530);
nor U10833 (N_10833,N_9197,N_10335);
or U10834 (N_10834,N_9654,N_9196);
nand U10835 (N_10835,N_10402,N_9809);
nor U10836 (N_10836,N_9508,N_9918);
and U10837 (N_10837,N_9964,N_9433);
and U10838 (N_10838,N_10225,N_9469);
nor U10839 (N_10839,N_9387,N_9456);
and U10840 (N_10840,N_10283,N_9126);
or U10841 (N_10841,N_9338,N_9898);
nand U10842 (N_10842,N_10034,N_10149);
or U10843 (N_10843,N_9307,N_9368);
or U10844 (N_10844,N_9462,N_10438);
or U10845 (N_10845,N_10414,N_9060);
nand U10846 (N_10846,N_9878,N_9253);
xor U10847 (N_10847,N_10093,N_9154);
and U10848 (N_10848,N_10359,N_9420);
nor U10849 (N_10849,N_9120,N_9942);
xnor U10850 (N_10850,N_9459,N_10384);
nand U10851 (N_10851,N_9135,N_10170);
xor U10852 (N_10852,N_9093,N_9231);
or U10853 (N_10853,N_9757,N_10431);
nand U10854 (N_10854,N_9842,N_9874);
and U10855 (N_10855,N_10069,N_9900);
nand U10856 (N_10856,N_9617,N_9616);
xor U10857 (N_10857,N_10082,N_9351);
and U10858 (N_10858,N_9869,N_9524);
nand U10859 (N_10859,N_10192,N_9077);
or U10860 (N_10860,N_9619,N_10318);
nor U10861 (N_10861,N_9427,N_9588);
nand U10862 (N_10862,N_9163,N_9413);
and U10863 (N_10863,N_9376,N_10117);
xor U10864 (N_10864,N_10162,N_9175);
nand U10865 (N_10865,N_9004,N_10140);
xor U10866 (N_10866,N_9709,N_9378);
and U10867 (N_10867,N_10104,N_10282);
nor U10868 (N_10868,N_10193,N_9225);
nor U10869 (N_10869,N_10142,N_9911);
or U10870 (N_10870,N_9123,N_10459);
nor U10871 (N_10871,N_9080,N_9340);
nor U10872 (N_10872,N_9465,N_9960);
or U10873 (N_10873,N_9262,N_10091);
nor U10874 (N_10874,N_9230,N_9783);
nor U10875 (N_10875,N_9272,N_10377);
nor U10876 (N_10876,N_10474,N_10290);
nor U10877 (N_10877,N_9845,N_10399);
nor U10878 (N_10878,N_9991,N_10157);
and U10879 (N_10879,N_9246,N_9337);
or U10880 (N_10880,N_9665,N_10155);
nor U10881 (N_10881,N_9547,N_9372);
xnor U10882 (N_10882,N_10443,N_9447);
and U10883 (N_10883,N_10485,N_10327);
or U10884 (N_10884,N_10216,N_9018);
nor U10885 (N_10885,N_10367,N_10138);
nand U10886 (N_10886,N_9994,N_9219);
nor U10887 (N_10887,N_10435,N_9944);
xnor U10888 (N_10888,N_9058,N_9226);
nand U10889 (N_10889,N_9831,N_9730);
and U10890 (N_10890,N_10068,N_10234);
and U10891 (N_10891,N_9770,N_9760);
and U10892 (N_10892,N_9054,N_9419);
and U10893 (N_10893,N_10233,N_9096);
or U10894 (N_10894,N_9651,N_9391);
nor U10895 (N_10895,N_9042,N_10492);
nand U10896 (N_10896,N_10413,N_10171);
or U10897 (N_10897,N_9807,N_9597);
and U10898 (N_10898,N_9582,N_9734);
or U10899 (N_10899,N_9426,N_9293);
or U10900 (N_10900,N_9330,N_9062);
or U10901 (N_10901,N_9303,N_9883);
and U10902 (N_10902,N_9475,N_9499);
xnor U10903 (N_10903,N_10345,N_9737);
and U10904 (N_10904,N_9265,N_10329);
nor U10905 (N_10905,N_9084,N_9183);
nand U10906 (N_10906,N_9704,N_9762);
xnor U10907 (N_10907,N_9794,N_10130);
nor U10908 (N_10908,N_9882,N_10241);
or U10909 (N_10909,N_9235,N_9116);
and U10910 (N_10910,N_9906,N_10397);
nor U10911 (N_10911,N_9923,N_9859);
and U10912 (N_10912,N_9208,N_9627);
xnor U10913 (N_10913,N_10045,N_9525);
and U10914 (N_10914,N_9345,N_9544);
and U10915 (N_10915,N_9571,N_9724);
and U10916 (N_10916,N_9686,N_9520);
xnor U10917 (N_10917,N_10124,N_9901);
or U10918 (N_10918,N_9990,N_9835);
and U10919 (N_10919,N_10083,N_9188);
and U10920 (N_10920,N_10264,N_9517);
or U10921 (N_10921,N_10372,N_9745);
nand U10922 (N_10922,N_9934,N_10253);
or U10923 (N_10923,N_9436,N_9152);
xnor U10924 (N_10924,N_9806,N_10185);
and U10925 (N_10925,N_9228,N_9117);
nand U10926 (N_10926,N_9868,N_9454);
nand U10927 (N_10927,N_10271,N_9170);
nand U10928 (N_10928,N_9585,N_9587);
nand U10929 (N_10929,N_9950,N_9255);
and U10930 (N_10930,N_9697,N_9072);
nand U10931 (N_10931,N_10230,N_9537);
and U10932 (N_10932,N_9353,N_9388);
and U10933 (N_10933,N_9746,N_9497);
nor U10934 (N_10934,N_9926,N_9494);
nand U10935 (N_10935,N_9955,N_9727);
nand U10936 (N_10936,N_10454,N_9329);
nor U10937 (N_10937,N_9083,N_10429);
or U10938 (N_10938,N_9119,N_9573);
and U10939 (N_10939,N_10351,N_9675);
or U10940 (N_10940,N_10148,N_10088);
nor U10941 (N_10941,N_9409,N_10035);
nor U10942 (N_10942,N_9239,N_9528);
nand U10943 (N_10943,N_9865,N_9731);
nor U10944 (N_10944,N_9234,N_9017);
nand U10945 (N_10945,N_9336,N_9184);
or U10946 (N_10946,N_10134,N_9818);
and U10947 (N_10947,N_9242,N_10487);
or U10948 (N_10948,N_10365,N_9192);
and U10949 (N_10949,N_9827,N_9678);
nand U10950 (N_10950,N_9412,N_9877);
or U10951 (N_10951,N_9324,N_10041);
nor U10952 (N_10952,N_9858,N_9889);
nor U10953 (N_10953,N_10215,N_10407);
or U10954 (N_10954,N_10265,N_10255);
xor U10955 (N_10955,N_10014,N_10154);
nor U10956 (N_10956,N_9607,N_9618);
or U10957 (N_10957,N_10087,N_9501);
and U10958 (N_10958,N_10004,N_9205);
xor U10959 (N_10959,N_9167,N_9808);
nand U10960 (N_10960,N_10394,N_9306);
nor U10961 (N_10961,N_10302,N_9129);
nor U10962 (N_10962,N_10294,N_10375);
nand U10963 (N_10963,N_9933,N_9396);
and U10964 (N_10964,N_9389,N_10224);
nor U10965 (N_10965,N_10449,N_10033);
and U10966 (N_10966,N_10003,N_9165);
xor U10967 (N_10967,N_9102,N_9108);
nand U10968 (N_10968,N_9064,N_9930);
and U10969 (N_10969,N_10199,N_10469);
nand U10970 (N_10970,N_9579,N_9407);
or U10971 (N_10971,N_9980,N_9824);
or U10972 (N_10972,N_10299,N_9512);
nand U10973 (N_10973,N_10477,N_10163);
nor U10974 (N_10974,N_9400,N_9157);
or U10975 (N_10975,N_9533,N_9173);
or U10976 (N_10976,N_9799,N_9156);
nand U10977 (N_10977,N_9902,N_10409);
and U10978 (N_10978,N_9626,N_10323);
nor U10979 (N_10979,N_9839,N_10121);
xor U10980 (N_10980,N_9252,N_10212);
or U10981 (N_10981,N_10310,N_10386);
or U10982 (N_10982,N_9591,N_9395);
nor U10983 (N_10983,N_9952,N_10432);
nor U10984 (N_10984,N_9784,N_9422);
nand U10985 (N_10985,N_9689,N_10235);
and U10986 (N_10986,N_10468,N_10055);
or U10987 (N_10987,N_9074,N_9128);
or U10988 (N_10988,N_9821,N_10051);
or U10989 (N_10989,N_10466,N_9812);
nand U10990 (N_10990,N_9811,N_9594);
and U10991 (N_10991,N_9790,N_9593);
or U10992 (N_10992,N_10179,N_9558);
xor U10993 (N_10993,N_10276,N_9771);
and U10994 (N_10994,N_9951,N_9646);
nand U10995 (N_10995,N_10122,N_9545);
nor U10996 (N_10996,N_10352,N_10077);
or U10997 (N_10997,N_9864,N_9814);
or U10998 (N_10998,N_10430,N_9138);
nor U10999 (N_10999,N_10220,N_9728);
and U11000 (N_11000,N_10451,N_9185);
or U11001 (N_11001,N_10426,N_9628);
nor U11002 (N_11002,N_10440,N_9629);
and U11003 (N_11003,N_10495,N_9575);
xor U11004 (N_11004,N_9045,N_10298);
and U11005 (N_11005,N_10109,N_9401);
xnor U11006 (N_11006,N_10221,N_10190);
and U11007 (N_11007,N_9736,N_9067);
nand U11008 (N_11008,N_10325,N_9823);
and U11009 (N_11009,N_10096,N_10047);
or U11010 (N_11010,N_10447,N_9632);
nor U11011 (N_11011,N_9250,N_9988);
or U11012 (N_11012,N_10049,N_9927);
or U11013 (N_11013,N_9633,N_9739);
and U11014 (N_11014,N_9268,N_9198);
and U11015 (N_11015,N_10341,N_9269);
or U11016 (N_11016,N_9039,N_9070);
nor U11017 (N_11017,N_10203,N_9503);
or U11018 (N_11018,N_9139,N_9073);
nor U11019 (N_11019,N_10465,N_9383);
or U11020 (N_11020,N_9207,N_9190);
nor U11021 (N_11021,N_9453,N_10135);
and U11022 (N_11022,N_10118,N_9872);
nor U11023 (N_11023,N_9992,N_9452);
or U11024 (N_11024,N_9648,N_10207);
xnor U11025 (N_11025,N_10369,N_9215);
nor U11026 (N_11026,N_9046,N_9304);
and U11027 (N_11027,N_9393,N_9725);
or U11028 (N_11028,N_9078,N_10328);
nor U11029 (N_11029,N_9369,N_9711);
nor U11030 (N_11030,N_9958,N_10133);
nand U11031 (N_11031,N_10305,N_9800);
nor U11032 (N_11032,N_9523,N_10422);
xor U11033 (N_11033,N_9343,N_9690);
or U11034 (N_11034,N_9394,N_10354);
and U11035 (N_11035,N_9143,N_10266);
nand U11036 (N_11036,N_9315,N_9999);
and U11037 (N_11037,N_10446,N_9995);
and U11038 (N_11038,N_9276,N_10489);
nor U11039 (N_11039,N_10347,N_9604);
or U11040 (N_11040,N_10187,N_9599);
and U11041 (N_11041,N_9418,N_10219);
nor U11042 (N_11042,N_10425,N_10374);
and U11043 (N_11043,N_9210,N_9966);
nand U11044 (N_11044,N_9245,N_9577);
nand U11045 (N_11045,N_10153,N_9759);
nor U11046 (N_11046,N_9257,N_9671);
or U11047 (N_11047,N_9201,N_9213);
nand U11048 (N_11048,N_10488,N_10396);
or U11049 (N_11049,N_9836,N_9560);
nor U11050 (N_11050,N_9982,N_9326);
xnor U11051 (N_11051,N_9975,N_9264);
nand U11052 (N_11052,N_9584,N_10473);
nor U11053 (N_11053,N_9888,N_10479);
or U11054 (N_11054,N_9033,N_9290);
nand U11055 (N_11055,N_10441,N_10147);
and U11056 (N_11056,N_10245,N_9886);
or U11057 (N_11057,N_9115,N_9114);
nor U11058 (N_11058,N_9962,N_9614);
or U11059 (N_11059,N_9908,N_9182);
nor U11060 (N_11060,N_9954,N_10462);
and U11061 (N_11061,N_10017,N_10141);
nor U11062 (N_11062,N_9473,N_9610);
nor U11063 (N_11063,N_9417,N_9359);
nand U11064 (N_11064,N_10239,N_9308);
and U11065 (N_11065,N_9317,N_9137);
nor U11066 (N_11066,N_9578,N_9392);
or U11067 (N_11067,N_9706,N_9750);
or U11068 (N_11068,N_10287,N_9692);
and U11069 (N_11069,N_9055,N_9305);
nor U11070 (N_11070,N_10139,N_9969);
nor U11071 (N_11071,N_9362,N_9820);
nand U11072 (N_11072,N_9887,N_9609);
or U11073 (N_11073,N_10267,N_9049);
xnor U11074 (N_11074,N_9623,N_10353);
nor U11075 (N_11075,N_9085,N_9068);
and U11076 (N_11076,N_9965,N_9130);
nor U11077 (N_11077,N_9174,N_10442);
nand U11078 (N_11078,N_9536,N_10380);
and U11079 (N_11079,N_10090,N_9012);
nor U11080 (N_11080,N_9589,N_9028);
nand U11081 (N_11081,N_9680,N_9311);
nor U11082 (N_11082,N_9637,N_10102);
nor U11083 (N_11083,N_9435,N_9803);
xor U11084 (N_11084,N_9470,N_10065);
nand U11085 (N_11085,N_9816,N_10333);
or U11086 (N_11086,N_9005,N_9707);
or U11087 (N_11087,N_9939,N_10458);
or U11088 (N_11088,N_9920,N_9656);
and U11089 (N_11089,N_9147,N_9403);
nor U11090 (N_11090,N_9014,N_9765);
or U11091 (N_11091,N_9364,N_9548);
or U11092 (N_11092,N_9026,N_10346);
or U11093 (N_11093,N_10010,N_9425);
and U11094 (N_11094,N_10408,N_9483);
and U11095 (N_11095,N_9546,N_10356);
and U11096 (N_11096,N_10496,N_10340);
nand U11097 (N_11097,N_9474,N_9327);
xor U11098 (N_11098,N_9718,N_10339);
or U11099 (N_11099,N_9961,N_9331);
nor U11100 (N_11100,N_9856,N_9460);
nor U11101 (N_11101,N_9006,N_9274);
or U11102 (N_11102,N_9057,N_9216);
nand U11103 (N_11103,N_9562,N_9445);
nand U11104 (N_11104,N_9733,N_10494);
or U11105 (N_11105,N_9267,N_9893);
xnor U11106 (N_11106,N_9476,N_10116);
nor U11107 (N_11107,N_9635,N_9615);
or U11108 (N_11108,N_9056,N_9968);
or U11109 (N_11109,N_10416,N_9260);
and U11110 (N_11110,N_9381,N_9630);
and U11111 (N_11111,N_10300,N_9467);
or U11112 (N_11112,N_9442,N_9029);
or U11113 (N_11113,N_9312,N_10424);
nand U11114 (N_11114,N_9489,N_10028);
nand U11115 (N_11115,N_9670,N_9561);
or U11116 (N_11116,N_9529,N_9710);
and U11117 (N_11117,N_9841,N_10227);
or U11118 (N_11118,N_10108,N_9292);
nor U11119 (N_11119,N_9498,N_10184);
or U11120 (N_11120,N_10232,N_9673);
nor U11121 (N_11121,N_10107,N_9510);
or U11122 (N_11122,N_9398,N_10293);
and U11123 (N_11123,N_9781,N_9935);
nand U11124 (N_11124,N_9020,N_10490);
xnor U11125 (N_11125,N_9193,N_10166);
xnor U11126 (N_11126,N_10022,N_9978);
and U11127 (N_11127,N_9048,N_9109);
nand U11128 (N_11128,N_9009,N_9377);
and U11129 (N_11129,N_9919,N_9667);
nand U11130 (N_11130,N_10201,N_9715);
or U11131 (N_11131,N_9249,N_9282);
xor U11132 (N_11132,N_9360,N_9166);
and U11133 (N_11133,N_9194,N_9441);
nand U11134 (N_11134,N_9238,N_10152);
and U11135 (N_11135,N_10295,N_9983);
nand U11136 (N_11136,N_9884,N_9957);
nor U11137 (N_11137,N_9729,N_10229);
nand U11138 (N_11138,N_9347,N_10168);
nor U11139 (N_11139,N_9310,N_9844);
nand U11140 (N_11140,N_9402,N_9550);
nor U11141 (N_11141,N_9301,N_9159);
and U11142 (N_11142,N_9322,N_10389);
nand U11143 (N_11143,N_9244,N_9112);
xor U11144 (N_11144,N_9200,N_10072);
and U11145 (N_11145,N_9313,N_9081);
nor U11146 (N_11146,N_10223,N_10455);
and U11147 (N_11147,N_9386,N_10101);
nand U11148 (N_11148,N_9176,N_10403);
nor U11149 (N_11149,N_9521,N_10286);
or U11150 (N_11150,N_9237,N_9370);
nor U11151 (N_11151,N_9768,N_10026);
and U11152 (N_11152,N_9602,N_9390);
nand U11153 (N_11153,N_9076,N_9158);
nand U11154 (N_11154,N_9259,N_10112);
nor U11155 (N_11155,N_10042,N_10291);
nand U11156 (N_11156,N_9041,N_10312);
or U11157 (N_11157,N_9450,N_9592);
nand U11158 (N_11158,N_9798,N_9828);
and U11159 (N_11159,N_9655,N_10064);
and U11160 (N_11160,N_9490,N_10086);
nand U11161 (N_11161,N_9947,N_9146);
nand U11162 (N_11162,N_9098,N_9851);
or U11163 (N_11163,N_10279,N_9764);
and U11164 (N_11164,N_9367,N_9241);
nor U11165 (N_11165,N_9694,N_9153);
nand U11166 (N_11166,N_9557,N_9202);
and U11167 (N_11167,N_9769,N_9500);
nand U11168 (N_11168,N_9003,N_9662);
xor U11169 (N_11169,N_10030,N_10321);
xor U11170 (N_11170,N_10381,N_10053);
nor U11171 (N_11171,N_9792,N_9365);
or U11172 (N_11172,N_10189,N_10210);
nand U11173 (N_11173,N_9342,N_9932);
and U11174 (N_11174,N_10498,N_9664);
nand U11175 (N_11175,N_9890,N_9861);
nor U11176 (N_11176,N_9956,N_10476);
or U11177 (N_11177,N_9810,N_10208);
nor U11178 (N_11178,N_10151,N_10129);
xnor U11179 (N_11179,N_9976,N_10012);
or U11180 (N_11180,N_10400,N_10002);
nand U11181 (N_11181,N_10311,N_9981);
and U11182 (N_11182,N_10126,N_9283);
nand U11183 (N_11183,N_9634,N_9682);
or U11184 (N_11184,N_9891,N_10268);
xor U11185 (N_11185,N_10344,N_9674);
and U11186 (N_11186,N_10385,N_9959);
nand U11187 (N_11187,N_10159,N_9979);
and U11188 (N_11188,N_9534,N_9279);
or U11189 (N_11189,N_9151,N_10103);
or U11190 (N_11190,N_10464,N_9240);
nor U11191 (N_11191,N_9701,N_10040);
nor U11192 (N_11192,N_9254,N_9862);
or U11193 (N_11193,N_9477,N_9031);
nand U11194 (N_11194,N_9251,N_9834);
or U11195 (N_11195,N_9127,N_9104);
or U11196 (N_11196,N_9027,N_9669);
nor U11197 (N_11197,N_9515,N_9432);
and U11198 (N_11198,N_10178,N_10304);
or U11199 (N_11199,N_10073,N_9748);
and U11200 (N_11200,N_10025,N_10452);
nand U11201 (N_11201,N_10194,N_9574);
nand U11202 (N_11202,N_9998,N_9287);
nor U11203 (N_11203,N_10095,N_9647);
nand U11204 (N_11204,N_9019,N_10337);
and U11205 (N_11205,N_10499,N_10368);
nor U11206 (N_11206,N_9929,N_9034);
and U11207 (N_11207,N_9482,N_9688);
or U11208 (N_11208,N_10478,N_9371);
or U11209 (N_11209,N_10324,N_9145);
xor U11210 (N_11210,N_9540,N_10111);
and U11211 (N_11211,N_9875,N_9023);
and U11212 (N_11212,N_9291,N_9937);
and U11213 (N_11213,N_9679,N_9502);
nand U11214 (N_11214,N_10127,N_10248);
and U11215 (N_11215,N_10173,N_9754);
xnor U11216 (N_11216,N_9486,N_9570);
or U11217 (N_11217,N_9542,N_9357);
and U11218 (N_11218,N_10421,N_9511);
or U11219 (N_11219,N_9945,N_10222);
nand U11220 (N_11220,N_9122,N_9698);
nand U11221 (N_11221,N_9977,N_9277);
or U11222 (N_11222,N_9796,N_9066);
and U11223 (N_11223,N_10475,N_10214);
nor U11224 (N_11224,N_9148,N_9171);
nor U11225 (N_11225,N_9464,N_9910);
nor U11226 (N_11226,N_9168,N_9914);
nor U11227 (N_11227,N_9172,N_9451);
xnor U11228 (N_11228,N_10254,N_9993);
nor U11229 (N_11229,N_9149,N_9702);
xor U11230 (N_11230,N_10274,N_9668);
nand U11231 (N_11231,N_9385,N_10023);
xor U11232 (N_11232,N_9299,N_9169);
or U11233 (N_11233,N_10262,N_9997);
nand U11234 (N_11234,N_9641,N_9967);
nand U11235 (N_11235,N_9411,N_9434);
xor U11236 (N_11236,N_10483,N_10355);
and U11237 (N_11237,N_9484,N_9429);
nand U11238 (N_11238,N_9606,N_9203);
or U11239 (N_11239,N_10467,N_10326);
or U11240 (N_11240,N_9430,N_9805);
and U11241 (N_11241,N_10437,N_9897);
nor U11242 (N_11242,N_9767,N_10410);
and U11243 (N_11243,N_10098,N_9379);
nor U11244 (N_11244,N_9323,N_10258);
nand U11245 (N_11245,N_9885,N_9263);
nand U11246 (N_11246,N_9774,N_9232);
and U11247 (N_11247,N_10057,N_9101);
xor U11248 (N_11248,N_9424,N_9572);
and U11249 (N_11249,N_10482,N_9069);
and U11250 (N_11250,N_9817,N_10455);
nor U11251 (N_11251,N_10063,N_9212);
or U11252 (N_11252,N_9344,N_9481);
nand U11253 (N_11253,N_9084,N_9414);
or U11254 (N_11254,N_10475,N_10199);
nor U11255 (N_11255,N_9022,N_9479);
nand U11256 (N_11256,N_9922,N_10140);
and U11257 (N_11257,N_9372,N_9343);
or U11258 (N_11258,N_9267,N_9951);
nor U11259 (N_11259,N_9104,N_9012);
and U11260 (N_11260,N_10468,N_9177);
nand U11261 (N_11261,N_9118,N_10201);
and U11262 (N_11262,N_10216,N_9347);
nand U11263 (N_11263,N_9751,N_9971);
nand U11264 (N_11264,N_9328,N_9804);
or U11265 (N_11265,N_9360,N_10241);
and U11266 (N_11266,N_9481,N_10257);
nand U11267 (N_11267,N_9706,N_9654);
or U11268 (N_11268,N_9107,N_10087);
xor U11269 (N_11269,N_9269,N_9301);
or U11270 (N_11270,N_9821,N_9564);
and U11271 (N_11271,N_9605,N_10085);
and U11272 (N_11272,N_10321,N_10363);
nand U11273 (N_11273,N_9440,N_10234);
nor U11274 (N_11274,N_9553,N_9596);
nand U11275 (N_11275,N_9485,N_9768);
nor U11276 (N_11276,N_9174,N_9352);
or U11277 (N_11277,N_10009,N_9083);
xor U11278 (N_11278,N_9070,N_9351);
and U11279 (N_11279,N_9637,N_9221);
xnor U11280 (N_11280,N_9632,N_9146);
and U11281 (N_11281,N_9093,N_9322);
nand U11282 (N_11282,N_10462,N_9114);
nor U11283 (N_11283,N_10458,N_10363);
nand U11284 (N_11284,N_9031,N_9874);
nand U11285 (N_11285,N_9965,N_10129);
and U11286 (N_11286,N_9042,N_10184);
nor U11287 (N_11287,N_9088,N_9455);
and U11288 (N_11288,N_9054,N_9220);
and U11289 (N_11289,N_10477,N_10488);
or U11290 (N_11290,N_10127,N_9511);
xor U11291 (N_11291,N_10143,N_9724);
nor U11292 (N_11292,N_9209,N_9736);
and U11293 (N_11293,N_10097,N_9284);
xnor U11294 (N_11294,N_9191,N_10412);
or U11295 (N_11295,N_10124,N_10237);
nor U11296 (N_11296,N_9360,N_9548);
nor U11297 (N_11297,N_9636,N_10026);
and U11298 (N_11298,N_9587,N_10417);
and U11299 (N_11299,N_10123,N_9121);
or U11300 (N_11300,N_9893,N_9753);
nand U11301 (N_11301,N_10488,N_9309);
and U11302 (N_11302,N_10206,N_9373);
xnor U11303 (N_11303,N_9126,N_10423);
nand U11304 (N_11304,N_9681,N_9063);
and U11305 (N_11305,N_9387,N_10266);
nand U11306 (N_11306,N_9897,N_9682);
nand U11307 (N_11307,N_9425,N_9316);
nand U11308 (N_11308,N_9401,N_10146);
xor U11309 (N_11309,N_9413,N_10070);
nor U11310 (N_11310,N_9086,N_9682);
or U11311 (N_11311,N_9478,N_9435);
nand U11312 (N_11312,N_9202,N_10072);
nand U11313 (N_11313,N_9717,N_9242);
xor U11314 (N_11314,N_9845,N_9274);
xnor U11315 (N_11315,N_9288,N_9462);
and U11316 (N_11316,N_9163,N_10427);
nand U11317 (N_11317,N_9831,N_9010);
nand U11318 (N_11318,N_10357,N_9635);
nor U11319 (N_11319,N_10199,N_10091);
nor U11320 (N_11320,N_10272,N_9308);
nor U11321 (N_11321,N_9221,N_9125);
nor U11322 (N_11322,N_10389,N_9299);
or U11323 (N_11323,N_10064,N_9838);
and U11324 (N_11324,N_9122,N_9463);
and U11325 (N_11325,N_9351,N_10335);
nand U11326 (N_11326,N_9801,N_9363);
and U11327 (N_11327,N_10436,N_9720);
and U11328 (N_11328,N_10117,N_9622);
or U11329 (N_11329,N_9709,N_10087);
xnor U11330 (N_11330,N_10215,N_9606);
nor U11331 (N_11331,N_9772,N_9412);
nand U11332 (N_11332,N_9715,N_9854);
and U11333 (N_11333,N_10208,N_9568);
and U11334 (N_11334,N_9851,N_9747);
and U11335 (N_11335,N_9665,N_10002);
nor U11336 (N_11336,N_10138,N_10102);
nand U11337 (N_11337,N_9516,N_10318);
nor U11338 (N_11338,N_10270,N_9977);
nand U11339 (N_11339,N_10189,N_9170);
nor U11340 (N_11340,N_9780,N_9790);
xnor U11341 (N_11341,N_9676,N_9654);
and U11342 (N_11342,N_10023,N_9588);
nor U11343 (N_11343,N_9315,N_9550);
nand U11344 (N_11344,N_10224,N_10490);
and U11345 (N_11345,N_9921,N_9618);
or U11346 (N_11346,N_10077,N_9951);
nor U11347 (N_11347,N_9771,N_9175);
nand U11348 (N_11348,N_9609,N_10328);
nand U11349 (N_11349,N_10031,N_10138);
nor U11350 (N_11350,N_9418,N_10299);
or U11351 (N_11351,N_10290,N_9697);
and U11352 (N_11352,N_9259,N_9658);
nor U11353 (N_11353,N_10109,N_9634);
nand U11354 (N_11354,N_9970,N_9238);
nor U11355 (N_11355,N_9875,N_10149);
nand U11356 (N_11356,N_10257,N_9253);
nand U11357 (N_11357,N_10461,N_10185);
nor U11358 (N_11358,N_10462,N_10139);
xor U11359 (N_11359,N_10122,N_9802);
nor U11360 (N_11360,N_9141,N_10471);
and U11361 (N_11361,N_9252,N_9020);
nand U11362 (N_11362,N_9911,N_10311);
or U11363 (N_11363,N_9261,N_9806);
xor U11364 (N_11364,N_10061,N_10250);
and U11365 (N_11365,N_10460,N_9913);
nor U11366 (N_11366,N_10469,N_9407);
or U11367 (N_11367,N_9560,N_10126);
and U11368 (N_11368,N_9041,N_9328);
nor U11369 (N_11369,N_9843,N_9186);
and U11370 (N_11370,N_10345,N_10330);
and U11371 (N_11371,N_9250,N_10386);
or U11372 (N_11372,N_10043,N_9786);
xnor U11373 (N_11373,N_9457,N_10362);
or U11374 (N_11374,N_9461,N_9253);
and U11375 (N_11375,N_9422,N_10264);
nor U11376 (N_11376,N_9432,N_10272);
or U11377 (N_11377,N_9623,N_9102);
and U11378 (N_11378,N_9099,N_9076);
nor U11379 (N_11379,N_9854,N_9055);
nand U11380 (N_11380,N_9472,N_9697);
nand U11381 (N_11381,N_9665,N_10233);
xor U11382 (N_11382,N_9937,N_9331);
or U11383 (N_11383,N_9794,N_9335);
nor U11384 (N_11384,N_10059,N_10182);
and U11385 (N_11385,N_9180,N_9187);
nand U11386 (N_11386,N_10282,N_10319);
nand U11387 (N_11387,N_9064,N_9626);
and U11388 (N_11388,N_10142,N_10469);
xor U11389 (N_11389,N_9267,N_9085);
nand U11390 (N_11390,N_9479,N_9730);
nand U11391 (N_11391,N_9264,N_10220);
nor U11392 (N_11392,N_9174,N_9124);
xor U11393 (N_11393,N_9264,N_10283);
or U11394 (N_11394,N_9816,N_9933);
nand U11395 (N_11395,N_9015,N_9149);
nor U11396 (N_11396,N_9933,N_9227);
nand U11397 (N_11397,N_9680,N_10310);
or U11398 (N_11398,N_9632,N_9538);
nor U11399 (N_11399,N_10121,N_9789);
xnor U11400 (N_11400,N_9240,N_9585);
nand U11401 (N_11401,N_9843,N_10242);
and U11402 (N_11402,N_9069,N_10224);
xor U11403 (N_11403,N_9564,N_9433);
nor U11404 (N_11404,N_10017,N_9157);
and U11405 (N_11405,N_9612,N_9792);
or U11406 (N_11406,N_10457,N_9754);
nor U11407 (N_11407,N_9257,N_10463);
nor U11408 (N_11408,N_9391,N_9086);
nor U11409 (N_11409,N_9073,N_9751);
xnor U11410 (N_11410,N_10194,N_9546);
and U11411 (N_11411,N_9354,N_10246);
or U11412 (N_11412,N_10182,N_9236);
nor U11413 (N_11413,N_10091,N_9493);
and U11414 (N_11414,N_9732,N_9968);
or U11415 (N_11415,N_10473,N_9661);
nor U11416 (N_11416,N_9534,N_9091);
nand U11417 (N_11417,N_10337,N_10287);
or U11418 (N_11418,N_10024,N_9177);
and U11419 (N_11419,N_9486,N_9078);
nor U11420 (N_11420,N_10317,N_10221);
xor U11421 (N_11421,N_9692,N_9156);
nor U11422 (N_11422,N_9607,N_10308);
nand U11423 (N_11423,N_10199,N_10024);
nand U11424 (N_11424,N_9555,N_10192);
nand U11425 (N_11425,N_9555,N_10092);
and U11426 (N_11426,N_10302,N_9151);
or U11427 (N_11427,N_9309,N_10240);
nor U11428 (N_11428,N_9953,N_9774);
nor U11429 (N_11429,N_10000,N_9336);
nand U11430 (N_11430,N_9759,N_10098);
or U11431 (N_11431,N_9659,N_9820);
and U11432 (N_11432,N_10086,N_10320);
and U11433 (N_11433,N_9934,N_9237);
and U11434 (N_11434,N_9228,N_9525);
nor U11435 (N_11435,N_10375,N_9705);
nor U11436 (N_11436,N_9006,N_10479);
and U11437 (N_11437,N_9923,N_9379);
or U11438 (N_11438,N_9961,N_9802);
and U11439 (N_11439,N_9580,N_9897);
and U11440 (N_11440,N_9041,N_9992);
and U11441 (N_11441,N_9170,N_10339);
and U11442 (N_11442,N_10236,N_10371);
nor U11443 (N_11443,N_9345,N_9225);
nand U11444 (N_11444,N_9304,N_10009);
nor U11445 (N_11445,N_9177,N_10390);
and U11446 (N_11446,N_9624,N_10228);
nor U11447 (N_11447,N_10429,N_9440);
nand U11448 (N_11448,N_9592,N_10092);
nor U11449 (N_11449,N_9225,N_10478);
nor U11450 (N_11450,N_9856,N_9576);
xor U11451 (N_11451,N_9556,N_9557);
or U11452 (N_11452,N_10125,N_9792);
xnor U11453 (N_11453,N_9984,N_10354);
and U11454 (N_11454,N_9116,N_9708);
xnor U11455 (N_11455,N_10448,N_10297);
nand U11456 (N_11456,N_10169,N_10171);
nand U11457 (N_11457,N_10222,N_9020);
nor U11458 (N_11458,N_9917,N_9810);
nand U11459 (N_11459,N_9835,N_10024);
and U11460 (N_11460,N_9304,N_9127);
nand U11461 (N_11461,N_9127,N_10473);
nand U11462 (N_11462,N_9008,N_9897);
nand U11463 (N_11463,N_10493,N_10066);
or U11464 (N_11464,N_9520,N_9920);
nand U11465 (N_11465,N_9446,N_9486);
nand U11466 (N_11466,N_9369,N_9450);
or U11467 (N_11467,N_9850,N_10384);
or U11468 (N_11468,N_10188,N_10112);
nor U11469 (N_11469,N_9500,N_9098);
or U11470 (N_11470,N_10294,N_9894);
or U11471 (N_11471,N_9883,N_10042);
nor U11472 (N_11472,N_10266,N_9965);
or U11473 (N_11473,N_9871,N_9180);
nand U11474 (N_11474,N_9340,N_10005);
and U11475 (N_11475,N_9484,N_10190);
xor U11476 (N_11476,N_9238,N_10307);
or U11477 (N_11477,N_9570,N_9946);
or U11478 (N_11478,N_9414,N_9117);
or U11479 (N_11479,N_10487,N_9579);
and U11480 (N_11480,N_9987,N_9016);
and U11481 (N_11481,N_9294,N_9557);
nor U11482 (N_11482,N_10420,N_10308);
nor U11483 (N_11483,N_10341,N_9266);
nand U11484 (N_11484,N_9681,N_9884);
or U11485 (N_11485,N_9350,N_10469);
nor U11486 (N_11486,N_9854,N_10173);
nor U11487 (N_11487,N_9005,N_9552);
nor U11488 (N_11488,N_10460,N_9533);
nor U11489 (N_11489,N_9989,N_9459);
and U11490 (N_11490,N_10269,N_10231);
nand U11491 (N_11491,N_9960,N_10093);
and U11492 (N_11492,N_10046,N_9516);
and U11493 (N_11493,N_10255,N_9408);
or U11494 (N_11494,N_9429,N_10112);
xor U11495 (N_11495,N_9515,N_10304);
or U11496 (N_11496,N_9792,N_10461);
nand U11497 (N_11497,N_9991,N_9788);
nor U11498 (N_11498,N_9568,N_9129);
xor U11499 (N_11499,N_9125,N_9171);
and U11500 (N_11500,N_10303,N_9380);
or U11501 (N_11501,N_9260,N_9663);
and U11502 (N_11502,N_10200,N_9433);
and U11503 (N_11503,N_10085,N_9665);
nor U11504 (N_11504,N_9452,N_9197);
or U11505 (N_11505,N_10318,N_9070);
and U11506 (N_11506,N_9355,N_10450);
and U11507 (N_11507,N_9470,N_9954);
xnor U11508 (N_11508,N_10483,N_10238);
nor U11509 (N_11509,N_10249,N_10014);
and U11510 (N_11510,N_10177,N_9775);
or U11511 (N_11511,N_9637,N_10238);
and U11512 (N_11512,N_9716,N_10018);
and U11513 (N_11513,N_10009,N_10376);
or U11514 (N_11514,N_9800,N_10244);
nor U11515 (N_11515,N_9404,N_9232);
and U11516 (N_11516,N_9103,N_9927);
nand U11517 (N_11517,N_10145,N_10363);
nor U11518 (N_11518,N_9949,N_9640);
and U11519 (N_11519,N_10157,N_9846);
or U11520 (N_11520,N_10373,N_9809);
nand U11521 (N_11521,N_9652,N_9548);
nor U11522 (N_11522,N_10183,N_10029);
nor U11523 (N_11523,N_10332,N_9074);
and U11524 (N_11524,N_10453,N_9649);
nor U11525 (N_11525,N_10050,N_9909);
or U11526 (N_11526,N_10200,N_9811);
or U11527 (N_11527,N_10402,N_9219);
nand U11528 (N_11528,N_9789,N_9966);
and U11529 (N_11529,N_10219,N_9252);
or U11530 (N_11530,N_10274,N_9992);
nor U11531 (N_11531,N_9355,N_10033);
nor U11532 (N_11532,N_9248,N_10357);
or U11533 (N_11533,N_9674,N_9586);
nor U11534 (N_11534,N_9687,N_9578);
or U11535 (N_11535,N_10214,N_10267);
and U11536 (N_11536,N_10297,N_10176);
nand U11537 (N_11537,N_9289,N_9590);
and U11538 (N_11538,N_10366,N_9494);
nand U11539 (N_11539,N_10490,N_9097);
nand U11540 (N_11540,N_9499,N_10327);
nor U11541 (N_11541,N_9034,N_9720);
and U11542 (N_11542,N_10245,N_9230);
nand U11543 (N_11543,N_10394,N_9956);
nor U11544 (N_11544,N_10320,N_10241);
or U11545 (N_11545,N_10248,N_9798);
and U11546 (N_11546,N_10018,N_9966);
nand U11547 (N_11547,N_9873,N_9567);
and U11548 (N_11548,N_9307,N_9196);
or U11549 (N_11549,N_9506,N_9229);
and U11550 (N_11550,N_9406,N_9339);
nor U11551 (N_11551,N_9226,N_9531);
nor U11552 (N_11552,N_9391,N_10089);
nand U11553 (N_11553,N_9222,N_9812);
and U11554 (N_11554,N_9533,N_9488);
nand U11555 (N_11555,N_9439,N_9091);
nor U11556 (N_11556,N_9194,N_9683);
and U11557 (N_11557,N_9647,N_10459);
nand U11558 (N_11558,N_9508,N_9098);
and U11559 (N_11559,N_9215,N_9014);
and U11560 (N_11560,N_9377,N_9065);
and U11561 (N_11561,N_9709,N_9475);
xor U11562 (N_11562,N_9168,N_9029);
nor U11563 (N_11563,N_9884,N_10011);
xor U11564 (N_11564,N_9739,N_9275);
nand U11565 (N_11565,N_9795,N_9397);
nand U11566 (N_11566,N_9247,N_9972);
nand U11567 (N_11567,N_9437,N_10172);
nor U11568 (N_11568,N_9392,N_10147);
or U11569 (N_11569,N_9499,N_9274);
or U11570 (N_11570,N_10453,N_10075);
xnor U11571 (N_11571,N_9684,N_9787);
and U11572 (N_11572,N_9839,N_10027);
xnor U11573 (N_11573,N_9523,N_9460);
xor U11574 (N_11574,N_9723,N_10420);
xor U11575 (N_11575,N_10183,N_9408);
or U11576 (N_11576,N_10159,N_10404);
xnor U11577 (N_11577,N_10352,N_9370);
nand U11578 (N_11578,N_9312,N_10105);
and U11579 (N_11579,N_9922,N_10219);
or U11580 (N_11580,N_10071,N_9493);
nor U11581 (N_11581,N_9146,N_10203);
nor U11582 (N_11582,N_10469,N_9925);
nor U11583 (N_11583,N_9739,N_9235);
nor U11584 (N_11584,N_10262,N_9833);
and U11585 (N_11585,N_9586,N_9652);
or U11586 (N_11586,N_9371,N_10171);
or U11587 (N_11587,N_10450,N_10362);
and U11588 (N_11588,N_9955,N_10040);
nand U11589 (N_11589,N_9199,N_9560);
or U11590 (N_11590,N_10415,N_9105);
nor U11591 (N_11591,N_9432,N_10189);
and U11592 (N_11592,N_9307,N_9593);
xor U11593 (N_11593,N_9582,N_9015);
and U11594 (N_11594,N_10094,N_9807);
nand U11595 (N_11595,N_10444,N_9580);
xnor U11596 (N_11596,N_9236,N_10451);
nand U11597 (N_11597,N_9213,N_10452);
or U11598 (N_11598,N_9275,N_9998);
and U11599 (N_11599,N_9589,N_10451);
or U11600 (N_11600,N_9082,N_9652);
and U11601 (N_11601,N_9989,N_9732);
and U11602 (N_11602,N_9313,N_10126);
nor U11603 (N_11603,N_9122,N_10339);
nand U11604 (N_11604,N_10345,N_10096);
or U11605 (N_11605,N_10468,N_9829);
or U11606 (N_11606,N_9508,N_10483);
nor U11607 (N_11607,N_10145,N_10004);
xnor U11608 (N_11608,N_10186,N_9222);
nand U11609 (N_11609,N_9259,N_9598);
nor U11610 (N_11610,N_9497,N_9124);
and U11611 (N_11611,N_10036,N_9662);
or U11612 (N_11612,N_9353,N_9438);
and U11613 (N_11613,N_10041,N_9511);
nand U11614 (N_11614,N_9277,N_9201);
and U11615 (N_11615,N_10080,N_10144);
nor U11616 (N_11616,N_9982,N_9401);
nor U11617 (N_11617,N_10306,N_9513);
and U11618 (N_11618,N_9222,N_10439);
xor U11619 (N_11619,N_9363,N_9134);
nor U11620 (N_11620,N_9754,N_10059);
and U11621 (N_11621,N_9739,N_9922);
or U11622 (N_11622,N_9537,N_9630);
nor U11623 (N_11623,N_9731,N_9423);
nor U11624 (N_11624,N_10241,N_9029);
nor U11625 (N_11625,N_10162,N_9565);
nand U11626 (N_11626,N_9259,N_10351);
nor U11627 (N_11627,N_10233,N_10337);
nand U11628 (N_11628,N_10266,N_9105);
and U11629 (N_11629,N_9727,N_9134);
xnor U11630 (N_11630,N_9266,N_10017);
nand U11631 (N_11631,N_10348,N_9508);
and U11632 (N_11632,N_9383,N_9651);
or U11633 (N_11633,N_10480,N_10372);
nand U11634 (N_11634,N_10443,N_10290);
or U11635 (N_11635,N_9914,N_10010);
nor U11636 (N_11636,N_9719,N_10067);
and U11637 (N_11637,N_9399,N_9731);
nand U11638 (N_11638,N_9637,N_9445);
nand U11639 (N_11639,N_10017,N_9073);
and U11640 (N_11640,N_10395,N_9211);
nand U11641 (N_11641,N_9527,N_9436);
or U11642 (N_11642,N_10073,N_9652);
or U11643 (N_11643,N_10201,N_10278);
nor U11644 (N_11644,N_9551,N_9043);
nand U11645 (N_11645,N_10346,N_9370);
nand U11646 (N_11646,N_9659,N_9679);
nor U11647 (N_11647,N_9147,N_10008);
or U11648 (N_11648,N_10445,N_10288);
xnor U11649 (N_11649,N_9435,N_9959);
xor U11650 (N_11650,N_9519,N_10163);
or U11651 (N_11651,N_10401,N_9983);
nor U11652 (N_11652,N_9584,N_9243);
and U11653 (N_11653,N_9374,N_10209);
and U11654 (N_11654,N_10411,N_10045);
nor U11655 (N_11655,N_9591,N_9692);
nand U11656 (N_11656,N_9031,N_9432);
and U11657 (N_11657,N_9554,N_10376);
or U11658 (N_11658,N_10299,N_10477);
nor U11659 (N_11659,N_9094,N_10119);
xor U11660 (N_11660,N_10383,N_9890);
and U11661 (N_11661,N_9177,N_9141);
or U11662 (N_11662,N_9310,N_9998);
and U11663 (N_11663,N_9061,N_9584);
nand U11664 (N_11664,N_9844,N_9929);
nand U11665 (N_11665,N_10287,N_9566);
xnor U11666 (N_11666,N_9539,N_9753);
or U11667 (N_11667,N_10041,N_9922);
and U11668 (N_11668,N_9767,N_10000);
or U11669 (N_11669,N_9196,N_9649);
nor U11670 (N_11670,N_9719,N_10237);
nor U11671 (N_11671,N_9973,N_9226);
or U11672 (N_11672,N_9318,N_10350);
or U11673 (N_11673,N_10319,N_9190);
nand U11674 (N_11674,N_10289,N_9045);
nor U11675 (N_11675,N_10307,N_9348);
or U11676 (N_11676,N_9145,N_9312);
nor U11677 (N_11677,N_9100,N_9533);
and U11678 (N_11678,N_9779,N_10309);
and U11679 (N_11679,N_9799,N_9329);
or U11680 (N_11680,N_10327,N_10212);
nor U11681 (N_11681,N_9168,N_10416);
or U11682 (N_11682,N_9393,N_9630);
nand U11683 (N_11683,N_10228,N_9657);
and U11684 (N_11684,N_10487,N_9572);
nor U11685 (N_11685,N_10029,N_9865);
nor U11686 (N_11686,N_9526,N_9321);
nor U11687 (N_11687,N_10165,N_10440);
or U11688 (N_11688,N_9582,N_10107);
nor U11689 (N_11689,N_9681,N_9832);
or U11690 (N_11690,N_9154,N_10337);
nor U11691 (N_11691,N_10428,N_9725);
and U11692 (N_11692,N_9602,N_9264);
and U11693 (N_11693,N_10354,N_9486);
xor U11694 (N_11694,N_10423,N_9819);
and U11695 (N_11695,N_9296,N_9880);
nand U11696 (N_11696,N_10381,N_9259);
or U11697 (N_11697,N_10461,N_10053);
or U11698 (N_11698,N_10291,N_9968);
or U11699 (N_11699,N_9654,N_9724);
nand U11700 (N_11700,N_9102,N_9947);
and U11701 (N_11701,N_10302,N_9087);
and U11702 (N_11702,N_9421,N_9314);
or U11703 (N_11703,N_9839,N_10123);
and U11704 (N_11704,N_9202,N_9148);
and U11705 (N_11705,N_10407,N_9616);
xor U11706 (N_11706,N_10031,N_9283);
nor U11707 (N_11707,N_10158,N_9896);
or U11708 (N_11708,N_9187,N_9594);
or U11709 (N_11709,N_9622,N_10339);
and U11710 (N_11710,N_9719,N_9933);
nand U11711 (N_11711,N_9697,N_9605);
or U11712 (N_11712,N_10082,N_9782);
nor U11713 (N_11713,N_9085,N_9020);
or U11714 (N_11714,N_9569,N_9467);
nand U11715 (N_11715,N_9785,N_9377);
and U11716 (N_11716,N_10187,N_10241);
or U11717 (N_11717,N_9579,N_9372);
nor U11718 (N_11718,N_9177,N_9737);
xor U11719 (N_11719,N_9563,N_9122);
and U11720 (N_11720,N_9078,N_9124);
xnor U11721 (N_11721,N_9578,N_10308);
nand U11722 (N_11722,N_9365,N_9337);
or U11723 (N_11723,N_9101,N_10233);
and U11724 (N_11724,N_9311,N_9398);
and U11725 (N_11725,N_10388,N_9492);
and U11726 (N_11726,N_10381,N_9366);
nand U11727 (N_11727,N_10287,N_9508);
xor U11728 (N_11728,N_9293,N_10201);
or U11729 (N_11729,N_9572,N_10152);
nand U11730 (N_11730,N_10100,N_10416);
nand U11731 (N_11731,N_9011,N_9303);
or U11732 (N_11732,N_9427,N_10189);
xnor U11733 (N_11733,N_9466,N_9981);
and U11734 (N_11734,N_10454,N_10316);
or U11735 (N_11735,N_9323,N_9436);
nand U11736 (N_11736,N_9068,N_9018);
or U11737 (N_11737,N_9418,N_9752);
and U11738 (N_11738,N_9263,N_9200);
and U11739 (N_11739,N_10493,N_9353);
and U11740 (N_11740,N_9680,N_9650);
xor U11741 (N_11741,N_10186,N_9779);
nand U11742 (N_11742,N_9875,N_9890);
nand U11743 (N_11743,N_9030,N_9685);
and U11744 (N_11744,N_10268,N_9984);
nor U11745 (N_11745,N_10300,N_9433);
and U11746 (N_11746,N_9612,N_10387);
nand U11747 (N_11747,N_9815,N_9265);
nor U11748 (N_11748,N_9661,N_9087);
and U11749 (N_11749,N_9881,N_10328);
nor U11750 (N_11750,N_10179,N_9948);
or U11751 (N_11751,N_9511,N_10115);
and U11752 (N_11752,N_10399,N_10434);
xnor U11753 (N_11753,N_9448,N_9811);
and U11754 (N_11754,N_9774,N_9285);
nand U11755 (N_11755,N_10218,N_10055);
xor U11756 (N_11756,N_9544,N_10239);
or U11757 (N_11757,N_10210,N_9578);
nor U11758 (N_11758,N_9913,N_10477);
nand U11759 (N_11759,N_9390,N_9268);
nor U11760 (N_11760,N_9334,N_9158);
or U11761 (N_11761,N_9914,N_10307);
nor U11762 (N_11762,N_9580,N_9791);
or U11763 (N_11763,N_9985,N_9221);
nor U11764 (N_11764,N_9400,N_9596);
nor U11765 (N_11765,N_10200,N_10098);
nor U11766 (N_11766,N_10140,N_9463);
or U11767 (N_11767,N_9501,N_9154);
or U11768 (N_11768,N_10155,N_9434);
and U11769 (N_11769,N_9644,N_9989);
nor U11770 (N_11770,N_9631,N_9539);
nand U11771 (N_11771,N_9768,N_9758);
nand U11772 (N_11772,N_9282,N_9196);
or U11773 (N_11773,N_10170,N_9331);
nand U11774 (N_11774,N_9010,N_9646);
nand U11775 (N_11775,N_9066,N_9857);
or U11776 (N_11776,N_10105,N_9474);
nand U11777 (N_11777,N_9519,N_9579);
nand U11778 (N_11778,N_10327,N_9547);
nand U11779 (N_11779,N_9258,N_9193);
nor U11780 (N_11780,N_9725,N_9415);
nor U11781 (N_11781,N_9256,N_9823);
xnor U11782 (N_11782,N_9276,N_10491);
xor U11783 (N_11783,N_9307,N_9424);
or U11784 (N_11784,N_10144,N_10167);
or U11785 (N_11785,N_9336,N_9475);
and U11786 (N_11786,N_10023,N_9346);
and U11787 (N_11787,N_9111,N_9633);
and U11788 (N_11788,N_10080,N_9553);
and U11789 (N_11789,N_10373,N_9154);
and U11790 (N_11790,N_9032,N_9746);
and U11791 (N_11791,N_9504,N_9752);
nor U11792 (N_11792,N_10324,N_10411);
or U11793 (N_11793,N_10436,N_10374);
or U11794 (N_11794,N_9676,N_9609);
or U11795 (N_11795,N_9116,N_9986);
nor U11796 (N_11796,N_9225,N_9365);
nor U11797 (N_11797,N_9293,N_9333);
and U11798 (N_11798,N_9718,N_10102);
nor U11799 (N_11799,N_10458,N_9533);
or U11800 (N_11800,N_10080,N_9365);
and U11801 (N_11801,N_10034,N_9975);
or U11802 (N_11802,N_9783,N_10213);
nor U11803 (N_11803,N_9120,N_10000);
and U11804 (N_11804,N_9880,N_10115);
and U11805 (N_11805,N_10424,N_9975);
or U11806 (N_11806,N_9563,N_9128);
or U11807 (N_11807,N_10470,N_9029);
nor U11808 (N_11808,N_9631,N_9945);
or U11809 (N_11809,N_9271,N_9625);
xor U11810 (N_11810,N_9031,N_10239);
nor U11811 (N_11811,N_9360,N_9160);
or U11812 (N_11812,N_9872,N_10275);
nand U11813 (N_11813,N_9976,N_9546);
nor U11814 (N_11814,N_10499,N_9095);
nand U11815 (N_11815,N_10245,N_10032);
nand U11816 (N_11816,N_9991,N_9548);
nand U11817 (N_11817,N_10038,N_10366);
and U11818 (N_11818,N_10396,N_9816);
nand U11819 (N_11819,N_9376,N_10048);
and U11820 (N_11820,N_10015,N_10338);
nor U11821 (N_11821,N_9186,N_10409);
nor U11822 (N_11822,N_9961,N_10365);
nand U11823 (N_11823,N_10181,N_9780);
nand U11824 (N_11824,N_9770,N_9749);
or U11825 (N_11825,N_9697,N_10076);
and U11826 (N_11826,N_9709,N_10214);
and U11827 (N_11827,N_10216,N_9288);
or U11828 (N_11828,N_9973,N_9005);
nor U11829 (N_11829,N_10107,N_10316);
or U11830 (N_11830,N_10115,N_9656);
nor U11831 (N_11831,N_9926,N_10028);
or U11832 (N_11832,N_9037,N_9554);
nand U11833 (N_11833,N_10138,N_10030);
or U11834 (N_11834,N_9906,N_10343);
nor U11835 (N_11835,N_9676,N_10241);
nand U11836 (N_11836,N_9319,N_9372);
or U11837 (N_11837,N_10387,N_9828);
or U11838 (N_11838,N_9054,N_9447);
or U11839 (N_11839,N_10335,N_10376);
nand U11840 (N_11840,N_10175,N_10313);
xnor U11841 (N_11841,N_9877,N_9919);
and U11842 (N_11842,N_10395,N_9174);
and U11843 (N_11843,N_9512,N_9143);
or U11844 (N_11844,N_10113,N_9943);
xor U11845 (N_11845,N_10072,N_9038);
nand U11846 (N_11846,N_9428,N_10240);
nor U11847 (N_11847,N_10263,N_9477);
or U11848 (N_11848,N_9815,N_10141);
and U11849 (N_11849,N_10112,N_9957);
nand U11850 (N_11850,N_10367,N_9827);
or U11851 (N_11851,N_9884,N_10400);
or U11852 (N_11852,N_9994,N_9222);
or U11853 (N_11853,N_9418,N_9540);
or U11854 (N_11854,N_9184,N_9635);
nor U11855 (N_11855,N_10423,N_9774);
and U11856 (N_11856,N_10228,N_9078);
nor U11857 (N_11857,N_9461,N_9043);
and U11858 (N_11858,N_9032,N_9869);
nor U11859 (N_11859,N_9977,N_9784);
xnor U11860 (N_11860,N_10220,N_9188);
or U11861 (N_11861,N_10218,N_9897);
or U11862 (N_11862,N_9832,N_9746);
and U11863 (N_11863,N_9715,N_10161);
nor U11864 (N_11864,N_10152,N_9048);
and U11865 (N_11865,N_10292,N_9493);
or U11866 (N_11866,N_10264,N_9193);
or U11867 (N_11867,N_9264,N_9714);
xor U11868 (N_11868,N_10103,N_9936);
and U11869 (N_11869,N_10292,N_9025);
nand U11870 (N_11870,N_9305,N_10305);
nor U11871 (N_11871,N_9907,N_9723);
xor U11872 (N_11872,N_9110,N_9238);
and U11873 (N_11873,N_9759,N_10382);
and U11874 (N_11874,N_9664,N_10039);
nand U11875 (N_11875,N_9051,N_9986);
or U11876 (N_11876,N_9193,N_9046);
nand U11877 (N_11877,N_10076,N_9279);
and U11878 (N_11878,N_10388,N_10396);
or U11879 (N_11879,N_9071,N_10344);
or U11880 (N_11880,N_10244,N_9459);
and U11881 (N_11881,N_9053,N_10350);
nand U11882 (N_11882,N_10230,N_10432);
nand U11883 (N_11883,N_10126,N_10350);
and U11884 (N_11884,N_9425,N_10436);
and U11885 (N_11885,N_10471,N_9377);
and U11886 (N_11886,N_10055,N_9888);
nand U11887 (N_11887,N_9244,N_9744);
or U11888 (N_11888,N_9364,N_10199);
nand U11889 (N_11889,N_9013,N_9378);
nand U11890 (N_11890,N_9694,N_10424);
nand U11891 (N_11891,N_10241,N_10088);
nand U11892 (N_11892,N_9961,N_9395);
and U11893 (N_11893,N_9502,N_10296);
or U11894 (N_11894,N_9004,N_10199);
or U11895 (N_11895,N_9534,N_10057);
and U11896 (N_11896,N_9828,N_9695);
or U11897 (N_11897,N_9096,N_10095);
nor U11898 (N_11898,N_9502,N_10250);
nor U11899 (N_11899,N_9548,N_9928);
nor U11900 (N_11900,N_10198,N_9280);
xor U11901 (N_11901,N_9468,N_9801);
or U11902 (N_11902,N_9198,N_10491);
nor U11903 (N_11903,N_9025,N_9939);
nor U11904 (N_11904,N_9764,N_9636);
nand U11905 (N_11905,N_9173,N_9322);
nand U11906 (N_11906,N_10272,N_9685);
or U11907 (N_11907,N_9612,N_9315);
xor U11908 (N_11908,N_9786,N_10345);
xor U11909 (N_11909,N_9182,N_9899);
nor U11910 (N_11910,N_9439,N_9307);
or U11911 (N_11911,N_9410,N_9515);
nand U11912 (N_11912,N_9085,N_10394);
and U11913 (N_11913,N_10149,N_9884);
nor U11914 (N_11914,N_9141,N_9973);
or U11915 (N_11915,N_9438,N_10312);
and U11916 (N_11916,N_9162,N_10085);
nand U11917 (N_11917,N_9671,N_9866);
and U11918 (N_11918,N_10370,N_9913);
and U11919 (N_11919,N_9477,N_10193);
nor U11920 (N_11920,N_10319,N_9314);
or U11921 (N_11921,N_9806,N_10081);
or U11922 (N_11922,N_9767,N_9286);
nor U11923 (N_11923,N_9204,N_9945);
xnor U11924 (N_11924,N_10361,N_9343);
or U11925 (N_11925,N_9685,N_10457);
and U11926 (N_11926,N_9928,N_9341);
nor U11927 (N_11927,N_9803,N_10478);
and U11928 (N_11928,N_10499,N_10384);
and U11929 (N_11929,N_9425,N_9400);
xor U11930 (N_11930,N_10064,N_9005);
nor U11931 (N_11931,N_9745,N_9416);
nand U11932 (N_11932,N_9332,N_10038);
nor U11933 (N_11933,N_10495,N_10243);
xor U11934 (N_11934,N_9560,N_9903);
or U11935 (N_11935,N_9961,N_9946);
and U11936 (N_11936,N_9432,N_9630);
nor U11937 (N_11937,N_9802,N_9596);
nand U11938 (N_11938,N_9537,N_10321);
or U11939 (N_11939,N_9873,N_9165);
or U11940 (N_11940,N_9233,N_9675);
xnor U11941 (N_11941,N_10349,N_9514);
and U11942 (N_11942,N_9468,N_10099);
and U11943 (N_11943,N_9327,N_9994);
nor U11944 (N_11944,N_10326,N_9570);
or U11945 (N_11945,N_10189,N_9827);
nor U11946 (N_11946,N_9830,N_9804);
nor U11947 (N_11947,N_10050,N_9069);
or U11948 (N_11948,N_9699,N_10020);
nand U11949 (N_11949,N_9858,N_10303);
and U11950 (N_11950,N_9072,N_10243);
nor U11951 (N_11951,N_9865,N_9352);
nand U11952 (N_11952,N_9674,N_10228);
nor U11953 (N_11953,N_9575,N_9912);
and U11954 (N_11954,N_9632,N_10251);
or U11955 (N_11955,N_10413,N_9697);
or U11956 (N_11956,N_9713,N_10296);
nand U11957 (N_11957,N_9191,N_10022);
nand U11958 (N_11958,N_9459,N_9041);
nand U11959 (N_11959,N_10342,N_10338);
nand U11960 (N_11960,N_9319,N_9825);
xnor U11961 (N_11961,N_9376,N_9966);
or U11962 (N_11962,N_9561,N_9609);
and U11963 (N_11963,N_9114,N_10215);
or U11964 (N_11964,N_9999,N_10057);
nand U11965 (N_11965,N_9670,N_10148);
or U11966 (N_11966,N_9883,N_10196);
nand U11967 (N_11967,N_9996,N_9746);
or U11968 (N_11968,N_9686,N_9738);
nand U11969 (N_11969,N_9557,N_10484);
xor U11970 (N_11970,N_9263,N_9614);
nor U11971 (N_11971,N_10462,N_9700);
nor U11972 (N_11972,N_9415,N_9377);
and U11973 (N_11973,N_9551,N_10408);
or U11974 (N_11974,N_9032,N_10040);
nor U11975 (N_11975,N_10010,N_10456);
and U11976 (N_11976,N_9165,N_9706);
nor U11977 (N_11977,N_10288,N_9336);
xnor U11978 (N_11978,N_10337,N_10254);
nor U11979 (N_11979,N_9583,N_9520);
and U11980 (N_11980,N_9872,N_9593);
nor U11981 (N_11981,N_10298,N_9458);
or U11982 (N_11982,N_9839,N_9773);
nand U11983 (N_11983,N_9374,N_9634);
and U11984 (N_11984,N_9552,N_10367);
nand U11985 (N_11985,N_9426,N_9759);
and U11986 (N_11986,N_9826,N_9878);
nor U11987 (N_11987,N_9403,N_9470);
nor U11988 (N_11988,N_9618,N_9288);
or U11989 (N_11989,N_9949,N_10331);
nand U11990 (N_11990,N_9662,N_10178);
xnor U11991 (N_11991,N_9676,N_10219);
and U11992 (N_11992,N_9435,N_9980);
nor U11993 (N_11993,N_9100,N_9847);
and U11994 (N_11994,N_9071,N_9374);
and U11995 (N_11995,N_9723,N_9646);
xor U11996 (N_11996,N_9420,N_9775);
or U11997 (N_11997,N_10395,N_9516);
xor U11998 (N_11998,N_10316,N_9271);
nor U11999 (N_11999,N_9908,N_10071);
or U12000 (N_12000,N_10673,N_11395);
and U12001 (N_12001,N_10536,N_10665);
or U12002 (N_12002,N_11869,N_11127);
and U12003 (N_12003,N_11842,N_10624);
or U12004 (N_12004,N_11578,N_10614);
nand U12005 (N_12005,N_11651,N_11447);
and U12006 (N_12006,N_10883,N_10630);
and U12007 (N_12007,N_11524,N_11915);
and U12008 (N_12008,N_11239,N_11260);
nand U12009 (N_12009,N_11604,N_11184);
or U12010 (N_12010,N_11032,N_11766);
nor U12011 (N_12011,N_10593,N_11954);
or U12012 (N_12012,N_11509,N_10518);
nor U12013 (N_12013,N_10544,N_11164);
or U12014 (N_12014,N_10520,N_11534);
and U12015 (N_12015,N_11416,N_10540);
nor U12016 (N_12016,N_10831,N_11219);
nor U12017 (N_12017,N_11332,N_10558);
and U12018 (N_12018,N_11659,N_11507);
and U12019 (N_12019,N_10873,N_11760);
and U12020 (N_12020,N_11500,N_10833);
and U12021 (N_12021,N_10539,N_10810);
and U12022 (N_12022,N_10804,N_11006);
nand U12023 (N_12023,N_11292,N_11863);
nor U12024 (N_12024,N_11872,N_10839);
nor U12025 (N_12025,N_11448,N_10638);
or U12026 (N_12026,N_10506,N_10745);
and U12027 (N_12027,N_10629,N_11345);
nand U12028 (N_12028,N_11820,N_11951);
and U12029 (N_12029,N_11404,N_11862);
nor U12030 (N_12030,N_10602,N_10815);
nand U12031 (N_12031,N_10578,N_11178);
xor U12032 (N_12032,N_10879,N_11564);
nor U12033 (N_12033,N_11901,N_11190);
nor U12034 (N_12034,N_10557,N_11704);
and U12035 (N_12035,N_11249,N_11344);
nand U12036 (N_12036,N_11061,N_11394);
nand U12037 (N_12037,N_10853,N_10798);
or U12038 (N_12038,N_11286,N_11603);
and U12039 (N_12039,N_11402,N_11986);
nor U12040 (N_12040,N_10513,N_10774);
nor U12041 (N_12041,N_11386,N_11070);
and U12042 (N_12042,N_10947,N_11014);
and U12043 (N_12043,N_11538,N_11479);
or U12044 (N_12044,N_11478,N_11972);
or U12045 (N_12045,N_11263,N_11827);
xor U12046 (N_12046,N_10546,N_11100);
and U12047 (N_12047,N_11497,N_11090);
nand U12048 (N_12048,N_11795,N_10646);
or U12049 (N_12049,N_11493,N_11905);
nand U12050 (N_12050,N_10928,N_10829);
nand U12051 (N_12051,N_11600,N_11949);
or U12052 (N_12052,N_10858,N_11126);
nand U12053 (N_12053,N_10662,N_11441);
and U12054 (N_12054,N_11072,N_11811);
or U12055 (N_12055,N_10961,N_11642);
and U12056 (N_12056,N_10940,N_11148);
or U12057 (N_12057,N_11728,N_11839);
xor U12058 (N_12058,N_11025,N_10837);
and U12059 (N_12059,N_11873,N_11012);
and U12060 (N_12060,N_11318,N_10505);
or U12061 (N_12061,N_11443,N_10827);
and U12062 (N_12062,N_11082,N_11287);
and U12063 (N_12063,N_11160,N_11158);
and U12064 (N_12064,N_10889,N_11699);
and U12065 (N_12065,N_10819,N_10507);
and U12066 (N_12066,N_11661,N_11555);
or U12067 (N_12067,N_11514,N_11806);
nand U12068 (N_12068,N_11266,N_11994);
nand U12069 (N_12069,N_10692,N_11676);
nor U12070 (N_12070,N_11510,N_11993);
or U12071 (N_12071,N_10852,N_10666);
nor U12072 (N_12072,N_11034,N_11698);
nor U12073 (N_12073,N_11282,N_11755);
nand U12074 (N_12074,N_11613,N_10533);
and U12075 (N_12075,N_10575,N_10969);
or U12076 (N_12076,N_10750,N_11902);
or U12077 (N_12077,N_11171,N_11081);
or U12078 (N_12078,N_11307,N_10741);
nor U12079 (N_12079,N_10886,N_10586);
nand U12080 (N_12080,N_10746,N_11789);
nand U12081 (N_12081,N_11189,N_10753);
nand U12082 (N_12082,N_11474,N_11162);
nor U12083 (N_12083,N_11211,N_10863);
nor U12084 (N_12084,N_10790,N_11357);
nor U12085 (N_12085,N_11914,N_11637);
and U12086 (N_12086,N_11480,N_11275);
nand U12087 (N_12087,N_10749,N_10892);
or U12088 (N_12088,N_10901,N_11226);
xor U12089 (N_12089,N_11312,N_10949);
nand U12090 (N_12090,N_11597,N_10604);
nor U12091 (N_12091,N_11970,N_11876);
xnor U12092 (N_12092,N_11655,N_11744);
nand U12093 (N_12093,N_11750,N_11335);
or U12094 (N_12094,N_11317,N_11022);
xnor U12095 (N_12095,N_11439,N_11131);
and U12096 (N_12096,N_11383,N_11172);
nor U12097 (N_12097,N_11229,N_10991);
xor U12098 (N_12098,N_11955,N_11544);
and U12099 (N_12099,N_10502,N_11742);
or U12100 (N_12100,N_11390,N_11518);
xnor U12101 (N_12101,N_10887,N_11215);
nand U12102 (N_12102,N_11531,N_10581);
and U12103 (N_12103,N_11537,N_10836);
xnor U12104 (N_12104,N_11315,N_11907);
xnor U12105 (N_12105,N_11831,N_10519);
or U12106 (N_12106,N_11000,N_11320);
or U12107 (N_12107,N_11977,N_10881);
nand U12108 (N_12108,N_11461,N_11325);
and U12109 (N_12109,N_11973,N_10948);
nor U12110 (N_12110,N_11028,N_11107);
nor U12111 (N_12111,N_11669,N_11417);
or U12112 (N_12112,N_11846,N_10973);
nand U12113 (N_12113,N_10868,N_10797);
nand U12114 (N_12114,N_11965,N_11513);
nor U12115 (N_12115,N_11477,N_10628);
and U12116 (N_12116,N_11415,N_10545);
or U12117 (N_12117,N_11738,N_11236);
nor U12118 (N_12118,N_11828,N_11272);
and U12119 (N_12119,N_11910,N_11176);
nand U12120 (N_12120,N_11289,N_11773);
nand U12121 (N_12121,N_10743,N_11297);
xnor U12122 (N_12122,N_11817,N_11576);
and U12123 (N_12123,N_10998,N_11206);
nand U12124 (N_12124,N_10688,N_11724);
or U12125 (N_12125,N_11129,N_11739);
nor U12126 (N_12126,N_10914,N_11792);
xnor U12127 (N_12127,N_11671,N_11024);
nand U12128 (N_12128,N_10936,N_10697);
nand U12129 (N_12129,N_11971,N_11339);
nand U12130 (N_12130,N_11529,N_11109);
nand U12131 (N_12131,N_11656,N_11888);
nor U12132 (N_12132,N_11179,N_11618);
nor U12133 (N_12133,N_10521,N_11051);
nand U12134 (N_12134,N_11912,N_11035);
xnor U12135 (N_12135,N_10656,N_10786);
or U12136 (N_12136,N_10951,N_10993);
nand U12137 (N_12137,N_10997,N_11660);
and U12138 (N_12138,N_11662,N_11165);
or U12139 (N_12139,N_10554,N_11645);
and U12140 (N_12140,N_11619,N_10670);
nor U12141 (N_12141,N_10678,N_11393);
nand U12142 (N_12142,N_11548,N_11861);
or U12143 (N_12143,N_10825,N_11231);
xor U12144 (N_12144,N_11076,N_11288);
or U12145 (N_12145,N_10919,N_11033);
and U12146 (N_12146,N_10588,N_11533);
nor U12147 (N_12147,N_10632,N_11328);
and U12148 (N_12148,N_10959,N_11877);
nor U12149 (N_12149,N_11694,N_11128);
and U12150 (N_12150,N_11643,N_11909);
nor U12151 (N_12151,N_11865,N_11673);
or U12152 (N_12152,N_10732,N_11468);
or U12153 (N_12153,N_11341,N_11354);
and U12154 (N_12154,N_11042,N_11711);
and U12155 (N_12155,N_11336,N_11470);
nor U12156 (N_12156,N_11530,N_11264);
and U12157 (N_12157,N_11298,N_11064);
nand U12158 (N_12158,N_11648,N_10585);
or U12159 (N_12159,N_11403,N_11830);
nor U12160 (N_12160,N_11136,N_11405);
nor U12161 (N_12161,N_11269,N_10535);
and U12162 (N_12162,N_11496,N_11149);
and U12163 (N_12163,N_11095,N_11551);
or U12164 (N_12164,N_11209,N_11759);
xor U12165 (N_12165,N_10555,N_10626);
nand U12166 (N_12166,N_10615,N_11367);
or U12167 (N_12167,N_11557,N_10950);
and U12168 (N_12168,N_11701,N_11208);
and U12169 (N_12169,N_10767,N_11440);
nor U12170 (N_12170,N_11372,N_11799);
nand U12171 (N_12171,N_11052,N_11472);
xnor U12172 (N_12172,N_10542,N_11890);
nand U12173 (N_12173,N_11875,N_11521);
or U12174 (N_12174,N_11844,N_11324);
or U12175 (N_12175,N_11293,N_10933);
or U12176 (N_12176,N_11098,N_11803);
nand U12177 (N_12177,N_11684,N_11020);
nand U12178 (N_12178,N_11499,N_11774);
nand U12179 (N_12179,N_10974,N_10922);
and U12180 (N_12180,N_10598,N_11784);
and U12181 (N_12181,N_10757,N_10595);
xor U12182 (N_12182,N_11240,N_10576);
nand U12183 (N_12183,N_11733,N_11895);
nand U12184 (N_12184,N_10864,N_11996);
xnor U12185 (N_12185,N_11366,N_10992);
nand U12186 (N_12186,N_11767,N_11522);
or U12187 (N_12187,N_11657,N_11234);
and U12188 (N_12188,N_10913,N_11543);
nand U12189 (N_12189,N_11770,N_11174);
and U12190 (N_12190,N_11953,N_10764);
xor U12191 (N_12191,N_10685,N_11958);
nor U12192 (N_12192,N_10801,N_11550);
xnor U12193 (N_12193,N_11837,N_10996);
nor U12194 (N_12194,N_10738,N_10891);
nor U12195 (N_12195,N_11968,N_10846);
nand U12196 (N_12196,N_11703,N_10800);
nor U12197 (N_12197,N_10809,N_11714);
nor U12198 (N_12198,N_10736,N_10989);
or U12199 (N_12199,N_11140,N_11438);
nand U12200 (N_12200,N_11255,N_11900);
nand U12201 (N_12201,N_10577,N_10986);
nand U12202 (N_12202,N_10861,N_10562);
xor U12203 (N_12203,N_10907,N_11425);
or U12204 (N_12204,N_10828,N_10556);
nor U12205 (N_12205,N_11175,N_11170);
nand U12206 (N_12206,N_11571,N_10882);
and U12207 (N_12207,N_11399,N_11195);
or U12208 (N_12208,N_10918,N_11331);
and U12209 (N_12209,N_11668,N_11545);
and U12210 (N_12210,N_11960,N_10664);
and U12211 (N_12211,N_11607,N_11593);
xnor U12212 (N_12212,N_11808,N_11541);
nand U12213 (N_12213,N_11116,N_11678);
xnor U12214 (N_12214,N_10740,N_11343);
nand U12215 (N_12215,N_11225,N_10672);
nand U12216 (N_12216,N_10636,N_11369);
nor U12217 (N_12217,N_11486,N_11836);
or U12218 (N_12218,N_11523,N_11663);
xnor U12219 (N_12219,N_10500,N_11717);
or U12220 (N_12220,N_11097,N_11420);
nand U12221 (N_12221,N_11365,N_11303);
and U12222 (N_12222,N_11429,N_10705);
and U12223 (N_12223,N_11152,N_11482);
nor U12224 (N_12224,N_11535,N_11316);
nor U12225 (N_12225,N_10690,N_10841);
and U12226 (N_12226,N_11279,N_10702);
or U12227 (N_12227,N_11221,N_11281);
nor U12228 (N_12228,N_11265,N_11892);
nor U12229 (N_12229,N_10761,N_10931);
and U12230 (N_12230,N_11062,N_10768);
or U12231 (N_12231,N_10669,N_11974);
nor U12232 (N_12232,N_10954,N_10938);
nor U12233 (N_12233,N_10843,N_11185);
nand U12234 (N_12234,N_11137,N_10600);
nor U12235 (N_12235,N_11682,N_11104);
nor U12236 (N_12236,N_11205,N_11007);
and U12237 (N_12237,N_10683,N_11670);
nor U12238 (N_12238,N_11692,N_10718);
or U12239 (N_12239,N_11031,N_10802);
nand U12240 (N_12240,N_10862,N_11797);
nand U12241 (N_12241,N_11822,N_11408);
xnor U12242 (N_12242,N_11815,N_11793);
nor U12243 (N_12243,N_11777,N_11248);
nand U12244 (N_12244,N_10869,N_11199);
or U12245 (N_12245,N_11086,N_11961);
and U12246 (N_12246,N_11962,N_11526);
nand U12247 (N_12247,N_10842,N_11740);
and U12248 (N_12248,N_10522,N_10701);
nand U12249 (N_12249,N_11825,N_10780);
or U12250 (N_12250,N_11009,N_11159);
nand U12251 (N_12251,N_11193,N_11102);
nand U12252 (N_12252,N_11736,N_11640);
or U12253 (N_12253,N_11304,N_11099);
or U12254 (N_12254,N_11926,N_11725);
or U12255 (N_12255,N_10773,N_10728);
nand U12256 (N_12256,N_11922,N_11566);
nand U12257 (N_12257,N_11885,N_11485);
or U12258 (N_12258,N_10932,N_11616);
nor U12259 (N_12259,N_10679,N_11823);
xnor U12260 (N_12260,N_11410,N_11731);
nor U12261 (N_12261,N_11683,N_11580);
nand U12262 (N_12262,N_11299,N_11338);
nand U12263 (N_12263,N_11748,N_11038);
nor U12264 (N_12264,N_10971,N_11984);
or U12265 (N_12265,N_10980,N_11540);
or U12266 (N_12266,N_11586,N_10503);
xnor U12267 (N_12267,N_11726,N_11419);
xor U12268 (N_12268,N_10633,N_11351);
nor U12269 (N_12269,N_11672,N_11105);
or U12270 (N_12270,N_11920,N_11644);
nor U12271 (N_12271,N_11492,N_11558);
or U12272 (N_12272,N_10592,N_10523);
and U12273 (N_12273,N_11749,N_11720);
and U12274 (N_12274,N_11730,N_11380);
or U12275 (N_12275,N_10693,N_11021);
nand U12276 (N_12276,N_11039,N_11244);
nor U12277 (N_12277,N_11133,N_11602);
nor U12278 (N_12278,N_10634,N_10821);
nand U12279 (N_12279,N_10720,N_10958);
nand U12280 (N_12280,N_11911,N_10684);
or U12281 (N_12281,N_11924,N_11918);
and U12282 (N_12282,N_11860,N_11707);
xor U12283 (N_12283,N_11069,N_11569);
or U12284 (N_12284,N_11110,N_11611);
and U12285 (N_12285,N_11306,N_11464);
nor U12286 (N_12286,N_10777,N_10657);
nand U12287 (N_12287,N_10511,N_10985);
and U12288 (N_12288,N_11641,N_11202);
nand U12289 (N_12289,N_11764,N_10714);
and U12290 (N_12290,N_10724,N_10621);
xor U12291 (N_12291,N_11400,N_11783);
nand U12292 (N_12292,N_11452,N_11563);
nand U12293 (N_12293,N_11928,N_10984);
xnor U12294 (N_12294,N_11268,N_11310);
nand U12295 (N_12295,N_11291,N_10706);
nand U12296 (N_12296,N_11952,N_10917);
and U12297 (N_12297,N_11917,N_11101);
and U12298 (N_12298,N_11300,N_11483);
xnor U12299 (N_12299,N_11243,N_11756);
or U12300 (N_12300,N_10651,N_11330);
xnor U12301 (N_12301,N_11595,N_11285);
or U12302 (N_12302,N_11758,N_11192);
nand U12303 (N_12303,N_10784,N_11594);
nor U12304 (N_12304,N_11976,N_10906);
nor U12305 (N_12305,N_10515,N_11992);
nand U12306 (N_12306,N_11864,N_11183);
xnor U12307 (N_12307,N_11732,N_11718);
nor U12308 (N_12308,N_10880,N_10874);
xnor U12309 (N_12309,N_11003,N_11630);
nand U12310 (N_12310,N_10549,N_11786);
nand U12311 (N_12311,N_11891,N_11494);
and U12312 (N_12312,N_11841,N_11713);
or U12313 (N_12313,N_10855,N_11796);
nand U12314 (N_12314,N_11041,N_11379);
and U12315 (N_12315,N_11450,N_11598);
and U12316 (N_12316,N_10721,N_11194);
nand U12317 (N_12317,N_10972,N_10699);
or U12318 (N_12318,N_11204,N_11445);
nand U12319 (N_12319,N_10856,N_10710);
nand U12320 (N_12320,N_11906,N_10758);
nor U12321 (N_12321,N_10711,N_10960);
xnor U12322 (N_12322,N_11987,N_11368);
and U12323 (N_12323,N_11005,N_10893);
or U12324 (N_12324,N_10579,N_10983);
nand U12325 (N_12325,N_10655,N_11451);
nand U12326 (N_12326,N_10723,N_11633);
xnor U12327 (N_12327,N_11868,N_11167);
and U12328 (N_12328,N_11456,N_11040);
nand U12329 (N_12329,N_10799,N_11791);
nand U12330 (N_12330,N_11089,N_11964);
or U12331 (N_12331,N_10899,N_10622);
nor U12332 (N_12332,N_11359,N_10647);
xor U12333 (N_12333,N_11180,N_11412);
xnor U12334 (N_12334,N_11916,N_11455);
and U12335 (N_12335,N_11201,N_10704);
nor U12336 (N_12336,N_10995,N_10652);
and U12337 (N_12337,N_11824,N_11322);
or U12338 (N_12338,N_11991,N_11181);
or U12339 (N_12339,N_11151,N_10717);
nand U12340 (N_12340,N_11702,N_10781);
xnor U12341 (N_12341,N_11037,N_11547);
nand U12342 (N_12342,N_11030,N_11527);
nand U12343 (N_12343,N_11460,N_10909);
nor U12344 (N_12344,N_11919,N_11056);
or U12345 (N_12345,N_10610,N_10559);
and U12346 (N_12346,N_11942,N_11940);
and U12347 (N_12347,N_11622,N_11621);
nand U12348 (N_12348,N_11074,N_11060);
or U12349 (N_12349,N_11246,N_10830);
nor U12350 (N_12350,N_11398,N_11145);
xnor U12351 (N_12351,N_11163,N_10766);
or U12352 (N_12352,N_10751,N_11929);
nor U12353 (N_12353,N_11442,N_10694);
or U12354 (N_12354,N_11884,N_11690);
nand U12355 (N_12355,N_10682,N_11536);
and U12356 (N_12356,N_10953,N_11011);
xnor U12357 (N_12357,N_11115,N_11491);
nand U12358 (N_12358,N_10979,N_11004);
nor U12359 (N_12359,N_11583,N_11838);
nor U12360 (N_12360,N_11511,N_11308);
nor U12361 (N_12361,N_10851,N_11375);
nand U12362 (N_12362,N_10796,N_11309);
xnor U12363 (N_12363,N_10845,N_10824);
or U12364 (N_12364,N_10528,N_11989);
nand U12365 (N_12365,N_11591,N_11363);
nand U12366 (N_12366,N_11782,N_11634);
or U12367 (N_12367,N_10903,N_10658);
nor U12368 (N_12368,N_10640,N_10916);
and U12369 (N_12369,N_11614,N_10580);
nor U12370 (N_12370,N_11883,N_10820);
or U12371 (N_12371,N_10510,N_10987);
nor U12372 (N_12372,N_11016,N_10512);
and U12373 (N_12373,N_11719,N_11223);
and U12374 (N_12374,N_11314,N_11788);
nor U12375 (N_12375,N_10982,N_10978);
nor U12376 (N_12376,N_11997,N_10573);
or U12377 (N_12377,N_10650,N_11270);
xor U12378 (N_12378,N_11138,N_11427);
xnor U12379 (N_12379,N_11818,N_10504);
nor U12380 (N_12380,N_10617,N_10517);
xnor U12381 (N_12381,N_10920,N_11675);
or U12382 (N_12382,N_11346,N_11801);
nor U12383 (N_12383,N_11388,N_10748);
nand U12384 (N_12384,N_11938,N_11761);
nor U12385 (N_12385,N_11465,N_11722);
nand U12386 (N_12386,N_11358,N_11232);
and U12387 (N_12387,N_11124,N_11401);
nor U12388 (N_12388,N_10832,N_11352);
nand U12389 (N_12389,N_10771,N_10812);
or U12390 (N_12390,N_11233,N_11988);
or U12391 (N_12391,N_11257,N_11027);
nand U12392 (N_12392,N_11577,N_11686);
nor U12393 (N_12393,N_10508,N_11666);
nand U12394 (N_12394,N_11498,N_11068);
or U12395 (N_12395,N_10875,N_10547);
or U12396 (N_12396,N_10779,N_10594);
or U12397 (N_12397,N_11995,N_10962);
xnor U12398 (N_12398,N_11191,N_11826);
or U12399 (N_12399,N_11407,N_11026);
or U12400 (N_12400,N_10726,N_10596);
nand U12401 (N_12401,N_11156,N_11975);
or U12402 (N_12402,N_11625,N_10625);
and U12403 (N_12403,N_10859,N_11857);
nand U12404 (N_12404,N_10788,N_10795);
nor U12405 (N_12405,N_11146,N_11866);
nand U12406 (N_12406,N_10737,N_11259);
or U12407 (N_12407,N_10927,N_11957);
or U12408 (N_12408,N_10955,N_11927);
xnor U12409 (N_12409,N_10713,N_10527);
nor U12410 (N_12410,N_11045,N_10791);
or U12411 (N_12411,N_11851,N_10923);
nor U12412 (N_12412,N_11409,N_10538);
and U12413 (N_12413,N_11652,N_11834);
nor U12414 (N_12414,N_11639,N_11627);
and U12415 (N_12415,N_11220,N_10794);
or U12416 (N_12416,N_10867,N_11542);
and U12417 (N_12417,N_11305,N_11921);
or U12418 (N_12418,N_11350,N_11517);
and U12419 (N_12419,N_10770,N_11879);
or U12420 (N_12420,N_11210,N_11475);
nor U12421 (N_12421,N_10541,N_10835);
nor U12422 (N_12422,N_11349,N_11273);
and U12423 (N_12423,N_10618,N_11476);
and U12424 (N_12424,N_10696,N_10912);
xor U12425 (N_12425,N_11983,N_10895);
and U12426 (N_12426,N_10719,N_10725);
nand U12427 (N_12427,N_11334,N_11903);
nand U12428 (N_12428,N_10548,N_11561);
or U12429 (N_12429,N_11941,N_11821);
xor U12430 (N_12430,N_10756,N_10915);
and U12431 (N_12431,N_11262,N_10840);
xor U12432 (N_12432,N_10675,N_11284);
nor U12433 (N_12433,N_11319,N_10731);
nor U12434 (N_12434,N_10988,N_10560);
and U12435 (N_12435,N_11665,N_11525);
and U12436 (N_12436,N_10660,N_10681);
xnor U12437 (N_12437,N_11679,N_10952);
or U12438 (N_12438,N_10807,N_11753);
and U12439 (N_12439,N_10564,N_10667);
and U12440 (N_12440,N_11710,N_11946);
and U12441 (N_12441,N_11370,N_10957);
nor U12442 (N_12442,N_11010,N_11512);
nor U12443 (N_12443,N_11638,N_11721);
and U12444 (N_12444,N_11812,N_11200);
nand U12445 (N_12445,N_11626,N_11242);
nor U12446 (N_12446,N_10772,N_11337);
xor U12447 (N_12447,N_10934,N_11814);
or U12448 (N_12448,N_11067,N_11065);
and U12449 (N_12449,N_10567,N_11833);
nor U12450 (N_12450,N_11241,N_11685);
nand U12451 (N_12451,N_10734,N_11810);
xor U12452 (N_12452,N_11177,N_11588);
or U12453 (N_12453,N_11371,N_11624);
nor U12454 (N_12454,N_10956,N_11709);
and U12455 (N_12455,N_10589,N_11469);
and U12456 (N_12456,N_11013,N_10930);
nor U12457 (N_12457,N_10994,N_11055);
or U12458 (N_12458,N_10551,N_11743);
nor U12459 (N_12459,N_10550,N_11426);
nor U12460 (N_12460,N_11406,N_11778);
nand U12461 (N_12461,N_11276,N_10942);
nor U12462 (N_12462,N_10689,N_11214);
or U12463 (N_12463,N_11790,N_11886);
or U12464 (N_12464,N_11935,N_11768);
nand U12465 (N_12465,N_11182,N_10803);
nor U12466 (N_12466,N_11723,N_11813);
nand U12467 (N_12467,N_11230,N_11658);
and U12468 (N_12468,N_10531,N_10848);
and U12469 (N_12469,N_11579,N_10911);
nor U12470 (N_12470,N_11646,N_11487);
nor U12471 (N_12471,N_11867,N_11423);
xor U12472 (N_12472,N_10762,N_11463);
nor U12473 (N_12473,N_11381,N_11213);
nor U12474 (N_12474,N_10663,N_11340);
and U12475 (N_12475,N_11677,N_11467);
or U12476 (N_12476,N_10811,N_11508);
xnor U12477 (N_12477,N_11939,N_11094);
and U12478 (N_12478,N_11198,N_11757);
and U12479 (N_12479,N_11224,N_11687);
nand U12480 (N_12480,N_10698,N_11364);
or U12481 (N_12481,N_11913,N_10653);
or U12482 (N_12482,N_10872,N_10501);
or U12483 (N_12483,N_10876,N_11391);
nand U12484 (N_12484,N_10695,N_10752);
nor U12485 (N_12485,N_11080,N_11169);
nor U12486 (N_12486,N_10739,N_11734);
or U12487 (N_12487,N_10970,N_10525);
xor U12488 (N_12488,N_11894,N_11835);
xnor U12489 (N_12489,N_11904,N_11392);
nand U12490 (N_12490,N_10990,N_11490);
nand U12491 (N_12491,N_10910,N_10643);
or U12492 (N_12492,N_11313,N_11945);
and U12493 (N_12493,N_10759,N_10613);
nand U12494 (N_12494,N_10529,N_10661);
and U12495 (N_12495,N_11329,N_11847);
xor U12496 (N_12496,N_11628,N_11413);
or U12497 (N_12497,N_11396,N_11804);
and U12498 (N_12498,N_11188,N_11431);
nand U12499 (N_12499,N_11780,N_11157);
nor U12500 (N_12500,N_10516,N_10783);
nor U12501 (N_12501,N_11096,N_11150);
xnor U12502 (N_12502,N_11252,N_11017);
xor U12503 (N_12503,N_11397,N_10999);
nand U12504 (N_12504,N_11277,N_11382);
nand U12505 (N_12505,N_10644,N_10537);
nor U12506 (N_12506,N_10964,N_11301);
nor U12507 (N_12507,N_10716,N_11125);
xnor U12508 (N_12508,N_10754,N_10715);
nand U12509 (N_12509,N_10654,N_11751);
nor U12510 (N_12510,N_11258,N_11111);
or U12511 (N_12511,N_11959,N_10926);
nor U12512 (N_12512,N_10543,N_10894);
xnor U12513 (N_12513,N_11610,N_10945);
nor U12514 (N_12514,N_11896,N_11850);
xor U12515 (N_12515,N_11930,N_11765);
nand U12516 (N_12516,N_11855,N_11084);
and U12517 (N_12517,N_11931,N_11389);
nor U12518 (N_12518,N_10561,N_10608);
or U12519 (N_12519,N_11132,N_10671);
nor U12520 (N_12520,N_11187,N_11173);
xor U12521 (N_12521,N_10870,N_11735);
xnor U12522 (N_12522,N_11166,N_11119);
nor U12523 (N_12523,N_11466,N_11745);
nor U12524 (N_12524,N_11573,N_11649);
nand U12525 (N_12525,N_11362,N_11141);
or U12526 (N_12526,N_11484,N_10601);
or U12527 (N_12527,N_11256,N_11650);
nor U12528 (N_12528,N_10871,N_11592);
nand U12529 (N_12529,N_11473,N_11969);
nor U12530 (N_12530,N_11852,N_11002);
nand U12531 (N_12531,N_11635,N_11462);
xnor U12532 (N_12532,N_11274,N_11356);
or U12533 (N_12533,N_11587,N_11963);
nand U12534 (N_12534,N_10981,N_10967);
nand U12535 (N_12535,N_11623,N_11809);
and U12536 (N_12536,N_11434,N_11321);
nand U12537 (N_12537,N_10787,N_11361);
nand U12538 (N_12538,N_11087,N_10865);
xor U12539 (N_12539,N_11430,N_10691);
nor U12540 (N_12540,N_10849,N_11874);
nor U12541 (N_12541,N_11218,N_11436);
nor U12542 (N_12542,N_10792,N_11505);
xnor U12543 (N_12543,N_11043,N_11763);
nand U12544 (N_12544,N_11212,N_10847);
nor U12545 (N_12545,N_11854,N_11539);
and U12546 (N_12546,N_10582,N_11144);
nor U12547 (N_12547,N_11785,N_11932);
and U12548 (N_12548,N_11546,N_11565);
nand U12549 (N_12549,N_11503,N_10707);
nor U12550 (N_12550,N_10612,N_11008);
and U12551 (N_12551,N_11428,N_11794);
nand U12552 (N_12552,N_11348,N_10727);
or U12553 (N_12553,N_10937,N_10509);
nor U12554 (N_12554,N_11762,N_11695);
or U12555 (N_12555,N_11376,N_11870);
nand U12556 (N_12556,N_11023,N_11075);
xnor U12557 (N_12557,N_10939,N_11222);
nor U12558 (N_12558,N_11433,N_10645);
or U12559 (N_12559,N_10823,N_11899);
nor U12560 (N_12560,N_11947,N_11471);
nand U12561 (N_12561,N_11059,N_11982);
or U12562 (N_12562,N_11807,N_10941);
nor U12563 (N_12563,N_11373,N_11437);
nor U12564 (N_12564,N_10778,N_11130);
and U12565 (N_12565,N_11489,N_11606);
or U12566 (N_12566,N_11934,N_11681);
or U12567 (N_12567,N_11050,N_10925);
xor U12568 (N_12568,N_10860,N_11424);
nor U12569 (N_12569,N_11845,N_11168);
or U12570 (N_12570,N_11680,N_11048);
xnor U12571 (N_12571,N_11567,N_11556);
or U12572 (N_12572,N_10921,N_11515);
or U12573 (N_12573,N_10782,N_11418);
and U12574 (N_12574,N_11881,N_11458);
and U12575 (N_12575,N_11856,N_11647);
or U12576 (N_12576,N_10850,N_11520);
nor U12577 (N_12577,N_10877,N_11018);
nand U12578 (N_12578,N_10844,N_11077);
nor U12579 (N_12579,N_11998,N_11333);
nor U12580 (N_12580,N_11631,N_10712);
nor U12581 (N_12581,N_10703,N_10944);
nand U12582 (N_12582,N_11360,N_11092);
and U12583 (N_12583,N_11245,N_11449);
and U12584 (N_12584,N_10709,N_11950);
and U12585 (N_12585,N_11135,N_11605);
and U12586 (N_12586,N_11700,N_11504);
xnor U12587 (N_12587,N_10620,N_10817);
or U12588 (N_12588,N_10793,N_11121);
nor U12589 (N_12589,N_11697,N_11582);
or U12590 (N_12590,N_11029,N_10587);
nor U12591 (N_12591,N_11155,N_11290);
nand U12592 (N_12592,N_11294,N_10603);
and U12593 (N_12593,N_11549,N_11250);
and U12594 (N_12594,N_11235,N_11729);
or U12595 (N_12595,N_11754,N_11203);
nor U12596 (N_12596,N_10552,N_11502);
or U12597 (N_12597,N_10805,N_11590);
and U12598 (N_12598,N_10606,N_11771);
nor U12599 (N_12599,N_11374,N_11053);
and U12600 (N_12600,N_11207,N_10900);
or U12601 (N_12601,N_10963,N_11715);
nor U12602 (N_12602,N_10763,N_10609);
and U12603 (N_12603,N_10929,N_10563);
nor U12604 (N_12604,N_11385,N_10722);
nor U12605 (N_12605,N_10631,N_10571);
or U12606 (N_12606,N_11302,N_11800);
nor U12607 (N_12607,N_11446,N_11779);
nand U12608 (N_12608,N_11046,N_10687);
nand U12609 (N_12609,N_11805,N_10553);
or U12610 (N_12610,N_11066,N_11015);
and U12611 (N_12611,N_11858,N_10599);
nor U12612 (N_12612,N_11057,N_10530);
nand U12613 (N_12613,N_10637,N_10591);
and U12614 (N_12614,N_10908,N_10924);
and U12615 (N_12615,N_10884,N_11481);
nor U12616 (N_12616,N_10566,N_11143);
nor U12617 (N_12617,N_10708,N_10905);
and U12618 (N_12618,N_11384,N_10649);
nand U12619 (N_12619,N_11599,N_11693);
nor U12620 (N_12620,N_10686,N_11716);
nor U12621 (N_12621,N_11562,N_10648);
or U12622 (N_12622,N_10744,N_11897);
or U12623 (N_12623,N_11880,N_11843);
or U12624 (N_12624,N_11091,N_11044);
and U12625 (N_12625,N_11444,N_10730);
nand U12626 (N_12626,N_11459,N_11083);
nand U12627 (N_12627,N_11893,N_11454);
or U12628 (N_12628,N_11832,N_10816);
nor U12629 (N_12629,N_11123,N_11769);
nor U12630 (N_12630,N_10977,N_11691);
and U12631 (N_12631,N_10635,N_11142);
or U12632 (N_12632,N_11103,N_11568);
nand U12633 (N_12633,N_11047,N_11848);
and U12634 (N_12634,N_10584,N_10888);
and U12635 (N_12635,N_11271,N_11327);
nor U12636 (N_12636,N_10574,N_11326);
or U12637 (N_12637,N_11937,N_11139);
nand U12638 (N_12638,N_11887,N_10659);
and U12639 (N_12639,N_11516,N_10838);
and U12640 (N_12640,N_10570,N_10946);
or U12641 (N_12641,N_10775,N_10619);
xor U12642 (N_12642,N_11574,N_11608);
nor U12643 (N_12643,N_11708,N_11978);
nor U12644 (N_12644,N_11553,N_11036);
nor U12645 (N_12645,N_10733,N_11114);
nand U12646 (N_12646,N_11596,N_11653);
and U12647 (N_12647,N_11253,N_11636);
nor U12648 (N_12648,N_10642,N_11859);
and U12649 (N_12649,N_11933,N_11217);
and U12650 (N_12650,N_11387,N_11570);
and U12651 (N_12651,N_10611,N_10668);
xnor U12652 (N_12652,N_11966,N_10976);
nand U12653 (N_12653,N_11923,N_11985);
nor U12654 (N_12654,N_11688,N_11705);
xor U12655 (N_12655,N_10826,N_10700);
nand U12656 (N_12656,N_10806,N_10904);
nand U12657 (N_12657,N_11088,N_10532);
or U12658 (N_12658,N_10943,N_11457);
nor U12659 (N_12659,N_11377,N_11323);
nor U12660 (N_12660,N_11063,N_11979);
and U12661 (N_12661,N_11122,N_10524);
nor U12662 (N_12662,N_11113,N_10755);
nor U12663 (N_12663,N_10674,N_11079);
or U12664 (N_12664,N_11689,N_11154);
or U12665 (N_12665,N_11421,N_11295);
and U12666 (N_12666,N_10623,N_11967);
and U12667 (N_12667,N_11889,N_11085);
xor U12668 (N_12668,N_11247,N_10765);
nor U12669 (N_12669,N_11196,N_10569);
nor U12670 (N_12670,N_11519,N_11422);
or U12671 (N_12671,N_10866,N_11106);
nor U12672 (N_12672,N_10742,N_10814);
nor U12673 (N_12673,N_11667,N_11560);
nor U12674 (N_12674,N_10785,N_11787);
and U12675 (N_12675,N_11501,N_10568);
or U12676 (N_12676,N_10776,N_11802);
nand U12677 (N_12677,N_11664,N_11153);
nand U12678 (N_12678,N_10968,N_11572);
or U12679 (N_12679,N_11712,N_11251);
or U12680 (N_12680,N_11296,N_11581);
nand U12681 (N_12681,N_11001,N_11706);
or U12682 (N_12682,N_11999,N_11620);
xnor U12683 (N_12683,N_11696,N_11411);
nor U12684 (N_12684,N_11819,N_11532);
nand U12685 (N_12685,N_11615,N_11898);
nand U12686 (N_12686,N_11980,N_11981);
or U12687 (N_12687,N_11674,N_11197);
and U12688 (N_12688,N_11228,N_11882);
and U12689 (N_12689,N_11654,N_11435);
xnor U12690 (N_12690,N_11775,N_11353);
and U12691 (N_12691,N_11071,N_11816);
and U12692 (N_12692,N_11798,N_10822);
and U12693 (N_12693,N_11355,N_11776);
nor U12694 (N_12694,N_11073,N_10890);
nor U12695 (N_12695,N_10680,N_11584);
xnor U12696 (N_12696,N_11585,N_11632);
nor U12697 (N_12697,N_11849,N_10769);
and U12698 (N_12698,N_10885,N_11781);
nand U12699 (N_12699,N_11453,N_11054);
or U12700 (N_12700,N_11589,N_10935);
and U12701 (N_12701,N_11752,N_10597);
and U12702 (N_12702,N_11528,N_11414);
nor U12703 (N_12703,N_10898,N_11216);
nand U12704 (N_12704,N_11948,N_10818);
nor U12705 (N_12705,N_11267,N_11254);
nor U12706 (N_12706,N_11342,N_10789);
nand U12707 (N_12707,N_11552,N_11747);
nor U12708 (N_12708,N_11829,N_10590);
xor U12709 (N_12709,N_10808,N_10627);
xnor U12710 (N_12710,N_10677,N_11117);
nand U12711 (N_12711,N_11956,N_10735);
and U12712 (N_12712,N_11601,N_11108);
nand U12713 (N_12713,N_10896,N_11280);
or U12714 (N_12714,N_10975,N_11283);
nor U12715 (N_12715,N_11093,N_11609);
and U12716 (N_12716,N_11078,N_10813);
and U12717 (N_12717,N_11227,N_11741);
and U12718 (N_12718,N_10514,N_10641);
nor U12719 (N_12719,N_11871,N_10966);
nor U12720 (N_12720,N_10534,N_11853);
and U12721 (N_12721,N_11737,N_11772);
and U12722 (N_12722,N_11990,N_10583);
nand U12723 (N_12723,N_10607,N_10605);
nand U12724 (N_12724,N_11840,N_11559);
nor U12725 (N_12725,N_11186,N_11554);
and U12726 (N_12726,N_11058,N_11925);
or U12727 (N_12727,N_11261,N_11878);
or U12728 (N_12728,N_11147,N_10965);
nand U12729 (N_12729,N_10572,N_10565);
nor U12730 (N_12730,N_10616,N_10526);
or U12731 (N_12731,N_11432,N_11347);
and U12732 (N_12732,N_11936,N_10729);
and U12733 (N_12733,N_11311,N_11488);
and U12734 (N_12734,N_11049,N_10747);
nand U12735 (N_12735,N_10676,N_11120);
and U12736 (N_12736,N_11944,N_11134);
or U12737 (N_12737,N_11617,N_11112);
nand U12738 (N_12738,N_11746,N_11506);
nand U12739 (N_12739,N_11612,N_11495);
and U12740 (N_12740,N_11019,N_11378);
nor U12741 (N_12741,N_11161,N_10854);
nor U12742 (N_12742,N_10897,N_10902);
nand U12743 (N_12743,N_11575,N_11118);
and U12744 (N_12744,N_10834,N_11237);
and U12745 (N_12745,N_10878,N_10857);
or U12746 (N_12746,N_11278,N_11238);
or U12747 (N_12747,N_11629,N_10639);
or U12748 (N_12748,N_11908,N_11727);
xor U12749 (N_12749,N_11943,N_10760);
nand U12750 (N_12750,N_10950,N_11099);
or U12751 (N_12751,N_10753,N_11452);
nand U12752 (N_12752,N_11616,N_10947);
nor U12753 (N_12753,N_10954,N_11027);
or U12754 (N_12754,N_10540,N_10717);
nor U12755 (N_12755,N_11583,N_11436);
or U12756 (N_12756,N_11918,N_11738);
or U12757 (N_12757,N_11574,N_10858);
or U12758 (N_12758,N_10580,N_11102);
nor U12759 (N_12759,N_11858,N_11582);
or U12760 (N_12760,N_11326,N_10968);
or U12761 (N_12761,N_11709,N_11833);
and U12762 (N_12762,N_10593,N_11648);
xor U12763 (N_12763,N_10544,N_11045);
nand U12764 (N_12764,N_11254,N_10954);
nand U12765 (N_12765,N_10678,N_11521);
and U12766 (N_12766,N_11524,N_11946);
nand U12767 (N_12767,N_10594,N_11795);
nor U12768 (N_12768,N_11644,N_10576);
nand U12769 (N_12769,N_10628,N_11842);
nor U12770 (N_12770,N_11979,N_10625);
xnor U12771 (N_12771,N_11306,N_11979);
or U12772 (N_12772,N_10652,N_10647);
xnor U12773 (N_12773,N_10676,N_11246);
nor U12774 (N_12774,N_10750,N_10548);
or U12775 (N_12775,N_11107,N_11880);
or U12776 (N_12776,N_11716,N_10758);
nand U12777 (N_12777,N_10914,N_10668);
nor U12778 (N_12778,N_11246,N_11807);
and U12779 (N_12779,N_11529,N_10714);
and U12780 (N_12780,N_11450,N_11026);
and U12781 (N_12781,N_11080,N_11751);
or U12782 (N_12782,N_10997,N_11774);
nor U12783 (N_12783,N_11744,N_11629);
and U12784 (N_12784,N_10521,N_10656);
nand U12785 (N_12785,N_11546,N_11589);
nor U12786 (N_12786,N_11198,N_11620);
or U12787 (N_12787,N_11243,N_11456);
and U12788 (N_12788,N_10504,N_11213);
and U12789 (N_12789,N_10665,N_10756);
nor U12790 (N_12790,N_11031,N_11909);
or U12791 (N_12791,N_11245,N_10869);
nor U12792 (N_12792,N_11140,N_11541);
xnor U12793 (N_12793,N_11785,N_11575);
or U12794 (N_12794,N_10807,N_11360);
nor U12795 (N_12795,N_11187,N_11115);
nor U12796 (N_12796,N_11670,N_10712);
and U12797 (N_12797,N_11872,N_10990);
xor U12798 (N_12798,N_11998,N_10536);
nand U12799 (N_12799,N_11658,N_11678);
and U12800 (N_12800,N_11063,N_11995);
nor U12801 (N_12801,N_11954,N_11299);
xor U12802 (N_12802,N_10944,N_11602);
or U12803 (N_12803,N_11741,N_11161);
nand U12804 (N_12804,N_10733,N_11122);
nor U12805 (N_12805,N_11963,N_10729);
nor U12806 (N_12806,N_11931,N_10774);
nand U12807 (N_12807,N_11304,N_10551);
nor U12808 (N_12808,N_10699,N_11049);
nand U12809 (N_12809,N_11708,N_10900);
nor U12810 (N_12810,N_11993,N_10988);
nor U12811 (N_12811,N_11739,N_11733);
nor U12812 (N_12812,N_11560,N_10546);
nor U12813 (N_12813,N_10634,N_11710);
or U12814 (N_12814,N_11543,N_11512);
and U12815 (N_12815,N_11206,N_11599);
xnor U12816 (N_12816,N_11014,N_11976);
and U12817 (N_12817,N_10544,N_10601);
nand U12818 (N_12818,N_11119,N_11464);
or U12819 (N_12819,N_11808,N_11077);
xor U12820 (N_12820,N_11621,N_11140);
nand U12821 (N_12821,N_11121,N_11974);
nand U12822 (N_12822,N_11338,N_11186);
nor U12823 (N_12823,N_11420,N_11960);
or U12824 (N_12824,N_11962,N_11092);
xor U12825 (N_12825,N_11068,N_10932);
nand U12826 (N_12826,N_11022,N_10564);
nor U12827 (N_12827,N_10817,N_11157);
nor U12828 (N_12828,N_11841,N_11553);
nand U12829 (N_12829,N_10898,N_10830);
and U12830 (N_12830,N_11674,N_10788);
nand U12831 (N_12831,N_11012,N_11207);
and U12832 (N_12832,N_10858,N_11660);
nand U12833 (N_12833,N_11405,N_10766);
and U12834 (N_12834,N_11403,N_10581);
nor U12835 (N_12835,N_11873,N_10533);
nand U12836 (N_12836,N_10596,N_11602);
nor U12837 (N_12837,N_11841,N_11637);
and U12838 (N_12838,N_11133,N_10853);
xnor U12839 (N_12839,N_11849,N_11820);
or U12840 (N_12840,N_10763,N_11135);
nor U12841 (N_12841,N_10874,N_10546);
nor U12842 (N_12842,N_11203,N_10827);
nand U12843 (N_12843,N_11846,N_10733);
nor U12844 (N_12844,N_11585,N_11034);
or U12845 (N_12845,N_10696,N_11537);
nor U12846 (N_12846,N_11500,N_11639);
xor U12847 (N_12847,N_11000,N_11015);
and U12848 (N_12848,N_11290,N_11879);
or U12849 (N_12849,N_11428,N_11633);
and U12850 (N_12850,N_11802,N_10538);
and U12851 (N_12851,N_10639,N_10692);
or U12852 (N_12852,N_11181,N_10522);
or U12853 (N_12853,N_10964,N_11412);
nor U12854 (N_12854,N_11708,N_10614);
nand U12855 (N_12855,N_11254,N_10805);
and U12856 (N_12856,N_11797,N_10557);
or U12857 (N_12857,N_11161,N_11226);
or U12858 (N_12858,N_10594,N_10790);
and U12859 (N_12859,N_11229,N_11839);
nand U12860 (N_12860,N_11206,N_11226);
and U12861 (N_12861,N_11691,N_11546);
and U12862 (N_12862,N_11154,N_10824);
nand U12863 (N_12863,N_11866,N_11745);
nor U12864 (N_12864,N_11114,N_10871);
or U12865 (N_12865,N_11416,N_11876);
nor U12866 (N_12866,N_11707,N_10867);
and U12867 (N_12867,N_10594,N_11329);
nor U12868 (N_12868,N_10712,N_10940);
and U12869 (N_12869,N_11743,N_11573);
nor U12870 (N_12870,N_11589,N_10844);
and U12871 (N_12871,N_10859,N_11691);
nor U12872 (N_12872,N_10912,N_11818);
nand U12873 (N_12873,N_10858,N_10896);
nor U12874 (N_12874,N_11382,N_11837);
and U12875 (N_12875,N_11700,N_11342);
and U12876 (N_12876,N_11132,N_11283);
and U12877 (N_12877,N_11009,N_10926);
or U12878 (N_12878,N_11705,N_11642);
and U12879 (N_12879,N_11218,N_10641);
or U12880 (N_12880,N_11458,N_10878);
nor U12881 (N_12881,N_11504,N_10808);
nand U12882 (N_12882,N_11781,N_11059);
nand U12883 (N_12883,N_10827,N_10899);
and U12884 (N_12884,N_11633,N_11084);
nor U12885 (N_12885,N_10709,N_11841);
nor U12886 (N_12886,N_10658,N_10958);
nand U12887 (N_12887,N_11619,N_10776);
nor U12888 (N_12888,N_10826,N_11596);
nand U12889 (N_12889,N_11940,N_11017);
or U12890 (N_12890,N_11105,N_10959);
and U12891 (N_12891,N_11014,N_11431);
xor U12892 (N_12892,N_11167,N_11663);
or U12893 (N_12893,N_10540,N_11561);
nor U12894 (N_12894,N_10644,N_11784);
and U12895 (N_12895,N_11286,N_10857);
nor U12896 (N_12896,N_10697,N_10983);
and U12897 (N_12897,N_11707,N_10857);
and U12898 (N_12898,N_11124,N_10635);
and U12899 (N_12899,N_11204,N_11985);
or U12900 (N_12900,N_11685,N_11060);
or U12901 (N_12901,N_10951,N_10745);
and U12902 (N_12902,N_11104,N_10845);
nor U12903 (N_12903,N_10632,N_11834);
and U12904 (N_12904,N_11466,N_11034);
nand U12905 (N_12905,N_10814,N_11338);
or U12906 (N_12906,N_10998,N_11320);
nor U12907 (N_12907,N_11840,N_10691);
or U12908 (N_12908,N_10823,N_11256);
or U12909 (N_12909,N_11304,N_10696);
nor U12910 (N_12910,N_10683,N_11586);
and U12911 (N_12911,N_11130,N_11016);
or U12912 (N_12912,N_10560,N_11385);
and U12913 (N_12913,N_11156,N_11580);
nor U12914 (N_12914,N_11591,N_11098);
xnor U12915 (N_12915,N_11729,N_11057);
nand U12916 (N_12916,N_10641,N_11697);
or U12917 (N_12917,N_10938,N_10795);
and U12918 (N_12918,N_11788,N_10789);
and U12919 (N_12919,N_11679,N_10787);
nor U12920 (N_12920,N_10813,N_11591);
and U12921 (N_12921,N_10563,N_11066);
or U12922 (N_12922,N_11533,N_11720);
or U12923 (N_12923,N_11307,N_11780);
and U12924 (N_12924,N_11667,N_10807);
nor U12925 (N_12925,N_10836,N_11494);
nand U12926 (N_12926,N_11727,N_10517);
nor U12927 (N_12927,N_10784,N_11126);
nor U12928 (N_12928,N_10514,N_11471);
nand U12929 (N_12929,N_11789,N_10523);
or U12930 (N_12930,N_10558,N_10826);
and U12931 (N_12931,N_10536,N_11299);
nand U12932 (N_12932,N_11912,N_11504);
and U12933 (N_12933,N_11218,N_10572);
or U12934 (N_12934,N_11659,N_10737);
xor U12935 (N_12935,N_11680,N_10707);
nor U12936 (N_12936,N_11370,N_11183);
nand U12937 (N_12937,N_11692,N_11850);
and U12938 (N_12938,N_11616,N_11572);
nor U12939 (N_12939,N_11501,N_10907);
or U12940 (N_12940,N_11388,N_11234);
and U12941 (N_12941,N_11679,N_11352);
and U12942 (N_12942,N_11168,N_11466);
and U12943 (N_12943,N_11642,N_10870);
or U12944 (N_12944,N_11071,N_11204);
nand U12945 (N_12945,N_11709,N_11102);
xnor U12946 (N_12946,N_11911,N_11544);
xor U12947 (N_12947,N_11439,N_11063);
or U12948 (N_12948,N_11269,N_10524);
and U12949 (N_12949,N_11118,N_11358);
nand U12950 (N_12950,N_10851,N_11007);
and U12951 (N_12951,N_10614,N_10578);
and U12952 (N_12952,N_10506,N_11479);
nor U12953 (N_12953,N_11086,N_11282);
nand U12954 (N_12954,N_10787,N_11349);
or U12955 (N_12955,N_11917,N_10501);
or U12956 (N_12956,N_10777,N_10846);
or U12957 (N_12957,N_11848,N_11055);
nor U12958 (N_12958,N_11320,N_10568);
nor U12959 (N_12959,N_11834,N_11179);
and U12960 (N_12960,N_11314,N_10790);
xnor U12961 (N_12961,N_10619,N_11404);
xor U12962 (N_12962,N_11755,N_10606);
or U12963 (N_12963,N_11818,N_11351);
and U12964 (N_12964,N_11883,N_11933);
and U12965 (N_12965,N_10858,N_11671);
nor U12966 (N_12966,N_11272,N_11302);
and U12967 (N_12967,N_11169,N_11781);
nor U12968 (N_12968,N_11861,N_10651);
or U12969 (N_12969,N_10704,N_11227);
or U12970 (N_12970,N_11025,N_11888);
or U12971 (N_12971,N_11866,N_11349);
nor U12972 (N_12972,N_11392,N_11917);
nor U12973 (N_12973,N_11997,N_11221);
nor U12974 (N_12974,N_11335,N_11847);
nor U12975 (N_12975,N_11137,N_10868);
or U12976 (N_12976,N_11308,N_11862);
or U12977 (N_12977,N_10804,N_11581);
or U12978 (N_12978,N_10604,N_11463);
nor U12979 (N_12979,N_11001,N_10652);
or U12980 (N_12980,N_11625,N_11256);
and U12981 (N_12981,N_10859,N_11145);
or U12982 (N_12982,N_10608,N_11693);
and U12983 (N_12983,N_11427,N_11144);
or U12984 (N_12984,N_11377,N_11585);
and U12985 (N_12985,N_11603,N_11484);
nor U12986 (N_12986,N_11544,N_11563);
nor U12987 (N_12987,N_11800,N_10712);
and U12988 (N_12988,N_10775,N_10907);
or U12989 (N_12989,N_10969,N_11949);
and U12990 (N_12990,N_10639,N_11801);
nand U12991 (N_12991,N_11781,N_11408);
and U12992 (N_12992,N_11199,N_10967);
and U12993 (N_12993,N_11248,N_10514);
and U12994 (N_12994,N_10926,N_10544);
and U12995 (N_12995,N_11484,N_11314);
and U12996 (N_12996,N_11768,N_11904);
nand U12997 (N_12997,N_10755,N_11104);
nor U12998 (N_12998,N_11330,N_10732);
or U12999 (N_12999,N_11815,N_11078);
xnor U13000 (N_13000,N_11534,N_11314);
nand U13001 (N_13001,N_11111,N_11819);
nand U13002 (N_13002,N_10619,N_10831);
xnor U13003 (N_13003,N_10909,N_11294);
nand U13004 (N_13004,N_10500,N_10882);
nor U13005 (N_13005,N_11177,N_11252);
nand U13006 (N_13006,N_11201,N_11242);
xnor U13007 (N_13007,N_11028,N_11735);
and U13008 (N_13008,N_11400,N_11349);
and U13009 (N_13009,N_10935,N_11104);
nand U13010 (N_13010,N_11612,N_11345);
xor U13011 (N_13011,N_11996,N_11959);
and U13012 (N_13012,N_11568,N_10565);
nand U13013 (N_13013,N_10862,N_11425);
nor U13014 (N_13014,N_11356,N_11780);
nand U13015 (N_13015,N_10681,N_11129);
or U13016 (N_13016,N_11344,N_10531);
and U13017 (N_13017,N_11003,N_11625);
nor U13018 (N_13018,N_10699,N_10958);
nand U13019 (N_13019,N_11385,N_11981);
or U13020 (N_13020,N_11066,N_11077);
nor U13021 (N_13021,N_11547,N_11771);
nand U13022 (N_13022,N_11788,N_11016);
nand U13023 (N_13023,N_10741,N_10726);
or U13024 (N_13024,N_10742,N_10657);
nor U13025 (N_13025,N_11904,N_10971);
and U13026 (N_13026,N_11941,N_11331);
and U13027 (N_13027,N_11090,N_10829);
or U13028 (N_13028,N_11397,N_11644);
and U13029 (N_13029,N_10864,N_10938);
or U13030 (N_13030,N_10758,N_11985);
and U13031 (N_13031,N_11135,N_10647);
or U13032 (N_13032,N_10913,N_11949);
and U13033 (N_13033,N_11502,N_10948);
nand U13034 (N_13034,N_10712,N_10871);
nand U13035 (N_13035,N_11372,N_11371);
or U13036 (N_13036,N_11311,N_11757);
nand U13037 (N_13037,N_11096,N_11828);
or U13038 (N_13038,N_11414,N_11125);
and U13039 (N_13039,N_11262,N_11187);
nor U13040 (N_13040,N_11433,N_11591);
and U13041 (N_13041,N_10607,N_11053);
and U13042 (N_13042,N_11916,N_11415);
nand U13043 (N_13043,N_10781,N_11479);
xnor U13044 (N_13044,N_11246,N_11652);
nor U13045 (N_13045,N_10810,N_10545);
nand U13046 (N_13046,N_11916,N_11693);
nand U13047 (N_13047,N_10579,N_11012);
or U13048 (N_13048,N_11815,N_10990);
nor U13049 (N_13049,N_11247,N_10861);
nor U13050 (N_13050,N_10996,N_11546);
and U13051 (N_13051,N_11717,N_11307);
and U13052 (N_13052,N_11924,N_10777);
xnor U13053 (N_13053,N_11995,N_11865);
and U13054 (N_13054,N_11389,N_11235);
nand U13055 (N_13055,N_11284,N_11878);
xnor U13056 (N_13056,N_10710,N_11206);
nand U13057 (N_13057,N_10555,N_10942);
nand U13058 (N_13058,N_11113,N_10642);
xor U13059 (N_13059,N_10725,N_11430);
and U13060 (N_13060,N_11317,N_11239);
and U13061 (N_13061,N_11277,N_10720);
or U13062 (N_13062,N_11447,N_11861);
nor U13063 (N_13063,N_11023,N_10632);
nor U13064 (N_13064,N_11256,N_10558);
nor U13065 (N_13065,N_11559,N_11419);
xor U13066 (N_13066,N_11993,N_11054);
xor U13067 (N_13067,N_11413,N_10971);
or U13068 (N_13068,N_11847,N_10518);
and U13069 (N_13069,N_11111,N_11108);
or U13070 (N_13070,N_11354,N_11100);
xnor U13071 (N_13071,N_11748,N_11541);
nor U13072 (N_13072,N_10812,N_11260);
nor U13073 (N_13073,N_11976,N_11077);
nand U13074 (N_13074,N_11310,N_10759);
and U13075 (N_13075,N_10641,N_10738);
nor U13076 (N_13076,N_11385,N_11051);
and U13077 (N_13077,N_11549,N_11777);
and U13078 (N_13078,N_11499,N_10824);
xnor U13079 (N_13079,N_11474,N_11079);
or U13080 (N_13080,N_10938,N_11903);
or U13081 (N_13081,N_11471,N_11024);
or U13082 (N_13082,N_11318,N_11613);
nand U13083 (N_13083,N_10979,N_11533);
nor U13084 (N_13084,N_11240,N_11794);
or U13085 (N_13085,N_10705,N_11186);
and U13086 (N_13086,N_10690,N_11555);
nor U13087 (N_13087,N_10770,N_10784);
xnor U13088 (N_13088,N_11953,N_11382);
nor U13089 (N_13089,N_10804,N_11414);
and U13090 (N_13090,N_11915,N_10995);
xnor U13091 (N_13091,N_10555,N_10551);
and U13092 (N_13092,N_10737,N_11312);
nor U13093 (N_13093,N_11532,N_11781);
nor U13094 (N_13094,N_10714,N_11121);
and U13095 (N_13095,N_10921,N_11875);
and U13096 (N_13096,N_11494,N_11436);
nand U13097 (N_13097,N_11234,N_10580);
and U13098 (N_13098,N_10666,N_11403);
nand U13099 (N_13099,N_11613,N_11180);
nor U13100 (N_13100,N_11631,N_10879);
nand U13101 (N_13101,N_10548,N_11911);
and U13102 (N_13102,N_10903,N_10515);
xnor U13103 (N_13103,N_11593,N_10955);
nor U13104 (N_13104,N_10548,N_11639);
or U13105 (N_13105,N_11587,N_11964);
and U13106 (N_13106,N_11503,N_11311);
and U13107 (N_13107,N_10796,N_11048);
nor U13108 (N_13108,N_11445,N_10985);
xor U13109 (N_13109,N_10840,N_10922);
or U13110 (N_13110,N_10585,N_10899);
or U13111 (N_13111,N_10570,N_11360);
or U13112 (N_13112,N_11483,N_11548);
nor U13113 (N_13113,N_11827,N_11914);
nor U13114 (N_13114,N_10874,N_10831);
nand U13115 (N_13115,N_10861,N_11725);
or U13116 (N_13116,N_11308,N_11935);
or U13117 (N_13117,N_11384,N_11024);
xnor U13118 (N_13118,N_11104,N_10768);
nor U13119 (N_13119,N_11059,N_10846);
nor U13120 (N_13120,N_11328,N_11061);
and U13121 (N_13121,N_11690,N_11002);
nor U13122 (N_13122,N_11180,N_10877);
nand U13123 (N_13123,N_11583,N_10835);
and U13124 (N_13124,N_10627,N_11305);
xnor U13125 (N_13125,N_10811,N_11037);
and U13126 (N_13126,N_10538,N_11119);
nand U13127 (N_13127,N_10643,N_10939);
nor U13128 (N_13128,N_11050,N_11830);
or U13129 (N_13129,N_11634,N_10955);
xnor U13130 (N_13130,N_10903,N_10569);
nand U13131 (N_13131,N_11305,N_11609);
or U13132 (N_13132,N_11490,N_11526);
or U13133 (N_13133,N_11106,N_10751);
nand U13134 (N_13134,N_10582,N_11086);
nand U13135 (N_13135,N_11380,N_11396);
or U13136 (N_13136,N_11051,N_10738);
and U13137 (N_13137,N_11069,N_11217);
nand U13138 (N_13138,N_11525,N_11942);
nor U13139 (N_13139,N_11990,N_10598);
or U13140 (N_13140,N_11202,N_10721);
xnor U13141 (N_13141,N_11597,N_11248);
and U13142 (N_13142,N_11018,N_11479);
and U13143 (N_13143,N_11425,N_11445);
nor U13144 (N_13144,N_10779,N_11533);
xnor U13145 (N_13145,N_11091,N_11473);
nor U13146 (N_13146,N_10561,N_10827);
nand U13147 (N_13147,N_10795,N_10530);
and U13148 (N_13148,N_10860,N_11960);
or U13149 (N_13149,N_11140,N_10892);
nor U13150 (N_13150,N_11089,N_11503);
or U13151 (N_13151,N_11677,N_11234);
nor U13152 (N_13152,N_11687,N_11704);
nand U13153 (N_13153,N_11741,N_10665);
nor U13154 (N_13154,N_11728,N_11381);
nor U13155 (N_13155,N_10556,N_11740);
nor U13156 (N_13156,N_11999,N_10973);
nor U13157 (N_13157,N_11106,N_10902);
nor U13158 (N_13158,N_10835,N_11162);
or U13159 (N_13159,N_10654,N_10895);
nor U13160 (N_13160,N_11261,N_10538);
nand U13161 (N_13161,N_11260,N_11979);
nand U13162 (N_13162,N_11150,N_11287);
or U13163 (N_13163,N_11247,N_11681);
nand U13164 (N_13164,N_11593,N_11544);
or U13165 (N_13165,N_11772,N_11126);
nand U13166 (N_13166,N_10769,N_11870);
nor U13167 (N_13167,N_11628,N_10851);
and U13168 (N_13168,N_11974,N_11450);
or U13169 (N_13169,N_11185,N_11314);
and U13170 (N_13170,N_11894,N_11319);
nand U13171 (N_13171,N_11915,N_10696);
nor U13172 (N_13172,N_10709,N_11646);
or U13173 (N_13173,N_11045,N_11752);
nand U13174 (N_13174,N_11951,N_11859);
and U13175 (N_13175,N_10641,N_11381);
or U13176 (N_13176,N_11607,N_11372);
xor U13177 (N_13177,N_10869,N_11558);
and U13178 (N_13178,N_11470,N_11869);
nor U13179 (N_13179,N_11254,N_10723);
nor U13180 (N_13180,N_10507,N_11423);
nor U13181 (N_13181,N_10646,N_11022);
xnor U13182 (N_13182,N_10638,N_11200);
and U13183 (N_13183,N_11778,N_10888);
nand U13184 (N_13184,N_11759,N_10607);
and U13185 (N_13185,N_10666,N_11720);
or U13186 (N_13186,N_11937,N_11482);
nand U13187 (N_13187,N_11412,N_10521);
nand U13188 (N_13188,N_11010,N_10505);
or U13189 (N_13189,N_11381,N_10532);
nand U13190 (N_13190,N_10831,N_11402);
nand U13191 (N_13191,N_10527,N_11499);
or U13192 (N_13192,N_11468,N_10801);
nor U13193 (N_13193,N_10731,N_11745);
and U13194 (N_13194,N_11213,N_11556);
and U13195 (N_13195,N_10829,N_10549);
and U13196 (N_13196,N_10550,N_11263);
and U13197 (N_13197,N_10916,N_11414);
or U13198 (N_13198,N_11142,N_10538);
xor U13199 (N_13199,N_11333,N_11689);
nand U13200 (N_13200,N_11061,N_11135);
nand U13201 (N_13201,N_11263,N_11526);
xor U13202 (N_13202,N_11220,N_11065);
nor U13203 (N_13203,N_11962,N_11462);
and U13204 (N_13204,N_11991,N_11020);
or U13205 (N_13205,N_10586,N_11497);
or U13206 (N_13206,N_11206,N_11575);
or U13207 (N_13207,N_11488,N_10529);
and U13208 (N_13208,N_10771,N_11129);
and U13209 (N_13209,N_10784,N_11698);
nand U13210 (N_13210,N_10970,N_11197);
and U13211 (N_13211,N_11062,N_10985);
or U13212 (N_13212,N_10731,N_11029);
nor U13213 (N_13213,N_11607,N_11974);
nor U13214 (N_13214,N_10989,N_10655);
nor U13215 (N_13215,N_11715,N_10889);
xor U13216 (N_13216,N_11931,N_11783);
nand U13217 (N_13217,N_10567,N_11279);
xor U13218 (N_13218,N_11569,N_10517);
xor U13219 (N_13219,N_11114,N_11109);
nand U13220 (N_13220,N_11378,N_11350);
nor U13221 (N_13221,N_10555,N_10780);
or U13222 (N_13222,N_11393,N_10735);
nand U13223 (N_13223,N_11724,N_11325);
and U13224 (N_13224,N_10607,N_11986);
nand U13225 (N_13225,N_11614,N_10860);
nand U13226 (N_13226,N_11094,N_11810);
and U13227 (N_13227,N_11700,N_11833);
nand U13228 (N_13228,N_10567,N_11099);
nor U13229 (N_13229,N_10804,N_11025);
nand U13230 (N_13230,N_11837,N_10819);
nor U13231 (N_13231,N_11581,N_11290);
nor U13232 (N_13232,N_10737,N_11067);
nand U13233 (N_13233,N_10883,N_11869);
and U13234 (N_13234,N_11036,N_11328);
nor U13235 (N_13235,N_11988,N_10874);
nor U13236 (N_13236,N_11450,N_11837);
nor U13237 (N_13237,N_10903,N_11123);
xor U13238 (N_13238,N_10593,N_11274);
nand U13239 (N_13239,N_11122,N_11892);
or U13240 (N_13240,N_11927,N_11236);
or U13241 (N_13241,N_11767,N_11029);
nand U13242 (N_13242,N_11679,N_10507);
and U13243 (N_13243,N_10635,N_11730);
xor U13244 (N_13244,N_10837,N_10624);
nor U13245 (N_13245,N_11853,N_11943);
or U13246 (N_13246,N_11391,N_11074);
and U13247 (N_13247,N_10514,N_11274);
nand U13248 (N_13248,N_11228,N_11620);
and U13249 (N_13249,N_11683,N_11714);
nand U13250 (N_13250,N_11998,N_11014);
or U13251 (N_13251,N_11758,N_11230);
or U13252 (N_13252,N_10853,N_11076);
nor U13253 (N_13253,N_11670,N_10761);
nor U13254 (N_13254,N_11630,N_10907);
and U13255 (N_13255,N_11127,N_11120);
xnor U13256 (N_13256,N_10714,N_10765);
or U13257 (N_13257,N_11254,N_10711);
nand U13258 (N_13258,N_11046,N_11896);
and U13259 (N_13259,N_11758,N_11585);
and U13260 (N_13260,N_11693,N_11565);
xor U13261 (N_13261,N_11419,N_11409);
xor U13262 (N_13262,N_11403,N_11688);
xnor U13263 (N_13263,N_11055,N_11299);
and U13264 (N_13264,N_10991,N_10825);
or U13265 (N_13265,N_11819,N_11444);
nand U13266 (N_13266,N_11968,N_11804);
or U13267 (N_13267,N_11104,N_11827);
nor U13268 (N_13268,N_11960,N_11783);
nor U13269 (N_13269,N_11153,N_10728);
and U13270 (N_13270,N_11309,N_10718);
and U13271 (N_13271,N_11679,N_11845);
nor U13272 (N_13272,N_11795,N_11542);
xor U13273 (N_13273,N_11939,N_11845);
or U13274 (N_13274,N_10725,N_11612);
or U13275 (N_13275,N_11461,N_10756);
or U13276 (N_13276,N_11066,N_10843);
and U13277 (N_13277,N_11766,N_11553);
nor U13278 (N_13278,N_10759,N_10629);
or U13279 (N_13279,N_10925,N_10905);
and U13280 (N_13280,N_11108,N_11246);
nand U13281 (N_13281,N_10500,N_11334);
nor U13282 (N_13282,N_11727,N_10511);
and U13283 (N_13283,N_11628,N_11289);
nand U13284 (N_13284,N_11415,N_11548);
nand U13285 (N_13285,N_11890,N_10859);
and U13286 (N_13286,N_10768,N_10844);
and U13287 (N_13287,N_11099,N_11204);
xor U13288 (N_13288,N_10899,N_11612);
nor U13289 (N_13289,N_11141,N_10536);
nor U13290 (N_13290,N_11743,N_10597);
or U13291 (N_13291,N_11830,N_10711);
xor U13292 (N_13292,N_11882,N_11660);
or U13293 (N_13293,N_10887,N_10610);
and U13294 (N_13294,N_10657,N_11703);
and U13295 (N_13295,N_10991,N_10526);
and U13296 (N_13296,N_11533,N_11267);
and U13297 (N_13297,N_11064,N_11759);
and U13298 (N_13298,N_10604,N_11908);
or U13299 (N_13299,N_10618,N_10850);
nor U13300 (N_13300,N_11951,N_11578);
and U13301 (N_13301,N_11572,N_11947);
nand U13302 (N_13302,N_11520,N_11327);
nand U13303 (N_13303,N_11467,N_11609);
nand U13304 (N_13304,N_11626,N_10653);
or U13305 (N_13305,N_11915,N_11215);
and U13306 (N_13306,N_11564,N_10688);
nand U13307 (N_13307,N_11665,N_10940);
xnor U13308 (N_13308,N_10993,N_11538);
nand U13309 (N_13309,N_11404,N_10539);
nand U13310 (N_13310,N_10976,N_10797);
nor U13311 (N_13311,N_11756,N_11012);
and U13312 (N_13312,N_11546,N_10886);
nand U13313 (N_13313,N_10981,N_10595);
nor U13314 (N_13314,N_11435,N_11527);
and U13315 (N_13315,N_11238,N_10508);
and U13316 (N_13316,N_11585,N_11537);
and U13317 (N_13317,N_11394,N_10518);
nor U13318 (N_13318,N_11672,N_11721);
nor U13319 (N_13319,N_11638,N_11247);
and U13320 (N_13320,N_11026,N_10722);
and U13321 (N_13321,N_10939,N_11290);
or U13322 (N_13322,N_11933,N_11269);
or U13323 (N_13323,N_11065,N_11406);
nor U13324 (N_13324,N_11381,N_11058);
nor U13325 (N_13325,N_11465,N_11127);
and U13326 (N_13326,N_10755,N_10605);
xor U13327 (N_13327,N_10892,N_11644);
xor U13328 (N_13328,N_11663,N_11250);
nand U13329 (N_13329,N_11144,N_11459);
nor U13330 (N_13330,N_11347,N_10981);
nand U13331 (N_13331,N_11658,N_11713);
and U13332 (N_13332,N_10677,N_11219);
nand U13333 (N_13333,N_11308,N_11254);
or U13334 (N_13334,N_10666,N_11270);
nor U13335 (N_13335,N_11400,N_11740);
and U13336 (N_13336,N_11390,N_10882);
and U13337 (N_13337,N_11650,N_11087);
or U13338 (N_13338,N_10927,N_11236);
and U13339 (N_13339,N_11583,N_11351);
nor U13340 (N_13340,N_10566,N_11258);
xor U13341 (N_13341,N_11541,N_11764);
and U13342 (N_13342,N_11772,N_10804);
or U13343 (N_13343,N_11218,N_11748);
xor U13344 (N_13344,N_10568,N_10941);
or U13345 (N_13345,N_10506,N_10750);
or U13346 (N_13346,N_10816,N_11858);
and U13347 (N_13347,N_11904,N_11622);
and U13348 (N_13348,N_10900,N_11922);
and U13349 (N_13349,N_11898,N_11764);
or U13350 (N_13350,N_11119,N_11064);
nand U13351 (N_13351,N_10996,N_11068);
nand U13352 (N_13352,N_11885,N_11177);
nand U13353 (N_13353,N_10755,N_10523);
nand U13354 (N_13354,N_10922,N_10530);
nand U13355 (N_13355,N_11537,N_11391);
or U13356 (N_13356,N_10704,N_11499);
nand U13357 (N_13357,N_10794,N_11512);
xnor U13358 (N_13358,N_10570,N_11142);
and U13359 (N_13359,N_11916,N_10815);
nor U13360 (N_13360,N_11031,N_11066);
nand U13361 (N_13361,N_11873,N_11186);
nand U13362 (N_13362,N_11774,N_10961);
nor U13363 (N_13363,N_11953,N_11294);
or U13364 (N_13364,N_11437,N_11924);
nand U13365 (N_13365,N_10902,N_11367);
and U13366 (N_13366,N_11411,N_11755);
xnor U13367 (N_13367,N_11858,N_11486);
and U13368 (N_13368,N_11825,N_11126);
nand U13369 (N_13369,N_11768,N_10594);
nand U13370 (N_13370,N_11470,N_11450);
nor U13371 (N_13371,N_11365,N_10831);
or U13372 (N_13372,N_11321,N_11780);
or U13373 (N_13373,N_10535,N_11132);
nand U13374 (N_13374,N_10990,N_11389);
and U13375 (N_13375,N_11048,N_10857);
xor U13376 (N_13376,N_11131,N_10852);
and U13377 (N_13377,N_11625,N_10682);
nor U13378 (N_13378,N_11090,N_10639);
xnor U13379 (N_13379,N_11708,N_11486);
or U13380 (N_13380,N_11089,N_11571);
nor U13381 (N_13381,N_11622,N_10784);
nor U13382 (N_13382,N_11166,N_10911);
and U13383 (N_13383,N_10677,N_11937);
xnor U13384 (N_13384,N_11327,N_11139);
and U13385 (N_13385,N_10856,N_11431);
nand U13386 (N_13386,N_11145,N_11042);
or U13387 (N_13387,N_11537,N_11433);
or U13388 (N_13388,N_11114,N_10530);
or U13389 (N_13389,N_10928,N_11539);
xnor U13390 (N_13390,N_11789,N_11716);
nand U13391 (N_13391,N_11853,N_10571);
or U13392 (N_13392,N_11112,N_11958);
xor U13393 (N_13393,N_10672,N_11697);
and U13394 (N_13394,N_10677,N_11684);
or U13395 (N_13395,N_10772,N_10918);
nor U13396 (N_13396,N_10878,N_10955);
and U13397 (N_13397,N_11151,N_10744);
and U13398 (N_13398,N_11137,N_10970);
nor U13399 (N_13399,N_11123,N_11507);
and U13400 (N_13400,N_11094,N_10684);
and U13401 (N_13401,N_10986,N_11035);
xnor U13402 (N_13402,N_11948,N_11572);
nand U13403 (N_13403,N_11476,N_11108);
and U13404 (N_13404,N_11772,N_11396);
and U13405 (N_13405,N_11413,N_11457);
nor U13406 (N_13406,N_11138,N_11715);
nor U13407 (N_13407,N_11406,N_10760);
nand U13408 (N_13408,N_11359,N_11128);
or U13409 (N_13409,N_10848,N_11842);
and U13410 (N_13410,N_11035,N_11508);
nor U13411 (N_13411,N_11296,N_11824);
or U13412 (N_13412,N_11991,N_11808);
or U13413 (N_13413,N_10943,N_11231);
or U13414 (N_13414,N_10901,N_11945);
nand U13415 (N_13415,N_11742,N_11554);
nor U13416 (N_13416,N_11351,N_11459);
nor U13417 (N_13417,N_11714,N_10640);
nor U13418 (N_13418,N_11940,N_10808);
nand U13419 (N_13419,N_10629,N_11650);
and U13420 (N_13420,N_10898,N_11672);
nor U13421 (N_13421,N_11196,N_10884);
nor U13422 (N_13422,N_10628,N_11770);
and U13423 (N_13423,N_11429,N_11178);
or U13424 (N_13424,N_10618,N_10844);
and U13425 (N_13425,N_10710,N_10754);
or U13426 (N_13426,N_10522,N_11294);
xor U13427 (N_13427,N_11543,N_10682);
nor U13428 (N_13428,N_10894,N_11862);
nand U13429 (N_13429,N_11214,N_11648);
and U13430 (N_13430,N_11321,N_11493);
nand U13431 (N_13431,N_11734,N_10747);
nand U13432 (N_13432,N_11572,N_11674);
and U13433 (N_13433,N_11231,N_11296);
nor U13434 (N_13434,N_10745,N_11881);
or U13435 (N_13435,N_11495,N_11223);
and U13436 (N_13436,N_11295,N_11494);
and U13437 (N_13437,N_11190,N_11460);
or U13438 (N_13438,N_10750,N_11636);
nand U13439 (N_13439,N_10580,N_10859);
nand U13440 (N_13440,N_11912,N_11946);
nand U13441 (N_13441,N_10772,N_11865);
or U13442 (N_13442,N_11611,N_11056);
and U13443 (N_13443,N_11847,N_10861);
nand U13444 (N_13444,N_10945,N_10506);
nor U13445 (N_13445,N_11264,N_10772);
or U13446 (N_13446,N_11971,N_10741);
nand U13447 (N_13447,N_11903,N_11080);
and U13448 (N_13448,N_10726,N_11798);
nand U13449 (N_13449,N_11497,N_11267);
or U13450 (N_13450,N_11771,N_11644);
or U13451 (N_13451,N_11132,N_11475);
nor U13452 (N_13452,N_11076,N_10769);
and U13453 (N_13453,N_11262,N_11652);
nand U13454 (N_13454,N_11648,N_11231);
and U13455 (N_13455,N_10672,N_10506);
or U13456 (N_13456,N_11414,N_10799);
or U13457 (N_13457,N_10659,N_11896);
nor U13458 (N_13458,N_11135,N_11770);
nor U13459 (N_13459,N_11787,N_11334);
nand U13460 (N_13460,N_10524,N_11293);
or U13461 (N_13461,N_11151,N_10963);
nor U13462 (N_13462,N_10605,N_11700);
and U13463 (N_13463,N_11204,N_11887);
and U13464 (N_13464,N_11974,N_11563);
nand U13465 (N_13465,N_11194,N_11496);
or U13466 (N_13466,N_10826,N_11561);
xnor U13467 (N_13467,N_10835,N_11497);
and U13468 (N_13468,N_11402,N_11179);
xnor U13469 (N_13469,N_11299,N_11302);
and U13470 (N_13470,N_11883,N_10521);
nand U13471 (N_13471,N_10676,N_11412);
and U13472 (N_13472,N_10638,N_11262);
nand U13473 (N_13473,N_10674,N_11112);
or U13474 (N_13474,N_11811,N_11407);
and U13475 (N_13475,N_10836,N_10657);
nor U13476 (N_13476,N_11935,N_10542);
nand U13477 (N_13477,N_11920,N_11775);
nor U13478 (N_13478,N_11510,N_11516);
or U13479 (N_13479,N_11578,N_10530);
or U13480 (N_13480,N_11219,N_11488);
nand U13481 (N_13481,N_10850,N_10621);
and U13482 (N_13482,N_10566,N_11146);
xnor U13483 (N_13483,N_10513,N_11207);
and U13484 (N_13484,N_11711,N_10873);
nor U13485 (N_13485,N_10891,N_10899);
and U13486 (N_13486,N_10893,N_11980);
nor U13487 (N_13487,N_10600,N_11433);
nor U13488 (N_13488,N_11649,N_11859);
nor U13489 (N_13489,N_11285,N_11998);
nor U13490 (N_13490,N_11861,N_10961);
and U13491 (N_13491,N_10706,N_11402);
nand U13492 (N_13492,N_10774,N_11045);
or U13493 (N_13493,N_11940,N_11648);
nor U13494 (N_13494,N_11705,N_11372);
or U13495 (N_13495,N_10815,N_11660);
nand U13496 (N_13496,N_10641,N_11436);
and U13497 (N_13497,N_10949,N_11085);
and U13498 (N_13498,N_11680,N_11560);
or U13499 (N_13499,N_11760,N_11074);
nor U13500 (N_13500,N_12975,N_12877);
or U13501 (N_13501,N_12440,N_12239);
or U13502 (N_13502,N_12065,N_12368);
nand U13503 (N_13503,N_13034,N_13336);
or U13504 (N_13504,N_13369,N_13470);
nand U13505 (N_13505,N_12100,N_13376);
and U13506 (N_13506,N_12494,N_13154);
nand U13507 (N_13507,N_12316,N_12081);
nor U13508 (N_13508,N_12578,N_12804);
and U13509 (N_13509,N_12745,N_12497);
nor U13510 (N_13510,N_12073,N_13035);
nor U13511 (N_13511,N_12312,N_12269);
and U13512 (N_13512,N_12459,N_13070);
nand U13513 (N_13513,N_13079,N_12600);
nand U13514 (N_13514,N_12551,N_12977);
nor U13515 (N_13515,N_12860,N_13298);
or U13516 (N_13516,N_12930,N_12714);
nand U13517 (N_13517,N_12950,N_12138);
nor U13518 (N_13518,N_13314,N_12470);
nand U13519 (N_13519,N_12691,N_12643);
and U13520 (N_13520,N_12722,N_12153);
nor U13521 (N_13521,N_12985,N_12094);
or U13522 (N_13522,N_13057,N_12658);
or U13523 (N_13523,N_13234,N_12781);
or U13524 (N_13524,N_12416,N_13211);
nor U13525 (N_13525,N_12549,N_12192);
nand U13526 (N_13526,N_12803,N_12102);
and U13527 (N_13527,N_13197,N_12926);
nor U13528 (N_13528,N_13022,N_12448);
nand U13529 (N_13529,N_12514,N_12965);
and U13530 (N_13530,N_12132,N_12788);
nand U13531 (N_13531,N_12822,N_13220);
nor U13532 (N_13532,N_13489,N_12488);
or U13533 (N_13533,N_12289,N_12990);
nor U13534 (N_13534,N_12762,N_12379);
and U13535 (N_13535,N_13253,N_12608);
and U13536 (N_13536,N_12642,N_13186);
xor U13537 (N_13537,N_12335,N_13128);
nor U13538 (N_13538,N_13026,N_12139);
nor U13539 (N_13539,N_12789,N_12082);
nor U13540 (N_13540,N_13260,N_12896);
and U13541 (N_13541,N_12807,N_12413);
nand U13542 (N_13542,N_12430,N_12765);
xor U13543 (N_13543,N_12566,N_12571);
nand U13544 (N_13544,N_12393,N_12227);
and U13545 (N_13545,N_13257,N_13464);
nand U13546 (N_13546,N_12253,N_13042);
or U13547 (N_13547,N_12882,N_12339);
and U13548 (N_13548,N_12115,N_12236);
nor U13549 (N_13549,N_12110,N_13181);
xnor U13550 (N_13550,N_12195,N_12796);
nor U13551 (N_13551,N_12888,N_12778);
and U13552 (N_13552,N_12212,N_12517);
nand U13553 (N_13553,N_12061,N_13475);
nand U13554 (N_13554,N_12500,N_12121);
nand U13555 (N_13555,N_13131,N_12189);
and U13556 (N_13556,N_12521,N_12180);
and U13557 (N_13557,N_13157,N_12895);
xor U13558 (N_13558,N_12006,N_12108);
or U13559 (N_13559,N_12098,N_13010);
nand U13560 (N_13560,N_13061,N_13139);
nor U13561 (N_13561,N_12943,N_12937);
and U13562 (N_13562,N_13067,N_12009);
or U13563 (N_13563,N_12951,N_12650);
and U13564 (N_13564,N_12162,N_12668);
nor U13565 (N_13565,N_12136,N_13142);
nand U13566 (N_13566,N_13280,N_12432);
nand U13567 (N_13567,N_12063,N_13043);
nand U13568 (N_13568,N_13469,N_12728);
nand U13569 (N_13569,N_12609,N_13435);
xor U13570 (N_13570,N_12768,N_12688);
nor U13571 (N_13571,N_12878,N_13462);
nor U13572 (N_13572,N_12099,N_13102);
or U13573 (N_13573,N_12387,N_13359);
nor U13574 (N_13574,N_13400,N_12334);
nand U13575 (N_13575,N_12629,N_12516);
xnor U13576 (N_13576,N_12855,N_12466);
and U13577 (N_13577,N_12265,N_13208);
nand U13578 (N_13578,N_12451,N_12423);
nor U13579 (N_13579,N_13416,N_12016);
nor U13580 (N_13580,N_12284,N_12815);
nor U13581 (N_13581,N_13311,N_12279);
or U13582 (N_13582,N_12574,N_12361);
or U13583 (N_13583,N_12767,N_12161);
nor U13584 (N_13584,N_13459,N_12321);
and U13585 (N_13585,N_13434,N_12071);
xor U13586 (N_13586,N_12601,N_12859);
nor U13587 (N_13587,N_13461,N_12823);
or U13588 (N_13588,N_12047,N_12193);
xor U13589 (N_13589,N_12570,N_12058);
and U13590 (N_13590,N_12587,N_13009);
nor U13591 (N_13591,N_12041,N_13219);
nand U13592 (N_13592,N_12680,N_12721);
and U13593 (N_13593,N_13347,N_13013);
or U13594 (N_13594,N_13136,N_12408);
or U13595 (N_13595,N_12087,N_12606);
or U13596 (N_13596,N_13091,N_13365);
and U13597 (N_13597,N_12511,N_13448);
or U13598 (N_13598,N_13151,N_12455);
or U13599 (N_13599,N_12305,N_12458);
nand U13600 (N_13600,N_12229,N_13072);
and U13601 (N_13601,N_13383,N_12175);
nor U13602 (N_13602,N_12824,N_13171);
xor U13603 (N_13603,N_12582,N_13198);
nand U13604 (N_13604,N_13317,N_12141);
or U13605 (N_13605,N_12693,N_12004);
nand U13606 (N_13606,N_12702,N_12909);
and U13607 (N_13607,N_12766,N_13279);
nand U13608 (N_13608,N_12954,N_13486);
and U13609 (N_13609,N_12320,N_12191);
nand U13610 (N_13610,N_12939,N_13269);
xnor U13611 (N_13611,N_13245,N_12631);
xnor U13612 (N_13612,N_12422,N_12522);
and U13613 (N_13613,N_12851,N_13120);
xnor U13614 (N_13614,N_13003,N_12346);
or U13615 (N_13615,N_12375,N_12306);
or U13616 (N_13616,N_13203,N_12929);
and U13617 (N_13617,N_12506,N_12317);
or U13618 (N_13618,N_12233,N_12275);
or U13619 (N_13619,N_13381,N_12736);
nor U13620 (N_13620,N_12509,N_12394);
nor U13621 (N_13621,N_12001,N_12104);
nand U13622 (N_13622,N_12769,N_12215);
or U13623 (N_13623,N_12901,N_13059);
nand U13624 (N_13624,N_12599,N_12739);
or U13625 (N_13625,N_12067,N_13296);
nand U13626 (N_13626,N_12559,N_12185);
nor U13627 (N_13627,N_12134,N_12278);
nand U13628 (N_13628,N_13485,N_12101);
and U13629 (N_13629,N_13146,N_12245);
or U13630 (N_13630,N_13321,N_13007);
nand U13631 (N_13631,N_12864,N_12124);
or U13632 (N_13632,N_12266,N_12217);
nor U13633 (N_13633,N_13421,N_12113);
or U13634 (N_13634,N_13152,N_12301);
nand U13635 (N_13635,N_13454,N_12190);
nor U13636 (N_13636,N_13479,N_12122);
or U13637 (N_13637,N_12567,N_12740);
and U13638 (N_13638,N_12095,N_13164);
nand U13639 (N_13639,N_12446,N_12857);
or U13640 (N_13640,N_12698,N_12628);
nand U13641 (N_13641,N_12294,N_12114);
or U13642 (N_13642,N_12130,N_13018);
nand U13643 (N_13643,N_12790,N_12120);
xor U13644 (N_13644,N_12591,N_12097);
or U13645 (N_13645,N_12223,N_13342);
nor U13646 (N_13646,N_12077,N_12750);
nor U13647 (N_13647,N_12250,N_13425);
or U13648 (N_13648,N_12228,N_13271);
nor U13649 (N_13649,N_12845,N_13442);
xnor U13650 (N_13650,N_12727,N_13327);
nand U13651 (N_13651,N_12593,N_12127);
and U13652 (N_13652,N_13101,N_13352);
nor U13653 (N_13653,N_12482,N_12263);
xnor U13654 (N_13654,N_12002,N_12350);
nand U13655 (N_13655,N_12978,N_13041);
and U13656 (N_13656,N_12048,N_12830);
xor U13657 (N_13657,N_13446,N_13318);
nand U13658 (N_13658,N_12219,N_12993);
and U13659 (N_13659,N_12816,N_13218);
nor U13660 (N_13660,N_12562,N_13239);
nand U13661 (N_13661,N_12307,N_13325);
or U13662 (N_13662,N_12103,N_13028);
xor U13663 (N_13663,N_13354,N_12270);
nor U13664 (N_13664,N_12079,N_12424);
xor U13665 (N_13665,N_13224,N_12057);
nand U13666 (N_13666,N_12826,N_12086);
or U13667 (N_13667,N_13375,N_12697);
or U13668 (N_13668,N_13230,N_12818);
and U13669 (N_13669,N_12873,N_13021);
and U13670 (N_13670,N_12771,N_12717);
and U13671 (N_13671,N_13020,N_12806);
nand U13672 (N_13672,N_13398,N_12831);
nand U13673 (N_13673,N_13005,N_13427);
nor U13674 (N_13674,N_13135,N_12282);
nand U13675 (N_13675,N_13452,N_12281);
nand U13676 (N_13676,N_13115,N_12479);
xor U13677 (N_13677,N_12991,N_12385);
nor U13678 (N_13678,N_12274,N_13247);
and U13679 (N_13679,N_12014,N_12142);
and U13680 (N_13680,N_12983,N_12208);
or U13681 (N_13681,N_13210,N_12676);
nand U13682 (N_13682,N_12123,N_12012);
and U13683 (N_13683,N_12777,N_12633);
nor U13684 (N_13684,N_13248,N_13453);
or U13685 (N_13685,N_13012,N_13086);
nor U13686 (N_13686,N_12331,N_13491);
nor U13687 (N_13687,N_13190,N_12996);
and U13688 (N_13688,N_12062,N_13049);
nor U13689 (N_13689,N_12475,N_12976);
or U13690 (N_13690,N_12992,N_13439);
nor U13691 (N_13691,N_12434,N_13265);
nor U13692 (N_13692,N_12537,N_12671);
xor U13693 (N_13693,N_13412,N_12283);
or U13694 (N_13694,N_13155,N_13037);
nor U13695 (N_13695,N_13490,N_12345);
and U13696 (N_13696,N_12246,N_12241);
nor U13697 (N_13697,N_12735,N_12119);
or U13698 (N_13698,N_12295,N_13196);
nand U13699 (N_13699,N_12495,N_12893);
and U13700 (N_13700,N_12442,N_12947);
or U13701 (N_13701,N_13444,N_13285);
nand U13702 (N_13702,N_12302,N_12042);
nor U13703 (N_13703,N_12743,N_12902);
nor U13704 (N_13704,N_13338,N_13329);
nor U13705 (N_13705,N_12799,N_12318);
nor U13706 (N_13706,N_13129,N_12213);
xor U13707 (N_13707,N_13306,N_12916);
xor U13708 (N_13708,N_12045,N_12453);
xnor U13709 (N_13709,N_13322,N_13056);
or U13710 (N_13710,N_12027,N_12971);
and U13711 (N_13711,N_13463,N_13428);
or U13712 (N_13712,N_12021,N_13258);
nor U13713 (N_13713,N_12936,N_13137);
or U13714 (N_13714,N_12010,N_13451);
or U13715 (N_13715,N_12372,N_13179);
nand U13716 (N_13716,N_13166,N_13341);
or U13717 (N_13717,N_12701,N_13346);
or U13718 (N_13718,N_13015,N_12832);
and U13719 (N_13719,N_12469,N_12209);
or U13720 (N_13720,N_12699,N_12946);
nand U13721 (N_13721,N_12614,N_12627);
nand U13722 (N_13722,N_12106,N_12805);
nand U13723 (N_13723,N_13033,N_13046);
nand U13724 (N_13724,N_12460,N_12272);
nand U13725 (N_13725,N_13403,N_13351);
or U13726 (N_13726,N_12310,N_12157);
nor U13727 (N_13727,N_13356,N_13368);
nor U13728 (N_13728,N_13432,N_13268);
or U13729 (N_13729,N_13417,N_12558);
and U13730 (N_13730,N_13187,N_12362);
nand U13731 (N_13731,N_12773,N_13293);
nand U13732 (N_13732,N_12922,N_12313);
or U13733 (N_13733,N_12941,N_12017);
and U13734 (N_13734,N_13273,N_12649);
nor U13735 (N_13735,N_13192,N_12586);
and U13736 (N_13736,N_13278,N_12222);
nor U13737 (N_13737,N_13367,N_13097);
or U13738 (N_13738,N_13156,N_12216);
nor U13739 (N_13739,N_13191,N_12812);
nand U13740 (N_13740,N_12581,N_12644);
nand U13741 (N_13741,N_13076,N_12373);
or U13742 (N_13742,N_12553,N_12746);
xnor U13743 (N_13743,N_12020,N_12724);
xnor U13744 (N_13744,N_12165,N_13083);
nand U13745 (N_13745,N_12204,N_12188);
nor U13746 (N_13746,N_12205,N_12224);
or U13747 (N_13747,N_12352,N_12530);
nor U13748 (N_13748,N_12641,N_12182);
nor U13749 (N_13749,N_12401,N_13431);
or U13750 (N_13750,N_13404,N_12967);
or U13751 (N_13751,N_13121,N_13343);
xnor U13752 (N_13752,N_12304,N_12705);
nand U13753 (N_13753,N_13094,N_13290);
xnor U13754 (N_13754,N_12592,N_13419);
nand U13755 (N_13755,N_12211,N_13002);
xor U13756 (N_13756,N_12894,N_12527);
nor U13757 (N_13757,N_12436,N_12982);
xnor U13758 (N_13758,N_12764,N_12054);
xor U13759 (N_13759,N_12092,N_12617);
nor U13760 (N_13760,N_12580,N_12646);
nor U13761 (N_13761,N_13313,N_12748);
nor U13762 (N_13762,N_12150,N_12912);
or U13763 (N_13763,N_13207,N_13466);
nand U13764 (N_13764,N_12149,N_12927);
xnor U13765 (N_13765,N_13051,N_12007);
xnor U13766 (N_13766,N_12602,N_12866);
nor U13767 (N_13767,N_12344,N_13487);
or U13768 (N_13768,N_13199,N_12478);
or U13769 (N_13769,N_13103,N_13402);
nor U13770 (N_13770,N_13324,N_12839);
nor U13771 (N_13771,N_13286,N_12809);
nor U13772 (N_13772,N_13482,N_12682);
nand U13773 (N_13773,N_12452,N_13232);
or U13774 (N_13774,N_13358,N_12322);
nand U13775 (N_13775,N_12653,N_13241);
and U13776 (N_13776,N_12164,N_12028);
and U13777 (N_13777,N_13240,N_12329);
nand U13778 (N_13778,N_13377,N_12226);
nor U13779 (N_13779,N_12908,N_12258);
and U13780 (N_13780,N_12986,N_13011);
and U13781 (N_13781,N_12520,N_12330);
nor U13782 (N_13782,N_12174,N_13393);
and U13783 (N_13783,N_12443,N_12022);
nor U13784 (N_13784,N_12607,N_13141);
and U13785 (N_13785,N_12252,N_13193);
or U13786 (N_13786,N_13478,N_12785);
or U13787 (N_13787,N_12238,N_12187);
or U13788 (N_13788,N_12536,N_12064);
nand U13789 (N_13789,N_13263,N_12315);
xnor U13790 (N_13790,N_13252,N_12111);
or U13791 (N_13791,N_12474,N_13214);
nand U13792 (N_13792,N_12358,N_12849);
nand U13793 (N_13793,N_12515,N_13483);
or U13794 (N_13794,N_12431,N_12367);
or U13795 (N_13795,N_12388,N_13226);
nand U13796 (N_13796,N_12585,N_13242);
nor U13797 (N_13797,N_12131,N_12490);
and U13798 (N_13798,N_12678,N_13017);
and U13799 (N_13799,N_12679,N_13223);
and U13800 (N_13800,N_12412,N_12417);
nor U13801 (N_13801,N_13050,N_12988);
xnor U13802 (N_13802,N_13205,N_13274);
nor U13803 (N_13803,N_13387,N_12659);
xnor U13804 (N_13804,N_12341,N_13426);
or U13805 (N_13805,N_12462,N_13294);
and U13806 (N_13806,N_13143,N_13016);
nand U13807 (N_13807,N_12090,N_12404);
or U13808 (N_13808,N_12645,N_12899);
xor U13809 (N_13809,N_12052,N_12801);
nand U13810 (N_13810,N_12683,N_13158);
nand U13811 (N_13811,N_12183,N_13437);
nor U13812 (N_13812,N_12512,N_12959);
nand U13813 (N_13813,N_12084,N_12342);
or U13814 (N_13814,N_13185,N_12963);
nand U13815 (N_13815,N_12874,N_12261);
or U13816 (N_13816,N_13385,N_12293);
and U13817 (N_13817,N_13071,N_13414);
nor U13818 (N_13818,N_12561,N_12221);
or U13819 (N_13819,N_12349,N_13484);
xnor U13820 (N_13820,N_12618,N_12210);
nor U13821 (N_13821,N_12962,N_12421);
nand U13822 (N_13822,N_12692,N_12793);
nor U13823 (N_13823,N_13264,N_12015);
or U13824 (N_13824,N_12030,N_12883);
nand U13825 (N_13825,N_12786,N_13477);
and U13826 (N_13826,N_13132,N_12526);
nor U13827 (N_13827,N_13073,N_13040);
or U13828 (N_13828,N_12240,N_13433);
nor U13829 (N_13829,N_12172,N_12176);
or U13830 (N_13830,N_13345,N_12532);
nand U13831 (N_13831,N_13254,N_12383);
nor U13832 (N_13832,N_12376,N_13436);
and U13833 (N_13833,N_13405,N_12670);
xnor U13834 (N_13834,N_13024,N_12489);
nor U13835 (N_13835,N_12657,N_12661);
nand U13836 (N_13836,N_12264,N_13093);
or U13837 (N_13837,N_12429,N_13379);
nand U13838 (N_13838,N_13289,N_12998);
or U13839 (N_13839,N_13008,N_13225);
nand U13840 (N_13840,N_12619,N_12378);
nand U13841 (N_13841,N_13114,N_12151);
and U13842 (N_13842,N_12972,N_13291);
nor U13843 (N_13843,N_13149,N_13335);
and U13844 (N_13844,N_13323,N_12598);
nor U13845 (N_13845,N_13334,N_12069);
nor U13846 (N_13846,N_13305,N_13267);
nand U13847 (N_13847,N_13209,N_12800);
and U13848 (N_13848,N_13288,N_12960);
xor U13849 (N_13849,N_12397,N_12589);
nor U13850 (N_13850,N_12477,N_12779);
and U13851 (N_13851,N_13100,N_12400);
and U13852 (N_13852,N_12763,N_12813);
nand U13853 (N_13853,N_12795,N_12684);
or U13854 (N_13854,N_12686,N_12439);
nand U13855 (N_13855,N_12406,N_12535);
or U13856 (N_13856,N_13457,N_12848);
xor U13857 (N_13857,N_12953,N_13045);
or U13858 (N_13858,N_12476,N_12999);
nor U13859 (N_13859,N_12243,N_13066);
or U13860 (N_13860,N_12863,N_13182);
xnor U13861 (N_13861,N_13283,N_13370);
nor U13862 (N_13862,N_13231,N_12552);
or U13863 (N_13863,N_12725,N_12053);
nor U13864 (N_13864,N_12481,N_12924);
xor U13865 (N_13865,N_12970,N_12635);
or U13866 (N_13866,N_12140,N_12220);
and U13867 (N_13867,N_12194,N_12524);
nor U13868 (N_13868,N_12887,N_12575);
nor U13869 (N_13869,N_12938,N_13389);
nand U13870 (N_13870,N_13212,N_13455);
or U13871 (N_13871,N_12889,N_12817);
or U13872 (N_13872,N_12355,N_12298);
nor U13873 (N_13873,N_12457,N_13409);
nand U13874 (N_13874,N_13481,N_12271);
nand U13875 (N_13875,N_12569,N_12198);
xor U13876 (N_13876,N_12303,N_13201);
nand U13877 (N_13877,N_13301,N_13440);
and U13878 (N_13878,N_13235,N_12925);
nand U13879 (N_13879,N_12904,N_12242);
nor U13880 (N_13880,N_13233,N_12531);
nand U13881 (N_13881,N_13054,N_13077);
and U13882 (N_13882,N_13118,N_12128);
xnor U13883 (N_13883,N_12518,N_12399);
nand U13884 (N_13884,N_12276,N_12471);
xnor U13885 (N_13885,N_12610,N_13087);
or U13886 (N_13886,N_12107,N_12534);
nor U13887 (N_13887,N_12038,N_12332);
or U13888 (N_13888,N_12170,N_13133);
or U13889 (N_13889,N_12995,N_12326);
nand U13890 (N_13890,N_12665,N_13423);
or U13891 (N_13891,N_12019,N_13213);
nor U13892 (N_13892,N_12961,N_13058);
or U13893 (N_13893,N_12923,N_12834);
nor U13894 (N_13894,N_12354,N_12538);
nor U13895 (N_13895,N_13062,N_12003);
nor U13896 (N_13896,N_12179,N_12666);
nor U13897 (N_13897,N_12050,N_12616);
nor U13898 (N_13898,N_12576,N_12821);
or U13899 (N_13899,N_12928,N_13309);
nand U13900 (N_13900,N_12523,N_12776);
nor U13901 (N_13901,N_12415,N_13328);
and U13902 (N_13902,N_12268,N_12677);
xnor U13903 (N_13903,N_12200,N_13460);
or U13904 (N_13904,N_12232,N_13188);
nand U13905 (N_13905,N_12742,N_13119);
nand U13906 (N_13906,N_13237,N_13085);
xor U13907 (N_13907,N_12381,N_12337);
nor U13908 (N_13908,N_13032,N_12262);
and U13909 (N_13909,N_12324,N_12528);
nor U13910 (N_13910,N_12835,N_13173);
nor U13911 (N_13911,N_12426,N_12148);
xnor U13912 (N_13912,N_13438,N_12749);
nor U13913 (N_13913,N_13052,N_13030);
or U13914 (N_13914,N_12914,N_13262);
nand U13915 (N_13915,N_12997,N_13410);
nor U13916 (N_13916,N_13472,N_12024);
nor U13917 (N_13917,N_13430,N_13467);
nor U13918 (N_13918,N_13172,N_12969);
or U13919 (N_13919,N_13238,N_12109);
nand U13920 (N_13920,N_12563,N_12147);
xor U13921 (N_13921,N_13471,N_12135);
xor U13922 (N_13922,N_12491,N_12709);
nor U13923 (N_13923,N_13331,N_12611);
nor U13924 (N_13924,N_13281,N_12498);
and U13925 (N_13925,N_12984,N_12726);
or U13926 (N_13926,N_13123,N_12395);
nand U13927 (N_13927,N_13168,N_12386);
xnor U13928 (N_13928,N_12720,N_13382);
and U13929 (N_13929,N_12186,N_12309);
and U13930 (N_13930,N_12449,N_12780);
and U13931 (N_13931,N_12144,N_12761);
xor U13932 (N_13932,N_12733,N_13029);
and U13933 (N_13933,N_12105,N_12025);
nand U13934 (N_13934,N_12484,N_12695);
nor U13935 (N_13935,N_12181,N_13222);
nor U13936 (N_13936,N_13019,N_12163);
or U13937 (N_13937,N_12710,N_12841);
or U13938 (N_13938,N_13063,N_12689);
nand U13939 (N_13939,N_13303,N_13177);
or U13940 (N_13940,N_12409,N_12507);
and U13941 (N_13941,N_12467,N_13497);
nand U13942 (N_13942,N_13195,N_12166);
nor U13943 (N_13943,N_12903,N_12093);
and U13944 (N_13944,N_13330,N_12129);
xnor U13945 (N_13945,N_13027,N_12356);
and U13946 (N_13946,N_13127,N_13320);
and U13947 (N_13947,N_13420,N_13380);
or U13948 (N_13948,N_12370,N_13122);
nor U13949 (N_13949,N_12405,N_13411);
and U13950 (N_13950,N_12913,N_13364);
or U13951 (N_13951,N_12359,N_13344);
xnor U13952 (N_13952,N_12729,N_13130);
nand U13953 (N_13953,N_13109,N_12177);
nor U13954 (N_13954,N_13144,N_12184);
nand U13955 (N_13955,N_12758,N_13308);
or U13956 (N_13956,N_13349,N_13270);
and U13957 (N_13957,N_12875,N_13493);
nand U13958 (N_13958,N_13332,N_12112);
nor U13959 (N_13959,N_12353,N_12700);
nor U13960 (N_13960,N_13084,N_12772);
nand U13961 (N_13961,N_13025,N_13355);
and U13962 (N_13962,N_13038,N_12744);
nor U13963 (N_13963,N_13340,N_12504);
nand U13964 (N_13964,N_12447,N_12502);
or U13965 (N_13965,N_13147,N_12753);
nor U13966 (N_13966,N_12133,N_13422);
and U13967 (N_13967,N_12323,N_12032);
nand U13968 (N_13968,N_13401,N_12008);
or U13969 (N_13969,N_12595,N_13069);
or U13970 (N_13970,N_12340,N_12300);
xnor U13971 (N_13971,N_12389,N_12357);
nor U13972 (N_13972,N_12572,N_12622);
nand U13973 (N_13973,N_12034,N_12811);
or U13974 (N_13974,N_12051,N_12059);
nand U13975 (N_13975,N_12256,N_12251);
and U13976 (N_13976,N_13112,N_13339);
nor U13977 (N_13977,N_12940,N_12225);
or U13978 (N_13978,N_13249,N_12203);
nor U13979 (N_13979,N_13441,N_12952);
nand U13980 (N_13980,N_12445,N_12377);
or U13981 (N_13981,N_12669,N_12468);
nor U13982 (N_13982,N_12525,N_13081);
and U13983 (N_13983,N_12510,N_13361);
nor U13984 (N_13984,N_12751,N_12934);
nor U13985 (N_13985,N_13053,N_13246);
nand U13986 (N_13986,N_12487,N_12070);
or U13987 (N_13987,N_12870,N_12199);
nand U13988 (N_13988,N_13215,N_12410);
nor U13989 (N_13989,N_12613,N_12674);
nor U13990 (N_13990,N_12651,N_13126);
or U13991 (N_13991,N_12694,N_12055);
nand U13992 (N_13992,N_13366,N_12931);
nor U13993 (N_13993,N_13170,N_12390);
nor U13994 (N_13994,N_12427,N_12391);
and U13995 (N_13995,N_12327,N_12757);
nand U13996 (N_13996,N_13396,N_12712);
nand U13997 (N_13997,N_12782,N_13036);
xnor U13998 (N_13998,N_13499,N_13039);
or U13999 (N_13999,N_12624,N_12308);
or U14000 (N_14000,N_12013,N_13064);
and U14001 (N_14001,N_12197,N_12955);
xnor U14002 (N_14002,N_12949,N_12837);
nand U14003 (N_14003,N_13319,N_12503);
nand U14004 (N_14004,N_13371,N_12783);
nor U14005 (N_14005,N_13384,N_12921);
xnor U14006 (N_14006,N_13250,N_12438);
nand U14007 (N_14007,N_12011,N_12656);
and U14008 (N_14008,N_12060,N_12068);
nand U14009 (N_14009,N_13299,N_12704);
and U14010 (N_14010,N_12456,N_12542);
and U14011 (N_14011,N_13312,N_12933);
nor U14012 (N_14012,N_12632,N_12096);
nand U14013 (N_14013,N_12548,N_12787);
nand U14014 (N_14014,N_13266,N_13413);
or U14015 (N_14015,N_12496,N_13078);
nand U14016 (N_14016,N_12555,N_13044);
or U14017 (N_14017,N_12218,N_13204);
and U14018 (N_14018,N_12273,N_12259);
nor U14019 (N_14019,N_12156,N_12437);
and U14020 (N_14020,N_13326,N_12620);
and U14021 (N_14021,N_12850,N_12557);
and U14022 (N_14022,N_12043,N_12248);
xor U14023 (N_14023,N_12827,N_12348);
and U14024 (N_14024,N_12685,N_12672);
and U14025 (N_14025,N_12637,N_12247);
or U14026 (N_14026,N_12828,N_12360);
nor U14027 (N_14027,N_13194,N_12037);
nor U14028 (N_14028,N_12754,N_13178);
or U14029 (N_14029,N_12973,N_13255);
and U14030 (N_14030,N_13113,N_12854);
and U14031 (N_14031,N_13159,N_12718);
nand U14032 (N_14032,N_13392,N_12169);
nand U14033 (N_14033,N_12056,N_12838);
nor U14034 (N_14034,N_12596,N_12152);
xnor U14035 (N_14035,N_12297,N_12154);
nand U14036 (N_14036,N_12737,N_13276);
nor U14037 (N_14037,N_12560,N_13161);
nand U14038 (N_14038,N_12505,N_12023);
nor U14039 (N_14039,N_13445,N_12989);
and U14040 (N_14040,N_13307,N_13099);
or U14041 (N_14041,N_12853,N_12756);
or U14042 (N_14042,N_12539,N_13406);
or U14043 (N_14043,N_12731,N_13105);
nor U14044 (N_14044,N_12286,N_12696);
or U14045 (N_14045,N_13167,N_12942);
xnor U14046 (N_14046,N_12820,N_12964);
nand U14047 (N_14047,N_12846,N_13150);
or U14048 (N_14048,N_12541,N_13337);
nand U14049 (N_14049,N_12747,N_12605);
and U14050 (N_14050,N_12640,N_12630);
nand U14051 (N_14051,N_13165,N_12664);
nand U14052 (N_14052,N_13399,N_13284);
nand U14053 (N_14053,N_12146,N_13145);
or U14054 (N_14054,N_13104,N_13111);
nand U14055 (N_14055,N_12621,N_12411);
or U14056 (N_14056,N_12291,N_13047);
nand U14057 (N_14057,N_12681,N_12842);
nand U14058 (N_14058,N_12615,N_13004);
nand U14059 (N_14059,N_12402,N_12483);
or U14060 (N_14060,N_12872,N_12196);
and U14061 (N_14061,N_12244,N_12380);
or U14062 (N_14062,N_12296,N_13390);
or U14063 (N_14063,N_12234,N_12026);
nand U14064 (N_14064,N_12255,N_12715);
and U14065 (N_14065,N_12647,N_12654);
nand U14066 (N_14066,N_12267,N_12480);
nor U14067 (N_14067,N_12074,N_12049);
and U14068 (N_14068,N_12636,N_12285);
nand U14069 (N_14069,N_13362,N_13304);
nand U14070 (N_14070,N_13180,N_13092);
or U14071 (N_14071,N_12472,N_12040);
xnor U14072 (N_14072,N_12871,N_13184);
nand U14073 (N_14073,N_13095,N_12492);
or U14074 (N_14074,N_12868,N_13060);
nand U14075 (N_14075,N_13474,N_12091);
or U14076 (N_14076,N_13229,N_12158);
xnor U14077 (N_14077,N_13080,N_13315);
nand U14078 (N_14078,N_12206,N_13125);
or U14079 (N_14079,N_13424,N_13216);
nor U14080 (N_14080,N_12867,N_12565);
xor U14081 (N_14081,N_12798,N_13031);
or U14082 (N_14082,N_13458,N_13175);
nor U14083 (N_14083,N_12987,N_12519);
nand U14084 (N_14084,N_12919,N_13162);
xnor U14085 (N_14085,N_13275,N_13251);
and U14086 (N_14086,N_12155,N_12738);
nand U14087 (N_14087,N_12588,N_12005);
and U14088 (N_14088,N_12966,N_12907);
and U14089 (N_14089,N_12957,N_13408);
nor U14090 (N_14090,N_12237,N_12825);
nor U14091 (N_14091,N_13106,N_13116);
nand U14092 (N_14092,N_12707,N_12336);
and U14093 (N_14093,N_12168,N_12556);
nand U14094 (N_14094,N_12703,N_12884);
and U14095 (N_14095,N_12968,N_12085);
nand U14096 (N_14096,N_12493,N_12072);
xnor U14097 (N_14097,N_12554,N_12829);
nand U14098 (N_14098,N_12711,N_12420);
nor U14099 (N_14099,N_12660,N_12910);
or U14100 (N_14100,N_12897,N_13480);
nand U14101 (N_14101,N_13244,N_12546);
or U14102 (N_14102,N_12891,N_12879);
nor U14103 (N_14103,N_12755,N_13282);
and U14104 (N_14104,N_12590,N_13140);
nor U14105 (N_14105,N_12869,N_13374);
nor U14106 (N_14106,N_12918,N_12143);
or U14107 (N_14107,N_12428,N_12364);
nand U14108 (N_14108,N_13297,N_12881);
and U14109 (N_14109,N_12719,N_12444);
nor U14110 (N_14110,N_12036,N_12862);
nand U14111 (N_14111,N_12403,N_12533);
xor U14112 (N_14112,N_13256,N_12171);
or U14113 (N_14113,N_12708,N_12915);
nand U14114 (N_14114,N_12260,N_12463);
nor U14115 (N_14115,N_12543,N_12441);
or U14116 (N_14116,N_12178,N_12464);
nand U14117 (N_14117,N_13449,N_12810);
and U14118 (N_14118,N_12145,N_12673);
nand U14119 (N_14119,N_12325,N_12235);
nor U14120 (N_14120,N_12775,N_13488);
and U14121 (N_14121,N_12652,N_13169);
nand U14122 (N_14122,N_12351,N_12944);
xor U14123 (N_14123,N_12277,N_12425);
nor U14124 (N_14124,N_13494,N_13498);
and U14125 (N_14125,N_12752,N_12407);
nor U14126 (N_14126,N_13407,N_13456);
nor U14127 (N_14127,N_12980,N_12540);
nand U14128 (N_14128,N_12382,N_12932);
or U14129 (N_14129,N_12981,N_12906);
and U14130 (N_14130,N_12465,N_12956);
nor U14131 (N_14131,N_12485,N_12876);
or U14132 (N_14132,N_12639,N_12343);
nor U14133 (N_14133,N_12435,N_12713);
and U14134 (N_14134,N_13014,N_12075);
nand U14135 (N_14135,N_13023,N_13394);
nand U14136 (N_14136,N_12892,N_13350);
and U14137 (N_14137,N_12230,N_13391);
xor U14138 (N_14138,N_12384,N_12935);
nor U14139 (N_14139,N_12573,N_12808);
and U14140 (N_14140,N_12254,N_12201);
and U14141 (N_14141,N_12662,N_12433);
nor U14142 (N_14142,N_13098,N_12486);
and U14143 (N_14143,N_12911,N_12945);
nand U14144 (N_14144,N_13006,N_12856);
nor U14145 (N_14145,N_12089,N_12333);
xnor U14146 (N_14146,N_13160,N_12890);
nor U14147 (N_14147,N_13117,N_12844);
nand U14148 (N_14148,N_12730,N_12774);
and U14149 (N_14149,N_12311,N_12508);
nand U14150 (N_14150,N_12039,N_12328);
and U14151 (N_14151,N_12833,N_12579);
and U14152 (N_14152,N_12723,N_13372);
or U14153 (N_14153,N_12499,N_13261);
nand U14154 (N_14154,N_13476,N_12675);
and U14155 (N_14155,N_12365,N_12794);
or U14156 (N_14156,N_12513,N_12638);
and U14157 (N_14157,N_12280,N_12257);
and U14158 (N_14158,N_12584,N_13418);
xor U14159 (N_14159,N_12398,N_12994);
nand U14160 (N_14160,N_13148,N_13206);
nor U14161 (N_14161,N_12690,N_13473);
and U14162 (N_14162,N_12116,N_12948);
or U14163 (N_14163,N_12414,N_12583);
nor U14164 (N_14164,N_13353,N_12080);
xor U14165 (N_14165,N_12160,N_13001);
xnor U14166 (N_14166,N_12861,N_12338);
or U14167 (N_14167,N_12917,N_12802);
nand U14168 (N_14168,N_12288,N_12419);
nor U14169 (N_14169,N_13348,N_12792);
nand U14170 (N_14170,N_12577,N_12031);
and U14171 (N_14171,N_12076,N_12687);
and U14172 (N_14172,N_13055,N_12231);
nor U14173 (N_14173,N_12655,N_12299);
and U14174 (N_14174,N_13090,N_12847);
xor U14175 (N_14175,N_12648,N_12920);
or U14176 (N_14176,N_13316,N_13447);
nand U14177 (N_14177,N_12568,N_13496);
and U14178 (N_14178,N_12900,N_12369);
xnor U14179 (N_14179,N_13221,N_12126);
xor U14180 (N_14180,N_12814,N_13465);
and U14181 (N_14181,N_13153,N_13075);
and U14182 (N_14182,N_12564,N_12202);
xnor U14183 (N_14183,N_13176,N_12759);
or U14184 (N_14184,N_12292,N_13138);
nor U14185 (N_14185,N_12366,N_12734);
nor U14186 (N_14186,N_12450,N_12760);
nand U14187 (N_14187,N_13357,N_12287);
nand U14188 (N_14188,N_12347,N_13000);
xnor U14189 (N_14189,N_13492,N_12454);
nand U14190 (N_14190,N_13259,N_12979);
nor U14191 (N_14191,N_12840,N_13202);
nor U14192 (N_14192,N_12604,N_13386);
nor U14193 (N_14193,N_13397,N_13292);
nor U14194 (N_14194,N_12905,N_13048);
nand U14195 (N_14195,N_12118,N_13333);
nand U14196 (N_14196,N_13450,N_13089);
or U14197 (N_14197,N_13065,N_13295);
or U14198 (N_14198,N_13082,N_13096);
or U14199 (N_14199,N_12249,N_12207);
or U14200 (N_14200,N_13300,N_12545);
nand U14201 (N_14201,N_12741,N_12716);
nor U14202 (N_14202,N_12865,N_12396);
nor U14203 (N_14203,N_12319,N_13217);
nor U14204 (N_14204,N_12797,N_12167);
or U14205 (N_14205,N_13415,N_12083);
and U14206 (N_14206,N_13108,N_12885);
nor U14207 (N_14207,N_13468,N_13189);
nand U14208 (N_14208,N_13134,N_13360);
nand U14209 (N_14209,N_12550,N_12880);
and U14210 (N_14210,N_12392,N_12858);
or U14211 (N_14211,N_13277,N_12290);
and U14212 (N_14212,N_13363,N_12770);
xor U14213 (N_14213,N_12363,N_12044);
or U14214 (N_14214,N_12018,N_12501);
or U14215 (N_14215,N_12088,N_12544);
nand U14216 (N_14216,N_13395,N_13243);
xnor U14217 (N_14217,N_13388,N_12547);
and U14218 (N_14218,N_12634,N_13088);
or U14219 (N_14219,N_12663,N_12125);
nand U14220 (N_14220,N_12214,N_12612);
or U14221 (N_14221,N_13110,N_12958);
and U14222 (N_14222,N_13272,N_12594);
nor U14223 (N_14223,N_12159,N_12418);
or U14224 (N_14224,N_12836,N_13068);
and U14225 (N_14225,N_12706,N_12625);
or U14226 (N_14226,N_13227,N_12374);
nand U14227 (N_14227,N_12078,N_12473);
and U14228 (N_14228,N_13429,N_12667);
and U14229 (N_14229,N_12974,N_12046);
and U14230 (N_14230,N_12033,N_13287);
and U14231 (N_14231,N_13074,N_13302);
or U14232 (N_14232,N_13200,N_12461);
and U14233 (N_14233,N_12371,N_12035);
nand U14234 (N_14234,N_12000,N_13228);
nand U14235 (N_14235,N_12843,N_13495);
or U14236 (N_14236,N_12791,N_12603);
or U14237 (N_14237,N_12597,N_13183);
and U14238 (N_14238,N_12117,N_13174);
nand U14239 (N_14239,N_13124,N_13236);
and U14240 (N_14240,N_12819,N_12623);
nor U14241 (N_14241,N_12173,N_12732);
nand U14242 (N_14242,N_12898,N_13107);
nor U14243 (N_14243,N_12029,N_13310);
or U14244 (N_14244,N_12852,N_13443);
or U14245 (N_14245,N_12784,N_12529);
xnor U14246 (N_14246,N_12137,N_12314);
xor U14247 (N_14247,N_13378,N_13163);
nand U14248 (N_14248,N_12066,N_13373);
or U14249 (N_14249,N_12886,N_12626);
or U14250 (N_14250,N_12797,N_12664);
or U14251 (N_14251,N_12316,N_12501);
nand U14252 (N_14252,N_12849,N_12597);
nand U14253 (N_14253,N_12862,N_12406);
xnor U14254 (N_14254,N_12210,N_12116);
xor U14255 (N_14255,N_12355,N_13101);
xnor U14256 (N_14256,N_12840,N_12542);
nand U14257 (N_14257,N_12036,N_12307);
and U14258 (N_14258,N_12514,N_13348);
nand U14259 (N_14259,N_12140,N_13483);
or U14260 (N_14260,N_12382,N_13334);
nor U14261 (N_14261,N_13176,N_12214);
or U14262 (N_14262,N_13485,N_12524);
nor U14263 (N_14263,N_12036,N_13136);
and U14264 (N_14264,N_12208,N_12393);
and U14265 (N_14265,N_12449,N_13302);
and U14266 (N_14266,N_13484,N_13152);
nor U14267 (N_14267,N_12833,N_13353);
nor U14268 (N_14268,N_13255,N_13089);
nand U14269 (N_14269,N_12130,N_13179);
nor U14270 (N_14270,N_12813,N_12000);
nand U14271 (N_14271,N_13389,N_13472);
nor U14272 (N_14272,N_12216,N_13107);
nand U14273 (N_14273,N_12377,N_12317);
and U14274 (N_14274,N_12584,N_12593);
nand U14275 (N_14275,N_12007,N_12640);
nor U14276 (N_14276,N_12117,N_12763);
or U14277 (N_14277,N_12374,N_12291);
or U14278 (N_14278,N_12825,N_12278);
nand U14279 (N_14279,N_13475,N_13126);
or U14280 (N_14280,N_12946,N_12738);
nand U14281 (N_14281,N_12560,N_12345);
or U14282 (N_14282,N_13453,N_12602);
and U14283 (N_14283,N_12662,N_12820);
nand U14284 (N_14284,N_13192,N_13028);
or U14285 (N_14285,N_12511,N_12654);
and U14286 (N_14286,N_12049,N_12466);
or U14287 (N_14287,N_12764,N_13191);
and U14288 (N_14288,N_12983,N_13275);
or U14289 (N_14289,N_12746,N_12969);
and U14290 (N_14290,N_13214,N_12749);
and U14291 (N_14291,N_13093,N_12817);
and U14292 (N_14292,N_12598,N_12969);
nand U14293 (N_14293,N_13182,N_12371);
and U14294 (N_14294,N_13385,N_12598);
nor U14295 (N_14295,N_12551,N_13291);
nand U14296 (N_14296,N_12012,N_12557);
nor U14297 (N_14297,N_12138,N_12680);
or U14298 (N_14298,N_13475,N_12548);
nand U14299 (N_14299,N_12176,N_12566);
or U14300 (N_14300,N_12634,N_13408);
nand U14301 (N_14301,N_12533,N_13266);
and U14302 (N_14302,N_12304,N_12735);
and U14303 (N_14303,N_12823,N_12367);
nand U14304 (N_14304,N_12556,N_13497);
nand U14305 (N_14305,N_12440,N_13254);
or U14306 (N_14306,N_12641,N_13267);
and U14307 (N_14307,N_12795,N_12694);
nand U14308 (N_14308,N_12972,N_13339);
and U14309 (N_14309,N_13402,N_12932);
nor U14310 (N_14310,N_13195,N_12349);
nand U14311 (N_14311,N_12060,N_12498);
nand U14312 (N_14312,N_12383,N_13300);
xor U14313 (N_14313,N_12074,N_12706);
or U14314 (N_14314,N_13245,N_12474);
nand U14315 (N_14315,N_12106,N_12851);
and U14316 (N_14316,N_13191,N_12921);
nand U14317 (N_14317,N_12919,N_13170);
nor U14318 (N_14318,N_12206,N_12014);
nand U14319 (N_14319,N_12481,N_13392);
nand U14320 (N_14320,N_12451,N_13149);
nand U14321 (N_14321,N_12043,N_12079);
xnor U14322 (N_14322,N_13478,N_12071);
or U14323 (N_14323,N_13307,N_13238);
or U14324 (N_14324,N_13167,N_13117);
and U14325 (N_14325,N_13433,N_12524);
or U14326 (N_14326,N_12847,N_13411);
and U14327 (N_14327,N_12934,N_13030);
and U14328 (N_14328,N_12589,N_12580);
nor U14329 (N_14329,N_13298,N_13253);
nor U14330 (N_14330,N_12239,N_12889);
nor U14331 (N_14331,N_12318,N_12472);
or U14332 (N_14332,N_12964,N_12396);
or U14333 (N_14333,N_13166,N_12749);
nor U14334 (N_14334,N_12759,N_13411);
xor U14335 (N_14335,N_13060,N_12152);
nand U14336 (N_14336,N_12660,N_12913);
or U14337 (N_14337,N_12413,N_13455);
or U14338 (N_14338,N_12630,N_12681);
or U14339 (N_14339,N_12749,N_12456);
and U14340 (N_14340,N_12445,N_13188);
nand U14341 (N_14341,N_12597,N_13490);
and U14342 (N_14342,N_12820,N_13461);
xnor U14343 (N_14343,N_12493,N_13237);
and U14344 (N_14344,N_12190,N_13032);
and U14345 (N_14345,N_12723,N_12414);
and U14346 (N_14346,N_13393,N_12605);
xor U14347 (N_14347,N_12500,N_13006);
xnor U14348 (N_14348,N_12446,N_12310);
and U14349 (N_14349,N_12120,N_12812);
xnor U14350 (N_14350,N_12838,N_13470);
and U14351 (N_14351,N_13084,N_12064);
nand U14352 (N_14352,N_12887,N_12974);
nor U14353 (N_14353,N_12042,N_13104);
nand U14354 (N_14354,N_12514,N_12164);
or U14355 (N_14355,N_12481,N_12828);
nand U14356 (N_14356,N_13128,N_13080);
nand U14357 (N_14357,N_13308,N_13087);
or U14358 (N_14358,N_12902,N_13484);
xor U14359 (N_14359,N_12081,N_12014);
or U14360 (N_14360,N_13185,N_13338);
nor U14361 (N_14361,N_13124,N_12413);
and U14362 (N_14362,N_12961,N_12212);
and U14363 (N_14363,N_13083,N_12513);
nor U14364 (N_14364,N_12000,N_12690);
nand U14365 (N_14365,N_13077,N_13004);
nor U14366 (N_14366,N_12497,N_12621);
and U14367 (N_14367,N_12368,N_12638);
nor U14368 (N_14368,N_13199,N_12141);
xor U14369 (N_14369,N_12133,N_13402);
nand U14370 (N_14370,N_12036,N_12612);
or U14371 (N_14371,N_12652,N_12844);
nor U14372 (N_14372,N_12799,N_12846);
nor U14373 (N_14373,N_12320,N_12118);
or U14374 (N_14374,N_12363,N_12256);
and U14375 (N_14375,N_13031,N_13071);
or U14376 (N_14376,N_12750,N_13091);
and U14377 (N_14377,N_12173,N_12245);
nand U14378 (N_14378,N_12276,N_12739);
nor U14379 (N_14379,N_12260,N_12266);
nor U14380 (N_14380,N_12489,N_13171);
or U14381 (N_14381,N_13117,N_12248);
nor U14382 (N_14382,N_12062,N_13069);
nor U14383 (N_14383,N_12387,N_13071);
nand U14384 (N_14384,N_13029,N_12571);
or U14385 (N_14385,N_12762,N_12184);
nor U14386 (N_14386,N_12543,N_12536);
or U14387 (N_14387,N_13073,N_13198);
or U14388 (N_14388,N_12000,N_12414);
nand U14389 (N_14389,N_12217,N_13227);
nand U14390 (N_14390,N_12008,N_13258);
nand U14391 (N_14391,N_12028,N_12063);
or U14392 (N_14392,N_12982,N_13469);
and U14393 (N_14393,N_12402,N_12064);
or U14394 (N_14394,N_13452,N_12207);
nor U14395 (N_14395,N_12159,N_13133);
or U14396 (N_14396,N_12286,N_12589);
and U14397 (N_14397,N_12012,N_12490);
or U14398 (N_14398,N_12616,N_12379);
nor U14399 (N_14399,N_13385,N_13294);
and U14400 (N_14400,N_12117,N_13348);
and U14401 (N_14401,N_13311,N_12561);
nand U14402 (N_14402,N_12158,N_12015);
and U14403 (N_14403,N_13087,N_12851);
nand U14404 (N_14404,N_12143,N_12132);
nor U14405 (N_14405,N_13307,N_12342);
nand U14406 (N_14406,N_13083,N_13004);
or U14407 (N_14407,N_12918,N_13342);
nor U14408 (N_14408,N_13129,N_13120);
or U14409 (N_14409,N_12010,N_12064);
nand U14410 (N_14410,N_13130,N_12724);
or U14411 (N_14411,N_12313,N_12416);
nand U14412 (N_14412,N_13203,N_13478);
nor U14413 (N_14413,N_12229,N_12100);
and U14414 (N_14414,N_12226,N_12337);
nor U14415 (N_14415,N_12681,N_13381);
nand U14416 (N_14416,N_13373,N_12772);
and U14417 (N_14417,N_12727,N_12297);
or U14418 (N_14418,N_12765,N_13120);
nor U14419 (N_14419,N_13120,N_12838);
nand U14420 (N_14420,N_12447,N_12753);
and U14421 (N_14421,N_13440,N_12441);
nor U14422 (N_14422,N_12596,N_12558);
nand U14423 (N_14423,N_12959,N_12462);
nor U14424 (N_14424,N_12439,N_12275);
nor U14425 (N_14425,N_13086,N_12337);
or U14426 (N_14426,N_13480,N_13250);
nor U14427 (N_14427,N_12307,N_12560);
and U14428 (N_14428,N_13162,N_13191);
nor U14429 (N_14429,N_13142,N_12925);
or U14430 (N_14430,N_12663,N_12814);
xor U14431 (N_14431,N_12645,N_12905);
or U14432 (N_14432,N_13130,N_12104);
or U14433 (N_14433,N_13416,N_12598);
nor U14434 (N_14434,N_12634,N_13373);
and U14435 (N_14435,N_12236,N_12463);
nand U14436 (N_14436,N_12255,N_13016);
nor U14437 (N_14437,N_13108,N_12340);
and U14438 (N_14438,N_13117,N_12474);
nand U14439 (N_14439,N_12003,N_12657);
or U14440 (N_14440,N_12642,N_13404);
nand U14441 (N_14441,N_13031,N_12664);
xor U14442 (N_14442,N_12800,N_13055);
nand U14443 (N_14443,N_13311,N_12016);
and U14444 (N_14444,N_12220,N_12993);
and U14445 (N_14445,N_12331,N_12814);
nand U14446 (N_14446,N_12937,N_12241);
or U14447 (N_14447,N_12630,N_12895);
nand U14448 (N_14448,N_12693,N_13211);
and U14449 (N_14449,N_13409,N_12949);
xnor U14450 (N_14450,N_12033,N_13129);
nor U14451 (N_14451,N_12729,N_12937);
nor U14452 (N_14452,N_12764,N_12218);
and U14453 (N_14453,N_12344,N_13415);
xnor U14454 (N_14454,N_13491,N_12263);
nand U14455 (N_14455,N_12236,N_12640);
or U14456 (N_14456,N_13493,N_12288);
nor U14457 (N_14457,N_12920,N_12849);
or U14458 (N_14458,N_13141,N_12318);
or U14459 (N_14459,N_12380,N_12852);
or U14460 (N_14460,N_12424,N_12249);
nand U14461 (N_14461,N_13059,N_12979);
nor U14462 (N_14462,N_12494,N_12679);
nor U14463 (N_14463,N_12800,N_12257);
and U14464 (N_14464,N_12153,N_12296);
and U14465 (N_14465,N_12760,N_12384);
xor U14466 (N_14466,N_12258,N_12153);
nor U14467 (N_14467,N_12527,N_12999);
nand U14468 (N_14468,N_12515,N_12019);
and U14469 (N_14469,N_12794,N_12012);
xor U14470 (N_14470,N_13306,N_12907);
nand U14471 (N_14471,N_12985,N_12736);
nor U14472 (N_14472,N_12275,N_12887);
nor U14473 (N_14473,N_12722,N_13499);
nor U14474 (N_14474,N_12990,N_13352);
and U14475 (N_14475,N_12666,N_12153);
and U14476 (N_14476,N_13420,N_12446);
xor U14477 (N_14477,N_13309,N_12395);
or U14478 (N_14478,N_12820,N_12213);
and U14479 (N_14479,N_13067,N_13419);
nand U14480 (N_14480,N_12876,N_13370);
nor U14481 (N_14481,N_12546,N_12176);
or U14482 (N_14482,N_12327,N_13029);
or U14483 (N_14483,N_12484,N_12138);
xor U14484 (N_14484,N_13218,N_12897);
nor U14485 (N_14485,N_12102,N_13377);
and U14486 (N_14486,N_13226,N_12357);
nand U14487 (N_14487,N_12360,N_12661);
nor U14488 (N_14488,N_13059,N_12502);
nor U14489 (N_14489,N_12547,N_12725);
or U14490 (N_14490,N_13133,N_12926);
and U14491 (N_14491,N_12892,N_13314);
and U14492 (N_14492,N_12779,N_12980);
nand U14493 (N_14493,N_12890,N_12752);
or U14494 (N_14494,N_12659,N_12999);
nand U14495 (N_14495,N_12633,N_13272);
nand U14496 (N_14496,N_12841,N_13146);
nor U14497 (N_14497,N_12401,N_13025);
or U14498 (N_14498,N_12160,N_13449);
and U14499 (N_14499,N_13244,N_13219);
nor U14500 (N_14500,N_12781,N_12806);
nor U14501 (N_14501,N_12580,N_12690);
nand U14502 (N_14502,N_12958,N_13459);
nor U14503 (N_14503,N_12686,N_12993);
nand U14504 (N_14504,N_13078,N_13268);
nand U14505 (N_14505,N_13416,N_12150);
or U14506 (N_14506,N_12670,N_12834);
or U14507 (N_14507,N_12211,N_12130);
nor U14508 (N_14508,N_13051,N_13129);
nor U14509 (N_14509,N_12898,N_12434);
nand U14510 (N_14510,N_12466,N_12374);
nor U14511 (N_14511,N_12072,N_12147);
or U14512 (N_14512,N_12743,N_12919);
and U14513 (N_14513,N_12468,N_12898);
and U14514 (N_14514,N_13389,N_12240);
nor U14515 (N_14515,N_12241,N_12498);
or U14516 (N_14516,N_12787,N_12112);
and U14517 (N_14517,N_13235,N_13275);
and U14518 (N_14518,N_12134,N_12585);
nand U14519 (N_14519,N_12610,N_12954);
nor U14520 (N_14520,N_13156,N_12812);
nand U14521 (N_14521,N_13344,N_12242);
nand U14522 (N_14522,N_12308,N_12377);
and U14523 (N_14523,N_12853,N_12397);
and U14524 (N_14524,N_13307,N_13226);
nor U14525 (N_14525,N_12915,N_13275);
nand U14526 (N_14526,N_12179,N_13137);
or U14527 (N_14527,N_13054,N_12042);
or U14528 (N_14528,N_12647,N_12963);
or U14529 (N_14529,N_13481,N_12399);
nor U14530 (N_14530,N_12646,N_13127);
nor U14531 (N_14531,N_12897,N_13190);
or U14532 (N_14532,N_12824,N_12143);
nand U14533 (N_14533,N_13489,N_12221);
nand U14534 (N_14534,N_12142,N_12767);
and U14535 (N_14535,N_12616,N_12099);
and U14536 (N_14536,N_12308,N_12025);
or U14537 (N_14537,N_13366,N_12081);
nor U14538 (N_14538,N_13183,N_12390);
nand U14539 (N_14539,N_12891,N_12338);
or U14540 (N_14540,N_12813,N_12273);
nand U14541 (N_14541,N_12640,N_12913);
and U14542 (N_14542,N_13243,N_12911);
nor U14543 (N_14543,N_12876,N_12209);
nor U14544 (N_14544,N_12440,N_12120);
or U14545 (N_14545,N_12030,N_12334);
nor U14546 (N_14546,N_12564,N_12628);
or U14547 (N_14547,N_13450,N_13061);
and U14548 (N_14548,N_13341,N_13449);
nand U14549 (N_14549,N_12718,N_12303);
or U14550 (N_14550,N_12254,N_12492);
or U14551 (N_14551,N_12070,N_12871);
nor U14552 (N_14552,N_12212,N_12981);
or U14553 (N_14553,N_12888,N_12499);
and U14554 (N_14554,N_13354,N_12983);
and U14555 (N_14555,N_12339,N_12718);
nand U14556 (N_14556,N_13331,N_12466);
xnor U14557 (N_14557,N_12897,N_13351);
or U14558 (N_14558,N_12897,N_12730);
and U14559 (N_14559,N_12587,N_13319);
or U14560 (N_14560,N_12242,N_12807);
or U14561 (N_14561,N_13272,N_12215);
xor U14562 (N_14562,N_12121,N_13344);
nor U14563 (N_14563,N_13101,N_12300);
or U14564 (N_14564,N_12277,N_12282);
nand U14565 (N_14565,N_12096,N_12437);
and U14566 (N_14566,N_13164,N_13303);
nand U14567 (N_14567,N_12422,N_12977);
nor U14568 (N_14568,N_13298,N_12208);
nand U14569 (N_14569,N_13027,N_13167);
and U14570 (N_14570,N_12098,N_12603);
and U14571 (N_14571,N_13124,N_12083);
and U14572 (N_14572,N_12162,N_12387);
or U14573 (N_14573,N_13162,N_12751);
and U14574 (N_14574,N_13489,N_12588);
and U14575 (N_14575,N_12347,N_12932);
nor U14576 (N_14576,N_12804,N_12853);
or U14577 (N_14577,N_12260,N_12559);
or U14578 (N_14578,N_12508,N_13439);
and U14579 (N_14579,N_13209,N_13172);
or U14580 (N_14580,N_12550,N_12626);
nand U14581 (N_14581,N_12440,N_12250);
nor U14582 (N_14582,N_12979,N_12789);
nand U14583 (N_14583,N_12307,N_12185);
or U14584 (N_14584,N_12345,N_12895);
nand U14585 (N_14585,N_12088,N_12542);
or U14586 (N_14586,N_12374,N_12789);
and U14587 (N_14587,N_13157,N_13259);
xor U14588 (N_14588,N_13426,N_12928);
and U14589 (N_14589,N_12851,N_12134);
and U14590 (N_14590,N_12708,N_12698);
and U14591 (N_14591,N_13305,N_12429);
nor U14592 (N_14592,N_13039,N_12906);
nor U14593 (N_14593,N_12866,N_12628);
or U14594 (N_14594,N_12292,N_12316);
nand U14595 (N_14595,N_13434,N_12420);
and U14596 (N_14596,N_13320,N_12929);
or U14597 (N_14597,N_13472,N_12784);
nand U14598 (N_14598,N_13264,N_12060);
or U14599 (N_14599,N_12335,N_13206);
or U14600 (N_14600,N_13444,N_12413);
or U14601 (N_14601,N_12866,N_12751);
nand U14602 (N_14602,N_13217,N_12210);
nor U14603 (N_14603,N_12820,N_12119);
xnor U14604 (N_14604,N_12368,N_12072);
nor U14605 (N_14605,N_12472,N_12597);
nor U14606 (N_14606,N_13006,N_12036);
nand U14607 (N_14607,N_12417,N_12896);
or U14608 (N_14608,N_12491,N_12359);
or U14609 (N_14609,N_12137,N_12311);
xor U14610 (N_14610,N_12166,N_12769);
and U14611 (N_14611,N_12924,N_13420);
nor U14612 (N_14612,N_12085,N_12293);
and U14613 (N_14613,N_12052,N_13037);
nor U14614 (N_14614,N_13374,N_13184);
nor U14615 (N_14615,N_12352,N_13233);
nand U14616 (N_14616,N_12042,N_13299);
nand U14617 (N_14617,N_12763,N_12966);
and U14618 (N_14618,N_12234,N_12350);
nor U14619 (N_14619,N_12109,N_12610);
nor U14620 (N_14620,N_12853,N_12310);
nor U14621 (N_14621,N_12340,N_12493);
nand U14622 (N_14622,N_12402,N_12997);
nor U14623 (N_14623,N_12912,N_12629);
or U14624 (N_14624,N_12145,N_12105);
or U14625 (N_14625,N_12991,N_12664);
or U14626 (N_14626,N_13172,N_12089);
and U14627 (N_14627,N_12245,N_13229);
or U14628 (N_14628,N_12406,N_12006);
nand U14629 (N_14629,N_12897,N_12029);
and U14630 (N_14630,N_12760,N_12952);
nand U14631 (N_14631,N_13269,N_13440);
or U14632 (N_14632,N_12300,N_12913);
nand U14633 (N_14633,N_12430,N_13254);
nor U14634 (N_14634,N_13065,N_13120);
and U14635 (N_14635,N_12542,N_13006);
and U14636 (N_14636,N_12965,N_13076);
nand U14637 (N_14637,N_12456,N_12082);
nor U14638 (N_14638,N_12278,N_12219);
or U14639 (N_14639,N_12147,N_12708);
or U14640 (N_14640,N_12786,N_12039);
nor U14641 (N_14641,N_12655,N_12858);
and U14642 (N_14642,N_13242,N_12248);
nor U14643 (N_14643,N_12992,N_12498);
nor U14644 (N_14644,N_12598,N_12359);
or U14645 (N_14645,N_13186,N_12773);
nand U14646 (N_14646,N_13452,N_12046);
and U14647 (N_14647,N_13340,N_13424);
or U14648 (N_14648,N_13486,N_13167);
nor U14649 (N_14649,N_12633,N_13277);
nand U14650 (N_14650,N_13050,N_12336);
and U14651 (N_14651,N_13058,N_12695);
nor U14652 (N_14652,N_12954,N_13391);
nand U14653 (N_14653,N_13051,N_12246);
nand U14654 (N_14654,N_13475,N_12530);
nor U14655 (N_14655,N_12700,N_12413);
and U14656 (N_14656,N_13147,N_12996);
nor U14657 (N_14657,N_12607,N_12810);
xnor U14658 (N_14658,N_12002,N_13001);
nand U14659 (N_14659,N_12398,N_12935);
and U14660 (N_14660,N_13487,N_13405);
and U14661 (N_14661,N_12568,N_12030);
and U14662 (N_14662,N_12825,N_13188);
nor U14663 (N_14663,N_13199,N_12172);
or U14664 (N_14664,N_12825,N_12213);
nor U14665 (N_14665,N_12927,N_12171);
or U14666 (N_14666,N_13493,N_12279);
nor U14667 (N_14667,N_13314,N_12314);
and U14668 (N_14668,N_12466,N_12559);
nand U14669 (N_14669,N_13000,N_13139);
nand U14670 (N_14670,N_13180,N_13350);
nand U14671 (N_14671,N_12504,N_12616);
and U14672 (N_14672,N_12346,N_12859);
nand U14673 (N_14673,N_12760,N_12089);
or U14674 (N_14674,N_13340,N_13409);
and U14675 (N_14675,N_13344,N_12054);
and U14676 (N_14676,N_12626,N_12712);
nand U14677 (N_14677,N_12715,N_12801);
nand U14678 (N_14678,N_13029,N_12795);
nand U14679 (N_14679,N_12156,N_12108);
nor U14680 (N_14680,N_13213,N_12593);
and U14681 (N_14681,N_13337,N_12295);
and U14682 (N_14682,N_13147,N_13297);
nand U14683 (N_14683,N_12773,N_12736);
xnor U14684 (N_14684,N_12514,N_12675);
or U14685 (N_14685,N_13267,N_12213);
nand U14686 (N_14686,N_12737,N_12243);
nor U14687 (N_14687,N_13127,N_12238);
nand U14688 (N_14688,N_13152,N_12504);
xor U14689 (N_14689,N_12361,N_13342);
and U14690 (N_14690,N_12152,N_12104);
and U14691 (N_14691,N_13413,N_13133);
nor U14692 (N_14692,N_12826,N_12750);
nand U14693 (N_14693,N_13431,N_13382);
nand U14694 (N_14694,N_12975,N_13495);
nand U14695 (N_14695,N_13349,N_13368);
nand U14696 (N_14696,N_13309,N_12582);
or U14697 (N_14697,N_13373,N_12114);
and U14698 (N_14698,N_12517,N_12494);
nor U14699 (N_14699,N_12022,N_13080);
or U14700 (N_14700,N_13089,N_12639);
or U14701 (N_14701,N_12484,N_12491);
nand U14702 (N_14702,N_12349,N_12192);
nor U14703 (N_14703,N_12090,N_12015);
nor U14704 (N_14704,N_12901,N_13091);
and U14705 (N_14705,N_12253,N_12072);
nand U14706 (N_14706,N_12438,N_12102);
and U14707 (N_14707,N_12415,N_12426);
nand U14708 (N_14708,N_13081,N_12972);
nor U14709 (N_14709,N_12340,N_13168);
and U14710 (N_14710,N_12426,N_12242);
nand U14711 (N_14711,N_12725,N_13472);
nand U14712 (N_14712,N_12187,N_12703);
nor U14713 (N_14713,N_12920,N_12234);
nor U14714 (N_14714,N_13205,N_12458);
nand U14715 (N_14715,N_12640,N_13344);
nand U14716 (N_14716,N_13064,N_12666);
nor U14717 (N_14717,N_13059,N_12873);
nand U14718 (N_14718,N_13090,N_13258);
nand U14719 (N_14719,N_12286,N_12910);
nor U14720 (N_14720,N_12453,N_13149);
nand U14721 (N_14721,N_12647,N_13463);
nand U14722 (N_14722,N_13043,N_12083);
and U14723 (N_14723,N_13483,N_12163);
and U14724 (N_14724,N_13382,N_13076);
nand U14725 (N_14725,N_12060,N_13196);
or U14726 (N_14726,N_12079,N_12826);
xnor U14727 (N_14727,N_12511,N_12438);
nand U14728 (N_14728,N_12605,N_12041);
nand U14729 (N_14729,N_12684,N_12767);
xor U14730 (N_14730,N_13235,N_12102);
xnor U14731 (N_14731,N_12450,N_13478);
nor U14732 (N_14732,N_13076,N_12374);
or U14733 (N_14733,N_12159,N_12124);
or U14734 (N_14734,N_12366,N_12362);
or U14735 (N_14735,N_12688,N_12067);
nand U14736 (N_14736,N_12289,N_13125);
and U14737 (N_14737,N_13439,N_13345);
and U14738 (N_14738,N_13278,N_13098);
nand U14739 (N_14739,N_12398,N_12640);
and U14740 (N_14740,N_12944,N_12664);
or U14741 (N_14741,N_13413,N_12442);
nand U14742 (N_14742,N_12011,N_12773);
or U14743 (N_14743,N_13318,N_12306);
nand U14744 (N_14744,N_13076,N_13209);
and U14745 (N_14745,N_12544,N_12733);
nand U14746 (N_14746,N_12112,N_12147);
and U14747 (N_14747,N_13430,N_12441);
and U14748 (N_14748,N_13320,N_13385);
or U14749 (N_14749,N_12516,N_12102);
xnor U14750 (N_14750,N_12150,N_12839);
nor U14751 (N_14751,N_12450,N_13312);
nor U14752 (N_14752,N_13452,N_13475);
nand U14753 (N_14753,N_12929,N_12396);
and U14754 (N_14754,N_12651,N_13177);
and U14755 (N_14755,N_12216,N_12376);
or U14756 (N_14756,N_12462,N_13042);
nor U14757 (N_14757,N_12723,N_12604);
and U14758 (N_14758,N_12799,N_12796);
nor U14759 (N_14759,N_13132,N_12871);
xor U14760 (N_14760,N_12322,N_13098);
nand U14761 (N_14761,N_12100,N_12895);
or U14762 (N_14762,N_12739,N_12094);
nor U14763 (N_14763,N_12729,N_13381);
xnor U14764 (N_14764,N_12777,N_13397);
and U14765 (N_14765,N_12976,N_12647);
nand U14766 (N_14766,N_12908,N_12737);
or U14767 (N_14767,N_13490,N_12711);
or U14768 (N_14768,N_12772,N_12952);
nand U14769 (N_14769,N_12638,N_12669);
or U14770 (N_14770,N_13358,N_12621);
nand U14771 (N_14771,N_13239,N_12474);
and U14772 (N_14772,N_12737,N_12550);
or U14773 (N_14773,N_12538,N_12743);
and U14774 (N_14774,N_13246,N_13047);
or U14775 (N_14775,N_12189,N_12350);
nand U14776 (N_14776,N_12450,N_12807);
xnor U14777 (N_14777,N_13471,N_12862);
xnor U14778 (N_14778,N_13233,N_12492);
nor U14779 (N_14779,N_13273,N_12344);
and U14780 (N_14780,N_12804,N_12222);
xor U14781 (N_14781,N_12841,N_12773);
or U14782 (N_14782,N_12486,N_13307);
nand U14783 (N_14783,N_13151,N_13366);
xor U14784 (N_14784,N_12080,N_12247);
nor U14785 (N_14785,N_12339,N_12366);
or U14786 (N_14786,N_12865,N_13084);
and U14787 (N_14787,N_13233,N_13002);
or U14788 (N_14788,N_13114,N_12125);
or U14789 (N_14789,N_12878,N_12347);
and U14790 (N_14790,N_12985,N_12228);
nor U14791 (N_14791,N_12906,N_12196);
and U14792 (N_14792,N_12530,N_12045);
or U14793 (N_14793,N_13306,N_13455);
and U14794 (N_14794,N_12043,N_12134);
nand U14795 (N_14795,N_12760,N_13030);
or U14796 (N_14796,N_12198,N_12271);
or U14797 (N_14797,N_12443,N_13203);
nor U14798 (N_14798,N_12825,N_13091);
nor U14799 (N_14799,N_12902,N_12460);
and U14800 (N_14800,N_12999,N_13000);
nand U14801 (N_14801,N_12895,N_13149);
or U14802 (N_14802,N_12808,N_12856);
and U14803 (N_14803,N_13010,N_12389);
and U14804 (N_14804,N_12764,N_13083);
nand U14805 (N_14805,N_12011,N_12152);
and U14806 (N_14806,N_12218,N_12943);
nand U14807 (N_14807,N_12478,N_12101);
and U14808 (N_14808,N_12872,N_13375);
nand U14809 (N_14809,N_13398,N_12764);
nor U14810 (N_14810,N_13091,N_12257);
and U14811 (N_14811,N_12807,N_12702);
and U14812 (N_14812,N_13146,N_12894);
or U14813 (N_14813,N_13295,N_13296);
nor U14814 (N_14814,N_13058,N_12989);
xor U14815 (N_14815,N_12114,N_12121);
xnor U14816 (N_14816,N_12042,N_12149);
or U14817 (N_14817,N_12726,N_12897);
nor U14818 (N_14818,N_13184,N_12152);
nor U14819 (N_14819,N_12771,N_12474);
nor U14820 (N_14820,N_12905,N_13327);
and U14821 (N_14821,N_13321,N_12578);
nor U14822 (N_14822,N_13198,N_13476);
or U14823 (N_14823,N_12887,N_13053);
nand U14824 (N_14824,N_12722,N_13075);
nor U14825 (N_14825,N_12562,N_12172);
or U14826 (N_14826,N_12097,N_12131);
xor U14827 (N_14827,N_12216,N_12634);
nand U14828 (N_14828,N_12946,N_12406);
nand U14829 (N_14829,N_12886,N_12960);
nand U14830 (N_14830,N_12035,N_12545);
nor U14831 (N_14831,N_12175,N_12711);
and U14832 (N_14832,N_12449,N_12485);
or U14833 (N_14833,N_12669,N_12537);
nor U14834 (N_14834,N_12838,N_13133);
nor U14835 (N_14835,N_12185,N_12804);
nor U14836 (N_14836,N_12867,N_12040);
and U14837 (N_14837,N_12147,N_12613);
and U14838 (N_14838,N_12155,N_12739);
xor U14839 (N_14839,N_13111,N_13368);
nor U14840 (N_14840,N_12302,N_12198);
or U14841 (N_14841,N_13322,N_12222);
nand U14842 (N_14842,N_12133,N_12268);
nor U14843 (N_14843,N_13065,N_13430);
nor U14844 (N_14844,N_12984,N_12954);
nor U14845 (N_14845,N_12903,N_12980);
nor U14846 (N_14846,N_12670,N_12106);
and U14847 (N_14847,N_13441,N_12510);
xnor U14848 (N_14848,N_12001,N_12127);
and U14849 (N_14849,N_12267,N_12646);
or U14850 (N_14850,N_12069,N_12656);
and U14851 (N_14851,N_12066,N_12830);
nor U14852 (N_14852,N_12458,N_12401);
nor U14853 (N_14853,N_12047,N_12149);
or U14854 (N_14854,N_13474,N_12245);
nor U14855 (N_14855,N_12605,N_13083);
nor U14856 (N_14856,N_12752,N_13473);
or U14857 (N_14857,N_12043,N_12496);
nor U14858 (N_14858,N_12073,N_12975);
and U14859 (N_14859,N_13015,N_12121);
and U14860 (N_14860,N_12888,N_12983);
nand U14861 (N_14861,N_12775,N_12809);
and U14862 (N_14862,N_12980,N_13332);
nand U14863 (N_14863,N_12480,N_13320);
and U14864 (N_14864,N_12645,N_12532);
nand U14865 (N_14865,N_12676,N_12546);
xnor U14866 (N_14866,N_13466,N_12815);
or U14867 (N_14867,N_12087,N_12932);
or U14868 (N_14868,N_12352,N_13134);
and U14869 (N_14869,N_13291,N_12742);
and U14870 (N_14870,N_12458,N_12532);
or U14871 (N_14871,N_12161,N_12095);
nand U14872 (N_14872,N_12555,N_12152);
nor U14873 (N_14873,N_12905,N_12926);
or U14874 (N_14874,N_12807,N_12256);
nand U14875 (N_14875,N_13054,N_13371);
xnor U14876 (N_14876,N_12352,N_13190);
nand U14877 (N_14877,N_12678,N_12552);
nor U14878 (N_14878,N_12912,N_13444);
nand U14879 (N_14879,N_13147,N_12197);
xnor U14880 (N_14880,N_12600,N_13162);
nor U14881 (N_14881,N_12222,N_12196);
nor U14882 (N_14882,N_12180,N_12439);
and U14883 (N_14883,N_12835,N_13350);
and U14884 (N_14884,N_12371,N_12080);
or U14885 (N_14885,N_13143,N_12120);
nand U14886 (N_14886,N_13060,N_12816);
nor U14887 (N_14887,N_12488,N_12378);
nand U14888 (N_14888,N_13211,N_13009);
and U14889 (N_14889,N_13060,N_13113);
nand U14890 (N_14890,N_12812,N_13417);
nand U14891 (N_14891,N_13358,N_12581);
xnor U14892 (N_14892,N_13397,N_12167);
nor U14893 (N_14893,N_12347,N_13057);
nand U14894 (N_14894,N_12418,N_13073);
nor U14895 (N_14895,N_12115,N_12178);
nand U14896 (N_14896,N_12486,N_12073);
nand U14897 (N_14897,N_12430,N_12584);
or U14898 (N_14898,N_12255,N_12729);
nand U14899 (N_14899,N_12298,N_12790);
nor U14900 (N_14900,N_12565,N_13472);
or U14901 (N_14901,N_13056,N_13201);
nand U14902 (N_14902,N_12065,N_13113);
or U14903 (N_14903,N_13420,N_13330);
nand U14904 (N_14904,N_12197,N_13178);
nand U14905 (N_14905,N_13054,N_13425);
nand U14906 (N_14906,N_12846,N_12725);
xor U14907 (N_14907,N_12429,N_12650);
nor U14908 (N_14908,N_12709,N_12608);
and U14909 (N_14909,N_13172,N_13444);
and U14910 (N_14910,N_12907,N_12507);
or U14911 (N_14911,N_12873,N_12816);
nor U14912 (N_14912,N_12099,N_12525);
nor U14913 (N_14913,N_12055,N_12401);
and U14914 (N_14914,N_12381,N_12794);
or U14915 (N_14915,N_12370,N_12387);
xnor U14916 (N_14916,N_12476,N_12106);
nor U14917 (N_14917,N_12755,N_13442);
nor U14918 (N_14918,N_12868,N_12982);
nand U14919 (N_14919,N_13455,N_12747);
nand U14920 (N_14920,N_12554,N_12051);
and U14921 (N_14921,N_13062,N_13329);
and U14922 (N_14922,N_12883,N_13497);
nand U14923 (N_14923,N_13497,N_12634);
and U14924 (N_14924,N_12166,N_12273);
and U14925 (N_14925,N_12846,N_13308);
nor U14926 (N_14926,N_12237,N_13029);
and U14927 (N_14927,N_13367,N_12463);
nand U14928 (N_14928,N_13411,N_12051);
and U14929 (N_14929,N_12283,N_12893);
nand U14930 (N_14930,N_13309,N_13467);
and U14931 (N_14931,N_12644,N_12238);
nand U14932 (N_14932,N_13304,N_12749);
or U14933 (N_14933,N_12154,N_13172);
or U14934 (N_14934,N_13019,N_13333);
nor U14935 (N_14935,N_12087,N_12575);
and U14936 (N_14936,N_12046,N_12278);
nand U14937 (N_14937,N_12204,N_13429);
or U14938 (N_14938,N_13469,N_13400);
xor U14939 (N_14939,N_12653,N_12684);
and U14940 (N_14940,N_13393,N_12972);
and U14941 (N_14941,N_13199,N_12888);
nand U14942 (N_14942,N_12359,N_12124);
nand U14943 (N_14943,N_12172,N_13083);
xnor U14944 (N_14944,N_12055,N_12398);
and U14945 (N_14945,N_12537,N_13340);
or U14946 (N_14946,N_12415,N_12609);
or U14947 (N_14947,N_12198,N_12215);
or U14948 (N_14948,N_12804,N_12456);
and U14949 (N_14949,N_12691,N_12298);
nor U14950 (N_14950,N_12454,N_13345);
and U14951 (N_14951,N_13418,N_12412);
nor U14952 (N_14952,N_12371,N_12892);
nand U14953 (N_14953,N_12516,N_12375);
or U14954 (N_14954,N_13089,N_12360);
or U14955 (N_14955,N_12197,N_13144);
and U14956 (N_14956,N_13141,N_12297);
or U14957 (N_14957,N_12927,N_13445);
nand U14958 (N_14958,N_13395,N_12807);
or U14959 (N_14959,N_13249,N_13462);
or U14960 (N_14960,N_13408,N_13379);
and U14961 (N_14961,N_13264,N_13275);
nor U14962 (N_14962,N_12670,N_13454);
nor U14963 (N_14963,N_12236,N_12960);
or U14964 (N_14964,N_13030,N_13159);
and U14965 (N_14965,N_13397,N_12875);
or U14966 (N_14966,N_13247,N_13024);
and U14967 (N_14967,N_12555,N_12627);
or U14968 (N_14968,N_12787,N_12969);
nor U14969 (N_14969,N_12728,N_12666);
or U14970 (N_14970,N_13237,N_13493);
or U14971 (N_14971,N_12054,N_12789);
nor U14972 (N_14972,N_12467,N_13105);
nand U14973 (N_14973,N_13458,N_13249);
xnor U14974 (N_14974,N_12808,N_12200);
nand U14975 (N_14975,N_13020,N_12564);
and U14976 (N_14976,N_12120,N_13041);
xnor U14977 (N_14977,N_13219,N_12586);
or U14978 (N_14978,N_12100,N_12173);
nor U14979 (N_14979,N_12476,N_12443);
nand U14980 (N_14980,N_13060,N_12199);
nor U14981 (N_14981,N_12051,N_12852);
nand U14982 (N_14982,N_13104,N_12312);
or U14983 (N_14983,N_12213,N_12395);
or U14984 (N_14984,N_13190,N_12703);
or U14985 (N_14985,N_12364,N_12133);
or U14986 (N_14986,N_12907,N_13302);
nor U14987 (N_14987,N_12857,N_12381);
and U14988 (N_14988,N_13164,N_12053);
or U14989 (N_14989,N_12701,N_13208);
nor U14990 (N_14990,N_12421,N_13209);
xnor U14991 (N_14991,N_12815,N_13073);
nor U14992 (N_14992,N_13244,N_13237);
nor U14993 (N_14993,N_12333,N_13400);
nor U14994 (N_14994,N_13176,N_13234);
nand U14995 (N_14995,N_12210,N_13117);
nor U14996 (N_14996,N_13040,N_12426);
nand U14997 (N_14997,N_12134,N_12574);
nand U14998 (N_14998,N_12080,N_12806);
or U14999 (N_14999,N_12318,N_12018);
or UO_0 (O_0,N_13763,N_14413);
and UO_1 (O_1,N_14865,N_14866);
nand UO_2 (O_2,N_13652,N_13944);
or UO_3 (O_3,N_14989,N_13642);
nor UO_4 (O_4,N_14256,N_14429);
or UO_5 (O_5,N_14059,N_13843);
and UO_6 (O_6,N_14625,N_14703);
and UO_7 (O_7,N_13627,N_13599);
nor UO_8 (O_8,N_14292,N_14245);
nand UO_9 (O_9,N_13903,N_13578);
or UO_10 (O_10,N_14313,N_14115);
nor UO_11 (O_11,N_14590,N_13616);
nand UO_12 (O_12,N_14636,N_13511);
or UO_13 (O_13,N_13746,N_14119);
nand UO_14 (O_14,N_14139,N_13505);
nor UO_15 (O_15,N_14459,N_14233);
nor UO_16 (O_16,N_13753,N_14649);
nand UO_17 (O_17,N_13919,N_13555);
and UO_18 (O_18,N_13653,N_13928);
nor UO_19 (O_19,N_13974,N_14318);
nand UO_20 (O_20,N_14263,N_14030);
and UO_21 (O_21,N_13906,N_14653);
nand UO_22 (O_22,N_14879,N_14394);
nand UO_23 (O_23,N_14380,N_13697);
or UO_24 (O_24,N_14358,N_14972);
nor UO_25 (O_25,N_13856,N_13647);
or UO_26 (O_26,N_14600,N_14261);
and UO_27 (O_27,N_14094,N_13829);
nor UO_28 (O_28,N_14721,N_14247);
or UO_29 (O_29,N_14795,N_14383);
xnor UO_30 (O_30,N_14714,N_14638);
and UO_31 (O_31,N_14813,N_14251);
nor UO_32 (O_32,N_13585,N_14164);
nand UO_33 (O_33,N_13727,N_14230);
or UO_34 (O_34,N_13503,N_13962);
nand UO_35 (O_35,N_13879,N_14116);
nand UO_36 (O_36,N_14319,N_13813);
or UO_37 (O_37,N_14569,N_13814);
nor UO_38 (O_38,N_14255,N_14466);
or UO_39 (O_39,N_13776,N_14817);
xnor UO_40 (O_40,N_13563,N_14389);
xnor UO_41 (O_41,N_14099,N_13633);
nor UO_42 (O_42,N_13560,N_14190);
or UO_43 (O_43,N_13923,N_14808);
nor UO_44 (O_44,N_14180,N_14936);
and UO_45 (O_45,N_14927,N_14840);
nor UO_46 (O_46,N_14104,N_14008);
and UO_47 (O_47,N_13989,N_14914);
or UO_48 (O_48,N_14494,N_14411);
or UO_49 (O_49,N_13828,N_14526);
or UO_50 (O_50,N_14107,N_14607);
or UO_51 (O_51,N_14532,N_14929);
nand UO_52 (O_52,N_14432,N_14705);
nor UO_53 (O_53,N_14558,N_14020);
and UO_54 (O_54,N_14129,N_13971);
nand UO_55 (O_55,N_13899,N_14542);
nor UO_56 (O_56,N_13537,N_14696);
nor UO_57 (O_57,N_13562,N_13773);
nand UO_58 (O_58,N_14563,N_14983);
or UO_59 (O_59,N_14125,N_14279);
and UO_60 (O_60,N_14382,N_13739);
nor UO_61 (O_61,N_14652,N_14923);
or UO_62 (O_62,N_14039,N_13832);
nor UO_63 (O_63,N_14407,N_13655);
nor UO_64 (O_64,N_14743,N_14484);
and UO_65 (O_65,N_13876,N_14599);
or UO_66 (O_66,N_14856,N_14199);
xor UO_67 (O_67,N_13536,N_13918);
and UO_68 (O_68,N_13663,N_13566);
nor UO_69 (O_69,N_14527,N_14662);
and UO_70 (O_70,N_13869,N_14715);
nand UO_71 (O_71,N_14659,N_14033);
and UO_72 (O_72,N_13927,N_14476);
and UO_73 (O_73,N_14651,N_14453);
and UO_74 (O_74,N_14804,N_13966);
or UO_75 (O_75,N_13981,N_14304);
xnor UO_76 (O_76,N_13625,N_14246);
and UO_77 (O_77,N_13991,N_14471);
or UO_78 (O_78,N_14712,N_14658);
and UO_79 (O_79,N_14240,N_14406);
xnor UO_80 (O_80,N_14043,N_14242);
and UO_81 (O_81,N_14968,N_14928);
or UO_82 (O_82,N_13573,N_14177);
nor UO_83 (O_83,N_14193,N_14814);
or UO_84 (O_84,N_14064,N_14618);
and UO_85 (O_85,N_14663,N_14924);
nand UO_86 (O_86,N_13878,N_13531);
nor UO_87 (O_87,N_13985,N_13975);
or UO_88 (O_88,N_14275,N_14617);
or UO_89 (O_89,N_14492,N_13941);
and UO_90 (O_90,N_14974,N_14788);
nor UO_91 (O_91,N_14470,N_13925);
nand UO_92 (O_92,N_14462,N_14481);
nor UO_93 (O_93,N_14421,N_13586);
nor UO_94 (O_94,N_14294,N_13839);
or UO_95 (O_95,N_14214,N_13707);
and UO_96 (O_96,N_14037,N_14202);
nor UO_97 (O_97,N_14175,N_14244);
or UO_98 (O_98,N_14055,N_14533);
or UO_99 (O_99,N_14784,N_13608);
nor UO_100 (O_100,N_14501,N_13862);
nand UO_101 (O_101,N_14521,N_14252);
or UO_102 (O_102,N_13917,N_13877);
nor UO_103 (O_103,N_13861,N_13557);
and UO_104 (O_104,N_14025,N_14755);
nand UO_105 (O_105,N_14356,N_14824);
or UO_106 (O_106,N_14642,N_14423);
nand UO_107 (O_107,N_13568,N_13582);
or UO_108 (O_108,N_14241,N_14379);
and UO_109 (O_109,N_14631,N_14591);
and UO_110 (O_110,N_13801,N_13820);
or UO_111 (O_111,N_13951,N_14078);
or UO_112 (O_112,N_13729,N_13853);
nand UO_113 (O_113,N_14523,N_14159);
or UO_114 (O_114,N_14325,N_13993);
nand UO_115 (O_115,N_13955,N_14567);
xor UO_116 (O_116,N_14616,N_14719);
nand UO_117 (O_117,N_13502,N_14189);
or UO_118 (O_118,N_14908,N_14352);
xor UO_119 (O_119,N_14282,N_13588);
nor UO_120 (O_120,N_14170,N_13796);
nor UO_121 (O_121,N_14666,N_14209);
nand UO_122 (O_122,N_14909,N_14769);
or UO_123 (O_123,N_13868,N_13807);
nand UO_124 (O_124,N_14745,N_13595);
xor UO_125 (O_125,N_13556,N_14153);
nor UO_126 (O_126,N_14003,N_14327);
nor UO_127 (O_127,N_14381,N_13534);
xnor UO_128 (O_128,N_14578,N_14932);
and UO_129 (O_129,N_13701,N_14031);
nor UO_130 (O_130,N_13851,N_13676);
or UO_131 (O_131,N_14106,N_14525);
nor UO_132 (O_132,N_13982,N_14150);
or UO_133 (O_133,N_14154,N_13772);
xnor UO_134 (O_134,N_14351,N_13591);
nand UO_135 (O_135,N_14451,N_13808);
xor UO_136 (O_136,N_14284,N_13947);
nand UO_137 (O_137,N_13614,N_14223);
or UO_138 (O_138,N_13852,N_14826);
nor UO_139 (O_139,N_14815,N_14508);
nor UO_140 (O_140,N_14372,N_14941);
nor UO_141 (O_141,N_14579,N_14041);
and UO_142 (O_142,N_14303,N_13969);
nor UO_143 (O_143,N_14390,N_14149);
nor UO_144 (O_144,N_13708,N_14683);
or UO_145 (O_145,N_14102,N_13995);
or UO_146 (O_146,N_14608,N_14518);
nand UO_147 (O_147,N_14321,N_13699);
xor UO_148 (O_148,N_14050,N_14782);
nor UO_149 (O_149,N_13538,N_14336);
nor UO_150 (O_150,N_14361,N_14408);
nand UO_151 (O_151,N_13574,N_14990);
nand UO_152 (O_152,N_13914,N_14821);
and UO_153 (O_153,N_14979,N_13964);
and UO_154 (O_154,N_13896,N_14790);
nand UO_155 (O_155,N_13620,N_14514);
and UO_156 (O_156,N_13775,N_14935);
nor UO_157 (O_157,N_13745,N_14353);
or UO_158 (O_158,N_13604,N_14225);
and UO_159 (O_159,N_14511,N_14004);
nand UO_160 (O_160,N_13520,N_13797);
nand UO_161 (O_161,N_14950,N_13605);
nand UO_162 (O_162,N_14961,N_13965);
nand UO_163 (O_163,N_14449,N_14269);
and UO_164 (O_164,N_13882,N_13968);
nand UO_165 (O_165,N_14845,N_14298);
nor UO_166 (O_166,N_13984,N_13806);
xor UO_167 (O_167,N_13810,N_14853);
and UO_168 (O_168,N_13835,N_14022);
nor UO_169 (O_169,N_14090,N_13979);
xnor UO_170 (O_170,N_14249,N_14016);
nand UO_171 (O_171,N_13705,N_14085);
or UO_172 (O_172,N_14925,N_14574);
nor UO_173 (O_173,N_14322,N_13897);
nand UO_174 (O_174,N_13680,N_14027);
nor UO_175 (O_175,N_14076,N_14777);
nor UO_176 (O_176,N_13683,N_13733);
nor UO_177 (O_177,N_14210,N_14046);
nor UO_178 (O_178,N_14458,N_14146);
nor UO_179 (O_179,N_13726,N_14506);
nor UO_180 (O_180,N_13724,N_14479);
and UO_181 (O_181,N_14759,N_14801);
nor UO_182 (O_182,N_13908,N_14748);
and UO_183 (O_183,N_13789,N_14185);
nor UO_184 (O_184,N_13512,N_14702);
nand UO_185 (O_185,N_14483,N_14461);
or UO_186 (O_186,N_13837,N_13936);
nor UO_187 (O_187,N_13514,N_14463);
or UO_188 (O_188,N_14898,N_14221);
nand UO_189 (O_189,N_14288,N_14689);
or UO_190 (O_190,N_14799,N_13528);
or UO_191 (O_191,N_13609,N_14477);
and UO_192 (O_192,N_13679,N_14945);
nor UO_193 (O_193,N_14348,N_14862);
nand UO_194 (O_194,N_14732,N_14727);
and UO_195 (O_195,N_14329,N_13501);
nand UO_196 (O_196,N_14171,N_13698);
nand UO_197 (O_197,N_14293,N_14678);
or UO_198 (O_198,N_14273,N_13695);
nor UO_199 (O_199,N_14015,N_14615);
nand UO_200 (O_200,N_13718,N_14215);
or UO_201 (O_201,N_14009,N_13794);
nor UO_202 (O_202,N_13983,N_14315);
nor UO_203 (O_203,N_14365,N_14392);
or UO_204 (O_204,N_14393,N_13823);
nor UO_205 (O_205,N_14758,N_14306);
nor UO_206 (O_206,N_13838,N_14543);
or UO_207 (O_207,N_13883,N_14786);
or UO_208 (O_208,N_13812,N_14061);
or UO_209 (O_209,N_14331,N_14664);
nor UO_210 (O_210,N_13715,N_14829);
or UO_211 (O_211,N_14167,N_14946);
and UO_212 (O_212,N_14264,N_14680);
or UO_213 (O_213,N_13874,N_13921);
nor UO_214 (O_214,N_14922,N_14074);
nor UO_215 (O_215,N_14770,N_13576);
and UO_216 (O_216,N_14378,N_14333);
nor UO_217 (O_217,N_13859,N_14627);
or UO_218 (O_218,N_14305,N_14317);
xor UO_219 (O_219,N_13976,N_14455);
nand UO_220 (O_220,N_14005,N_14836);
and UO_221 (O_221,N_14060,N_13518);
or UO_222 (O_222,N_13544,N_14165);
nand UO_223 (O_223,N_13959,N_14573);
nor UO_224 (O_224,N_14783,N_13630);
nand UO_225 (O_225,N_14101,N_14930);
nand UO_226 (O_226,N_13957,N_13910);
nand UO_227 (O_227,N_14988,N_14776);
xnor UO_228 (O_228,N_13833,N_13543);
xnor UO_229 (O_229,N_13722,N_14117);
nor UO_230 (O_230,N_14552,N_13997);
and UO_231 (O_231,N_13811,N_13622);
and UO_232 (O_232,N_13546,N_13567);
nand UO_233 (O_233,N_13803,N_13783);
or UO_234 (O_234,N_14540,N_14848);
xor UO_235 (O_235,N_14822,N_14291);
and UO_236 (O_236,N_13788,N_14595);
nor UO_237 (O_237,N_14529,N_13559);
nand UO_238 (O_238,N_13703,N_14869);
nor UO_239 (O_239,N_14539,N_13629);
or UO_240 (O_240,N_13948,N_14958);
nand UO_241 (O_241,N_13623,N_14274);
and UO_242 (O_242,N_14984,N_14896);
nand UO_243 (O_243,N_13597,N_13858);
or UO_244 (O_244,N_14384,N_13782);
and UO_245 (O_245,N_14203,N_13749);
nand UO_246 (O_246,N_14105,N_14975);
nor UO_247 (O_247,N_14992,N_13880);
xnor UO_248 (O_248,N_14837,N_14360);
nand UO_249 (O_249,N_14536,N_14554);
and UO_250 (O_250,N_13545,N_14730);
nor UO_251 (O_251,N_14229,N_13717);
and UO_252 (O_252,N_14111,N_14442);
or UO_253 (O_253,N_14596,N_14272);
xor UO_254 (O_254,N_14987,N_14688);
or UO_255 (O_255,N_14326,N_14187);
nand UO_256 (O_256,N_14524,N_13561);
nand UO_257 (O_257,N_14802,N_13755);
nor UO_258 (O_258,N_14919,N_14609);
nor UO_259 (O_259,N_13674,N_14956);
and UO_260 (O_260,N_14414,N_14805);
nand UO_261 (O_261,N_14647,N_14726);
or UO_262 (O_262,N_14420,N_14537);
nand UO_263 (O_263,N_14827,N_14340);
nor UO_264 (O_264,N_13953,N_14771);
and UO_265 (O_265,N_14307,N_14387);
and UO_266 (O_266,N_14335,N_13890);
nor UO_267 (O_267,N_14838,N_14472);
nand UO_268 (O_268,N_13774,N_14849);
nor UO_269 (O_269,N_14359,N_14547);
or UO_270 (O_270,N_14014,N_13934);
nor UO_271 (O_271,N_14964,N_14338);
and UO_272 (O_272,N_13684,N_14347);
or UO_273 (O_273,N_14169,N_14575);
nand UO_274 (O_274,N_14118,N_14309);
nand UO_275 (O_275,N_13909,N_14986);
nand UO_276 (O_276,N_14422,N_13681);
nand UO_277 (O_277,N_13894,N_14488);
and UO_278 (O_278,N_14138,N_13641);
nor UO_279 (O_279,N_14174,N_13670);
nand UO_280 (O_280,N_14095,N_13624);
and UO_281 (O_281,N_13777,N_14897);
nor UO_282 (O_282,N_13665,N_13954);
nand UO_283 (O_283,N_14092,N_14088);
nor UO_284 (O_284,N_14280,N_14940);
nor UO_285 (O_285,N_14747,N_13667);
nor UO_286 (O_286,N_14966,N_14551);
nand UO_287 (O_287,N_14713,N_14067);
xor UO_288 (O_288,N_14486,N_14868);
nand UO_289 (O_289,N_14978,N_14495);
and UO_290 (O_290,N_13860,N_14254);
and UO_291 (O_291,N_14522,N_13815);
and UO_292 (O_292,N_13564,N_13817);
nor UO_293 (O_293,N_14646,N_13792);
nand UO_294 (O_294,N_13902,N_14895);
nor UO_295 (O_295,N_13617,N_13607);
nor UO_296 (O_296,N_14789,N_14195);
xnor UO_297 (O_297,N_14339,N_14723);
or UO_298 (O_298,N_13760,N_14023);
nand UO_299 (O_299,N_14639,N_14226);
nor UO_300 (O_300,N_14676,N_14391);
nor UO_301 (O_301,N_14120,N_13907);
nor UO_302 (O_302,N_14228,N_14768);
and UO_303 (O_303,N_14910,N_14235);
nand UO_304 (O_304,N_14000,N_14700);
and UO_305 (O_305,N_14672,N_14456);
and UO_306 (O_306,N_13887,N_14130);
and UO_307 (O_307,N_14873,N_14892);
and UO_308 (O_308,N_14820,N_13643);
or UO_309 (O_309,N_14913,N_14510);
or UO_310 (O_310,N_14468,N_14640);
and UO_311 (O_311,N_14911,N_14841);
and UO_312 (O_312,N_14754,N_14490);
nand UO_313 (O_313,N_14548,N_14103);
and UO_314 (O_314,N_14860,N_14373);
or UO_315 (O_315,N_14752,N_13704);
nor UO_316 (O_316,N_14981,N_13922);
and UO_317 (O_317,N_13945,N_14823);
or UO_318 (O_318,N_14962,N_14204);
and UO_319 (O_319,N_14580,N_13799);
or UO_320 (O_320,N_14762,N_14236);
and UO_321 (O_321,N_13873,N_14643);
xnor UO_322 (O_322,N_14670,N_14475);
nand UO_323 (O_323,N_14035,N_14262);
or UO_324 (O_324,N_13687,N_14891);
and UO_325 (O_325,N_14781,N_14127);
nor UO_326 (O_326,N_13986,N_14875);
xnor UO_327 (O_327,N_13834,N_14894);
or UO_328 (O_328,N_13584,N_14545);
xnor UO_329 (O_329,N_14613,N_13553);
nor UO_330 (O_330,N_14857,N_14943);
nor UO_331 (O_331,N_14734,N_14415);
or UO_332 (O_332,N_14342,N_14629);
nand UO_333 (O_333,N_13677,N_13736);
nand UO_334 (O_334,N_13762,N_14257);
nand UO_335 (O_335,N_14780,N_14083);
nand UO_336 (O_336,N_13875,N_14316);
nand UO_337 (O_337,N_13693,N_13872);
nand UO_338 (O_338,N_14132,N_14809);
xnor UO_339 (O_339,N_13891,N_14725);
or UO_340 (O_340,N_14655,N_14872);
and UO_341 (O_341,N_14560,N_14626);
nor UO_342 (O_342,N_14208,N_14660);
and UO_343 (O_343,N_13734,N_13972);
nand UO_344 (O_344,N_14998,N_13657);
nand UO_345 (O_345,N_14556,N_14354);
and UO_346 (O_346,N_14370,N_14912);
nand UO_347 (O_347,N_14811,N_14893);
and UO_348 (O_348,N_14281,N_13541);
or UO_349 (O_349,N_13529,N_14502);
nand UO_350 (O_350,N_14753,N_13949);
nand UO_351 (O_351,N_13594,N_14544);
or UO_352 (O_352,N_13800,N_14564);
nor UO_353 (O_353,N_13650,N_14681);
nor UO_354 (O_354,N_13513,N_14830);
xnor UO_355 (O_355,N_14054,N_14007);
and UO_356 (O_356,N_13721,N_14546);
and UO_357 (O_357,N_13600,N_13754);
and UO_358 (O_358,N_14534,N_13805);
or UO_359 (O_359,N_14160,N_14299);
nor UO_360 (O_360,N_14620,N_14864);
or UO_361 (O_361,N_13827,N_14143);
and UO_362 (O_362,N_14363,N_14168);
and UO_363 (O_363,N_14124,N_13539);
and UO_364 (O_364,N_13626,N_14377);
and UO_365 (O_365,N_13731,N_13678);
nor UO_366 (O_366,N_14368,N_14601);
or UO_367 (O_367,N_14399,N_14973);
or UO_368 (O_368,N_14375,N_14561);
and UO_369 (O_369,N_14576,N_14312);
xor UO_370 (O_370,N_14260,N_14188);
nor UO_371 (O_371,N_13870,N_14970);
nor UO_372 (O_372,N_14641,N_13532);
xor UO_373 (O_373,N_14289,N_14855);
nor UO_374 (O_374,N_14634,N_14870);
or UO_375 (O_375,N_14211,N_14213);
and UO_376 (O_376,N_14694,N_14996);
nand UO_377 (O_377,N_14571,N_14833);
nand UO_378 (O_378,N_13885,N_13589);
nor UO_379 (O_379,N_14707,N_13929);
and UO_380 (O_380,N_13510,N_13732);
xor UO_381 (O_381,N_14675,N_14419);
nor UO_382 (O_382,N_14942,N_14566);
nor UO_383 (O_383,N_14152,N_13649);
nor UO_384 (O_384,N_14186,N_13990);
nand UO_385 (O_385,N_14276,N_14902);
xor UO_386 (O_386,N_14901,N_13523);
and UO_387 (O_387,N_14109,N_14760);
xnor UO_388 (O_388,N_14012,N_13973);
nand UO_389 (O_389,N_14265,N_14819);
xnor UO_390 (O_390,N_14982,N_13577);
and UO_391 (O_391,N_13744,N_14343);
nand UO_392 (O_392,N_14491,N_14598);
nand UO_393 (O_393,N_14267,N_14045);
and UO_394 (O_394,N_14021,N_13593);
and UO_395 (O_395,N_13844,N_14767);
and UO_396 (O_396,N_13992,N_14011);
or UO_397 (O_397,N_14583,N_14497);
or UO_398 (O_398,N_14019,N_14320);
and UO_399 (O_399,N_14155,N_14948);
and UO_400 (O_400,N_14917,N_13780);
xor UO_401 (O_401,N_14397,N_14428);
or UO_402 (O_402,N_14557,N_13713);
nand UO_403 (O_403,N_14158,N_13842);
nor UO_404 (O_404,N_14916,N_14141);
nor UO_405 (O_405,N_13530,N_14711);
and UO_406 (O_406,N_13634,N_13849);
nor UO_407 (O_407,N_13850,N_13527);
or UO_408 (O_408,N_14594,N_13765);
nor UO_409 (O_409,N_14905,N_14877);
nand UO_410 (O_410,N_14114,N_13666);
or UO_411 (O_411,N_14454,N_14503);
nor UO_412 (O_412,N_13672,N_13958);
nor UO_413 (O_413,N_13864,N_14409);
nor UO_414 (O_414,N_14296,N_13793);
nor UO_415 (O_415,N_14075,N_14328);
and UO_416 (O_416,N_14947,N_14048);
and UO_417 (O_417,N_14796,N_14586);
or UO_418 (O_418,N_14427,N_13950);
nand UO_419 (O_419,N_13506,N_13540);
nand UO_420 (O_420,N_14509,N_14417);
and UO_421 (O_421,N_13824,N_14512);
nor UO_422 (O_422,N_14904,N_14787);
nand UO_423 (O_423,N_14955,N_13654);
or UO_424 (O_424,N_14433,N_13504);
and UO_425 (O_425,N_14485,N_14851);
nand UO_426 (O_426,N_13987,N_14997);
nor UO_427 (O_427,N_14400,N_14073);
or UO_428 (O_428,N_14098,N_14038);
or UO_429 (O_429,N_14398,N_14216);
nand UO_430 (O_430,N_13549,N_14746);
xor UO_431 (O_431,N_14969,N_13618);
xnor UO_432 (O_432,N_13615,N_14121);
nand UO_433 (O_433,N_14582,N_13848);
or UO_434 (O_434,N_13524,N_14430);
nand UO_435 (O_435,N_13889,N_14049);
nor UO_436 (O_436,N_14765,N_14234);
or UO_437 (O_437,N_13943,N_14581);
nor UO_438 (O_438,N_13669,N_14763);
nor UO_439 (O_439,N_13911,N_14425);
nand UO_440 (O_440,N_14344,N_14460);
or UO_441 (O_441,N_14622,N_13728);
nor UO_442 (O_442,N_14062,N_14029);
or UO_443 (O_443,N_13551,N_14178);
or UO_444 (O_444,N_14562,N_14100);
or UO_445 (O_445,N_14716,N_14549);
nand UO_446 (O_446,N_13994,N_14385);
or UO_447 (O_447,N_14938,N_13688);
or UO_448 (O_448,N_14065,N_14219);
nand UO_449 (O_449,N_14535,N_14624);
or UO_450 (O_450,N_14126,N_14248);
xnor UO_451 (O_451,N_14699,N_14283);
nand UO_452 (O_452,N_14816,N_14800);
nor UO_453 (O_453,N_14954,N_14565);
or UO_454 (O_454,N_14122,N_14710);
or UO_455 (O_455,N_13522,N_14093);
or UO_456 (O_456,N_14825,N_14018);
nand UO_457 (O_457,N_14131,N_14297);
nor UO_458 (O_458,N_13961,N_13719);
nor UO_459 (O_459,N_14403,N_14314);
nor UO_460 (O_460,N_13686,N_14779);
nor UO_461 (O_461,N_13795,N_13583);
nor UO_462 (O_462,N_14323,N_13580);
nand UO_463 (O_463,N_13764,N_13931);
nand UO_464 (O_464,N_13596,N_14224);
nand UO_465 (O_465,N_13871,N_14220);
or UO_466 (O_466,N_13579,N_13977);
and UO_467 (O_467,N_13933,N_13602);
and UO_468 (O_468,N_14418,N_14637);
xnor UO_469 (O_469,N_14531,N_14402);
and UO_470 (O_470,N_13786,N_13587);
nor UO_471 (O_471,N_14028,N_14890);
nor UO_472 (O_472,N_14903,N_14271);
nor UO_473 (O_473,N_13516,N_13779);
and UO_474 (O_474,N_14863,N_14587);
and UO_475 (O_475,N_13747,N_14704);
nor UO_476 (O_476,N_14071,N_14493);
nor UO_477 (O_477,N_14589,N_14010);
and UO_478 (O_478,N_13572,N_13770);
xor UO_479 (O_479,N_14024,N_14302);
nand UO_480 (O_480,N_14474,N_14412);
xor UO_481 (O_481,N_14112,N_14135);
xor UO_482 (O_482,N_14349,N_14051);
nor UO_483 (O_483,N_13613,N_14775);
nand UO_484 (O_484,N_14404,N_13846);
xnor UO_485 (O_485,N_13926,N_14741);
and UO_486 (O_486,N_14985,N_13610);
nor UO_487 (O_487,N_14794,N_13939);
and UO_488 (O_488,N_14737,N_13716);
or UO_489 (O_489,N_14729,N_13750);
xor UO_490 (O_490,N_13865,N_14184);
nand UO_491 (O_491,N_14846,N_13571);
nor UO_492 (O_492,N_14362,N_13825);
or UO_493 (O_493,N_14268,N_14553);
and UO_494 (O_494,N_13507,N_14270);
nor UO_495 (O_495,N_13645,N_13863);
nand UO_496 (O_496,N_14134,N_13898);
nor UO_497 (O_497,N_13691,N_14087);
nor UO_498 (O_498,N_14173,N_14395);
nand UO_499 (O_499,N_13533,N_14738);
and UO_500 (O_500,N_14610,N_13508);
and UO_501 (O_501,N_14791,N_14069);
nor UO_502 (O_502,N_14648,N_13740);
nor UO_503 (O_503,N_14081,N_14232);
nand UO_504 (O_504,N_14971,N_14239);
and UO_505 (O_505,N_13798,N_14405);
xor UO_506 (O_506,N_13900,N_14137);
nor UO_507 (O_507,N_14888,N_14332);
or UO_508 (O_508,N_13970,N_13590);
nor UO_509 (O_509,N_14937,N_14570);
and UO_510 (O_510,N_14357,N_14706);
nor UO_511 (O_511,N_14697,N_13659);
or UO_512 (O_512,N_13552,N_14350);
or UO_513 (O_513,N_14500,N_14113);
nor UO_514 (O_514,N_14907,N_14528);
xor UO_515 (O_515,N_13816,N_14341);
nand UO_516 (O_516,N_13500,N_14147);
or UO_517 (O_517,N_14926,N_13720);
xor UO_518 (O_518,N_14369,N_13662);
and UO_519 (O_519,N_13636,N_14084);
and UO_520 (O_520,N_14717,N_13565);
xnor UO_521 (O_521,N_13841,N_14222);
nand UO_522 (O_522,N_14123,N_13867);
nand UO_523 (O_523,N_14396,N_14597);
and UO_524 (O_524,N_13826,N_14728);
and UO_525 (O_525,N_14757,N_14834);
nor UO_526 (O_526,N_14207,N_14182);
nand UO_527 (O_527,N_13742,N_13924);
nor UO_528 (O_528,N_14682,N_14761);
nand UO_529 (O_529,N_13696,N_14161);
xor UO_530 (O_530,N_13857,N_14921);
xor UO_531 (O_531,N_14237,N_14218);
or UO_532 (O_532,N_13905,N_14447);
nand UO_533 (O_533,N_14792,N_14630);
or UO_534 (O_534,N_14108,N_14496);
nand UO_535 (O_535,N_14733,N_14977);
nor UO_536 (O_536,N_14036,N_13996);
and UO_537 (O_537,N_14559,N_13621);
nand UO_538 (O_538,N_14967,N_14355);
nand UO_539 (O_539,N_14803,N_13912);
nand UO_540 (O_540,N_13606,N_14136);
nand UO_541 (O_541,N_14883,N_13836);
nand UO_542 (O_542,N_14931,N_14847);
nor UO_543 (O_543,N_14330,N_13738);
nand UO_544 (O_544,N_14951,N_14842);
nand UO_545 (O_545,N_14040,N_14079);
and UO_546 (O_546,N_14957,N_14243);
nor UO_547 (O_547,N_14450,N_14915);
nand UO_548 (O_548,N_14778,N_14489);
xor UO_549 (O_549,N_14685,N_13575);
and UO_550 (O_550,N_13661,N_14538);
or UO_551 (O_551,N_13638,N_14690);
and UO_552 (O_552,N_13692,N_14166);
nor UO_553 (O_553,N_14259,N_14089);
and UO_554 (O_554,N_13639,N_13637);
nor UO_555 (O_555,N_14963,N_13980);
nor UO_556 (O_556,N_14959,N_13767);
and UO_557 (O_557,N_14818,N_14623);
and UO_558 (O_558,N_14424,N_13998);
or UO_559 (O_559,N_14513,N_14797);
nand UO_560 (O_560,N_13821,N_14295);
nand UO_561 (O_561,N_14197,N_13847);
nand UO_562 (O_562,N_14920,N_14656);
nor UO_563 (O_563,N_13904,N_14605);
and UO_564 (O_564,N_14217,N_14068);
or UO_565 (O_565,N_14588,N_14032);
and UO_566 (O_566,N_14645,N_14310);
nand UO_567 (O_567,N_14091,N_14774);
xnor UO_568 (O_568,N_13525,N_14722);
or UO_569 (O_569,N_14691,N_14070);
nor UO_570 (O_570,N_13668,N_14568);
and UO_571 (O_571,N_14654,N_14673);
nor UO_572 (O_572,N_14906,N_14258);
or UO_573 (O_573,N_14133,N_14692);
or UO_574 (O_574,N_14619,N_14324);
nor UO_575 (O_575,N_14452,N_14441);
and UO_576 (O_576,N_14667,N_14480);
and UO_577 (O_577,N_14650,N_14077);
nand UO_578 (O_578,N_13752,N_14438);
xor UO_579 (O_579,N_14671,N_14157);
or UO_580 (O_580,N_14426,N_14006);
nand UO_581 (O_581,N_13644,N_13822);
nor UO_582 (O_582,N_13656,N_14530);
or UO_583 (O_583,N_13978,N_13581);
and UO_584 (O_584,N_14611,N_13769);
or UO_585 (O_585,N_14487,N_13930);
nor UO_586 (O_586,N_14467,N_13700);
and UO_587 (O_587,N_14072,N_14918);
nor UO_588 (O_588,N_14621,N_14482);
nor UO_589 (O_589,N_14346,N_14162);
nor UO_590 (O_590,N_14047,N_14677);
and UO_591 (O_591,N_13913,N_14934);
nor UO_592 (O_592,N_13673,N_14172);
nor UO_593 (O_593,N_14810,N_13612);
or UO_594 (O_594,N_13915,N_14364);
or UO_595 (O_595,N_13702,N_14205);
nand UO_596 (O_596,N_14465,N_14437);
xnor UO_597 (O_597,N_13818,N_13632);
xor UO_598 (O_598,N_14498,N_14718);
nand UO_599 (O_599,N_14944,N_14519);
nor UO_600 (O_600,N_13967,N_14861);
or UO_601 (O_601,N_13570,N_14614);
and UO_602 (O_602,N_14832,N_14156);
nor UO_603 (O_603,N_13723,N_14401);
nand UO_604 (O_604,N_13804,N_14740);
nor UO_605 (O_605,N_14687,N_14798);
or UO_606 (O_606,N_14878,N_14749);
nand UO_607 (O_607,N_14665,N_13711);
nor UO_608 (O_608,N_14933,N_13855);
or UO_609 (O_609,N_13757,N_13558);
or UO_610 (O_610,N_13664,N_14835);
and UO_611 (O_611,N_14416,N_13940);
nand UO_612 (O_612,N_13542,N_14148);
xnor UO_613 (O_613,N_14082,N_14504);
or UO_614 (O_614,N_13694,N_13547);
nor UO_615 (O_615,N_14785,N_13675);
or UO_616 (O_616,N_14812,N_13866);
or UO_617 (O_617,N_13840,N_13631);
or UO_618 (O_618,N_14806,N_14231);
nor UO_619 (O_619,N_13785,N_14086);
nand UO_620 (O_620,N_14277,N_14953);
or UO_621 (O_621,N_14446,N_13690);
nand UO_622 (O_622,N_14478,N_14334);
nor UO_623 (O_623,N_14854,N_14541);
or UO_624 (O_624,N_14628,N_14201);
nand UO_625 (O_625,N_14644,N_13598);
nand UO_626 (O_626,N_14444,N_14080);
and UO_627 (O_627,N_14876,N_14867);
or UO_628 (O_628,N_13535,N_14176);
nor UO_629 (O_629,N_14772,N_14026);
nand UO_630 (O_630,N_13946,N_14844);
nand UO_631 (O_631,N_13761,N_14744);
nor UO_632 (O_632,N_14448,N_14163);
xor UO_633 (O_633,N_13601,N_14939);
or UO_634 (O_634,N_14739,N_14577);
nand UO_635 (O_635,N_13956,N_13759);
xnor UO_636 (O_636,N_14515,N_14034);
and UO_637 (O_637,N_14555,N_14828);
nor UO_638 (O_638,N_14337,N_14880);
and UO_639 (O_639,N_14592,N_13743);
or UO_640 (O_640,N_14013,N_14440);
nor UO_641 (O_641,N_14097,N_14686);
or UO_642 (O_642,N_14999,N_13658);
and UO_643 (O_643,N_14612,N_14731);
xnor UO_644 (O_644,N_14751,N_14572);
xnor UO_645 (O_645,N_13960,N_13519);
and UO_646 (O_646,N_14439,N_14238);
and UO_647 (O_647,N_14191,N_14001);
and UO_648 (O_648,N_14674,N_14991);
nand UO_649 (O_649,N_14301,N_13845);
nor UO_650 (O_650,N_13942,N_14517);
xor UO_651 (O_651,N_14473,N_14053);
nor UO_652 (O_652,N_14550,N_14764);
and UO_653 (O_653,N_14874,N_13712);
or UO_654 (O_654,N_14858,N_14657);
nor UO_655 (O_655,N_14308,N_14850);
nor UO_656 (O_656,N_13888,N_14507);
and UO_657 (O_657,N_14843,N_14183);
or UO_658 (O_658,N_14859,N_14285);
and UO_659 (O_659,N_13938,N_14096);
or UO_660 (O_660,N_13778,N_14388);
or UO_661 (O_661,N_14899,N_13714);
or UO_662 (O_662,N_14766,N_13706);
nor UO_663 (O_663,N_14371,N_14290);
nand UO_664 (O_664,N_13730,N_13790);
and UO_665 (O_665,N_14128,N_14196);
and UO_666 (O_666,N_13628,N_14684);
or UO_667 (O_667,N_13509,N_14058);
nor UO_668 (O_668,N_14952,N_13569);
nor UO_669 (O_669,N_14720,N_13640);
and UO_670 (O_670,N_14052,N_14661);
and UO_671 (O_671,N_14593,N_14374);
or UO_672 (O_672,N_13685,N_14735);
nor UO_673 (O_673,N_13999,N_14278);
nand UO_674 (O_674,N_13766,N_14469);
nand UO_675 (O_675,N_14287,N_13526);
xnor UO_676 (O_676,N_13802,N_14993);
and UO_677 (O_677,N_13648,N_14900);
and UO_678 (O_678,N_14724,N_13881);
or UO_679 (O_679,N_13787,N_13854);
nor UO_680 (O_680,N_14994,N_14516);
or UO_681 (O_681,N_14366,N_14063);
and UO_682 (O_682,N_13916,N_13550);
nand UO_683 (O_683,N_13932,N_14750);
xor UO_684 (O_684,N_13521,N_14839);
nand UO_685 (O_685,N_14632,N_14633);
nand UO_686 (O_686,N_14695,N_14889);
nand UO_687 (O_687,N_13988,N_14949);
and UO_688 (O_688,N_14367,N_14708);
nand UO_689 (O_689,N_14585,N_14807);
nor UO_690 (O_690,N_14110,N_14793);
and UO_691 (O_691,N_14756,N_14017);
xor UO_692 (O_692,N_14443,N_14668);
xnor UO_693 (O_693,N_14057,N_14499);
nand UO_694 (O_694,N_14584,N_13660);
and UO_695 (O_695,N_14882,N_14181);
nor UO_696 (O_696,N_14831,N_14693);
nor UO_697 (O_697,N_14192,N_13884);
nor UO_698 (O_698,N_13741,N_14410);
nand UO_699 (O_699,N_14709,N_13517);
and UO_700 (O_700,N_13554,N_13646);
nor UO_701 (O_701,N_13819,N_14604);
or UO_702 (O_702,N_13920,N_13603);
or UO_703 (O_703,N_14194,N_13895);
and UO_704 (O_704,N_13901,N_14436);
and UO_705 (O_705,N_13682,N_13737);
and UO_706 (O_706,N_14995,N_14965);
xor UO_707 (O_707,N_14431,N_14881);
nor UO_708 (O_708,N_14142,N_14635);
nor UO_709 (O_709,N_14445,N_13935);
nand UO_710 (O_710,N_13892,N_13651);
and UO_711 (O_711,N_13830,N_14679);
nand UO_712 (O_712,N_14435,N_13893);
and UO_713 (O_713,N_14980,N_13710);
and UO_714 (O_714,N_14044,N_14464);
nand UO_715 (O_715,N_13781,N_13611);
and UO_716 (O_716,N_14698,N_14140);
nand UO_717 (O_717,N_13725,N_14198);
nor UO_718 (O_718,N_14311,N_13748);
and UO_719 (O_719,N_13619,N_14887);
nand UO_720 (O_720,N_13791,N_14002);
nand UO_721 (O_721,N_14885,N_13886);
nand UO_722 (O_722,N_14253,N_13756);
or UO_723 (O_723,N_14742,N_13937);
or UO_724 (O_724,N_14286,N_14227);
and UO_725 (O_725,N_13515,N_14960);
and UO_726 (O_726,N_14520,N_14434);
and UO_727 (O_727,N_14200,N_14066);
or UO_728 (O_728,N_14250,N_14151);
and UO_729 (O_729,N_14505,N_14871);
or UO_730 (O_730,N_14212,N_14386);
nand UO_731 (O_731,N_13963,N_13548);
and UO_732 (O_732,N_14345,N_14206);
nor UO_733 (O_733,N_14852,N_14376);
and UO_734 (O_734,N_14603,N_14602);
and UO_735 (O_735,N_13671,N_13831);
and UO_736 (O_736,N_13735,N_13758);
nor UO_737 (O_737,N_13768,N_14042);
nand UO_738 (O_738,N_13635,N_14145);
xor UO_739 (O_739,N_14884,N_13709);
nor UO_740 (O_740,N_13751,N_14886);
or UO_741 (O_741,N_13689,N_13809);
and UO_742 (O_742,N_14606,N_14457);
nor UO_743 (O_743,N_14701,N_14179);
and UO_744 (O_744,N_14056,N_14976);
or UO_745 (O_745,N_14736,N_13784);
xor UO_746 (O_746,N_14144,N_14773);
nand UO_747 (O_747,N_13771,N_13592);
xnor UO_748 (O_748,N_14669,N_14266);
nor UO_749 (O_749,N_14300,N_13952);
nor UO_750 (O_750,N_14043,N_14160);
xnor UO_751 (O_751,N_14116,N_13786);
nand UO_752 (O_752,N_14561,N_13799);
xor UO_753 (O_753,N_14845,N_14703);
or UO_754 (O_754,N_13984,N_14615);
and UO_755 (O_755,N_14634,N_14540);
nor UO_756 (O_756,N_14494,N_14255);
or UO_757 (O_757,N_14521,N_13896);
or UO_758 (O_758,N_14352,N_14864);
and UO_759 (O_759,N_14771,N_13546);
and UO_760 (O_760,N_13538,N_14289);
or UO_761 (O_761,N_13573,N_14163);
nand UO_762 (O_762,N_13846,N_14766);
and UO_763 (O_763,N_14212,N_14582);
nor UO_764 (O_764,N_14361,N_14446);
and UO_765 (O_765,N_14524,N_14873);
and UO_766 (O_766,N_13733,N_14757);
nor UO_767 (O_767,N_14618,N_14600);
nand UO_768 (O_768,N_14549,N_14292);
nand UO_769 (O_769,N_14558,N_13758);
and UO_770 (O_770,N_13573,N_14985);
nand UO_771 (O_771,N_14017,N_14703);
or UO_772 (O_772,N_14206,N_14895);
or UO_773 (O_773,N_13652,N_14234);
and UO_774 (O_774,N_14197,N_13886);
xor UO_775 (O_775,N_14527,N_13901);
and UO_776 (O_776,N_13672,N_13802);
or UO_777 (O_777,N_14015,N_14569);
or UO_778 (O_778,N_14264,N_13589);
or UO_779 (O_779,N_14743,N_14577);
or UO_780 (O_780,N_13943,N_13609);
nand UO_781 (O_781,N_13899,N_14594);
nand UO_782 (O_782,N_14790,N_13892);
nor UO_783 (O_783,N_13553,N_14173);
or UO_784 (O_784,N_14467,N_14178);
nor UO_785 (O_785,N_13555,N_14023);
xor UO_786 (O_786,N_14206,N_14587);
nand UO_787 (O_787,N_14292,N_14017);
and UO_788 (O_788,N_14584,N_13712);
nor UO_789 (O_789,N_14281,N_13760);
nor UO_790 (O_790,N_13752,N_14611);
and UO_791 (O_791,N_13595,N_14506);
and UO_792 (O_792,N_14743,N_13578);
nor UO_793 (O_793,N_14310,N_14409);
and UO_794 (O_794,N_14634,N_13567);
and UO_795 (O_795,N_14248,N_14558);
xnor UO_796 (O_796,N_14306,N_14572);
xor UO_797 (O_797,N_14208,N_13571);
nand UO_798 (O_798,N_14376,N_14583);
and UO_799 (O_799,N_14116,N_14384);
xor UO_800 (O_800,N_13766,N_14690);
nor UO_801 (O_801,N_14245,N_14341);
nor UO_802 (O_802,N_14080,N_13998);
or UO_803 (O_803,N_13642,N_14978);
nor UO_804 (O_804,N_14353,N_14393);
and UO_805 (O_805,N_13649,N_13532);
nor UO_806 (O_806,N_13656,N_13628);
nand UO_807 (O_807,N_14392,N_14132);
and UO_808 (O_808,N_14545,N_14772);
or UO_809 (O_809,N_14463,N_14834);
and UO_810 (O_810,N_14312,N_14622);
nor UO_811 (O_811,N_13839,N_14529);
nor UO_812 (O_812,N_13852,N_13770);
and UO_813 (O_813,N_13906,N_13787);
nor UO_814 (O_814,N_13545,N_14681);
xor UO_815 (O_815,N_14444,N_14638);
nor UO_816 (O_816,N_14111,N_14876);
nand UO_817 (O_817,N_13813,N_13556);
nor UO_818 (O_818,N_13815,N_14368);
and UO_819 (O_819,N_14461,N_14828);
or UO_820 (O_820,N_14790,N_14630);
nand UO_821 (O_821,N_14420,N_13758);
nor UO_822 (O_822,N_14398,N_13607);
or UO_823 (O_823,N_14118,N_14816);
xor UO_824 (O_824,N_14356,N_13527);
nand UO_825 (O_825,N_14602,N_14662);
nand UO_826 (O_826,N_14175,N_13585);
nor UO_827 (O_827,N_13806,N_14544);
and UO_828 (O_828,N_14191,N_13879);
or UO_829 (O_829,N_14055,N_13668);
or UO_830 (O_830,N_14439,N_14214);
or UO_831 (O_831,N_14787,N_14713);
xnor UO_832 (O_832,N_14115,N_14504);
nand UO_833 (O_833,N_14908,N_14650);
nand UO_834 (O_834,N_14863,N_14324);
and UO_835 (O_835,N_14762,N_14942);
or UO_836 (O_836,N_14427,N_14169);
nand UO_837 (O_837,N_13659,N_14190);
nor UO_838 (O_838,N_13800,N_14195);
xor UO_839 (O_839,N_14193,N_13776);
xnor UO_840 (O_840,N_13797,N_14289);
or UO_841 (O_841,N_13878,N_14486);
nand UO_842 (O_842,N_14484,N_14003);
or UO_843 (O_843,N_14045,N_14041);
nand UO_844 (O_844,N_13605,N_14026);
nand UO_845 (O_845,N_14950,N_14339);
nor UO_846 (O_846,N_13900,N_14096);
nor UO_847 (O_847,N_14589,N_14634);
nor UO_848 (O_848,N_14522,N_14222);
or UO_849 (O_849,N_13520,N_13807);
or UO_850 (O_850,N_14493,N_14922);
or UO_851 (O_851,N_13873,N_14536);
nor UO_852 (O_852,N_14841,N_14595);
xor UO_853 (O_853,N_13833,N_14617);
and UO_854 (O_854,N_14671,N_14866);
nor UO_855 (O_855,N_14493,N_14408);
or UO_856 (O_856,N_14411,N_14851);
and UO_857 (O_857,N_14500,N_14695);
nor UO_858 (O_858,N_14842,N_14105);
or UO_859 (O_859,N_14522,N_13555);
xnor UO_860 (O_860,N_14296,N_14201);
or UO_861 (O_861,N_14825,N_14004);
xnor UO_862 (O_862,N_14427,N_13643);
nand UO_863 (O_863,N_14620,N_14639);
and UO_864 (O_864,N_14733,N_14743);
and UO_865 (O_865,N_14430,N_14896);
and UO_866 (O_866,N_14276,N_14636);
or UO_867 (O_867,N_14938,N_14698);
or UO_868 (O_868,N_14299,N_14618);
or UO_869 (O_869,N_14004,N_14590);
and UO_870 (O_870,N_13654,N_14303);
nand UO_871 (O_871,N_13975,N_14457);
or UO_872 (O_872,N_13813,N_14691);
nand UO_873 (O_873,N_14217,N_14370);
or UO_874 (O_874,N_14350,N_14462);
and UO_875 (O_875,N_14842,N_14183);
nand UO_876 (O_876,N_13998,N_13745);
or UO_877 (O_877,N_14445,N_13832);
nor UO_878 (O_878,N_14422,N_14541);
or UO_879 (O_879,N_14112,N_14013);
nand UO_880 (O_880,N_14913,N_14020);
and UO_881 (O_881,N_13731,N_14184);
nor UO_882 (O_882,N_14818,N_14840);
xor UO_883 (O_883,N_13783,N_13527);
nor UO_884 (O_884,N_13501,N_14201);
nand UO_885 (O_885,N_14062,N_13720);
nor UO_886 (O_886,N_14831,N_13833);
or UO_887 (O_887,N_14015,N_14322);
nand UO_888 (O_888,N_14456,N_13900);
and UO_889 (O_889,N_14500,N_13714);
and UO_890 (O_890,N_14579,N_14245);
and UO_891 (O_891,N_14904,N_14159);
nand UO_892 (O_892,N_14716,N_14961);
nor UO_893 (O_893,N_13815,N_14545);
nand UO_894 (O_894,N_14139,N_14103);
and UO_895 (O_895,N_14467,N_13870);
nand UO_896 (O_896,N_14762,N_14005);
or UO_897 (O_897,N_13652,N_14202);
nand UO_898 (O_898,N_13939,N_14838);
nand UO_899 (O_899,N_13546,N_13794);
and UO_900 (O_900,N_14232,N_13530);
or UO_901 (O_901,N_14846,N_13829);
and UO_902 (O_902,N_13933,N_14648);
and UO_903 (O_903,N_13852,N_14911);
nor UO_904 (O_904,N_14924,N_14280);
and UO_905 (O_905,N_14729,N_13864);
or UO_906 (O_906,N_13604,N_14250);
and UO_907 (O_907,N_14271,N_14402);
nor UO_908 (O_908,N_13884,N_14775);
nor UO_909 (O_909,N_14710,N_14726);
nand UO_910 (O_910,N_14419,N_14634);
nand UO_911 (O_911,N_14761,N_14532);
or UO_912 (O_912,N_14693,N_14929);
xor UO_913 (O_913,N_13823,N_13648);
nor UO_914 (O_914,N_14461,N_14685);
nand UO_915 (O_915,N_13554,N_14834);
and UO_916 (O_916,N_13549,N_14095);
or UO_917 (O_917,N_14476,N_14955);
and UO_918 (O_918,N_14903,N_13831);
nand UO_919 (O_919,N_13702,N_13646);
and UO_920 (O_920,N_13894,N_14926);
nand UO_921 (O_921,N_14870,N_14756);
or UO_922 (O_922,N_14904,N_14669);
or UO_923 (O_923,N_14907,N_14608);
nand UO_924 (O_924,N_14438,N_14689);
xnor UO_925 (O_925,N_14695,N_14810);
xor UO_926 (O_926,N_14715,N_14879);
nor UO_927 (O_927,N_13503,N_14229);
xnor UO_928 (O_928,N_14957,N_13660);
xor UO_929 (O_929,N_14605,N_13744);
and UO_930 (O_930,N_14096,N_13648);
or UO_931 (O_931,N_13976,N_13796);
or UO_932 (O_932,N_14925,N_14190);
nor UO_933 (O_933,N_13657,N_14366);
nand UO_934 (O_934,N_14191,N_14564);
nor UO_935 (O_935,N_14495,N_14712);
and UO_936 (O_936,N_14263,N_14075);
nor UO_937 (O_937,N_14245,N_14524);
nand UO_938 (O_938,N_14272,N_14497);
nand UO_939 (O_939,N_13623,N_14843);
or UO_940 (O_940,N_14704,N_13626);
nand UO_941 (O_941,N_14738,N_13892);
nand UO_942 (O_942,N_14682,N_13841);
xnor UO_943 (O_943,N_13724,N_13795);
nand UO_944 (O_944,N_14136,N_14117);
and UO_945 (O_945,N_14392,N_13551);
nor UO_946 (O_946,N_14483,N_14528);
or UO_947 (O_947,N_14323,N_13977);
xnor UO_948 (O_948,N_14642,N_14428);
xnor UO_949 (O_949,N_14895,N_14025);
and UO_950 (O_950,N_13702,N_13752);
and UO_951 (O_951,N_13547,N_14861);
nand UO_952 (O_952,N_14481,N_14310);
and UO_953 (O_953,N_14135,N_14924);
or UO_954 (O_954,N_14915,N_14430);
and UO_955 (O_955,N_14346,N_14562);
xnor UO_956 (O_956,N_14967,N_13978);
nor UO_957 (O_957,N_14235,N_14801);
or UO_958 (O_958,N_14316,N_14661);
nand UO_959 (O_959,N_13837,N_13590);
and UO_960 (O_960,N_13700,N_14073);
nor UO_961 (O_961,N_14654,N_13727);
nand UO_962 (O_962,N_14658,N_14629);
and UO_963 (O_963,N_13673,N_14939);
or UO_964 (O_964,N_13703,N_14956);
nor UO_965 (O_965,N_13992,N_14778);
and UO_966 (O_966,N_14645,N_14494);
or UO_967 (O_967,N_14449,N_14882);
and UO_968 (O_968,N_14719,N_14724);
or UO_969 (O_969,N_14492,N_13857);
or UO_970 (O_970,N_14810,N_14062);
nand UO_971 (O_971,N_13744,N_14310);
nor UO_972 (O_972,N_14385,N_14542);
or UO_973 (O_973,N_13932,N_14224);
nor UO_974 (O_974,N_14186,N_14833);
or UO_975 (O_975,N_14087,N_14163);
or UO_976 (O_976,N_13520,N_14896);
and UO_977 (O_977,N_14269,N_14384);
or UO_978 (O_978,N_14563,N_14345);
or UO_979 (O_979,N_13970,N_14022);
and UO_980 (O_980,N_13727,N_14763);
nand UO_981 (O_981,N_14337,N_14975);
or UO_982 (O_982,N_13912,N_13648);
nand UO_983 (O_983,N_13845,N_14417);
xnor UO_984 (O_984,N_13700,N_14327);
or UO_985 (O_985,N_14251,N_13630);
nor UO_986 (O_986,N_14375,N_14339);
nand UO_987 (O_987,N_13593,N_14633);
nor UO_988 (O_988,N_14858,N_13589);
or UO_989 (O_989,N_13616,N_14829);
and UO_990 (O_990,N_13738,N_14856);
or UO_991 (O_991,N_14452,N_14033);
or UO_992 (O_992,N_13860,N_14902);
and UO_993 (O_993,N_13985,N_14302);
nor UO_994 (O_994,N_14141,N_14908);
nor UO_995 (O_995,N_14556,N_14882);
or UO_996 (O_996,N_14259,N_13950);
or UO_997 (O_997,N_14176,N_14895);
nor UO_998 (O_998,N_14556,N_13664);
nor UO_999 (O_999,N_14899,N_14534);
and UO_1000 (O_1000,N_14766,N_13963);
and UO_1001 (O_1001,N_14168,N_13556);
and UO_1002 (O_1002,N_13805,N_14675);
and UO_1003 (O_1003,N_13665,N_14757);
nand UO_1004 (O_1004,N_13671,N_14081);
nand UO_1005 (O_1005,N_14973,N_14769);
xor UO_1006 (O_1006,N_14006,N_14908);
or UO_1007 (O_1007,N_14247,N_14848);
nor UO_1008 (O_1008,N_13912,N_14194);
and UO_1009 (O_1009,N_13819,N_13507);
or UO_1010 (O_1010,N_14133,N_14082);
nand UO_1011 (O_1011,N_13591,N_13769);
nor UO_1012 (O_1012,N_14342,N_14158);
nand UO_1013 (O_1013,N_13703,N_14553);
nor UO_1014 (O_1014,N_13738,N_14285);
and UO_1015 (O_1015,N_14749,N_14571);
and UO_1016 (O_1016,N_13524,N_14860);
or UO_1017 (O_1017,N_13831,N_13991);
nor UO_1018 (O_1018,N_13763,N_14132);
nand UO_1019 (O_1019,N_14999,N_14200);
xor UO_1020 (O_1020,N_14010,N_14888);
nand UO_1021 (O_1021,N_14481,N_14844);
or UO_1022 (O_1022,N_14453,N_14690);
nor UO_1023 (O_1023,N_13553,N_14221);
and UO_1024 (O_1024,N_14617,N_14873);
or UO_1025 (O_1025,N_13595,N_13698);
xor UO_1026 (O_1026,N_14443,N_13560);
and UO_1027 (O_1027,N_13915,N_13863);
xor UO_1028 (O_1028,N_14904,N_13956);
xnor UO_1029 (O_1029,N_13585,N_13769);
or UO_1030 (O_1030,N_13781,N_14275);
nand UO_1031 (O_1031,N_14800,N_13806);
nand UO_1032 (O_1032,N_14557,N_13718);
and UO_1033 (O_1033,N_13537,N_14062);
nor UO_1034 (O_1034,N_13565,N_14333);
nand UO_1035 (O_1035,N_14976,N_13613);
and UO_1036 (O_1036,N_13973,N_14322);
and UO_1037 (O_1037,N_13928,N_14987);
xnor UO_1038 (O_1038,N_14536,N_13506);
or UO_1039 (O_1039,N_14956,N_14475);
nand UO_1040 (O_1040,N_14689,N_13961);
nor UO_1041 (O_1041,N_14599,N_14994);
or UO_1042 (O_1042,N_13763,N_14325);
or UO_1043 (O_1043,N_13592,N_13956);
nor UO_1044 (O_1044,N_13594,N_14481);
xor UO_1045 (O_1045,N_14073,N_14634);
or UO_1046 (O_1046,N_14713,N_14097);
xor UO_1047 (O_1047,N_14789,N_14683);
and UO_1048 (O_1048,N_13965,N_13997);
nor UO_1049 (O_1049,N_13615,N_14719);
or UO_1050 (O_1050,N_13769,N_14154);
nand UO_1051 (O_1051,N_14716,N_14747);
xor UO_1052 (O_1052,N_14122,N_14899);
nor UO_1053 (O_1053,N_14170,N_14330);
nand UO_1054 (O_1054,N_13551,N_13601);
or UO_1055 (O_1055,N_14621,N_13817);
or UO_1056 (O_1056,N_13717,N_14433);
nand UO_1057 (O_1057,N_14166,N_14576);
xor UO_1058 (O_1058,N_14300,N_13891);
or UO_1059 (O_1059,N_13634,N_13737);
nor UO_1060 (O_1060,N_14109,N_14457);
and UO_1061 (O_1061,N_14271,N_14619);
and UO_1062 (O_1062,N_14278,N_13903);
nand UO_1063 (O_1063,N_13741,N_13620);
nand UO_1064 (O_1064,N_14100,N_14067);
nor UO_1065 (O_1065,N_14996,N_14628);
xor UO_1066 (O_1066,N_13656,N_14379);
or UO_1067 (O_1067,N_14171,N_13652);
nor UO_1068 (O_1068,N_14345,N_14057);
and UO_1069 (O_1069,N_13896,N_14407);
and UO_1070 (O_1070,N_14766,N_14238);
and UO_1071 (O_1071,N_14854,N_14881);
nand UO_1072 (O_1072,N_14842,N_13640);
nor UO_1073 (O_1073,N_13644,N_13662);
and UO_1074 (O_1074,N_14085,N_14933);
nand UO_1075 (O_1075,N_14029,N_13643);
nand UO_1076 (O_1076,N_14236,N_13529);
and UO_1077 (O_1077,N_13853,N_14565);
nor UO_1078 (O_1078,N_13815,N_14821);
nand UO_1079 (O_1079,N_13547,N_13524);
and UO_1080 (O_1080,N_13544,N_14217);
nor UO_1081 (O_1081,N_14788,N_13937);
xnor UO_1082 (O_1082,N_14902,N_14790);
or UO_1083 (O_1083,N_14866,N_14922);
and UO_1084 (O_1084,N_13864,N_13750);
or UO_1085 (O_1085,N_13812,N_14553);
nor UO_1086 (O_1086,N_14305,N_14418);
nor UO_1087 (O_1087,N_14188,N_13892);
nor UO_1088 (O_1088,N_13541,N_14733);
nand UO_1089 (O_1089,N_13786,N_13788);
or UO_1090 (O_1090,N_13596,N_13962);
nor UO_1091 (O_1091,N_14120,N_13832);
nand UO_1092 (O_1092,N_14750,N_14241);
nand UO_1093 (O_1093,N_13995,N_14411);
nand UO_1094 (O_1094,N_14196,N_14099);
or UO_1095 (O_1095,N_14707,N_14110);
xnor UO_1096 (O_1096,N_14190,N_14306);
or UO_1097 (O_1097,N_14445,N_14417);
xor UO_1098 (O_1098,N_14648,N_13782);
or UO_1099 (O_1099,N_13801,N_13874);
or UO_1100 (O_1100,N_13500,N_14735);
nor UO_1101 (O_1101,N_13688,N_14979);
nor UO_1102 (O_1102,N_14308,N_14445);
nand UO_1103 (O_1103,N_14687,N_14287);
or UO_1104 (O_1104,N_14023,N_13539);
and UO_1105 (O_1105,N_14917,N_14760);
nand UO_1106 (O_1106,N_14866,N_13688);
nand UO_1107 (O_1107,N_13591,N_14304);
xor UO_1108 (O_1108,N_14791,N_13719);
nor UO_1109 (O_1109,N_14055,N_14228);
nand UO_1110 (O_1110,N_13968,N_14345);
nor UO_1111 (O_1111,N_14760,N_14706);
or UO_1112 (O_1112,N_14035,N_13989);
nand UO_1113 (O_1113,N_14732,N_14102);
nor UO_1114 (O_1114,N_13683,N_14159);
nor UO_1115 (O_1115,N_14367,N_13953);
or UO_1116 (O_1116,N_14703,N_14086);
and UO_1117 (O_1117,N_14331,N_14553);
and UO_1118 (O_1118,N_13781,N_14099);
or UO_1119 (O_1119,N_14503,N_14664);
nor UO_1120 (O_1120,N_14430,N_14776);
xor UO_1121 (O_1121,N_13820,N_14678);
and UO_1122 (O_1122,N_14122,N_14024);
and UO_1123 (O_1123,N_13939,N_13828);
nand UO_1124 (O_1124,N_14762,N_14624);
nand UO_1125 (O_1125,N_13656,N_13575);
and UO_1126 (O_1126,N_13552,N_14252);
nor UO_1127 (O_1127,N_14355,N_14849);
or UO_1128 (O_1128,N_13533,N_13717);
nand UO_1129 (O_1129,N_14658,N_14191);
nor UO_1130 (O_1130,N_13688,N_13691);
and UO_1131 (O_1131,N_14200,N_14228);
or UO_1132 (O_1132,N_14183,N_14316);
and UO_1133 (O_1133,N_14949,N_13620);
or UO_1134 (O_1134,N_14963,N_14129);
or UO_1135 (O_1135,N_13942,N_14624);
nor UO_1136 (O_1136,N_13746,N_14281);
or UO_1137 (O_1137,N_13972,N_14838);
nor UO_1138 (O_1138,N_14418,N_13837);
nor UO_1139 (O_1139,N_14798,N_14768);
and UO_1140 (O_1140,N_14885,N_14497);
nand UO_1141 (O_1141,N_14848,N_14752);
nand UO_1142 (O_1142,N_14780,N_14358);
and UO_1143 (O_1143,N_14284,N_14555);
xnor UO_1144 (O_1144,N_13573,N_14485);
and UO_1145 (O_1145,N_14880,N_13852);
xnor UO_1146 (O_1146,N_13989,N_14484);
xor UO_1147 (O_1147,N_13666,N_14321);
nor UO_1148 (O_1148,N_13902,N_14433);
xnor UO_1149 (O_1149,N_13626,N_13935);
nor UO_1150 (O_1150,N_14717,N_14935);
or UO_1151 (O_1151,N_14638,N_13689);
nor UO_1152 (O_1152,N_14156,N_14477);
nand UO_1153 (O_1153,N_13685,N_13670);
nand UO_1154 (O_1154,N_13527,N_13730);
and UO_1155 (O_1155,N_13550,N_14908);
nand UO_1156 (O_1156,N_14316,N_13997);
or UO_1157 (O_1157,N_14680,N_14726);
nand UO_1158 (O_1158,N_14504,N_14212);
nand UO_1159 (O_1159,N_14005,N_14673);
and UO_1160 (O_1160,N_14478,N_14373);
xnor UO_1161 (O_1161,N_14885,N_13950);
nand UO_1162 (O_1162,N_14953,N_14397);
nand UO_1163 (O_1163,N_14295,N_13941);
xnor UO_1164 (O_1164,N_14903,N_13887);
nand UO_1165 (O_1165,N_14158,N_14323);
or UO_1166 (O_1166,N_14698,N_14412);
nor UO_1167 (O_1167,N_14979,N_14942);
nor UO_1168 (O_1168,N_14006,N_14320);
nor UO_1169 (O_1169,N_14228,N_14676);
nor UO_1170 (O_1170,N_14682,N_14184);
nor UO_1171 (O_1171,N_13996,N_14775);
and UO_1172 (O_1172,N_14591,N_14425);
or UO_1173 (O_1173,N_14645,N_14773);
nand UO_1174 (O_1174,N_14268,N_14540);
nor UO_1175 (O_1175,N_13756,N_14256);
nand UO_1176 (O_1176,N_14196,N_13836);
nor UO_1177 (O_1177,N_14507,N_13912);
or UO_1178 (O_1178,N_14474,N_14122);
xor UO_1179 (O_1179,N_14127,N_14333);
nand UO_1180 (O_1180,N_14444,N_13992);
nand UO_1181 (O_1181,N_13708,N_13867);
or UO_1182 (O_1182,N_13953,N_13755);
and UO_1183 (O_1183,N_14437,N_14787);
and UO_1184 (O_1184,N_14942,N_14650);
nand UO_1185 (O_1185,N_13832,N_13918);
xnor UO_1186 (O_1186,N_14576,N_14266);
or UO_1187 (O_1187,N_14500,N_13801);
and UO_1188 (O_1188,N_14802,N_14902);
nand UO_1189 (O_1189,N_14542,N_14189);
or UO_1190 (O_1190,N_13883,N_13661);
nor UO_1191 (O_1191,N_13821,N_14211);
or UO_1192 (O_1192,N_13545,N_13784);
and UO_1193 (O_1193,N_14262,N_13566);
nor UO_1194 (O_1194,N_13873,N_13968);
and UO_1195 (O_1195,N_14879,N_14718);
and UO_1196 (O_1196,N_14655,N_14810);
xor UO_1197 (O_1197,N_14189,N_14799);
or UO_1198 (O_1198,N_14413,N_13536);
nand UO_1199 (O_1199,N_13775,N_14738);
xor UO_1200 (O_1200,N_14410,N_14114);
nor UO_1201 (O_1201,N_13861,N_14475);
or UO_1202 (O_1202,N_13720,N_14352);
or UO_1203 (O_1203,N_14742,N_14178);
or UO_1204 (O_1204,N_13777,N_14944);
and UO_1205 (O_1205,N_14327,N_13980);
or UO_1206 (O_1206,N_14471,N_14627);
or UO_1207 (O_1207,N_13914,N_14581);
nor UO_1208 (O_1208,N_14537,N_14329);
nor UO_1209 (O_1209,N_14505,N_14117);
or UO_1210 (O_1210,N_14936,N_14949);
nand UO_1211 (O_1211,N_14516,N_14612);
xnor UO_1212 (O_1212,N_14850,N_14549);
and UO_1213 (O_1213,N_14524,N_13790);
and UO_1214 (O_1214,N_13733,N_14690);
and UO_1215 (O_1215,N_14483,N_13855);
nor UO_1216 (O_1216,N_14406,N_14256);
nor UO_1217 (O_1217,N_13916,N_14961);
or UO_1218 (O_1218,N_14609,N_14157);
or UO_1219 (O_1219,N_13839,N_13962);
or UO_1220 (O_1220,N_14406,N_13946);
and UO_1221 (O_1221,N_13950,N_14890);
and UO_1222 (O_1222,N_14258,N_13971);
nor UO_1223 (O_1223,N_14621,N_14635);
and UO_1224 (O_1224,N_14028,N_13624);
xor UO_1225 (O_1225,N_14678,N_13758);
or UO_1226 (O_1226,N_14061,N_13823);
and UO_1227 (O_1227,N_13582,N_13807);
and UO_1228 (O_1228,N_13994,N_14925);
nand UO_1229 (O_1229,N_13652,N_13946);
nor UO_1230 (O_1230,N_14809,N_14037);
nand UO_1231 (O_1231,N_14464,N_14095);
and UO_1232 (O_1232,N_14479,N_14358);
nor UO_1233 (O_1233,N_14811,N_14114);
or UO_1234 (O_1234,N_13637,N_14026);
nor UO_1235 (O_1235,N_13986,N_14848);
xor UO_1236 (O_1236,N_14809,N_14990);
and UO_1237 (O_1237,N_14866,N_13629);
or UO_1238 (O_1238,N_14253,N_14294);
nand UO_1239 (O_1239,N_13525,N_13684);
or UO_1240 (O_1240,N_14872,N_14286);
nand UO_1241 (O_1241,N_13977,N_13754);
nand UO_1242 (O_1242,N_14240,N_14596);
xnor UO_1243 (O_1243,N_13948,N_14454);
xor UO_1244 (O_1244,N_14525,N_13691);
xor UO_1245 (O_1245,N_14273,N_13769);
nand UO_1246 (O_1246,N_14794,N_14407);
xnor UO_1247 (O_1247,N_13716,N_14736);
or UO_1248 (O_1248,N_14842,N_13746);
and UO_1249 (O_1249,N_13510,N_14973);
or UO_1250 (O_1250,N_13706,N_14001);
xnor UO_1251 (O_1251,N_13745,N_14422);
and UO_1252 (O_1252,N_14456,N_14453);
nor UO_1253 (O_1253,N_14471,N_14954);
or UO_1254 (O_1254,N_13924,N_14328);
or UO_1255 (O_1255,N_14896,N_13937);
and UO_1256 (O_1256,N_14623,N_13789);
and UO_1257 (O_1257,N_14722,N_14833);
nand UO_1258 (O_1258,N_13802,N_14917);
and UO_1259 (O_1259,N_14093,N_13786);
nor UO_1260 (O_1260,N_14999,N_13756);
or UO_1261 (O_1261,N_13918,N_14487);
nor UO_1262 (O_1262,N_14672,N_13923);
nor UO_1263 (O_1263,N_13652,N_14148);
nand UO_1264 (O_1264,N_13509,N_14426);
nor UO_1265 (O_1265,N_14349,N_14489);
and UO_1266 (O_1266,N_14186,N_14028);
nand UO_1267 (O_1267,N_13782,N_13662);
nand UO_1268 (O_1268,N_14488,N_13728);
nand UO_1269 (O_1269,N_13795,N_14664);
nand UO_1270 (O_1270,N_14172,N_14161);
and UO_1271 (O_1271,N_13544,N_13879);
and UO_1272 (O_1272,N_13967,N_14833);
xnor UO_1273 (O_1273,N_14666,N_13546);
or UO_1274 (O_1274,N_14454,N_14176);
nand UO_1275 (O_1275,N_14219,N_14922);
nand UO_1276 (O_1276,N_14852,N_14217);
xor UO_1277 (O_1277,N_13663,N_14650);
nand UO_1278 (O_1278,N_13692,N_14841);
nor UO_1279 (O_1279,N_14603,N_14795);
and UO_1280 (O_1280,N_14831,N_13611);
xor UO_1281 (O_1281,N_14651,N_14648);
nor UO_1282 (O_1282,N_13681,N_14489);
nand UO_1283 (O_1283,N_13859,N_14652);
nand UO_1284 (O_1284,N_14898,N_14528);
and UO_1285 (O_1285,N_14384,N_13940);
or UO_1286 (O_1286,N_14679,N_13670);
or UO_1287 (O_1287,N_13774,N_13757);
nor UO_1288 (O_1288,N_13622,N_14365);
and UO_1289 (O_1289,N_14541,N_14617);
or UO_1290 (O_1290,N_14651,N_14978);
nand UO_1291 (O_1291,N_14924,N_13766);
nor UO_1292 (O_1292,N_14346,N_14766);
nand UO_1293 (O_1293,N_14710,N_14035);
or UO_1294 (O_1294,N_14947,N_14031);
nand UO_1295 (O_1295,N_14637,N_14554);
or UO_1296 (O_1296,N_14158,N_14306);
and UO_1297 (O_1297,N_13980,N_14532);
and UO_1298 (O_1298,N_13833,N_14107);
and UO_1299 (O_1299,N_13982,N_14195);
xnor UO_1300 (O_1300,N_14831,N_14164);
or UO_1301 (O_1301,N_14114,N_14210);
nand UO_1302 (O_1302,N_14366,N_14077);
nor UO_1303 (O_1303,N_13696,N_14971);
nor UO_1304 (O_1304,N_14453,N_14222);
nor UO_1305 (O_1305,N_13698,N_14307);
nor UO_1306 (O_1306,N_14293,N_14928);
nor UO_1307 (O_1307,N_13832,N_13755);
or UO_1308 (O_1308,N_13524,N_14936);
nand UO_1309 (O_1309,N_13987,N_14394);
nand UO_1310 (O_1310,N_13824,N_13652);
or UO_1311 (O_1311,N_13714,N_14818);
or UO_1312 (O_1312,N_14178,N_13783);
and UO_1313 (O_1313,N_14149,N_14635);
or UO_1314 (O_1314,N_14433,N_13745);
and UO_1315 (O_1315,N_14988,N_14212);
nor UO_1316 (O_1316,N_14959,N_13706);
nor UO_1317 (O_1317,N_14315,N_14577);
nand UO_1318 (O_1318,N_14542,N_14658);
nor UO_1319 (O_1319,N_14830,N_14334);
nand UO_1320 (O_1320,N_14761,N_13685);
nand UO_1321 (O_1321,N_14427,N_14215);
or UO_1322 (O_1322,N_14349,N_14235);
and UO_1323 (O_1323,N_14894,N_14886);
or UO_1324 (O_1324,N_13821,N_13827);
nor UO_1325 (O_1325,N_14776,N_13961);
xor UO_1326 (O_1326,N_14058,N_14586);
xor UO_1327 (O_1327,N_13637,N_14814);
nor UO_1328 (O_1328,N_14790,N_13559);
nand UO_1329 (O_1329,N_13815,N_14089);
nand UO_1330 (O_1330,N_14749,N_13973);
and UO_1331 (O_1331,N_14488,N_13977);
xor UO_1332 (O_1332,N_14911,N_13756);
xnor UO_1333 (O_1333,N_13946,N_14507);
nor UO_1334 (O_1334,N_14069,N_13923);
xnor UO_1335 (O_1335,N_14754,N_13663);
and UO_1336 (O_1336,N_14268,N_13650);
xor UO_1337 (O_1337,N_14953,N_14797);
nand UO_1338 (O_1338,N_14593,N_14818);
and UO_1339 (O_1339,N_13588,N_13568);
or UO_1340 (O_1340,N_14439,N_14778);
nor UO_1341 (O_1341,N_14947,N_14328);
or UO_1342 (O_1342,N_14669,N_13658);
or UO_1343 (O_1343,N_13739,N_14398);
nor UO_1344 (O_1344,N_14426,N_14142);
nand UO_1345 (O_1345,N_14658,N_14711);
or UO_1346 (O_1346,N_13706,N_13830);
nand UO_1347 (O_1347,N_13786,N_13936);
xnor UO_1348 (O_1348,N_14624,N_13903);
or UO_1349 (O_1349,N_14007,N_13684);
and UO_1350 (O_1350,N_14942,N_13508);
nor UO_1351 (O_1351,N_14458,N_14752);
nand UO_1352 (O_1352,N_13883,N_13701);
nor UO_1353 (O_1353,N_13816,N_13971);
and UO_1354 (O_1354,N_13795,N_13738);
nor UO_1355 (O_1355,N_14698,N_14664);
or UO_1356 (O_1356,N_14736,N_14745);
xor UO_1357 (O_1357,N_14205,N_14854);
nor UO_1358 (O_1358,N_13671,N_13837);
and UO_1359 (O_1359,N_14375,N_14655);
xor UO_1360 (O_1360,N_14370,N_14162);
nand UO_1361 (O_1361,N_13554,N_14315);
nand UO_1362 (O_1362,N_14127,N_13521);
nor UO_1363 (O_1363,N_14514,N_14947);
nand UO_1364 (O_1364,N_13676,N_14291);
or UO_1365 (O_1365,N_14720,N_13774);
and UO_1366 (O_1366,N_14845,N_13635);
nor UO_1367 (O_1367,N_14859,N_14434);
and UO_1368 (O_1368,N_14910,N_14752);
and UO_1369 (O_1369,N_13742,N_13867);
nand UO_1370 (O_1370,N_14616,N_14970);
or UO_1371 (O_1371,N_14414,N_13869);
or UO_1372 (O_1372,N_14057,N_13628);
or UO_1373 (O_1373,N_14706,N_14988);
nor UO_1374 (O_1374,N_13735,N_13677);
nor UO_1375 (O_1375,N_13517,N_14982);
nor UO_1376 (O_1376,N_14881,N_13706);
nand UO_1377 (O_1377,N_14215,N_14113);
nand UO_1378 (O_1378,N_14792,N_14054);
and UO_1379 (O_1379,N_14843,N_14678);
nand UO_1380 (O_1380,N_13826,N_14516);
nor UO_1381 (O_1381,N_14696,N_14527);
or UO_1382 (O_1382,N_13655,N_14948);
or UO_1383 (O_1383,N_13669,N_14583);
or UO_1384 (O_1384,N_13954,N_13787);
nand UO_1385 (O_1385,N_14106,N_14666);
nand UO_1386 (O_1386,N_13869,N_13707);
and UO_1387 (O_1387,N_14591,N_13618);
nor UO_1388 (O_1388,N_14383,N_13837);
or UO_1389 (O_1389,N_13514,N_14258);
and UO_1390 (O_1390,N_14692,N_14866);
nand UO_1391 (O_1391,N_14550,N_13666);
nand UO_1392 (O_1392,N_14943,N_14482);
or UO_1393 (O_1393,N_13513,N_13932);
and UO_1394 (O_1394,N_14210,N_14031);
or UO_1395 (O_1395,N_14847,N_13843);
nor UO_1396 (O_1396,N_13892,N_14066);
nor UO_1397 (O_1397,N_14626,N_14934);
and UO_1398 (O_1398,N_14539,N_13544);
nand UO_1399 (O_1399,N_14050,N_14338);
nand UO_1400 (O_1400,N_14303,N_14990);
and UO_1401 (O_1401,N_14457,N_14572);
and UO_1402 (O_1402,N_13736,N_14167);
xnor UO_1403 (O_1403,N_14522,N_14134);
or UO_1404 (O_1404,N_13531,N_13922);
xnor UO_1405 (O_1405,N_14032,N_14621);
nand UO_1406 (O_1406,N_14360,N_13838);
or UO_1407 (O_1407,N_13924,N_13613);
or UO_1408 (O_1408,N_14278,N_14167);
nor UO_1409 (O_1409,N_13981,N_14231);
and UO_1410 (O_1410,N_14040,N_14254);
and UO_1411 (O_1411,N_14624,N_14274);
or UO_1412 (O_1412,N_13970,N_14852);
and UO_1413 (O_1413,N_14144,N_13920);
nand UO_1414 (O_1414,N_13505,N_13799);
nand UO_1415 (O_1415,N_14732,N_14458);
nor UO_1416 (O_1416,N_14643,N_13825);
nand UO_1417 (O_1417,N_13661,N_14880);
and UO_1418 (O_1418,N_14089,N_14764);
nand UO_1419 (O_1419,N_14898,N_14768);
nand UO_1420 (O_1420,N_14341,N_14771);
nor UO_1421 (O_1421,N_14291,N_14259);
and UO_1422 (O_1422,N_14665,N_14518);
or UO_1423 (O_1423,N_13724,N_14654);
or UO_1424 (O_1424,N_14081,N_13548);
xnor UO_1425 (O_1425,N_14604,N_14950);
nand UO_1426 (O_1426,N_14262,N_14554);
or UO_1427 (O_1427,N_14339,N_14104);
nor UO_1428 (O_1428,N_14036,N_14131);
or UO_1429 (O_1429,N_13851,N_14334);
nor UO_1430 (O_1430,N_14814,N_13912);
or UO_1431 (O_1431,N_14698,N_13799);
nand UO_1432 (O_1432,N_14020,N_14448);
nor UO_1433 (O_1433,N_13815,N_14969);
or UO_1434 (O_1434,N_13854,N_13745);
xor UO_1435 (O_1435,N_14992,N_13926);
nand UO_1436 (O_1436,N_13724,N_14351);
nand UO_1437 (O_1437,N_14849,N_14767);
and UO_1438 (O_1438,N_14087,N_14660);
nor UO_1439 (O_1439,N_13605,N_14266);
or UO_1440 (O_1440,N_14714,N_14479);
or UO_1441 (O_1441,N_13920,N_14282);
nand UO_1442 (O_1442,N_13809,N_14703);
or UO_1443 (O_1443,N_14114,N_14497);
nor UO_1444 (O_1444,N_13814,N_14471);
nor UO_1445 (O_1445,N_13677,N_14711);
or UO_1446 (O_1446,N_14319,N_14544);
and UO_1447 (O_1447,N_14432,N_13540);
xor UO_1448 (O_1448,N_14225,N_14908);
and UO_1449 (O_1449,N_14104,N_14800);
nand UO_1450 (O_1450,N_14189,N_14365);
nand UO_1451 (O_1451,N_13659,N_14343);
nor UO_1452 (O_1452,N_13822,N_14238);
nor UO_1453 (O_1453,N_13640,N_14032);
and UO_1454 (O_1454,N_13849,N_13770);
nand UO_1455 (O_1455,N_14692,N_14084);
nand UO_1456 (O_1456,N_14945,N_13925);
nand UO_1457 (O_1457,N_14548,N_14606);
or UO_1458 (O_1458,N_14944,N_14101);
and UO_1459 (O_1459,N_14337,N_14165);
nand UO_1460 (O_1460,N_14115,N_14956);
nor UO_1461 (O_1461,N_14207,N_13863);
or UO_1462 (O_1462,N_14186,N_14638);
nor UO_1463 (O_1463,N_13803,N_14794);
and UO_1464 (O_1464,N_14025,N_14956);
and UO_1465 (O_1465,N_13572,N_13938);
nand UO_1466 (O_1466,N_13502,N_14767);
and UO_1467 (O_1467,N_13755,N_14091);
and UO_1468 (O_1468,N_13600,N_14104);
nand UO_1469 (O_1469,N_13513,N_14475);
and UO_1470 (O_1470,N_14427,N_13961);
xor UO_1471 (O_1471,N_13887,N_13691);
or UO_1472 (O_1472,N_14016,N_14833);
xnor UO_1473 (O_1473,N_13766,N_13598);
nand UO_1474 (O_1474,N_14775,N_13667);
or UO_1475 (O_1475,N_13827,N_13527);
or UO_1476 (O_1476,N_14870,N_13694);
and UO_1477 (O_1477,N_14996,N_14061);
nor UO_1478 (O_1478,N_14027,N_13713);
nor UO_1479 (O_1479,N_13809,N_14036);
nor UO_1480 (O_1480,N_14216,N_13793);
xor UO_1481 (O_1481,N_13864,N_14906);
and UO_1482 (O_1482,N_14959,N_14722);
or UO_1483 (O_1483,N_13757,N_14202);
and UO_1484 (O_1484,N_14829,N_13935);
and UO_1485 (O_1485,N_13522,N_13591);
xor UO_1486 (O_1486,N_14858,N_14558);
and UO_1487 (O_1487,N_14047,N_13837);
xnor UO_1488 (O_1488,N_13573,N_14342);
xor UO_1489 (O_1489,N_13573,N_13509);
xor UO_1490 (O_1490,N_14321,N_14453);
nor UO_1491 (O_1491,N_14723,N_13645);
and UO_1492 (O_1492,N_14623,N_14445);
nor UO_1493 (O_1493,N_14855,N_14486);
and UO_1494 (O_1494,N_13574,N_14187);
nand UO_1495 (O_1495,N_14685,N_14978);
nor UO_1496 (O_1496,N_13606,N_13547);
nor UO_1497 (O_1497,N_13691,N_14300);
nor UO_1498 (O_1498,N_14340,N_14529);
nand UO_1499 (O_1499,N_14657,N_14595);
nor UO_1500 (O_1500,N_14708,N_14226);
nor UO_1501 (O_1501,N_14146,N_14287);
or UO_1502 (O_1502,N_14920,N_14190);
or UO_1503 (O_1503,N_13829,N_14208);
nor UO_1504 (O_1504,N_13723,N_13523);
nand UO_1505 (O_1505,N_14119,N_14910);
or UO_1506 (O_1506,N_13507,N_13571);
and UO_1507 (O_1507,N_13508,N_13780);
nor UO_1508 (O_1508,N_14121,N_14980);
or UO_1509 (O_1509,N_13859,N_13611);
or UO_1510 (O_1510,N_14477,N_14319);
nand UO_1511 (O_1511,N_13841,N_14707);
or UO_1512 (O_1512,N_13516,N_13672);
or UO_1513 (O_1513,N_13826,N_14716);
or UO_1514 (O_1514,N_14203,N_14550);
and UO_1515 (O_1515,N_14011,N_14044);
and UO_1516 (O_1516,N_14327,N_14343);
xnor UO_1517 (O_1517,N_13617,N_14404);
nand UO_1518 (O_1518,N_14399,N_14128);
and UO_1519 (O_1519,N_13886,N_14749);
nand UO_1520 (O_1520,N_13836,N_13734);
and UO_1521 (O_1521,N_14882,N_14429);
and UO_1522 (O_1522,N_14840,N_13558);
or UO_1523 (O_1523,N_14850,N_13501);
or UO_1524 (O_1524,N_13504,N_13559);
or UO_1525 (O_1525,N_14671,N_13851);
and UO_1526 (O_1526,N_13654,N_14520);
nor UO_1527 (O_1527,N_13915,N_14830);
or UO_1528 (O_1528,N_14273,N_14216);
nor UO_1529 (O_1529,N_14918,N_13592);
or UO_1530 (O_1530,N_14159,N_14527);
or UO_1531 (O_1531,N_13834,N_13835);
nor UO_1532 (O_1532,N_13829,N_13781);
or UO_1533 (O_1533,N_14153,N_14381);
and UO_1534 (O_1534,N_14024,N_13995);
and UO_1535 (O_1535,N_14179,N_13604);
and UO_1536 (O_1536,N_13577,N_14054);
or UO_1537 (O_1537,N_14205,N_14089);
and UO_1538 (O_1538,N_14949,N_13990);
and UO_1539 (O_1539,N_13895,N_14822);
and UO_1540 (O_1540,N_14074,N_13626);
xnor UO_1541 (O_1541,N_13739,N_13747);
nand UO_1542 (O_1542,N_13730,N_14668);
or UO_1543 (O_1543,N_14976,N_14689);
or UO_1544 (O_1544,N_14025,N_14264);
nor UO_1545 (O_1545,N_14319,N_14745);
and UO_1546 (O_1546,N_14838,N_13562);
or UO_1547 (O_1547,N_13762,N_14538);
nor UO_1548 (O_1548,N_13819,N_14565);
or UO_1549 (O_1549,N_13776,N_14234);
or UO_1550 (O_1550,N_13660,N_13786);
and UO_1551 (O_1551,N_13636,N_14116);
nor UO_1552 (O_1552,N_13813,N_14563);
nand UO_1553 (O_1553,N_14824,N_14778);
or UO_1554 (O_1554,N_13902,N_13768);
or UO_1555 (O_1555,N_14012,N_13644);
or UO_1556 (O_1556,N_14298,N_13874);
and UO_1557 (O_1557,N_13528,N_14894);
nor UO_1558 (O_1558,N_13863,N_13763);
nand UO_1559 (O_1559,N_14382,N_13659);
nor UO_1560 (O_1560,N_13755,N_14876);
and UO_1561 (O_1561,N_14194,N_14448);
nand UO_1562 (O_1562,N_14895,N_14810);
xor UO_1563 (O_1563,N_14479,N_14436);
xor UO_1564 (O_1564,N_13828,N_14915);
nand UO_1565 (O_1565,N_14304,N_13822);
or UO_1566 (O_1566,N_14858,N_14515);
nand UO_1567 (O_1567,N_14680,N_13679);
and UO_1568 (O_1568,N_14383,N_14943);
and UO_1569 (O_1569,N_14111,N_13795);
nand UO_1570 (O_1570,N_14036,N_14955);
nand UO_1571 (O_1571,N_14243,N_14305);
xnor UO_1572 (O_1572,N_14368,N_13599);
or UO_1573 (O_1573,N_14457,N_14139);
or UO_1574 (O_1574,N_14072,N_14796);
nor UO_1575 (O_1575,N_13831,N_14093);
nand UO_1576 (O_1576,N_14050,N_13917);
and UO_1577 (O_1577,N_13682,N_13542);
xnor UO_1578 (O_1578,N_14902,N_14457);
or UO_1579 (O_1579,N_14499,N_14440);
and UO_1580 (O_1580,N_13856,N_13823);
or UO_1581 (O_1581,N_14921,N_14873);
nand UO_1582 (O_1582,N_14799,N_14872);
nand UO_1583 (O_1583,N_14275,N_14610);
nor UO_1584 (O_1584,N_14962,N_13705);
nor UO_1585 (O_1585,N_14611,N_13929);
xor UO_1586 (O_1586,N_14890,N_14949);
or UO_1587 (O_1587,N_14068,N_14240);
nand UO_1588 (O_1588,N_14134,N_14515);
nor UO_1589 (O_1589,N_14954,N_14660);
nand UO_1590 (O_1590,N_14700,N_14323);
nor UO_1591 (O_1591,N_14418,N_13682);
or UO_1592 (O_1592,N_14719,N_14375);
nand UO_1593 (O_1593,N_14869,N_13684);
and UO_1594 (O_1594,N_14089,N_14559);
and UO_1595 (O_1595,N_14613,N_14645);
and UO_1596 (O_1596,N_14975,N_14518);
nor UO_1597 (O_1597,N_13580,N_13586);
and UO_1598 (O_1598,N_14852,N_14201);
or UO_1599 (O_1599,N_13756,N_13613);
or UO_1600 (O_1600,N_14373,N_14515);
nor UO_1601 (O_1601,N_13683,N_14757);
or UO_1602 (O_1602,N_13738,N_14287);
and UO_1603 (O_1603,N_14133,N_14395);
nor UO_1604 (O_1604,N_13704,N_14906);
nand UO_1605 (O_1605,N_13921,N_14001);
nor UO_1606 (O_1606,N_14743,N_14152);
and UO_1607 (O_1607,N_14188,N_14644);
nand UO_1608 (O_1608,N_13537,N_14896);
and UO_1609 (O_1609,N_13849,N_14820);
xnor UO_1610 (O_1610,N_14469,N_14455);
nor UO_1611 (O_1611,N_13769,N_13887);
or UO_1612 (O_1612,N_13563,N_14948);
and UO_1613 (O_1613,N_13615,N_14696);
and UO_1614 (O_1614,N_14569,N_13522);
or UO_1615 (O_1615,N_14465,N_13588);
nand UO_1616 (O_1616,N_14121,N_13622);
nand UO_1617 (O_1617,N_14865,N_14060);
nand UO_1618 (O_1618,N_13733,N_14639);
nor UO_1619 (O_1619,N_14764,N_14101);
or UO_1620 (O_1620,N_13773,N_14289);
nand UO_1621 (O_1621,N_14443,N_14061);
or UO_1622 (O_1622,N_14569,N_13930);
xor UO_1623 (O_1623,N_14983,N_13929);
nor UO_1624 (O_1624,N_14649,N_14107);
nor UO_1625 (O_1625,N_14805,N_13564);
nand UO_1626 (O_1626,N_13984,N_14699);
nand UO_1627 (O_1627,N_13783,N_14778);
and UO_1628 (O_1628,N_13545,N_14951);
and UO_1629 (O_1629,N_14020,N_14243);
nand UO_1630 (O_1630,N_14614,N_14741);
and UO_1631 (O_1631,N_13924,N_14090);
nand UO_1632 (O_1632,N_14738,N_13500);
nor UO_1633 (O_1633,N_14685,N_14540);
and UO_1634 (O_1634,N_13758,N_14948);
nor UO_1635 (O_1635,N_14615,N_14991);
or UO_1636 (O_1636,N_14976,N_13723);
xnor UO_1637 (O_1637,N_13959,N_14860);
and UO_1638 (O_1638,N_13748,N_13693);
nor UO_1639 (O_1639,N_14387,N_13553);
nor UO_1640 (O_1640,N_14245,N_13567);
nand UO_1641 (O_1641,N_14361,N_14032);
nor UO_1642 (O_1642,N_14957,N_14549);
and UO_1643 (O_1643,N_13683,N_14728);
nand UO_1644 (O_1644,N_14053,N_13855);
or UO_1645 (O_1645,N_14898,N_14961);
or UO_1646 (O_1646,N_14319,N_14283);
nand UO_1647 (O_1647,N_14627,N_14794);
or UO_1648 (O_1648,N_14393,N_14448);
and UO_1649 (O_1649,N_14717,N_13651);
or UO_1650 (O_1650,N_14168,N_14980);
or UO_1651 (O_1651,N_14707,N_14849);
or UO_1652 (O_1652,N_13511,N_14752);
nand UO_1653 (O_1653,N_14237,N_13718);
nor UO_1654 (O_1654,N_14119,N_14568);
or UO_1655 (O_1655,N_13902,N_14309);
and UO_1656 (O_1656,N_14096,N_13525);
nand UO_1657 (O_1657,N_14398,N_14091);
nor UO_1658 (O_1658,N_14182,N_14533);
nor UO_1659 (O_1659,N_14662,N_13838);
and UO_1660 (O_1660,N_14562,N_14082);
and UO_1661 (O_1661,N_14975,N_14113);
and UO_1662 (O_1662,N_14710,N_14228);
xnor UO_1663 (O_1663,N_14106,N_14025);
and UO_1664 (O_1664,N_14385,N_13975);
nor UO_1665 (O_1665,N_14113,N_13514);
or UO_1666 (O_1666,N_14015,N_14065);
and UO_1667 (O_1667,N_14871,N_14154);
nand UO_1668 (O_1668,N_14203,N_14803);
nor UO_1669 (O_1669,N_14439,N_14311);
nor UO_1670 (O_1670,N_14865,N_13511);
or UO_1671 (O_1671,N_13807,N_13590);
or UO_1672 (O_1672,N_13822,N_14206);
and UO_1673 (O_1673,N_14997,N_14583);
nor UO_1674 (O_1674,N_13969,N_14385);
nand UO_1675 (O_1675,N_13914,N_14470);
and UO_1676 (O_1676,N_14904,N_13809);
nor UO_1677 (O_1677,N_13529,N_13767);
and UO_1678 (O_1678,N_14666,N_14614);
and UO_1679 (O_1679,N_13694,N_14639);
and UO_1680 (O_1680,N_14153,N_13976);
or UO_1681 (O_1681,N_14544,N_14408);
and UO_1682 (O_1682,N_14624,N_14476);
nor UO_1683 (O_1683,N_14117,N_13689);
nor UO_1684 (O_1684,N_14425,N_14876);
and UO_1685 (O_1685,N_14070,N_14426);
or UO_1686 (O_1686,N_14674,N_14831);
xnor UO_1687 (O_1687,N_14413,N_13955);
or UO_1688 (O_1688,N_14257,N_14155);
or UO_1689 (O_1689,N_13774,N_13738);
nand UO_1690 (O_1690,N_14795,N_14600);
xnor UO_1691 (O_1691,N_13892,N_14676);
and UO_1692 (O_1692,N_14475,N_14635);
and UO_1693 (O_1693,N_14521,N_14485);
and UO_1694 (O_1694,N_14905,N_13537);
or UO_1695 (O_1695,N_13650,N_14285);
nor UO_1696 (O_1696,N_13838,N_13742);
and UO_1697 (O_1697,N_14733,N_14304);
nand UO_1698 (O_1698,N_14559,N_14799);
and UO_1699 (O_1699,N_14568,N_14723);
or UO_1700 (O_1700,N_13647,N_13812);
xor UO_1701 (O_1701,N_13772,N_13524);
and UO_1702 (O_1702,N_14982,N_14443);
nand UO_1703 (O_1703,N_14403,N_14213);
and UO_1704 (O_1704,N_14435,N_14447);
or UO_1705 (O_1705,N_13513,N_14756);
or UO_1706 (O_1706,N_14767,N_13609);
nand UO_1707 (O_1707,N_13720,N_13859);
or UO_1708 (O_1708,N_14287,N_14308);
and UO_1709 (O_1709,N_14533,N_13915);
nand UO_1710 (O_1710,N_14523,N_14370);
or UO_1711 (O_1711,N_14946,N_14010);
nand UO_1712 (O_1712,N_14348,N_13864);
or UO_1713 (O_1713,N_14963,N_14834);
and UO_1714 (O_1714,N_14490,N_14186);
and UO_1715 (O_1715,N_14010,N_13776);
and UO_1716 (O_1716,N_14855,N_13673);
or UO_1717 (O_1717,N_14927,N_14898);
and UO_1718 (O_1718,N_13888,N_14579);
and UO_1719 (O_1719,N_13530,N_14564);
nand UO_1720 (O_1720,N_14676,N_13505);
or UO_1721 (O_1721,N_14942,N_14157);
and UO_1722 (O_1722,N_13873,N_13831);
nor UO_1723 (O_1723,N_14178,N_14789);
nand UO_1724 (O_1724,N_14404,N_14580);
and UO_1725 (O_1725,N_14821,N_14283);
nand UO_1726 (O_1726,N_14346,N_14583);
or UO_1727 (O_1727,N_14221,N_13605);
nand UO_1728 (O_1728,N_14925,N_13933);
and UO_1729 (O_1729,N_13773,N_13747);
and UO_1730 (O_1730,N_14041,N_14717);
or UO_1731 (O_1731,N_14275,N_13598);
nor UO_1732 (O_1732,N_13858,N_14643);
or UO_1733 (O_1733,N_13770,N_14354);
xor UO_1734 (O_1734,N_13804,N_14852);
nand UO_1735 (O_1735,N_14412,N_14459);
and UO_1736 (O_1736,N_14973,N_13644);
and UO_1737 (O_1737,N_14862,N_14887);
nand UO_1738 (O_1738,N_14353,N_14304);
nand UO_1739 (O_1739,N_14684,N_14021);
nand UO_1740 (O_1740,N_14778,N_13987);
nand UO_1741 (O_1741,N_14474,N_13600);
or UO_1742 (O_1742,N_14264,N_14895);
and UO_1743 (O_1743,N_14145,N_13956);
and UO_1744 (O_1744,N_14323,N_14609);
nand UO_1745 (O_1745,N_14730,N_14881);
and UO_1746 (O_1746,N_14307,N_13647);
nor UO_1747 (O_1747,N_14461,N_13889);
nor UO_1748 (O_1748,N_14589,N_14427);
and UO_1749 (O_1749,N_13564,N_14982);
or UO_1750 (O_1750,N_14988,N_14580);
and UO_1751 (O_1751,N_14694,N_14850);
or UO_1752 (O_1752,N_14437,N_14620);
nor UO_1753 (O_1753,N_14454,N_13629);
or UO_1754 (O_1754,N_14111,N_13737);
nand UO_1755 (O_1755,N_13750,N_13939);
xor UO_1756 (O_1756,N_14768,N_14022);
or UO_1757 (O_1757,N_14046,N_13866);
or UO_1758 (O_1758,N_14250,N_14643);
and UO_1759 (O_1759,N_14955,N_14538);
xor UO_1760 (O_1760,N_14334,N_14999);
or UO_1761 (O_1761,N_14700,N_14168);
xor UO_1762 (O_1762,N_13790,N_14375);
nand UO_1763 (O_1763,N_14053,N_14413);
nor UO_1764 (O_1764,N_14799,N_13787);
xor UO_1765 (O_1765,N_14887,N_14853);
nor UO_1766 (O_1766,N_14696,N_13504);
or UO_1767 (O_1767,N_14168,N_14809);
or UO_1768 (O_1768,N_14162,N_13536);
and UO_1769 (O_1769,N_14276,N_14807);
or UO_1770 (O_1770,N_14651,N_14598);
or UO_1771 (O_1771,N_13882,N_14104);
xor UO_1772 (O_1772,N_13721,N_13825);
and UO_1773 (O_1773,N_14214,N_14688);
nand UO_1774 (O_1774,N_13832,N_14492);
xnor UO_1775 (O_1775,N_14433,N_14719);
or UO_1776 (O_1776,N_13878,N_14409);
nand UO_1777 (O_1777,N_14825,N_13867);
or UO_1778 (O_1778,N_14012,N_13694);
or UO_1779 (O_1779,N_14783,N_13691);
nor UO_1780 (O_1780,N_13514,N_13852);
and UO_1781 (O_1781,N_14059,N_13545);
or UO_1782 (O_1782,N_14430,N_14511);
nor UO_1783 (O_1783,N_13673,N_14705);
nand UO_1784 (O_1784,N_14847,N_14307);
nand UO_1785 (O_1785,N_13717,N_14122);
nor UO_1786 (O_1786,N_13713,N_14026);
nor UO_1787 (O_1787,N_14368,N_14283);
nor UO_1788 (O_1788,N_14117,N_13828);
nand UO_1789 (O_1789,N_14068,N_14950);
nor UO_1790 (O_1790,N_14920,N_14041);
nor UO_1791 (O_1791,N_14158,N_14590);
and UO_1792 (O_1792,N_13749,N_13790);
or UO_1793 (O_1793,N_14185,N_14253);
or UO_1794 (O_1794,N_14026,N_14192);
xnor UO_1795 (O_1795,N_14223,N_13516);
and UO_1796 (O_1796,N_14963,N_13900);
nor UO_1797 (O_1797,N_14081,N_13871);
nand UO_1798 (O_1798,N_13907,N_13954);
xor UO_1799 (O_1799,N_13916,N_14740);
nor UO_1800 (O_1800,N_13890,N_14683);
nand UO_1801 (O_1801,N_13601,N_14915);
nand UO_1802 (O_1802,N_14466,N_14220);
nor UO_1803 (O_1803,N_14279,N_13579);
nand UO_1804 (O_1804,N_13505,N_13608);
and UO_1805 (O_1805,N_13672,N_14022);
or UO_1806 (O_1806,N_13753,N_13834);
nor UO_1807 (O_1807,N_13504,N_13887);
and UO_1808 (O_1808,N_14791,N_13579);
and UO_1809 (O_1809,N_14722,N_13999);
xor UO_1810 (O_1810,N_14787,N_14829);
nor UO_1811 (O_1811,N_14121,N_14144);
nor UO_1812 (O_1812,N_14366,N_14413);
nand UO_1813 (O_1813,N_14824,N_14276);
nor UO_1814 (O_1814,N_14559,N_14823);
and UO_1815 (O_1815,N_14295,N_14588);
xor UO_1816 (O_1816,N_14629,N_14732);
and UO_1817 (O_1817,N_14510,N_14991);
nand UO_1818 (O_1818,N_14473,N_14901);
nand UO_1819 (O_1819,N_14161,N_14007);
and UO_1820 (O_1820,N_14902,N_13768);
or UO_1821 (O_1821,N_14473,N_13543);
nand UO_1822 (O_1822,N_14738,N_13821);
nand UO_1823 (O_1823,N_13534,N_14826);
and UO_1824 (O_1824,N_13878,N_14473);
nand UO_1825 (O_1825,N_13958,N_13617);
nand UO_1826 (O_1826,N_14279,N_14424);
nand UO_1827 (O_1827,N_13814,N_13542);
nor UO_1828 (O_1828,N_14148,N_13601);
nand UO_1829 (O_1829,N_14260,N_14782);
xnor UO_1830 (O_1830,N_13881,N_14851);
nor UO_1831 (O_1831,N_14576,N_14455);
nand UO_1832 (O_1832,N_13748,N_14228);
nand UO_1833 (O_1833,N_14419,N_13746);
nand UO_1834 (O_1834,N_14342,N_14614);
and UO_1835 (O_1835,N_14602,N_14854);
nand UO_1836 (O_1836,N_14510,N_14457);
and UO_1837 (O_1837,N_13601,N_14929);
and UO_1838 (O_1838,N_14497,N_13938);
nand UO_1839 (O_1839,N_14285,N_14246);
and UO_1840 (O_1840,N_14917,N_14305);
nor UO_1841 (O_1841,N_14196,N_13745);
and UO_1842 (O_1842,N_14945,N_14799);
nor UO_1843 (O_1843,N_13896,N_14966);
nor UO_1844 (O_1844,N_14071,N_14637);
or UO_1845 (O_1845,N_14973,N_14763);
nand UO_1846 (O_1846,N_13709,N_14123);
and UO_1847 (O_1847,N_14007,N_14718);
nand UO_1848 (O_1848,N_13895,N_13896);
and UO_1849 (O_1849,N_13774,N_14339);
nor UO_1850 (O_1850,N_14954,N_13741);
or UO_1851 (O_1851,N_14334,N_14675);
nand UO_1852 (O_1852,N_13650,N_13813);
xnor UO_1853 (O_1853,N_14674,N_13756);
nand UO_1854 (O_1854,N_13968,N_13695);
xor UO_1855 (O_1855,N_14319,N_14452);
nor UO_1856 (O_1856,N_14389,N_13824);
or UO_1857 (O_1857,N_14427,N_14014);
nand UO_1858 (O_1858,N_14430,N_14143);
and UO_1859 (O_1859,N_13534,N_14884);
or UO_1860 (O_1860,N_14048,N_13875);
nor UO_1861 (O_1861,N_14574,N_14621);
and UO_1862 (O_1862,N_14692,N_14808);
and UO_1863 (O_1863,N_13512,N_13801);
nand UO_1864 (O_1864,N_14089,N_14244);
nor UO_1865 (O_1865,N_14260,N_14247);
xor UO_1866 (O_1866,N_13780,N_13620);
nor UO_1867 (O_1867,N_14959,N_14839);
and UO_1868 (O_1868,N_14287,N_14667);
or UO_1869 (O_1869,N_14879,N_14963);
nand UO_1870 (O_1870,N_14706,N_13965);
nand UO_1871 (O_1871,N_14437,N_14337);
or UO_1872 (O_1872,N_13594,N_14934);
nand UO_1873 (O_1873,N_14787,N_14626);
nand UO_1874 (O_1874,N_13602,N_14965);
and UO_1875 (O_1875,N_14908,N_14729);
or UO_1876 (O_1876,N_13713,N_14495);
and UO_1877 (O_1877,N_13812,N_13780);
xor UO_1878 (O_1878,N_14692,N_13619);
nor UO_1879 (O_1879,N_14711,N_14010);
or UO_1880 (O_1880,N_14651,N_13968);
nor UO_1881 (O_1881,N_13757,N_14512);
xor UO_1882 (O_1882,N_14938,N_13570);
nand UO_1883 (O_1883,N_14946,N_14185);
or UO_1884 (O_1884,N_14100,N_13534);
xor UO_1885 (O_1885,N_14041,N_14798);
and UO_1886 (O_1886,N_14731,N_13865);
nor UO_1887 (O_1887,N_14317,N_13685);
or UO_1888 (O_1888,N_14977,N_14882);
or UO_1889 (O_1889,N_14009,N_14699);
nor UO_1890 (O_1890,N_14882,N_14949);
or UO_1891 (O_1891,N_13549,N_13550);
and UO_1892 (O_1892,N_14651,N_14573);
or UO_1893 (O_1893,N_14353,N_13834);
and UO_1894 (O_1894,N_13932,N_14948);
or UO_1895 (O_1895,N_13734,N_13647);
and UO_1896 (O_1896,N_14132,N_14948);
nor UO_1897 (O_1897,N_14519,N_14390);
and UO_1898 (O_1898,N_14850,N_13526);
or UO_1899 (O_1899,N_13715,N_13635);
and UO_1900 (O_1900,N_14119,N_14887);
or UO_1901 (O_1901,N_14190,N_13648);
or UO_1902 (O_1902,N_14127,N_14691);
and UO_1903 (O_1903,N_14196,N_13965);
nor UO_1904 (O_1904,N_14515,N_14956);
xnor UO_1905 (O_1905,N_14536,N_13640);
xnor UO_1906 (O_1906,N_14654,N_13766);
or UO_1907 (O_1907,N_14595,N_13784);
nand UO_1908 (O_1908,N_14574,N_14012);
or UO_1909 (O_1909,N_14436,N_14767);
nor UO_1910 (O_1910,N_14000,N_14037);
and UO_1911 (O_1911,N_13609,N_14224);
and UO_1912 (O_1912,N_14250,N_13977);
nor UO_1913 (O_1913,N_13712,N_14360);
xnor UO_1914 (O_1914,N_14415,N_14098);
nor UO_1915 (O_1915,N_14283,N_13693);
nand UO_1916 (O_1916,N_14700,N_14470);
nand UO_1917 (O_1917,N_14347,N_13743);
nor UO_1918 (O_1918,N_14535,N_13690);
and UO_1919 (O_1919,N_13783,N_14977);
nand UO_1920 (O_1920,N_13784,N_14162);
nor UO_1921 (O_1921,N_13963,N_13580);
nor UO_1922 (O_1922,N_13621,N_14232);
nor UO_1923 (O_1923,N_13838,N_13974);
nand UO_1924 (O_1924,N_14120,N_14532);
or UO_1925 (O_1925,N_13869,N_14647);
nand UO_1926 (O_1926,N_14306,N_13519);
nor UO_1927 (O_1927,N_14256,N_14337);
nand UO_1928 (O_1928,N_13696,N_14621);
nor UO_1929 (O_1929,N_14903,N_14664);
or UO_1930 (O_1930,N_13826,N_14343);
nor UO_1931 (O_1931,N_13842,N_14275);
or UO_1932 (O_1932,N_13671,N_14387);
nand UO_1933 (O_1933,N_14527,N_14564);
nor UO_1934 (O_1934,N_14008,N_13810);
nor UO_1935 (O_1935,N_14635,N_14193);
or UO_1936 (O_1936,N_13913,N_13678);
nand UO_1937 (O_1937,N_13722,N_13796);
nand UO_1938 (O_1938,N_14340,N_14272);
xnor UO_1939 (O_1939,N_14363,N_14207);
nand UO_1940 (O_1940,N_14000,N_14976);
nand UO_1941 (O_1941,N_14385,N_14076);
and UO_1942 (O_1942,N_13679,N_13832);
nand UO_1943 (O_1943,N_14731,N_14126);
nor UO_1944 (O_1944,N_14571,N_14731);
nor UO_1945 (O_1945,N_13888,N_14918);
or UO_1946 (O_1946,N_13677,N_14908);
nand UO_1947 (O_1947,N_14271,N_14945);
nor UO_1948 (O_1948,N_14455,N_14422);
and UO_1949 (O_1949,N_14817,N_14155);
nor UO_1950 (O_1950,N_14834,N_13563);
nand UO_1951 (O_1951,N_14097,N_14803);
nand UO_1952 (O_1952,N_14989,N_14146);
nor UO_1953 (O_1953,N_14522,N_14032);
xnor UO_1954 (O_1954,N_14065,N_13659);
nand UO_1955 (O_1955,N_14894,N_14364);
nand UO_1956 (O_1956,N_14979,N_14466);
nand UO_1957 (O_1957,N_14624,N_14276);
and UO_1958 (O_1958,N_14997,N_14032);
nand UO_1959 (O_1959,N_13983,N_13670);
or UO_1960 (O_1960,N_14120,N_14320);
nand UO_1961 (O_1961,N_14978,N_14285);
nor UO_1962 (O_1962,N_14362,N_14218);
and UO_1963 (O_1963,N_14986,N_14466);
and UO_1964 (O_1964,N_14476,N_14319);
nor UO_1965 (O_1965,N_14060,N_14663);
or UO_1966 (O_1966,N_14283,N_13689);
and UO_1967 (O_1967,N_14723,N_14591);
nor UO_1968 (O_1968,N_13657,N_13800);
or UO_1969 (O_1969,N_14390,N_13560);
nor UO_1970 (O_1970,N_14507,N_14679);
nand UO_1971 (O_1971,N_13833,N_13832);
nor UO_1972 (O_1972,N_13955,N_14386);
or UO_1973 (O_1973,N_14537,N_14243);
xnor UO_1974 (O_1974,N_13622,N_14823);
nor UO_1975 (O_1975,N_14033,N_13624);
nor UO_1976 (O_1976,N_14608,N_13700);
nor UO_1977 (O_1977,N_13622,N_14689);
xnor UO_1978 (O_1978,N_14678,N_14980);
nor UO_1979 (O_1979,N_14320,N_13720);
nand UO_1980 (O_1980,N_14153,N_14669);
nand UO_1981 (O_1981,N_13615,N_14146);
nand UO_1982 (O_1982,N_14959,N_14286);
or UO_1983 (O_1983,N_13800,N_14694);
xor UO_1984 (O_1984,N_14688,N_14280);
and UO_1985 (O_1985,N_14411,N_14904);
and UO_1986 (O_1986,N_14682,N_14694);
nor UO_1987 (O_1987,N_13760,N_14430);
and UO_1988 (O_1988,N_13868,N_14830);
or UO_1989 (O_1989,N_13800,N_14920);
nand UO_1990 (O_1990,N_14254,N_13930);
or UO_1991 (O_1991,N_14268,N_14999);
nor UO_1992 (O_1992,N_14883,N_14291);
xor UO_1993 (O_1993,N_14784,N_13798);
nor UO_1994 (O_1994,N_13975,N_13627);
xnor UO_1995 (O_1995,N_14101,N_13885);
xnor UO_1996 (O_1996,N_14792,N_14383);
nand UO_1997 (O_1997,N_14986,N_14685);
or UO_1998 (O_1998,N_13576,N_13767);
and UO_1999 (O_1999,N_13608,N_14597);
endmodule