module basic_3000_30000_3500_5_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_1552,In_408);
or U1 (N_1,In_775,In_2959);
nor U2 (N_2,In_2230,In_69);
nand U3 (N_3,In_2141,In_2008);
nand U4 (N_4,In_1788,In_101);
nor U5 (N_5,In_2923,In_2796);
nor U6 (N_6,In_1791,In_710);
nor U7 (N_7,In_1012,In_584);
xnor U8 (N_8,In_2561,In_426);
xor U9 (N_9,In_1695,In_898);
nor U10 (N_10,In_171,In_2709);
and U11 (N_11,In_2397,In_981);
xnor U12 (N_12,In_2569,In_2202);
or U13 (N_13,In_83,In_2805);
nor U14 (N_14,In_1747,In_1795);
or U15 (N_15,In_1206,In_2079);
or U16 (N_16,In_2224,In_749);
and U17 (N_17,In_1245,In_2034);
xnor U18 (N_18,In_1323,In_60);
and U19 (N_19,In_1238,In_2045);
nor U20 (N_20,In_354,In_319);
nand U21 (N_21,In_890,In_64);
or U22 (N_22,In_1311,In_827);
nor U23 (N_23,In_429,In_1366);
or U24 (N_24,In_1852,In_2490);
and U25 (N_25,In_2904,In_1900);
or U26 (N_26,In_2739,In_869);
nor U27 (N_27,In_629,In_1251);
nand U28 (N_28,In_2924,In_2716);
and U29 (N_29,In_957,In_811);
or U30 (N_30,In_2506,In_2910);
xor U31 (N_31,In_624,In_352);
or U32 (N_32,In_1254,In_2591);
nor U33 (N_33,In_262,In_2855);
nor U34 (N_34,In_2846,In_282);
nor U35 (N_35,In_1765,In_2766);
nor U36 (N_36,In_2710,In_1225);
and U37 (N_37,In_1044,In_1588);
nand U38 (N_38,In_654,In_2121);
and U39 (N_39,In_1802,In_2654);
and U40 (N_40,In_2953,In_335);
and U41 (N_41,In_2936,In_125);
nand U42 (N_42,In_2351,In_2056);
nand U43 (N_43,In_1369,In_250);
nand U44 (N_44,In_1589,In_2930);
nor U45 (N_45,In_1689,In_1841);
nand U46 (N_46,In_615,In_2815);
nor U47 (N_47,In_1719,In_2961);
xnor U48 (N_48,In_1202,In_186);
or U49 (N_49,In_2195,In_216);
nor U50 (N_50,In_2852,In_1106);
xor U51 (N_51,In_1313,In_2279);
and U52 (N_52,In_882,In_2266);
and U53 (N_53,In_540,In_265);
and U54 (N_54,In_2402,In_2257);
xor U55 (N_55,In_2334,In_2154);
and U56 (N_56,In_1129,In_314);
nor U57 (N_57,In_2986,In_2577);
nor U58 (N_58,In_1616,In_2259);
xor U59 (N_59,In_1343,In_2782);
or U60 (N_60,In_505,In_2363);
nand U61 (N_61,In_2631,In_2164);
xnor U62 (N_62,In_512,In_2730);
or U63 (N_63,In_1718,In_2832);
nand U64 (N_64,In_2295,In_1091);
nand U65 (N_65,In_2851,In_2228);
xnor U66 (N_66,In_2160,In_557);
nand U67 (N_67,In_1836,In_1108);
nor U68 (N_68,In_233,In_1997);
nor U69 (N_69,In_1347,In_391);
or U70 (N_70,In_80,In_2450);
nor U71 (N_71,In_1723,In_658);
and U72 (N_72,In_90,In_1565);
and U73 (N_73,In_2774,In_338);
and U74 (N_74,In_1321,In_1391);
and U75 (N_75,In_2128,In_2408);
nand U76 (N_76,In_1069,In_2212);
or U77 (N_77,In_2773,In_1165);
xor U78 (N_78,In_2042,In_87);
or U79 (N_79,In_1601,In_1891);
nor U80 (N_80,In_1591,In_681);
and U81 (N_81,In_145,In_579);
or U82 (N_82,In_2401,In_107);
nand U83 (N_83,In_2482,In_247);
xor U84 (N_84,In_594,In_1410);
and U85 (N_85,In_1483,In_884);
or U86 (N_86,In_2179,In_643);
or U87 (N_87,In_1354,In_2229);
nand U88 (N_88,In_460,In_1965);
nor U89 (N_89,In_178,In_337);
and U90 (N_90,In_2542,In_565);
nor U91 (N_91,In_2433,In_2955);
nand U92 (N_92,In_2949,In_2248);
and U93 (N_93,In_1112,In_2338);
and U94 (N_94,In_1527,In_1444);
xor U95 (N_95,In_430,In_2013);
nand U96 (N_96,In_1966,In_2666);
or U97 (N_97,In_2557,In_1692);
or U98 (N_98,In_2349,In_2938);
and U99 (N_99,In_301,In_2153);
and U100 (N_100,In_2135,In_1503);
nand U101 (N_101,In_2918,In_721);
nor U102 (N_102,In_1549,In_2864);
nor U103 (N_103,In_183,In_2399);
nor U104 (N_104,In_1389,In_2052);
nand U105 (N_105,In_649,In_1574);
or U106 (N_106,In_238,In_745);
nand U107 (N_107,In_1412,In_672);
xnor U108 (N_108,In_1640,In_2607);
and U109 (N_109,In_2753,In_1083);
nor U110 (N_110,In_2734,In_1801);
and U111 (N_111,In_809,In_1385);
nand U112 (N_112,In_1631,In_2385);
nand U113 (N_113,In_2544,In_381);
and U114 (N_114,In_1517,In_1257);
nor U115 (N_115,In_2728,In_1660);
nor U116 (N_116,In_986,In_187);
or U117 (N_117,In_397,In_1865);
nand U118 (N_118,In_225,In_2817);
or U119 (N_119,In_2637,In_2995);
nand U120 (N_120,In_835,In_1538);
xnor U121 (N_121,In_1562,In_2795);
xnor U122 (N_122,In_2359,In_2198);
xor U123 (N_123,In_1162,In_872);
nand U124 (N_124,In_2346,In_2209);
nand U125 (N_125,In_2190,In_613);
or U126 (N_126,In_2092,In_2232);
or U127 (N_127,In_257,In_201);
xor U128 (N_128,In_824,In_1013);
xor U129 (N_129,In_815,In_2260);
nor U130 (N_130,In_2322,In_2458);
or U131 (N_131,In_1701,In_1994);
or U132 (N_132,In_2786,In_481);
and U133 (N_133,In_523,In_437);
nor U134 (N_134,In_756,In_205);
nand U135 (N_135,In_611,In_895);
or U136 (N_136,In_1330,In_1753);
xor U137 (N_137,In_1773,In_1744);
and U138 (N_138,In_2278,In_2388);
xor U139 (N_139,In_1636,In_398);
nor U140 (N_140,In_2593,In_1109);
and U141 (N_141,In_1397,In_581);
xnor U142 (N_142,In_1024,In_1009);
or U143 (N_143,In_2496,In_637);
and U144 (N_144,In_1693,In_1264);
and U145 (N_145,In_2847,In_2374);
and U146 (N_146,In_375,In_976);
and U147 (N_147,In_192,In_2438);
or U148 (N_148,In_2941,In_419);
xor U149 (N_149,In_683,In_1346);
and U150 (N_150,In_2174,In_1700);
and U151 (N_151,In_1134,In_2344);
and U152 (N_152,In_2800,In_1996);
or U153 (N_153,In_794,In_2810);
or U154 (N_154,In_2062,In_963);
or U155 (N_155,In_1702,In_1748);
nand U156 (N_156,In_1222,In_1688);
and U157 (N_157,In_2263,In_1668);
nand U158 (N_158,In_1992,In_2067);
nand U159 (N_159,In_1539,In_38);
xor U160 (N_160,In_1178,In_1957);
and U161 (N_161,In_1099,In_2777);
nand U162 (N_162,In_59,In_2811);
nand U163 (N_163,In_1945,In_2380);
nor U164 (N_164,In_2240,In_1156);
nor U165 (N_165,In_1087,In_830);
nand U166 (N_166,In_2389,In_2188);
xnor U167 (N_167,In_1819,In_1644);
nor U168 (N_168,In_2614,In_1821);
or U169 (N_169,In_1460,In_243);
xor U170 (N_170,In_1886,In_742);
or U171 (N_171,In_2732,In_2724);
or U172 (N_172,In_1405,In_1734);
nor U173 (N_173,In_1512,In_2479);
nand U174 (N_174,In_2481,In_2601);
nor U175 (N_175,In_1316,In_1642);
and U176 (N_176,In_2306,In_2406);
and U177 (N_177,In_1058,In_2199);
and U178 (N_178,In_2100,In_2533);
or U179 (N_179,In_2030,In_1356);
and U180 (N_180,In_170,In_1256);
or U181 (N_181,In_1671,In_96);
nor U182 (N_182,In_2894,In_266);
xor U183 (N_183,In_1486,In_2510);
nand U184 (N_184,In_2234,In_2831);
nor U185 (N_185,In_1745,In_2933);
xor U186 (N_186,In_1741,In_2221);
and U187 (N_187,In_212,In_610);
nor U188 (N_188,In_932,In_274);
nor U189 (N_189,In_256,In_340);
nand U190 (N_190,In_25,In_2973);
nor U191 (N_191,In_2435,In_1095);
nand U192 (N_192,In_1000,In_1426);
and U193 (N_193,In_2583,In_2527);
nand U194 (N_194,In_2524,In_2634);
nor U195 (N_195,In_1414,In_22);
xnor U196 (N_196,In_2116,In_1501);
and U197 (N_197,In_731,In_1573);
nor U198 (N_198,In_1423,In_150);
or U199 (N_199,In_893,In_2405);
nand U200 (N_200,In_2391,In_1203);
nor U201 (N_201,In_2083,In_1577);
xnor U202 (N_202,In_934,In_1157);
xor U203 (N_203,In_1011,In_312);
xnor U204 (N_204,In_1510,In_387);
or U205 (N_205,In_1492,In_1319);
or U206 (N_206,In_1951,In_191);
and U207 (N_207,In_2350,In_878);
nand U208 (N_208,In_29,In_1384);
or U209 (N_209,In_2792,In_1296);
or U210 (N_210,In_2778,In_1285);
xnor U211 (N_211,In_940,In_1986);
and U212 (N_212,In_120,In_577);
nor U213 (N_213,In_2589,In_26);
or U214 (N_214,In_2967,In_1059);
or U215 (N_215,In_1300,In_5);
nor U216 (N_216,In_133,In_2017);
and U217 (N_217,In_966,In_2403);
nor U218 (N_218,In_871,In_2468);
xnor U219 (N_219,In_1533,In_1046);
or U220 (N_220,In_147,In_907);
nand U221 (N_221,In_867,In_908);
nand U222 (N_222,In_676,In_2371);
xnor U223 (N_223,In_2485,In_2537);
xor U224 (N_224,In_2144,In_1694);
xnor U225 (N_225,In_1553,In_2964);
nor U226 (N_226,In_328,In_2844);
nor U227 (N_227,In_1709,In_172);
or U228 (N_228,In_1567,In_635);
nor U229 (N_229,In_2685,In_678);
nand U230 (N_230,In_595,In_355);
or U231 (N_231,In_2898,In_2222);
and U232 (N_232,In_1793,In_1943);
nor U233 (N_233,In_772,In_2020);
nor U234 (N_234,In_2097,In_1131);
or U235 (N_235,In_1635,In_1895);
nand U236 (N_236,In_933,In_2422);
or U237 (N_237,In_42,In_628);
or U238 (N_238,In_1955,In_1430);
or U239 (N_239,In_2578,In_2860);
nand U240 (N_240,In_630,In_1164);
or U241 (N_241,In_331,In_2281);
or U242 (N_242,In_1602,In_776);
nor U243 (N_243,In_290,In_740);
xnor U244 (N_244,In_1449,In_2563);
and U245 (N_245,In_1094,In_121);
nand U246 (N_246,In_1896,In_982);
or U247 (N_247,In_2297,In_1828);
nand U248 (N_248,In_2980,In_11);
nor U249 (N_249,In_1085,In_1546);
xnor U250 (N_250,In_1172,In_313);
xor U251 (N_251,In_558,In_2090);
nor U252 (N_252,In_1357,In_1055);
nand U253 (N_253,In_2797,In_747);
xor U254 (N_254,In_1580,In_1931);
or U255 (N_255,In_200,In_2241);
or U256 (N_256,In_1732,In_356);
and U257 (N_257,In_1839,In_1278);
nand U258 (N_258,In_1142,In_1089);
nor U259 (N_259,In_1267,In_2515);
xor U260 (N_260,In_894,In_2880);
nand U261 (N_261,In_999,In_2893);
xor U262 (N_262,In_929,In_2623);
nor U263 (N_263,In_2977,In_652);
and U264 (N_264,In_10,In_1542);
and U265 (N_265,In_1736,In_727);
nor U266 (N_266,In_1604,In_2075);
and U267 (N_267,In_1715,In_488);
nand U268 (N_268,In_2663,In_1757);
xnor U269 (N_269,In_539,In_1863);
nand U270 (N_270,In_675,In_655);
and U271 (N_271,In_2615,In_1246);
nand U272 (N_272,In_1376,In_2719);
nor U273 (N_273,In_2095,In_1353);
nor U274 (N_274,In_1790,In_547);
nand U275 (N_275,In_2437,In_805);
xnor U276 (N_276,In_2084,In_1842);
nand U277 (N_277,In_126,In_2000);
or U278 (N_278,In_164,In_2721);
xor U279 (N_279,In_1958,In_1678);
xor U280 (N_280,In_2197,In_2501);
nor U281 (N_281,In_1440,In_332);
xor U282 (N_282,In_2798,In_2512);
and U283 (N_283,In_1607,In_850);
nand U284 (N_284,In_1811,In_57);
nor U285 (N_285,In_228,In_2249);
nand U286 (N_286,In_1088,In_1283);
or U287 (N_287,In_1023,In_1073);
nand U288 (N_288,In_1787,In_816);
nand U289 (N_289,In_1443,In_1864);
and U290 (N_290,In_21,In_1505);
or U291 (N_291,In_2413,In_1208);
or U292 (N_292,In_1594,In_2142);
and U293 (N_293,In_1010,In_777);
xor U294 (N_294,In_1808,In_1956);
xor U295 (N_295,In_1402,In_2304);
nand U296 (N_296,In_1455,In_2236);
and U297 (N_297,In_2219,In_2504);
xor U298 (N_298,In_267,In_2856);
nand U299 (N_299,In_226,In_369);
nand U300 (N_300,In_1703,In_2101);
nand U301 (N_301,In_1673,In_779);
nand U302 (N_302,In_2047,In_2518);
and U303 (N_303,In_153,In_2627);
and U304 (N_304,In_2319,In_1663);
or U305 (N_305,In_881,In_2985);
xnor U306 (N_306,In_1603,In_665);
nand U307 (N_307,In_1868,In_1239);
nand U308 (N_308,In_1328,In_2169);
nand U309 (N_309,In_1596,In_2963);
or U310 (N_310,In_707,In_2550);
and U311 (N_311,In_2731,In_971);
xnor U312 (N_312,In_2655,In_2091);
xnor U313 (N_313,In_2760,In_1698);
nor U314 (N_314,In_728,In_1163);
nor U315 (N_315,In_2088,In_2046);
nor U316 (N_316,In_2011,In_2168);
or U317 (N_317,In_1447,In_2184);
xnor U318 (N_318,In_466,In_489);
or U319 (N_319,In_964,In_2282);
and U320 (N_320,In_946,In_833);
nand U321 (N_321,In_1027,In_2929);
and U322 (N_322,In_694,In_2036);
or U323 (N_323,In_325,In_295);
nand U324 (N_324,In_996,In_263);
nand U325 (N_325,In_2521,In_1248);
and U326 (N_326,In_1092,In_2261);
and U327 (N_327,In_464,In_660);
and U328 (N_328,In_2919,In_1775);
or U329 (N_329,In_717,In_1530);
or U330 (N_330,In_795,In_1479);
nor U331 (N_331,In_468,In_1439);
or U332 (N_332,In_1071,In_2425);
and U333 (N_333,In_2744,In_2992);
nor U334 (N_334,In_602,In_249);
or U335 (N_335,In_1261,In_2684);
and U336 (N_336,In_1817,In_1471);
and U337 (N_337,In_2635,In_75);
nor U338 (N_338,In_2837,In_457);
nor U339 (N_339,In_2451,In_807);
nand U340 (N_340,In_2722,In_2911);
nor U341 (N_341,In_2983,In_2843);
xnor U342 (N_342,In_1597,In_1298);
or U343 (N_343,In_2806,In_2386);
or U344 (N_344,In_403,In_1103);
xor U345 (N_345,In_2447,In_729);
nand U346 (N_346,In_2947,In_1712);
or U347 (N_347,In_545,In_2010);
and U348 (N_348,In_2838,In_2393);
nor U349 (N_349,In_700,In_1525);
xor U350 (N_350,In_1626,In_1595);
nand U351 (N_351,In_2839,In_2769);
nand U352 (N_352,In_2147,In_2493);
xnor U353 (N_353,In_2492,In_2429);
nand U354 (N_354,In_1560,In_2455);
or U355 (N_355,In_1432,In_1054);
nor U356 (N_356,In_253,In_497);
and U357 (N_357,In_968,In_2368);
and U358 (N_358,In_2177,In_2816);
nor U359 (N_359,In_166,In_1335);
or U360 (N_360,In_115,In_808);
or U361 (N_361,In_1262,In_1104);
or U362 (N_362,In_2874,In_689);
xnor U363 (N_363,In_2982,In_767);
and U364 (N_364,In_65,In_56);
nand U365 (N_365,In_2511,In_852);
nor U366 (N_366,In_2625,In_1643);
or U367 (N_367,In_1329,In_2794);
or U368 (N_368,In_715,In_774);
or U369 (N_369,In_318,In_2531);
xnor U370 (N_370,In_942,In_1535);
and U371 (N_371,In_716,In_917);
or U372 (N_372,In_2300,In_280);
xor U373 (N_373,In_2891,In_2957);
nand U374 (N_374,In_1143,In_1491);
nand U375 (N_375,In_124,In_1659);
nand U376 (N_376,In_1875,In_2361);
or U377 (N_377,In_157,In_2476);
and U378 (N_378,In_2061,In_2252);
or U379 (N_379,In_1854,In_451);
nand U380 (N_380,In_1537,In_2106);
xor U381 (N_381,In_1777,In_904);
or U382 (N_382,In_1252,In_555);
or U383 (N_383,In_251,In_1504);
or U384 (N_384,In_1170,In_443);
or U385 (N_385,In_1666,In_1381);
nor U386 (N_386,In_2421,In_1566);
or U387 (N_387,In_203,In_1799);
or U388 (N_388,In_347,In_84);
nor U389 (N_389,In_2896,In_1062);
nor U390 (N_390,In_1291,In_708);
or U391 (N_391,In_2137,In_360);
nand U392 (N_392,In_1302,In_1665);
or U393 (N_393,In_2867,In_394);
nor U394 (N_394,In_1998,In_2662);
or U395 (N_395,In_2002,In_1282);
xor U396 (N_396,In_82,In_568);
nor U397 (N_397,In_2581,In_405);
nand U398 (N_398,In_718,In_2376);
xnor U399 (N_399,In_2089,In_1196);
and U400 (N_400,In_308,In_2284);
nor U401 (N_401,In_2159,In_1870);
or U402 (N_402,In_1185,In_2431);
or U403 (N_403,In_1060,In_1758);
and U404 (N_404,In_972,In_1582);
xor U405 (N_405,In_2922,In_149);
nand U406 (N_406,In_1242,In_958);
xor U407 (N_407,In_2579,In_1590);
nand U408 (N_408,In_2348,In_255);
xnor U409 (N_409,In_1968,In_1434);
or U410 (N_410,In_955,In_1287);
or U411 (N_411,In_1217,In_1789);
or U412 (N_412,In_784,In_483);
and U413 (N_413,In_1331,In_1794);
nand U414 (N_414,In_1770,In_193);
or U415 (N_415,In_2277,In_2672);
and U416 (N_416,In_47,In_1524);
or U417 (N_417,In_2801,In_1128);
xor U418 (N_418,In_889,In_2283);
and U419 (N_419,In_736,In_826);
nor U420 (N_420,In_1326,In_2331);
nand U421 (N_421,In_494,In_161);
nor U422 (N_422,In_1212,In_902);
nand U423 (N_423,In_2328,In_977);
and U424 (N_424,In_2019,In_1684);
and U425 (N_425,In_2342,In_2661);
nor U426 (N_426,In_1834,In_603);
and U427 (N_427,In_2446,In_2937);
and U428 (N_428,In_2733,In_2701);
or U429 (N_429,In_642,In_2939);
and U430 (N_430,In_1395,In_2616);
or U431 (N_431,In_693,In_832);
xnor U432 (N_432,In_661,In_303);
nand U433 (N_433,In_1547,In_1180);
xnor U434 (N_434,In_1738,In_2823);
nor U435 (N_435,In_2649,In_99);
nor U436 (N_436,In_1141,In_2339);
and U437 (N_437,In_2993,In_2119);
or U438 (N_438,In_2314,In_536);
nand U439 (N_439,In_2469,In_1976);
xor U440 (N_440,In_983,In_130);
and U441 (N_441,In_1314,In_1379);
nor U442 (N_442,In_905,In_1872);
xnor U443 (N_443,In_1639,In_813);
and U444 (N_444,In_1127,In_1428);
and U445 (N_445,In_1920,In_2237);
xnor U446 (N_446,In_2560,In_551);
xor U447 (N_447,In_350,In_1457);
xnor U448 (N_448,In_353,In_2271);
nand U449 (N_449,In_2657,In_73);
or U450 (N_450,In_1883,In_1615);
nor U451 (N_451,In_1598,In_991);
xnor U452 (N_452,In_1076,In_1493);
or U453 (N_453,In_2364,In_1482);
nor U454 (N_454,In_1605,In_1362);
xor U455 (N_455,In_2044,In_839);
nor U456 (N_456,In_2785,In_1559);
or U457 (N_457,In_1396,In_1056);
or U458 (N_458,In_563,In_2396);
or U459 (N_459,In_2747,In_2706);
nand U460 (N_460,In_1214,In_1725);
or U461 (N_461,In_897,In_1324);
xnor U462 (N_462,In_634,In_1531);
xnor U463 (N_463,In_2804,In_1761);
nand U464 (N_464,In_1276,In_2);
or U465 (N_465,In_1583,In_1950);
nand U466 (N_466,In_2238,In_2610);
and U467 (N_467,In_657,In_1407);
or U468 (N_468,In_2807,In_261);
and U469 (N_469,In_1080,In_2650);
or U470 (N_470,In_1617,In_2070);
or U471 (N_471,In_2575,In_287);
nor U472 (N_472,In_362,In_2185);
or U473 (N_473,In_412,In_173);
and U474 (N_474,In_2862,In_2016);
nor U475 (N_475,In_778,In_324);
nand U476 (N_476,In_2671,In_623);
and U477 (N_477,In_2183,In_44);
xor U478 (N_478,In_1610,In_2580);
and U479 (N_479,In_2203,In_384);
nor U480 (N_480,In_1942,In_632);
and U481 (N_481,In_2568,In_1030);
nor U482 (N_482,In_2480,In_1911);
xnor U483 (N_483,In_639,In_2419);
xor U484 (N_484,In_349,In_1520);
xor U485 (N_485,In_1048,In_825);
and U486 (N_486,In_2660,In_2265);
nor U487 (N_487,In_1614,In_1004);
or U488 (N_488,In_2473,In_781);
or U489 (N_489,In_1277,In_947);
xnor U490 (N_490,In_2704,In_670);
nor U491 (N_491,In_651,In_1498);
xor U492 (N_492,In_591,In_662);
nand U493 (N_493,In_414,In_1686);
and U494 (N_494,In_561,In_39);
nand U495 (N_495,In_724,In_341);
nand U496 (N_496,In_485,In_1915);
nand U497 (N_497,In_2695,In_1892);
xnor U498 (N_498,In_664,In_1954);
nand U499 (N_499,In_1848,In_2094);
and U500 (N_500,In_1377,In_703);
xnor U501 (N_501,In_713,In_2166);
nand U502 (N_502,In_844,In_2771);
nand U503 (N_503,In_2107,In_1200);
xnor U504 (N_504,In_239,In_2598);
or U505 (N_505,In_679,In_2167);
xor U506 (N_506,In_2384,In_520);
or U507 (N_507,In_773,In_1053);
or U508 (N_508,In_1980,In_901);
nand U509 (N_509,In_723,In_1473);
nand U510 (N_510,In_411,In_455);
or U511 (N_511,In_196,In_1105);
nor U512 (N_512,In_875,In_420);
nor U513 (N_513,In_2756,In_2115);
nand U514 (N_514,In_2656,In_2445);
and U515 (N_515,In_1767,In_1554);
xor U516 (N_516,In_2841,In_479);
and U517 (N_517,In_2471,In_2256);
or U518 (N_518,In_1940,In_2576);
nor U519 (N_519,In_1189,In_2516);
nor U520 (N_520,In_685,In_873);
and U521 (N_521,In_589,In_1806);
nor U522 (N_522,In_2758,In_2848);
xnor U523 (N_523,In_1456,In_2741);
nor U524 (N_524,In_111,In_2943);
xor U525 (N_525,In_2617,In_2270);
nand U526 (N_526,In_1348,In_1184);
nor U527 (N_527,In_49,In_1993);
nor U528 (N_528,In_969,In_2602);
nand U529 (N_529,In_837,In_2900);
nand U530 (N_530,In_962,In_572);
xor U531 (N_531,In_725,In_469);
xor U532 (N_532,In_2600,In_622);
nand U533 (N_533,In_1052,In_1146);
nor U534 (N_534,In_2307,In_2629);
nand U535 (N_535,In_1228,In_2976);
xnor U536 (N_536,In_519,In_526);
or U537 (N_537,In_1823,In_2157);
and U538 (N_538,In_407,In_2658);
xor U539 (N_539,In_1477,In_364);
and U540 (N_540,In_0,In_2545);
and U541 (N_541,In_1754,In_2054);
xor U542 (N_542,In_1878,In_790);
nand U543 (N_543,In_2194,In_1392);
nor U544 (N_544,In_2031,In_2329);
nor U545 (N_545,In_599,In_2783);
or U546 (N_546,In_2311,In_151);
or U547 (N_547,In_1973,In_614);
nor U548 (N_548,In_677,In_2665);
xor U549 (N_549,In_2503,In_2987);
xnor U550 (N_550,In_2633,In_1514);
nand U551 (N_551,In_231,In_1962);
nor U552 (N_552,In_2098,In_220);
nor U553 (N_553,In_2039,In_386);
nand U554 (N_554,In_1101,In_2621);
nor U555 (N_555,In_33,In_1630);
and U556 (N_556,In_2522,In_363);
xor U557 (N_557,In_1880,In_1273);
or U558 (N_558,In_1241,In_1327);
or U559 (N_559,In_1265,In_1809);
xnor U560 (N_560,In_686,In_1341);
or U561 (N_561,In_1031,In_2225);
nand U562 (N_562,In_2436,In_2849);
nor U563 (N_563,In_447,In_2032);
and U564 (N_564,In_272,In_2155);
xnor U565 (N_565,In_1067,In_2309);
xnor U566 (N_566,In_346,In_58);
nor U567 (N_567,In_938,In_1959);
and U568 (N_568,In_2233,In_2427);
nor U569 (N_569,In_2752,In_2049);
nor U570 (N_570,In_242,In_2564);
or U571 (N_571,In_993,In_1778);
or U572 (N_572,In_390,In_2004);
xor U573 (N_573,In_417,In_1953);
xor U574 (N_574,In_527,In_53);
and U575 (N_575,In_2173,In_617);
xnor U576 (N_576,In_2373,In_2928);
nor U577 (N_577,In_155,In_1413);
nand U578 (N_578,In_590,In_1484);
xnor U579 (N_579,In_1687,In_2776);
nand U580 (N_580,In_2305,In_2907);
nor U581 (N_581,In_2041,In_2285);
xnor U582 (N_582,In_1268,In_1042);
or U583 (N_583,In_2337,In_1064);
and U584 (N_584,In_1970,In_70);
and U585 (N_585,In_2268,In_1967);
and U586 (N_586,In_292,In_549);
nor U587 (N_587,In_307,In_2347);
and U588 (N_588,In_2746,In_2651);
or U589 (N_589,In_1798,In_1881);
nor U590 (N_590,In_900,In_1825);
nor U591 (N_591,In_2740,In_2392);
or U592 (N_592,In_2999,In_27);
xnor U593 (N_593,In_1908,In_754);
or U594 (N_594,In_24,In_2387);
nor U595 (N_595,In_587,In_382);
nor U596 (N_596,In_2033,In_1037);
nor U597 (N_597,In_1213,In_2833);
and U598 (N_598,In_1174,In_1051);
or U599 (N_599,In_2390,In_1084);
xor U600 (N_600,In_1318,In_2077);
or U601 (N_601,In_66,In_2291);
and U602 (N_602,In_2877,In_480);
nand U603 (N_603,In_103,In_1867);
xor U604 (N_604,In_2432,In_618);
or U605 (N_605,In_2597,In_1);
xor U606 (N_606,In_918,In_915);
xnor U607 (N_607,In_237,In_525);
nand U608 (N_608,In_1132,In_1846);
nor U609 (N_609,In_2472,In_554);
nor U610 (N_610,In_1082,In_2245);
nor U611 (N_611,In_2357,In_1496);
xor U612 (N_612,In_2883,In_692);
nor U613 (N_613,In_2178,In_1137);
or U614 (N_614,In_348,In_1057);
and U615 (N_615,In_385,In_221);
or U616 (N_616,In_2854,In_2069);
nand U617 (N_617,In_698,In_2876);
and U618 (N_618,In_682,In_1107);
or U619 (N_619,In_36,In_788);
nor U620 (N_620,In_1193,In_1662);
xnor U621 (N_621,In_2680,In_1608);
and U622 (N_622,In_769,In_2486);
nor U623 (N_623,In_323,In_102);
or U624 (N_624,In_230,In_1295);
and U625 (N_625,In_486,In_104);
xor U626 (N_626,In_719,In_477);
nand U627 (N_627,In_2356,In_2381);
nand U628 (N_628,In_2958,In_2821);
xor U629 (N_629,In_949,In_176);
nor U630 (N_630,In_1086,In_2921);
or U631 (N_631,In_2514,In_2038);
xor U632 (N_632,In_1522,In_858);
and U633 (N_633,In_2587,In_1495);
or U634 (N_634,In_416,In_1303);
nand U635 (N_635,In_516,In_298);
or U636 (N_636,In_1974,In_2333);
nand U637 (N_637,In_179,In_2175);
and U638 (N_638,In_1373,In_2738);
xnor U639 (N_639,In_2824,In_2592);
or U640 (N_640,In_1890,In_1018);
or U641 (N_641,In_1415,In_2235);
nor U642 (N_642,In_1850,In_1721);
nand U643 (N_643,In_892,In_1181);
and U644 (N_644,In_691,In_1047);
or U645 (N_645,In_1857,In_1333);
nor U646 (N_646,In_1985,In_2647);
nor U647 (N_647,In_640,In_400);
or U648 (N_648,In_2463,In_2726);
nand U649 (N_649,In_2382,In_797);
or U650 (N_650,In_1451,In_156);
nor U651 (N_651,In_2736,In_1509);
and U652 (N_652,In_2156,In_2808);
and U653 (N_653,In_739,In_1628);
or U654 (N_654,In_2763,In_2780);
xnor U655 (N_655,In_2541,In_1450);
xor U656 (N_656,In_606,In_2683);
xor U657 (N_657,In_2086,In_765);
and U658 (N_658,In_2632,In_1783);
xor U659 (N_659,In_1036,In_559);
nor U660 (N_660,In_1194,In_2055);
nand U661 (N_661,In_1914,In_2462);
nor U662 (N_662,In_383,In_1874);
or U663 (N_663,In_1280,In_108);
nand U664 (N_664,In_2430,In_2335);
xnor U665 (N_665,In_1680,In_366);
nand U666 (N_666,In_1894,In_2288);
xnor U667 (N_667,In_2878,In_2417);
xor U668 (N_668,In_2951,In_1065);
xor U669 (N_669,In_1730,In_785);
and U670 (N_670,In_1759,In_1126);
and U671 (N_671,In_1987,In_1115);
and U672 (N_672,In_1726,In_2692);
nor U673 (N_673,In_2573,In_1461);
and U674 (N_674,In_2791,In_2254);
xnor U675 (N_675,In_2646,In_1877);
xnor U676 (N_676,In_647,In_2151);
nand U677 (N_677,In_1147,In_1576);
and U678 (N_678,In_140,In_493);
nand U679 (N_679,In_1814,In_41);
xor U680 (N_680,In_2588,In_286);
and U681 (N_681,In_528,In_2372);
nand U682 (N_682,In_2689,In_2505);
nand U683 (N_683,In_94,In_2915);
and U684 (N_684,In_2916,In_1960);
nand U685 (N_685,In_2085,In_1928);
nand U686 (N_686,In_1835,In_518);
or U687 (N_687,In_1130,In_449);
xor U688 (N_688,In_1551,In_264);
and U689 (N_689,In_2192,In_1079);
or U690 (N_690,In_1469,In_2302);
xnor U691 (N_691,In_1930,In_1627);
xor U692 (N_692,In_667,In_1435);
or U693 (N_693,In_802,In_2324);
or U694 (N_694,In_849,In_76);
or U695 (N_695,In_1480,In_2273);
xor U696 (N_696,In_2749,In_2962);
nor U697 (N_697,In_798,In_206);
nand U698 (N_698,In_2415,In_2781);
nor U699 (N_699,In_1507,In_1236);
xnor U700 (N_700,In_829,In_2946);
or U701 (N_701,In_284,In_2676);
or U702 (N_702,In_1796,In_2822);
nor U703 (N_703,In_78,In_2909);
or U704 (N_704,In_1829,In_2218);
or U705 (N_705,In_1215,In_2714);
and U706 (N_706,In_702,In_1979);
nand U707 (N_707,In_1187,In_515);
nand U708 (N_708,In_529,In_1478);
or U709 (N_709,In_848,In_40);
and U710 (N_710,In_1714,In_586);
xor U711 (N_711,In_733,In_2014);
xor U712 (N_712,In_1648,In_329);
and U713 (N_713,In_2711,In_1177);
and U714 (N_714,In_2819,In_1679);
and U715 (N_715,In_1437,In_215);
or U716 (N_716,In_2132,In_1145);
and U717 (N_717,In_1229,In_2507);
xnor U718 (N_718,In_388,In_1699);
nand U719 (N_719,In_1843,In_2718);
and U720 (N_720,In_68,In_758);
nor U721 (N_721,In_1305,In_1074);
xnor U722 (N_722,In_2870,In_2605);
or U723 (N_723,In_1912,In_513);
nor U724 (N_724,In_2125,In_841);
nand U725 (N_725,In_291,In_1292);
or U726 (N_726,In_2158,In_48);
nor U727 (N_727,In_2426,In_2024);
or U728 (N_728,In_2751,In_1370);
and U729 (N_729,In_2444,In_2723);
or U730 (N_730,In_861,In_1197);
nand U731 (N_731,In_1532,In_2772);
xor U732 (N_732,In_2200,In_1233);
and U733 (N_733,In_521,In_845);
nand U734 (N_734,In_2443,In_1035);
nor U735 (N_735,In_1800,In_2926);
nor U736 (N_736,In_2063,In_1223);
xor U737 (N_737,In_439,In_1521);
and U738 (N_738,In_1816,In_2139);
xor U739 (N_739,In_463,In_165);
xor U740 (N_740,In_456,In_2035);
xor U741 (N_741,In_2836,In_2975);
and U742 (N_742,In_985,In_2978);
nand U743 (N_743,In_1400,In_1269);
nor U744 (N_744,In_926,In_2562);
nand U745 (N_745,In_863,In_2294);
or U746 (N_746,In_656,In_607);
xor U747 (N_747,In_973,In_2250);
and U748 (N_748,In_1306,In_1199);
nand U749 (N_749,In_2935,In_434);
or U750 (N_750,In_2483,In_1188);
or U751 (N_751,In_1155,In_1981);
xnor U752 (N_752,In_1016,In_533);
or U753 (N_753,In_1116,In_441);
nand U754 (N_754,In_210,In_552);
or U755 (N_755,In_2176,In_2764);
or U756 (N_756,In_1288,In_753);
and U757 (N_757,In_1481,In_2196);
xor U758 (N_758,In_1653,In_2096);
nand U759 (N_759,In_2470,In_2585);
and U760 (N_760,In_37,In_1349);
nor U761 (N_761,In_2532,In_2636);
or U762 (N_762,In_1459,In_2713);
xor U763 (N_763,In_163,In_831);
and U764 (N_764,In_2080,In_2950);
xnor U765 (N_765,In_1453,In_1244);
or U766 (N_766,In_936,In_2280);
xor U767 (N_767,In_1536,In_1632);
xor U768 (N_768,In_1139,In_259);
nand U769 (N_769,In_368,In_859);
xnor U770 (N_770,In_2696,In_244);
or U771 (N_771,In_2182,In_380);
or U772 (N_772,In_2863,In_1952);
nand U773 (N_773,In_2316,In_1465);
nand U774 (N_774,In_1171,In_1740);
xor U775 (N_775,In_2336,In_2948);
and U776 (N_776,In_2912,In_766);
xnor U777 (N_777,In_1364,In_2110);
or U778 (N_778,In_234,In_1258);
nor U779 (N_779,In_1097,In_1613);
nand U780 (N_780,In_2673,In_2027);
xnor U781 (N_781,In_1338,In_1383);
xnor U782 (N_782,In_761,In_1166);
nor U783 (N_783,In_160,In_548);
and U784 (N_784,In_473,In_1022);
nor U785 (N_785,In_1682,In_320);
or U786 (N_786,In_1216,In_2565);
and U787 (N_787,In_168,In_1063);
nand U788 (N_788,In_1792,In_1933);
xnor U789 (N_789,In_1408,In_159);
and U790 (N_790,In_2996,In_365);
nor U791 (N_791,In_913,In_1923);
nor U792 (N_792,In_541,In_8);
nand U793 (N_793,In_2885,In_1971);
or U794 (N_794,In_2494,In_1149);
xor U795 (N_795,In_804,In_567);
xor U796 (N_796,In_1905,In_134);
and U797 (N_797,In_1609,In_1919);
nor U798 (N_798,In_1742,In_2136);
nand U799 (N_799,In_110,In_28);
xor U800 (N_800,In_2534,In_2551);
xor U801 (N_801,In_2220,In_2465);
nor U802 (N_802,In_2353,In_2081);
nor U803 (N_803,In_2082,In_2205);
or U804 (N_804,In_1681,In_2189);
or U805 (N_805,In_574,In_2775);
xor U806 (N_806,In_2186,In_2457);
and U807 (N_807,In_227,In_1876);
nand U808 (N_808,In_1209,In_596);
nand U809 (N_809,In_137,In_1367);
nand U810 (N_810,In_1893,In_496);
and U811 (N_811,In_714,In_570);
or U812 (N_812,In_1485,In_2835);
and U813 (N_813,In_294,In_213);
nand U814 (N_814,In_874,In_885);
nand U815 (N_815,In_1167,In_462);
or U816 (N_816,In_2879,In_1763);
xor U817 (N_817,In_1334,In_1342);
xnor U818 (N_818,In_2148,In_2858);
nand U819 (N_819,In_2076,In_1488);
nand U820 (N_820,In_1906,In_2050);
nor U821 (N_821,In_812,In_621);
nand U822 (N_822,In_2247,In_2813);
nor U823 (N_823,In_680,In_2640);
nor U824 (N_824,In_2475,In_4);
and U825 (N_825,In_1255,In_1490);
nand U826 (N_826,In_820,In_2866);
nand U827 (N_827,In_1409,In_669);
xor U828 (N_828,In_2608,In_931);
nand U829 (N_829,In_2466,In_1374);
xor U830 (N_830,In_1072,In_1849);
nor U831 (N_831,In_880,In_598);
and U832 (N_832,In_306,In_1690);
nor U833 (N_833,In_899,In_395);
and U834 (N_834,In_2497,In_1117);
xnor U835 (N_835,In_2513,In_1186);
xnor U836 (N_836,In_1122,In_177);
or U837 (N_837,In_2697,In_342);
nand U838 (N_838,In_2354,In_413);
xor U839 (N_839,In_2884,In_1387);
nand U840 (N_840,In_311,In_935);
or U841 (N_841,In_1403,In_1984);
nor U842 (N_842,In_732,In_2743);
nor U843 (N_843,In_2966,In_1641);
nand U844 (N_844,In_2029,In_2217);
or U845 (N_845,In_18,In_2554);
xor U846 (N_846,In_2789,In_326);
nor U847 (N_847,In_1308,In_1898);
nand U848 (N_848,In_2246,In_2694);
and U849 (N_849,In_276,In_2897);
xor U850 (N_850,In_309,In_843);
nand U851 (N_851,In_2418,In_2264);
xnor U852 (N_852,In_232,In_1847);
nand U853 (N_853,In_2407,In_2913);
nor U854 (N_854,In_223,In_866);
or U855 (N_855,In_2882,In_2326);
nor U856 (N_856,In_2133,In_2613);
and U857 (N_857,In_1077,In_1578);
or U858 (N_858,In_2691,In_726);
nor U859 (N_859,In_2286,In_975);
or U860 (N_860,In_928,In_2377);
nand U861 (N_861,In_1029,In_888);
and U862 (N_862,In_2688,In_2308);
xor U863 (N_863,In_2708,In_2187);
nor U864 (N_864,In_2301,In_438);
nand U865 (N_865,In_1339,In_1964);
or U866 (N_866,In_696,In_1768);
nor U867 (N_867,In_2509,In_1568);
and U868 (N_868,In_1002,In_277);
and U869 (N_869,In_2065,In_1393);
and U870 (N_870,In_268,In_1487);
xor U871 (N_871,In_1526,In_1475);
xnor U872 (N_872,In_1360,In_1275);
and U873 (N_873,In_2626,In_620);
or U874 (N_874,In_1380,In_2165);
nand U875 (N_875,In_2845,In_569);
and U876 (N_876,In_2355,In_674);
nor U877 (N_877,In_503,In_2123);
and U878 (N_878,In_2028,In_61);
xnor U879 (N_879,In_1049,In_452);
xnor U880 (N_880,In_2586,In_1885);
xor U881 (N_881,In_2216,In_990);
and U882 (N_882,In_357,In_2566);
nor U883 (N_883,In_52,In_1776);
nand U884 (N_884,In_77,In_241);
nor U885 (N_885,In_653,In_2720);
and U886 (N_886,In_1683,In_46);
nor U887 (N_887,In_699,In_2888);
xnor U888 (N_888,In_296,In_592);
and U889 (N_889,In_43,In_2068);
xor U890 (N_890,In_791,In_978);
and U891 (N_891,In_476,In_644);
nor U892 (N_892,In_1625,In_989);
and U893 (N_893,In_2037,In_370);
or U894 (N_894,In_914,In_743);
or U895 (N_895,In_491,In_20);
or U896 (N_896,In_1230,In_97);
and U897 (N_897,In_1999,In_690);
or U898 (N_898,In_2315,In_641);
or U899 (N_899,In_1003,In_2213);
nand U900 (N_900,In_289,In_1805);
nand U901 (N_901,In_1210,In_2001);
nand U902 (N_902,In_1118,In_2395);
and U903 (N_903,In_1090,In_402);
nand U904 (N_904,In_2681,In_2143);
or U905 (N_905,In_616,In_1654);
nor U906 (N_906,In_217,In_2784);
or U907 (N_907,In_1458,In_2276);
xor U908 (N_908,In_2619,In_1050);
and U909 (N_909,In_911,In_738);
xor U910 (N_910,In_2204,In_910);
nor U911 (N_911,In_393,In_1207);
nor U912 (N_912,In_2677,In_2064);
or U913 (N_913,In_2448,In_2111);
or U914 (N_914,In_2873,In_909);
or U915 (N_915,In_2765,In_2802);
nor U916 (N_916,In_143,In_1340);
nand U917 (N_917,In_275,In_2243);
or U918 (N_918,In_2005,In_1175);
nand U919 (N_919,In_1624,In_792);
or U920 (N_920,In_162,In_2679);
xnor U921 (N_921,In_939,In_2970);
xor U922 (N_922,In_787,In_1845);
nor U923 (N_923,In_514,In_2026);
nand U924 (N_924,In_1544,In_1934);
or U925 (N_925,In_142,In_1961);
xor U926 (N_926,In_1903,In_1516);
nand U927 (N_927,In_358,In_1871);
xor U928 (N_928,In_2994,In_465);
xor U929 (N_929,In_9,In_79);
and U930 (N_930,In_870,In_2299);
xnor U931 (N_931,In_1325,In_144);
nand U932 (N_932,In_2814,In_1224);
xor U933 (N_933,In_1889,In_1579);
xnor U934 (N_934,In_482,In_1211);
nand U935 (N_935,In_1438,In_2612);
nand U936 (N_936,In_269,In_376);
nand U937 (N_937,In_1148,In_1826);
nand U938 (N_938,In_2118,In_2767);
or U939 (N_939,In_13,In_2416);
nand U940 (N_940,In_508,In_1824);
and U941 (N_941,In_461,In_2499);
or U942 (N_942,In_1350,In_2539);
xnor U943 (N_943,In_2275,In_2715);
xnor U944 (N_944,In_1832,In_705);
and U945 (N_945,In_1833,In_1144);
nor U946 (N_946,In_50,In_2461);
xor U947 (N_947,In_522,In_442);
nor U948 (N_948,In_1810,In_2488);
nand U949 (N_949,In_2829,In_2595);
or U950 (N_950,In_2523,In_1158);
or U951 (N_951,In_1634,In_299);
and U952 (N_952,In_1807,In_2440);
nand U953 (N_953,In_1466,In_2321);
xnor U954 (N_954,In_2456,In_1837);
or U955 (N_955,In_974,In_2093);
nor U956 (N_956,In_945,In_605);
and U957 (N_957,In_2484,In_1110);
nor U958 (N_958,In_1421,In_2606);
or U959 (N_959,In_1812,In_2330);
or U960 (N_960,In_1669,In_2942);
or U961 (N_961,In_2686,In_1017);
and U962 (N_962,In_2369,In_980);
and U963 (N_963,In_474,In_1728);
xor U964 (N_964,In_2768,In_1474);
or U965 (N_965,In_1704,In_1183);
nand U966 (N_966,In_2231,In_2520);
or U967 (N_967,In_1028,In_472);
nor U968 (N_968,In_2303,In_190);
xnor U969 (N_969,In_789,In_2972);
and U970 (N_970,In_182,In_960);
nand U971 (N_971,In_1154,In_2886);
or U972 (N_972,In_2172,In_448);
xnor U973 (N_973,In_202,In_2664);
nand U974 (N_974,In_1581,In_2717);
nand U975 (N_975,In_1936,In_1926);
xor U976 (N_976,In_2495,In_937);
xor U977 (N_977,In_1873,In_2474);
nand U978 (N_978,In_454,In_1822);
nand U979 (N_979,In_648,In_2920);
or U980 (N_980,In_1618,In_2312);
xor U981 (N_981,In_106,In_532);
nor U982 (N_982,In_806,In_379);
nor U983 (N_983,In_2508,In_2669);
or U984 (N_984,In_1070,In_810);
or U985 (N_985,In_2362,In_2358);
nor U986 (N_986,In_2622,In_609);
and U987 (N_987,In_270,In_673);
xor U988 (N_988,In_374,In_1015);
and U989 (N_989,In_912,In_1785);
nand U990 (N_990,In_2830,In_2434);
xor U991 (N_991,In_502,In_2850);
nor U992 (N_992,In_1293,In_2690);
nand U993 (N_993,In_627,In_1921);
and U994 (N_994,In_139,In_1021);
or U995 (N_995,In_744,In_2163);
nor U996 (N_996,In_119,In_1433);
xnor U997 (N_997,In_2193,In_793);
and U998 (N_998,In_300,In_1534);
xnor U999 (N_999,In_1901,In_687);
nor U1000 (N_1000,In_2687,In_2558);
nor U1001 (N_1001,In_1651,In_1173);
and U1002 (N_1002,In_1813,In_1541);
nand U1003 (N_1003,In_1352,In_1198);
and U1004 (N_1004,In_1645,In_1918);
and U1005 (N_1005,In_2145,In_32);
or U1006 (N_1006,In_1556,In_1722);
nand U1007 (N_1007,In_1995,In_1937);
nand U1008 (N_1008,In_959,In_2552);
nor U1009 (N_1009,In_763,In_1191);
or U1010 (N_1010,In_2809,In_2770);
or U1011 (N_1011,In_638,In_2414);
nor U1012 (N_1012,In_2908,In_207);
nor U1013 (N_1013,In_566,In_2394);
or U1014 (N_1014,In_2678,In_961);
nor U1015 (N_1015,In_406,In_1545);
or U1016 (N_1016,In_214,In_2428);
nand U1017 (N_1017,In_1075,In_2825);
and U1018 (N_1018,In_2931,In_2639);
and U1019 (N_1019,In_1941,In_1043);
nand U1020 (N_1020,In_1026,In_2296);
nor U1021 (N_1021,In_1231,In_30);
and U1022 (N_1022,In_351,In_1192);
nand U1023 (N_1023,In_51,In_2181);
nor U1024 (N_1024,In_89,In_2409);
nand U1025 (N_1025,In_511,In_344);
or U1026 (N_1026,In_2452,In_1337);
nand U1027 (N_1027,In_281,In_2099);
and U1028 (N_1028,In_500,In_1160);
nor U1029 (N_1029,In_2058,In_2310);
xnor U1030 (N_1030,In_2954,In_152);
xnor U1031 (N_1031,In_389,In_2129);
nand U1032 (N_1032,In_2754,In_1253);
xor U1033 (N_1033,In_1869,In_560);
and U1034 (N_1034,In_2102,In_116);
and U1035 (N_1035,In_2827,In_538);
nor U1036 (N_1036,In_697,In_321);
nand U1037 (N_1037,In_650,In_1515);
and U1038 (N_1038,In_1119,In_2120);
or U1039 (N_1039,In_1270,In_1032);
and U1040 (N_1040,In_2023,In_55);
nand U1041 (N_1041,In_1713,In_546);
nand U1042 (N_1042,In_2826,In_1935);
or U1043 (N_1043,In_14,In_1902);
nand U1044 (N_1044,In_2779,In_746);
xor U1045 (N_1045,In_712,In_1696);
xor U1046 (N_1046,In_373,In_2906);
nor U1047 (N_1047,In_1446,In_1983);
and U1048 (N_1048,In_941,In_2620);
xor U1049 (N_1049,In_2464,In_2645);
and U1050 (N_1050,In_1113,In_2536);
nand U1051 (N_1051,In_951,In_2914);
xor U1052 (N_1052,In_305,In_16);
xor U1053 (N_1053,In_2917,In_734);
xor U1054 (N_1054,In_2727,In_919);
or U1055 (N_1055,In_1658,In_608);
nor U1056 (N_1056,In_1944,In_1499);
nor U1057 (N_1057,In_2652,In_1564);
nor U1058 (N_1058,In_1452,In_248);
nand U1059 (N_1059,In_573,In_2126);
nand U1060 (N_1060,In_2925,In_2559);
or U1061 (N_1061,In_1840,In_671);
nand U1062 (N_1062,In_1502,In_1250);
xor U1063 (N_1063,In_2674,In_2945);
xor U1064 (N_1064,In_2298,In_1125);
or U1065 (N_1065,In_2423,In_85);
nand U1066 (N_1066,In_425,In_967);
and U1067 (N_1067,In_1468,In_730);
xnor U1068 (N_1068,In_1661,In_2124);
nand U1069 (N_1069,In_1332,In_2146);
xnor U1070 (N_1070,In_2644,In_2971);
or U1071 (N_1071,In_2991,In_1897);
or U1072 (N_1072,In_2548,In_1769);
xor U1073 (N_1073,In_1780,In_2881);
nor U1074 (N_1074,In_593,In_1724);
or U1075 (N_1075,In_1670,In_840);
nor U1076 (N_1076,In_2729,In_123);
nor U1077 (N_1077,In_1649,In_224);
nor U1078 (N_1078,In_1234,In_1416);
or U1079 (N_1079,In_1226,In_317);
nor U1080 (N_1080,In_684,In_2828);
and U1081 (N_1081,In_471,In_62);
nor U1082 (N_1082,In_2705,In_799);
xnor U1083 (N_1083,In_2998,In_631);
and U1084 (N_1084,In_2725,In_2206);
or U1085 (N_1085,In_1657,In_2293);
or U1086 (N_1086,In_2820,In_189);
nand U1087 (N_1087,In_506,In_148);
and U1088 (N_1088,In_278,In_2343);
and U1089 (N_1089,In_601,In_2021);
nor U1090 (N_1090,In_1638,In_194);
nand U1091 (N_1091,In_2528,In_1345);
or U1092 (N_1092,In_814,In_2134);
or U1093 (N_1093,In_1569,In_2059);
nand U1094 (N_1094,In_1497,In_67);
or U1095 (N_1095,In_1691,In_1297);
and U1096 (N_1096,In_984,In_1411);
or U1097 (N_1097,In_1424,In_1006);
nor U1098 (N_1098,In_1612,In_2262);
or U1099 (N_1099,In_2890,In_877);
nand U1100 (N_1100,In_1038,In_459);
nor U1101 (N_1101,In_421,In_2223);
xor U1102 (N_1102,In_432,In_2762);
and U1103 (N_1103,In_2984,In_1472);
and U1104 (N_1104,In_865,In_1831);
xnor U1105 (N_1105,In_54,In_100);
and U1106 (N_1106,In_757,In_854);
nand U1107 (N_1107,In_1221,In_847);
nor U1108 (N_1108,In_2378,In_1623);
or U1109 (N_1109,In_1746,In_1907);
and U1110 (N_1110,In_659,In_95);
or U1111 (N_1111,In_752,In_467);
nand U1112 (N_1112,In_2327,In_2899);
or U1113 (N_1113,In_2968,In_2411);
nor U1114 (N_1114,In_2477,In_2340);
and U1115 (N_1115,In_1528,In_1399);
nor U1116 (N_1116,In_92,In_1762);
or U1117 (N_1117,In_2404,In_2750);
xor U1118 (N_1118,In_2556,In_372);
xor U1119 (N_1119,In_1851,In_440);
or U1120 (N_1120,In_953,In_1672);
nor U1121 (N_1121,In_2960,In_1093);
xor U1122 (N_1122,In_1039,In_564);
nand U1123 (N_1123,In_1150,In_1420);
nand U1124 (N_1124,In_127,In_2491);
xor U1125 (N_1125,In_1135,In_7);
xnor U1126 (N_1126,In_1570,In_2370);
nor U1127 (N_1127,In_2703,In_2865);
xor U1128 (N_1128,In_2365,In_2582);
and U1129 (N_1129,In_1543,In_834);
nand U1130 (N_1130,In_1938,In_737);
xor U1131 (N_1131,In_842,In_2267);
nor U1132 (N_1132,In_1593,In_2745);
nor U1133 (N_1133,In_1916,In_19);
or U1134 (N_1134,In_891,In_501);
nor U1135 (N_1135,In_1856,In_1804);
nor U1136 (N_1136,In_1818,In_1219);
or U1137 (N_1137,In_141,In_478);
or U1138 (N_1138,In_625,In_1007);
nor U1139 (N_1139,In_2905,In_1540);
or U1140 (N_1140,In_336,In_1417);
xor U1141 (N_1141,In_1735,In_444);
nor U1142 (N_1142,In_1201,In_2127);
xnor U1143 (N_1143,In_1917,In_876);
or U1144 (N_1144,In_1739,In_198);
and U1145 (N_1145,In_131,In_1290);
xnor U1146 (N_1146,In_987,In_2323);
nor U1147 (N_1147,In_2965,In_1422);
nand U1148 (N_1148,In_2105,In_544);
nor U1149 (N_1149,In_1884,In_2944);
nand U1150 (N_1150,In_2707,In_63);
xor U1151 (N_1151,In_258,In_297);
or U1152 (N_1152,In_2969,In_1390);
and U1153 (N_1153,In_2670,In_2072);
or U1154 (N_1154,In_404,In_345);
xor U1155 (N_1155,In_924,In_2113);
nand U1156 (N_1156,In_72,In_175);
nor U1157 (N_1157,In_822,In_2790);
xor U1158 (N_1158,In_271,In_2269);
or U1159 (N_1159,In_2009,In_1508);
and U1160 (N_1160,In_1513,In_1677);
xnor U1161 (N_1161,In_1169,In_2489);
nor U1162 (N_1162,In_1558,In_2149);
and U1163 (N_1163,In_199,In_801);
nand U1164 (N_1164,In_786,In_31);
nor U1165 (N_1165,In_2834,In_1924);
nand U1166 (N_1166,In_2572,In_921);
xor U1167 (N_1167,In_1153,In_1910);
nor U1168 (N_1168,In_1862,In_1045);
nand U1169 (N_1169,In_1674,In_783);
nor U1170 (N_1170,In_1858,In_1394);
or U1171 (N_1171,In_246,In_2025);
nand U1172 (N_1172,In_181,In_1946);
and U1173 (N_1173,In_2526,In_1494);
xnor U1174 (N_1174,In_2317,In_2546);
nand U1175 (N_1175,In_2700,In_1519);
nand U1176 (N_1176,In_2150,In_988);
nor U1177 (N_1177,In_1425,In_1005);
nand U1178 (N_1178,In_2757,In_304);
xor U1179 (N_1179,In_896,In_2609);
xnor U1180 (N_1180,In_887,In_1120);
xor U1181 (N_1181,In_1310,In_129);
and U1182 (N_1182,In_1078,In_2454);
nand U1183 (N_1183,In_1351,In_1243);
nand U1184 (N_1184,In_334,In_431);
or U1185 (N_1185,In_1529,In_2478);
and U1186 (N_1186,In_764,In_2152);
xor U1187 (N_1187,In_1299,In_185);
xor U1188 (N_1188,In_1707,In_1136);
xnor U1189 (N_1189,In_1204,In_2140);
or U1190 (N_1190,In_583,In_1336);
and U1191 (N_1191,In_531,In_2162);
and U1192 (N_1192,In_2051,In_2793);
nand U1193 (N_1193,In_316,In_701);
xor U1194 (N_1194,In_612,In_998);
xnor U1195 (N_1195,In_735,In_1463);
nand U1196 (N_1196,In_818,In_2040);
nand U1197 (N_1197,In_862,In_1830);
nand U1198 (N_1198,In_1815,In_1727);
and U1199 (N_1199,In_17,In_741);
or U1200 (N_1200,In_2997,In_1571);
nor U1201 (N_1201,In_1675,In_1041);
or U1202 (N_1202,In_1034,In_1098);
nor U1203 (N_1203,In_113,In_2360);
and U1204 (N_1204,In_2712,In_952);
or U1205 (N_1205,In_1281,In_534);
xnor U1206 (N_1206,In_750,In_879);
and U1207 (N_1207,In_2060,In_2078);
nor U1208 (N_1208,In_34,In_2109);
or U1209 (N_1209,In_2227,In_1020);
and U1210 (N_1210,In_1646,In_1445);
xnor U1211 (N_1211,In_821,In_2643);
xor U1212 (N_1212,In_2748,In_720);
and U1213 (N_1213,In_1827,In_2682);
xnor U1214 (N_1214,In_136,In_167);
nor U1215 (N_1215,In_2803,In_1969);
and U1216 (N_1216,In_285,In_755);
and U1217 (N_1217,In_2667,In_1025);
nand U1218 (N_1218,In_853,In_1750);
or U1219 (N_1219,In_2903,In_2255);
nor U1220 (N_1220,In_1304,In_433);
nand U1221 (N_1221,In_883,In_1899);
nor U1222 (N_1222,In_2057,In_504);
and U1223 (N_1223,In_1733,In_470);
and U1224 (N_1224,In_315,In_1121);
xor U1225 (N_1225,In_1772,In_510);
or U1226 (N_1226,In_1710,In_1557);
or U1227 (N_1227,In_1755,In_1887);
nor U1228 (N_1228,In_2161,In_2927);
or U1229 (N_1229,In_2074,In_582);
or U1230 (N_1230,In_1227,In_3);
or U1231 (N_1231,In_188,In_965);
and U1232 (N_1232,In_836,In_1922);
nor U1233 (N_1233,In_2871,In_1637);
or U1234 (N_1234,In_128,In_600);
and U1235 (N_1235,In_1249,In_711);
nor U1236 (N_1236,In_235,In_1195);
nand U1237 (N_1237,In_98,In_2799);
or U1238 (N_1238,In_392,In_860);
or U1239 (N_1239,In_2668,In_828);
or U1240 (N_1240,In_1448,In_435);
and U1241 (N_1241,In_948,In_760);
nand U1242 (N_1242,In_1368,In_1464);
xor U1243 (N_1243,In_1441,In_1140);
nor U1244 (N_1244,In_1365,In_695);
and U1245 (N_1245,In_45,In_2742);
xor U1246 (N_1246,In_2759,In_575);
or U1247 (N_1247,In_2439,In_283);
nand U1248 (N_1248,In_2498,In_1382);
nand U1249 (N_1249,In_636,In_2517);
nand U1250 (N_1250,In_1774,In_1205);
or U1251 (N_1251,In_2053,In_1442);
xor U1252 (N_1252,In_1592,In_922);
or U1253 (N_1253,In_475,In_2618);
xor U1254 (N_1254,In_1322,In_122);
xor U1255 (N_1255,In_856,In_1518);
or U1256 (N_1256,In_1989,In_800);
xnor U1257 (N_1257,In_2341,In_796);
nand U1258 (N_1258,In_2540,In_2574);
nor U1259 (N_1259,In_722,In_2400);
xor U1260 (N_1260,In_2114,In_2367);
or U1261 (N_1261,In_2383,In_1102);
nand U1262 (N_1262,In_604,In_436);
xor U1263 (N_1263,In_2989,In_2242);
nor U1264 (N_1264,In_2868,In_252);
or U1265 (N_1265,In_86,In_1949);
and U1266 (N_1266,In_367,In_762);
and U1267 (N_1267,In_1685,In_117);
nand U1268 (N_1268,In_154,In_542);
xor U1269 (N_1269,In_254,In_1371);
and U1270 (N_1270,In_709,In_1550);
and U1271 (N_1271,In_2934,In_1932);
nand U1272 (N_1272,In_1406,In_1317);
and U1273 (N_1273,In_2979,In_1358);
xor U1274 (N_1274,In_1470,In_619);
nor U1275 (N_1275,In_2015,In_1925);
or U1276 (N_1276,In_704,In_343);
xnor U1277 (N_1277,In_427,In_327);
nand U1278 (N_1278,In_2842,In_1743);
nand U1279 (N_1279,In_1182,In_994);
or U1280 (N_1280,In_1100,In_1629);
nor U1281 (N_1281,In_1860,In_1600);
or U1282 (N_1282,In_91,In_1611);
or U1283 (N_1283,In_1982,In_1301);
nand U1284 (N_1284,In_1749,In_424);
nand U1285 (N_1285,In_1585,In_2594);
xor U1286 (N_1286,In_2584,In_868);
xor U1287 (N_1287,In_2253,In_208);
or U1288 (N_1288,In_535,In_1844);
nor U1289 (N_1289,In_2332,In_1375);
and U1290 (N_1290,In_236,In_174);
nand U1291 (N_1291,In_1259,In_759);
nand U1292 (N_1292,In_2693,In_1697);
or U1293 (N_1293,In_2549,In_1711);
and U1294 (N_1294,In_245,In_1561);
nor U1295 (N_1295,In_1584,In_954);
xnor U1296 (N_1296,In_1781,In_1904);
and U1297 (N_1297,In_1133,In_322);
or U1298 (N_1298,In_2642,In_537);
nor U1299 (N_1299,In_1237,In_2872);
nor U1300 (N_1300,In_748,In_2379);
or U1301 (N_1301,In_2226,In_1401);
and U1302 (N_1302,In_2412,In_371);
nor U1303 (N_1303,In_2251,In_288);
nand U1304 (N_1304,In_920,In_2932);
and U1305 (N_1305,In_2112,In_553);
nor U1306 (N_1306,In_2735,In_517);
and U1307 (N_1307,In_333,In_1927);
nand U1308 (N_1308,In_1359,In_1068);
xor U1309 (N_1309,In_930,In_851);
and U1310 (N_1310,In_2500,In_2502);
nor U1311 (N_1311,In_1882,In_1760);
nand U1312 (N_1312,In_838,In_2244);
xnor U1313 (N_1313,In_1797,In_2007);
or U1314 (N_1314,In_180,In_1467);
nor U1315 (N_1315,In_817,In_507);
xor U1316 (N_1316,In_293,In_2207);
nor U1317 (N_1317,In_580,In_1853);
or U1318 (N_1318,In_2487,In_428);
xor U1319 (N_1319,In_1523,In_571);
nand U1320 (N_1320,In_2018,In_1752);
xor U1321 (N_1321,In_2320,In_2274);
nand U1322 (N_1322,In_823,In_706);
and U1323 (N_1323,In_1320,In_2453);
and U1324 (N_1324,In_135,In_1756);
xnor U1325 (N_1325,In_2974,In_1271);
nand U1326 (N_1326,In_409,In_864);
xnor U1327 (N_1327,In_1586,In_1489);
nand U1328 (N_1328,In_2659,In_1650);
xor U1329 (N_1329,In_992,In_1284);
or U1330 (N_1330,In_2006,In_2638);
xnor U1331 (N_1331,In_260,In_2043);
or U1332 (N_1332,In_633,In_2289);
xor U1333 (N_1333,In_1294,In_487);
or U1334 (N_1334,In_1427,In_1168);
xor U1335 (N_1335,In_1235,In_15);
xnor U1336 (N_1336,In_1655,In_1652);
xnor U1337 (N_1337,In_1190,In_2375);
xor U1338 (N_1338,In_2988,In_484);
or U1339 (N_1339,In_1633,In_1247);
or U1340 (N_1340,In_279,In_1861);
nand U1341 (N_1341,In_446,In_229);
or U1342 (N_1342,In_1081,In_1737);
or U1343 (N_1343,In_2048,In_1289);
xor U1344 (N_1344,In_1388,In_1312);
nor U1345 (N_1345,In_1764,In_2130);
nor U1346 (N_1346,In_576,In_1124);
or U1347 (N_1347,In_1240,In_118);
xnor U1348 (N_1348,In_2675,In_146);
xor U1349 (N_1349,In_1138,In_2287);
or U1350 (N_1350,In_1344,In_2171);
nor U1351 (N_1351,In_2345,In_222);
and U1352 (N_1352,In_903,In_2138);
and U1353 (N_1353,In_1220,In_2325);
or U1354 (N_1354,In_2108,In_2818);
nor U1355 (N_1355,In_2087,In_423);
xnor U1356 (N_1356,In_916,In_1040);
or U1357 (N_1357,In_1978,In_1751);
nor U1358 (N_1358,In_495,In_410);
and U1359 (N_1359,In_2956,In_1272);
and U1360 (N_1360,In_2170,In_2981);
nand U1361 (N_1361,In_1972,In_2952);
nor U1362 (N_1362,In_71,In_2857);
or U1363 (N_1363,In_2467,In_1548);
xnor U1364 (N_1364,In_688,In_132);
nand U1365 (N_1365,In_498,In_1454);
nand U1366 (N_1366,In_219,In_1307);
nand U1367 (N_1367,In_626,In_2571);
nand U1368 (N_1368,In_1888,In_2547);
xor U1369 (N_1369,In_768,In_2122);
nor U1370 (N_1370,In_2887,In_1647);
or U1371 (N_1371,In_1123,In_1436);
and U1372 (N_1372,In_2889,In_2012);
xor U1373 (N_1373,In_2459,In_1429);
nand U1374 (N_1374,In_1622,In_543);
nand U1375 (N_1375,In_2529,In_1355);
or U1376 (N_1376,In_1717,In_6);
nor U1377 (N_1377,In_524,In_2313);
and U1378 (N_1378,In_1476,In_1664);
and U1379 (N_1379,In_2117,In_556);
nand U1380 (N_1380,In_184,In_925);
nor U1381 (N_1381,In_109,In_1948);
nor U1382 (N_1382,In_418,In_1909);
and U1383 (N_1383,In_2628,In_1731);
xor U1384 (N_1384,In_944,In_1061);
xnor U1385 (N_1385,In_2103,In_1988);
nor U1386 (N_1386,In_2525,In_956);
nand U1387 (N_1387,In_751,In_2901);
and U1388 (N_1388,In_2641,In_2940);
or U1389 (N_1389,In_2698,In_1363);
and U1390 (N_1390,In_158,In_490);
nor U1391 (N_1391,In_1782,In_211);
xor U1392 (N_1392,In_422,In_2853);
and U1393 (N_1393,In_2449,In_2590);
nor U1394 (N_1394,In_2570,In_780);
nor U1395 (N_1395,In_562,In_273);
nor U1396 (N_1396,In_1372,In_204);
or U1397 (N_1397,In_886,In_1606);
nor U1398 (N_1398,In_401,In_1621);
xnor U1399 (N_1399,In_1286,In_1218);
or U1400 (N_1400,In_339,In_2201);
or U1401 (N_1401,In_1990,In_1232);
or U1402 (N_1402,In_2022,In_2624);
nand U1403 (N_1403,In_2191,In_1511);
or U1404 (N_1404,In_1977,In_23);
nor U1405 (N_1405,In_197,In_1161);
and U1406 (N_1406,In_2073,In_209);
nor U1407 (N_1407,In_1555,In_2787);
nand U1408 (N_1408,In_492,In_1575);
and U1409 (N_1409,In_1705,In_169);
and U1410 (N_1410,In_2410,In_1263);
nand U1411 (N_1411,In_377,In_819);
and U1412 (N_1412,In_2460,In_2596);
nor U1413 (N_1413,In_923,In_499);
and U1414 (N_1414,In_88,In_970);
or U1415 (N_1415,In_310,In_1708);
or U1416 (N_1416,In_2352,In_1378);
xnor U1417 (N_1417,In_2239,In_1398);
xnor U1418 (N_1418,In_1676,In_1176);
nand U1419 (N_1419,In_2424,In_2180);
nor U1420 (N_1420,In_2131,In_2258);
or U1421 (N_1421,In_1803,In_2519);
nor U1422 (N_1422,In_2902,In_2208);
xnor U1423 (N_1423,In_1963,In_2699);
nor U1424 (N_1424,In_458,In_1975);
and U1425 (N_1425,In_666,In_2895);
and U1426 (N_1426,In_1019,In_74);
nor U1427 (N_1427,In_646,In_218);
and U1428 (N_1428,In_1260,In_782);
or U1429 (N_1429,In_240,In_2290);
nor U1430 (N_1430,In_1786,In_1014);
or U1431 (N_1431,In_979,In_1500);
nor U1432 (N_1432,In_1599,In_1309);
nand U1433 (N_1433,In_2420,In_2648);
or U1434 (N_1434,In_1001,In_1855);
nor U1435 (N_1435,In_302,In_2366);
nor U1436 (N_1436,In_578,In_415);
nor U1437 (N_1437,In_1361,In_927);
xnor U1438 (N_1438,In_585,In_2861);
xnor U1439 (N_1439,In_2788,In_2071);
nor U1440 (N_1440,In_2875,In_1418);
nor U1441 (N_1441,In_453,In_1114);
xor U1442 (N_1442,In_1587,In_1152);
or U1443 (N_1443,In_771,In_1667);
and U1444 (N_1444,In_399,In_645);
nor U1445 (N_1445,In_906,In_1939);
xor U1446 (N_1446,In_950,In_1913);
and U1447 (N_1447,In_1879,In_35);
nand U1448 (N_1448,In_1506,In_1315);
or U1449 (N_1449,In_2398,In_1386);
nor U1450 (N_1450,In_2630,In_855);
xor U1451 (N_1451,In_2442,In_2215);
nand U1452 (N_1452,In_2211,In_1066);
and U1453 (N_1453,In_2210,In_846);
nor U1454 (N_1454,In_2553,In_1779);
nand U1455 (N_1455,In_509,In_943);
nand U1456 (N_1456,In_1729,In_668);
xnor U1457 (N_1457,In_2603,In_2737);
and U1458 (N_1458,In_997,In_1274);
or U1459 (N_1459,In_1947,In_2003);
and U1460 (N_1460,In_2812,In_1620);
and U1461 (N_1461,In_1179,In_1159);
or U1462 (N_1462,In_450,In_1838);
and U1463 (N_1463,In_2538,In_445);
and U1464 (N_1464,In_1404,In_330);
and U1465 (N_1465,In_2292,In_1279);
nor U1466 (N_1466,In_803,In_2543);
nor U1467 (N_1467,In_114,In_378);
xor U1468 (N_1468,In_138,In_1706);
or U1469 (N_1469,In_2555,In_1008);
nor U1470 (N_1470,In_1656,In_1859);
nor U1471 (N_1471,In_1820,In_1619);
or U1472 (N_1472,In_2066,In_2214);
or U1473 (N_1473,In_2611,In_361);
xor U1474 (N_1474,In_1716,In_396);
xnor U1475 (N_1475,In_1462,In_2761);
and U1476 (N_1476,In_1431,In_2599);
or U1477 (N_1477,In_2567,In_1033);
or U1478 (N_1478,In_770,In_12);
and U1479 (N_1479,In_1419,In_1266);
nand U1480 (N_1480,In_857,In_2840);
xor U1481 (N_1481,In_1720,In_359);
and U1482 (N_1482,In_2104,In_663);
nor U1483 (N_1483,In_1096,In_597);
or U1484 (N_1484,In_2530,In_1563);
or U1485 (N_1485,In_2604,In_112);
xnor U1486 (N_1486,In_1929,In_81);
or U1487 (N_1487,In_1771,In_2702);
xnor U1488 (N_1488,In_1766,In_93);
xor U1489 (N_1489,In_550,In_1111);
or U1490 (N_1490,In_2535,In_2441);
nor U1491 (N_1491,In_530,In_105);
and U1492 (N_1492,In_588,In_2869);
and U1493 (N_1493,In_1572,In_1784);
xnor U1494 (N_1494,In_1151,In_2755);
nor U1495 (N_1495,In_2653,In_2318);
and U1496 (N_1496,In_995,In_195);
or U1497 (N_1497,In_2859,In_1991);
and U1498 (N_1498,In_1866,In_2990);
nand U1499 (N_1499,In_2892,In_2272);
or U1500 (N_1500,In_667,In_2512);
nor U1501 (N_1501,In_592,In_1303);
and U1502 (N_1502,In_1740,In_1454);
nor U1503 (N_1503,In_2667,In_671);
xor U1504 (N_1504,In_2468,In_245);
and U1505 (N_1505,In_2472,In_1505);
nand U1506 (N_1506,In_1304,In_2787);
xnor U1507 (N_1507,In_1764,In_575);
xor U1508 (N_1508,In_739,In_2354);
xor U1509 (N_1509,In_60,In_316);
nand U1510 (N_1510,In_953,In_548);
nor U1511 (N_1511,In_1355,In_2730);
xnor U1512 (N_1512,In_172,In_878);
nand U1513 (N_1513,In_2482,In_1733);
and U1514 (N_1514,In_1657,In_118);
xor U1515 (N_1515,In_2064,In_1);
nor U1516 (N_1516,In_1646,In_473);
nor U1517 (N_1517,In_357,In_1283);
xor U1518 (N_1518,In_432,In_1512);
nor U1519 (N_1519,In_2925,In_1135);
nor U1520 (N_1520,In_2687,In_1947);
xor U1521 (N_1521,In_498,In_1249);
xor U1522 (N_1522,In_860,In_386);
nand U1523 (N_1523,In_1297,In_2268);
and U1524 (N_1524,In_2921,In_2110);
nand U1525 (N_1525,In_10,In_2772);
and U1526 (N_1526,In_323,In_37);
or U1527 (N_1527,In_1985,In_1001);
and U1528 (N_1528,In_2983,In_454);
nor U1529 (N_1529,In_164,In_1651);
nor U1530 (N_1530,In_2779,In_2941);
or U1531 (N_1531,In_892,In_264);
and U1532 (N_1532,In_2567,In_1607);
or U1533 (N_1533,In_1265,In_679);
and U1534 (N_1534,In_485,In_2569);
xnor U1535 (N_1535,In_1901,In_2994);
nor U1536 (N_1536,In_1553,In_263);
nor U1537 (N_1537,In_363,In_1677);
and U1538 (N_1538,In_30,In_1467);
nand U1539 (N_1539,In_2687,In_452);
nand U1540 (N_1540,In_1616,In_1460);
and U1541 (N_1541,In_1430,In_1983);
and U1542 (N_1542,In_690,In_2623);
nand U1543 (N_1543,In_1923,In_1730);
or U1544 (N_1544,In_2312,In_2140);
nand U1545 (N_1545,In_2163,In_1777);
nor U1546 (N_1546,In_438,In_1113);
or U1547 (N_1547,In_1384,In_2369);
nand U1548 (N_1548,In_943,In_2021);
nand U1549 (N_1549,In_1771,In_609);
xnor U1550 (N_1550,In_1097,In_31);
xnor U1551 (N_1551,In_1614,In_2455);
nor U1552 (N_1552,In_804,In_279);
nor U1553 (N_1553,In_43,In_354);
or U1554 (N_1554,In_2471,In_1470);
xnor U1555 (N_1555,In_908,In_1416);
nor U1556 (N_1556,In_2871,In_488);
or U1557 (N_1557,In_2708,In_70);
and U1558 (N_1558,In_2785,In_1293);
and U1559 (N_1559,In_262,In_1732);
or U1560 (N_1560,In_1547,In_1346);
and U1561 (N_1561,In_2242,In_677);
and U1562 (N_1562,In_142,In_855);
nand U1563 (N_1563,In_995,In_552);
nor U1564 (N_1564,In_2423,In_2007);
and U1565 (N_1565,In_23,In_907);
xor U1566 (N_1566,In_1590,In_2927);
and U1567 (N_1567,In_1285,In_1361);
or U1568 (N_1568,In_993,In_1690);
nor U1569 (N_1569,In_1748,In_262);
and U1570 (N_1570,In_1638,In_924);
nand U1571 (N_1571,In_1224,In_2889);
xor U1572 (N_1572,In_1498,In_1745);
nand U1573 (N_1573,In_2547,In_2662);
and U1574 (N_1574,In_976,In_1198);
xnor U1575 (N_1575,In_2331,In_245);
and U1576 (N_1576,In_1207,In_2386);
and U1577 (N_1577,In_1760,In_2310);
and U1578 (N_1578,In_2751,In_1941);
or U1579 (N_1579,In_416,In_345);
xor U1580 (N_1580,In_436,In_2599);
and U1581 (N_1581,In_2520,In_1098);
or U1582 (N_1582,In_2685,In_1768);
and U1583 (N_1583,In_352,In_1571);
nor U1584 (N_1584,In_2537,In_850);
nor U1585 (N_1585,In_45,In_1393);
or U1586 (N_1586,In_187,In_2466);
nand U1587 (N_1587,In_2422,In_584);
nor U1588 (N_1588,In_308,In_1251);
xor U1589 (N_1589,In_2894,In_175);
and U1590 (N_1590,In_1236,In_1543);
nor U1591 (N_1591,In_2466,In_2962);
or U1592 (N_1592,In_300,In_2372);
or U1593 (N_1593,In_778,In_1752);
and U1594 (N_1594,In_289,In_492);
xor U1595 (N_1595,In_119,In_2811);
nor U1596 (N_1596,In_50,In_2820);
nand U1597 (N_1597,In_954,In_2180);
xor U1598 (N_1598,In_2849,In_1159);
nor U1599 (N_1599,In_1397,In_2482);
xnor U1600 (N_1600,In_1412,In_662);
and U1601 (N_1601,In_770,In_2649);
or U1602 (N_1602,In_1520,In_454);
or U1603 (N_1603,In_437,In_2709);
and U1604 (N_1604,In_2826,In_1047);
nor U1605 (N_1605,In_2312,In_587);
or U1606 (N_1606,In_381,In_2393);
xor U1607 (N_1607,In_1731,In_110);
nand U1608 (N_1608,In_1703,In_780);
nand U1609 (N_1609,In_790,In_2148);
or U1610 (N_1610,In_2278,In_668);
or U1611 (N_1611,In_2787,In_696);
xor U1612 (N_1612,In_2451,In_1895);
xor U1613 (N_1613,In_1914,In_2052);
or U1614 (N_1614,In_1970,In_2011);
nor U1615 (N_1615,In_2614,In_2730);
xor U1616 (N_1616,In_2626,In_500);
nand U1617 (N_1617,In_2546,In_211);
and U1618 (N_1618,In_2037,In_1635);
or U1619 (N_1619,In_827,In_873);
or U1620 (N_1620,In_1343,In_2608);
and U1621 (N_1621,In_2953,In_863);
nor U1622 (N_1622,In_1458,In_595);
nand U1623 (N_1623,In_2792,In_2027);
or U1624 (N_1624,In_904,In_497);
nor U1625 (N_1625,In_1397,In_1744);
or U1626 (N_1626,In_126,In_304);
and U1627 (N_1627,In_11,In_1037);
nand U1628 (N_1628,In_2730,In_508);
or U1629 (N_1629,In_1435,In_1178);
nor U1630 (N_1630,In_469,In_695);
or U1631 (N_1631,In_1282,In_81);
or U1632 (N_1632,In_2060,In_255);
nand U1633 (N_1633,In_1814,In_2507);
and U1634 (N_1634,In_1103,In_1205);
xnor U1635 (N_1635,In_1454,In_439);
or U1636 (N_1636,In_115,In_1568);
and U1637 (N_1637,In_664,In_1355);
xor U1638 (N_1638,In_631,In_2089);
and U1639 (N_1639,In_294,In_2840);
nor U1640 (N_1640,In_1368,In_1858);
and U1641 (N_1641,In_885,In_2591);
or U1642 (N_1642,In_656,In_996);
and U1643 (N_1643,In_2038,In_1381);
and U1644 (N_1644,In_420,In_2850);
nor U1645 (N_1645,In_2456,In_2487);
xnor U1646 (N_1646,In_848,In_1133);
nor U1647 (N_1647,In_1306,In_832);
nor U1648 (N_1648,In_92,In_821);
and U1649 (N_1649,In_602,In_146);
and U1650 (N_1650,In_1827,In_998);
nor U1651 (N_1651,In_1107,In_1497);
and U1652 (N_1652,In_2852,In_2357);
and U1653 (N_1653,In_1682,In_1005);
or U1654 (N_1654,In_1424,In_2597);
or U1655 (N_1655,In_378,In_2241);
xnor U1656 (N_1656,In_1861,In_239);
or U1657 (N_1657,In_501,In_2579);
nand U1658 (N_1658,In_1598,In_2515);
nand U1659 (N_1659,In_321,In_347);
or U1660 (N_1660,In_1989,In_2998);
nor U1661 (N_1661,In_2855,In_1889);
and U1662 (N_1662,In_989,In_88);
or U1663 (N_1663,In_1621,In_391);
nor U1664 (N_1664,In_2717,In_90);
and U1665 (N_1665,In_562,In_2012);
or U1666 (N_1666,In_1163,In_2817);
xor U1667 (N_1667,In_2280,In_2975);
nand U1668 (N_1668,In_977,In_2804);
nor U1669 (N_1669,In_2566,In_779);
or U1670 (N_1670,In_2185,In_215);
nor U1671 (N_1671,In_2950,In_1811);
xnor U1672 (N_1672,In_1122,In_2078);
xor U1673 (N_1673,In_1322,In_1796);
xor U1674 (N_1674,In_528,In_144);
and U1675 (N_1675,In_2401,In_1012);
nand U1676 (N_1676,In_464,In_2577);
or U1677 (N_1677,In_943,In_2341);
and U1678 (N_1678,In_1941,In_792);
or U1679 (N_1679,In_319,In_306);
nor U1680 (N_1680,In_1940,In_2178);
nor U1681 (N_1681,In_605,In_1291);
xor U1682 (N_1682,In_2696,In_2078);
nand U1683 (N_1683,In_888,In_1360);
xnor U1684 (N_1684,In_702,In_2250);
xor U1685 (N_1685,In_914,In_1321);
nand U1686 (N_1686,In_536,In_192);
nand U1687 (N_1687,In_715,In_204);
nand U1688 (N_1688,In_59,In_1047);
and U1689 (N_1689,In_2983,In_362);
nor U1690 (N_1690,In_1988,In_1722);
xor U1691 (N_1691,In_1537,In_98);
or U1692 (N_1692,In_2302,In_906);
nand U1693 (N_1693,In_1983,In_1982);
or U1694 (N_1694,In_1138,In_610);
xnor U1695 (N_1695,In_2516,In_43);
nand U1696 (N_1696,In_1744,In_788);
nand U1697 (N_1697,In_851,In_2000);
xnor U1698 (N_1698,In_1703,In_2982);
nand U1699 (N_1699,In_1498,In_1557);
and U1700 (N_1700,In_2115,In_392);
xor U1701 (N_1701,In_1814,In_377);
nor U1702 (N_1702,In_763,In_2747);
xnor U1703 (N_1703,In_474,In_1085);
and U1704 (N_1704,In_1017,In_1657);
nand U1705 (N_1705,In_959,In_516);
xor U1706 (N_1706,In_783,In_1331);
nor U1707 (N_1707,In_2470,In_2817);
and U1708 (N_1708,In_2164,In_1892);
or U1709 (N_1709,In_829,In_2299);
nor U1710 (N_1710,In_873,In_1171);
or U1711 (N_1711,In_502,In_737);
nor U1712 (N_1712,In_2945,In_22);
or U1713 (N_1713,In_1768,In_1636);
or U1714 (N_1714,In_2425,In_2914);
or U1715 (N_1715,In_440,In_1776);
or U1716 (N_1716,In_804,In_1465);
xnor U1717 (N_1717,In_1993,In_231);
or U1718 (N_1718,In_309,In_152);
and U1719 (N_1719,In_38,In_188);
xnor U1720 (N_1720,In_745,In_72);
and U1721 (N_1721,In_118,In_2441);
or U1722 (N_1722,In_2722,In_2452);
and U1723 (N_1723,In_2655,In_1900);
nand U1724 (N_1724,In_1654,In_2384);
xnor U1725 (N_1725,In_572,In_2423);
or U1726 (N_1726,In_356,In_2179);
or U1727 (N_1727,In_1389,In_1734);
nor U1728 (N_1728,In_1608,In_279);
nor U1729 (N_1729,In_1186,In_760);
nand U1730 (N_1730,In_2398,In_2224);
or U1731 (N_1731,In_1437,In_1729);
or U1732 (N_1732,In_1217,In_1771);
nand U1733 (N_1733,In_2597,In_2867);
xor U1734 (N_1734,In_729,In_2318);
and U1735 (N_1735,In_735,In_362);
and U1736 (N_1736,In_2210,In_1384);
or U1737 (N_1737,In_979,In_1789);
nand U1738 (N_1738,In_2590,In_2074);
nor U1739 (N_1739,In_412,In_1067);
nand U1740 (N_1740,In_2423,In_2909);
nand U1741 (N_1741,In_1555,In_1855);
nor U1742 (N_1742,In_1376,In_2896);
nor U1743 (N_1743,In_1482,In_605);
nor U1744 (N_1744,In_2125,In_1923);
nor U1745 (N_1745,In_1592,In_2363);
and U1746 (N_1746,In_2803,In_658);
xor U1747 (N_1747,In_193,In_879);
and U1748 (N_1748,In_2041,In_1301);
xor U1749 (N_1749,In_2253,In_2363);
nand U1750 (N_1750,In_2508,In_2213);
or U1751 (N_1751,In_1994,In_2224);
nor U1752 (N_1752,In_2651,In_2825);
or U1753 (N_1753,In_508,In_1431);
xnor U1754 (N_1754,In_2684,In_2541);
or U1755 (N_1755,In_1341,In_323);
nor U1756 (N_1756,In_669,In_1989);
xor U1757 (N_1757,In_2248,In_205);
xor U1758 (N_1758,In_618,In_1947);
and U1759 (N_1759,In_1889,In_297);
nand U1760 (N_1760,In_2274,In_1404);
or U1761 (N_1761,In_2333,In_2555);
nand U1762 (N_1762,In_1831,In_1222);
and U1763 (N_1763,In_1384,In_79);
or U1764 (N_1764,In_1137,In_997);
nand U1765 (N_1765,In_1781,In_2336);
nor U1766 (N_1766,In_791,In_2841);
nand U1767 (N_1767,In_2284,In_1065);
xnor U1768 (N_1768,In_593,In_362);
and U1769 (N_1769,In_1783,In_851);
nor U1770 (N_1770,In_1352,In_37);
and U1771 (N_1771,In_525,In_1130);
and U1772 (N_1772,In_131,In_1208);
nor U1773 (N_1773,In_806,In_2656);
and U1774 (N_1774,In_969,In_1412);
nor U1775 (N_1775,In_504,In_898);
xnor U1776 (N_1776,In_1288,In_1083);
or U1777 (N_1777,In_2726,In_2471);
xor U1778 (N_1778,In_2547,In_2326);
or U1779 (N_1779,In_85,In_83);
or U1780 (N_1780,In_2772,In_2950);
and U1781 (N_1781,In_806,In_6);
xnor U1782 (N_1782,In_2656,In_629);
nand U1783 (N_1783,In_90,In_1256);
nand U1784 (N_1784,In_138,In_294);
xnor U1785 (N_1785,In_750,In_316);
or U1786 (N_1786,In_1434,In_1671);
and U1787 (N_1787,In_1836,In_64);
or U1788 (N_1788,In_2269,In_406);
and U1789 (N_1789,In_2640,In_554);
nand U1790 (N_1790,In_2573,In_2692);
or U1791 (N_1791,In_1955,In_1537);
and U1792 (N_1792,In_594,In_595);
or U1793 (N_1793,In_1507,In_1624);
nand U1794 (N_1794,In_2480,In_1728);
or U1795 (N_1795,In_914,In_2689);
nor U1796 (N_1796,In_2844,In_1164);
xor U1797 (N_1797,In_346,In_2421);
xor U1798 (N_1798,In_1456,In_2213);
xnor U1799 (N_1799,In_1825,In_1858);
and U1800 (N_1800,In_2249,In_916);
or U1801 (N_1801,In_2964,In_2928);
xnor U1802 (N_1802,In_1398,In_546);
nand U1803 (N_1803,In_2849,In_2025);
xnor U1804 (N_1804,In_672,In_1301);
and U1805 (N_1805,In_846,In_2758);
or U1806 (N_1806,In_2076,In_340);
nor U1807 (N_1807,In_1544,In_2480);
nand U1808 (N_1808,In_1647,In_1655);
or U1809 (N_1809,In_315,In_2611);
nand U1810 (N_1810,In_2906,In_1739);
nor U1811 (N_1811,In_262,In_2707);
or U1812 (N_1812,In_58,In_754);
xor U1813 (N_1813,In_2302,In_320);
or U1814 (N_1814,In_2614,In_149);
xor U1815 (N_1815,In_641,In_1423);
nand U1816 (N_1816,In_1689,In_979);
and U1817 (N_1817,In_2111,In_1348);
or U1818 (N_1818,In_2136,In_2497);
xnor U1819 (N_1819,In_214,In_2027);
xnor U1820 (N_1820,In_2111,In_740);
or U1821 (N_1821,In_2795,In_2142);
or U1822 (N_1822,In_2158,In_1053);
xnor U1823 (N_1823,In_946,In_2802);
nand U1824 (N_1824,In_2687,In_2349);
xor U1825 (N_1825,In_1241,In_2531);
xnor U1826 (N_1826,In_2423,In_478);
nor U1827 (N_1827,In_1447,In_1317);
xnor U1828 (N_1828,In_2898,In_1558);
or U1829 (N_1829,In_2039,In_1098);
nand U1830 (N_1830,In_1418,In_2186);
nor U1831 (N_1831,In_2295,In_1616);
or U1832 (N_1832,In_860,In_1241);
and U1833 (N_1833,In_2541,In_2275);
nor U1834 (N_1834,In_577,In_2956);
nor U1835 (N_1835,In_460,In_842);
or U1836 (N_1836,In_2857,In_2443);
nand U1837 (N_1837,In_1018,In_1617);
or U1838 (N_1838,In_2166,In_226);
nor U1839 (N_1839,In_1268,In_2532);
nor U1840 (N_1840,In_1836,In_511);
nand U1841 (N_1841,In_566,In_181);
and U1842 (N_1842,In_2291,In_1829);
nor U1843 (N_1843,In_2779,In_1044);
or U1844 (N_1844,In_1814,In_2814);
or U1845 (N_1845,In_2752,In_1975);
xnor U1846 (N_1846,In_1467,In_1669);
xnor U1847 (N_1847,In_2073,In_2812);
or U1848 (N_1848,In_2816,In_1994);
or U1849 (N_1849,In_1423,In_449);
and U1850 (N_1850,In_1240,In_419);
and U1851 (N_1851,In_2012,In_1635);
nor U1852 (N_1852,In_2861,In_382);
and U1853 (N_1853,In_166,In_846);
and U1854 (N_1854,In_1800,In_434);
nor U1855 (N_1855,In_2901,In_1518);
and U1856 (N_1856,In_1384,In_1647);
nor U1857 (N_1857,In_1313,In_2706);
or U1858 (N_1858,In_1197,In_1895);
nor U1859 (N_1859,In_1669,In_746);
nand U1860 (N_1860,In_2352,In_1241);
and U1861 (N_1861,In_406,In_1471);
nor U1862 (N_1862,In_2806,In_271);
xor U1863 (N_1863,In_710,In_1914);
and U1864 (N_1864,In_492,In_722);
and U1865 (N_1865,In_2985,In_317);
or U1866 (N_1866,In_2808,In_2164);
nor U1867 (N_1867,In_1873,In_1909);
and U1868 (N_1868,In_1671,In_498);
and U1869 (N_1869,In_997,In_1536);
or U1870 (N_1870,In_2125,In_926);
nand U1871 (N_1871,In_812,In_1351);
nand U1872 (N_1872,In_1792,In_2452);
and U1873 (N_1873,In_2375,In_2880);
or U1874 (N_1874,In_971,In_358);
and U1875 (N_1875,In_666,In_1311);
or U1876 (N_1876,In_1572,In_2119);
or U1877 (N_1877,In_2297,In_654);
nand U1878 (N_1878,In_623,In_1388);
xor U1879 (N_1879,In_2858,In_1409);
or U1880 (N_1880,In_2555,In_2801);
or U1881 (N_1881,In_1845,In_14);
xnor U1882 (N_1882,In_865,In_2480);
and U1883 (N_1883,In_820,In_60);
and U1884 (N_1884,In_1819,In_958);
and U1885 (N_1885,In_2677,In_1820);
and U1886 (N_1886,In_1856,In_2081);
and U1887 (N_1887,In_2890,In_1541);
nand U1888 (N_1888,In_67,In_79);
or U1889 (N_1889,In_1039,In_2919);
and U1890 (N_1890,In_1337,In_1246);
and U1891 (N_1891,In_1867,In_1714);
nor U1892 (N_1892,In_2907,In_136);
nor U1893 (N_1893,In_352,In_2089);
xnor U1894 (N_1894,In_1962,In_403);
nand U1895 (N_1895,In_2662,In_1203);
xor U1896 (N_1896,In_1061,In_2510);
nor U1897 (N_1897,In_2909,In_1968);
xnor U1898 (N_1898,In_229,In_1222);
nand U1899 (N_1899,In_2858,In_2234);
xnor U1900 (N_1900,In_2981,In_2153);
nor U1901 (N_1901,In_1170,In_2361);
and U1902 (N_1902,In_1659,In_783);
or U1903 (N_1903,In_874,In_189);
nand U1904 (N_1904,In_2834,In_1085);
nor U1905 (N_1905,In_1312,In_2974);
nand U1906 (N_1906,In_586,In_1972);
or U1907 (N_1907,In_1904,In_113);
nand U1908 (N_1908,In_1344,In_342);
xor U1909 (N_1909,In_2523,In_1153);
or U1910 (N_1910,In_2046,In_1228);
or U1911 (N_1911,In_95,In_332);
nor U1912 (N_1912,In_1548,In_497);
and U1913 (N_1913,In_1556,In_511);
nand U1914 (N_1914,In_713,In_2677);
nor U1915 (N_1915,In_1322,In_1467);
nor U1916 (N_1916,In_1594,In_1867);
and U1917 (N_1917,In_1864,In_93);
or U1918 (N_1918,In_1976,In_1209);
nand U1919 (N_1919,In_536,In_588);
nand U1920 (N_1920,In_2633,In_1755);
xor U1921 (N_1921,In_325,In_1437);
nor U1922 (N_1922,In_1605,In_328);
nand U1923 (N_1923,In_1186,In_1981);
and U1924 (N_1924,In_1711,In_1908);
nor U1925 (N_1925,In_1922,In_2124);
nand U1926 (N_1926,In_161,In_275);
and U1927 (N_1927,In_2523,In_1396);
xnor U1928 (N_1928,In_945,In_2744);
nand U1929 (N_1929,In_2662,In_2669);
xnor U1930 (N_1930,In_2203,In_1402);
nor U1931 (N_1931,In_619,In_1853);
nor U1932 (N_1932,In_2733,In_748);
xor U1933 (N_1933,In_1852,In_2934);
or U1934 (N_1934,In_1022,In_709);
nand U1935 (N_1935,In_6,In_247);
nand U1936 (N_1936,In_459,In_2606);
xor U1937 (N_1937,In_212,In_1907);
xnor U1938 (N_1938,In_1102,In_2781);
or U1939 (N_1939,In_1962,In_2344);
nand U1940 (N_1940,In_244,In_341);
nor U1941 (N_1941,In_1594,In_2806);
nor U1942 (N_1942,In_1760,In_2869);
and U1943 (N_1943,In_2167,In_1372);
nor U1944 (N_1944,In_2874,In_2689);
and U1945 (N_1945,In_2742,In_2643);
or U1946 (N_1946,In_1251,In_757);
xor U1947 (N_1947,In_1173,In_890);
nand U1948 (N_1948,In_2268,In_1719);
nor U1949 (N_1949,In_911,In_178);
or U1950 (N_1950,In_1478,In_1810);
xor U1951 (N_1951,In_2245,In_2592);
nand U1952 (N_1952,In_2615,In_769);
nor U1953 (N_1953,In_2772,In_2832);
xnor U1954 (N_1954,In_1855,In_1545);
and U1955 (N_1955,In_1742,In_657);
and U1956 (N_1956,In_1145,In_2082);
nor U1957 (N_1957,In_388,In_501);
and U1958 (N_1958,In_2299,In_2103);
nor U1959 (N_1959,In_1573,In_1594);
nor U1960 (N_1960,In_1099,In_2645);
and U1961 (N_1961,In_1993,In_579);
nand U1962 (N_1962,In_5,In_2151);
or U1963 (N_1963,In_2878,In_206);
and U1964 (N_1964,In_1508,In_1470);
xnor U1965 (N_1965,In_2421,In_1574);
and U1966 (N_1966,In_2150,In_1592);
nand U1967 (N_1967,In_2282,In_315);
nor U1968 (N_1968,In_278,In_1372);
and U1969 (N_1969,In_1987,In_433);
and U1970 (N_1970,In_1142,In_1863);
and U1971 (N_1971,In_2394,In_1763);
nor U1972 (N_1972,In_2533,In_484);
and U1973 (N_1973,In_1695,In_734);
xnor U1974 (N_1974,In_630,In_948);
nand U1975 (N_1975,In_1376,In_1808);
and U1976 (N_1976,In_2281,In_1487);
and U1977 (N_1977,In_2413,In_2150);
xor U1978 (N_1978,In_692,In_2842);
nand U1979 (N_1979,In_1968,In_2646);
xor U1980 (N_1980,In_2089,In_378);
xnor U1981 (N_1981,In_1131,In_2927);
and U1982 (N_1982,In_1595,In_692);
nor U1983 (N_1983,In_1425,In_1725);
xnor U1984 (N_1984,In_2162,In_1356);
nand U1985 (N_1985,In_1778,In_97);
nand U1986 (N_1986,In_735,In_611);
or U1987 (N_1987,In_1019,In_2623);
xor U1988 (N_1988,In_1481,In_292);
and U1989 (N_1989,In_1099,In_1046);
xor U1990 (N_1990,In_1257,In_1832);
nor U1991 (N_1991,In_2218,In_1142);
xor U1992 (N_1992,In_1891,In_1976);
xnor U1993 (N_1993,In_132,In_1255);
xor U1994 (N_1994,In_6,In_2556);
and U1995 (N_1995,In_1352,In_1285);
xnor U1996 (N_1996,In_2144,In_1961);
and U1997 (N_1997,In_2875,In_105);
or U1998 (N_1998,In_1656,In_886);
xor U1999 (N_1999,In_274,In_1606);
xor U2000 (N_2000,In_1478,In_1489);
and U2001 (N_2001,In_2957,In_946);
and U2002 (N_2002,In_2636,In_1625);
and U2003 (N_2003,In_1348,In_100);
and U2004 (N_2004,In_475,In_2440);
xnor U2005 (N_2005,In_795,In_1739);
and U2006 (N_2006,In_981,In_2812);
and U2007 (N_2007,In_1015,In_1773);
xor U2008 (N_2008,In_2224,In_2255);
nand U2009 (N_2009,In_1935,In_2995);
xor U2010 (N_2010,In_2724,In_1093);
nor U2011 (N_2011,In_1491,In_2539);
nor U2012 (N_2012,In_773,In_1880);
nor U2013 (N_2013,In_1481,In_2119);
nand U2014 (N_2014,In_608,In_628);
and U2015 (N_2015,In_1926,In_1927);
nor U2016 (N_2016,In_1363,In_2298);
xor U2017 (N_2017,In_1738,In_2356);
nor U2018 (N_2018,In_2872,In_1641);
nand U2019 (N_2019,In_1819,In_69);
and U2020 (N_2020,In_935,In_2594);
xnor U2021 (N_2021,In_1004,In_321);
and U2022 (N_2022,In_1750,In_1865);
and U2023 (N_2023,In_2623,In_638);
nand U2024 (N_2024,In_2492,In_1318);
or U2025 (N_2025,In_131,In_1489);
and U2026 (N_2026,In_252,In_2753);
xnor U2027 (N_2027,In_776,In_1778);
xnor U2028 (N_2028,In_473,In_1371);
and U2029 (N_2029,In_96,In_2924);
nand U2030 (N_2030,In_449,In_1750);
nor U2031 (N_2031,In_842,In_1309);
nand U2032 (N_2032,In_1354,In_2772);
xor U2033 (N_2033,In_2945,In_431);
and U2034 (N_2034,In_1236,In_1295);
xor U2035 (N_2035,In_756,In_773);
or U2036 (N_2036,In_1841,In_641);
nand U2037 (N_2037,In_1603,In_679);
or U2038 (N_2038,In_1723,In_193);
and U2039 (N_2039,In_2117,In_2306);
nand U2040 (N_2040,In_1851,In_736);
and U2041 (N_2041,In_2854,In_842);
and U2042 (N_2042,In_2602,In_850);
and U2043 (N_2043,In_1690,In_187);
and U2044 (N_2044,In_2878,In_686);
and U2045 (N_2045,In_2981,In_1743);
or U2046 (N_2046,In_856,In_1704);
and U2047 (N_2047,In_1649,In_2671);
nand U2048 (N_2048,In_1931,In_1481);
nand U2049 (N_2049,In_482,In_1571);
and U2050 (N_2050,In_849,In_2788);
or U2051 (N_2051,In_1842,In_1723);
nor U2052 (N_2052,In_1348,In_212);
or U2053 (N_2053,In_1464,In_1184);
or U2054 (N_2054,In_517,In_2845);
nand U2055 (N_2055,In_1866,In_671);
and U2056 (N_2056,In_879,In_1662);
and U2057 (N_2057,In_1515,In_2325);
nor U2058 (N_2058,In_1091,In_1251);
and U2059 (N_2059,In_2399,In_1771);
xor U2060 (N_2060,In_2562,In_2111);
xor U2061 (N_2061,In_2714,In_2097);
or U2062 (N_2062,In_2774,In_717);
or U2063 (N_2063,In_1519,In_2273);
xnor U2064 (N_2064,In_1036,In_2150);
nor U2065 (N_2065,In_682,In_2223);
nand U2066 (N_2066,In_2123,In_2637);
xnor U2067 (N_2067,In_504,In_331);
or U2068 (N_2068,In_479,In_2740);
or U2069 (N_2069,In_2869,In_2727);
or U2070 (N_2070,In_1811,In_2923);
xnor U2071 (N_2071,In_2493,In_2048);
nor U2072 (N_2072,In_1502,In_519);
xnor U2073 (N_2073,In_160,In_1784);
and U2074 (N_2074,In_2722,In_2561);
nor U2075 (N_2075,In_2537,In_698);
nor U2076 (N_2076,In_607,In_2685);
nor U2077 (N_2077,In_2767,In_2092);
or U2078 (N_2078,In_847,In_559);
or U2079 (N_2079,In_2861,In_1353);
nand U2080 (N_2080,In_1685,In_580);
nand U2081 (N_2081,In_1429,In_356);
xnor U2082 (N_2082,In_1232,In_975);
xor U2083 (N_2083,In_1236,In_896);
nor U2084 (N_2084,In_608,In_1731);
or U2085 (N_2085,In_2074,In_2739);
nor U2086 (N_2086,In_1661,In_75);
xor U2087 (N_2087,In_2239,In_778);
nand U2088 (N_2088,In_2544,In_861);
nand U2089 (N_2089,In_2379,In_489);
and U2090 (N_2090,In_401,In_435);
nor U2091 (N_2091,In_843,In_2807);
nor U2092 (N_2092,In_441,In_2569);
nand U2093 (N_2093,In_1366,In_2316);
nand U2094 (N_2094,In_723,In_2716);
or U2095 (N_2095,In_1833,In_926);
and U2096 (N_2096,In_272,In_417);
or U2097 (N_2097,In_1432,In_1184);
xnor U2098 (N_2098,In_1909,In_2120);
or U2099 (N_2099,In_467,In_37);
and U2100 (N_2100,In_1782,In_1995);
or U2101 (N_2101,In_1676,In_1388);
nor U2102 (N_2102,In_2351,In_1572);
xor U2103 (N_2103,In_1446,In_2712);
and U2104 (N_2104,In_215,In_2449);
or U2105 (N_2105,In_1848,In_2478);
nand U2106 (N_2106,In_2937,In_2355);
or U2107 (N_2107,In_476,In_174);
xnor U2108 (N_2108,In_1290,In_720);
nor U2109 (N_2109,In_1460,In_1543);
nor U2110 (N_2110,In_564,In_2192);
and U2111 (N_2111,In_2823,In_1741);
and U2112 (N_2112,In_2302,In_1509);
or U2113 (N_2113,In_1836,In_2741);
or U2114 (N_2114,In_680,In_958);
nor U2115 (N_2115,In_605,In_2962);
and U2116 (N_2116,In_660,In_686);
xor U2117 (N_2117,In_537,In_1982);
nor U2118 (N_2118,In_381,In_2047);
nand U2119 (N_2119,In_726,In_926);
nor U2120 (N_2120,In_213,In_70);
and U2121 (N_2121,In_749,In_2526);
or U2122 (N_2122,In_1893,In_1662);
or U2123 (N_2123,In_2415,In_1096);
nand U2124 (N_2124,In_1003,In_2183);
xnor U2125 (N_2125,In_291,In_2449);
xnor U2126 (N_2126,In_2616,In_2751);
and U2127 (N_2127,In_1793,In_1851);
nand U2128 (N_2128,In_546,In_256);
xnor U2129 (N_2129,In_2730,In_1499);
and U2130 (N_2130,In_565,In_908);
nand U2131 (N_2131,In_2974,In_1505);
xnor U2132 (N_2132,In_2490,In_2666);
nor U2133 (N_2133,In_2915,In_1334);
or U2134 (N_2134,In_484,In_2310);
and U2135 (N_2135,In_1585,In_1175);
or U2136 (N_2136,In_1267,In_541);
nor U2137 (N_2137,In_230,In_2803);
nand U2138 (N_2138,In_512,In_2173);
and U2139 (N_2139,In_1358,In_2106);
and U2140 (N_2140,In_1469,In_2837);
nand U2141 (N_2141,In_255,In_2012);
nand U2142 (N_2142,In_715,In_2561);
xnor U2143 (N_2143,In_2183,In_265);
nand U2144 (N_2144,In_2923,In_1415);
and U2145 (N_2145,In_1420,In_946);
or U2146 (N_2146,In_2996,In_2391);
xor U2147 (N_2147,In_869,In_1570);
and U2148 (N_2148,In_2860,In_2835);
xor U2149 (N_2149,In_2300,In_1566);
and U2150 (N_2150,In_1248,In_472);
or U2151 (N_2151,In_1150,In_393);
xor U2152 (N_2152,In_1763,In_2548);
and U2153 (N_2153,In_1941,In_408);
and U2154 (N_2154,In_1648,In_914);
nand U2155 (N_2155,In_1833,In_2798);
nor U2156 (N_2156,In_914,In_1943);
or U2157 (N_2157,In_1700,In_1118);
and U2158 (N_2158,In_2314,In_609);
and U2159 (N_2159,In_1233,In_2640);
nor U2160 (N_2160,In_2991,In_196);
nor U2161 (N_2161,In_904,In_2984);
and U2162 (N_2162,In_1290,In_1661);
or U2163 (N_2163,In_2819,In_1587);
nand U2164 (N_2164,In_1193,In_393);
nand U2165 (N_2165,In_1083,In_994);
nor U2166 (N_2166,In_1850,In_1690);
nor U2167 (N_2167,In_2035,In_1863);
nand U2168 (N_2168,In_1309,In_1972);
nor U2169 (N_2169,In_41,In_1622);
nor U2170 (N_2170,In_725,In_2212);
or U2171 (N_2171,In_2528,In_1576);
and U2172 (N_2172,In_1219,In_1166);
and U2173 (N_2173,In_1645,In_2430);
nand U2174 (N_2174,In_852,In_1848);
nand U2175 (N_2175,In_2663,In_1883);
nand U2176 (N_2176,In_546,In_1380);
and U2177 (N_2177,In_1936,In_1593);
or U2178 (N_2178,In_1942,In_2760);
or U2179 (N_2179,In_1276,In_725);
or U2180 (N_2180,In_187,In_1069);
xor U2181 (N_2181,In_1800,In_962);
nor U2182 (N_2182,In_2540,In_153);
nand U2183 (N_2183,In_421,In_2022);
or U2184 (N_2184,In_1840,In_1957);
xnor U2185 (N_2185,In_1008,In_2266);
and U2186 (N_2186,In_2539,In_2165);
nand U2187 (N_2187,In_1174,In_496);
and U2188 (N_2188,In_184,In_1780);
nand U2189 (N_2189,In_378,In_578);
and U2190 (N_2190,In_1292,In_2621);
nor U2191 (N_2191,In_2450,In_2674);
nand U2192 (N_2192,In_297,In_2604);
and U2193 (N_2193,In_967,In_2223);
and U2194 (N_2194,In_2861,In_590);
nor U2195 (N_2195,In_2428,In_749);
xor U2196 (N_2196,In_471,In_1072);
xnor U2197 (N_2197,In_1220,In_2221);
nor U2198 (N_2198,In_2008,In_888);
nor U2199 (N_2199,In_666,In_2838);
nand U2200 (N_2200,In_1680,In_174);
and U2201 (N_2201,In_1221,In_2591);
or U2202 (N_2202,In_917,In_2443);
or U2203 (N_2203,In_2322,In_1259);
xor U2204 (N_2204,In_1268,In_2048);
xnor U2205 (N_2205,In_1888,In_2043);
and U2206 (N_2206,In_2404,In_189);
xor U2207 (N_2207,In_2428,In_2714);
nor U2208 (N_2208,In_525,In_1921);
and U2209 (N_2209,In_2751,In_920);
and U2210 (N_2210,In_775,In_1008);
or U2211 (N_2211,In_1084,In_1298);
nor U2212 (N_2212,In_1239,In_101);
nor U2213 (N_2213,In_567,In_629);
and U2214 (N_2214,In_2743,In_2637);
nor U2215 (N_2215,In_2962,In_329);
nand U2216 (N_2216,In_1404,In_2712);
nand U2217 (N_2217,In_2123,In_1844);
and U2218 (N_2218,In_2452,In_1666);
or U2219 (N_2219,In_1456,In_1366);
nand U2220 (N_2220,In_2337,In_302);
and U2221 (N_2221,In_155,In_2402);
nand U2222 (N_2222,In_703,In_1109);
xnor U2223 (N_2223,In_2960,In_2760);
xnor U2224 (N_2224,In_626,In_345);
xnor U2225 (N_2225,In_1990,In_2275);
nand U2226 (N_2226,In_2455,In_1551);
nand U2227 (N_2227,In_1333,In_1461);
and U2228 (N_2228,In_2658,In_2375);
or U2229 (N_2229,In_1708,In_1524);
xor U2230 (N_2230,In_809,In_2346);
or U2231 (N_2231,In_1786,In_2555);
xor U2232 (N_2232,In_1452,In_1456);
or U2233 (N_2233,In_2865,In_467);
nand U2234 (N_2234,In_1913,In_791);
and U2235 (N_2235,In_2739,In_2003);
and U2236 (N_2236,In_1453,In_1139);
nand U2237 (N_2237,In_398,In_618);
nor U2238 (N_2238,In_554,In_1483);
xor U2239 (N_2239,In_2500,In_987);
or U2240 (N_2240,In_1846,In_662);
xor U2241 (N_2241,In_2806,In_1004);
or U2242 (N_2242,In_746,In_370);
or U2243 (N_2243,In_1166,In_1920);
and U2244 (N_2244,In_2733,In_1252);
xnor U2245 (N_2245,In_189,In_145);
and U2246 (N_2246,In_613,In_12);
nand U2247 (N_2247,In_399,In_1469);
xor U2248 (N_2248,In_1009,In_403);
nand U2249 (N_2249,In_1618,In_2980);
and U2250 (N_2250,In_2944,In_2355);
or U2251 (N_2251,In_1153,In_1044);
nand U2252 (N_2252,In_1541,In_2328);
nand U2253 (N_2253,In_486,In_2930);
xnor U2254 (N_2254,In_2771,In_1482);
and U2255 (N_2255,In_2796,In_1320);
nand U2256 (N_2256,In_1636,In_558);
or U2257 (N_2257,In_1349,In_2762);
nor U2258 (N_2258,In_2417,In_2007);
nor U2259 (N_2259,In_1375,In_259);
nor U2260 (N_2260,In_490,In_1740);
and U2261 (N_2261,In_1462,In_333);
nand U2262 (N_2262,In_596,In_979);
or U2263 (N_2263,In_1964,In_572);
xor U2264 (N_2264,In_15,In_2970);
xnor U2265 (N_2265,In_2678,In_581);
or U2266 (N_2266,In_1349,In_10);
nand U2267 (N_2267,In_2415,In_578);
nand U2268 (N_2268,In_2660,In_654);
and U2269 (N_2269,In_1785,In_2226);
nor U2270 (N_2270,In_2883,In_1382);
xnor U2271 (N_2271,In_2420,In_1176);
and U2272 (N_2272,In_2113,In_2524);
nand U2273 (N_2273,In_350,In_2585);
xor U2274 (N_2274,In_2559,In_40);
nor U2275 (N_2275,In_1276,In_440);
or U2276 (N_2276,In_998,In_38);
or U2277 (N_2277,In_1748,In_2164);
nor U2278 (N_2278,In_2971,In_2548);
xor U2279 (N_2279,In_2806,In_49);
nand U2280 (N_2280,In_801,In_132);
xnor U2281 (N_2281,In_2099,In_1011);
or U2282 (N_2282,In_232,In_2651);
xnor U2283 (N_2283,In_799,In_245);
xnor U2284 (N_2284,In_649,In_1532);
xnor U2285 (N_2285,In_2358,In_2344);
nand U2286 (N_2286,In_1157,In_570);
nand U2287 (N_2287,In_2725,In_298);
xnor U2288 (N_2288,In_1942,In_1971);
or U2289 (N_2289,In_1561,In_2637);
nand U2290 (N_2290,In_695,In_647);
and U2291 (N_2291,In_935,In_2557);
nor U2292 (N_2292,In_2133,In_1127);
and U2293 (N_2293,In_1161,In_32);
xor U2294 (N_2294,In_653,In_775);
nand U2295 (N_2295,In_498,In_36);
or U2296 (N_2296,In_484,In_2458);
nor U2297 (N_2297,In_1520,In_2231);
xnor U2298 (N_2298,In_2948,In_2506);
xnor U2299 (N_2299,In_534,In_2609);
nand U2300 (N_2300,In_1899,In_2188);
nand U2301 (N_2301,In_1625,In_2640);
nor U2302 (N_2302,In_1832,In_1108);
nand U2303 (N_2303,In_1071,In_978);
nand U2304 (N_2304,In_2460,In_800);
or U2305 (N_2305,In_2524,In_2191);
and U2306 (N_2306,In_945,In_964);
nand U2307 (N_2307,In_1116,In_2954);
or U2308 (N_2308,In_433,In_2173);
and U2309 (N_2309,In_817,In_155);
xor U2310 (N_2310,In_2533,In_690);
nand U2311 (N_2311,In_2588,In_1883);
or U2312 (N_2312,In_2650,In_849);
nor U2313 (N_2313,In_2863,In_938);
and U2314 (N_2314,In_2314,In_1393);
or U2315 (N_2315,In_1549,In_879);
nor U2316 (N_2316,In_1996,In_1416);
or U2317 (N_2317,In_2462,In_872);
nand U2318 (N_2318,In_910,In_2081);
nor U2319 (N_2319,In_439,In_2858);
xnor U2320 (N_2320,In_196,In_2216);
nand U2321 (N_2321,In_2930,In_2088);
and U2322 (N_2322,In_2475,In_2260);
nand U2323 (N_2323,In_2417,In_240);
or U2324 (N_2324,In_885,In_1078);
xnor U2325 (N_2325,In_1189,In_890);
and U2326 (N_2326,In_1957,In_1334);
or U2327 (N_2327,In_2578,In_1813);
or U2328 (N_2328,In_1184,In_133);
and U2329 (N_2329,In_320,In_1199);
and U2330 (N_2330,In_1612,In_1595);
nand U2331 (N_2331,In_751,In_1045);
xnor U2332 (N_2332,In_1997,In_416);
or U2333 (N_2333,In_1327,In_905);
xor U2334 (N_2334,In_1471,In_1374);
and U2335 (N_2335,In_1904,In_501);
and U2336 (N_2336,In_507,In_1155);
nand U2337 (N_2337,In_2122,In_2413);
nand U2338 (N_2338,In_1610,In_251);
or U2339 (N_2339,In_2804,In_1359);
or U2340 (N_2340,In_2704,In_1731);
nand U2341 (N_2341,In_196,In_994);
and U2342 (N_2342,In_2125,In_2206);
nand U2343 (N_2343,In_869,In_597);
xnor U2344 (N_2344,In_763,In_2361);
xor U2345 (N_2345,In_2874,In_120);
and U2346 (N_2346,In_1780,In_1551);
nand U2347 (N_2347,In_1666,In_540);
or U2348 (N_2348,In_800,In_165);
or U2349 (N_2349,In_1896,In_570);
nor U2350 (N_2350,In_1687,In_1207);
or U2351 (N_2351,In_2307,In_2692);
or U2352 (N_2352,In_690,In_1699);
nor U2353 (N_2353,In_2227,In_75);
nand U2354 (N_2354,In_259,In_2886);
nor U2355 (N_2355,In_2394,In_351);
xnor U2356 (N_2356,In_2620,In_492);
nor U2357 (N_2357,In_2718,In_972);
xnor U2358 (N_2358,In_228,In_990);
nor U2359 (N_2359,In_394,In_2077);
xor U2360 (N_2360,In_1599,In_335);
nand U2361 (N_2361,In_1316,In_2277);
or U2362 (N_2362,In_27,In_2801);
nand U2363 (N_2363,In_1266,In_1680);
xor U2364 (N_2364,In_752,In_1347);
xnor U2365 (N_2365,In_741,In_1035);
or U2366 (N_2366,In_2500,In_1233);
xnor U2367 (N_2367,In_1863,In_1862);
xnor U2368 (N_2368,In_1366,In_2396);
nand U2369 (N_2369,In_2782,In_2272);
xor U2370 (N_2370,In_2329,In_171);
nor U2371 (N_2371,In_521,In_2357);
nor U2372 (N_2372,In_2595,In_11);
xor U2373 (N_2373,In_1441,In_578);
or U2374 (N_2374,In_2384,In_1804);
nor U2375 (N_2375,In_1506,In_1162);
nand U2376 (N_2376,In_2942,In_2966);
nor U2377 (N_2377,In_11,In_2331);
xor U2378 (N_2378,In_261,In_792);
xor U2379 (N_2379,In_2528,In_1927);
xnor U2380 (N_2380,In_1204,In_1542);
xnor U2381 (N_2381,In_2411,In_2762);
xnor U2382 (N_2382,In_1252,In_1634);
nor U2383 (N_2383,In_400,In_438);
or U2384 (N_2384,In_670,In_673);
nor U2385 (N_2385,In_2960,In_1753);
nor U2386 (N_2386,In_1402,In_129);
nand U2387 (N_2387,In_102,In_228);
and U2388 (N_2388,In_1985,In_1203);
or U2389 (N_2389,In_1695,In_947);
nand U2390 (N_2390,In_2832,In_1294);
xnor U2391 (N_2391,In_2821,In_1600);
nor U2392 (N_2392,In_380,In_1777);
or U2393 (N_2393,In_2323,In_1601);
nor U2394 (N_2394,In_1230,In_1126);
and U2395 (N_2395,In_1269,In_2509);
nand U2396 (N_2396,In_2283,In_2556);
nor U2397 (N_2397,In_2887,In_1269);
or U2398 (N_2398,In_423,In_699);
xor U2399 (N_2399,In_1785,In_38);
nand U2400 (N_2400,In_187,In_1213);
and U2401 (N_2401,In_2271,In_312);
nor U2402 (N_2402,In_534,In_1485);
nor U2403 (N_2403,In_1173,In_581);
nand U2404 (N_2404,In_1173,In_2841);
nor U2405 (N_2405,In_1963,In_131);
xnor U2406 (N_2406,In_998,In_573);
nand U2407 (N_2407,In_2362,In_444);
and U2408 (N_2408,In_1203,In_2083);
xor U2409 (N_2409,In_1139,In_1268);
and U2410 (N_2410,In_1409,In_2412);
nor U2411 (N_2411,In_2171,In_2883);
or U2412 (N_2412,In_456,In_774);
nand U2413 (N_2413,In_1555,In_2530);
nor U2414 (N_2414,In_2566,In_474);
xor U2415 (N_2415,In_2153,In_2912);
and U2416 (N_2416,In_907,In_985);
xnor U2417 (N_2417,In_643,In_2086);
nand U2418 (N_2418,In_2232,In_1919);
or U2419 (N_2419,In_1366,In_2427);
and U2420 (N_2420,In_1847,In_598);
xnor U2421 (N_2421,In_1329,In_1964);
and U2422 (N_2422,In_1510,In_434);
nor U2423 (N_2423,In_1571,In_1504);
xor U2424 (N_2424,In_149,In_610);
nand U2425 (N_2425,In_68,In_262);
or U2426 (N_2426,In_2365,In_1458);
nand U2427 (N_2427,In_2906,In_30);
nand U2428 (N_2428,In_494,In_2793);
nand U2429 (N_2429,In_2801,In_1158);
or U2430 (N_2430,In_2914,In_2466);
xnor U2431 (N_2431,In_1753,In_2149);
and U2432 (N_2432,In_250,In_2835);
nand U2433 (N_2433,In_292,In_2701);
or U2434 (N_2434,In_1431,In_2271);
and U2435 (N_2435,In_2191,In_1294);
nor U2436 (N_2436,In_1382,In_1153);
and U2437 (N_2437,In_788,In_92);
nand U2438 (N_2438,In_1540,In_749);
nor U2439 (N_2439,In_738,In_1776);
xnor U2440 (N_2440,In_1279,In_1958);
xor U2441 (N_2441,In_1684,In_475);
and U2442 (N_2442,In_2901,In_663);
xor U2443 (N_2443,In_2497,In_37);
nand U2444 (N_2444,In_916,In_161);
or U2445 (N_2445,In_1537,In_858);
nor U2446 (N_2446,In_795,In_1204);
nor U2447 (N_2447,In_430,In_1906);
xnor U2448 (N_2448,In_2857,In_1448);
and U2449 (N_2449,In_64,In_1662);
nand U2450 (N_2450,In_1200,In_2730);
xnor U2451 (N_2451,In_2947,In_985);
and U2452 (N_2452,In_621,In_915);
nand U2453 (N_2453,In_240,In_153);
nor U2454 (N_2454,In_2416,In_2337);
xor U2455 (N_2455,In_135,In_105);
nor U2456 (N_2456,In_361,In_877);
nor U2457 (N_2457,In_765,In_2545);
nand U2458 (N_2458,In_756,In_1967);
nor U2459 (N_2459,In_2773,In_2670);
and U2460 (N_2460,In_1060,In_1260);
nand U2461 (N_2461,In_954,In_2431);
or U2462 (N_2462,In_1548,In_2797);
xor U2463 (N_2463,In_1681,In_1334);
nand U2464 (N_2464,In_2991,In_173);
xnor U2465 (N_2465,In_1362,In_2717);
nand U2466 (N_2466,In_2194,In_2059);
or U2467 (N_2467,In_709,In_2067);
nand U2468 (N_2468,In_2216,In_1011);
nand U2469 (N_2469,In_1627,In_1128);
xor U2470 (N_2470,In_1751,In_2285);
and U2471 (N_2471,In_1846,In_1121);
nor U2472 (N_2472,In_1971,In_537);
nor U2473 (N_2473,In_2674,In_1300);
xor U2474 (N_2474,In_1931,In_192);
or U2475 (N_2475,In_889,In_1484);
and U2476 (N_2476,In_598,In_1670);
or U2477 (N_2477,In_307,In_212);
xnor U2478 (N_2478,In_184,In_755);
nand U2479 (N_2479,In_62,In_2162);
nor U2480 (N_2480,In_770,In_1780);
nor U2481 (N_2481,In_1921,In_1394);
and U2482 (N_2482,In_2916,In_839);
nand U2483 (N_2483,In_1266,In_406);
or U2484 (N_2484,In_12,In_2015);
nand U2485 (N_2485,In_461,In_1202);
or U2486 (N_2486,In_1185,In_2806);
nor U2487 (N_2487,In_2137,In_743);
nor U2488 (N_2488,In_1772,In_2638);
and U2489 (N_2489,In_2147,In_1224);
nand U2490 (N_2490,In_206,In_327);
and U2491 (N_2491,In_2488,In_2740);
nand U2492 (N_2492,In_88,In_295);
xor U2493 (N_2493,In_2657,In_2842);
nand U2494 (N_2494,In_843,In_525);
and U2495 (N_2495,In_1091,In_889);
and U2496 (N_2496,In_2701,In_1602);
xnor U2497 (N_2497,In_1789,In_1339);
and U2498 (N_2498,In_1990,In_2501);
nor U2499 (N_2499,In_2137,In_2387);
and U2500 (N_2500,In_789,In_1553);
or U2501 (N_2501,In_1315,In_1340);
xor U2502 (N_2502,In_849,In_2866);
or U2503 (N_2503,In_2692,In_1565);
xnor U2504 (N_2504,In_1982,In_419);
xnor U2505 (N_2505,In_1912,In_2765);
nor U2506 (N_2506,In_481,In_1675);
and U2507 (N_2507,In_1348,In_2555);
nor U2508 (N_2508,In_575,In_872);
xnor U2509 (N_2509,In_474,In_2251);
xnor U2510 (N_2510,In_2042,In_496);
or U2511 (N_2511,In_2470,In_1602);
xnor U2512 (N_2512,In_2656,In_2474);
or U2513 (N_2513,In_2715,In_1934);
xor U2514 (N_2514,In_192,In_79);
xnor U2515 (N_2515,In_1986,In_1684);
xnor U2516 (N_2516,In_896,In_2431);
xnor U2517 (N_2517,In_1091,In_1004);
or U2518 (N_2518,In_737,In_921);
and U2519 (N_2519,In_2675,In_966);
or U2520 (N_2520,In_1276,In_163);
xor U2521 (N_2521,In_419,In_586);
nor U2522 (N_2522,In_1119,In_2500);
nand U2523 (N_2523,In_1729,In_1198);
xnor U2524 (N_2524,In_2369,In_147);
and U2525 (N_2525,In_1002,In_1086);
nand U2526 (N_2526,In_1078,In_1937);
and U2527 (N_2527,In_1749,In_2348);
or U2528 (N_2528,In_1813,In_266);
nand U2529 (N_2529,In_2834,In_635);
nor U2530 (N_2530,In_511,In_103);
nand U2531 (N_2531,In_2995,In_2790);
xor U2532 (N_2532,In_458,In_424);
and U2533 (N_2533,In_419,In_1825);
nand U2534 (N_2534,In_1963,In_758);
and U2535 (N_2535,In_2173,In_1066);
xnor U2536 (N_2536,In_2053,In_2250);
xor U2537 (N_2537,In_1523,In_1327);
nand U2538 (N_2538,In_2893,In_260);
nand U2539 (N_2539,In_2877,In_2287);
and U2540 (N_2540,In_508,In_1964);
xor U2541 (N_2541,In_388,In_487);
and U2542 (N_2542,In_383,In_1675);
or U2543 (N_2543,In_2685,In_2238);
or U2544 (N_2544,In_1527,In_120);
and U2545 (N_2545,In_1657,In_141);
or U2546 (N_2546,In_1275,In_2974);
nand U2547 (N_2547,In_2691,In_2365);
or U2548 (N_2548,In_1533,In_1305);
or U2549 (N_2549,In_391,In_2689);
nor U2550 (N_2550,In_2845,In_2219);
or U2551 (N_2551,In_2449,In_1039);
xnor U2552 (N_2552,In_2729,In_1431);
and U2553 (N_2553,In_1730,In_2023);
and U2554 (N_2554,In_249,In_2243);
xnor U2555 (N_2555,In_1443,In_796);
nand U2556 (N_2556,In_2241,In_1768);
and U2557 (N_2557,In_1059,In_64);
and U2558 (N_2558,In_1144,In_1824);
nor U2559 (N_2559,In_2036,In_878);
and U2560 (N_2560,In_638,In_255);
or U2561 (N_2561,In_930,In_2048);
nand U2562 (N_2562,In_1653,In_2631);
nand U2563 (N_2563,In_2422,In_861);
xor U2564 (N_2564,In_2413,In_2728);
or U2565 (N_2565,In_2501,In_1586);
or U2566 (N_2566,In_859,In_233);
xnor U2567 (N_2567,In_2275,In_224);
or U2568 (N_2568,In_666,In_442);
nor U2569 (N_2569,In_560,In_2857);
or U2570 (N_2570,In_2475,In_1671);
or U2571 (N_2571,In_1963,In_1426);
nor U2572 (N_2572,In_1032,In_247);
nor U2573 (N_2573,In_1499,In_2770);
nand U2574 (N_2574,In_2715,In_1000);
and U2575 (N_2575,In_1207,In_2175);
xor U2576 (N_2576,In_1880,In_452);
nand U2577 (N_2577,In_2836,In_2721);
xnor U2578 (N_2578,In_463,In_699);
nor U2579 (N_2579,In_588,In_1593);
and U2580 (N_2580,In_539,In_1975);
xnor U2581 (N_2581,In_859,In_2572);
or U2582 (N_2582,In_528,In_1626);
nor U2583 (N_2583,In_1622,In_1750);
nor U2584 (N_2584,In_2646,In_2107);
and U2585 (N_2585,In_1795,In_2927);
nor U2586 (N_2586,In_799,In_2457);
nor U2587 (N_2587,In_2109,In_1078);
nor U2588 (N_2588,In_2511,In_2603);
and U2589 (N_2589,In_2561,In_826);
nand U2590 (N_2590,In_15,In_87);
nand U2591 (N_2591,In_1077,In_1819);
nor U2592 (N_2592,In_2635,In_1469);
or U2593 (N_2593,In_2852,In_1545);
xnor U2594 (N_2594,In_462,In_1597);
xor U2595 (N_2595,In_1216,In_2938);
xnor U2596 (N_2596,In_2960,In_2941);
and U2597 (N_2597,In_1219,In_2341);
nand U2598 (N_2598,In_2291,In_1276);
nor U2599 (N_2599,In_11,In_2658);
xor U2600 (N_2600,In_2739,In_2101);
nand U2601 (N_2601,In_860,In_892);
xnor U2602 (N_2602,In_2450,In_82);
xnor U2603 (N_2603,In_1958,In_2096);
and U2604 (N_2604,In_1319,In_1955);
and U2605 (N_2605,In_2543,In_1646);
nand U2606 (N_2606,In_292,In_1555);
xor U2607 (N_2607,In_216,In_2123);
and U2608 (N_2608,In_789,In_1426);
or U2609 (N_2609,In_403,In_634);
and U2610 (N_2610,In_751,In_2713);
nand U2611 (N_2611,In_320,In_350);
or U2612 (N_2612,In_185,In_1703);
nand U2613 (N_2613,In_1179,In_2685);
nor U2614 (N_2614,In_1220,In_1563);
or U2615 (N_2615,In_2778,In_1913);
or U2616 (N_2616,In_2424,In_2821);
nor U2617 (N_2617,In_2555,In_421);
xnor U2618 (N_2618,In_2822,In_929);
nor U2619 (N_2619,In_2988,In_831);
or U2620 (N_2620,In_1972,In_155);
xor U2621 (N_2621,In_755,In_1184);
nand U2622 (N_2622,In_1539,In_1506);
nor U2623 (N_2623,In_2783,In_385);
nor U2624 (N_2624,In_1894,In_345);
xnor U2625 (N_2625,In_599,In_293);
or U2626 (N_2626,In_412,In_2834);
and U2627 (N_2627,In_609,In_1905);
or U2628 (N_2628,In_2561,In_565);
nand U2629 (N_2629,In_1939,In_2081);
or U2630 (N_2630,In_939,In_2585);
or U2631 (N_2631,In_1389,In_1701);
and U2632 (N_2632,In_2540,In_2216);
nand U2633 (N_2633,In_1037,In_552);
nor U2634 (N_2634,In_2638,In_1263);
or U2635 (N_2635,In_2701,In_412);
and U2636 (N_2636,In_2099,In_1699);
nand U2637 (N_2637,In_1794,In_1445);
nand U2638 (N_2638,In_2788,In_1342);
or U2639 (N_2639,In_988,In_1045);
xnor U2640 (N_2640,In_2623,In_333);
and U2641 (N_2641,In_2927,In_873);
and U2642 (N_2642,In_1195,In_1341);
and U2643 (N_2643,In_1461,In_2146);
xnor U2644 (N_2644,In_1157,In_1404);
and U2645 (N_2645,In_39,In_1161);
nand U2646 (N_2646,In_912,In_1730);
and U2647 (N_2647,In_87,In_199);
nor U2648 (N_2648,In_267,In_1098);
nand U2649 (N_2649,In_444,In_1982);
nand U2650 (N_2650,In_1743,In_260);
and U2651 (N_2651,In_2214,In_2978);
or U2652 (N_2652,In_1427,In_1363);
nand U2653 (N_2653,In_2208,In_1942);
xor U2654 (N_2654,In_940,In_315);
nor U2655 (N_2655,In_2721,In_1993);
xor U2656 (N_2656,In_167,In_1252);
or U2657 (N_2657,In_619,In_750);
and U2658 (N_2658,In_2361,In_1485);
xnor U2659 (N_2659,In_2081,In_1379);
and U2660 (N_2660,In_1903,In_971);
nand U2661 (N_2661,In_1142,In_633);
and U2662 (N_2662,In_2267,In_1859);
xor U2663 (N_2663,In_1338,In_1697);
or U2664 (N_2664,In_1205,In_1440);
nand U2665 (N_2665,In_1683,In_2578);
and U2666 (N_2666,In_1587,In_2319);
or U2667 (N_2667,In_47,In_1115);
or U2668 (N_2668,In_2149,In_2907);
xor U2669 (N_2669,In_201,In_818);
and U2670 (N_2670,In_2828,In_2166);
and U2671 (N_2671,In_291,In_2613);
xor U2672 (N_2672,In_2855,In_1432);
xor U2673 (N_2673,In_440,In_2745);
nand U2674 (N_2674,In_1852,In_109);
xor U2675 (N_2675,In_2632,In_1478);
nor U2676 (N_2676,In_736,In_2341);
nand U2677 (N_2677,In_215,In_2506);
and U2678 (N_2678,In_846,In_189);
or U2679 (N_2679,In_392,In_538);
or U2680 (N_2680,In_643,In_1922);
or U2681 (N_2681,In_864,In_554);
and U2682 (N_2682,In_951,In_2016);
nand U2683 (N_2683,In_378,In_888);
nor U2684 (N_2684,In_2100,In_2198);
or U2685 (N_2685,In_2265,In_1303);
or U2686 (N_2686,In_2374,In_2795);
nor U2687 (N_2687,In_2119,In_1942);
or U2688 (N_2688,In_1615,In_1921);
or U2689 (N_2689,In_2738,In_1586);
and U2690 (N_2690,In_2080,In_852);
and U2691 (N_2691,In_2348,In_1885);
nor U2692 (N_2692,In_448,In_1307);
xnor U2693 (N_2693,In_1807,In_2148);
xor U2694 (N_2694,In_2754,In_1885);
xnor U2695 (N_2695,In_667,In_2259);
and U2696 (N_2696,In_2372,In_2988);
or U2697 (N_2697,In_1616,In_1360);
and U2698 (N_2698,In_150,In_703);
or U2699 (N_2699,In_74,In_473);
nand U2700 (N_2700,In_748,In_2508);
and U2701 (N_2701,In_1281,In_364);
nand U2702 (N_2702,In_537,In_1335);
nor U2703 (N_2703,In_434,In_222);
and U2704 (N_2704,In_2351,In_637);
and U2705 (N_2705,In_2526,In_2984);
nand U2706 (N_2706,In_1722,In_398);
xor U2707 (N_2707,In_2123,In_1782);
or U2708 (N_2708,In_1517,In_920);
nand U2709 (N_2709,In_44,In_203);
and U2710 (N_2710,In_2989,In_1728);
and U2711 (N_2711,In_2970,In_2270);
and U2712 (N_2712,In_891,In_256);
or U2713 (N_2713,In_601,In_1517);
and U2714 (N_2714,In_2001,In_2708);
nor U2715 (N_2715,In_933,In_2192);
xnor U2716 (N_2716,In_817,In_947);
or U2717 (N_2717,In_2319,In_1012);
nand U2718 (N_2718,In_145,In_479);
and U2719 (N_2719,In_744,In_1822);
xnor U2720 (N_2720,In_137,In_1306);
and U2721 (N_2721,In_2273,In_2846);
and U2722 (N_2722,In_2542,In_2844);
nor U2723 (N_2723,In_500,In_1010);
nand U2724 (N_2724,In_2400,In_2012);
nand U2725 (N_2725,In_902,In_803);
nor U2726 (N_2726,In_2217,In_1839);
and U2727 (N_2727,In_167,In_2496);
xor U2728 (N_2728,In_1803,In_2426);
nor U2729 (N_2729,In_405,In_953);
and U2730 (N_2730,In_2983,In_1232);
nor U2731 (N_2731,In_244,In_162);
and U2732 (N_2732,In_2205,In_168);
xnor U2733 (N_2733,In_1172,In_637);
or U2734 (N_2734,In_1857,In_2699);
xor U2735 (N_2735,In_577,In_2178);
or U2736 (N_2736,In_2939,In_2776);
xor U2737 (N_2737,In_2589,In_2720);
and U2738 (N_2738,In_1732,In_660);
nor U2739 (N_2739,In_615,In_927);
xor U2740 (N_2740,In_810,In_2294);
or U2741 (N_2741,In_2684,In_945);
nand U2742 (N_2742,In_2808,In_2073);
xnor U2743 (N_2743,In_2084,In_255);
xor U2744 (N_2744,In_175,In_1674);
nor U2745 (N_2745,In_938,In_2427);
nor U2746 (N_2746,In_1907,In_2673);
nor U2747 (N_2747,In_2397,In_2791);
and U2748 (N_2748,In_2084,In_348);
nand U2749 (N_2749,In_2170,In_2293);
xnor U2750 (N_2750,In_1133,In_1234);
nor U2751 (N_2751,In_1751,In_141);
or U2752 (N_2752,In_1199,In_1920);
xor U2753 (N_2753,In_120,In_1896);
nor U2754 (N_2754,In_2077,In_504);
nor U2755 (N_2755,In_2040,In_1320);
xor U2756 (N_2756,In_1557,In_821);
and U2757 (N_2757,In_2265,In_1626);
nor U2758 (N_2758,In_2257,In_546);
and U2759 (N_2759,In_2415,In_126);
nor U2760 (N_2760,In_874,In_1242);
nor U2761 (N_2761,In_2922,In_221);
nand U2762 (N_2762,In_985,In_2012);
xor U2763 (N_2763,In_2618,In_1149);
xnor U2764 (N_2764,In_2870,In_817);
nor U2765 (N_2765,In_1833,In_1904);
nand U2766 (N_2766,In_1605,In_1549);
xor U2767 (N_2767,In_1041,In_1668);
xnor U2768 (N_2768,In_1477,In_2228);
nor U2769 (N_2769,In_546,In_1761);
or U2770 (N_2770,In_1073,In_1908);
and U2771 (N_2771,In_2753,In_1616);
and U2772 (N_2772,In_2516,In_1313);
xor U2773 (N_2773,In_2675,In_2786);
nand U2774 (N_2774,In_946,In_1617);
and U2775 (N_2775,In_1748,In_2770);
nand U2776 (N_2776,In_2435,In_2780);
or U2777 (N_2777,In_163,In_51);
xnor U2778 (N_2778,In_1983,In_116);
and U2779 (N_2779,In_2068,In_64);
xor U2780 (N_2780,In_1011,In_1216);
and U2781 (N_2781,In_1237,In_2315);
nor U2782 (N_2782,In_695,In_2562);
xor U2783 (N_2783,In_1952,In_984);
or U2784 (N_2784,In_2729,In_1988);
nand U2785 (N_2785,In_1860,In_398);
xor U2786 (N_2786,In_2005,In_2922);
xor U2787 (N_2787,In_845,In_1689);
nand U2788 (N_2788,In_1708,In_1789);
or U2789 (N_2789,In_2057,In_195);
xor U2790 (N_2790,In_1325,In_862);
xor U2791 (N_2791,In_2910,In_2316);
or U2792 (N_2792,In_2319,In_56);
or U2793 (N_2793,In_391,In_2263);
and U2794 (N_2794,In_2431,In_1260);
xnor U2795 (N_2795,In_1062,In_879);
and U2796 (N_2796,In_2864,In_636);
nand U2797 (N_2797,In_1000,In_1623);
and U2798 (N_2798,In_1797,In_958);
xor U2799 (N_2799,In_916,In_2023);
nor U2800 (N_2800,In_1924,In_1969);
or U2801 (N_2801,In_2414,In_118);
nand U2802 (N_2802,In_2375,In_1450);
nand U2803 (N_2803,In_2504,In_646);
xnor U2804 (N_2804,In_1214,In_1854);
nand U2805 (N_2805,In_2556,In_1337);
and U2806 (N_2806,In_1339,In_0);
and U2807 (N_2807,In_1476,In_751);
nand U2808 (N_2808,In_520,In_2840);
nor U2809 (N_2809,In_1632,In_404);
nand U2810 (N_2810,In_2280,In_871);
nor U2811 (N_2811,In_398,In_2604);
xnor U2812 (N_2812,In_983,In_2045);
or U2813 (N_2813,In_797,In_1849);
xor U2814 (N_2814,In_2032,In_212);
or U2815 (N_2815,In_677,In_2974);
nand U2816 (N_2816,In_1135,In_2804);
or U2817 (N_2817,In_1137,In_465);
nand U2818 (N_2818,In_1132,In_818);
xnor U2819 (N_2819,In_712,In_848);
xor U2820 (N_2820,In_292,In_2164);
or U2821 (N_2821,In_366,In_1285);
nor U2822 (N_2822,In_306,In_2281);
xnor U2823 (N_2823,In_1258,In_467);
and U2824 (N_2824,In_1769,In_2425);
nor U2825 (N_2825,In_947,In_1052);
and U2826 (N_2826,In_711,In_782);
nand U2827 (N_2827,In_40,In_422);
xnor U2828 (N_2828,In_2916,In_1280);
xor U2829 (N_2829,In_903,In_323);
and U2830 (N_2830,In_2264,In_2746);
or U2831 (N_2831,In_2826,In_2728);
xor U2832 (N_2832,In_2414,In_2604);
and U2833 (N_2833,In_1462,In_2285);
nor U2834 (N_2834,In_1414,In_2137);
xnor U2835 (N_2835,In_1013,In_2073);
xor U2836 (N_2836,In_521,In_2453);
nand U2837 (N_2837,In_2152,In_618);
nor U2838 (N_2838,In_2699,In_636);
nand U2839 (N_2839,In_465,In_2068);
xnor U2840 (N_2840,In_1338,In_2805);
xnor U2841 (N_2841,In_1752,In_661);
xnor U2842 (N_2842,In_1259,In_2353);
or U2843 (N_2843,In_2260,In_1903);
nand U2844 (N_2844,In_1041,In_319);
nand U2845 (N_2845,In_1981,In_2696);
nor U2846 (N_2846,In_282,In_2180);
xor U2847 (N_2847,In_1725,In_1541);
or U2848 (N_2848,In_2751,In_2875);
nand U2849 (N_2849,In_1262,In_2523);
and U2850 (N_2850,In_792,In_1469);
and U2851 (N_2851,In_1498,In_701);
or U2852 (N_2852,In_2626,In_101);
or U2853 (N_2853,In_2703,In_503);
xnor U2854 (N_2854,In_1402,In_611);
and U2855 (N_2855,In_1372,In_1563);
nand U2856 (N_2856,In_1225,In_2338);
or U2857 (N_2857,In_328,In_342);
nor U2858 (N_2858,In_2196,In_173);
and U2859 (N_2859,In_2984,In_2575);
and U2860 (N_2860,In_2343,In_2306);
nor U2861 (N_2861,In_1101,In_356);
and U2862 (N_2862,In_2430,In_2286);
or U2863 (N_2863,In_2439,In_938);
or U2864 (N_2864,In_1682,In_1031);
nand U2865 (N_2865,In_606,In_1386);
nand U2866 (N_2866,In_1564,In_2839);
nand U2867 (N_2867,In_1543,In_2336);
xnor U2868 (N_2868,In_1741,In_1985);
or U2869 (N_2869,In_2752,In_1061);
xor U2870 (N_2870,In_2680,In_291);
and U2871 (N_2871,In_1865,In_346);
nor U2872 (N_2872,In_1640,In_1970);
nor U2873 (N_2873,In_339,In_1458);
and U2874 (N_2874,In_1770,In_1797);
nand U2875 (N_2875,In_53,In_478);
nand U2876 (N_2876,In_2171,In_2676);
nor U2877 (N_2877,In_2088,In_1526);
nand U2878 (N_2878,In_726,In_326);
nor U2879 (N_2879,In_889,In_1101);
or U2880 (N_2880,In_2186,In_2471);
and U2881 (N_2881,In_2675,In_313);
nand U2882 (N_2882,In_1482,In_2916);
and U2883 (N_2883,In_2921,In_1151);
xor U2884 (N_2884,In_301,In_2236);
xnor U2885 (N_2885,In_2540,In_465);
xor U2886 (N_2886,In_1864,In_1162);
and U2887 (N_2887,In_1430,In_1504);
and U2888 (N_2888,In_2511,In_2619);
or U2889 (N_2889,In_1492,In_1956);
xor U2890 (N_2890,In_2411,In_2509);
xnor U2891 (N_2891,In_1253,In_2328);
xnor U2892 (N_2892,In_608,In_1135);
and U2893 (N_2893,In_1512,In_1471);
nand U2894 (N_2894,In_329,In_2081);
nand U2895 (N_2895,In_983,In_1781);
xnor U2896 (N_2896,In_474,In_2516);
and U2897 (N_2897,In_174,In_1848);
or U2898 (N_2898,In_1155,In_2552);
xnor U2899 (N_2899,In_1700,In_2610);
or U2900 (N_2900,In_938,In_1860);
xnor U2901 (N_2901,In_637,In_946);
and U2902 (N_2902,In_1765,In_1062);
xor U2903 (N_2903,In_708,In_982);
or U2904 (N_2904,In_1958,In_2932);
xnor U2905 (N_2905,In_1771,In_955);
nor U2906 (N_2906,In_1410,In_2547);
xor U2907 (N_2907,In_1332,In_1949);
and U2908 (N_2908,In_1668,In_1046);
and U2909 (N_2909,In_711,In_2277);
nor U2910 (N_2910,In_2832,In_1634);
and U2911 (N_2911,In_944,In_2106);
and U2912 (N_2912,In_1325,In_1553);
xor U2913 (N_2913,In_1976,In_2939);
or U2914 (N_2914,In_1754,In_1618);
nand U2915 (N_2915,In_685,In_1664);
and U2916 (N_2916,In_2948,In_575);
xor U2917 (N_2917,In_1426,In_131);
or U2918 (N_2918,In_1184,In_1842);
nand U2919 (N_2919,In_2985,In_709);
xor U2920 (N_2920,In_1301,In_2181);
and U2921 (N_2921,In_1602,In_1567);
nor U2922 (N_2922,In_126,In_1697);
nor U2923 (N_2923,In_647,In_736);
nor U2924 (N_2924,In_1021,In_2438);
nand U2925 (N_2925,In_893,In_1637);
xor U2926 (N_2926,In_1993,In_266);
nor U2927 (N_2927,In_1455,In_1704);
xnor U2928 (N_2928,In_169,In_1970);
nor U2929 (N_2929,In_17,In_810);
or U2930 (N_2930,In_2268,In_541);
and U2931 (N_2931,In_1277,In_1201);
nand U2932 (N_2932,In_2502,In_1119);
nand U2933 (N_2933,In_607,In_2760);
nor U2934 (N_2934,In_759,In_720);
nand U2935 (N_2935,In_608,In_2415);
xnor U2936 (N_2936,In_2943,In_273);
or U2937 (N_2937,In_1584,In_1116);
nor U2938 (N_2938,In_2800,In_2799);
nand U2939 (N_2939,In_2804,In_2595);
nand U2940 (N_2940,In_1413,In_1764);
and U2941 (N_2941,In_775,In_524);
nand U2942 (N_2942,In_2802,In_2377);
or U2943 (N_2943,In_985,In_95);
nand U2944 (N_2944,In_462,In_2853);
nor U2945 (N_2945,In_2937,In_294);
or U2946 (N_2946,In_2446,In_2501);
nor U2947 (N_2947,In_420,In_461);
xor U2948 (N_2948,In_962,In_2220);
nor U2949 (N_2949,In_1665,In_2412);
nor U2950 (N_2950,In_812,In_1697);
xor U2951 (N_2951,In_2266,In_2026);
or U2952 (N_2952,In_1131,In_987);
and U2953 (N_2953,In_58,In_946);
or U2954 (N_2954,In_86,In_2890);
xor U2955 (N_2955,In_1093,In_2113);
or U2956 (N_2956,In_1225,In_2014);
xnor U2957 (N_2957,In_1312,In_2023);
and U2958 (N_2958,In_2158,In_1104);
and U2959 (N_2959,In_963,In_173);
or U2960 (N_2960,In_734,In_1036);
nor U2961 (N_2961,In_2481,In_473);
xnor U2962 (N_2962,In_1286,In_2224);
nand U2963 (N_2963,In_176,In_2647);
nand U2964 (N_2964,In_227,In_800);
nor U2965 (N_2965,In_2533,In_2633);
xor U2966 (N_2966,In_2328,In_2720);
nand U2967 (N_2967,In_1639,In_1513);
xnor U2968 (N_2968,In_2969,In_1189);
and U2969 (N_2969,In_1253,In_869);
xor U2970 (N_2970,In_2953,In_17);
xnor U2971 (N_2971,In_620,In_697);
nand U2972 (N_2972,In_872,In_346);
xor U2973 (N_2973,In_2092,In_1840);
nor U2974 (N_2974,In_2370,In_2223);
nor U2975 (N_2975,In_227,In_2681);
xnor U2976 (N_2976,In_1789,In_2192);
xnor U2977 (N_2977,In_2061,In_2392);
nand U2978 (N_2978,In_88,In_1874);
and U2979 (N_2979,In_959,In_2041);
nor U2980 (N_2980,In_2091,In_1939);
or U2981 (N_2981,In_299,In_1800);
xor U2982 (N_2982,In_1806,In_2881);
or U2983 (N_2983,In_571,In_1310);
xnor U2984 (N_2984,In_1224,In_298);
and U2985 (N_2985,In_2808,In_664);
and U2986 (N_2986,In_430,In_414);
or U2987 (N_2987,In_1501,In_920);
xnor U2988 (N_2988,In_1082,In_2513);
nand U2989 (N_2989,In_2734,In_1377);
or U2990 (N_2990,In_2517,In_2526);
or U2991 (N_2991,In_2396,In_2677);
xor U2992 (N_2992,In_2678,In_1241);
or U2993 (N_2993,In_1535,In_661);
nand U2994 (N_2994,In_1295,In_1461);
or U2995 (N_2995,In_192,In_1348);
and U2996 (N_2996,In_1322,In_1281);
or U2997 (N_2997,In_920,In_437);
and U2998 (N_2998,In_1102,In_244);
nand U2999 (N_2999,In_1793,In_2041);
or U3000 (N_3000,In_2188,In_17);
nor U3001 (N_3001,In_2580,In_1789);
and U3002 (N_3002,In_102,In_1707);
nor U3003 (N_3003,In_1040,In_694);
or U3004 (N_3004,In_2302,In_365);
xor U3005 (N_3005,In_973,In_1134);
xor U3006 (N_3006,In_2551,In_509);
nand U3007 (N_3007,In_1534,In_182);
and U3008 (N_3008,In_2113,In_1944);
nand U3009 (N_3009,In_2234,In_550);
or U3010 (N_3010,In_267,In_2509);
nor U3011 (N_3011,In_1667,In_2899);
nor U3012 (N_3012,In_2356,In_65);
or U3013 (N_3013,In_69,In_1990);
nand U3014 (N_3014,In_1911,In_29);
and U3015 (N_3015,In_1060,In_2402);
xnor U3016 (N_3016,In_295,In_2240);
and U3017 (N_3017,In_1161,In_2301);
or U3018 (N_3018,In_1756,In_1420);
nand U3019 (N_3019,In_1747,In_2196);
nor U3020 (N_3020,In_1670,In_1075);
nor U3021 (N_3021,In_2374,In_1344);
xor U3022 (N_3022,In_1231,In_930);
and U3023 (N_3023,In_391,In_289);
and U3024 (N_3024,In_1485,In_2718);
and U3025 (N_3025,In_2125,In_2523);
and U3026 (N_3026,In_1141,In_2374);
and U3027 (N_3027,In_700,In_573);
nor U3028 (N_3028,In_2308,In_2039);
and U3029 (N_3029,In_667,In_725);
xor U3030 (N_3030,In_1687,In_2428);
or U3031 (N_3031,In_2406,In_1261);
nor U3032 (N_3032,In_2635,In_800);
and U3033 (N_3033,In_236,In_1954);
xnor U3034 (N_3034,In_876,In_2029);
and U3035 (N_3035,In_946,In_2099);
and U3036 (N_3036,In_453,In_344);
or U3037 (N_3037,In_1001,In_2122);
nand U3038 (N_3038,In_1264,In_2361);
nor U3039 (N_3039,In_1524,In_104);
nor U3040 (N_3040,In_1719,In_1543);
xor U3041 (N_3041,In_2684,In_911);
or U3042 (N_3042,In_2934,In_1315);
and U3043 (N_3043,In_2861,In_1486);
or U3044 (N_3044,In_1107,In_2331);
nor U3045 (N_3045,In_685,In_798);
or U3046 (N_3046,In_899,In_174);
nor U3047 (N_3047,In_1543,In_2797);
and U3048 (N_3048,In_2478,In_510);
nand U3049 (N_3049,In_1702,In_2110);
nor U3050 (N_3050,In_2797,In_292);
nor U3051 (N_3051,In_969,In_804);
xnor U3052 (N_3052,In_2939,In_736);
nand U3053 (N_3053,In_1013,In_2809);
xor U3054 (N_3054,In_2466,In_1356);
or U3055 (N_3055,In_229,In_165);
or U3056 (N_3056,In_1770,In_2584);
xnor U3057 (N_3057,In_1617,In_2736);
nand U3058 (N_3058,In_254,In_953);
nor U3059 (N_3059,In_2410,In_1653);
and U3060 (N_3060,In_1429,In_2871);
and U3061 (N_3061,In_2906,In_1114);
nor U3062 (N_3062,In_1426,In_1528);
nand U3063 (N_3063,In_2008,In_206);
or U3064 (N_3064,In_2491,In_1950);
or U3065 (N_3065,In_2013,In_767);
nand U3066 (N_3066,In_317,In_464);
and U3067 (N_3067,In_1753,In_401);
xor U3068 (N_3068,In_1181,In_134);
xnor U3069 (N_3069,In_2854,In_2722);
nand U3070 (N_3070,In_2374,In_754);
nand U3071 (N_3071,In_2744,In_1499);
or U3072 (N_3072,In_241,In_1093);
or U3073 (N_3073,In_1069,In_1116);
nand U3074 (N_3074,In_2006,In_149);
and U3075 (N_3075,In_2229,In_1099);
nor U3076 (N_3076,In_1340,In_1101);
nor U3077 (N_3077,In_1607,In_486);
xor U3078 (N_3078,In_641,In_937);
nor U3079 (N_3079,In_2030,In_1049);
xor U3080 (N_3080,In_1819,In_1470);
xnor U3081 (N_3081,In_25,In_765);
nand U3082 (N_3082,In_2124,In_1669);
nand U3083 (N_3083,In_2484,In_1247);
nor U3084 (N_3084,In_2049,In_2164);
nand U3085 (N_3085,In_2470,In_2619);
nand U3086 (N_3086,In_915,In_2116);
and U3087 (N_3087,In_2364,In_838);
or U3088 (N_3088,In_771,In_1098);
and U3089 (N_3089,In_2792,In_325);
and U3090 (N_3090,In_38,In_2020);
nor U3091 (N_3091,In_2174,In_1885);
nor U3092 (N_3092,In_242,In_1071);
or U3093 (N_3093,In_1025,In_2990);
and U3094 (N_3094,In_1140,In_316);
or U3095 (N_3095,In_1150,In_2487);
xor U3096 (N_3096,In_1865,In_442);
or U3097 (N_3097,In_2445,In_1755);
nor U3098 (N_3098,In_54,In_2497);
nand U3099 (N_3099,In_2656,In_537);
or U3100 (N_3100,In_2499,In_113);
or U3101 (N_3101,In_513,In_2668);
nor U3102 (N_3102,In_790,In_309);
xnor U3103 (N_3103,In_2635,In_2445);
or U3104 (N_3104,In_1092,In_2772);
xnor U3105 (N_3105,In_2317,In_1429);
nor U3106 (N_3106,In_2452,In_2547);
xnor U3107 (N_3107,In_366,In_2567);
xor U3108 (N_3108,In_1772,In_237);
and U3109 (N_3109,In_2294,In_2349);
xor U3110 (N_3110,In_2790,In_1124);
nand U3111 (N_3111,In_1576,In_2205);
and U3112 (N_3112,In_1345,In_1933);
nand U3113 (N_3113,In_203,In_803);
or U3114 (N_3114,In_2207,In_1874);
or U3115 (N_3115,In_2664,In_1685);
xnor U3116 (N_3116,In_182,In_213);
nor U3117 (N_3117,In_518,In_457);
and U3118 (N_3118,In_1100,In_2462);
nand U3119 (N_3119,In_2846,In_1868);
xor U3120 (N_3120,In_1469,In_151);
nor U3121 (N_3121,In_986,In_1017);
xnor U3122 (N_3122,In_2825,In_1365);
xnor U3123 (N_3123,In_231,In_2091);
and U3124 (N_3124,In_953,In_2594);
nor U3125 (N_3125,In_256,In_864);
xor U3126 (N_3126,In_50,In_2633);
nand U3127 (N_3127,In_1176,In_998);
nor U3128 (N_3128,In_1259,In_1401);
nor U3129 (N_3129,In_1291,In_845);
or U3130 (N_3130,In_367,In_917);
nor U3131 (N_3131,In_694,In_1891);
nor U3132 (N_3132,In_763,In_1723);
or U3133 (N_3133,In_1688,In_364);
xnor U3134 (N_3134,In_2010,In_2091);
xnor U3135 (N_3135,In_1107,In_2075);
and U3136 (N_3136,In_1460,In_2519);
or U3137 (N_3137,In_899,In_832);
nand U3138 (N_3138,In_963,In_1726);
and U3139 (N_3139,In_423,In_1623);
and U3140 (N_3140,In_2329,In_809);
xor U3141 (N_3141,In_1469,In_858);
nand U3142 (N_3142,In_2496,In_852);
or U3143 (N_3143,In_105,In_2903);
nand U3144 (N_3144,In_1133,In_2124);
or U3145 (N_3145,In_1528,In_43);
nor U3146 (N_3146,In_2580,In_2380);
xor U3147 (N_3147,In_906,In_2277);
nand U3148 (N_3148,In_2091,In_1710);
and U3149 (N_3149,In_2060,In_123);
nor U3150 (N_3150,In_1208,In_139);
nor U3151 (N_3151,In_1536,In_1213);
nor U3152 (N_3152,In_2483,In_1773);
and U3153 (N_3153,In_777,In_137);
xor U3154 (N_3154,In_2880,In_1391);
or U3155 (N_3155,In_820,In_490);
nor U3156 (N_3156,In_426,In_855);
nor U3157 (N_3157,In_103,In_1122);
xor U3158 (N_3158,In_186,In_1209);
or U3159 (N_3159,In_760,In_934);
nand U3160 (N_3160,In_2406,In_1334);
and U3161 (N_3161,In_1714,In_634);
and U3162 (N_3162,In_479,In_1623);
and U3163 (N_3163,In_2478,In_340);
and U3164 (N_3164,In_1187,In_909);
nand U3165 (N_3165,In_1839,In_1292);
and U3166 (N_3166,In_1877,In_85);
nand U3167 (N_3167,In_1317,In_633);
or U3168 (N_3168,In_1117,In_87);
nand U3169 (N_3169,In_2673,In_2460);
nor U3170 (N_3170,In_1741,In_2931);
nand U3171 (N_3171,In_100,In_2914);
and U3172 (N_3172,In_839,In_2268);
and U3173 (N_3173,In_2857,In_1827);
or U3174 (N_3174,In_2475,In_1085);
xnor U3175 (N_3175,In_121,In_2791);
or U3176 (N_3176,In_452,In_2041);
or U3177 (N_3177,In_1328,In_2182);
xor U3178 (N_3178,In_2123,In_2154);
nor U3179 (N_3179,In_2128,In_365);
and U3180 (N_3180,In_1680,In_2531);
nor U3181 (N_3181,In_2727,In_71);
or U3182 (N_3182,In_2408,In_1241);
or U3183 (N_3183,In_783,In_1664);
nor U3184 (N_3184,In_526,In_710);
nand U3185 (N_3185,In_2111,In_2137);
nand U3186 (N_3186,In_386,In_2255);
or U3187 (N_3187,In_41,In_2792);
nor U3188 (N_3188,In_1624,In_23);
nand U3189 (N_3189,In_1265,In_2183);
nor U3190 (N_3190,In_1284,In_1282);
or U3191 (N_3191,In_1656,In_2870);
nor U3192 (N_3192,In_2528,In_1233);
nor U3193 (N_3193,In_383,In_1237);
xnor U3194 (N_3194,In_2600,In_731);
xnor U3195 (N_3195,In_2600,In_1997);
and U3196 (N_3196,In_958,In_698);
or U3197 (N_3197,In_2128,In_1025);
xnor U3198 (N_3198,In_2414,In_1750);
and U3199 (N_3199,In_372,In_338);
nand U3200 (N_3200,In_1853,In_2662);
and U3201 (N_3201,In_1968,In_1017);
xor U3202 (N_3202,In_1700,In_977);
or U3203 (N_3203,In_1732,In_247);
xor U3204 (N_3204,In_1058,In_1012);
and U3205 (N_3205,In_1784,In_2028);
xor U3206 (N_3206,In_2119,In_2694);
nand U3207 (N_3207,In_2237,In_886);
or U3208 (N_3208,In_667,In_284);
nor U3209 (N_3209,In_2045,In_2537);
and U3210 (N_3210,In_1549,In_2472);
nand U3211 (N_3211,In_2403,In_2018);
and U3212 (N_3212,In_2911,In_2651);
nand U3213 (N_3213,In_172,In_1221);
xnor U3214 (N_3214,In_2871,In_834);
or U3215 (N_3215,In_758,In_208);
and U3216 (N_3216,In_1845,In_2302);
nand U3217 (N_3217,In_2637,In_2934);
nor U3218 (N_3218,In_2256,In_1127);
or U3219 (N_3219,In_2968,In_85);
and U3220 (N_3220,In_62,In_1807);
and U3221 (N_3221,In_1166,In_2486);
nand U3222 (N_3222,In_138,In_1429);
nor U3223 (N_3223,In_2465,In_2375);
xnor U3224 (N_3224,In_1531,In_2175);
nor U3225 (N_3225,In_2231,In_989);
nor U3226 (N_3226,In_755,In_503);
xor U3227 (N_3227,In_2298,In_945);
or U3228 (N_3228,In_2092,In_2488);
nand U3229 (N_3229,In_1427,In_1566);
and U3230 (N_3230,In_1528,In_1392);
and U3231 (N_3231,In_587,In_1238);
and U3232 (N_3232,In_1140,In_997);
and U3233 (N_3233,In_1314,In_2665);
xnor U3234 (N_3234,In_2482,In_1740);
nand U3235 (N_3235,In_2779,In_1849);
nor U3236 (N_3236,In_2722,In_1428);
nand U3237 (N_3237,In_213,In_653);
or U3238 (N_3238,In_1991,In_1444);
nor U3239 (N_3239,In_2553,In_2622);
xor U3240 (N_3240,In_2218,In_1080);
nor U3241 (N_3241,In_1400,In_2711);
and U3242 (N_3242,In_786,In_495);
and U3243 (N_3243,In_2341,In_1857);
xnor U3244 (N_3244,In_2823,In_2506);
and U3245 (N_3245,In_560,In_2097);
nor U3246 (N_3246,In_2172,In_2496);
or U3247 (N_3247,In_61,In_1149);
xor U3248 (N_3248,In_1444,In_2067);
or U3249 (N_3249,In_672,In_1038);
and U3250 (N_3250,In_309,In_2290);
or U3251 (N_3251,In_2607,In_2099);
or U3252 (N_3252,In_2364,In_1172);
nor U3253 (N_3253,In_779,In_307);
nor U3254 (N_3254,In_2131,In_2590);
xnor U3255 (N_3255,In_2679,In_982);
or U3256 (N_3256,In_2458,In_731);
and U3257 (N_3257,In_2435,In_1300);
nor U3258 (N_3258,In_1127,In_2136);
nor U3259 (N_3259,In_2080,In_1500);
or U3260 (N_3260,In_1153,In_1590);
or U3261 (N_3261,In_568,In_1082);
xor U3262 (N_3262,In_1726,In_891);
xor U3263 (N_3263,In_2432,In_1144);
nand U3264 (N_3264,In_521,In_2108);
xnor U3265 (N_3265,In_2289,In_88);
xnor U3266 (N_3266,In_742,In_441);
nor U3267 (N_3267,In_2649,In_2365);
nand U3268 (N_3268,In_542,In_2001);
and U3269 (N_3269,In_1617,In_2115);
or U3270 (N_3270,In_1086,In_2113);
and U3271 (N_3271,In_2147,In_960);
xor U3272 (N_3272,In_2943,In_409);
xor U3273 (N_3273,In_2753,In_1930);
and U3274 (N_3274,In_245,In_2995);
xor U3275 (N_3275,In_743,In_962);
xnor U3276 (N_3276,In_111,In_1190);
and U3277 (N_3277,In_1994,In_2347);
nand U3278 (N_3278,In_2987,In_2052);
xnor U3279 (N_3279,In_169,In_2825);
nor U3280 (N_3280,In_1069,In_989);
nor U3281 (N_3281,In_2390,In_2358);
or U3282 (N_3282,In_966,In_633);
or U3283 (N_3283,In_1345,In_1755);
or U3284 (N_3284,In_2742,In_2169);
or U3285 (N_3285,In_662,In_1253);
and U3286 (N_3286,In_1960,In_233);
and U3287 (N_3287,In_1279,In_1801);
nor U3288 (N_3288,In_2919,In_398);
or U3289 (N_3289,In_2189,In_239);
nor U3290 (N_3290,In_2519,In_136);
nor U3291 (N_3291,In_641,In_2485);
nor U3292 (N_3292,In_1710,In_1720);
and U3293 (N_3293,In_450,In_2549);
and U3294 (N_3294,In_531,In_1841);
xnor U3295 (N_3295,In_1394,In_1666);
nor U3296 (N_3296,In_494,In_1352);
or U3297 (N_3297,In_518,In_355);
nand U3298 (N_3298,In_1412,In_145);
or U3299 (N_3299,In_2604,In_1671);
xnor U3300 (N_3300,In_741,In_1029);
xor U3301 (N_3301,In_915,In_2983);
or U3302 (N_3302,In_1048,In_2010);
nand U3303 (N_3303,In_227,In_2887);
nor U3304 (N_3304,In_1231,In_1853);
nand U3305 (N_3305,In_1606,In_672);
or U3306 (N_3306,In_1680,In_1970);
and U3307 (N_3307,In_376,In_1991);
xnor U3308 (N_3308,In_2816,In_708);
xnor U3309 (N_3309,In_692,In_1053);
nor U3310 (N_3310,In_1571,In_2345);
nor U3311 (N_3311,In_2243,In_2724);
or U3312 (N_3312,In_1825,In_2988);
or U3313 (N_3313,In_1296,In_598);
and U3314 (N_3314,In_1003,In_285);
and U3315 (N_3315,In_2108,In_136);
or U3316 (N_3316,In_2442,In_383);
nand U3317 (N_3317,In_2961,In_1544);
nor U3318 (N_3318,In_2936,In_1738);
nor U3319 (N_3319,In_2301,In_2617);
nor U3320 (N_3320,In_2484,In_637);
xnor U3321 (N_3321,In_2863,In_2357);
or U3322 (N_3322,In_2528,In_2453);
xor U3323 (N_3323,In_2422,In_1627);
or U3324 (N_3324,In_1674,In_2506);
or U3325 (N_3325,In_1366,In_112);
nand U3326 (N_3326,In_303,In_1867);
or U3327 (N_3327,In_1086,In_2809);
and U3328 (N_3328,In_2139,In_706);
nor U3329 (N_3329,In_2010,In_1055);
nand U3330 (N_3330,In_984,In_1760);
or U3331 (N_3331,In_1464,In_960);
xnor U3332 (N_3332,In_501,In_330);
xnor U3333 (N_3333,In_441,In_1352);
nand U3334 (N_3334,In_1883,In_561);
or U3335 (N_3335,In_2444,In_44);
nand U3336 (N_3336,In_380,In_812);
nor U3337 (N_3337,In_240,In_634);
xor U3338 (N_3338,In_1709,In_2976);
or U3339 (N_3339,In_1627,In_306);
and U3340 (N_3340,In_2726,In_1387);
nand U3341 (N_3341,In_1522,In_1008);
xnor U3342 (N_3342,In_2437,In_2249);
nor U3343 (N_3343,In_2333,In_1700);
nand U3344 (N_3344,In_2902,In_1258);
nor U3345 (N_3345,In_228,In_64);
or U3346 (N_3346,In_2182,In_240);
and U3347 (N_3347,In_391,In_2223);
or U3348 (N_3348,In_2969,In_2341);
xor U3349 (N_3349,In_2154,In_2013);
and U3350 (N_3350,In_186,In_2813);
nand U3351 (N_3351,In_533,In_2796);
nand U3352 (N_3352,In_2659,In_2099);
and U3353 (N_3353,In_250,In_2124);
and U3354 (N_3354,In_1036,In_1174);
xor U3355 (N_3355,In_1959,In_2756);
nor U3356 (N_3356,In_2717,In_1224);
xor U3357 (N_3357,In_271,In_174);
and U3358 (N_3358,In_842,In_1058);
nand U3359 (N_3359,In_2112,In_1649);
nand U3360 (N_3360,In_2746,In_2480);
nand U3361 (N_3361,In_546,In_350);
nand U3362 (N_3362,In_1027,In_2675);
xor U3363 (N_3363,In_2935,In_1247);
and U3364 (N_3364,In_2699,In_2871);
nor U3365 (N_3365,In_260,In_1571);
nand U3366 (N_3366,In_1004,In_1917);
or U3367 (N_3367,In_1018,In_864);
xor U3368 (N_3368,In_951,In_1506);
xnor U3369 (N_3369,In_2713,In_1526);
or U3370 (N_3370,In_547,In_2286);
and U3371 (N_3371,In_1387,In_835);
nor U3372 (N_3372,In_86,In_2820);
xnor U3373 (N_3373,In_1554,In_1075);
or U3374 (N_3374,In_2537,In_1006);
nor U3375 (N_3375,In_1611,In_1658);
or U3376 (N_3376,In_457,In_2416);
or U3377 (N_3377,In_1342,In_2309);
xnor U3378 (N_3378,In_2152,In_212);
xnor U3379 (N_3379,In_1525,In_2636);
or U3380 (N_3380,In_2930,In_875);
nor U3381 (N_3381,In_2656,In_1471);
and U3382 (N_3382,In_1998,In_980);
nor U3383 (N_3383,In_2967,In_1865);
nand U3384 (N_3384,In_2866,In_1868);
or U3385 (N_3385,In_666,In_316);
or U3386 (N_3386,In_1115,In_1218);
and U3387 (N_3387,In_1685,In_2074);
and U3388 (N_3388,In_312,In_1016);
and U3389 (N_3389,In_883,In_2309);
and U3390 (N_3390,In_834,In_668);
or U3391 (N_3391,In_2149,In_1329);
nor U3392 (N_3392,In_2340,In_197);
and U3393 (N_3393,In_2466,In_1603);
nand U3394 (N_3394,In_946,In_328);
xnor U3395 (N_3395,In_1781,In_660);
nor U3396 (N_3396,In_1759,In_2898);
or U3397 (N_3397,In_696,In_2681);
or U3398 (N_3398,In_1012,In_1218);
and U3399 (N_3399,In_1101,In_2916);
and U3400 (N_3400,In_2330,In_2181);
nand U3401 (N_3401,In_2225,In_2865);
and U3402 (N_3402,In_70,In_2191);
nand U3403 (N_3403,In_2655,In_1279);
xnor U3404 (N_3404,In_1261,In_1484);
and U3405 (N_3405,In_2164,In_1934);
and U3406 (N_3406,In_2350,In_133);
or U3407 (N_3407,In_2582,In_314);
xor U3408 (N_3408,In_749,In_1318);
nor U3409 (N_3409,In_2883,In_552);
and U3410 (N_3410,In_891,In_591);
nand U3411 (N_3411,In_1900,In_1446);
or U3412 (N_3412,In_1368,In_2187);
or U3413 (N_3413,In_868,In_2974);
and U3414 (N_3414,In_859,In_1950);
nand U3415 (N_3415,In_668,In_621);
and U3416 (N_3416,In_1885,In_1611);
xnor U3417 (N_3417,In_350,In_960);
or U3418 (N_3418,In_2949,In_2186);
and U3419 (N_3419,In_2228,In_2094);
and U3420 (N_3420,In_721,In_1157);
nand U3421 (N_3421,In_1540,In_1204);
nor U3422 (N_3422,In_1833,In_1951);
nor U3423 (N_3423,In_2234,In_492);
or U3424 (N_3424,In_364,In_323);
xor U3425 (N_3425,In_697,In_1088);
and U3426 (N_3426,In_2075,In_1257);
nand U3427 (N_3427,In_1024,In_1201);
and U3428 (N_3428,In_905,In_651);
nor U3429 (N_3429,In_2592,In_825);
nand U3430 (N_3430,In_71,In_205);
xor U3431 (N_3431,In_581,In_109);
and U3432 (N_3432,In_1769,In_1997);
and U3433 (N_3433,In_2982,In_736);
or U3434 (N_3434,In_1023,In_1632);
and U3435 (N_3435,In_2243,In_902);
nand U3436 (N_3436,In_1010,In_2958);
and U3437 (N_3437,In_207,In_209);
xnor U3438 (N_3438,In_1327,In_337);
nand U3439 (N_3439,In_460,In_1084);
nand U3440 (N_3440,In_617,In_2189);
nand U3441 (N_3441,In_115,In_2781);
or U3442 (N_3442,In_592,In_1835);
xnor U3443 (N_3443,In_2978,In_2086);
nor U3444 (N_3444,In_2748,In_150);
or U3445 (N_3445,In_1568,In_1765);
or U3446 (N_3446,In_2484,In_881);
or U3447 (N_3447,In_1685,In_2496);
nor U3448 (N_3448,In_2352,In_2300);
xor U3449 (N_3449,In_2290,In_1189);
and U3450 (N_3450,In_1829,In_1661);
xnor U3451 (N_3451,In_1763,In_2294);
xnor U3452 (N_3452,In_1996,In_523);
nand U3453 (N_3453,In_2662,In_860);
or U3454 (N_3454,In_382,In_249);
nor U3455 (N_3455,In_1571,In_544);
nand U3456 (N_3456,In_2550,In_242);
xnor U3457 (N_3457,In_647,In_1038);
xnor U3458 (N_3458,In_792,In_1890);
and U3459 (N_3459,In_2137,In_1642);
nand U3460 (N_3460,In_2314,In_2259);
or U3461 (N_3461,In_276,In_321);
nor U3462 (N_3462,In_1058,In_2247);
and U3463 (N_3463,In_1177,In_2557);
nor U3464 (N_3464,In_1932,In_608);
xnor U3465 (N_3465,In_2823,In_1887);
and U3466 (N_3466,In_2749,In_1980);
or U3467 (N_3467,In_1193,In_98);
xnor U3468 (N_3468,In_2076,In_465);
and U3469 (N_3469,In_2580,In_152);
or U3470 (N_3470,In_2371,In_2236);
or U3471 (N_3471,In_2063,In_2073);
nand U3472 (N_3472,In_2437,In_2673);
or U3473 (N_3473,In_2650,In_2714);
nand U3474 (N_3474,In_1930,In_874);
or U3475 (N_3475,In_2480,In_2993);
and U3476 (N_3476,In_1152,In_1541);
nand U3477 (N_3477,In_465,In_881);
or U3478 (N_3478,In_2313,In_2464);
nor U3479 (N_3479,In_922,In_440);
nand U3480 (N_3480,In_1483,In_2756);
nand U3481 (N_3481,In_2739,In_2184);
nand U3482 (N_3482,In_632,In_2391);
or U3483 (N_3483,In_286,In_2100);
xnor U3484 (N_3484,In_71,In_762);
and U3485 (N_3485,In_209,In_863);
xnor U3486 (N_3486,In_2267,In_1414);
nand U3487 (N_3487,In_1448,In_1862);
nand U3488 (N_3488,In_198,In_2653);
and U3489 (N_3489,In_2294,In_2118);
nand U3490 (N_3490,In_1130,In_1959);
nor U3491 (N_3491,In_160,In_1410);
or U3492 (N_3492,In_964,In_2110);
nor U3493 (N_3493,In_1844,In_604);
or U3494 (N_3494,In_2404,In_229);
nor U3495 (N_3495,In_867,In_2093);
nand U3496 (N_3496,In_1109,In_2876);
or U3497 (N_3497,In_17,In_319);
nor U3498 (N_3498,In_2244,In_1186);
xnor U3499 (N_3499,In_2808,In_1124);
or U3500 (N_3500,In_1941,In_1301);
nor U3501 (N_3501,In_2218,In_105);
nand U3502 (N_3502,In_1264,In_360);
xnor U3503 (N_3503,In_2946,In_1476);
or U3504 (N_3504,In_1259,In_517);
or U3505 (N_3505,In_449,In_2648);
xnor U3506 (N_3506,In_801,In_1959);
and U3507 (N_3507,In_2442,In_797);
xnor U3508 (N_3508,In_2274,In_1225);
and U3509 (N_3509,In_506,In_2344);
or U3510 (N_3510,In_490,In_2639);
or U3511 (N_3511,In_100,In_362);
nand U3512 (N_3512,In_1825,In_2224);
or U3513 (N_3513,In_2128,In_1048);
nor U3514 (N_3514,In_2158,In_2455);
nand U3515 (N_3515,In_2252,In_299);
and U3516 (N_3516,In_2574,In_2717);
nand U3517 (N_3517,In_1937,In_430);
nor U3518 (N_3518,In_2628,In_2414);
xor U3519 (N_3519,In_1452,In_478);
and U3520 (N_3520,In_882,In_1982);
and U3521 (N_3521,In_1831,In_66);
nand U3522 (N_3522,In_1871,In_942);
nand U3523 (N_3523,In_2845,In_695);
nand U3524 (N_3524,In_1548,In_644);
or U3525 (N_3525,In_1048,In_1065);
nand U3526 (N_3526,In_464,In_2486);
and U3527 (N_3527,In_1487,In_2023);
nand U3528 (N_3528,In_153,In_1700);
xor U3529 (N_3529,In_2106,In_966);
xnor U3530 (N_3530,In_1101,In_314);
or U3531 (N_3531,In_720,In_604);
nand U3532 (N_3532,In_2135,In_590);
nor U3533 (N_3533,In_561,In_427);
xor U3534 (N_3534,In_2086,In_2680);
nor U3535 (N_3535,In_983,In_2097);
or U3536 (N_3536,In_2816,In_1003);
or U3537 (N_3537,In_423,In_2677);
or U3538 (N_3538,In_1298,In_146);
xnor U3539 (N_3539,In_156,In_1498);
and U3540 (N_3540,In_2205,In_160);
nor U3541 (N_3541,In_2242,In_732);
nand U3542 (N_3542,In_264,In_1066);
nor U3543 (N_3543,In_2016,In_1207);
nand U3544 (N_3544,In_606,In_1654);
or U3545 (N_3545,In_1899,In_2168);
nand U3546 (N_3546,In_187,In_2185);
and U3547 (N_3547,In_2055,In_553);
or U3548 (N_3548,In_237,In_1955);
or U3549 (N_3549,In_56,In_1228);
and U3550 (N_3550,In_2861,In_837);
nor U3551 (N_3551,In_2473,In_1203);
xnor U3552 (N_3552,In_203,In_1502);
xor U3553 (N_3553,In_2858,In_1930);
xor U3554 (N_3554,In_2234,In_2230);
or U3555 (N_3555,In_877,In_2773);
xnor U3556 (N_3556,In_991,In_1900);
nand U3557 (N_3557,In_477,In_317);
nor U3558 (N_3558,In_1918,In_1892);
xnor U3559 (N_3559,In_2445,In_2420);
nor U3560 (N_3560,In_385,In_2074);
xor U3561 (N_3561,In_299,In_2482);
xnor U3562 (N_3562,In_1612,In_2738);
and U3563 (N_3563,In_1520,In_1315);
xor U3564 (N_3564,In_47,In_972);
nand U3565 (N_3565,In_103,In_876);
nand U3566 (N_3566,In_1367,In_774);
and U3567 (N_3567,In_706,In_2307);
nor U3568 (N_3568,In_2018,In_1324);
nand U3569 (N_3569,In_2926,In_2578);
xor U3570 (N_3570,In_1670,In_1889);
nor U3571 (N_3571,In_987,In_1967);
xnor U3572 (N_3572,In_1952,In_440);
and U3573 (N_3573,In_393,In_1275);
or U3574 (N_3574,In_340,In_470);
nor U3575 (N_3575,In_2642,In_1596);
or U3576 (N_3576,In_611,In_1465);
or U3577 (N_3577,In_846,In_1499);
xor U3578 (N_3578,In_2902,In_1559);
nand U3579 (N_3579,In_2828,In_2322);
xnor U3580 (N_3580,In_2065,In_2928);
xnor U3581 (N_3581,In_921,In_931);
nor U3582 (N_3582,In_2012,In_601);
and U3583 (N_3583,In_2186,In_2062);
or U3584 (N_3584,In_632,In_2279);
nand U3585 (N_3585,In_152,In_1876);
nand U3586 (N_3586,In_2482,In_1496);
xor U3587 (N_3587,In_1522,In_568);
or U3588 (N_3588,In_21,In_538);
or U3589 (N_3589,In_47,In_2120);
and U3590 (N_3590,In_2528,In_181);
nand U3591 (N_3591,In_1575,In_1025);
xor U3592 (N_3592,In_1284,In_624);
or U3593 (N_3593,In_2995,In_909);
nand U3594 (N_3594,In_1120,In_575);
or U3595 (N_3595,In_2745,In_1541);
nand U3596 (N_3596,In_623,In_611);
nor U3597 (N_3597,In_882,In_1743);
and U3598 (N_3598,In_11,In_1584);
nand U3599 (N_3599,In_2962,In_2366);
nand U3600 (N_3600,In_183,In_700);
or U3601 (N_3601,In_779,In_121);
nand U3602 (N_3602,In_2968,In_302);
nor U3603 (N_3603,In_2890,In_1061);
nand U3604 (N_3604,In_1593,In_1265);
nand U3605 (N_3605,In_1950,In_37);
xor U3606 (N_3606,In_929,In_2621);
and U3607 (N_3607,In_910,In_357);
nor U3608 (N_3608,In_663,In_1344);
nor U3609 (N_3609,In_560,In_2982);
and U3610 (N_3610,In_1391,In_1576);
nor U3611 (N_3611,In_94,In_998);
nand U3612 (N_3612,In_1867,In_1512);
nand U3613 (N_3613,In_2018,In_2910);
or U3614 (N_3614,In_68,In_725);
xor U3615 (N_3615,In_1923,In_2966);
and U3616 (N_3616,In_656,In_402);
or U3617 (N_3617,In_1154,In_1812);
xnor U3618 (N_3618,In_528,In_2719);
xnor U3619 (N_3619,In_2032,In_374);
nor U3620 (N_3620,In_1138,In_1581);
nor U3621 (N_3621,In_940,In_662);
xnor U3622 (N_3622,In_1624,In_2488);
or U3623 (N_3623,In_716,In_721);
nand U3624 (N_3624,In_770,In_1411);
nor U3625 (N_3625,In_2404,In_1669);
nand U3626 (N_3626,In_344,In_1236);
and U3627 (N_3627,In_2977,In_1277);
or U3628 (N_3628,In_2914,In_584);
or U3629 (N_3629,In_2999,In_2323);
nor U3630 (N_3630,In_1264,In_2023);
nand U3631 (N_3631,In_2689,In_2892);
nand U3632 (N_3632,In_1889,In_1007);
nand U3633 (N_3633,In_46,In_1347);
and U3634 (N_3634,In_1648,In_2839);
xnor U3635 (N_3635,In_2083,In_2391);
nand U3636 (N_3636,In_106,In_2488);
nand U3637 (N_3637,In_2277,In_2001);
and U3638 (N_3638,In_2643,In_1313);
xor U3639 (N_3639,In_1791,In_1042);
xnor U3640 (N_3640,In_2669,In_2155);
and U3641 (N_3641,In_1943,In_2628);
nand U3642 (N_3642,In_1927,In_492);
nand U3643 (N_3643,In_984,In_2762);
or U3644 (N_3644,In_671,In_1277);
xnor U3645 (N_3645,In_189,In_836);
nor U3646 (N_3646,In_1812,In_473);
and U3647 (N_3647,In_2126,In_704);
nor U3648 (N_3648,In_253,In_2126);
or U3649 (N_3649,In_2150,In_536);
xor U3650 (N_3650,In_832,In_319);
nor U3651 (N_3651,In_2582,In_2192);
and U3652 (N_3652,In_2444,In_1189);
nand U3653 (N_3653,In_1788,In_1687);
nand U3654 (N_3654,In_2600,In_1384);
and U3655 (N_3655,In_164,In_195);
nand U3656 (N_3656,In_2669,In_140);
nor U3657 (N_3657,In_1503,In_2553);
nor U3658 (N_3658,In_728,In_861);
xnor U3659 (N_3659,In_236,In_2365);
nor U3660 (N_3660,In_3,In_1555);
nor U3661 (N_3661,In_2330,In_1883);
or U3662 (N_3662,In_762,In_2699);
xnor U3663 (N_3663,In_1794,In_76);
and U3664 (N_3664,In_2085,In_1103);
xnor U3665 (N_3665,In_1322,In_1359);
xnor U3666 (N_3666,In_1404,In_1907);
or U3667 (N_3667,In_2700,In_1943);
nand U3668 (N_3668,In_1014,In_1605);
nor U3669 (N_3669,In_2873,In_387);
nand U3670 (N_3670,In_1054,In_2644);
nor U3671 (N_3671,In_1065,In_960);
nand U3672 (N_3672,In_2051,In_2792);
or U3673 (N_3673,In_1669,In_1415);
or U3674 (N_3674,In_176,In_1328);
nor U3675 (N_3675,In_2450,In_2483);
or U3676 (N_3676,In_2166,In_683);
nor U3677 (N_3677,In_2981,In_1464);
and U3678 (N_3678,In_2644,In_2197);
and U3679 (N_3679,In_412,In_885);
and U3680 (N_3680,In_2781,In_438);
xnor U3681 (N_3681,In_481,In_234);
and U3682 (N_3682,In_1447,In_2259);
and U3683 (N_3683,In_2958,In_2990);
nand U3684 (N_3684,In_1609,In_2468);
nor U3685 (N_3685,In_1346,In_1410);
nor U3686 (N_3686,In_2798,In_1419);
and U3687 (N_3687,In_435,In_2999);
xor U3688 (N_3688,In_2625,In_1180);
nand U3689 (N_3689,In_1000,In_1240);
nand U3690 (N_3690,In_415,In_250);
nor U3691 (N_3691,In_372,In_231);
and U3692 (N_3692,In_1773,In_627);
nand U3693 (N_3693,In_1827,In_1880);
nand U3694 (N_3694,In_535,In_2367);
or U3695 (N_3695,In_2228,In_2490);
and U3696 (N_3696,In_955,In_2158);
and U3697 (N_3697,In_1139,In_2520);
nor U3698 (N_3698,In_223,In_2695);
xor U3699 (N_3699,In_1068,In_2132);
and U3700 (N_3700,In_2180,In_1328);
nor U3701 (N_3701,In_853,In_2151);
or U3702 (N_3702,In_770,In_572);
nor U3703 (N_3703,In_1288,In_2539);
or U3704 (N_3704,In_2027,In_1271);
or U3705 (N_3705,In_2571,In_1053);
nand U3706 (N_3706,In_2592,In_947);
nand U3707 (N_3707,In_2271,In_1822);
and U3708 (N_3708,In_2398,In_2881);
nor U3709 (N_3709,In_2120,In_1593);
nand U3710 (N_3710,In_1757,In_358);
xor U3711 (N_3711,In_1966,In_2271);
nor U3712 (N_3712,In_2230,In_435);
nand U3713 (N_3713,In_2586,In_704);
nor U3714 (N_3714,In_2894,In_2668);
or U3715 (N_3715,In_420,In_2211);
nor U3716 (N_3716,In_2682,In_1515);
nand U3717 (N_3717,In_1399,In_2556);
nor U3718 (N_3718,In_869,In_2324);
nand U3719 (N_3719,In_2130,In_2897);
or U3720 (N_3720,In_1347,In_1918);
xor U3721 (N_3721,In_1781,In_2621);
and U3722 (N_3722,In_2939,In_1773);
or U3723 (N_3723,In_1674,In_1173);
and U3724 (N_3724,In_1555,In_736);
xor U3725 (N_3725,In_1533,In_2236);
or U3726 (N_3726,In_658,In_55);
or U3727 (N_3727,In_2336,In_256);
or U3728 (N_3728,In_2610,In_1378);
xnor U3729 (N_3729,In_1327,In_174);
xnor U3730 (N_3730,In_2468,In_1428);
or U3731 (N_3731,In_53,In_849);
and U3732 (N_3732,In_1791,In_1767);
or U3733 (N_3733,In_973,In_1864);
and U3734 (N_3734,In_1541,In_2740);
xnor U3735 (N_3735,In_2776,In_356);
nand U3736 (N_3736,In_1976,In_1615);
or U3737 (N_3737,In_1320,In_2320);
xnor U3738 (N_3738,In_1208,In_179);
or U3739 (N_3739,In_722,In_458);
xnor U3740 (N_3740,In_21,In_574);
xor U3741 (N_3741,In_2506,In_2068);
xor U3742 (N_3742,In_2992,In_1369);
nand U3743 (N_3743,In_371,In_31);
xor U3744 (N_3744,In_2435,In_542);
xnor U3745 (N_3745,In_2292,In_1300);
or U3746 (N_3746,In_207,In_1428);
nand U3747 (N_3747,In_699,In_1474);
or U3748 (N_3748,In_2081,In_826);
xor U3749 (N_3749,In_1864,In_1284);
nand U3750 (N_3750,In_1395,In_2145);
or U3751 (N_3751,In_2638,In_2443);
nor U3752 (N_3752,In_93,In_55);
xnor U3753 (N_3753,In_1469,In_987);
nand U3754 (N_3754,In_20,In_1600);
and U3755 (N_3755,In_1783,In_2787);
nand U3756 (N_3756,In_285,In_381);
and U3757 (N_3757,In_1770,In_2090);
and U3758 (N_3758,In_158,In_1051);
and U3759 (N_3759,In_2613,In_2216);
nor U3760 (N_3760,In_1241,In_2960);
nand U3761 (N_3761,In_1001,In_2685);
or U3762 (N_3762,In_2513,In_2733);
xnor U3763 (N_3763,In_2720,In_1538);
nand U3764 (N_3764,In_2238,In_1160);
and U3765 (N_3765,In_1011,In_1515);
and U3766 (N_3766,In_1627,In_2893);
or U3767 (N_3767,In_2155,In_2909);
nor U3768 (N_3768,In_231,In_1343);
nand U3769 (N_3769,In_806,In_1442);
or U3770 (N_3770,In_2960,In_1099);
or U3771 (N_3771,In_293,In_906);
nor U3772 (N_3772,In_1883,In_1173);
nand U3773 (N_3773,In_2408,In_2814);
nand U3774 (N_3774,In_785,In_1198);
or U3775 (N_3775,In_427,In_2989);
nor U3776 (N_3776,In_1951,In_1409);
xnor U3777 (N_3777,In_2914,In_692);
nand U3778 (N_3778,In_1343,In_2117);
nor U3779 (N_3779,In_219,In_2142);
nor U3780 (N_3780,In_90,In_808);
nor U3781 (N_3781,In_1704,In_1506);
and U3782 (N_3782,In_1245,In_800);
and U3783 (N_3783,In_2219,In_76);
and U3784 (N_3784,In_337,In_1690);
xnor U3785 (N_3785,In_774,In_2269);
nor U3786 (N_3786,In_57,In_750);
nand U3787 (N_3787,In_821,In_2663);
or U3788 (N_3788,In_2456,In_1146);
and U3789 (N_3789,In_1204,In_2199);
or U3790 (N_3790,In_1628,In_1828);
xnor U3791 (N_3791,In_2094,In_2498);
and U3792 (N_3792,In_1991,In_534);
nor U3793 (N_3793,In_1888,In_1949);
xor U3794 (N_3794,In_2260,In_249);
and U3795 (N_3795,In_2222,In_2382);
nor U3796 (N_3796,In_2663,In_1923);
nand U3797 (N_3797,In_1187,In_851);
xor U3798 (N_3798,In_1970,In_1223);
nor U3799 (N_3799,In_2884,In_459);
nand U3800 (N_3800,In_1979,In_2840);
or U3801 (N_3801,In_553,In_350);
xnor U3802 (N_3802,In_2808,In_2944);
and U3803 (N_3803,In_1529,In_2681);
nor U3804 (N_3804,In_2452,In_1445);
xor U3805 (N_3805,In_411,In_1713);
or U3806 (N_3806,In_2122,In_2394);
nor U3807 (N_3807,In_1003,In_1773);
nand U3808 (N_3808,In_1315,In_2593);
nand U3809 (N_3809,In_2003,In_1589);
or U3810 (N_3810,In_655,In_1607);
or U3811 (N_3811,In_130,In_106);
and U3812 (N_3812,In_184,In_1737);
nor U3813 (N_3813,In_465,In_1093);
nand U3814 (N_3814,In_650,In_75);
or U3815 (N_3815,In_2248,In_422);
or U3816 (N_3816,In_2112,In_876);
nand U3817 (N_3817,In_1829,In_2428);
or U3818 (N_3818,In_1876,In_1064);
nor U3819 (N_3819,In_2724,In_2397);
or U3820 (N_3820,In_2432,In_2970);
nor U3821 (N_3821,In_2929,In_148);
xnor U3822 (N_3822,In_2153,In_2585);
nor U3823 (N_3823,In_585,In_2687);
nor U3824 (N_3824,In_1228,In_880);
nor U3825 (N_3825,In_372,In_2897);
nor U3826 (N_3826,In_131,In_482);
or U3827 (N_3827,In_1530,In_1465);
or U3828 (N_3828,In_1974,In_960);
xor U3829 (N_3829,In_2171,In_905);
nand U3830 (N_3830,In_274,In_1489);
xor U3831 (N_3831,In_2636,In_2212);
or U3832 (N_3832,In_551,In_2639);
xor U3833 (N_3833,In_1301,In_710);
or U3834 (N_3834,In_2172,In_2830);
or U3835 (N_3835,In_2947,In_2611);
or U3836 (N_3836,In_818,In_780);
nand U3837 (N_3837,In_677,In_1611);
nor U3838 (N_3838,In_1080,In_2843);
or U3839 (N_3839,In_1505,In_2323);
and U3840 (N_3840,In_169,In_2324);
or U3841 (N_3841,In_2309,In_1150);
and U3842 (N_3842,In_1263,In_996);
or U3843 (N_3843,In_638,In_1398);
or U3844 (N_3844,In_2533,In_1089);
nor U3845 (N_3845,In_1990,In_1117);
nand U3846 (N_3846,In_2200,In_1836);
and U3847 (N_3847,In_699,In_169);
nand U3848 (N_3848,In_646,In_1262);
nor U3849 (N_3849,In_987,In_58);
and U3850 (N_3850,In_1762,In_2078);
or U3851 (N_3851,In_63,In_711);
or U3852 (N_3852,In_1543,In_201);
nor U3853 (N_3853,In_1414,In_2380);
or U3854 (N_3854,In_1786,In_527);
nand U3855 (N_3855,In_2027,In_2411);
xor U3856 (N_3856,In_1475,In_784);
or U3857 (N_3857,In_1404,In_1044);
or U3858 (N_3858,In_1841,In_958);
and U3859 (N_3859,In_594,In_801);
xor U3860 (N_3860,In_609,In_1984);
and U3861 (N_3861,In_577,In_2983);
xor U3862 (N_3862,In_1499,In_980);
nor U3863 (N_3863,In_2764,In_771);
nor U3864 (N_3864,In_1963,In_1682);
and U3865 (N_3865,In_1010,In_319);
nor U3866 (N_3866,In_2152,In_2498);
xor U3867 (N_3867,In_2925,In_715);
or U3868 (N_3868,In_1,In_1074);
nand U3869 (N_3869,In_246,In_280);
and U3870 (N_3870,In_1437,In_52);
xor U3871 (N_3871,In_2273,In_243);
or U3872 (N_3872,In_2766,In_1664);
and U3873 (N_3873,In_383,In_310);
nand U3874 (N_3874,In_1990,In_1754);
or U3875 (N_3875,In_1674,In_2360);
or U3876 (N_3876,In_2750,In_843);
nand U3877 (N_3877,In_1176,In_291);
xor U3878 (N_3878,In_813,In_2754);
nand U3879 (N_3879,In_1380,In_2715);
and U3880 (N_3880,In_2069,In_682);
nand U3881 (N_3881,In_2949,In_1470);
xnor U3882 (N_3882,In_1862,In_2330);
nand U3883 (N_3883,In_2844,In_606);
and U3884 (N_3884,In_902,In_2311);
or U3885 (N_3885,In_2839,In_1988);
xor U3886 (N_3886,In_1332,In_2819);
nor U3887 (N_3887,In_2147,In_865);
nand U3888 (N_3888,In_1674,In_1397);
nand U3889 (N_3889,In_1824,In_2270);
nor U3890 (N_3890,In_1919,In_766);
xor U3891 (N_3891,In_1182,In_654);
xnor U3892 (N_3892,In_2902,In_1669);
nor U3893 (N_3893,In_2915,In_945);
xor U3894 (N_3894,In_1851,In_2800);
and U3895 (N_3895,In_628,In_613);
nor U3896 (N_3896,In_606,In_1736);
nand U3897 (N_3897,In_402,In_2338);
xor U3898 (N_3898,In_1239,In_867);
xor U3899 (N_3899,In_2565,In_1668);
nor U3900 (N_3900,In_500,In_99);
nor U3901 (N_3901,In_2385,In_112);
or U3902 (N_3902,In_2546,In_683);
nor U3903 (N_3903,In_1124,In_266);
nand U3904 (N_3904,In_1226,In_1477);
or U3905 (N_3905,In_1958,In_1580);
nor U3906 (N_3906,In_1286,In_2097);
nor U3907 (N_3907,In_2988,In_1409);
nor U3908 (N_3908,In_151,In_1260);
nor U3909 (N_3909,In_1201,In_1905);
xor U3910 (N_3910,In_2340,In_1424);
nand U3911 (N_3911,In_2883,In_2730);
nor U3912 (N_3912,In_2031,In_2844);
nand U3913 (N_3913,In_1585,In_476);
nor U3914 (N_3914,In_2149,In_8);
xor U3915 (N_3915,In_2395,In_2399);
and U3916 (N_3916,In_2390,In_381);
and U3917 (N_3917,In_2058,In_951);
and U3918 (N_3918,In_630,In_1616);
xnor U3919 (N_3919,In_358,In_1558);
or U3920 (N_3920,In_2204,In_969);
xor U3921 (N_3921,In_2177,In_784);
nor U3922 (N_3922,In_2937,In_2079);
xor U3923 (N_3923,In_2301,In_2846);
nand U3924 (N_3924,In_2438,In_154);
or U3925 (N_3925,In_2914,In_2307);
and U3926 (N_3926,In_2458,In_2878);
or U3927 (N_3927,In_2927,In_1491);
xor U3928 (N_3928,In_2347,In_2932);
nor U3929 (N_3929,In_1465,In_197);
nand U3930 (N_3930,In_493,In_1081);
nor U3931 (N_3931,In_269,In_2900);
nor U3932 (N_3932,In_1682,In_1203);
nor U3933 (N_3933,In_1517,In_1792);
and U3934 (N_3934,In_534,In_1791);
nand U3935 (N_3935,In_680,In_2883);
or U3936 (N_3936,In_261,In_1357);
and U3937 (N_3937,In_1001,In_635);
xnor U3938 (N_3938,In_1837,In_2778);
or U3939 (N_3939,In_1722,In_131);
nor U3940 (N_3940,In_1387,In_322);
and U3941 (N_3941,In_2455,In_1602);
nor U3942 (N_3942,In_629,In_1627);
and U3943 (N_3943,In_795,In_350);
or U3944 (N_3944,In_522,In_1727);
and U3945 (N_3945,In_1392,In_2264);
nand U3946 (N_3946,In_2290,In_206);
or U3947 (N_3947,In_447,In_689);
xor U3948 (N_3948,In_199,In_94);
or U3949 (N_3949,In_799,In_2726);
nor U3950 (N_3950,In_704,In_1316);
nand U3951 (N_3951,In_1062,In_268);
or U3952 (N_3952,In_779,In_151);
xor U3953 (N_3953,In_73,In_1345);
xnor U3954 (N_3954,In_1766,In_2948);
xor U3955 (N_3955,In_2560,In_2451);
xnor U3956 (N_3956,In_2228,In_1118);
nand U3957 (N_3957,In_2941,In_2099);
or U3958 (N_3958,In_2823,In_883);
and U3959 (N_3959,In_1328,In_1145);
xor U3960 (N_3960,In_2969,In_100);
nand U3961 (N_3961,In_1837,In_709);
nor U3962 (N_3962,In_1405,In_735);
xnor U3963 (N_3963,In_1523,In_1193);
or U3964 (N_3964,In_790,In_771);
or U3965 (N_3965,In_2123,In_1933);
and U3966 (N_3966,In_439,In_2211);
xor U3967 (N_3967,In_390,In_536);
nand U3968 (N_3968,In_1911,In_2796);
nand U3969 (N_3969,In_2573,In_641);
nor U3970 (N_3970,In_2066,In_936);
or U3971 (N_3971,In_1829,In_2921);
nor U3972 (N_3972,In_2933,In_174);
xor U3973 (N_3973,In_2689,In_2472);
and U3974 (N_3974,In_477,In_4);
nand U3975 (N_3975,In_2611,In_1741);
nor U3976 (N_3976,In_2055,In_1985);
and U3977 (N_3977,In_2060,In_1226);
nand U3978 (N_3978,In_2344,In_2470);
nand U3979 (N_3979,In_1476,In_2708);
or U3980 (N_3980,In_2386,In_2900);
and U3981 (N_3981,In_2829,In_1441);
nor U3982 (N_3982,In_2471,In_2045);
and U3983 (N_3983,In_2048,In_782);
and U3984 (N_3984,In_2410,In_522);
and U3985 (N_3985,In_1060,In_2153);
and U3986 (N_3986,In_2274,In_546);
nor U3987 (N_3987,In_123,In_1290);
nor U3988 (N_3988,In_2629,In_1789);
and U3989 (N_3989,In_1834,In_1666);
nand U3990 (N_3990,In_1917,In_606);
and U3991 (N_3991,In_479,In_564);
nand U3992 (N_3992,In_186,In_653);
or U3993 (N_3993,In_696,In_462);
nand U3994 (N_3994,In_818,In_947);
nand U3995 (N_3995,In_2667,In_1296);
or U3996 (N_3996,In_242,In_2518);
xnor U3997 (N_3997,In_1660,In_1232);
xnor U3998 (N_3998,In_1649,In_439);
xnor U3999 (N_3999,In_1785,In_2842);
or U4000 (N_4000,In_650,In_1995);
nand U4001 (N_4001,In_2355,In_1374);
nor U4002 (N_4002,In_2471,In_1705);
nand U4003 (N_4003,In_1860,In_282);
nor U4004 (N_4004,In_2520,In_1878);
nor U4005 (N_4005,In_326,In_2819);
nor U4006 (N_4006,In_1053,In_2279);
nor U4007 (N_4007,In_1400,In_1848);
and U4008 (N_4008,In_1664,In_2652);
nor U4009 (N_4009,In_273,In_1303);
and U4010 (N_4010,In_1117,In_2443);
or U4011 (N_4011,In_2663,In_1260);
nor U4012 (N_4012,In_1246,In_1800);
or U4013 (N_4013,In_1645,In_2363);
and U4014 (N_4014,In_207,In_1564);
nor U4015 (N_4015,In_2526,In_403);
nor U4016 (N_4016,In_1595,In_2339);
xnor U4017 (N_4017,In_2972,In_2981);
or U4018 (N_4018,In_900,In_2763);
xnor U4019 (N_4019,In_2290,In_1936);
or U4020 (N_4020,In_2564,In_943);
xnor U4021 (N_4021,In_1008,In_1398);
or U4022 (N_4022,In_1960,In_946);
and U4023 (N_4023,In_928,In_2477);
nor U4024 (N_4024,In_2940,In_2296);
and U4025 (N_4025,In_2040,In_2107);
nor U4026 (N_4026,In_470,In_2994);
xor U4027 (N_4027,In_1822,In_130);
nor U4028 (N_4028,In_510,In_2015);
nor U4029 (N_4029,In_13,In_2357);
or U4030 (N_4030,In_490,In_2238);
nand U4031 (N_4031,In_2866,In_1249);
nand U4032 (N_4032,In_2693,In_1959);
xor U4033 (N_4033,In_1375,In_291);
nand U4034 (N_4034,In_164,In_2472);
nor U4035 (N_4035,In_1009,In_2262);
nand U4036 (N_4036,In_663,In_1723);
and U4037 (N_4037,In_520,In_2211);
xor U4038 (N_4038,In_992,In_1409);
or U4039 (N_4039,In_2694,In_1278);
or U4040 (N_4040,In_338,In_74);
nor U4041 (N_4041,In_2078,In_1141);
xor U4042 (N_4042,In_745,In_2442);
xnor U4043 (N_4043,In_1196,In_695);
and U4044 (N_4044,In_1741,In_1794);
nor U4045 (N_4045,In_2656,In_198);
xnor U4046 (N_4046,In_171,In_1910);
nor U4047 (N_4047,In_283,In_74);
nor U4048 (N_4048,In_2677,In_62);
or U4049 (N_4049,In_2322,In_1860);
nor U4050 (N_4050,In_1553,In_811);
and U4051 (N_4051,In_2088,In_2807);
nor U4052 (N_4052,In_2243,In_2539);
nor U4053 (N_4053,In_1347,In_1446);
and U4054 (N_4054,In_405,In_1029);
nand U4055 (N_4055,In_1822,In_1946);
nor U4056 (N_4056,In_743,In_1414);
nand U4057 (N_4057,In_817,In_2533);
nor U4058 (N_4058,In_2126,In_2994);
nor U4059 (N_4059,In_1219,In_657);
xor U4060 (N_4060,In_315,In_725);
xnor U4061 (N_4061,In_136,In_2589);
and U4062 (N_4062,In_688,In_1999);
nand U4063 (N_4063,In_1317,In_754);
nor U4064 (N_4064,In_1208,In_2830);
nand U4065 (N_4065,In_2325,In_1505);
nor U4066 (N_4066,In_987,In_1155);
and U4067 (N_4067,In_1125,In_152);
and U4068 (N_4068,In_700,In_685);
xor U4069 (N_4069,In_983,In_2472);
and U4070 (N_4070,In_2299,In_1918);
or U4071 (N_4071,In_2951,In_2010);
nor U4072 (N_4072,In_185,In_93);
xor U4073 (N_4073,In_343,In_2726);
xor U4074 (N_4074,In_2820,In_4);
xnor U4075 (N_4075,In_1541,In_2140);
xor U4076 (N_4076,In_2348,In_137);
nand U4077 (N_4077,In_268,In_2918);
or U4078 (N_4078,In_2753,In_1867);
nand U4079 (N_4079,In_1875,In_1273);
xnor U4080 (N_4080,In_986,In_2300);
nor U4081 (N_4081,In_2198,In_1515);
nand U4082 (N_4082,In_2671,In_954);
xnor U4083 (N_4083,In_1970,In_1609);
nor U4084 (N_4084,In_1524,In_181);
xor U4085 (N_4085,In_342,In_481);
or U4086 (N_4086,In_559,In_1604);
xnor U4087 (N_4087,In_2051,In_969);
nor U4088 (N_4088,In_2627,In_1094);
nand U4089 (N_4089,In_181,In_322);
or U4090 (N_4090,In_851,In_1492);
nor U4091 (N_4091,In_2977,In_1852);
nand U4092 (N_4092,In_1538,In_1632);
nand U4093 (N_4093,In_808,In_1928);
or U4094 (N_4094,In_2673,In_989);
or U4095 (N_4095,In_2767,In_1349);
and U4096 (N_4096,In_1615,In_1443);
nand U4097 (N_4097,In_1668,In_1677);
xor U4098 (N_4098,In_2285,In_287);
xnor U4099 (N_4099,In_2491,In_987);
or U4100 (N_4100,In_1889,In_855);
nand U4101 (N_4101,In_2627,In_926);
xnor U4102 (N_4102,In_2175,In_2810);
nor U4103 (N_4103,In_1202,In_364);
or U4104 (N_4104,In_484,In_282);
nor U4105 (N_4105,In_2721,In_2481);
or U4106 (N_4106,In_913,In_1849);
nand U4107 (N_4107,In_252,In_2257);
nor U4108 (N_4108,In_1877,In_1737);
or U4109 (N_4109,In_2047,In_1975);
nand U4110 (N_4110,In_1293,In_1088);
and U4111 (N_4111,In_1168,In_2814);
xnor U4112 (N_4112,In_1301,In_1066);
xor U4113 (N_4113,In_782,In_2134);
xor U4114 (N_4114,In_838,In_1252);
or U4115 (N_4115,In_1086,In_841);
nor U4116 (N_4116,In_705,In_1314);
or U4117 (N_4117,In_1171,In_2284);
xor U4118 (N_4118,In_2395,In_521);
xor U4119 (N_4119,In_500,In_15);
xnor U4120 (N_4120,In_1904,In_2171);
or U4121 (N_4121,In_1518,In_1905);
nor U4122 (N_4122,In_1292,In_593);
or U4123 (N_4123,In_2317,In_2398);
nand U4124 (N_4124,In_2695,In_12);
and U4125 (N_4125,In_435,In_193);
nor U4126 (N_4126,In_2145,In_404);
nand U4127 (N_4127,In_1421,In_1229);
nor U4128 (N_4128,In_1652,In_2207);
and U4129 (N_4129,In_2568,In_2976);
xnor U4130 (N_4130,In_2195,In_1863);
nor U4131 (N_4131,In_76,In_1418);
and U4132 (N_4132,In_971,In_2319);
or U4133 (N_4133,In_2460,In_657);
nor U4134 (N_4134,In_1156,In_2692);
nand U4135 (N_4135,In_2567,In_1237);
xor U4136 (N_4136,In_1775,In_1732);
or U4137 (N_4137,In_1288,In_2031);
xnor U4138 (N_4138,In_802,In_299);
or U4139 (N_4139,In_1290,In_351);
nor U4140 (N_4140,In_630,In_10);
nand U4141 (N_4141,In_1491,In_1606);
xnor U4142 (N_4142,In_2646,In_2296);
or U4143 (N_4143,In_1707,In_2777);
or U4144 (N_4144,In_2961,In_2182);
nand U4145 (N_4145,In_1775,In_2641);
nand U4146 (N_4146,In_1285,In_751);
or U4147 (N_4147,In_1767,In_1370);
nand U4148 (N_4148,In_843,In_1770);
and U4149 (N_4149,In_2911,In_1044);
xnor U4150 (N_4150,In_1087,In_1040);
nor U4151 (N_4151,In_1042,In_92);
xor U4152 (N_4152,In_2434,In_242);
nor U4153 (N_4153,In_2095,In_2660);
nor U4154 (N_4154,In_1115,In_651);
nor U4155 (N_4155,In_2117,In_1561);
nand U4156 (N_4156,In_1443,In_1588);
and U4157 (N_4157,In_1063,In_1166);
nor U4158 (N_4158,In_1366,In_548);
or U4159 (N_4159,In_1969,In_1606);
nand U4160 (N_4160,In_1527,In_2499);
nand U4161 (N_4161,In_552,In_473);
or U4162 (N_4162,In_1756,In_967);
xnor U4163 (N_4163,In_1351,In_2712);
and U4164 (N_4164,In_1671,In_2788);
xor U4165 (N_4165,In_2246,In_765);
and U4166 (N_4166,In_2321,In_589);
nand U4167 (N_4167,In_2603,In_2800);
nand U4168 (N_4168,In_647,In_836);
and U4169 (N_4169,In_357,In_781);
or U4170 (N_4170,In_987,In_2614);
nor U4171 (N_4171,In_1834,In_2023);
and U4172 (N_4172,In_694,In_118);
xnor U4173 (N_4173,In_2195,In_2258);
nor U4174 (N_4174,In_2359,In_368);
nand U4175 (N_4175,In_412,In_1280);
xnor U4176 (N_4176,In_2575,In_2429);
xnor U4177 (N_4177,In_56,In_204);
and U4178 (N_4178,In_1280,In_1297);
xor U4179 (N_4179,In_974,In_1016);
or U4180 (N_4180,In_1415,In_2053);
nor U4181 (N_4181,In_1232,In_1641);
and U4182 (N_4182,In_474,In_417);
and U4183 (N_4183,In_2802,In_1117);
or U4184 (N_4184,In_863,In_2163);
nand U4185 (N_4185,In_1711,In_1271);
nand U4186 (N_4186,In_2717,In_1657);
xor U4187 (N_4187,In_2931,In_1488);
or U4188 (N_4188,In_2803,In_2166);
xnor U4189 (N_4189,In_153,In_2169);
xor U4190 (N_4190,In_1686,In_6);
xnor U4191 (N_4191,In_2313,In_715);
and U4192 (N_4192,In_2067,In_514);
or U4193 (N_4193,In_1499,In_1271);
and U4194 (N_4194,In_2677,In_300);
nand U4195 (N_4195,In_2860,In_2799);
and U4196 (N_4196,In_1864,In_2715);
nor U4197 (N_4197,In_442,In_1299);
nor U4198 (N_4198,In_991,In_338);
xnor U4199 (N_4199,In_1750,In_2075);
nand U4200 (N_4200,In_698,In_1743);
nor U4201 (N_4201,In_768,In_893);
and U4202 (N_4202,In_1728,In_27);
nand U4203 (N_4203,In_1960,In_669);
xor U4204 (N_4204,In_1055,In_1832);
or U4205 (N_4205,In_1737,In_2917);
nand U4206 (N_4206,In_2220,In_1547);
xor U4207 (N_4207,In_2011,In_57);
xor U4208 (N_4208,In_2170,In_2010);
or U4209 (N_4209,In_2875,In_2165);
nand U4210 (N_4210,In_2943,In_1185);
or U4211 (N_4211,In_1459,In_266);
xor U4212 (N_4212,In_2132,In_958);
xnor U4213 (N_4213,In_143,In_2324);
nand U4214 (N_4214,In_947,In_2570);
or U4215 (N_4215,In_2877,In_970);
xor U4216 (N_4216,In_2936,In_2860);
and U4217 (N_4217,In_1644,In_241);
nor U4218 (N_4218,In_2239,In_748);
nor U4219 (N_4219,In_793,In_470);
xor U4220 (N_4220,In_2575,In_397);
nor U4221 (N_4221,In_1707,In_1143);
or U4222 (N_4222,In_1908,In_535);
or U4223 (N_4223,In_1665,In_586);
xnor U4224 (N_4224,In_816,In_493);
and U4225 (N_4225,In_2547,In_2907);
or U4226 (N_4226,In_2587,In_2071);
nor U4227 (N_4227,In_870,In_659);
nor U4228 (N_4228,In_2635,In_1940);
nor U4229 (N_4229,In_1832,In_2701);
or U4230 (N_4230,In_1214,In_2517);
xor U4231 (N_4231,In_2561,In_690);
nor U4232 (N_4232,In_480,In_2741);
nand U4233 (N_4233,In_2234,In_1514);
and U4234 (N_4234,In_1006,In_2074);
xor U4235 (N_4235,In_145,In_2385);
nor U4236 (N_4236,In_2953,In_837);
or U4237 (N_4237,In_1847,In_1652);
nand U4238 (N_4238,In_1723,In_2640);
and U4239 (N_4239,In_1632,In_1512);
or U4240 (N_4240,In_198,In_2528);
xnor U4241 (N_4241,In_2434,In_602);
nor U4242 (N_4242,In_2711,In_0);
and U4243 (N_4243,In_2010,In_327);
and U4244 (N_4244,In_1837,In_2106);
nor U4245 (N_4245,In_391,In_225);
nand U4246 (N_4246,In_2408,In_832);
xnor U4247 (N_4247,In_296,In_1241);
xor U4248 (N_4248,In_2048,In_2186);
and U4249 (N_4249,In_141,In_243);
nor U4250 (N_4250,In_903,In_2596);
xnor U4251 (N_4251,In_2240,In_2641);
nor U4252 (N_4252,In_2734,In_1054);
and U4253 (N_4253,In_1590,In_241);
or U4254 (N_4254,In_68,In_1748);
nor U4255 (N_4255,In_1394,In_1417);
nand U4256 (N_4256,In_2671,In_2288);
xor U4257 (N_4257,In_1790,In_683);
xnor U4258 (N_4258,In_547,In_1086);
or U4259 (N_4259,In_1460,In_2073);
or U4260 (N_4260,In_707,In_2617);
xnor U4261 (N_4261,In_63,In_1014);
or U4262 (N_4262,In_398,In_905);
or U4263 (N_4263,In_1247,In_1177);
nor U4264 (N_4264,In_1053,In_1411);
nor U4265 (N_4265,In_1281,In_183);
nand U4266 (N_4266,In_2361,In_2780);
or U4267 (N_4267,In_735,In_1177);
or U4268 (N_4268,In_149,In_1471);
nor U4269 (N_4269,In_543,In_2861);
or U4270 (N_4270,In_2782,In_1670);
or U4271 (N_4271,In_942,In_1111);
nor U4272 (N_4272,In_2452,In_839);
xnor U4273 (N_4273,In_715,In_1555);
or U4274 (N_4274,In_1442,In_1224);
xor U4275 (N_4275,In_2615,In_2758);
nor U4276 (N_4276,In_2377,In_592);
and U4277 (N_4277,In_2777,In_1540);
nand U4278 (N_4278,In_1858,In_879);
xor U4279 (N_4279,In_1019,In_634);
and U4280 (N_4280,In_309,In_1002);
or U4281 (N_4281,In_2687,In_836);
nor U4282 (N_4282,In_2157,In_1613);
nand U4283 (N_4283,In_1775,In_2901);
nand U4284 (N_4284,In_193,In_2069);
and U4285 (N_4285,In_214,In_1234);
or U4286 (N_4286,In_2168,In_377);
nand U4287 (N_4287,In_768,In_1916);
and U4288 (N_4288,In_321,In_19);
nand U4289 (N_4289,In_2621,In_983);
and U4290 (N_4290,In_10,In_1838);
or U4291 (N_4291,In_1276,In_1804);
xnor U4292 (N_4292,In_2830,In_2370);
or U4293 (N_4293,In_2991,In_1232);
nor U4294 (N_4294,In_2453,In_222);
and U4295 (N_4295,In_2846,In_1499);
nand U4296 (N_4296,In_1020,In_2202);
and U4297 (N_4297,In_1784,In_1088);
or U4298 (N_4298,In_2534,In_0);
nand U4299 (N_4299,In_929,In_2313);
nand U4300 (N_4300,In_926,In_2828);
and U4301 (N_4301,In_2188,In_1422);
and U4302 (N_4302,In_649,In_2178);
nand U4303 (N_4303,In_989,In_1890);
nand U4304 (N_4304,In_2820,In_1917);
and U4305 (N_4305,In_916,In_2510);
or U4306 (N_4306,In_590,In_843);
nor U4307 (N_4307,In_557,In_1773);
and U4308 (N_4308,In_2046,In_1397);
nor U4309 (N_4309,In_2131,In_131);
or U4310 (N_4310,In_894,In_200);
nor U4311 (N_4311,In_1960,In_1744);
or U4312 (N_4312,In_193,In_2705);
nand U4313 (N_4313,In_809,In_308);
or U4314 (N_4314,In_2844,In_2880);
or U4315 (N_4315,In_293,In_1008);
xnor U4316 (N_4316,In_1173,In_1730);
nor U4317 (N_4317,In_1346,In_1439);
nor U4318 (N_4318,In_861,In_64);
xor U4319 (N_4319,In_910,In_176);
nor U4320 (N_4320,In_2209,In_2906);
nor U4321 (N_4321,In_304,In_424);
or U4322 (N_4322,In_2570,In_2269);
and U4323 (N_4323,In_2978,In_2647);
or U4324 (N_4324,In_2750,In_1753);
nand U4325 (N_4325,In_299,In_33);
nor U4326 (N_4326,In_1455,In_387);
nor U4327 (N_4327,In_2193,In_1995);
nor U4328 (N_4328,In_2005,In_1975);
and U4329 (N_4329,In_1476,In_2387);
and U4330 (N_4330,In_152,In_2851);
or U4331 (N_4331,In_1057,In_2225);
xor U4332 (N_4332,In_1291,In_2231);
or U4333 (N_4333,In_2533,In_1496);
xnor U4334 (N_4334,In_2213,In_2093);
xnor U4335 (N_4335,In_1873,In_863);
and U4336 (N_4336,In_484,In_1692);
nor U4337 (N_4337,In_1376,In_2947);
nor U4338 (N_4338,In_1874,In_367);
nor U4339 (N_4339,In_865,In_2046);
nor U4340 (N_4340,In_2803,In_1721);
or U4341 (N_4341,In_2275,In_1452);
nor U4342 (N_4342,In_448,In_1514);
and U4343 (N_4343,In_771,In_2247);
and U4344 (N_4344,In_1647,In_1635);
nand U4345 (N_4345,In_864,In_2267);
nand U4346 (N_4346,In_555,In_1896);
and U4347 (N_4347,In_306,In_1072);
nor U4348 (N_4348,In_734,In_53);
and U4349 (N_4349,In_2964,In_164);
nand U4350 (N_4350,In_1333,In_1230);
and U4351 (N_4351,In_101,In_1046);
or U4352 (N_4352,In_1435,In_575);
xnor U4353 (N_4353,In_2942,In_506);
and U4354 (N_4354,In_938,In_2404);
nand U4355 (N_4355,In_868,In_2364);
xor U4356 (N_4356,In_624,In_2161);
nand U4357 (N_4357,In_172,In_2515);
and U4358 (N_4358,In_2164,In_1800);
nand U4359 (N_4359,In_1272,In_1143);
nand U4360 (N_4360,In_1749,In_2060);
nand U4361 (N_4361,In_1148,In_2798);
nor U4362 (N_4362,In_1366,In_2710);
nand U4363 (N_4363,In_639,In_145);
or U4364 (N_4364,In_1755,In_669);
xor U4365 (N_4365,In_767,In_2083);
nor U4366 (N_4366,In_1410,In_1856);
nor U4367 (N_4367,In_1693,In_564);
xor U4368 (N_4368,In_2602,In_1722);
nand U4369 (N_4369,In_2472,In_2853);
nand U4370 (N_4370,In_1412,In_1291);
and U4371 (N_4371,In_497,In_1648);
xnor U4372 (N_4372,In_209,In_1531);
xnor U4373 (N_4373,In_113,In_72);
nand U4374 (N_4374,In_644,In_893);
or U4375 (N_4375,In_2502,In_2730);
or U4376 (N_4376,In_1358,In_529);
xor U4377 (N_4377,In_2997,In_90);
nor U4378 (N_4378,In_2476,In_547);
nand U4379 (N_4379,In_2706,In_2258);
nand U4380 (N_4380,In_2414,In_2841);
nor U4381 (N_4381,In_2394,In_2503);
nand U4382 (N_4382,In_1305,In_2278);
nor U4383 (N_4383,In_251,In_2743);
xor U4384 (N_4384,In_618,In_1492);
nor U4385 (N_4385,In_920,In_2952);
and U4386 (N_4386,In_2302,In_986);
nand U4387 (N_4387,In_915,In_1538);
or U4388 (N_4388,In_2329,In_2848);
nand U4389 (N_4389,In_2439,In_269);
xnor U4390 (N_4390,In_1781,In_605);
nand U4391 (N_4391,In_819,In_1369);
nand U4392 (N_4392,In_482,In_1543);
nor U4393 (N_4393,In_2739,In_1501);
nand U4394 (N_4394,In_652,In_2549);
nor U4395 (N_4395,In_621,In_150);
or U4396 (N_4396,In_934,In_2383);
nor U4397 (N_4397,In_436,In_1344);
nand U4398 (N_4398,In_207,In_1982);
nand U4399 (N_4399,In_1464,In_26);
xor U4400 (N_4400,In_2950,In_845);
xor U4401 (N_4401,In_2277,In_323);
nor U4402 (N_4402,In_2621,In_1081);
xor U4403 (N_4403,In_2846,In_2619);
nor U4404 (N_4404,In_2507,In_942);
or U4405 (N_4405,In_2900,In_1594);
nor U4406 (N_4406,In_663,In_1925);
and U4407 (N_4407,In_1609,In_2014);
or U4408 (N_4408,In_396,In_1159);
and U4409 (N_4409,In_1915,In_2231);
nor U4410 (N_4410,In_805,In_1165);
and U4411 (N_4411,In_363,In_212);
nand U4412 (N_4412,In_1625,In_879);
xor U4413 (N_4413,In_634,In_2294);
or U4414 (N_4414,In_2724,In_1371);
or U4415 (N_4415,In_2391,In_210);
nand U4416 (N_4416,In_1387,In_2838);
nand U4417 (N_4417,In_342,In_1103);
or U4418 (N_4418,In_357,In_1731);
xnor U4419 (N_4419,In_1121,In_1114);
or U4420 (N_4420,In_664,In_2712);
xor U4421 (N_4421,In_640,In_2026);
or U4422 (N_4422,In_1992,In_2662);
nand U4423 (N_4423,In_1769,In_1345);
nor U4424 (N_4424,In_645,In_1014);
nor U4425 (N_4425,In_2277,In_1458);
or U4426 (N_4426,In_2297,In_1251);
xnor U4427 (N_4427,In_2015,In_2122);
nor U4428 (N_4428,In_467,In_1046);
xor U4429 (N_4429,In_2549,In_2092);
nor U4430 (N_4430,In_2651,In_2088);
nand U4431 (N_4431,In_2306,In_448);
or U4432 (N_4432,In_2747,In_2031);
and U4433 (N_4433,In_960,In_2895);
nand U4434 (N_4434,In_2849,In_420);
and U4435 (N_4435,In_2300,In_2813);
nor U4436 (N_4436,In_1447,In_1111);
and U4437 (N_4437,In_1108,In_2947);
or U4438 (N_4438,In_470,In_884);
nand U4439 (N_4439,In_1857,In_812);
or U4440 (N_4440,In_656,In_870);
nor U4441 (N_4441,In_1749,In_1608);
nor U4442 (N_4442,In_2435,In_927);
or U4443 (N_4443,In_643,In_511);
and U4444 (N_4444,In_1149,In_2595);
xnor U4445 (N_4445,In_1251,In_349);
nor U4446 (N_4446,In_2509,In_717);
and U4447 (N_4447,In_1191,In_861);
xor U4448 (N_4448,In_2407,In_1587);
or U4449 (N_4449,In_648,In_2555);
xnor U4450 (N_4450,In_1792,In_2701);
and U4451 (N_4451,In_1229,In_1006);
xnor U4452 (N_4452,In_174,In_2562);
nor U4453 (N_4453,In_1019,In_650);
xor U4454 (N_4454,In_1486,In_907);
nor U4455 (N_4455,In_367,In_1787);
xnor U4456 (N_4456,In_304,In_218);
nor U4457 (N_4457,In_1939,In_2389);
or U4458 (N_4458,In_920,In_244);
or U4459 (N_4459,In_982,In_527);
nand U4460 (N_4460,In_1033,In_919);
nor U4461 (N_4461,In_2349,In_2767);
or U4462 (N_4462,In_2948,In_1858);
or U4463 (N_4463,In_1077,In_981);
xor U4464 (N_4464,In_2936,In_1138);
and U4465 (N_4465,In_71,In_2762);
and U4466 (N_4466,In_782,In_2841);
xnor U4467 (N_4467,In_2670,In_528);
and U4468 (N_4468,In_128,In_122);
or U4469 (N_4469,In_1882,In_2337);
nor U4470 (N_4470,In_2079,In_680);
and U4471 (N_4471,In_725,In_1884);
xor U4472 (N_4472,In_1786,In_32);
or U4473 (N_4473,In_1939,In_1986);
xor U4474 (N_4474,In_1208,In_997);
nor U4475 (N_4475,In_2654,In_2889);
and U4476 (N_4476,In_392,In_2824);
or U4477 (N_4477,In_1008,In_1144);
and U4478 (N_4478,In_2446,In_2212);
nor U4479 (N_4479,In_1347,In_2738);
nand U4480 (N_4480,In_2592,In_128);
and U4481 (N_4481,In_395,In_2608);
or U4482 (N_4482,In_1394,In_1407);
or U4483 (N_4483,In_349,In_910);
nor U4484 (N_4484,In_1162,In_1884);
xnor U4485 (N_4485,In_2725,In_1108);
or U4486 (N_4486,In_2626,In_2975);
and U4487 (N_4487,In_500,In_1155);
nand U4488 (N_4488,In_1835,In_1314);
nand U4489 (N_4489,In_2176,In_1644);
nor U4490 (N_4490,In_473,In_851);
xnor U4491 (N_4491,In_1202,In_1200);
nor U4492 (N_4492,In_2759,In_1109);
xnor U4493 (N_4493,In_559,In_1942);
nand U4494 (N_4494,In_313,In_135);
xnor U4495 (N_4495,In_1605,In_2016);
or U4496 (N_4496,In_1919,In_325);
xor U4497 (N_4497,In_738,In_2778);
nand U4498 (N_4498,In_1037,In_664);
xnor U4499 (N_4499,In_2350,In_752);
and U4500 (N_4500,In_2407,In_2453);
or U4501 (N_4501,In_1744,In_1734);
xor U4502 (N_4502,In_1443,In_335);
xnor U4503 (N_4503,In_481,In_879);
nor U4504 (N_4504,In_850,In_1715);
or U4505 (N_4505,In_2322,In_374);
xor U4506 (N_4506,In_2860,In_2870);
and U4507 (N_4507,In_921,In_1146);
or U4508 (N_4508,In_1267,In_917);
nor U4509 (N_4509,In_62,In_1969);
and U4510 (N_4510,In_2264,In_321);
nand U4511 (N_4511,In_2926,In_644);
and U4512 (N_4512,In_1508,In_397);
and U4513 (N_4513,In_2434,In_2773);
nand U4514 (N_4514,In_2010,In_177);
nand U4515 (N_4515,In_1109,In_2928);
and U4516 (N_4516,In_1751,In_2701);
nor U4517 (N_4517,In_1093,In_1702);
nand U4518 (N_4518,In_694,In_617);
xor U4519 (N_4519,In_1551,In_1013);
nand U4520 (N_4520,In_2539,In_1920);
nand U4521 (N_4521,In_2535,In_1718);
and U4522 (N_4522,In_2255,In_294);
and U4523 (N_4523,In_2741,In_365);
xor U4524 (N_4524,In_1557,In_1463);
nor U4525 (N_4525,In_965,In_778);
xor U4526 (N_4526,In_223,In_2145);
or U4527 (N_4527,In_127,In_780);
nor U4528 (N_4528,In_1730,In_1527);
nand U4529 (N_4529,In_2475,In_2055);
and U4530 (N_4530,In_1424,In_903);
nand U4531 (N_4531,In_2222,In_2162);
nor U4532 (N_4532,In_1752,In_2886);
or U4533 (N_4533,In_2296,In_323);
xor U4534 (N_4534,In_523,In_929);
and U4535 (N_4535,In_1920,In_756);
xnor U4536 (N_4536,In_2714,In_2649);
xnor U4537 (N_4537,In_1168,In_2533);
and U4538 (N_4538,In_1117,In_1810);
nor U4539 (N_4539,In_1299,In_2624);
nor U4540 (N_4540,In_1579,In_86);
or U4541 (N_4541,In_2982,In_2012);
nand U4542 (N_4542,In_575,In_2985);
nor U4543 (N_4543,In_2,In_346);
nand U4544 (N_4544,In_1715,In_1212);
xor U4545 (N_4545,In_553,In_1133);
nand U4546 (N_4546,In_2015,In_770);
and U4547 (N_4547,In_2626,In_2235);
xor U4548 (N_4548,In_2386,In_1206);
nand U4549 (N_4549,In_1013,In_1754);
nor U4550 (N_4550,In_1390,In_2709);
and U4551 (N_4551,In_2256,In_2153);
xnor U4552 (N_4552,In_436,In_1374);
or U4553 (N_4553,In_639,In_853);
nand U4554 (N_4554,In_2368,In_2007);
or U4555 (N_4555,In_1834,In_1238);
or U4556 (N_4556,In_1518,In_2998);
nand U4557 (N_4557,In_1706,In_204);
and U4558 (N_4558,In_1095,In_724);
and U4559 (N_4559,In_1677,In_1038);
nand U4560 (N_4560,In_806,In_1890);
or U4561 (N_4561,In_2876,In_2439);
nand U4562 (N_4562,In_2907,In_2905);
nor U4563 (N_4563,In_2572,In_829);
xor U4564 (N_4564,In_2364,In_2582);
and U4565 (N_4565,In_822,In_1850);
nand U4566 (N_4566,In_1120,In_2633);
nor U4567 (N_4567,In_1395,In_1142);
xor U4568 (N_4568,In_616,In_2307);
and U4569 (N_4569,In_2395,In_1465);
xnor U4570 (N_4570,In_943,In_2057);
nand U4571 (N_4571,In_2649,In_2894);
or U4572 (N_4572,In_2635,In_244);
or U4573 (N_4573,In_1096,In_682);
or U4574 (N_4574,In_748,In_2833);
or U4575 (N_4575,In_745,In_470);
nand U4576 (N_4576,In_1062,In_2059);
and U4577 (N_4577,In_2947,In_2642);
nand U4578 (N_4578,In_2833,In_293);
nand U4579 (N_4579,In_282,In_1137);
nand U4580 (N_4580,In_2891,In_2748);
xor U4581 (N_4581,In_130,In_1146);
nand U4582 (N_4582,In_1323,In_2001);
xnor U4583 (N_4583,In_2333,In_217);
or U4584 (N_4584,In_2204,In_1393);
nand U4585 (N_4585,In_1732,In_823);
xnor U4586 (N_4586,In_2023,In_2612);
xnor U4587 (N_4587,In_843,In_2800);
or U4588 (N_4588,In_1800,In_1729);
and U4589 (N_4589,In_702,In_372);
or U4590 (N_4590,In_352,In_78);
or U4591 (N_4591,In_1081,In_2840);
nor U4592 (N_4592,In_2124,In_1786);
and U4593 (N_4593,In_579,In_1841);
nand U4594 (N_4594,In_1719,In_2168);
nor U4595 (N_4595,In_1985,In_2012);
xor U4596 (N_4596,In_1515,In_999);
nand U4597 (N_4597,In_2137,In_2493);
xnor U4598 (N_4598,In_2329,In_2968);
nor U4599 (N_4599,In_1938,In_0);
xnor U4600 (N_4600,In_157,In_2841);
xnor U4601 (N_4601,In_680,In_833);
nand U4602 (N_4602,In_1511,In_2828);
xor U4603 (N_4603,In_70,In_159);
or U4604 (N_4604,In_2503,In_144);
and U4605 (N_4605,In_1874,In_1985);
or U4606 (N_4606,In_2592,In_1229);
nand U4607 (N_4607,In_1261,In_828);
and U4608 (N_4608,In_2691,In_2728);
xor U4609 (N_4609,In_607,In_245);
nand U4610 (N_4610,In_1915,In_1319);
nor U4611 (N_4611,In_1939,In_2640);
nand U4612 (N_4612,In_1981,In_2889);
and U4613 (N_4613,In_2774,In_738);
nand U4614 (N_4614,In_1405,In_1448);
xnor U4615 (N_4615,In_97,In_295);
nor U4616 (N_4616,In_1366,In_2114);
nor U4617 (N_4617,In_2356,In_2139);
and U4618 (N_4618,In_1585,In_366);
xnor U4619 (N_4619,In_1175,In_1671);
and U4620 (N_4620,In_132,In_637);
and U4621 (N_4621,In_742,In_411);
xnor U4622 (N_4622,In_1399,In_990);
nor U4623 (N_4623,In_2079,In_1469);
and U4624 (N_4624,In_1806,In_1922);
nor U4625 (N_4625,In_2834,In_262);
or U4626 (N_4626,In_48,In_220);
nand U4627 (N_4627,In_1276,In_2908);
and U4628 (N_4628,In_2808,In_2935);
nor U4629 (N_4629,In_54,In_427);
nor U4630 (N_4630,In_2669,In_2647);
or U4631 (N_4631,In_2858,In_1062);
nor U4632 (N_4632,In_2369,In_1066);
nor U4633 (N_4633,In_1903,In_1136);
nor U4634 (N_4634,In_1194,In_1979);
xnor U4635 (N_4635,In_2593,In_1047);
or U4636 (N_4636,In_2049,In_2262);
nor U4637 (N_4637,In_1079,In_1913);
or U4638 (N_4638,In_1548,In_2796);
xor U4639 (N_4639,In_133,In_1194);
nand U4640 (N_4640,In_827,In_1080);
nor U4641 (N_4641,In_755,In_460);
or U4642 (N_4642,In_2835,In_2971);
nor U4643 (N_4643,In_2733,In_1930);
or U4644 (N_4644,In_2768,In_1815);
or U4645 (N_4645,In_2884,In_2035);
nand U4646 (N_4646,In_2680,In_641);
xnor U4647 (N_4647,In_2173,In_2460);
and U4648 (N_4648,In_1658,In_317);
nand U4649 (N_4649,In_345,In_505);
nor U4650 (N_4650,In_1792,In_252);
xnor U4651 (N_4651,In_2684,In_1842);
nor U4652 (N_4652,In_2339,In_988);
nor U4653 (N_4653,In_145,In_1898);
nor U4654 (N_4654,In_7,In_1321);
xor U4655 (N_4655,In_2317,In_2402);
xor U4656 (N_4656,In_2101,In_1446);
nor U4657 (N_4657,In_2573,In_2156);
nor U4658 (N_4658,In_457,In_1993);
nand U4659 (N_4659,In_1803,In_2452);
xor U4660 (N_4660,In_2741,In_236);
xnor U4661 (N_4661,In_2554,In_1059);
or U4662 (N_4662,In_1870,In_583);
nand U4663 (N_4663,In_2352,In_1563);
and U4664 (N_4664,In_1587,In_836);
nand U4665 (N_4665,In_1106,In_1176);
nor U4666 (N_4666,In_604,In_2829);
or U4667 (N_4667,In_2300,In_2026);
and U4668 (N_4668,In_1061,In_1744);
or U4669 (N_4669,In_2887,In_2933);
xnor U4670 (N_4670,In_16,In_2052);
xnor U4671 (N_4671,In_547,In_2387);
xnor U4672 (N_4672,In_2031,In_1600);
and U4673 (N_4673,In_1699,In_549);
xnor U4674 (N_4674,In_7,In_1842);
nand U4675 (N_4675,In_2557,In_612);
nor U4676 (N_4676,In_1409,In_1455);
nand U4677 (N_4677,In_2225,In_1974);
nand U4678 (N_4678,In_423,In_41);
or U4679 (N_4679,In_1734,In_483);
nand U4680 (N_4680,In_571,In_1055);
and U4681 (N_4681,In_170,In_81);
xor U4682 (N_4682,In_1177,In_2721);
and U4683 (N_4683,In_426,In_1399);
nor U4684 (N_4684,In_184,In_416);
or U4685 (N_4685,In_1158,In_1220);
xnor U4686 (N_4686,In_1161,In_90);
nor U4687 (N_4687,In_800,In_2479);
xnor U4688 (N_4688,In_989,In_2761);
and U4689 (N_4689,In_1958,In_1913);
nand U4690 (N_4690,In_1622,In_1581);
or U4691 (N_4691,In_499,In_1194);
nand U4692 (N_4692,In_967,In_156);
nor U4693 (N_4693,In_983,In_1611);
and U4694 (N_4694,In_1732,In_2232);
nand U4695 (N_4695,In_395,In_2286);
xor U4696 (N_4696,In_2692,In_2506);
nor U4697 (N_4697,In_2688,In_341);
nand U4698 (N_4698,In_1572,In_746);
or U4699 (N_4699,In_197,In_427);
nand U4700 (N_4700,In_318,In_2774);
nor U4701 (N_4701,In_2487,In_1749);
nand U4702 (N_4702,In_208,In_2791);
xnor U4703 (N_4703,In_375,In_690);
nor U4704 (N_4704,In_1969,In_1509);
nand U4705 (N_4705,In_2679,In_1724);
or U4706 (N_4706,In_98,In_758);
and U4707 (N_4707,In_2423,In_971);
and U4708 (N_4708,In_2217,In_3);
xnor U4709 (N_4709,In_1738,In_855);
nand U4710 (N_4710,In_2785,In_606);
nor U4711 (N_4711,In_1208,In_277);
or U4712 (N_4712,In_2518,In_342);
and U4713 (N_4713,In_2086,In_1887);
xor U4714 (N_4714,In_1344,In_789);
nor U4715 (N_4715,In_859,In_1635);
xor U4716 (N_4716,In_1675,In_1621);
nand U4717 (N_4717,In_1894,In_1788);
and U4718 (N_4718,In_2811,In_2531);
xnor U4719 (N_4719,In_1300,In_1604);
nor U4720 (N_4720,In_2882,In_1281);
or U4721 (N_4721,In_609,In_1079);
xor U4722 (N_4722,In_1800,In_2912);
nand U4723 (N_4723,In_2753,In_2331);
nand U4724 (N_4724,In_2699,In_1530);
nor U4725 (N_4725,In_210,In_2615);
xnor U4726 (N_4726,In_1602,In_1672);
or U4727 (N_4727,In_2563,In_1851);
nand U4728 (N_4728,In_2296,In_2878);
and U4729 (N_4729,In_1469,In_1754);
and U4730 (N_4730,In_467,In_2243);
nand U4731 (N_4731,In_714,In_2403);
and U4732 (N_4732,In_1626,In_2655);
or U4733 (N_4733,In_1185,In_501);
xnor U4734 (N_4734,In_2267,In_768);
or U4735 (N_4735,In_202,In_1081);
nor U4736 (N_4736,In_1993,In_2321);
or U4737 (N_4737,In_1059,In_1905);
xor U4738 (N_4738,In_981,In_1139);
or U4739 (N_4739,In_879,In_1203);
or U4740 (N_4740,In_197,In_2156);
xnor U4741 (N_4741,In_1592,In_299);
and U4742 (N_4742,In_284,In_1983);
nand U4743 (N_4743,In_1394,In_706);
nand U4744 (N_4744,In_2668,In_2710);
nor U4745 (N_4745,In_2100,In_276);
or U4746 (N_4746,In_1272,In_1035);
and U4747 (N_4747,In_2709,In_579);
or U4748 (N_4748,In_2616,In_3);
and U4749 (N_4749,In_2468,In_2914);
and U4750 (N_4750,In_671,In_757);
nand U4751 (N_4751,In_2629,In_2082);
nand U4752 (N_4752,In_573,In_1006);
xnor U4753 (N_4753,In_1267,In_2281);
nand U4754 (N_4754,In_2137,In_2913);
xor U4755 (N_4755,In_2079,In_2393);
and U4756 (N_4756,In_1360,In_2512);
or U4757 (N_4757,In_1610,In_816);
xnor U4758 (N_4758,In_819,In_1481);
xor U4759 (N_4759,In_143,In_2020);
or U4760 (N_4760,In_2148,In_2896);
and U4761 (N_4761,In_2,In_175);
nand U4762 (N_4762,In_390,In_1362);
nor U4763 (N_4763,In_1012,In_519);
or U4764 (N_4764,In_1005,In_2460);
nand U4765 (N_4765,In_1155,In_2429);
and U4766 (N_4766,In_450,In_1714);
nor U4767 (N_4767,In_341,In_1421);
nor U4768 (N_4768,In_462,In_979);
or U4769 (N_4769,In_2405,In_475);
nand U4770 (N_4770,In_2157,In_1422);
and U4771 (N_4771,In_823,In_2954);
xnor U4772 (N_4772,In_2786,In_741);
xnor U4773 (N_4773,In_210,In_2601);
nor U4774 (N_4774,In_284,In_1253);
nor U4775 (N_4775,In_125,In_2660);
or U4776 (N_4776,In_1678,In_2715);
xnor U4777 (N_4777,In_2727,In_2710);
or U4778 (N_4778,In_1361,In_4);
nand U4779 (N_4779,In_2553,In_1217);
xor U4780 (N_4780,In_266,In_124);
and U4781 (N_4781,In_1321,In_1098);
and U4782 (N_4782,In_2473,In_1545);
and U4783 (N_4783,In_2046,In_2023);
nor U4784 (N_4784,In_2162,In_340);
nand U4785 (N_4785,In_202,In_1840);
nand U4786 (N_4786,In_1449,In_1978);
or U4787 (N_4787,In_2104,In_1135);
nand U4788 (N_4788,In_2129,In_2294);
nor U4789 (N_4789,In_2320,In_4);
xor U4790 (N_4790,In_1391,In_908);
and U4791 (N_4791,In_1597,In_1134);
nor U4792 (N_4792,In_1685,In_2205);
xor U4793 (N_4793,In_242,In_1493);
xor U4794 (N_4794,In_1699,In_510);
nand U4795 (N_4795,In_1143,In_2515);
or U4796 (N_4796,In_565,In_2058);
xnor U4797 (N_4797,In_1797,In_2510);
and U4798 (N_4798,In_1592,In_2924);
xor U4799 (N_4799,In_413,In_2360);
and U4800 (N_4800,In_1573,In_2227);
nor U4801 (N_4801,In_1441,In_2885);
nor U4802 (N_4802,In_2047,In_1908);
or U4803 (N_4803,In_2418,In_309);
xor U4804 (N_4804,In_873,In_2479);
xnor U4805 (N_4805,In_2521,In_1273);
xnor U4806 (N_4806,In_1354,In_1513);
xor U4807 (N_4807,In_1576,In_2397);
or U4808 (N_4808,In_2769,In_2518);
nand U4809 (N_4809,In_641,In_2208);
nor U4810 (N_4810,In_1081,In_862);
or U4811 (N_4811,In_850,In_1398);
nand U4812 (N_4812,In_2647,In_1075);
xor U4813 (N_4813,In_2236,In_2229);
and U4814 (N_4814,In_1324,In_2119);
and U4815 (N_4815,In_876,In_1891);
xor U4816 (N_4816,In_1380,In_2663);
nand U4817 (N_4817,In_504,In_807);
or U4818 (N_4818,In_2143,In_1022);
xnor U4819 (N_4819,In_2947,In_2581);
nor U4820 (N_4820,In_2622,In_451);
nand U4821 (N_4821,In_2915,In_924);
or U4822 (N_4822,In_1063,In_1784);
and U4823 (N_4823,In_151,In_464);
nor U4824 (N_4824,In_980,In_99);
and U4825 (N_4825,In_311,In_2348);
or U4826 (N_4826,In_1293,In_2709);
xnor U4827 (N_4827,In_1072,In_956);
xnor U4828 (N_4828,In_2731,In_1670);
nand U4829 (N_4829,In_1989,In_2019);
or U4830 (N_4830,In_875,In_1065);
and U4831 (N_4831,In_2214,In_783);
nor U4832 (N_4832,In_2459,In_234);
or U4833 (N_4833,In_1166,In_2543);
xnor U4834 (N_4834,In_1550,In_2511);
and U4835 (N_4835,In_286,In_2531);
nor U4836 (N_4836,In_252,In_2989);
and U4837 (N_4837,In_1072,In_1019);
or U4838 (N_4838,In_2913,In_683);
and U4839 (N_4839,In_438,In_2616);
or U4840 (N_4840,In_513,In_550);
and U4841 (N_4841,In_1817,In_2032);
xor U4842 (N_4842,In_2374,In_2081);
or U4843 (N_4843,In_2015,In_694);
nor U4844 (N_4844,In_1173,In_2639);
xor U4845 (N_4845,In_1824,In_946);
and U4846 (N_4846,In_1152,In_322);
nand U4847 (N_4847,In_828,In_2497);
or U4848 (N_4848,In_207,In_1391);
xor U4849 (N_4849,In_705,In_2283);
nand U4850 (N_4850,In_377,In_2589);
nor U4851 (N_4851,In_2504,In_549);
nor U4852 (N_4852,In_104,In_1202);
or U4853 (N_4853,In_2256,In_1831);
xor U4854 (N_4854,In_2377,In_2798);
xnor U4855 (N_4855,In_1285,In_2093);
nor U4856 (N_4856,In_314,In_1399);
or U4857 (N_4857,In_2620,In_2244);
nor U4858 (N_4858,In_327,In_1104);
or U4859 (N_4859,In_285,In_1335);
and U4860 (N_4860,In_1877,In_909);
nand U4861 (N_4861,In_1647,In_1767);
xnor U4862 (N_4862,In_2783,In_1760);
or U4863 (N_4863,In_1266,In_1707);
or U4864 (N_4864,In_1840,In_2937);
nand U4865 (N_4865,In_1227,In_2801);
nor U4866 (N_4866,In_668,In_10);
xor U4867 (N_4867,In_1306,In_1245);
xnor U4868 (N_4868,In_1975,In_84);
nand U4869 (N_4869,In_814,In_262);
or U4870 (N_4870,In_1502,In_471);
or U4871 (N_4871,In_1448,In_8);
xnor U4872 (N_4872,In_400,In_1208);
nand U4873 (N_4873,In_121,In_1297);
nand U4874 (N_4874,In_429,In_2821);
and U4875 (N_4875,In_2689,In_156);
xor U4876 (N_4876,In_1790,In_503);
nand U4877 (N_4877,In_2341,In_2639);
xor U4878 (N_4878,In_1150,In_2512);
nand U4879 (N_4879,In_1787,In_2643);
xnor U4880 (N_4880,In_969,In_950);
and U4881 (N_4881,In_2487,In_2577);
xor U4882 (N_4882,In_2464,In_2517);
xnor U4883 (N_4883,In_2381,In_1432);
nand U4884 (N_4884,In_163,In_2080);
or U4885 (N_4885,In_1572,In_2590);
and U4886 (N_4886,In_2029,In_2671);
nand U4887 (N_4887,In_79,In_541);
xnor U4888 (N_4888,In_766,In_1699);
or U4889 (N_4889,In_890,In_2676);
xnor U4890 (N_4890,In_1473,In_1528);
and U4891 (N_4891,In_120,In_2216);
nand U4892 (N_4892,In_555,In_1);
and U4893 (N_4893,In_704,In_2060);
and U4894 (N_4894,In_818,In_493);
nand U4895 (N_4895,In_1353,In_665);
nand U4896 (N_4896,In_2656,In_2258);
xor U4897 (N_4897,In_1630,In_44);
nand U4898 (N_4898,In_1796,In_2992);
xor U4899 (N_4899,In_2680,In_2910);
and U4900 (N_4900,In_2842,In_1745);
and U4901 (N_4901,In_1433,In_2204);
nand U4902 (N_4902,In_769,In_332);
nand U4903 (N_4903,In_2494,In_2808);
nand U4904 (N_4904,In_1043,In_1234);
or U4905 (N_4905,In_2088,In_1542);
xor U4906 (N_4906,In_98,In_2454);
nor U4907 (N_4907,In_21,In_619);
or U4908 (N_4908,In_1495,In_1639);
and U4909 (N_4909,In_142,In_1418);
xor U4910 (N_4910,In_2527,In_2808);
or U4911 (N_4911,In_1861,In_707);
nand U4912 (N_4912,In_344,In_832);
and U4913 (N_4913,In_1625,In_63);
or U4914 (N_4914,In_1359,In_2915);
or U4915 (N_4915,In_2633,In_2122);
nor U4916 (N_4916,In_1107,In_2559);
nor U4917 (N_4917,In_1681,In_1104);
nor U4918 (N_4918,In_1648,In_1157);
nand U4919 (N_4919,In_2569,In_2932);
nand U4920 (N_4920,In_842,In_538);
or U4921 (N_4921,In_1842,In_2750);
nor U4922 (N_4922,In_255,In_661);
nand U4923 (N_4923,In_1988,In_882);
xor U4924 (N_4924,In_2325,In_907);
and U4925 (N_4925,In_2468,In_2318);
xnor U4926 (N_4926,In_2726,In_1845);
and U4927 (N_4927,In_2430,In_1730);
and U4928 (N_4928,In_785,In_1830);
nor U4929 (N_4929,In_1473,In_493);
nand U4930 (N_4930,In_1154,In_2416);
nand U4931 (N_4931,In_2993,In_825);
and U4932 (N_4932,In_1142,In_2613);
xor U4933 (N_4933,In_2298,In_1606);
and U4934 (N_4934,In_2197,In_999);
nand U4935 (N_4935,In_1311,In_2669);
or U4936 (N_4936,In_1628,In_1739);
and U4937 (N_4937,In_342,In_37);
nor U4938 (N_4938,In_151,In_2939);
nor U4939 (N_4939,In_1995,In_1144);
nor U4940 (N_4940,In_429,In_2288);
xor U4941 (N_4941,In_2998,In_576);
or U4942 (N_4942,In_941,In_817);
nand U4943 (N_4943,In_2970,In_2844);
nand U4944 (N_4944,In_2883,In_1122);
nor U4945 (N_4945,In_395,In_1956);
nand U4946 (N_4946,In_1214,In_2264);
xor U4947 (N_4947,In_1215,In_559);
nor U4948 (N_4948,In_999,In_2890);
nor U4949 (N_4949,In_2433,In_1925);
xor U4950 (N_4950,In_2647,In_897);
nor U4951 (N_4951,In_78,In_2125);
nand U4952 (N_4952,In_1329,In_2948);
xnor U4953 (N_4953,In_2771,In_1419);
nand U4954 (N_4954,In_758,In_1499);
and U4955 (N_4955,In_1910,In_2196);
or U4956 (N_4956,In_34,In_2738);
and U4957 (N_4957,In_1985,In_2067);
and U4958 (N_4958,In_278,In_1655);
nor U4959 (N_4959,In_270,In_417);
or U4960 (N_4960,In_1913,In_2632);
or U4961 (N_4961,In_2991,In_1035);
nand U4962 (N_4962,In_2509,In_1902);
nand U4963 (N_4963,In_2835,In_2772);
and U4964 (N_4964,In_782,In_486);
and U4965 (N_4965,In_1793,In_1989);
nor U4966 (N_4966,In_1522,In_2643);
nand U4967 (N_4967,In_2364,In_1019);
or U4968 (N_4968,In_1447,In_1296);
and U4969 (N_4969,In_1032,In_2749);
nor U4970 (N_4970,In_2269,In_1034);
xor U4971 (N_4971,In_2,In_1533);
nand U4972 (N_4972,In_2343,In_662);
nand U4973 (N_4973,In_200,In_82);
xnor U4974 (N_4974,In_1720,In_1210);
nand U4975 (N_4975,In_2010,In_1167);
xnor U4976 (N_4976,In_1284,In_935);
xor U4977 (N_4977,In_2852,In_2984);
nand U4978 (N_4978,In_540,In_2065);
nand U4979 (N_4979,In_1592,In_2484);
nor U4980 (N_4980,In_43,In_304);
nor U4981 (N_4981,In_2319,In_1213);
and U4982 (N_4982,In_1515,In_2313);
and U4983 (N_4983,In_2700,In_2533);
xor U4984 (N_4984,In_2408,In_1947);
nand U4985 (N_4985,In_620,In_340);
nor U4986 (N_4986,In_1552,In_2912);
or U4987 (N_4987,In_657,In_1629);
nand U4988 (N_4988,In_2076,In_2005);
xor U4989 (N_4989,In_1167,In_774);
xnor U4990 (N_4990,In_2692,In_1645);
nand U4991 (N_4991,In_913,In_2534);
nor U4992 (N_4992,In_1386,In_2220);
nor U4993 (N_4993,In_2631,In_2661);
and U4994 (N_4994,In_2832,In_1064);
and U4995 (N_4995,In_1583,In_444);
or U4996 (N_4996,In_267,In_62);
xnor U4997 (N_4997,In_2955,In_1605);
and U4998 (N_4998,In_1187,In_928);
nand U4999 (N_4999,In_184,In_853);
and U5000 (N_5000,In_483,In_661);
nand U5001 (N_5001,In_2644,In_573);
or U5002 (N_5002,In_1472,In_288);
nand U5003 (N_5003,In_653,In_2637);
nand U5004 (N_5004,In_2266,In_30);
or U5005 (N_5005,In_2833,In_792);
and U5006 (N_5006,In_2224,In_910);
or U5007 (N_5007,In_696,In_661);
or U5008 (N_5008,In_1351,In_2247);
nand U5009 (N_5009,In_2270,In_1633);
or U5010 (N_5010,In_2468,In_2152);
xnor U5011 (N_5011,In_2340,In_2171);
nor U5012 (N_5012,In_400,In_2445);
nor U5013 (N_5013,In_93,In_305);
or U5014 (N_5014,In_1612,In_166);
or U5015 (N_5015,In_345,In_2104);
or U5016 (N_5016,In_2022,In_2798);
xor U5017 (N_5017,In_2758,In_830);
or U5018 (N_5018,In_1878,In_1980);
and U5019 (N_5019,In_0,In_1785);
or U5020 (N_5020,In_403,In_626);
or U5021 (N_5021,In_216,In_1683);
and U5022 (N_5022,In_2012,In_622);
and U5023 (N_5023,In_1021,In_700);
and U5024 (N_5024,In_2564,In_1770);
nand U5025 (N_5025,In_1187,In_1584);
and U5026 (N_5026,In_2577,In_730);
or U5027 (N_5027,In_2292,In_77);
nand U5028 (N_5028,In_204,In_166);
xor U5029 (N_5029,In_2669,In_174);
nand U5030 (N_5030,In_2045,In_102);
nand U5031 (N_5031,In_1768,In_2115);
nand U5032 (N_5032,In_412,In_428);
nand U5033 (N_5033,In_1214,In_1230);
xor U5034 (N_5034,In_2054,In_1248);
or U5035 (N_5035,In_2736,In_1646);
nand U5036 (N_5036,In_1097,In_2134);
nand U5037 (N_5037,In_1443,In_2274);
and U5038 (N_5038,In_1509,In_1408);
nor U5039 (N_5039,In_1156,In_2797);
nor U5040 (N_5040,In_2350,In_1330);
or U5041 (N_5041,In_1068,In_1780);
xor U5042 (N_5042,In_1665,In_1891);
or U5043 (N_5043,In_2292,In_1779);
and U5044 (N_5044,In_2601,In_374);
nand U5045 (N_5045,In_2860,In_2597);
xor U5046 (N_5046,In_1537,In_794);
nand U5047 (N_5047,In_1595,In_277);
or U5048 (N_5048,In_1898,In_527);
xnor U5049 (N_5049,In_1958,In_1378);
xnor U5050 (N_5050,In_2384,In_2992);
or U5051 (N_5051,In_2092,In_1681);
nand U5052 (N_5052,In_708,In_157);
or U5053 (N_5053,In_986,In_996);
nand U5054 (N_5054,In_1411,In_1364);
or U5055 (N_5055,In_1227,In_2494);
and U5056 (N_5056,In_5,In_1952);
xor U5057 (N_5057,In_2752,In_1421);
xnor U5058 (N_5058,In_1903,In_13);
and U5059 (N_5059,In_1700,In_2053);
xnor U5060 (N_5060,In_274,In_1187);
nand U5061 (N_5061,In_716,In_43);
or U5062 (N_5062,In_1975,In_626);
nand U5063 (N_5063,In_2917,In_2525);
and U5064 (N_5064,In_370,In_245);
nand U5065 (N_5065,In_2097,In_1996);
and U5066 (N_5066,In_392,In_2603);
nor U5067 (N_5067,In_745,In_1499);
and U5068 (N_5068,In_1374,In_2868);
or U5069 (N_5069,In_2640,In_2822);
or U5070 (N_5070,In_2501,In_703);
nand U5071 (N_5071,In_518,In_1774);
and U5072 (N_5072,In_1958,In_2158);
nor U5073 (N_5073,In_2739,In_2646);
xnor U5074 (N_5074,In_704,In_965);
or U5075 (N_5075,In_1770,In_826);
nor U5076 (N_5076,In_2203,In_578);
nand U5077 (N_5077,In_2497,In_229);
nor U5078 (N_5078,In_2859,In_2841);
xor U5079 (N_5079,In_1686,In_2033);
xor U5080 (N_5080,In_1382,In_411);
xnor U5081 (N_5081,In_687,In_2592);
xor U5082 (N_5082,In_2473,In_676);
and U5083 (N_5083,In_1749,In_1184);
nand U5084 (N_5084,In_690,In_2677);
or U5085 (N_5085,In_1527,In_1802);
or U5086 (N_5086,In_480,In_2495);
xor U5087 (N_5087,In_1838,In_38);
and U5088 (N_5088,In_2189,In_1870);
nand U5089 (N_5089,In_422,In_1098);
nand U5090 (N_5090,In_2804,In_2702);
nor U5091 (N_5091,In_156,In_2213);
nor U5092 (N_5092,In_2177,In_134);
nand U5093 (N_5093,In_2672,In_1059);
and U5094 (N_5094,In_1631,In_1814);
nand U5095 (N_5095,In_929,In_2842);
nor U5096 (N_5096,In_1691,In_1390);
and U5097 (N_5097,In_53,In_296);
nor U5098 (N_5098,In_2661,In_881);
and U5099 (N_5099,In_1781,In_1039);
xnor U5100 (N_5100,In_1991,In_1487);
or U5101 (N_5101,In_1505,In_752);
nand U5102 (N_5102,In_2079,In_2014);
xnor U5103 (N_5103,In_1132,In_2828);
nand U5104 (N_5104,In_2881,In_2131);
and U5105 (N_5105,In_1969,In_1838);
nor U5106 (N_5106,In_2731,In_1549);
or U5107 (N_5107,In_561,In_1065);
xor U5108 (N_5108,In_1279,In_2727);
nor U5109 (N_5109,In_1123,In_180);
nor U5110 (N_5110,In_1320,In_915);
nor U5111 (N_5111,In_2251,In_2996);
nor U5112 (N_5112,In_620,In_770);
and U5113 (N_5113,In_677,In_1727);
xnor U5114 (N_5114,In_1510,In_2149);
and U5115 (N_5115,In_2005,In_2209);
nand U5116 (N_5116,In_1271,In_293);
nor U5117 (N_5117,In_2876,In_140);
nand U5118 (N_5118,In_79,In_2517);
xor U5119 (N_5119,In_2658,In_232);
nor U5120 (N_5120,In_1385,In_1535);
nor U5121 (N_5121,In_86,In_2699);
nand U5122 (N_5122,In_958,In_529);
or U5123 (N_5123,In_823,In_2665);
nand U5124 (N_5124,In_2848,In_2048);
or U5125 (N_5125,In_2815,In_1187);
or U5126 (N_5126,In_1439,In_305);
or U5127 (N_5127,In_856,In_2256);
nor U5128 (N_5128,In_267,In_2530);
or U5129 (N_5129,In_1095,In_1619);
xnor U5130 (N_5130,In_1233,In_984);
nand U5131 (N_5131,In_432,In_2075);
nor U5132 (N_5132,In_18,In_2416);
or U5133 (N_5133,In_2148,In_1217);
or U5134 (N_5134,In_2945,In_917);
or U5135 (N_5135,In_618,In_2084);
nand U5136 (N_5136,In_2075,In_1988);
nand U5137 (N_5137,In_2935,In_2954);
nand U5138 (N_5138,In_616,In_2294);
nand U5139 (N_5139,In_1831,In_2596);
or U5140 (N_5140,In_2437,In_771);
and U5141 (N_5141,In_1734,In_214);
or U5142 (N_5142,In_2363,In_1831);
xnor U5143 (N_5143,In_700,In_1041);
xnor U5144 (N_5144,In_1342,In_578);
xnor U5145 (N_5145,In_468,In_1701);
or U5146 (N_5146,In_2555,In_741);
nor U5147 (N_5147,In_1930,In_254);
nand U5148 (N_5148,In_1112,In_392);
or U5149 (N_5149,In_1178,In_1034);
xnor U5150 (N_5150,In_510,In_668);
and U5151 (N_5151,In_255,In_187);
xnor U5152 (N_5152,In_2076,In_1634);
nand U5153 (N_5153,In_2020,In_1835);
or U5154 (N_5154,In_2802,In_1764);
nor U5155 (N_5155,In_816,In_93);
and U5156 (N_5156,In_1382,In_2334);
and U5157 (N_5157,In_415,In_1101);
or U5158 (N_5158,In_300,In_1725);
nor U5159 (N_5159,In_1788,In_291);
or U5160 (N_5160,In_2642,In_473);
and U5161 (N_5161,In_1668,In_1643);
or U5162 (N_5162,In_1464,In_2372);
nand U5163 (N_5163,In_2082,In_900);
xor U5164 (N_5164,In_417,In_2653);
nor U5165 (N_5165,In_2493,In_2009);
nand U5166 (N_5166,In_1244,In_2939);
xor U5167 (N_5167,In_2020,In_1107);
and U5168 (N_5168,In_1552,In_327);
and U5169 (N_5169,In_716,In_1437);
nand U5170 (N_5170,In_2252,In_1939);
and U5171 (N_5171,In_803,In_2727);
nor U5172 (N_5172,In_530,In_2273);
nand U5173 (N_5173,In_92,In_716);
and U5174 (N_5174,In_2497,In_1245);
and U5175 (N_5175,In_1522,In_1643);
nand U5176 (N_5176,In_1327,In_2343);
nor U5177 (N_5177,In_428,In_789);
or U5178 (N_5178,In_2905,In_2284);
or U5179 (N_5179,In_2357,In_659);
xnor U5180 (N_5180,In_2400,In_2536);
and U5181 (N_5181,In_1274,In_656);
and U5182 (N_5182,In_2157,In_1402);
or U5183 (N_5183,In_1310,In_1317);
nand U5184 (N_5184,In_1544,In_1785);
nand U5185 (N_5185,In_796,In_2811);
or U5186 (N_5186,In_2666,In_244);
and U5187 (N_5187,In_1492,In_694);
nand U5188 (N_5188,In_2212,In_1055);
nor U5189 (N_5189,In_250,In_2852);
or U5190 (N_5190,In_1117,In_1366);
nor U5191 (N_5191,In_1100,In_443);
or U5192 (N_5192,In_909,In_324);
xor U5193 (N_5193,In_420,In_768);
or U5194 (N_5194,In_1852,In_1008);
nand U5195 (N_5195,In_2801,In_2682);
nand U5196 (N_5196,In_791,In_1800);
and U5197 (N_5197,In_1542,In_2988);
xor U5198 (N_5198,In_590,In_1026);
nand U5199 (N_5199,In_2300,In_973);
nand U5200 (N_5200,In_901,In_1118);
or U5201 (N_5201,In_1160,In_1588);
xor U5202 (N_5202,In_511,In_2138);
xor U5203 (N_5203,In_2290,In_2489);
nor U5204 (N_5204,In_2500,In_71);
xor U5205 (N_5205,In_2044,In_1187);
xor U5206 (N_5206,In_2838,In_2526);
nor U5207 (N_5207,In_1179,In_1823);
nand U5208 (N_5208,In_2897,In_1400);
nor U5209 (N_5209,In_982,In_276);
and U5210 (N_5210,In_1298,In_9);
nand U5211 (N_5211,In_338,In_810);
and U5212 (N_5212,In_915,In_963);
or U5213 (N_5213,In_2309,In_555);
xor U5214 (N_5214,In_2120,In_1581);
nor U5215 (N_5215,In_1010,In_44);
or U5216 (N_5216,In_1851,In_913);
nor U5217 (N_5217,In_1512,In_440);
nand U5218 (N_5218,In_812,In_618);
or U5219 (N_5219,In_749,In_1539);
or U5220 (N_5220,In_2463,In_2695);
nand U5221 (N_5221,In_1148,In_1603);
or U5222 (N_5222,In_2789,In_2825);
nand U5223 (N_5223,In_2116,In_907);
nor U5224 (N_5224,In_764,In_881);
xnor U5225 (N_5225,In_720,In_315);
nand U5226 (N_5226,In_2933,In_1239);
nand U5227 (N_5227,In_894,In_2296);
nor U5228 (N_5228,In_1738,In_2575);
nor U5229 (N_5229,In_1441,In_1012);
and U5230 (N_5230,In_987,In_373);
or U5231 (N_5231,In_2530,In_650);
or U5232 (N_5232,In_1468,In_1533);
nand U5233 (N_5233,In_587,In_1638);
nor U5234 (N_5234,In_1629,In_442);
xnor U5235 (N_5235,In_2138,In_1659);
or U5236 (N_5236,In_1520,In_2965);
or U5237 (N_5237,In_528,In_54);
xor U5238 (N_5238,In_1081,In_1008);
and U5239 (N_5239,In_392,In_124);
or U5240 (N_5240,In_2871,In_617);
xor U5241 (N_5241,In_686,In_1932);
xor U5242 (N_5242,In_1247,In_1832);
xnor U5243 (N_5243,In_1145,In_2526);
nand U5244 (N_5244,In_1964,In_86);
and U5245 (N_5245,In_49,In_1061);
and U5246 (N_5246,In_97,In_2211);
or U5247 (N_5247,In_604,In_1395);
nand U5248 (N_5248,In_593,In_702);
nor U5249 (N_5249,In_1313,In_251);
xnor U5250 (N_5250,In_259,In_1966);
and U5251 (N_5251,In_2974,In_1251);
and U5252 (N_5252,In_981,In_893);
xor U5253 (N_5253,In_256,In_2063);
nand U5254 (N_5254,In_40,In_1946);
nor U5255 (N_5255,In_1818,In_2967);
xnor U5256 (N_5256,In_1278,In_101);
nand U5257 (N_5257,In_393,In_799);
and U5258 (N_5258,In_1974,In_1731);
nand U5259 (N_5259,In_2512,In_803);
nor U5260 (N_5260,In_2327,In_1060);
xor U5261 (N_5261,In_1387,In_1674);
xnor U5262 (N_5262,In_2683,In_1651);
nand U5263 (N_5263,In_2602,In_1860);
or U5264 (N_5264,In_580,In_1675);
or U5265 (N_5265,In_107,In_1254);
nand U5266 (N_5266,In_469,In_297);
nand U5267 (N_5267,In_1502,In_929);
nand U5268 (N_5268,In_1849,In_1824);
nor U5269 (N_5269,In_269,In_224);
nand U5270 (N_5270,In_2709,In_236);
nor U5271 (N_5271,In_1353,In_2385);
or U5272 (N_5272,In_557,In_168);
xor U5273 (N_5273,In_1040,In_1606);
or U5274 (N_5274,In_2367,In_1063);
nand U5275 (N_5275,In_1946,In_576);
or U5276 (N_5276,In_1068,In_499);
xor U5277 (N_5277,In_1064,In_148);
xnor U5278 (N_5278,In_2858,In_68);
xnor U5279 (N_5279,In_2177,In_2626);
or U5280 (N_5280,In_2779,In_127);
or U5281 (N_5281,In_468,In_1009);
nand U5282 (N_5282,In_1259,In_1375);
or U5283 (N_5283,In_2636,In_2553);
nor U5284 (N_5284,In_579,In_123);
nor U5285 (N_5285,In_1361,In_1328);
nor U5286 (N_5286,In_367,In_2389);
xnor U5287 (N_5287,In_1018,In_2238);
and U5288 (N_5288,In_309,In_2276);
nor U5289 (N_5289,In_515,In_414);
xor U5290 (N_5290,In_1038,In_2791);
xnor U5291 (N_5291,In_2472,In_2069);
nor U5292 (N_5292,In_411,In_493);
xor U5293 (N_5293,In_1237,In_1604);
or U5294 (N_5294,In_1803,In_2942);
xnor U5295 (N_5295,In_500,In_1360);
and U5296 (N_5296,In_800,In_2780);
xnor U5297 (N_5297,In_2027,In_2445);
and U5298 (N_5298,In_912,In_1717);
and U5299 (N_5299,In_285,In_183);
nor U5300 (N_5300,In_989,In_925);
or U5301 (N_5301,In_31,In_642);
or U5302 (N_5302,In_772,In_744);
or U5303 (N_5303,In_1336,In_351);
xor U5304 (N_5304,In_2772,In_745);
and U5305 (N_5305,In_2463,In_1638);
and U5306 (N_5306,In_665,In_2222);
nand U5307 (N_5307,In_996,In_2311);
nor U5308 (N_5308,In_1039,In_2787);
nor U5309 (N_5309,In_2540,In_185);
and U5310 (N_5310,In_2157,In_2362);
and U5311 (N_5311,In_767,In_1082);
and U5312 (N_5312,In_2315,In_1532);
xnor U5313 (N_5313,In_2777,In_841);
xor U5314 (N_5314,In_2221,In_1138);
nand U5315 (N_5315,In_1076,In_1274);
and U5316 (N_5316,In_723,In_389);
xnor U5317 (N_5317,In_102,In_809);
nand U5318 (N_5318,In_2141,In_1790);
nand U5319 (N_5319,In_209,In_284);
and U5320 (N_5320,In_805,In_439);
xnor U5321 (N_5321,In_1541,In_2975);
or U5322 (N_5322,In_182,In_2619);
nand U5323 (N_5323,In_2584,In_2945);
and U5324 (N_5324,In_718,In_1434);
or U5325 (N_5325,In_1021,In_758);
or U5326 (N_5326,In_2418,In_2303);
nor U5327 (N_5327,In_2967,In_2620);
or U5328 (N_5328,In_1227,In_1491);
nand U5329 (N_5329,In_2943,In_1176);
xnor U5330 (N_5330,In_841,In_914);
and U5331 (N_5331,In_1071,In_1803);
and U5332 (N_5332,In_2856,In_410);
or U5333 (N_5333,In_1361,In_2711);
or U5334 (N_5334,In_374,In_2299);
or U5335 (N_5335,In_1891,In_2891);
nand U5336 (N_5336,In_423,In_2609);
nor U5337 (N_5337,In_1577,In_1434);
nand U5338 (N_5338,In_2428,In_578);
nor U5339 (N_5339,In_2659,In_1992);
or U5340 (N_5340,In_2483,In_2962);
nor U5341 (N_5341,In_1260,In_2279);
xnor U5342 (N_5342,In_1551,In_1499);
nor U5343 (N_5343,In_1817,In_1760);
nand U5344 (N_5344,In_1481,In_2628);
and U5345 (N_5345,In_1865,In_2810);
and U5346 (N_5346,In_2594,In_100);
nand U5347 (N_5347,In_1659,In_819);
or U5348 (N_5348,In_2977,In_2756);
nand U5349 (N_5349,In_1091,In_1821);
nand U5350 (N_5350,In_738,In_204);
xor U5351 (N_5351,In_1351,In_1747);
nor U5352 (N_5352,In_1616,In_1492);
nand U5353 (N_5353,In_2126,In_255);
nand U5354 (N_5354,In_1624,In_391);
xnor U5355 (N_5355,In_658,In_417);
nor U5356 (N_5356,In_1917,In_1579);
xnor U5357 (N_5357,In_2386,In_2975);
nand U5358 (N_5358,In_73,In_2931);
xnor U5359 (N_5359,In_1577,In_1024);
nand U5360 (N_5360,In_1427,In_2903);
xor U5361 (N_5361,In_2624,In_792);
and U5362 (N_5362,In_1702,In_2671);
nand U5363 (N_5363,In_2600,In_329);
nor U5364 (N_5364,In_999,In_2724);
and U5365 (N_5365,In_2831,In_1503);
xnor U5366 (N_5366,In_1858,In_1273);
xnor U5367 (N_5367,In_1051,In_2595);
nand U5368 (N_5368,In_2897,In_148);
nor U5369 (N_5369,In_6,In_2439);
and U5370 (N_5370,In_142,In_1492);
nand U5371 (N_5371,In_611,In_394);
nand U5372 (N_5372,In_477,In_236);
xnor U5373 (N_5373,In_2339,In_2749);
nor U5374 (N_5374,In_1953,In_2962);
xnor U5375 (N_5375,In_1490,In_2329);
nor U5376 (N_5376,In_1264,In_1021);
xor U5377 (N_5377,In_1085,In_1346);
or U5378 (N_5378,In_1110,In_1468);
nor U5379 (N_5379,In_2530,In_97);
and U5380 (N_5380,In_61,In_562);
xnor U5381 (N_5381,In_1275,In_2609);
or U5382 (N_5382,In_341,In_1613);
or U5383 (N_5383,In_1922,In_924);
xnor U5384 (N_5384,In_1014,In_1741);
or U5385 (N_5385,In_152,In_138);
nor U5386 (N_5386,In_216,In_2274);
nor U5387 (N_5387,In_2006,In_2501);
nor U5388 (N_5388,In_2535,In_946);
nor U5389 (N_5389,In_2456,In_2039);
or U5390 (N_5390,In_687,In_1442);
and U5391 (N_5391,In_307,In_2553);
nor U5392 (N_5392,In_1494,In_2684);
nand U5393 (N_5393,In_2212,In_686);
xor U5394 (N_5394,In_1630,In_1858);
and U5395 (N_5395,In_275,In_1930);
nor U5396 (N_5396,In_2338,In_2446);
or U5397 (N_5397,In_151,In_2254);
nor U5398 (N_5398,In_2799,In_714);
nor U5399 (N_5399,In_690,In_1432);
nand U5400 (N_5400,In_577,In_148);
nor U5401 (N_5401,In_2580,In_2374);
and U5402 (N_5402,In_1504,In_1203);
nor U5403 (N_5403,In_502,In_1026);
or U5404 (N_5404,In_2104,In_276);
nand U5405 (N_5405,In_1988,In_2591);
nor U5406 (N_5406,In_1799,In_1013);
nand U5407 (N_5407,In_2944,In_3);
xor U5408 (N_5408,In_2772,In_2476);
nand U5409 (N_5409,In_1903,In_2968);
xnor U5410 (N_5410,In_1462,In_1000);
nor U5411 (N_5411,In_1772,In_2343);
nand U5412 (N_5412,In_2777,In_2304);
and U5413 (N_5413,In_1380,In_2633);
nor U5414 (N_5414,In_299,In_1263);
xnor U5415 (N_5415,In_2114,In_2694);
nand U5416 (N_5416,In_870,In_335);
nor U5417 (N_5417,In_1916,In_755);
nand U5418 (N_5418,In_1066,In_142);
nand U5419 (N_5419,In_2603,In_108);
nor U5420 (N_5420,In_1930,In_415);
nand U5421 (N_5421,In_2368,In_1094);
nand U5422 (N_5422,In_2572,In_2939);
xnor U5423 (N_5423,In_1710,In_1094);
and U5424 (N_5424,In_2672,In_2593);
and U5425 (N_5425,In_2070,In_2208);
and U5426 (N_5426,In_1787,In_2727);
nor U5427 (N_5427,In_2633,In_402);
or U5428 (N_5428,In_897,In_2767);
xor U5429 (N_5429,In_944,In_432);
nor U5430 (N_5430,In_1249,In_2420);
and U5431 (N_5431,In_841,In_2301);
nor U5432 (N_5432,In_2606,In_851);
xnor U5433 (N_5433,In_2875,In_894);
nor U5434 (N_5434,In_2439,In_2326);
nand U5435 (N_5435,In_1672,In_1940);
or U5436 (N_5436,In_1394,In_947);
nor U5437 (N_5437,In_693,In_1028);
or U5438 (N_5438,In_1936,In_2540);
xor U5439 (N_5439,In_1927,In_790);
xnor U5440 (N_5440,In_158,In_738);
or U5441 (N_5441,In_2971,In_2972);
and U5442 (N_5442,In_2339,In_1190);
nand U5443 (N_5443,In_1989,In_2653);
or U5444 (N_5444,In_2778,In_2356);
nand U5445 (N_5445,In_2441,In_2151);
nor U5446 (N_5446,In_1256,In_2939);
nor U5447 (N_5447,In_2457,In_1765);
xnor U5448 (N_5448,In_1044,In_2273);
nand U5449 (N_5449,In_1323,In_1525);
and U5450 (N_5450,In_738,In_1197);
or U5451 (N_5451,In_615,In_1485);
nor U5452 (N_5452,In_783,In_2173);
nor U5453 (N_5453,In_1119,In_2644);
and U5454 (N_5454,In_981,In_2087);
nand U5455 (N_5455,In_2294,In_179);
nand U5456 (N_5456,In_2433,In_457);
nand U5457 (N_5457,In_2080,In_1445);
nand U5458 (N_5458,In_1038,In_559);
nand U5459 (N_5459,In_2469,In_1102);
nand U5460 (N_5460,In_2378,In_1725);
and U5461 (N_5461,In_2992,In_1422);
xor U5462 (N_5462,In_724,In_190);
or U5463 (N_5463,In_581,In_2473);
xor U5464 (N_5464,In_1272,In_102);
nor U5465 (N_5465,In_1617,In_1641);
or U5466 (N_5466,In_2536,In_2360);
nand U5467 (N_5467,In_673,In_2114);
and U5468 (N_5468,In_2117,In_1947);
nand U5469 (N_5469,In_2978,In_765);
nand U5470 (N_5470,In_635,In_2700);
or U5471 (N_5471,In_2064,In_1226);
nand U5472 (N_5472,In_1183,In_1031);
and U5473 (N_5473,In_2115,In_502);
or U5474 (N_5474,In_508,In_2923);
or U5475 (N_5475,In_1115,In_124);
nor U5476 (N_5476,In_44,In_2404);
nand U5477 (N_5477,In_228,In_2061);
or U5478 (N_5478,In_1744,In_158);
and U5479 (N_5479,In_2100,In_1722);
nand U5480 (N_5480,In_1222,In_2542);
or U5481 (N_5481,In_1376,In_1640);
nor U5482 (N_5482,In_1759,In_726);
nand U5483 (N_5483,In_324,In_536);
xnor U5484 (N_5484,In_2988,In_352);
and U5485 (N_5485,In_2941,In_65);
and U5486 (N_5486,In_2760,In_115);
and U5487 (N_5487,In_2916,In_1323);
xnor U5488 (N_5488,In_118,In_2123);
or U5489 (N_5489,In_1908,In_182);
xor U5490 (N_5490,In_1576,In_1370);
xnor U5491 (N_5491,In_1317,In_454);
nand U5492 (N_5492,In_2544,In_2527);
xor U5493 (N_5493,In_2983,In_1904);
and U5494 (N_5494,In_2548,In_2919);
and U5495 (N_5495,In_2298,In_223);
xor U5496 (N_5496,In_2080,In_2564);
or U5497 (N_5497,In_1499,In_526);
xnor U5498 (N_5498,In_2916,In_211);
and U5499 (N_5499,In_904,In_885);
xnor U5500 (N_5500,In_1612,In_2040);
and U5501 (N_5501,In_2834,In_1033);
or U5502 (N_5502,In_1600,In_1862);
xor U5503 (N_5503,In_2375,In_762);
xnor U5504 (N_5504,In_240,In_486);
and U5505 (N_5505,In_1390,In_371);
or U5506 (N_5506,In_179,In_2431);
and U5507 (N_5507,In_1759,In_57);
or U5508 (N_5508,In_1057,In_1458);
and U5509 (N_5509,In_486,In_1372);
xnor U5510 (N_5510,In_1012,In_2141);
nand U5511 (N_5511,In_928,In_1893);
and U5512 (N_5512,In_1217,In_2210);
nor U5513 (N_5513,In_111,In_792);
xnor U5514 (N_5514,In_935,In_787);
nand U5515 (N_5515,In_2061,In_2161);
or U5516 (N_5516,In_2733,In_230);
nor U5517 (N_5517,In_2401,In_2077);
or U5518 (N_5518,In_1257,In_2819);
or U5519 (N_5519,In_1253,In_1670);
or U5520 (N_5520,In_683,In_2455);
xnor U5521 (N_5521,In_2491,In_123);
or U5522 (N_5522,In_2224,In_2522);
nor U5523 (N_5523,In_1215,In_247);
xnor U5524 (N_5524,In_256,In_412);
or U5525 (N_5525,In_1088,In_610);
nor U5526 (N_5526,In_2022,In_1904);
and U5527 (N_5527,In_953,In_13);
or U5528 (N_5528,In_1480,In_1875);
nor U5529 (N_5529,In_1414,In_448);
or U5530 (N_5530,In_2714,In_231);
or U5531 (N_5531,In_1703,In_2428);
and U5532 (N_5532,In_454,In_1024);
nor U5533 (N_5533,In_804,In_1092);
and U5534 (N_5534,In_476,In_709);
nor U5535 (N_5535,In_816,In_667);
nor U5536 (N_5536,In_2712,In_647);
or U5537 (N_5537,In_2511,In_1612);
nand U5538 (N_5538,In_716,In_2917);
nor U5539 (N_5539,In_1651,In_1536);
nor U5540 (N_5540,In_1437,In_244);
xor U5541 (N_5541,In_1534,In_2260);
xnor U5542 (N_5542,In_831,In_764);
or U5543 (N_5543,In_1208,In_1342);
xnor U5544 (N_5544,In_1408,In_2130);
xor U5545 (N_5545,In_491,In_2653);
nand U5546 (N_5546,In_465,In_1211);
and U5547 (N_5547,In_513,In_207);
or U5548 (N_5548,In_2905,In_581);
nor U5549 (N_5549,In_2035,In_1199);
xor U5550 (N_5550,In_2963,In_1620);
xnor U5551 (N_5551,In_633,In_2170);
or U5552 (N_5552,In_43,In_1054);
xnor U5553 (N_5553,In_666,In_311);
or U5554 (N_5554,In_1791,In_227);
xnor U5555 (N_5555,In_2076,In_1733);
nor U5556 (N_5556,In_1689,In_859);
nor U5557 (N_5557,In_2428,In_1191);
nand U5558 (N_5558,In_1355,In_2636);
xor U5559 (N_5559,In_1398,In_2784);
and U5560 (N_5560,In_56,In_1207);
xnor U5561 (N_5561,In_2390,In_504);
or U5562 (N_5562,In_1343,In_516);
nand U5563 (N_5563,In_1439,In_132);
and U5564 (N_5564,In_2995,In_117);
nor U5565 (N_5565,In_2601,In_1998);
or U5566 (N_5566,In_29,In_317);
and U5567 (N_5567,In_189,In_2571);
nor U5568 (N_5568,In_940,In_1476);
nor U5569 (N_5569,In_1927,In_2064);
or U5570 (N_5570,In_1160,In_1007);
nand U5571 (N_5571,In_157,In_911);
and U5572 (N_5572,In_2611,In_1009);
and U5573 (N_5573,In_2239,In_1372);
nor U5574 (N_5574,In_1128,In_1722);
or U5575 (N_5575,In_278,In_2430);
or U5576 (N_5576,In_1117,In_1572);
or U5577 (N_5577,In_2431,In_2916);
nand U5578 (N_5578,In_1876,In_433);
or U5579 (N_5579,In_276,In_1045);
or U5580 (N_5580,In_609,In_2134);
nand U5581 (N_5581,In_1451,In_1466);
and U5582 (N_5582,In_1702,In_873);
or U5583 (N_5583,In_1113,In_2550);
nand U5584 (N_5584,In_1856,In_647);
and U5585 (N_5585,In_408,In_2797);
or U5586 (N_5586,In_1690,In_2910);
or U5587 (N_5587,In_644,In_482);
or U5588 (N_5588,In_2547,In_1220);
nor U5589 (N_5589,In_2458,In_471);
and U5590 (N_5590,In_1685,In_2621);
nor U5591 (N_5591,In_1356,In_323);
nor U5592 (N_5592,In_2528,In_1591);
and U5593 (N_5593,In_1771,In_181);
or U5594 (N_5594,In_2514,In_2804);
or U5595 (N_5595,In_569,In_212);
nor U5596 (N_5596,In_287,In_1678);
nor U5597 (N_5597,In_1301,In_2491);
and U5598 (N_5598,In_367,In_328);
or U5599 (N_5599,In_646,In_1226);
xnor U5600 (N_5600,In_67,In_1248);
or U5601 (N_5601,In_2537,In_424);
nand U5602 (N_5602,In_1488,In_95);
nand U5603 (N_5603,In_77,In_517);
nand U5604 (N_5604,In_2403,In_1460);
nand U5605 (N_5605,In_473,In_982);
xor U5606 (N_5606,In_786,In_2052);
nand U5607 (N_5607,In_613,In_687);
nor U5608 (N_5608,In_312,In_2530);
nor U5609 (N_5609,In_1648,In_2231);
nor U5610 (N_5610,In_537,In_1805);
nor U5611 (N_5611,In_410,In_961);
nand U5612 (N_5612,In_2211,In_587);
nand U5613 (N_5613,In_819,In_2781);
xnor U5614 (N_5614,In_1726,In_1738);
nor U5615 (N_5615,In_1439,In_2688);
nand U5616 (N_5616,In_2422,In_642);
or U5617 (N_5617,In_2777,In_452);
nand U5618 (N_5618,In_380,In_1160);
and U5619 (N_5619,In_2542,In_1633);
or U5620 (N_5620,In_1481,In_777);
xor U5621 (N_5621,In_1450,In_1553);
nor U5622 (N_5622,In_1217,In_512);
xnor U5623 (N_5623,In_1547,In_766);
nand U5624 (N_5624,In_455,In_1721);
nand U5625 (N_5625,In_1203,In_2802);
or U5626 (N_5626,In_2130,In_804);
nor U5627 (N_5627,In_1443,In_441);
nor U5628 (N_5628,In_1132,In_2565);
or U5629 (N_5629,In_527,In_98);
xnor U5630 (N_5630,In_761,In_1819);
and U5631 (N_5631,In_147,In_886);
and U5632 (N_5632,In_1938,In_2342);
or U5633 (N_5633,In_966,In_294);
nand U5634 (N_5634,In_2221,In_1364);
xnor U5635 (N_5635,In_84,In_721);
xnor U5636 (N_5636,In_427,In_2354);
nor U5637 (N_5637,In_1884,In_1431);
nor U5638 (N_5638,In_2740,In_2867);
nor U5639 (N_5639,In_2583,In_1620);
nand U5640 (N_5640,In_1678,In_2904);
and U5641 (N_5641,In_1392,In_2514);
nor U5642 (N_5642,In_286,In_1489);
xnor U5643 (N_5643,In_2529,In_835);
nand U5644 (N_5644,In_2234,In_2057);
and U5645 (N_5645,In_1185,In_1731);
xnor U5646 (N_5646,In_605,In_159);
nand U5647 (N_5647,In_498,In_1864);
and U5648 (N_5648,In_18,In_2971);
xnor U5649 (N_5649,In_378,In_1844);
nor U5650 (N_5650,In_2163,In_1631);
nor U5651 (N_5651,In_495,In_2298);
nor U5652 (N_5652,In_790,In_1694);
and U5653 (N_5653,In_877,In_1842);
xnor U5654 (N_5654,In_1892,In_152);
and U5655 (N_5655,In_233,In_1787);
xor U5656 (N_5656,In_1303,In_1498);
and U5657 (N_5657,In_2610,In_96);
nor U5658 (N_5658,In_2566,In_1191);
and U5659 (N_5659,In_2559,In_1907);
nand U5660 (N_5660,In_613,In_2226);
or U5661 (N_5661,In_1397,In_410);
or U5662 (N_5662,In_678,In_1879);
xnor U5663 (N_5663,In_2074,In_489);
nor U5664 (N_5664,In_2100,In_2206);
nand U5665 (N_5665,In_1327,In_572);
xnor U5666 (N_5666,In_1341,In_1503);
or U5667 (N_5667,In_45,In_2634);
nand U5668 (N_5668,In_2324,In_1994);
and U5669 (N_5669,In_2201,In_2336);
and U5670 (N_5670,In_778,In_32);
and U5671 (N_5671,In_242,In_748);
or U5672 (N_5672,In_109,In_146);
nand U5673 (N_5673,In_490,In_453);
xor U5674 (N_5674,In_2303,In_668);
nor U5675 (N_5675,In_1105,In_2117);
or U5676 (N_5676,In_2796,In_22);
and U5677 (N_5677,In_811,In_670);
nor U5678 (N_5678,In_2890,In_1803);
or U5679 (N_5679,In_2736,In_2193);
nand U5680 (N_5680,In_2523,In_2051);
nand U5681 (N_5681,In_2275,In_1991);
xor U5682 (N_5682,In_514,In_2399);
nand U5683 (N_5683,In_913,In_890);
nand U5684 (N_5684,In_2980,In_1950);
and U5685 (N_5685,In_1430,In_2964);
nand U5686 (N_5686,In_921,In_2703);
nand U5687 (N_5687,In_1527,In_588);
nor U5688 (N_5688,In_1472,In_1815);
or U5689 (N_5689,In_478,In_1355);
or U5690 (N_5690,In_1582,In_1855);
nand U5691 (N_5691,In_2233,In_2927);
or U5692 (N_5692,In_1528,In_108);
nor U5693 (N_5693,In_325,In_583);
nand U5694 (N_5694,In_35,In_1650);
and U5695 (N_5695,In_1486,In_1999);
or U5696 (N_5696,In_2550,In_2103);
and U5697 (N_5697,In_634,In_1162);
nand U5698 (N_5698,In_2958,In_355);
and U5699 (N_5699,In_1947,In_820);
or U5700 (N_5700,In_2323,In_561);
xnor U5701 (N_5701,In_1972,In_1874);
nor U5702 (N_5702,In_2525,In_505);
xnor U5703 (N_5703,In_626,In_1112);
nor U5704 (N_5704,In_1178,In_2082);
and U5705 (N_5705,In_1383,In_180);
or U5706 (N_5706,In_391,In_795);
xor U5707 (N_5707,In_1220,In_2864);
or U5708 (N_5708,In_2816,In_709);
or U5709 (N_5709,In_1344,In_1379);
nand U5710 (N_5710,In_1453,In_2618);
nand U5711 (N_5711,In_832,In_614);
or U5712 (N_5712,In_329,In_1684);
and U5713 (N_5713,In_1806,In_1978);
xor U5714 (N_5714,In_2776,In_1297);
nor U5715 (N_5715,In_1981,In_250);
and U5716 (N_5716,In_2220,In_1667);
nor U5717 (N_5717,In_2736,In_219);
xor U5718 (N_5718,In_2145,In_2850);
nand U5719 (N_5719,In_1267,In_721);
xnor U5720 (N_5720,In_1940,In_2226);
nor U5721 (N_5721,In_2452,In_2646);
nand U5722 (N_5722,In_408,In_716);
and U5723 (N_5723,In_2227,In_888);
or U5724 (N_5724,In_1372,In_2904);
nor U5725 (N_5725,In_143,In_1665);
and U5726 (N_5726,In_2377,In_2689);
xnor U5727 (N_5727,In_2002,In_855);
and U5728 (N_5728,In_218,In_2012);
xnor U5729 (N_5729,In_2452,In_1579);
xor U5730 (N_5730,In_385,In_1139);
and U5731 (N_5731,In_2107,In_2183);
or U5732 (N_5732,In_2722,In_698);
nor U5733 (N_5733,In_1186,In_2785);
or U5734 (N_5734,In_2113,In_408);
or U5735 (N_5735,In_230,In_2558);
and U5736 (N_5736,In_210,In_1110);
and U5737 (N_5737,In_2607,In_2549);
xnor U5738 (N_5738,In_2675,In_264);
nor U5739 (N_5739,In_2566,In_1047);
nor U5740 (N_5740,In_1784,In_689);
and U5741 (N_5741,In_656,In_1566);
or U5742 (N_5742,In_2854,In_1129);
or U5743 (N_5743,In_1885,In_1866);
xor U5744 (N_5744,In_1842,In_260);
or U5745 (N_5745,In_2384,In_2886);
and U5746 (N_5746,In_2296,In_948);
and U5747 (N_5747,In_1233,In_1271);
or U5748 (N_5748,In_2111,In_287);
nor U5749 (N_5749,In_476,In_2811);
and U5750 (N_5750,In_515,In_2512);
nor U5751 (N_5751,In_308,In_1316);
xnor U5752 (N_5752,In_1082,In_79);
nand U5753 (N_5753,In_65,In_70);
or U5754 (N_5754,In_2736,In_1639);
xor U5755 (N_5755,In_1539,In_787);
or U5756 (N_5756,In_606,In_1283);
nand U5757 (N_5757,In_800,In_2257);
nor U5758 (N_5758,In_2138,In_1703);
nand U5759 (N_5759,In_2050,In_2666);
nand U5760 (N_5760,In_2049,In_1439);
and U5761 (N_5761,In_1474,In_355);
or U5762 (N_5762,In_423,In_2655);
nor U5763 (N_5763,In_2351,In_2061);
xor U5764 (N_5764,In_1708,In_1196);
or U5765 (N_5765,In_441,In_1258);
nand U5766 (N_5766,In_216,In_1960);
nand U5767 (N_5767,In_2511,In_1976);
xor U5768 (N_5768,In_963,In_506);
or U5769 (N_5769,In_1765,In_298);
or U5770 (N_5770,In_464,In_2368);
and U5771 (N_5771,In_2805,In_1415);
or U5772 (N_5772,In_1627,In_2622);
nand U5773 (N_5773,In_460,In_318);
nand U5774 (N_5774,In_2727,In_2096);
and U5775 (N_5775,In_91,In_2338);
and U5776 (N_5776,In_84,In_667);
or U5777 (N_5777,In_650,In_669);
nor U5778 (N_5778,In_394,In_2930);
nor U5779 (N_5779,In_2597,In_1347);
and U5780 (N_5780,In_282,In_778);
nand U5781 (N_5781,In_2913,In_2906);
nor U5782 (N_5782,In_800,In_126);
nand U5783 (N_5783,In_2626,In_81);
and U5784 (N_5784,In_1419,In_1561);
or U5785 (N_5785,In_1628,In_2898);
or U5786 (N_5786,In_1986,In_433);
xor U5787 (N_5787,In_1804,In_1347);
xor U5788 (N_5788,In_2752,In_2822);
xor U5789 (N_5789,In_24,In_1225);
xor U5790 (N_5790,In_2025,In_1636);
nand U5791 (N_5791,In_2568,In_1538);
xor U5792 (N_5792,In_2197,In_2946);
and U5793 (N_5793,In_361,In_2201);
or U5794 (N_5794,In_1009,In_1867);
or U5795 (N_5795,In_996,In_1791);
nand U5796 (N_5796,In_1214,In_1321);
nand U5797 (N_5797,In_809,In_2344);
nand U5798 (N_5798,In_2344,In_2668);
or U5799 (N_5799,In_951,In_231);
nand U5800 (N_5800,In_433,In_1310);
xor U5801 (N_5801,In_2814,In_1402);
and U5802 (N_5802,In_1537,In_515);
and U5803 (N_5803,In_2653,In_1625);
nand U5804 (N_5804,In_258,In_1989);
xor U5805 (N_5805,In_998,In_2336);
and U5806 (N_5806,In_2574,In_787);
nand U5807 (N_5807,In_2660,In_1478);
and U5808 (N_5808,In_1427,In_2418);
and U5809 (N_5809,In_2525,In_2488);
xnor U5810 (N_5810,In_980,In_355);
xor U5811 (N_5811,In_866,In_2075);
or U5812 (N_5812,In_2010,In_2462);
nand U5813 (N_5813,In_681,In_2166);
and U5814 (N_5814,In_1130,In_1098);
xor U5815 (N_5815,In_1010,In_2446);
and U5816 (N_5816,In_2656,In_547);
or U5817 (N_5817,In_2489,In_257);
xor U5818 (N_5818,In_1250,In_2768);
or U5819 (N_5819,In_862,In_526);
and U5820 (N_5820,In_2504,In_320);
and U5821 (N_5821,In_1331,In_749);
nand U5822 (N_5822,In_2014,In_740);
nor U5823 (N_5823,In_1559,In_2141);
xor U5824 (N_5824,In_2403,In_601);
nor U5825 (N_5825,In_2099,In_96);
and U5826 (N_5826,In_1192,In_661);
or U5827 (N_5827,In_100,In_2540);
or U5828 (N_5828,In_1566,In_2798);
or U5829 (N_5829,In_928,In_1015);
xnor U5830 (N_5830,In_1793,In_388);
xnor U5831 (N_5831,In_1056,In_625);
xor U5832 (N_5832,In_587,In_2383);
xnor U5833 (N_5833,In_2434,In_266);
nor U5834 (N_5834,In_2481,In_456);
or U5835 (N_5835,In_554,In_759);
nor U5836 (N_5836,In_373,In_2058);
and U5837 (N_5837,In_716,In_1278);
nor U5838 (N_5838,In_408,In_2198);
nor U5839 (N_5839,In_1529,In_2854);
and U5840 (N_5840,In_536,In_2092);
and U5841 (N_5841,In_198,In_753);
nor U5842 (N_5842,In_335,In_687);
nor U5843 (N_5843,In_1445,In_1878);
and U5844 (N_5844,In_2487,In_81);
nand U5845 (N_5845,In_2459,In_2969);
xor U5846 (N_5846,In_916,In_945);
nand U5847 (N_5847,In_2702,In_2232);
and U5848 (N_5848,In_2950,In_1015);
xnor U5849 (N_5849,In_101,In_922);
nand U5850 (N_5850,In_1431,In_170);
or U5851 (N_5851,In_1556,In_2486);
xnor U5852 (N_5852,In_1659,In_758);
nor U5853 (N_5853,In_804,In_1610);
or U5854 (N_5854,In_1001,In_2960);
nor U5855 (N_5855,In_1434,In_2571);
nor U5856 (N_5856,In_1859,In_1583);
nand U5857 (N_5857,In_2064,In_2243);
xnor U5858 (N_5858,In_2840,In_2206);
and U5859 (N_5859,In_2963,In_756);
nand U5860 (N_5860,In_174,In_1782);
xor U5861 (N_5861,In_1888,In_267);
xnor U5862 (N_5862,In_110,In_873);
and U5863 (N_5863,In_1362,In_2522);
or U5864 (N_5864,In_2194,In_2629);
nand U5865 (N_5865,In_2823,In_326);
nor U5866 (N_5866,In_551,In_2439);
xnor U5867 (N_5867,In_2746,In_2386);
nor U5868 (N_5868,In_1514,In_2758);
nand U5869 (N_5869,In_2669,In_361);
nand U5870 (N_5870,In_2393,In_1391);
or U5871 (N_5871,In_2799,In_2910);
or U5872 (N_5872,In_569,In_2179);
or U5873 (N_5873,In_1092,In_1861);
nand U5874 (N_5874,In_1217,In_2281);
xor U5875 (N_5875,In_970,In_2857);
or U5876 (N_5876,In_1830,In_762);
nand U5877 (N_5877,In_2938,In_1377);
xor U5878 (N_5878,In_2751,In_218);
nor U5879 (N_5879,In_162,In_701);
nor U5880 (N_5880,In_228,In_1479);
nor U5881 (N_5881,In_1105,In_2328);
and U5882 (N_5882,In_496,In_233);
nor U5883 (N_5883,In_2913,In_2114);
nand U5884 (N_5884,In_1651,In_1001);
and U5885 (N_5885,In_715,In_456);
nor U5886 (N_5886,In_2191,In_876);
nand U5887 (N_5887,In_2747,In_930);
nand U5888 (N_5888,In_316,In_1590);
or U5889 (N_5889,In_1212,In_1815);
or U5890 (N_5890,In_361,In_2775);
and U5891 (N_5891,In_1233,In_2526);
or U5892 (N_5892,In_1810,In_1578);
nor U5893 (N_5893,In_1296,In_1374);
nor U5894 (N_5894,In_1935,In_1789);
xor U5895 (N_5895,In_2657,In_1702);
or U5896 (N_5896,In_2716,In_2096);
nand U5897 (N_5897,In_1045,In_1729);
and U5898 (N_5898,In_528,In_1460);
nor U5899 (N_5899,In_1581,In_2735);
nand U5900 (N_5900,In_2760,In_1340);
and U5901 (N_5901,In_185,In_2852);
or U5902 (N_5902,In_1800,In_1375);
and U5903 (N_5903,In_754,In_878);
nor U5904 (N_5904,In_958,In_2296);
or U5905 (N_5905,In_124,In_1003);
nand U5906 (N_5906,In_2686,In_2196);
xor U5907 (N_5907,In_77,In_2420);
nor U5908 (N_5908,In_163,In_1833);
and U5909 (N_5909,In_64,In_2455);
nand U5910 (N_5910,In_1572,In_211);
or U5911 (N_5911,In_88,In_1146);
xor U5912 (N_5912,In_2394,In_1551);
nand U5913 (N_5913,In_116,In_516);
and U5914 (N_5914,In_566,In_2391);
nand U5915 (N_5915,In_2635,In_503);
nor U5916 (N_5916,In_2446,In_694);
nand U5917 (N_5917,In_240,In_1071);
xor U5918 (N_5918,In_2207,In_1934);
nor U5919 (N_5919,In_2488,In_1070);
nor U5920 (N_5920,In_2685,In_1770);
nand U5921 (N_5921,In_2319,In_2635);
xnor U5922 (N_5922,In_748,In_1148);
or U5923 (N_5923,In_1936,In_2261);
or U5924 (N_5924,In_2305,In_2831);
or U5925 (N_5925,In_2154,In_575);
nor U5926 (N_5926,In_1645,In_1843);
nand U5927 (N_5927,In_2362,In_2704);
and U5928 (N_5928,In_1447,In_1753);
or U5929 (N_5929,In_8,In_334);
xnor U5930 (N_5930,In_516,In_1313);
nor U5931 (N_5931,In_422,In_2874);
nor U5932 (N_5932,In_2206,In_677);
and U5933 (N_5933,In_291,In_471);
or U5934 (N_5934,In_743,In_2098);
nor U5935 (N_5935,In_2393,In_1548);
nor U5936 (N_5936,In_2682,In_1453);
and U5937 (N_5937,In_2650,In_646);
nand U5938 (N_5938,In_530,In_2549);
nand U5939 (N_5939,In_2807,In_1437);
nor U5940 (N_5940,In_948,In_1864);
or U5941 (N_5941,In_1487,In_2210);
nand U5942 (N_5942,In_490,In_2099);
nor U5943 (N_5943,In_140,In_577);
nand U5944 (N_5944,In_1792,In_993);
xnor U5945 (N_5945,In_1334,In_35);
nand U5946 (N_5946,In_440,In_2096);
nand U5947 (N_5947,In_1079,In_2880);
or U5948 (N_5948,In_1061,In_1331);
or U5949 (N_5949,In_2434,In_1297);
xor U5950 (N_5950,In_240,In_2981);
or U5951 (N_5951,In_2984,In_1153);
xnor U5952 (N_5952,In_509,In_2631);
xnor U5953 (N_5953,In_2678,In_685);
nor U5954 (N_5954,In_1230,In_2519);
nand U5955 (N_5955,In_1949,In_1508);
xor U5956 (N_5956,In_2933,In_429);
or U5957 (N_5957,In_2127,In_1285);
nand U5958 (N_5958,In_1318,In_1669);
or U5959 (N_5959,In_1389,In_2096);
nor U5960 (N_5960,In_2145,In_1215);
nor U5961 (N_5961,In_443,In_1501);
or U5962 (N_5962,In_1849,In_1518);
and U5963 (N_5963,In_2701,In_2560);
nand U5964 (N_5964,In_55,In_2637);
and U5965 (N_5965,In_2770,In_81);
nor U5966 (N_5966,In_1507,In_2163);
xnor U5967 (N_5967,In_1224,In_2457);
and U5968 (N_5968,In_1782,In_2665);
or U5969 (N_5969,In_2790,In_1089);
xnor U5970 (N_5970,In_832,In_121);
and U5971 (N_5971,In_1677,In_853);
xor U5972 (N_5972,In_1341,In_2286);
xor U5973 (N_5973,In_2623,In_1075);
and U5974 (N_5974,In_1560,In_1415);
xor U5975 (N_5975,In_2976,In_2312);
and U5976 (N_5976,In_2941,In_1365);
or U5977 (N_5977,In_1518,In_1394);
or U5978 (N_5978,In_2834,In_63);
xor U5979 (N_5979,In_1978,In_2321);
nand U5980 (N_5980,In_590,In_1183);
and U5981 (N_5981,In_2891,In_2474);
xor U5982 (N_5982,In_2898,In_2195);
xnor U5983 (N_5983,In_2340,In_1580);
nand U5984 (N_5984,In_1166,In_120);
or U5985 (N_5985,In_2645,In_1412);
xnor U5986 (N_5986,In_2157,In_444);
nor U5987 (N_5987,In_2427,In_1874);
or U5988 (N_5988,In_589,In_458);
xnor U5989 (N_5989,In_1851,In_1542);
or U5990 (N_5990,In_2701,In_2730);
xnor U5991 (N_5991,In_250,In_365);
and U5992 (N_5992,In_316,In_1959);
nand U5993 (N_5993,In_1123,In_1286);
or U5994 (N_5994,In_2680,In_1351);
nand U5995 (N_5995,In_2484,In_2968);
nor U5996 (N_5996,In_2124,In_106);
nand U5997 (N_5997,In_1082,In_140);
xnor U5998 (N_5998,In_1698,In_2335);
or U5999 (N_5999,In_2284,In_1897);
nand U6000 (N_6000,N_1090,N_5029);
nand U6001 (N_6001,N_2443,N_2244);
nor U6002 (N_6002,N_5680,N_3595);
nor U6003 (N_6003,N_2552,N_5043);
or U6004 (N_6004,N_1532,N_2966);
nor U6005 (N_6005,N_4520,N_317);
and U6006 (N_6006,N_3556,N_2239);
nand U6007 (N_6007,N_4564,N_405);
nor U6008 (N_6008,N_2070,N_3210);
or U6009 (N_6009,N_3923,N_5417);
and U6010 (N_6010,N_1740,N_4353);
xor U6011 (N_6011,N_4134,N_4169);
nor U6012 (N_6012,N_5487,N_446);
nand U6013 (N_6013,N_4957,N_4468);
xnor U6014 (N_6014,N_156,N_4918);
and U6015 (N_6015,N_1683,N_3120);
or U6016 (N_6016,N_66,N_2488);
or U6017 (N_6017,N_4195,N_4724);
or U6018 (N_6018,N_973,N_353);
xnor U6019 (N_6019,N_5096,N_4962);
nand U6020 (N_6020,N_2585,N_2571);
and U6021 (N_6021,N_153,N_2687);
nand U6022 (N_6022,N_5789,N_3925);
nand U6023 (N_6023,N_3788,N_679);
nand U6024 (N_6024,N_4793,N_283);
or U6025 (N_6025,N_3344,N_5194);
xor U6026 (N_6026,N_2883,N_724);
nand U6027 (N_6027,N_4624,N_2406);
or U6028 (N_6028,N_2914,N_1878);
or U6029 (N_6029,N_306,N_218);
xnor U6030 (N_6030,N_1169,N_239);
and U6031 (N_6031,N_2516,N_1926);
and U6032 (N_6032,N_986,N_4083);
or U6033 (N_6033,N_2996,N_2984);
xnor U6034 (N_6034,N_5059,N_108);
nand U6035 (N_6035,N_597,N_5617);
nand U6036 (N_6036,N_115,N_5757);
nor U6037 (N_6037,N_1453,N_3578);
or U6038 (N_6038,N_269,N_681);
nand U6039 (N_6039,N_733,N_3101);
nor U6040 (N_6040,N_318,N_3500);
xor U6041 (N_6041,N_1902,N_2731);
or U6042 (N_6042,N_772,N_3453);
xor U6043 (N_6043,N_3276,N_3811);
nand U6044 (N_6044,N_3449,N_1216);
or U6045 (N_6045,N_596,N_532);
nand U6046 (N_6046,N_1513,N_3954);
and U6047 (N_6047,N_492,N_2232);
xnor U6048 (N_6048,N_5798,N_3837);
nand U6049 (N_6049,N_5449,N_1019);
nand U6050 (N_6050,N_5703,N_4227);
nand U6051 (N_6051,N_1806,N_59);
xnor U6052 (N_6052,N_638,N_3367);
nor U6053 (N_6053,N_3743,N_3744);
or U6054 (N_6054,N_5512,N_2617);
nand U6055 (N_6055,N_3405,N_5038);
and U6056 (N_6056,N_5346,N_4985);
and U6057 (N_6057,N_2051,N_5685);
nand U6058 (N_6058,N_2638,N_1613);
nor U6059 (N_6059,N_2475,N_1150);
or U6060 (N_6060,N_5636,N_3422);
or U6061 (N_6061,N_4408,N_4410);
nand U6062 (N_6062,N_263,N_2316);
nor U6063 (N_6063,N_1097,N_3293);
nand U6064 (N_6064,N_1448,N_1257);
and U6065 (N_6065,N_721,N_1509);
nand U6066 (N_6066,N_4429,N_5375);
or U6067 (N_6067,N_2682,N_3263);
nand U6068 (N_6068,N_4750,N_4033);
xor U6069 (N_6069,N_932,N_803);
and U6070 (N_6070,N_1711,N_5764);
nor U6071 (N_6071,N_4805,N_383);
and U6072 (N_6072,N_5927,N_5161);
and U6073 (N_6073,N_4505,N_1096);
nor U6074 (N_6074,N_1720,N_2485);
or U6075 (N_6075,N_1722,N_579);
and U6076 (N_6076,N_1560,N_4635);
xnor U6077 (N_6077,N_5706,N_5788);
or U6078 (N_6078,N_5594,N_4010);
xor U6079 (N_6079,N_2343,N_5190);
xor U6080 (N_6080,N_1574,N_478);
and U6081 (N_6081,N_1591,N_1116);
nand U6082 (N_6082,N_3428,N_5571);
nand U6083 (N_6083,N_1788,N_3051);
and U6084 (N_6084,N_2945,N_3860);
xnor U6085 (N_6085,N_4200,N_2245);
nand U6086 (N_6086,N_2203,N_5524);
and U6087 (N_6087,N_2725,N_4725);
xor U6088 (N_6088,N_1551,N_3304);
xor U6089 (N_6089,N_3141,N_3127);
or U6090 (N_6090,N_4153,N_899);
and U6091 (N_6091,N_41,N_5835);
or U6092 (N_6092,N_1395,N_5276);
xnor U6093 (N_6093,N_5162,N_3721);
xor U6094 (N_6094,N_3368,N_3458);
or U6095 (N_6095,N_3711,N_5005);
or U6096 (N_6096,N_3203,N_1502);
or U6097 (N_6097,N_4229,N_104);
and U6098 (N_6098,N_4166,N_2860);
or U6099 (N_6099,N_4361,N_631);
nor U6100 (N_6100,N_1083,N_4614);
nand U6101 (N_6101,N_5255,N_5983);
and U6102 (N_6102,N_2065,N_3270);
or U6103 (N_6103,N_3738,N_4285);
and U6104 (N_6104,N_3661,N_1995);
nor U6105 (N_6105,N_5037,N_1203);
or U6106 (N_6106,N_2098,N_2761);
xnor U6107 (N_6107,N_4015,N_4509);
and U6108 (N_6108,N_4478,N_1317);
and U6109 (N_6109,N_3968,N_1311);
and U6110 (N_6110,N_5955,N_3482);
or U6111 (N_6111,N_1005,N_4781);
nand U6112 (N_6112,N_628,N_4995);
and U6113 (N_6113,N_2390,N_4312);
and U6114 (N_6114,N_3286,N_3872);
nand U6115 (N_6115,N_4922,N_731);
nand U6116 (N_6116,N_2364,N_3255);
nand U6117 (N_6117,N_1316,N_357);
xnor U6118 (N_6118,N_2877,N_5482);
nand U6119 (N_6119,N_1079,N_2523);
nand U6120 (N_6120,N_4121,N_3946);
or U6121 (N_6121,N_5692,N_5605);
nor U6122 (N_6122,N_1155,N_5966);
nand U6123 (N_6123,N_1534,N_3810);
nand U6124 (N_6124,N_321,N_5995);
nand U6125 (N_6125,N_309,N_3414);
or U6126 (N_6126,N_3671,N_2438);
nor U6127 (N_6127,N_1309,N_3608);
xnor U6128 (N_6128,N_940,N_100);
nand U6129 (N_6129,N_3532,N_5198);
xnor U6130 (N_6130,N_4540,N_1397);
nor U6131 (N_6131,N_1181,N_4946);
xor U6132 (N_6132,N_3506,N_3717);
nand U6133 (N_6133,N_4059,N_1458);
or U6134 (N_6134,N_3436,N_5374);
and U6135 (N_6135,N_268,N_1567);
nor U6136 (N_6136,N_4496,N_621);
nand U6137 (N_6137,N_1086,N_2896);
or U6138 (N_6138,N_3582,N_1685);
or U6139 (N_6139,N_4549,N_5174);
and U6140 (N_6140,N_5717,N_2224);
and U6141 (N_6141,N_3729,N_1709);
nor U6142 (N_6142,N_5290,N_5765);
nor U6143 (N_6143,N_4825,N_1295);
and U6144 (N_6144,N_5117,N_942);
xor U6145 (N_6145,N_3512,N_2282);
xnor U6146 (N_6146,N_5484,N_5182);
xor U6147 (N_6147,N_4425,N_5993);
and U6148 (N_6148,N_5971,N_3611);
nand U6149 (N_6149,N_4937,N_3497);
and U6150 (N_6150,N_3409,N_189);
nor U6151 (N_6151,N_2985,N_3621);
or U6152 (N_6152,N_4899,N_5508);
or U6153 (N_6153,N_5628,N_2085);
and U6154 (N_6154,N_5886,N_3131);
nor U6155 (N_6155,N_4284,N_4642);
and U6156 (N_6156,N_725,N_1290);
nand U6157 (N_6157,N_5091,N_4903);
xor U6158 (N_6158,N_686,N_869);
and U6159 (N_6159,N_1307,N_5552);
nor U6160 (N_6160,N_476,N_5268);
or U6161 (N_6161,N_3266,N_3845);
nand U6162 (N_6162,N_3797,N_5180);
or U6163 (N_6163,N_4666,N_378);
or U6164 (N_6164,N_2919,N_2878);
nand U6165 (N_6165,N_3378,N_5607);
nor U6166 (N_6166,N_3979,N_2466);
nor U6167 (N_6167,N_3577,N_5420);
nor U6168 (N_6168,N_1990,N_4542);
nor U6169 (N_6169,N_5267,N_2833);
nand U6170 (N_6170,N_1872,N_3106);
nor U6171 (N_6171,N_374,N_2901);
or U6172 (N_6172,N_1134,N_984);
or U6173 (N_6173,N_4859,N_1426);
and U6174 (N_6174,N_4902,N_2223);
nand U6175 (N_6175,N_1218,N_171);
xnor U6176 (N_6176,N_2327,N_3990);
nor U6177 (N_6177,N_4287,N_5774);
nand U6178 (N_6178,N_530,N_3960);
xor U6179 (N_6179,N_1931,N_3767);
and U6180 (N_6180,N_1456,N_1300);
and U6181 (N_6181,N_3487,N_878);
or U6182 (N_6182,N_2118,N_2353);
and U6183 (N_6183,N_3292,N_800);
and U6184 (N_6184,N_2369,N_2315);
or U6185 (N_6185,N_5304,N_5228);
and U6186 (N_6186,N_2658,N_2605);
nand U6187 (N_6187,N_2884,N_3275);
or U6188 (N_6188,N_4440,N_5170);
nor U6189 (N_6189,N_35,N_5700);
xnor U6190 (N_6190,N_1254,N_4317);
nor U6191 (N_6191,N_4352,N_4406);
xnor U6192 (N_6192,N_692,N_3514);
nor U6193 (N_6193,N_2125,N_4749);
nor U6194 (N_6194,N_4430,N_5310);
and U6195 (N_6195,N_2717,N_2242);
and U6196 (N_6196,N_3065,N_4192);
xnor U6197 (N_6197,N_1006,N_2854);
xnor U6198 (N_6198,N_3321,N_2791);
and U6199 (N_6199,N_3701,N_4180);
nand U6200 (N_6200,N_3319,N_2291);
nand U6201 (N_6201,N_210,N_3978);
or U6202 (N_6202,N_4808,N_1620);
nand U6203 (N_6203,N_4163,N_1576);
and U6204 (N_6204,N_4584,N_3124);
nand U6205 (N_6205,N_635,N_5477);
nand U6206 (N_6206,N_1894,N_5000);
xor U6207 (N_6207,N_3572,N_1879);
nand U6208 (N_6208,N_1399,N_1583);
nand U6209 (N_6209,N_2181,N_4209);
nand U6210 (N_6210,N_824,N_4242);
and U6211 (N_6211,N_1377,N_5601);
xnor U6212 (N_6212,N_4865,N_4215);
nor U6213 (N_6213,N_3570,N_5762);
nand U6214 (N_6214,N_1819,N_4127);
or U6215 (N_6215,N_1248,N_5192);
nand U6216 (N_6216,N_418,N_4024);
and U6217 (N_6217,N_5961,N_190);
or U6218 (N_6218,N_4745,N_1626);
nor U6219 (N_6219,N_1111,N_5796);
nand U6220 (N_6220,N_3333,N_2418);
nand U6221 (N_6221,N_3308,N_3305);
nor U6222 (N_6222,N_2890,N_2066);
or U6223 (N_6223,N_1929,N_2231);
or U6224 (N_6224,N_3236,N_2861);
and U6225 (N_6225,N_1544,N_3650);
xnor U6226 (N_6226,N_4398,N_3518);
nand U6227 (N_6227,N_197,N_5207);
or U6228 (N_6228,N_5036,N_5328);
xnor U6229 (N_6229,N_2851,N_4692);
and U6230 (N_6230,N_4225,N_5218);
nor U6231 (N_6231,N_1052,N_207);
and U6232 (N_6232,N_4090,N_3223);
xnor U6233 (N_6233,N_4456,N_5407);
xor U6234 (N_6234,N_649,N_1635);
xor U6235 (N_6235,N_4543,N_1588);
or U6236 (N_6236,N_5933,N_5083);
nand U6237 (N_6237,N_1563,N_1174);
or U6238 (N_6238,N_3080,N_2718);
or U6239 (N_6239,N_3774,N_380);
xor U6240 (N_6240,N_3312,N_1144);
or U6241 (N_6241,N_521,N_2057);
xnor U6242 (N_6242,N_2139,N_348);
and U6243 (N_6243,N_4139,N_565);
or U6244 (N_6244,N_5224,N_2772);
xor U6245 (N_6245,N_1507,N_1496);
or U6246 (N_6246,N_4332,N_697);
and U6247 (N_6247,N_4265,N_624);
or U6248 (N_6248,N_4880,N_212);
nor U6249 (N_6249,N_5184,N_2416);
and U6250 (N_6250,N_425,N_2991);
nor U6251 (N_6251,N_3730,N_4816);
xor U6252 (N_6252,N_4885,N_1557);
xor U6253 (N_6253,N_422,N_4518);
and U6254 (N_6254,N_5677,N_3664);
or U6255 (N_6255,N_2587,N_1897);
or U6256 (N_6256,N_4940,N_2374);
or U6257 (N_6257,N_4858,N_4275);
or U6258 (N_6258,N_5656,N_1113);
xnor U6259 (N_6259,N_7,N_2659);
and U6260 (N_6260,N_2569,N_2649);
or U6261 (N_6261,N_1302,N_3163);
nand U6262 (N_6262,N_1278,N_905);
nor U6263 (N_6263,N_3259,N_567);
nand U6264 (N_6264,N_428,N_2113);
or U6265 (N_6265,N_2848,N_5592);
nor U6266 (N_6266,N_327,N_5748);
nand U6267 (N_6267,N_4882,N_322);
nand U6268 (N_6268,N_4446,N_355);
nand U6269 (N_6269,N_3583,N_1266);
or U6270 (N_6270,N_4841,N_2820);
or U6271 (N_6271,N_768,N_4789);
nand U6272 (N_6272,N_959,N_1895);
or U6273 (N_6273,N_3814,N_4016);
nor U6274 (N_6274,N_4092,N_541);
nor U6275 (N_6275,N_3113,N_4393);
xnor U6276 (N_6276,N_3165,N_2253);
nor U6277 (N_6277,N_1958,N_3665);
xor U6278 (N_6278,N_4826,N_735);
xor U6279 (N_6279,N_688,N_3193);
and U6280 (N_6280,N_2227,N_149);
nor U6281 (N_6281,N_782,N_3053);
and U6282 (N_6282,N_2800,N_3808);
nor U6283 (N_6283,N_2467,N_4704);
and U6284 (N_6284,N_3426,N_2235);
xor U6285 (N_6285,N_5196,N_2686);
nor U6286 (N_6286,N_2367,N_3361);
or U6287 (N_6287,N_3546,N_1130);
xor U6288 (N_6288,N_421,N_2236);
and U6289 (N_6289,N_4277,N_417);
xnor U6290 (N_6290,N_5265,N_4757);
and U6291 (N_6291,N_2171,N_3600);
xnor U6292 (N_6292,N_102,N_2805);
and U6293 (N_6293,N_2908,N_3416);
nand U6294 (N_6294,N_2603,N_527);
xor U6295 (N_6295,N_4649,N_2272);
nor U6296 (N_6296,N_2373,N_3406);
nor U6297 (N_6297,N_1340,N_3930);
nand U6298 (N_6298,N_3098,N_1285);
xor U6299 (N_6299,N_3676,N_2332);
nand U6300 (N_6300,N_882,N_1310);
and U6301 (N_6301,N_5900,N_4339);
and U6302 (N_6302,N_561,N_1240);
nor U6303 (N_6303,N_5894,N_5042);
xor U6304 (N_6304,N_2850,N_3160);
or U6305 (N_6305,N_5092,N_2238);
nand U6306 (N_6306,N_3874,N_5377);
nand U6307 (N_6307,N_3599,N_627);
and U6308 (N_6308,N_2082,N_4143);
or U6309 (N_6309,N_461,N_1189);
nor U6310 (N_6310,N_5047,N_2193);
or U6311 (N_6311,N_5220,N_3474);
nand U6312 (N_6312,N_1071,N_5572);
or U6313 (N_6313,N_918,N_4994);
or U6314 (N_6314,N_4422,N_4038);
and U6315 (N_6315,N_3508,N_1183);
or U6316 (N_6316,N_840,N_4727);
or U6317 (N_6317,N_896,N_3002);
and U6318 (N_6318,N_562,N_4924);
or U6319 (N_6319,N_3015,N_3287);
xor U6320 (N_6320,N_3176,N_702);
and U6321 (N_6321,N_2305,N_2789);
or U6322 (N_6322,N_929,N_4335);
or U6323 (N_6323,N_491,N_664);
nor U6324 (N_6324,N_3742,N_3456);
xor U6325 (N_6325,N_1444,N_2034);
xor U6326 (N_6326,N_1959,N_658);
nand U6327 (N_6327,N_3951,N_2500);
nor U6328 (N_6328,N_4778,N_3554);
xor U6329 (N_6329,N_5274,N_2565);
nor U6330 (N_6330,N_5028,N_2149);
nor U6331 (N_6331,N_689,N_246);
nand U6332 (N_6332,N_2133,N_2625);
or U6333 (N_6333,N_5133,N_3828);
nor U6334 (N_6334,N_1371,N_5926);
nand U6335 (N_6335,N_162,N_4917);
or U6336 (N_6336,N_4787,N_1360);
and U6337 (N_6337,N_3039,N_4098);
nand U6338 (N_6338,N_2976,N_1853);
xor U6339 (N_6339,N_719,N_4157);
or U6340 (N_6340,N_2929,N_1691);
nand U6341 (N_6341,N_1949,N_1801);
xnor U6342 (N_6342,N_332,N_5734);
xnor U6343 (N_6343,N_2216,N_2463);
or U6344 (N_6344,N_4401,N_2351);
xnor U6345 (N_6345,N_3912,N_2176);
and U6346 (N_6346,N_501,N_5011);
xnor U6347 (N_6347,N_5881,N_2795);
xnor U6348 (N_6348,N_2511,N_2226);
or U6349 (N_6349,N_3649,N_2698);
nor U6350 (N_6350,N_1575,N_5053);
xor U6351 (N_6351,N_5786,N_1766);
and U6352 (N_6352,N_651,N_3782);
xor U6353 (N_6353,N_4258,N_933);
or U6354 (N_6354,N_5625,N_5464);
xnor U6355 (N_6355,N_3465,N_3069);
xnor U6356 (N_6356,N_2397,N_4610);
nand U6357 (N_6357,N_4751,N_3964);
nor U6358 (N_6358,N_1651,N_26);
nor U6359 (N_6359,N_2811,N_2492);
nand U6360 (N_6360,N_5749,N_3061);
xnor U6361 (N_6361,N_186,N_4276);
or U6362 (N_6362,N_1112,N_1478);
nor U6363 (N_6363,N_1412,N_141);
and U6364 (N_6364,N_533,N_3815);
nor U6365 (N_6365,N_356,N_3237);
xnor U6366 (N_6366,N_487,N_1775);
nor U6367 (N_6367,N_4367,N_1736);
nor U6368 (N_6368,N_4007,N_1392);
nor U6369 (N_6369,N_1343,N_2147);
xor U6370 (N_6370,N_715,N_1463);
xor U6371 (N_6371,N_2283,N_5880);
nor U6372 (N_6372,N_3753,N_4253);
nor U6373 (N_6373,N_3396,N_1188);
xnor U6374 (N_6374,N_3343,N_2408);
and U6375 (N_6375,N_4554,N_748);
or U6376 (N_6376,N_3168,N_5175);
or U6377 (N_6377,N_5299,N_1027);
xor U6378 (N_6378,N_5266,N_3706);
or U6379 (N_6379,N_470,N_3358);
xnor U6380 (N_6380,N_390,N_5861);
nor U6381 (N_6381,N_1900,N_5666);
and U6382 (N_6382,N_5538,N_1986);
nor U6383 (N_6383,N_13,N_3088);
nand U6384 (N_6384,N_249,N_598);
or U6385 (N_6385,N_3220,N_3598);
nand U6386 (N_6386,N_3454,N_1579);
or U6387 (N_6387,N_9,N_3626);
nor U6388 (N_6388,N_5869,N_3023);
xor U6389 (N_6389,N_3330,N_4949);
nor U6390 (N_6390,N_2997,N_2348);
or U6391 (N_6391,N_2869,N_647);
and U6392 (N_6392,N_2513,N_1105);
nand U6393 (N_6393,N_2295,N_548);
nor U6394 (N_6394,N_93,N_4346);
and U6395 (N_6395,N_4026,N_625);
nand U6396 (N_6396,N_1061,N_4741);
nand U6397 (N_6397,N_836,N_489);
and U6398 (N_6398,N_4099,N_2602);
nand U6399 (N_6399,N_5370,N_2323);
nand U6400 (N_6400,N_415,N_4034);
xor U6401 (N_6401,N_915,N_996);
nand U6402 (N_6402,N_2208,N_2304);
nor U6403 (N_6403,N_4055,N_2963);
or U6404 (N_6404,N_1401,N_3843);
and U6405 (N_6405,N_1919,N_1157);
nand U6406 (N_6406,N_240,N_1941);
nand U6407 (N_6407,N_2872,N_5221);
and U6408 (N_6408,N_5506,N_4879);
nor U6409 (N_6409,N_570,N_1264);
and U6410 (N_6410,N_3250,N_1523);
nor U6411 (N_6411,N_3760,N_5159);
xnor U6412 (N_6412,N_5390,N_366);
nand U6413 (N_6413,N_5223,N_5819);
and U6414 (N_6414,N_2473,N_3579);
and U6415 (N_6415,N_1535,N_5132);
or U6416 (N_6416,N_5637,N_1622);
xor U6417 (N_6417,N_3256,N_2944);
nor U6418 (N_6418,N_566,N_3639);
xor U6419 (N_6419,N_2897,N_759);
or U6420 (N_6420,N_904,N_2881);
and U6421 (N_6421,N_4115,N_3261);
nand U6422 (N_6422,N_2331,N_4457);
nand U6423 (N_6423,N_1000,N_4194);
nor U6424 (N_6424,N_5782,N_507);
nand U6425 (N_6425,N_769,N_1383);
nand U6426 (N_6426,N_480,N_1272);
xnor U6427 (N_6427,N_4417,N_3686);
nand U6428 (N_6428,N_3102,N_4113);
and U6429 (N_6429,N_11,N_5609);
xor U6430 (N_6430,N_4293,N_2469);
xnor U6431 (N_6431,N_5815,N_3629);
or U6432 (N_6432,N_3823,N_3432);
nor U6433 (N_6433,N_5459,N_2240);
nor U6434 (N_6434,N_1693,N_1245);
or U6435 (N_6435,N_2254,N_2298);
nor U6436 (N_6436,N_4598,N_5082);
nand U6437 (N_6437,N_4118,N_510);
or U6438 (N_6438,N_4535,N_3590);
or U6439 (N_6439,N_75,N_3971);
and U6440 (N_6440,N_4204,N_3317);
nand U6441 (N_6441,N_4498,N_4782);
or U6442 (N_6442,N_3094,N_5416);
xnor U6443 (N_6443,N_3737,N_773);
nand U6444 (N_6444,N_1356,N_4548);
or U6445 (N_6445,N_2197,N_3638);
and U6446 (N_6446,N_1283,N_2655);
or U6447 (N_6447,N_3682,N_4892);
xnor U6448 (N_6448,N_2818,N_219);
nand U6449 (N_6449,N_276,N_3152);
nand U6450 (N_6450,N_4824,N_2542);
nor U6451 (N_6451,N_4510,N_610);
nor U6452 (N_6452,N_2062,N_4264);
nand U6453 (N_6453,N_5535,N_3566);
nor U6454 (N_6454,N_5289,N_1963);
and U6455 (N_6455,N_1742,N_76);
nor U6456 (N_6456,N_4883,N_5746);
nor U6457 (N_6457,N_1639,N_4951);
and U6458 (N_6458,N_4474,N_4183);
or U6459 (N_6459,N_3589,N_3181);
and U6460 (N_6460,N_5797,N_4578);
and U6461 (N_6461,N_2968,N_5118);
and U6462 (N_6462,N_743,N_1794);
and U6463 (N_6463,N_5325,N_1488);
nand U6464 (N_6464,N_3509,N_4222);
and U6465 (N_6465,N_2180,N_555);
and U6466 (N_6466,N_5022,N_3313);
nor U6467 (N_6467,N_4168,N_4057);
xor U6468 (N_6468,N_3043,N_3792);
or U6469 (N_6469,N_2407,N_3014);
and U6470 (N_6470,N_4066,N_3194);
xnor U6471 (N_6471,N_3145,N_5766);
or U6472 (N_6472,N_1199,N_1748);
nand U6473 (N_6473,N_5629,N_3515);
nand U6474 (N_6474,N_675,N_161);
nor U6475 (N_6475,N_4680,N_3271);
nand U6476 (N_6476,N_1539,N_2145);
or U6477 (N_6477,N_3662,N_2915);
xnor U6478 (N_6478,N_1614,N_4095);
or U6479 (N_6479,N_738,N_4976);
or U6480 (N_6480,N_3784,N_1674);
or U6481 (N_6481,N_5451,N_2219);
xnor U6482 (N_6482,N_320,N_238);
nor U6483 (N_6483,N_2150,N_5439);
nor U6484 (N_6484,N_3614,N_3602);
xor U6485 (N_6485,N_4071,N_1476);
nor U6486 (N_6486,N_3530,N_1924);
xnor U6487 (N_6487,N_922,N_2217);
xnor U6488 (N_6488,N_2312,N_4839);
nor U6489 (N_6489,N_2678,N_1612);
xor U6490 (N_6490,N_1844,N_5492);
and U6491 (N_6491,N_2849,N_4615);
and U6492 (N_6492,N_3592,N_395);
nand U6493 (N_6493,N_1547,N_294);
xnor U6494 (N_6494,N_4077,N_1044);
and U6495 (N_6495,N_3349,N_2421);
nor U6496 (N_6496,N_994,N_3175);
xor U6497 (N_6497,N_3408,N_3427);
nor U6498 (N_6498,N_116,N_1351);
xnor U6499 (N_6499,N_3001,N_581);
nand U6500 (N_6500,N_4923,N_2358);
and U6501 (N_6501,N_975,N_2105);
nor U6502 (N_6502,N_4492,N_3699);
nand U6503 (N_6503,N_5751,N_1676);
nand U6504 (N_6504,N_5795,N_912);
xor U6505 (N_6505,N_1885,N_794);
xor U6506 (N_6506,N_1190,N_3574);
nand U6507 (N_6507,N_1214,N_5347);
xnor U6508 (N_6508,N_4573,N_131);
xor U6509 (N_6509,N_5496,N_4357);
xor U6510 (N_6510,N_5204,N_1602);
nand U6511 (N_6511,N_4330,N_1684);
nand U6512 (N_6512,N_3955,N_2285);
xor U6513 (N_6513,N_5684,N_5831);
nand U6514 (N_6514,N_5147,N_5001);
nand U6515 (N_6515,N_534,N_4605);
xnor U6516 (N_6516,N_1881,N_1700);
nand U6517 (N_6517,N_4980,N_832);
xnor U6518 (N_6518,N_2898,N_4864);
and U6519 (N_6519,N_5879,N_90);
nor U6520 (N_6520,N_713,N_1255);
nand U6521 (N_6521,N_4999,N_3214);
nand U6522 (N_6522,N_3460,N_2828);
or U6523 (N_6523,N_2071,N_2159);
xor U6524 (N_6524,N_5309,N_3603);
nand U6525 (N_6525,N_2187,N_613);
nor U6526 (N_6526,N_2114,N_4145);
nor U6527 (N_6527,N_5587,N_2391);
or U6528 (N_6528,N_5154,N_5682);
nand U6529 (N_6529,N_2940,N_3331);
and U6530 (N_6530,N_2271,N_4586);
and U6531 (N_6531,N_698,N_5079);
nor U6532 (N_6532,N_1652,N_1370);
nand U6533 (N_6533,N_3318,N_1981);
xor U6534 (N_6534,N_4319,N_4633);
xnor U6535 (N_6535,N_1129,N_1455);
xor U6536 (N_6536,N_5596,N_946);
nand U6537 (N_6537,N_256,N_2797);
or U6538 (N_6538,N_1994,N_5504);
nand U6539 (N_6539,N_3419,N_5997);
or U6540 (N_6540,N_2465,N_2221);
xor U6541 (N_6541,N_12,N_4851);
xnor U6542 (N_6542,N_122,N_3804);
nand U6543 (N_6543,N_1018,N_2646);
or U6544 (N_6544,N_5131,N_808);
and U6545 (N_6545,N_682,N_1841);
nand U6546 (N_6546,N_1127,N_3550);
nand U6547 (N_6547,N_5604,N_92);
or U6548 (N_6548,N_2441,N_410);
or U6549 (N_6549,N_2478,N_5217);
nor U6550 (N_6550,N_3136,N_1493);
and U6551 (N_6551,N_1462,N_5686);
and U6552 (N_6552,N_5052,N_3242);
and U6553 (N_6553,N_2262,N_5622);
nand U6554 (N_6554,N_802,N_2243);
and U6555 (N_6555,N_3545,N_3529);
xor U6556 (N_6556,N_4022,N_2430);
and U6557 (N_6557,N_5713,N_4416);
nor U6558 (N_6558,N_1067,N_298);
nor U6559 (N_6559,N_1039,N_5776);
xnor U6560 (N_6560,N_1718,N_5583);
nand U6561 (N_6561,N_4551,N_2371);
xor U6562 (N_6562,N_5485,N_693);
nand U6563 (N_6563,N_63,N_5094);
and U6564 (N_6564,N_4792,N_1553);
xor U6565 (N_6565,N_4512,N_5424);
or U6566 (N_6566,N_220,N_5657);
or U6567 (N_6567,N_1091,N_4640);
nor U6568 (N_6568,N_4131,N_4819);
and U6569 (N_6569,N_1843,N_2049);
and U6570 (N_6570,N_5292,N_5303);
nand U6571 (N_6571,N_1184,N_1654);
and U6572 (N_6572,N_3437,N_3710);
or U6573 (N_6573,N_2589,N_4511);
and U6574 (N_6574,N_2429,N_1584);
xnor U6575 (N_6575,N_148,N_1874);
nor U6576 (N_6576,N_5191,N_4343);
or U6577 (N_6577,N_3221,N_4128);
and U6578 (N_6578,N_2887,N_3169);
and U6579 (N_6579,N_4658,N_1056);
or U6580 (N_6580,N_1605,N_4958);
nor U6581 (N_6581,N_351,N_1855);
and U6582 (N_6582,N_3423,N_17);
nor U6583 (N_6583,N_2733,N_2675);
and U6584 (N_6584,N_314,N_5662);
nand U6585 (N_6585,N_1793,N_4028);
or U6586 (N_6586,N_5856,N_1439);
xor U6587 (N_6587,N_1969,N_4075);
or U6588 (N_6588,N_1314,N_1274);
nand U6589 (N_6589,N_5651,N_2975);
xnor U6590 (N_6590,N_5306,N_1768);
nor U6591 (N_6591,N_5984,N_4506);
and U6592 (N_6592,N_2266,N_4004);
or U6593 (N_6593,N_1944,N_399);
and U6594 (N_6594,N_2606,N_1447);
nor U6595 (N_6595,N_74,N_1103);
nand U6596 (N_6596,N_5939,N_1518);
nor U6597 (N_6597,N_1012,N_5702);
and U6598 (N_6598,N_790,N_3790);
and U6599 (N_6599,N_2684,N_4291);
xor U6600 (N_6600,N_5233,N_4931);
nor U6601 (N_6601,N_1207,N_1480);
xnor U6602 (N_6602,N_1298,N_2752);
xor U6603 (N_6603,N_1580,N_438);
xnor U6604 (N_6604,N_224,N_3447);
xor U6605 (N_6605,N_4837,N_2444);
nand U6606 (N_6606,N_2460,N_4964);
nor U6607 (N_6607,N_465,N_2209);
and U6608 (N_6608,N_1373,N_5985);
nor U6609 (N_6609,N_4581,N_1242);
nor U6610 (N_6610,N_3931,N_4556);
nor U6611 (N_6611,N_1530,N_2503);
xnor U6612 (N_6612,N_5273,N_5020);
or U6613 (N_6613,N_5863,N_3854);
or U6614 (N_6614,N_3763,N_164);
or U6615 (N_6615,N_5495,N_2892);
xnor U6616 (N_6616,N_5072,N_2679);
or U6617 (N_6617,N_2609,N_5623);
nor U6618 (N_6618,N_1938,N_4973);
nand U6619 (N_6619,N_2889,N_2362);
nor U6620 (N_6620,N_3435,N_5804);
and U6621 (N_6621,N_3997,N_1331);
and U6622 (N_6622,N_5380,N_1032);
or U6623 (N_6623,N_537,N_4555);
or U6624 (N_6624,N_890,N_1824);
xor U6625 (N_6625,N_4762,N_1890);
nor U6626 (N_6626,N_5839,N_4453);
nor U6627 (N_6627,N_3620,N_3452);
nor U6628 (N_6628,N_5836,N_5383);
and U6629 (N_6629,N_5923,N_3462);
or U6630 (N_6630,N_602,N_1671);
and U6631 (N_6631,N_5802,N_3553);
or U6632 (N_6632,N_146,N_3996);
or U6633 (N_6633,N_5531,N_5603);
and U6634 (N_6634,N_1960,N_4613);
nor U6635 (N_6635,N_2981,N_4847);
and U6636 (N_6636,N_2959,N_1407);
and U6637 (N_6637,N_4173,N_4821);
nor U6638 (N_6638,N_2179,N_3666);
or U6639 (N_6639,N_5807,N_919);
nor U6640 (N_6640,N_3593,N_1440);
nand U6641 (N_6641,N_1643,N_1767);
or U6642 (N_6642,N_1870,N_985);
nor U6643 (N_6643,N_5248,N_3898);
xnor U6644 (N_6644,N_4685,N_4273);
nand U6645 (N_6645,N_2656,N_4728);
xor U6646 (N_6646,N_2263,N_3480);
or U6647 (N_6647,N_5210,N_228);
xnor U6648 (N_6648,N_538,N_1686);
nor U6649 (N_6649,N_4220,N_2763);
nor U6650 (N_6650,N_2228,N_5387);
or U6651 (N_6651,N_5376,N_2307);
or U6652 (N_6652,N_135,N_4673);
xnor U6653 (N_6653,N_3888,N_3148);
and U6654 (N_6654,N_2581,N_4412);
nor U6655 (N_6655,N_870,N_2626);
nor U6656 (N_6656,N_5647,N_5429);
nor U6657 (N_6657,N_1782,N_2624);
nor U6658 (N_6658,N_407,N_586);
nand U6659 (N_6659,N_5723,N_2001);
or U6660 (N_6660,N_2121,N_4775);
or U6661 (N_6661,N_2200,N_4539);
xor U6662 (N_6662,N_2056,N_1727);
nand U6663 (N_6663,N_1047,N_4230);
nor U6664 (N_6664,N_1756,N_577);
and U6665 (N_6665,N_5278,N_2726);
nor U6666 (N_6666,N_2019,N_4694);
or U6667 (N_6667,N_1372,N_4739);
nor U6668 (N_6668,N_5433,N_4829);
xor U6669 (N_6669,N_4914,N_4419);
xnor U6670 (N_6670,N_5171,N_5924);
xor U6671 (N_6671,N_1306,N_616);
nand U6672 (N_6672,N_368,N_467);
xor U6673 (N_6673,N_546,N_170);
and U6674 (N_6674,N_3869,N_2029);
nor U6675 (N_6675,N_1861,N_3660);
or U6676 (N_6676,N_3958,N_4027);
nand U6677 (N_6677,N_301,N_3768);
nor U6678 (N_6678,N_3643,N_1549);
or U6679 (N_6679,N_2470,N_1470);
nor U6680 (N_6680,N_2012,N_3778);
or U6681 (N_6681,N_179,N_5744);
nor U6682 (N_6682,N_1858,N_1644);
and U6683 (N_6683,N_3571,N_4175);
and U6684 (N_6684,N_3268,N_2947);
or U6685 (N_6685,N_3502,N_4959);
nor U6686 (N_6686,N_5458,N_2086);
nor U6687 (N_6687,N_1378,N_5260);
nand U6688 (N_6688,N_2637,N_4405);
xnor U6689 (N_6689,N_5741,N_3994);
and U6690 (N_6690,N_4513,N_954);
nor U6691 (N_6691,N_494,N_4934);
nand U6692 (N_6692,N_1491,N_1080);
xor U6693 (N_6693,N_916,N_603);
xor U6694 (N_6694,N_1212,N_5876);
xnor U6695 (N_6695,N_5483,N_4526);
nor U6696 (N_6696,N_4399,N_2876);
nand U6697 (N_6697,N_4376,N_1765);
xnor U6698 (N_6698,N_637,N_3689);
xor U6699 (N_6699,N_3455,N_2858);
and U6700 (N_6700,N_1821,N_4085);
nor U6701 (N_6701,N_1585,N_2598);
nand U6702 (N_6702,N_4262,N_2337);
and U6703 (N_6703,N_2928,N_1800);
or U6704 (N_6704,N_403,N_826);
nand U6705 (N_6705,N_2506,N_2786);
nor U6706 (N_6706,N_1481,N_3212);
nand U6707 (N_6707,N_2045,N_917);
and U6708 (N_6708,N_496,N_4479);
and U6709 (N_6709,N_2296,N_1318);
xnor U6710 (N_6710,N_5003,N_457);
nor U6711 (N_6711,N_2146,N_3787);
or U6712 (N_6712,N_5203,N_3354);
xor U6713 (N_6713,N_1754,N_483);
or U6714 (N_6714,N_2387,N_3952);
nand U6715 (N_6715,N_5873,N_3071);
or U6716 (N_6716,N_5699,N_1349);
nor U6717 (N_6717,N_1839,N_3272);
nand U6718 (N_6718,N_2932,N_1508);
nor U6719 (N_6719,N_1007,N_44);
nor U6720 (N_6720,N_3693,N_2411);
or U6721 (N_6721,N_622,N_1556);
nor U6722 (N_6722,N_5659,N_113);
xor U6723 (N_6723,N_3617,N_4340);
nor U6724 (N_6724,N_4476,N_4001);
and U6725 (N_6725,N_1128,N_2508);
nor U6726 (N_6726,N_4008,N_4094);
xor U6727 (N_6727,N_456,N_3902);
or U6728 (N_6728,N_2053,N_5676);
xor U6729 (N_6729,N_3531,N_3704);
nand U6730 (N_6730,N_2110,N_4919);
or U6731 (N_6731,N_1603,N_4280);
nor U6732 (N_6732,N_2946,N_4720);
or U6733 (N_6733,N_5409,N_5382);
or U6734 (N_6734,N_4871,N_3842);
nor U6735 (N_6735,N_4256,N_3832);
xnor U6736 (N_6736,N_2462,N_2412);
or U6737 (N_6737,N_1659,N_3327);
or U6738 (N_6738,N_5206,N_3457);
xor U6739 (N_6739,N_4254,N_4645);
and U6740 (N_6740,N_4203,N_1177);
nor U6741 (N_6741,N_5404,N_3526);
and U6742 (N_6742,N_39,N_771);
xor U6743 (N_6743,N_2050,N_2680);
xor U6744 (N_6744,N_5148,N_4961);
xor U6745 (N_6745,N_2455,N_3000);
nor U6746 (N_6746,N_1978,N_742);
nand U6747 (N_6747,N_237,N_4072);
nor U6748 (N_6748,N_1002,N_969);
nor U6749 (N_6749,N_392,N_3848);
and U6750 (N_6750,N_411,N_5414);
and U6751 (N_6751,N_5358,N_1543);
xnor U6752 (N_6752,N_2995,N_1382);
and U6753 (N_6753,N_1152,N_5398);
and U6754 (N_6754,N_4671,N_1410);
nand U6755 (N_6755,N_4122,N_2611);
nor U6756 (N_6756,N_4091,N_5178);
or U6757 (N_6757,N_126,N_3332);
nor U6758 (N_6758,N_3935,N_3555);
and U6759 (N_6759,N_3161,N_2629);
nor U6760 (N_6760,N_4259,N_2924);
nor U6761 (N_6761,N_3026,N_5335);
nand U6762 (N_6762,N_1436,N_230);
and U6763 (N_6763,N_2987,N_868);
nor U6764 (N_6764,N_1664,N_4979);
or U6765 (N_6765,N_4972,N_4799);
nor U6766 (N_6766,N_5491,N_2835);
xnor U6767 (N_6767,N_750,N_1419);
xnor U6768 (N_6768,N_888,N_3190);
or U6769 (N_6769,N_3260,N_5550);
and U6770 (N_6770,N_4852,N_2192);
and U6771 (N_6771,N_1914,N_5724);
nor U6772 (N_6772,N_1609,N_3981);
and U6773 (N_6773,N_5039,N_2433);
nor U6774 (N_6774,N_4870,N_1637);
xnor U6775 (N_6775,N_3393,N_4849);
xnor U6776 (N_6776,N_1252,N_1650);
xnor U6777 (N_6777,N_1831,N_389);
nor U6778 (N_6778,N_163,N_343);
xor U6779 (N_6779,N_1390,N_807);
and U6780 (N_6780,N_4358,N_2061);
xor U6781 (N_6781,N_2135,N_1961);
or U6782 (N_6782,N_3215,N_4191);
nand U6783 (N_6783,N_5754,N_2895);
nand U6784 (N_6784,N_4060,N_4233);
or U6785 (N_6785,N_3865,N_902);
nand U6786 (N_6786,N_3179,N_2198);
and U6787 (N_6787,N_542,N_4497);
xnor U6788 (N_6788,N_5738,N_2955);
nand U6789 (N_6789,N_3722,N_3995);
and U6790 (N_6790,N_1016,N_2158);
nand U6791 (N_6791,N_1171,N_4014);
nand U6792 (N_6792,N_2837,N_1822);
and U6793 (N_6793,N_2368,N_2038);
or U6794 (N_6794,N_4521,N_5542);
xor U6795 (N_6795,N_2130,N_5031);
nand U6796 (N_6796,N_3122,N_1089);
xor U6797 (N_6797,N_1799,N_1421);
nor U6798 (N_6798,N_2359,N_3688);
and U6799 (N_6799,N_5639,N_3387);
or U6800 (N_6800,N_493,N_183);
xor U6801 (N_6801,N_387,N_5081);
xor U6802 (N_6802,N_4895,N_887);
nor U6803 (N_6803,N_5826,N_4449);
nand U6804 (N_6804,N_2865,N_4350);
nand U6805 (N_6805,N_924,N_880);
nand U6806 (N_6806,N_1696,N_3873);
or U6807 (N_6807,N_2740,N_3541);
xnor U6808 (N_6808,N_1702,N_1132);
xnor U6809 (N_6809,N_3905,N_1732);
and U6810 (N_6810,N_1838,N_1342);
or U6811 (N_6811,N_594,N_4000);
xnor U6812 (N_6812,N_5912,N_4913);
or U6813 (N_6813,N_5286,N_3834);
and U6814 (N_6814,N_347,N_5714);
and U6815 (N_6815,N_3383,N_5388);
xnor U6816 (N_6816,N_3177,N_3024);
or U6817 (N_6817,N_2360,N_1780);
xor U6818 (N_6818,N_5127,N_4431);
or U6819 (N_6819,N_1863,N_2402);
xnor U6820 (N_6820,N_589,N_599);
and U6821 (N_6821,N_229,N_3974);
or U6822 (N_6822,N_3476,N_4846);
nand U6823 (N_6823,N_3950,N_334);
xor U6824 (N_6824,N_1784,N_5155);
xor U6825 (N_6825,N_2302,N_1149);
or U6826 (N_6826,N_2035,N_3709);
nor U6827 (N_6827,N_4356,N_233);
nor U6828 (N_6828,N_5264,N_1260);
xor U6829 (N_6829,N_3404,N_5084);
or U6830 (N_6830,N_335,N_5988);
and U6831 (N_6831,N_3539,N_3533);
and U6832 (N_6832,N_4427,N_1186);
or U6833 (N_6833,N_947,N_3696);
xor U6834 (N_6834,N_3381,N_587);
nor U6835 (N_6835,N_1850,N_1570);
xnor U6836 (N_6836,N_1076,N_5421);
xor U6837 (N_6837,N_2037,N_5410);
and U6838 (N_6838,N_2691,N_3929);
xor U6839 (N_6839,N_3133,N_2212);
or U6840 (N_6840,N_2810,N_3745);
or U6841 (N_6841,N_1675,N_453);
nand U6842 (N_6842,N_5152,N_5413);
or U6843 (N_6843,N_5940,N_4659);
nand U6844 (N_6844,N_4046,N_5513);
xor U6845 (N_6845,N_2688,N_4011);
xor U6846 (N_6846,N_2592,N_4828);
or U6847 (N_6847,N_1167,N_3619);
nor U6848 (N_6848,N_2151,N_1231);
nor U6849 (N_6849,N_214,N_4908);
xor U6850 (N_6850,N_4652,N_3382);
nor U6851 (N_6851,N_974,N_2422);
xor U6852 (N_6852,N_2471,N_4900);
xor U6853 (N_6853,N_4714,N_2826);
nor U6854 (N_6854,N_818,N_5794);
nand U6855 (N_6855,N_2090,N_4838);
xnor U6856 (N_6856,N_1077,N_2671);
or U6857 (N_6857,N_1966,N_31);
or U6858 (N_6858,N_4770,N_1369);
nand U6859 (N_6859,N_4968,N_1474);
xor U6860 (N_6860,N_2785,N_3669);
and U6861 (N_6861,N_2823,N_1928);
or U6862 (N_6862,N_4984,N_3524);
xor U6863 (N_6863,N_5235,N_2261);
and U6864 (N_6864,N_2426,N_4550);
nand U6865 (N_6865,N_4351,N_3940);
or U6866 (N_6866,N_2410,N_3780);
nand U6867 (N_6867,N_4928,N_4300);
and U6868 (N_6868,N_962,N_1517);
xnor U6869 (N_6869,N_949,N_3459);
xnor U6870 (N_6870,N_206,N_671);
and U6871 (N_6871,N_391,N_5418);
and U6872 (N_6872,N_73,N_1847);
or U6873 (N_6873,N_3967,N_5891);
and U6874 (N_6874,N_4684,N_3939);
xor U6875 (N_6875,N_945,N_5750);
nand U6876 (N_6876,N_5101,N_5990);
xnor U6877 (N_6877,N_2095,N_1689);
and U6878 (N_6878,N_1725,N_4068);
or U6879 (N_6879,N_3254,N_1569);
xor U6880 (N_6880,N_3280,N_4706);
nor U6881 (N_6881,N_4911,N_372);
or U6882 (N_6882,N_2248,N_5867);
xnor U6883 (N_6883,N_1717,N_866);
xor U6884 (N_6884,N_5500,N_2917);
and U6885 (N_6885,N_2002,N_2880);
nand U6886 (N_6886,N_56,N_1363);
or U6887 (N_6887,N_4019,N_5199);
xor U6888 (N_6888,N_2619,N_536);
and U6889 (N_6889,N_1037,N_1942);
or U6890 (N_6890,N_4662,N_5002);
and U6891 (N_6891,N_4665,N_176);
nand U6892 (N_6892,N_4198,N_5241);
and U6893 (N_6893,N_2322,N_5440);
nor U6894 (N_6894,N_5360,N_3496);
xnor U6895 (N_6895,N_3403,N_563);
or U6896 (N_6896,N_3913,N_703);
and U6897 (N_6897,N_5396,N_462);
xnor U6898 (N_6898,N_3062,N_316);
or U6899 (N_6899,N_4460,N_2532);
nand U6900 (N_6900,N_4664,N_4411);
xnor U6901 (N_6901,N_5883,N_5120);
xnor U6902 (N_6902,N_779,N_5143);
xnor U6903 (N_6903,N_812,N_4423);
nand U6904 (N_6904,N_1505,N_5030);
and U6905 (N_6905,N_5465,N_87);
and U6906 (N_6906,N_3209,N_3316);
and U6907 (N_6907,N_1380,N_4981);
and U6908 (N_6908,N_5818,N_690);
nand U6909 (N_6909,N_3827,N_1542);
nand U6910 (N_6910,N_5935,N_1625);
xnor U6911 (N_6911,N_1122,N_4948);
or U6912 (N_6912,N_4246,N_4688);
nand U6913 (N_6913,N_1294,N_2798);
nor U6914 (N_6914,N_4184,N_2132);
xnor U6915 (N_6915,N_4676,N_5551);
nand U6916 (N_6916,N_3424,N_3892);
or U6917 (N_6917,N_2702,N_5478);
xnor U6918 (N_6918,N_311,N_5785);
and U6919 (N_6919,N_2714,N_2827);
nand U6920 (N_6920,N_5105,N_5050);
nand U6921 (N_6921,N_1522,N_1940);
or U6922 (N_6922,N_2127,N_4631);
xor U6923 (N_6923,N_1098,N_4036);
xor U6924 (N_6924,N_508,N_5044);
nor U6925 (N_6925,N_2148,N_5259);
nand U6926 (N_6926,N_4217,N_3297);
and U6927 (N_6927,N_2561,N_660);
nand U6928 (N_6928,N_1734,N_3575);
nand U6929 (N_6929,N_1494,N_2573);
xor U6930 (N_6930,N_5124,N_3623);
xnor U6931 (N_6931,N_4061,N_2925);
and U6932 (N_6932,N_1472,N_4176);
nand U6933 (N_6933,N_1085,N_5648);
nand U6934 (N_6934,N_221,N_3471);
and U6935 (N_6935,N_1368,N_2891);
or U6936 (N_6936,N_5564,N_528);
nor U6937 (N_6937,N_753,N_2366);
nor U6938 (N_6938,N_2083,N_2610);
or U6939 (N_6939,N_3109,N_1910);
xnor U6940 (N_6940,N_2616,N_2549);
or U6941 (N_6941,N_4243,N_720);
nand U6942 (N_6942,N_3045,N_661);
nor U6943 (N_6943,N_5896,N_2768);
nand U6944 (N_6944,N_3521,N_2935);
nor U6945 (N_6945,N_1361,N_5026);
or U6946 (N_6946,N_3850,N_612);
or U6947 (N_6947,N_696,N_1108);
nor U6948 (N_6948,N_2445,N_4773);
nand U6949 (N_6949,N_265,N_3056);
nor U6950 (N_6950,N_3228,N_4593);
nand U6951 (N_6951,N_4767,N_1922);
xnor U6952 (N_6952,N_5557,N_4630);
nor U6953 (N_6953,N_1348,N_2535);
nor U6954 (N_6954,N_495,N_3117);
or U6955 (N_6955,N_5582,N_4251);
xor U6956 (N_6956,N_4969,N_4383);
xor U6957 (N_6957,N_1589,N_1814);
or U6958 (N_6958,N_3733,N_2623);
nor U6959 (N_6959,N_3055,N_2449);
xnor U6960 (N_6960,N_1172,N_3021);
or U6961 (N_6961,N_2456,N_3295);
or U6962 (N_6962,N_152,N_977);
nor U6963 (N_6963,N_861,N_3948);
or U6964 (N_6964,N_3833,N_4833);
or U6965 (N_6965,N_2140,N_1891);
and U6966 (N_6966,N_3352,N_2222);
xnor U6967 (N_6967,N_5113,N_4611);
nor U6968 (N_6968,N_2009,N_535);
nand U6969 (N_6969,N_2068,N_3284);
nor U6970 (N_6970,N_4044,N_2423);
and U6971 (N_6971,N_1078,N_4623);
nand U6972 (N_6972,N_497,N_4618);
nand U6973 (N_6973,N_5817,N_1345);
nand U6974 (N_6974,N_3921,N_77);
nand U6975 (N_6975,N_4616,N_234);
nor U6976 (N_6976,N_103,N_4407);
nand U6977 (N_6977,N_3656,N_4796);
nand U6978 (N_6978,N_5716,N_1572);
nor U6979 (N_6979,N_2269,N_5518);
nor U6980 (N_6980,N_4103,N_5431);
xor U6981 (N_6981,N_3817,N_5709);
and U6982 (N_6982,N_1437,N_2712);
and U6983 (N_6983,N_3648,N_5242);
xnor U6984 (N_6984,N_1706,N_4037);
nor U6985 (N_6985,N_381,N_3357);
xnor U6986 (N_6986,N_2059,N_2375);
nand U6987 (N_6987,N_1912,N_5457);
nor U6988 (N_6988,N_3060,N_3551);
and U6989 (N_6989,N_5996,N_4360);
and U6990 (N_6990,N_5394,N_3520);
xor U6991 (N_6991,N_1564,N_2273);
nand U6992 (N_6992,N_1715,N_3486);
or U6993 (N_6993,N_4179,N_5627);
nand U6994 (N_6994,N_615,N_3245);
or U6995 (N_6995,N_5488,N_1297);
xnor U6996 (N_6996,N_5010,N_3251);
nor U6997 (N_6997,N_798,N_3200);
xnor U6998 (N_6998,N_5930,N_1516);
xnor U6999 (N_6999,N_303,N_3339);
nand U7000 (N_7000,N_350,N_2807);
or U7001 (N_7001,N_5066,N_2910);
nor U7002 (N_7002,N_3442,N_5690);
or U7003 (N_7003,N_3003,N_5618);
nor U7004 (N_7004,N_3594,N_5517);
nand U7005 (N_7005,N_3334,N_5858);
nand U7006 (N_7006,N_1856,N_4190);
xnor U7007 (N_7007,N_1989,N_3273);
xnor U7008 (N_7008,N_155,N_325);
xnor U7009 (N_7009,N_3347,N_1082);
and U7010 (N_7010,N_4832,N_1417);
xnor U7011 (N_7011,N_1156,N_4310);
nor U7012 (N_7012,N_5379,N_4172);
nor U7013 (N_7013,N_27,N_2695);
or U7014 (N_7014,N_5450,N_5910);
nor U7015 (N_7015,N_5922,N_3887);
xor U7016 (N_7016,N_3969,N_5139);
or U7017 (N_7017,N_3895,N_642);
nor U7018 (N_7018,N_2326,N_4784);
or U7019 (N_7019,N_4448,N_1434);
nor U7020 (N_7020,N_5959,N_1611);
nand U7021 (N_7021,N_4532,N_4005);
or U7022 (N_7022,N_241,N_2742);
and U7023 (N_7023,N_3824,N_5430);
xnor U7024 (N_7024,N_3877,N_1514);
xor U7025 (N_7025,N_5674,N_2381);
or U7026 (N_7026,N_550,N_5875);
nor U7027 (N_7027,N_3732,N_5576);
nand U7028 (N_7028,N_4647,N_2885);
xnor U7029 (N_7029,N_3727,N_1692);
and U7030 (N_7030,N_5791,N_2138);
and U7031 (N_7031,N_1956,N_1999);
xor U7032 (N_7032,N_3868,N_4588);
and U7033 (N_7033,N_3234,N_4653);
nand U7034 (N_7034,N_1058,N_5872);
nor U7035 (N_7035,N_64,N_3646);
nand U7036 (N_7036,N_2864,N_2276);
or U7037 (N_7037,N_1915,N_3795);
nand U7038 (N_7038,N_5434,N_5511);
nor U7039 (N_7039,N_5405,N_5855);
and U7040 (N_7040,N_4996,N_1951);
or U7041 (N_7041,N_2284,N_5962);
and U7042 (N_7042,N_1420,N_2949);
nand U7043 (N_7043,N_4488,N_5825);
nor U7044 (N_7044,N_4558,N_30);
nor U7045 (N_7045,N_3751,N_2525);
nor U7046 (N_7046,N_2186,N_142);
xor U7047 (N_7047,N_1497,N_678);
and U7048 (N_7048,N_150,N_1606);
nand U7049 (N_7049,N_3822,N_1649);
and U7050 (N_7050,N_1680,N_1276);
nand U7051 (N_7051,N_4644,N_1192);
nor U7052 (N_7052,N_4487,N_5140);
or U7053 (N_7053,N_36,N_2496);
xor U7054 (N_7054,N_1029,N_3963);
nand U7055 (N_7055,N_4294,N_3791);
xnor U7056 (N_7056,N_4561,N_4777);
or U7057 (N_7057,N_5172,N_1304);
nor U7058 (N_7058,N_4585,N_2859);
xnor U7059 (N_7059,N_582,N_2521);
and U7060 (N_7060,N_4544,N_300);
xnor U7061 (N_7061,N_2094,N_3705);
and U7062 (N_7062,N_2184,N_2648);
xnor U7063 (N_7063,N_2013,N_1561);
nor U7064 (N_7064,N_5077,N_4566);
and U7065 (N_7065,N_1498,N_5247);
xnor U7066 (N_7066,N_1251,N_2336);
or U7067 (N_7067,N_4729,N_1694);
nor U7068 (N_7068,N_444,N_2612);
nand U7069 (N_7069,N_5761,N_2417);
xor U7070 (N_7070,N_3915,N_2642);
or U7071 (N_7071,N_4189,N_2540);
xor U7072 (N_7072,N_1424,N_1893);
or U7073 (N_7073,N_2155,N_2153);
nor U7074 (N_7074,N_1735,N_3988);
and U7075 (N_7075,N_3536,N_185);
and U7076 (N_7076,N_761,N_4041);
nand U7077 (N_7077,N_1808,N_120);
and U7078 (N_7078,N_5558,N_2994);
nand U7079 (N_7079,N_5045,N_683);
and U7080 (N_7080,N_2667,N_2074);
and U7081 (N_7081,N_502,N_5938);
xnor U7082 (N_7082,N_5994,N_5725);
or U7083 (N_7083,N_3034,N_4413);
nor U7084 (N_7084,N_2386,N_3859);
and U7085 (N_7085,N_3985,N_3206);
xnor U7086 (N_7086,N_2017,N_3641);
or U7087 (N_7087,N_3973,N_2972);
or U7088 (N_7088,N_4056,N_1327);
nand U7089 (N_7089,N_3323,N_367);
or U7090 (N_7090,N_5874,N_3776);
nor U7091 (N_7091,N_5792,N_1341);
xnor U7092 (N_7092,N_2566,N_2527);
and U7093 (N_7093,N_1287,N_5668);
nand U7094 (N_7094,N_46,N_5320);
nand U7095 (N_7095,N_2732,N_5463);
nand U7096 (N_7096,N_471,N_1244);
xor U7097 (N_7097,N_22,N_3813);
xor U7098 (N_7098,N_956,N_2292);
xor U7099 (N_7099,N_5978,N_2518);
or U7100 (N_7100,N_2233,N_3903);
and U7101 (N_7101,N_3785,N_4261);
or U7102 (N_7102,N_2808,N_2683);
nor U7103 (N_7103,N_5441,N_1852);
xor U7104 (N_7104,N_5909,N_5701);
nand U7105 (N_7105,N_5362,N_5510);
and U7106 (N_7106,N_4536,N_4458);
nand U7107 (N_7107,N_2737,N_5580);
nor U7108 (N_7108,N_2681,N_1751);
or U7109 (N_7109,N_5689,N_3401);
nor U7110 (N_7110,N_3796,N_5486);
and U7111 (N_7111,N_2363,N_3607);
and U7112 (N_7112,N_2847,N_4313);
or U7113 (N_7113,N_3446,N_3634);
nor U7114 (N_7114,N_1074,N_2863);
nand U7115 (N_7115,N_583,N_1663);
nand U7116 (N_7116,N_2930,N_4737);
and U7117 (N_7117,N_1170,N_4455);
nor U7118 (N_7118,N_4516,N_5344);
xnor U7119 (N_7119,N_4212,N_2088);
and U7120 (N_7120,N_2904,N_1066);
or U7121 (N_7121,N_2129,N_4905);
nor U7122 (N_7122,N_3097,N_4252);
and U7123 (N_7123,N_980,N_3581);
nor U7124 (N_7124,N_3340,N_3451);
nand U7125 (N_7125,N_3461,N_1063);
and U7126 (N_7126,N_4205,N_3067);
nand U7127 (N_7127,N_3998,N_5693);
xnor U7128 (N_7128,N_3324,N_4089);
xor U7129 (N_7129,N_4648,N_3517);
nand U7130 (N_7130,N_3841,N_5770);
nor U7131 (N_7131,N_310,N_3941);
or U7132 (N_7132,N_5357,N_3070);
and U7133 (N_7133,N_3882,N_3830);
nand U7134 (N_7134,N_854,N_2663);
and U7135 (N_7135,N_944,N_1191);
or U7136 (N_7136,N_1143,N_3105);
nand U7137 (N_7137,N_1536,N_4876);
nand U7138 (N_7138,N_1404,N_5633);
nand U7139 (N_7139,N_1690,N_1641);
nor U7140 (N_7140,N_2196,N_2644);
and U7141 (N_7141,N_3932,N_460);
and U7142 (N_7142,N_2657,N_2100);
and U7143 (N_7143,N_416,N_1288);
nand U7144 (N_7144,N_1059,N_910);
nand U7145 (N_7145,N_4454,N_3198);
nand U7146 (N_7146,N_3360,N_1355);
xor U7147 (N_7147,N_404,N_2309);
xor U7148 (N_7148,N_3836,N_451);
or U7149 (N_7149,N_2738,N_5279);
xor U7150 (N_7150,N_5777,N_2841);
or U7151 (N_7151,N_2128,N_3018);
nand U7152 (N_7152,N_3908,N_668);
and U7153 (N_7153,N_4503,N_1776);
xnor U7154 (N_7154,N_1202,N_1393);
or U7155 (N_7155,N_645,N_4124);
xnor U7156 (N_7156,N_4154,N_2365);
or U7157 (N_7157,N_1215,N_5381);
nand U7158 (N_7158,N_3137,N_788);
and U7159 (N_7159,N_1050,N_828);
nand U7160 (N_7160,N_4569,N_4904);
or U7161 (N_7161,N_5019,N_5004);
nand U7162 (N_7162,N_2666,N_5115);
nand U7163 (N_7163,N_5048,N_1357);
and U7164 (N_7164,N_1219,N_4626);
nor U7165 (N_7165,N_2318,N_295);
nor U7166 (N_7166,N_2134,N_4743);
nand U7167 (N_7167,N_1749,N_2690);
or U7168 (N_7168,N_192,N_2782);
xnor U7169 (N_7169,N_2956,N_302);
and U7170 (N_7170,N_1592,N_2600);
nor U7171 (N_7171,N_255,N_1827);
xnor U7172 (N_7172,N_3042,N_2790);
or U7173 (N_7173,N_5696,N_4384);
nor U7174 (N_7174,N_5800,N_1595);
or U7175 (N_7175,N_5809,N_2308);
and U7176 (N_7176,N_2764,N_5915);
nor U7177 (N_7177,N_3548,N_5600);
or U7178 (N_7178,N_1471,N_2152);
and U7179 (N_7179,N_5111,N_2893);
xor U7180 (N_7180,N_2933,N_2705);
and U7181 (N_7181,N_4178,N_763);
nor U7182 (N_7182,N_4811,N_3922);
or U7183 (N_7183,N_3373,N_2344);
xor U7184 (N_7184,N_2464,N_4249);
nor U7185 (N_7185,N_2766,N_271);
nor U7186 (N_7186,N_1423,N_4491);
nand U7187 (N_7187,N_147,N_3522);
or U7188 (N_7188,N_1770,N_4834);
nor U7189 (N_7189,N_5902,N_4935);
nor U7190 (N_7190,N_2108,N_906);
xnor U7191 (N_7191,N_5866,N_4221);
xnor U7192 (N_7192,N_4297,N_3329);
nor U7193 (N_7193,N_4954,N_3740);
xnor U7194 (N_7194,N_3899,N_2734);
nand U7195 (N_7195,N_5342,N_3289);
nor U7196 (N_7196,N_2595,N_3170);
nor U7197 (N_7197,N_913,N_5525);
nor U7198 (N_7198,N_2225,N_1927);
xnor U7199 (N_7199,N_5112,N_4464);
or U7200 (N_7200,N_4840,N_2916);
xor U7201 (N_7201,N_5426,N_4538);
nand U7202 (N_7202,N_2545,N_620);
nand U7203 (N_7203,N_1003,N_5107);
xor U7204 (N_7204,N_281,N_1807);
or U7205 (N_7205,N_5135,N_3298);
xnor U7206 (N_7206,N_3306,N_2819);
or U7207 (N_7207,N_1594,N_5354);
nand U7208 (N_7208,N_1427,N_3528);
nor U7209 (N_7209,N_3473,N_571);
and U7210 (N_7210,N_4281,N_260);
nor U7211 (N_7211,N_5803,N_5183);
and U7212 (N_7212,N_3875,N_503);
xor U7213 (N_7213,N_4199,N_1418);
nor U7214 (N_7214,N_726,N_5730);
xnor U7215 (N_7215,N_3155,N_5372);
or U7216 (N_7216,N_655,N_3746);
or U7217 (N_7217,N_1933,N_5691);
or U7218 (N_7218,N_3011,N_4656);
xor U7219 (N_7219,N_1991,N_2514);
or U7220 (N_7220,N_5917,N_5168);
nand U7221 (N_7221,N_5537,N_3208);
or U7222 (N_7222,N_1328,N_4240);
nand U7223 (N_7223,N_5138,N_5969);
xor U7224 (N_7224,N_823,N_892);
nand U7225 (N_7225,N_1632,N_1173);
or U7226 (N_7226,N_3376,N_5116);
xor U7227 (N_7227,N_1501,N_2921);
nand U7228 (N_7228,N_4021,N_6);
xor U7229 (N_7229,N_4687,N_2746);
xnor U7230 (N_7230,N_2483,N_4670);
xnor U7231 (N_7231,N_412,N_3444);
or U7232 (N_7232,N_3725,N_509);
or U7233 (N_7233,N_3748,N_1586);
nor U7234 (N_7234,N_4185,N_512);
nand U7235 (N_7235,N_2758,N_5121);
or U7236 (N_7236,N_3219,N_3752);
nand U7237 (N_7237,N_2167,N_2191);
or U7238 (N_7238,N_1842,N_2378);
or U7239 (N_7239,N_3597,N_2993);
nand U7240 (N_7240,N_3694,N_4887);
nand U7241 (N_7241,N_3944,N_601);
nand U7242 (N_7242,N_40,N_1515);
xor U7243 (N_7243,N_4161,N_1225);
and U7244 (N_7244,N_3366,N_3510);
nand U7245 (N_7245,N_3847,N_2607);
nand U7246 (N_7246,N_4370,N_5675);
or U7247 (N_7247,N_2970,N_1333);
and U7248 (N_7248,N_4155,N_2489);
and U7249 (N_7249,N_1224,N_2404);
xnor U7250 (N_7250,N_4211,N_716);
xor U7251 (N_7251,N_402,N_4866);
or U7252 (N_7252,N_137,N_2264);
xor U7253 (N_7253,N_2102,N_4069);
xnor U7254 (N_7254,N_694,N_4967);
or U7255 (N_7255,N_557,N_4078);
nor U7256 (N_7256,N_3394,N_3498);
xnor U7257 (N_7257,N_2579,N_3100);
xor U7258 (N_7258,N_2459,N_4070);
nand U7259 (N_7259,N_1428,N_2306);
and U7260 (N_7260,N_4126,N_2393);
nor U7261 (N_7261,N_1980,N_2384);
and U7262 (N_7262,N_2560,N_209);
xor U7263 (N_7263,N_225,N_5213);
nor U7264 (N_7264,N_3303,N_2515);
nand U7265 (N_7265,N_511,N_1757);
nand U7266 (N_7266,N_2010,N_4369);
or U7267 (N_7267,N_1565,N_3647);
and U7268 (N_7268,N_680,N_3421);
or U7269 (N_7269,N_1289,N_4862);
nand U7270 (N_7270,N_3691,N_712);
nand U7271 (N_7271,N_3314,N_5340);
xor U7272 (N_7272,N_4752,N_5104);
nand U7273 (N_7273,N_1187,N_4855);
xnor U7274 (N_7274,N_5934,N_134);
xor U7275 (N_7275,N_4086,N_248);
or U7276 (N_7276,N_3362,N_2632);
and U7277 (N_7277,N_1092,N_5727);
xnor U7278 (N_7278,N_4500,N_1973);
nand U7279 (N_7279,N_1618,N_3196);
nand U7280 (N_7280,N_853,N_5842);
xor U7281 (N_7281,N_1468,N_3150);
and U7282 (N_7282,N_5964,N_3402);
or U7283 (N_7283,N_4991,N_5307);
nor U7284 (N_7284,N_5015,N_4170);
xor U7285 (N_7285,N_2982,N_5694);
nand U7286 (N_7286,N_1627,N_4907);
and U7287 (N_7287,N_2376,N_2042);
and U7288 (N_7288,N_549,N_1972);
nor U7289 (N_7289,N_2647,N_3519);
xnor U7290 (N_7290,N_3173,N_4674);
and U7291 (N_7291,N_5324,N_5158);
or U7292 (N_7292,N_5554,N_5932);
nand U7293 (N_7293,N_308,N_2802);
nand U7294 (N_7294,N_3672,N_3491);
nor U7295 (N_7295,N_1701,N_3274);
or U7296 (N_7296,N_3992,N_2170);
nor U7297 (N_7297,N_4920,N_2286);
nand U7298 (N_7298,N_2943,N_964);
nand U7299 (N_7299,N_195,N_5621);
xnor U7300 (N_7300,N_3685,N_1487);
and U7301 (N_7301,N_2836,N_128);
nand U7302 (N_7302,N_1182,N_4324);
nand U7303 (N_7303,N_4290,N_1597);
and U7304 (N_7304,N_2023,N_1001);
or U7305 (N_7305,N_5968,N_4990);
xnor U7306 (N_7306,N_3277,N_2693);
or U7307 (N_7307,N_5157,N_1510);
nand U7308 (N_7308,N_3893,N_5569);
nor U7309 (N_7309,N_4404,N_5638);
or U7310 (N_7310,N_5363,N_140);
nor U7311 (N_7311,N_1554,N_2722);
or U7312 (N_7312,N_2330,N_618);
nand U7313 (N_7313,N_4668,N_1804);
nor U7314 (N_7314,N_4266,N_3418);
and U7315 (N_7315,N_413,N_3914);
nand U7316 (N_7316,N_1267,N_4975);
nor U7317 (N_7317,N_5688,N_2776);
or U7318 (N_7318,N_3856,N_953);
and U7319 (N_7319,N_4715,N_1975);
and U7320 (N_7320,N_2538,N_5811);
and U7321 (N_7321,N_5540,N_4323);
or U7322 (N_7322,N_5254,N_4705);
nand U7323 (N_7323,N_1140,N_2188);
xnor U7324 (N_7324,N_607,N_3966);
xnor U7325 (N_7325,N_3675,N_2447);
nand U7326 (N_7326,N_1035,N_5888);
or U7327 (N_7327,N_1110,N_3677);
nor U7328 (N_7328,N_1227,N_2101);
nor U7329 (N_7329,N_1280,N_3047);
nor U7330 (N_7330,N_1273,N_2104);
or U7331 (N_7331,N_3064,N_1239);
or U7332 (N_7332,N_2008,N_1120);
nor U7333 (N_7333,N_4591,N_1967);
xnor U7334 (N_7334,N_2544,N_4486);
and U7335 (N_7335,N_4053,N_4686);
and U7336 (N_7336,N_2249,N_463);
and U7337 (N_7337,N_1647,N_262);
nor U7338 (N_7338,N_1011,N_5645);
nor U7339 (N_7339,N_3775,N_3479);
or U7340 (N_7340,N_3557,N_2461);
nand U7341 (N_7341,N_5270,N_687);
and U7342 (N_7342,N_5967,N_5415);
nor U7343 (N_7343,N_1010,N_834);
or U7344 (N_7344,N_5333,N_1398);
or U7345 (N_7345,N_4006,N_2792);
xnor U7346 (N_7346,N_3678,N_514);
nand U7347 (N_7347,N_3900,N_4533);
nand U7348 (N_7348,N_5733,N_2413);
and U7349 (N_7349,N_4395,N_1452);
or U7350 (N_7350,N_2165,N_1993);
nand U7351 (N_7351,N_3534,N_4599);
xor U7352 (N_7352,N_1811,N_1125);
or U7353 (N_7353,N_3601,N_1738);
nor U7354 (N_7354,N_409,N_1653);
nand U7355 (N_7355,N_5122,N_540);
nand U7356 (N_7356,N_5944,N_3720);
nand U7357 (N_7357,N_5246,N_2618);
xnor U7358 (N_7358,N_5163,N_4912);
or U7359 (N_7359,N_1087,N_2613);
or U7360 (N_7360,N_951,N_3037);
or U7361 (N_7361,N_893,N_4164);
or U7362 (N_7362,N_3700,N_5169);
and U7363 (N_7363,N_1697,N_741);
nor U7364 (N_7364,N_3038,N_4519);
nor U7365 (N_7365,N_865,N_1889);
nor U7366 (N_7366,N_1223,N_4804);
xnor U7367 (N_7367,N_1828,N_4884);
and U7368 (N_7368,N_5920,N_5249);
or U7369 (N_7369,N_1562,N_2572);
or U7370 (N_7370,N_4269,N_1728);
and U7371 (N_7371,N_2247,N_5230);
xnor U7372 (N_7372,N_3027,N_365);
or U7373 (N_7373,N_643,N_4755);
or U7374 (N_7374,N_1578,N_1906);
and U7375 (N_7375,N_3195,N_3389);
nand U7376 (N_7376,N_2866,N_1305);
or U7377 (N_7377,N_5998,N_5743);
and U7378 (N_7378,N_5298,N_1303);
nor U7379 (N_7379,N_3211,N_5893);
or U7380 (N_7380,N_2015,N_3226);
or U7381 (N_7381,N_1763,N_1004);
nor U7382 (N_7382,N_2674,N_5176);
nand U7383 (N_7383,N_623,N_1862);
nand U7384 (N_7384,N_858,N_98);
nand U7385 (N_7385,N_2174,N_5720);
xor U7386 (N_7386,N_3159,N_5987);
and U7387 (N_7387,N_2380,N_4400);
xor U7388 (N_7388,N_2570,N_4791);
nand U7389 (N_7389,N_3013,N_4943);
xnor U7390 (N_7390,N_3494,N_4587);
nand U7391 (N_7391,N_859,N_3140);
and U7392 (N_7392,N_4490,N_717);
nor U7393 (N_7393,N_5715,N_4162);
and U7394 (N_7394,N_3390,N_101);
nand U7395 (N_7395,N_4726,N_3463);
nand U7396 (N_7396,N_795,N_1974);
and U7397 (N_7397,N_3852,N_5661);
or U7398 (N_7398,N_5125,N_943);
or U7399 (N_7399,N_2172,N_903);
nand U7400 (N_7400,N_4759,N_490);
nand U7401 (N_7401,N_4326,N_989);
or U7402 (N_7402,N_5514,N_1262);
nor U7403 (N_7403,N_5642,N_816);
and U7404 (N_7404,N_4442,N_86);
xnor U7405 (N_7405,N_5945,N_4875);
or U7406 (N_7406,N_5799,N_1908);
nor U7407 (N_7407,N_5275,N_5099);
and U7408 (N_7408,N_4790,N_5852);
xor U7409 (N_7409,N_5177,N_5767);
and U7410 (N_7410,N_5824,N_874);
nor U7411 (N_7411,N_1930,N_3723);
nor U7412 (N_7412,N_2379,N_3041);
xor U7413 (N_7413,N_923,N_5573);
and U7414 (N_7414,N_2568,N_3513);
nor U7415 (N_7415,N_3269,N_646);
nor U7416 (N_7416,N_5400,N_5614);
and U7417 (N_7417,N_2458,N_5589);
and U7418 (N_7418,N_1646,N_2967);
nand U7419 (N_7419,N_1787,N_4756);
and U7420 (N_7420,N_2979,N_2389);
nand U7421 (N_7421,N_5041,N_5384);
or U7422 (N_7422,N_1099,N_2750);
nor U7423 (N_7423,N_5958,N_3695);
xor U7424 (N_7424,N_3185,N_1781);
xnor U7425 (N_7425,N_4344,N_1818);
xor U7426 (N_7426,N_1771,N_2120);
nor U7427 (N_7427,N_4388,N_701);
or U7428 (N_7428,N_1733,N_2124);
nand U7429 (N_7429,N_213,N_481);
nand U7430 (N_7430,N_4965,N_930);
and U7431 (N_7431,N_3819,N_1162);
nor U7432 (N_7432,N_4950,N_1492);
nand U7433 (N_7433,N_3636,N_5545);
xnor U7434 (N_7434,N_2951,N_732);
nand U7435 (N_7435,N_5356,N_474);
nand U7436 (N_7436,N_4553,N_2633);
and U7437 (N_7437,N_5301,N_217);
nor U7438 (N_7438,N_1422,N_2804);
or U7439 (N_7439,N_5868,N_3005);
nor U7440 (N_7440,N_5533,N_3911);
xnor U7441 (N_7441,N_4608,N_4354);
nand U7442 (N_7442,N_2937,N_4271);
nand U7443 (N_7443,N_296,N_3816);
and U7444 (N_7444,N_4397,N_4299);
nor U7445 (N_7445,N_42,N_737);
nand U7446 (N_7446,N_1166,N_4672);
and U7447 (N_7447,N_5840,N_3143);
nor U7448 (N_7448,N_477,N_2361);
nand U7449 (N_7449,N_3077,N_1511);
nor U7450 (N_7450,N_657,N_2528);
nor U7451 (N_7451,N_3559,N_2097);
and U7452 (N_7452,N_3674,N_3802);
and U7453 (N_7453,N_2730,N_4434);
nand U7454 (N_7454,N_5942,N_2435);
xnor U7455 (N_7455,N_691,N_723);
or U7456 (N_7456,N_3991,N_4836);
nor U7457 (N_7457,N_551,N_443);
and U7458 (N_7458,N_2747,N_53);
xor U7459 (N_7459,N_2297,N_1209);
or U7460 (N_7460,N_2052,N_5392);
nor U7461 (N_7461,N_558,N_5365);
or U7462 (N_7462,N_4282,N_2334);
and U7463 (N_7463,N_2472,N_2021);
and U7464 (N_7464,N_2530,N_4325);
xor U7465 (N_7465,N_3591,N_3564);
xor U7466 (N_7466,N_1925,N_2564);
or U7467 (N_7467,N_5683,N_831);
and U7468 (N_7468,N_2962,N_952);
nor U7469 (N_7469,N_2636,N_3484);
nor U7470 (N_7470,N_2321,N_4110);
nand U7471 (N_7471,N_5865,N_5064);
and U7472 (N_7472,N_3030,N_3073);
or U7473 (N_7473,N_1848,N_226);
xor U7474 (N_7474,N_5361,N_2329);
and U7475 (N_7475,N_1911,N_1779);
nand U7476 (N_7476,N_2495,N_3095);
xor U7477 (N_7477,N_1634,N_3412);
xor U7478 (N_7478,N_590,N_5821);
or U7479 (N_7479,N_3240,N_420);
xor U7480 (N_7480,N_3906,N_1950);
or U7481 (N_7481,N_3162,N_49);
nor U7482 (N_7482,N_3146,N_5890);
and U7483 (N_7483,N_4603,N_529);
xor U7484 (N_7484,N_4682,N_1277);
and U7485 (N_7485,N_1920,N_4363);
and U7486 (N_7486,N_3035,N_5918);
nor U7487 (N_7487,N_4886,N_71);
nor U7488 (N_7488,N_5768,N_2621);
nand U7489 (N_7489,N_963,N_5035);
or U7490 (N_7490,N_4697,N_3341);
xnor U7491 (N_7491,N_264,N_4663);
nand U7492 (N_7492,N_4568,N_2558);
xor U7493 (N_7493,N_4080,N_1467);
or U7494 (N_7494,N_2450,N_1987);
and U7495 (N_7495,N_2436,N_3448);
nand U7496 (N_7496,N_2706,N_3712);
or U7497 (N_7497,N_3156,N_4120);
or U7498 (N_7498,N_5128,N_2157);
xor U7499 (N_7499,N_5351,N_5102);
xor U7500 (N_7500,N_3806,N_3835);
xnor U7501 (N_7501,N_4156,N_2548);
nand U7502 (N_7502,N_2517,N_4385);
or U7503 (N_7503,N_5186,N_3040);
nor U7504 (N_7504,N_3884,N_2482);
nand U7505 (N_7505,N_5919,N_3586);
or U7506 (N_7506,N_862,N_4202);
nand U7507 (N_7507,N_3464,N_3659);
or U7508 (N_7508,N_2809,N_2559);
nand U7509 (N_7509,N_1234,N_4797);
or U7510 (N_7510,N_1997,N_4003);
nand U7511 (N_7511,N_3468,N_939);
or U7512 (N_7512,N_82,N_815);
nand U7513 (N_7513,N_5460,N_5948);
nand U7514 (N_7514,N_193,N_4480);
nand U7515 (N_7515,N_4927,N_5046);
xnor U7516 (N_7516,N_5151,N_1258);
or U7517 (N_7517,N_1443,N_4054);
xnor U7518 (N_7518,N_1558,N_5728);
and U7519 (N_7519,N_1541,N_846);
nand U7520 (N_7520,N_4575,N_5529);
or U7521 (N_7521,N_1604,N_525);
nand U7522 (N_7522,N_5075,N_1062);
and U7523 (N_7523,N_1334,N_4753);
nand U7524 (N_7524,N_1475,N_2069);
and U7525 (N_7525,N_3119,N_2028);
and U7526 (N_7526,N_117,N_172);
nor U7527 (N_7527,N_1196,N_5581);
and U7528 (N_7528,N_4629,N_1322);
or U7529 (N_7529,N_1965,N_4807);
nor U7530 (N_7530,N_4765,N_3076);
nand U7531 (N_7531,N_4292,N_786);
and U7532 (N_7532,N_377,N_4783);
xor U7533 (N_7533,N_4048,N_4130);
or U7534 (N_7534,N_4888,N_5773);
or U7535 (N_7535,N_2575,N_95);
and U7536 (N_7536,N_4636,N_4655);
and U7537 (N_7537,N_4696,N_5747);
and U7538 (N_7538,N_4930,N_5574);
nand U7539 (N_7539,N_965,N_4529);
nor U7540 (N_7540,N_5051,N_5833);
nor U7541 (N_7541,N_4571,N_5681);
and U7542 (N_7542,N_2829,N_2160);
or U7543 (N_7543,N_4079,N_633);
and U7544 (N_7544,N_838,N_3871);
nor U7545 (N_7545,N_3075,N_313);
xnor U7546 (N_7546,N_3670,N_3082);
nor U7547 (N_7547,N_3052,N_1031);
and U7548 (N_7548,N_4723,N_3972);
nor U7549 (N_7549,N_4868,N_1825);
and U7550 (N_7550,N_4541,N_632);
nand U7551 (N_7551,N_1338,N_3663);
nand U7552 (N_7552,N_5137,N_4806);
or U7553 (N_7553,N_5566,N_2394);
or U7554 (N_7554,N_799,N_1983);
nor U7555 (N_7555,N_2164,N_5801);
nor U7556 (N_7556,N_5444,N_1060);
xor U7557 (N_7557,N_5490,N_2067);
nand U7558 (N_7558,N_997,N_1433);
or U7559 (N_7559,N_5016,N_747);
xor U7560 (N_7560,N_3605,N_652);
nor U7561 (N_7561,N_3439,N_3779);
and U7562 (N_7562,N_2428,N_2765);
or U7563 (N_7563,N_1408,N_1785);
or U7564 (N_7564,N_81,N_5085);
nor U7565 (N_7565,N_109,N_67);
xnor U7566 (N_7566,N_2615,N_1238);
or U7567 (N_7567,N_5871,N_235);
nor U7568 (N_7568,N_5205,N_1815);
nor U7569 (N_7569,N_2112,N_3821);
xnor U7570 (N_7570,N_5911,N_3217);
nor U7571 (N_7571,N_1326,N_3558);
nor U7572 (N_7572,N_5368,N_4942);
xor U7573 (N_7573,N_1201,N_1450);
and U7574 (N_7574,N_2781,N_107);
xnor U7575 (N_7575,N_4901,N_10);
or U7576 (N_7576,N_4241,N_5497);
nor U7577 (N_7577,N_4776,N_4744);
or U7578 (N_7578,N_2392,N_3719);
or U7579 (N_7579,N_3483,N_3290);
nand U7580 (N_7580,N_4764,N_3880);
xnor U7581 (N_7581,N_0,N_3063);
nor U7582 (N_7582,N_1737,N_1859);
and U7583 (N_7583,N_3407,N_730);
xor U7584 (N_7584,N_4364,N_4960);
or U7585 (N_7585,N_718,N_3235);
and U7586 (N_7586,N_950,N_55);
or U7587 (N_7587,N_3167,N_3562);
nand U7588 (N_7588,N_1817,N_4810);
xnor U7589 (N_7589,N_5232,N_3262);
nor U7590 (N_7590,N_3501,N_414);
xor U7591 (N_7591,N_4580,N_4355);
nor U7592 (N_7592,N_5813,N_2320);
xnor U7593 (N_7593,N_1425,N_4362);
or U7594 (N_7594,N_1607,N_1114);
xnor U7595 (N_7595,N_5611,N_2230);
and U7596 (N_7596,N_5468,N_4174);
or U7597 (N_7597,N_3036,N_4067);
xnor U7598 (N_7598,N_1213,N_2886);
or U7599 (N_7599,N_2520,N_2409);
nand U7600 (N_7600,N_2630,N_5308);
xnor U7601 (N_7601,N_960,N_1301);
xor U7602 (N_7602,N_324,N_2965);
xor U7603 (N_7603,N_243,N_20);
or U7604 (N_7604,N_4159,N_187);
xor U7605 (N_7605,N_1753,N_5479);
nor U7606 (N_7606,N_5916,N_3129);
nand U7607 (N_7607,N_1045,N_2255);
nand U7608 (N_7608,N_5236,N_5391);
nor U7609 (N_7609,N_1464,N_482);
and U7610 (N_7610,N_2770,N_545);
and U7611 (N_7611,N_2163,N_762);
and U7612 (N_7612,N_2287,N_4470);
xnor U7613 (N_7613,N_3878,N_3505);
xnor U7614 (N_7614,N_4747,N_5759);
xnor U7615 (N_7615,N_3540,N_4238);
xnor U7616 (N_7616,N_2580,N_2669);
nand U7617 (N_7617,N_1628,N_5349);
nor U7618 (N_7618,N_605,N_346);
xnor U7619 (N_7619,N_5074,N_4643);
and U7620 (N_7620,N_1724,N_3134);
nand U7621 (N_7621,N_722,N_3535);
or U7622 (N_7622,N_1710,N_851);
or U7623 (N_7623,N_970,N_1708);
xor U7624 (N_7624,N_4177,N_4301);
nand U7625 (N_7625,N_3747,N_5585);
or U7626 (N_7626,N_5188,N_1587);
or U7627 (N_7627,N_4443,N_4432);
nor U7628 (N_7628,N_3320,N_388);
xnor U7629 (N_7629,N_5,N_1743);
and U7630 (N_7630,N_1883,N_3511);
xnor U7631 (N_7631,N_1261,N_118);
and U7632 (N_7632,N_4827,N_2510);
nor U7633 (N_7633,N_5315,N_850);
nand U7634 (N_7634,N_955,N_5021);
nor U7635 (N_7635,N_2354,N_4409);
xnor U7636 (N_7636,N_1048,N_2080);
and U7637 (N_7637,N_5284,N_5291);
nand U7638 (N_7638,N_886,N_4108);
nor U7639 (N_7639,N_5195,N_2723);
nand U7640 (N_7640,N_2662,N_4589);
nor U7641 (N_7641,N_4771,N_5179);
and U7642 (N_7642,N_1854,N_3862);
nor U7643 (N_7643,N_341,N_979);
and U7644 (N_7644,N_791,N_5584);
or U7645 (N_7645,N_921,N_5438);
and U7646 (N_7646,N_5503,N_3032);
nor U7647 (N_7647,N_4823,N_2741);
nor U7648 (N_7648,N_3777,N_136);
or U7649 (N_7649,N_2703,N_3202);
and U7650 (N_7650,N_5598,N_165);
or U7651 (N_7651,N_2838,N_2383);
or U7652 (N_7652,N_151,N_1241);
nand U7653 (N_7653,N_2154,N_4379);
xor U7654 (N_7654,N_5698,N_5277);
nand U7655 (N_7655,N_4257,N_236);
or U7656 (N_7656,N_5025,N_4896);
nand U7657 (N_7657,N_3085,N_3769);
and U7658 (N_7658,N_4627,N_5054);
nand U7659 (N_7659,N_3,N_885);
and U7660 (N_7660,N_4105,N_3385);
or U7661 (N_7661,N_1538,N_5812);
or U7662 (N_7662,N_1119,N_216);
and U7663 (N_7663,N_2793,N_360);
xor U7664 (N_7664,N_4146,N_5745);
xnor U7665 (N_7665,N_111,N_852);
nor U7666 (N_7666,N_3379,N_5753);
xor U7667 (N_7667,N_4140,N_2004);
nor U7668 (N_7668,N_1746,N_1324);
or U7669 (N_7669,N_5466,N_1133);
or U7670 (N_7670,N_3258,N_5626);
nor U7671 (N_7671,N_4795,N_3881);
xor U7672 (N_7672,N_282,N_242);
xnor U7673 (N_7673,N_4435,N_5664);
and U7674 (N_7674,N_2096,N_5480);
or U7675 (N_7675,N_5311,N_516);
and U7676 (N_7676,N_358,N_648);
or U7677 (N_7677,N_4612,N_273);
xnor U7678 (N_7678,N_606,N_119);
xnor U7679 (N_7679,N_3395,N_4889);
xor U7680 (N_7680,N_3764,N_5832);
or U7681 (N_7681,N_2562,N_5251);
xnor U7682 (N_7682,N_1519,N_5222);
xnor U7683 (N_7683,N_5781,N_1745);
xnor U7684 (N_7684,N_3355,N_5521);
or U7685 (N_7685,N_3761,N_809);
nand U7686 (N_7686,N_4473,N_4318);
xor U7687 (N_7687,N_177,N_5018);
and U7688 (N_7688,N_364,N_1741);
xnor U7689 (N_7689,N_1107,N_5722);
nor U7690 (N_7690,N_4231,N_4853);
and U7691 (N_7691,N_133,N_1747);
nor U7692 (N_7692,N_1069,N_909);
and U7693 (N_7693,N_3680,N_677);
and U7694 (N_7694,N_3369,N_5397);
xnor U7695 (N_7695,N_1988,N_4933);
and U7696 (N_7696,N_5318,N_94);
and U7697 (N_7697,N_4527,N_2778);
or U7698 (N_7698,N_4484,N_2754);
or U7699 (N_7699,N_4708,N_2787);
nor U7700 (N_7700,N_406,N_3467);
xor U7701 (N_7701,N_2185,N_4493);
xor U7702 (N_7702,N_5523,N_5772);
nand U7703 (N_7703,N_158,N_1179);
and U7704 (N_7704,N_4906,N_4447);
or U7705 (N_7705,N_1750,N_5505);
nor U7706 (N_7706,N_3786,N_1249);
or U7707 (N_7707,N_4574,N_3961);
nand U7708 (N_7708,N_3049,N_5568);
nor U7709 (N_7709,N_4845,N_3702);
or U7710 (N_7710,N_569,N_778);
and U7711 (N_7711,N_199,N_2676);
nand U7712 (N_7712,N_2474,N_5323);
and U7713 (N_7713,N_5878,N_2063);
and U7714 (N_7714,N_4660,N_1109);
xor U7715 (N_7715,N_1158,N_4881);
and U7716 (N_7716,N_3231,N_1036);
nand U7717 (N_7717,N_143,N_3999);
nand U7718 (N_7718,N_2773,N_3301);
or U7719 (N_7719,N_1014,N_4394);
or U7720 (N_7720,N_2806,N_18);
xor U7721 (N_7721,N_4366,N_125);
nor U7722 (N_7722,N_1389,N_3803);
nand U7723 (N_7723,N_928,N_5252);
xnor U7724 (N_7724,N_829,N_375);
and U7725 (N_7725,N_4813,N_670);
nor U7726 (N_7726,N_1164,N_1506);
nor U7727 (N_7727,N_4766,N_3844);
nor U7728 (N_7728,N_2241,N_4815);
nand U7729 (N_7729,N_4522,N_4689);
and U7730 (N_7730,N_5654,N_4515);
nor U7731 (N_7731,N_4012,N_5336);
nand U7732 (N_7732,N_4274,N_2634);
nand U7733 (N_7733,N_4445,N_634);
nor U7734 (N_7734,N_58,N_2719);
xor U7735 (N_7735,N_307,N_4785);
nand U7736 (N_7736,N_5126,N_5974);
or U7737 (N_7737,N_5498,N_5882);
or U7738 (N_7738,N_2346,N_3901);
nand U7739 (N_7739,N_3115,N_3855);
or U7740 (N_7740,N_1526,N_3121);
xnor U7741 (N_7741,N_2989,N_4414);
xor U7742 (N_7742,N_175,N_464);
or U7743 (N_7743,N_4165,N_5455);
xor U7744 (N_7744,N_5783,N_2779);
xor U7745 (N_7745,N_1153,N_2092);
nor U7746 (N_7746,N_5156,N_2652);
and U7747 (N_7747,N_5160,N_3563);
nand U7748 (N_7748,N_5032,N_1865);
nand U7749 (N_7749,N_5543,N_1445);
and U7750 (N_7750,N_3697,N_3716);
and U7751 (N_7751,N_1352,N_336);
and U7752 (N_7752,N_2926,N_5612);
or U7753 (N_7753,N_5049,N_2599);
or U7754 (N_7754,N_5847,N_2938);
xnor U7755 (N_7755,N_363,N_3440);
nand U7756 (N_7756,N_3805,N_4481);
and U7757 (N_7757,N_5989,N_2341);
nor U7758 (N_7758,N_4794,N_3947);
nand U7759 (N_7759,N_4272,N_958);
nand U7760 (N_7760,N_352,N_2757);
nor U7761 (N_7761,N_3857,N_1473);
and U7762 (N_7762,N_711,N_4971);
xor U7763 (N_7763,N_1846,N_757);
nand U7764 (N_7764,N_3916,N_517);
nand U7765 (N_7765,N_1270,N_4822);
and U7766 (N_7766,N_2106,N_5058);
or U7767 (N_7767,N_4698,N_5403);
and U7768 (N_7768,N_4974,N_3089);
or U7769 (N_7769,N_21,N_1124);
nor U7770 (N_7770,N_972,N_5946);
xnor U7771 (N_7771,N_710,N_4062);
xnor U7772 (N_7772,N_5763,N_4043);
xnor U7773 (N_7773,N_2,N_1759);
xnor U7774 (N_7774,N_1790,N_4228);
and U7775 (N_7775,N_4915,N_5007);
or U7776 (N_7776,N_5089,N_2141);
and U7777 (N_7777,N_1193,N_498);
and U7778 (N_7778,N_168,N_4334);
or U7779 (N_7779,N_5652,N_3799);
nor U7780 (N_7780,N_4263,N_931);
nand U7781 (N_7781,N_5544,N_600);
nand U7782 (N_7782,N_2457,N_105);
nor U7783 (N_7783,N_2775,N_3490);
xor U7784 (N_7784,N_5914,N_1875);
nand U7785 (N_7785,N_3989,N_592);
or U7786 (N_7786,N_4798,N_2952);
or U7787 (N_7787,N_4576,N_900);
xor U7788 (N_7788,N_4137,N_3384);
nand U7789 (N_7789,N_1714,N_4594);
and U7790 (N_7790,N_3758,N_2064);
xnor U7791 (N_7791,N_5950,N_839);
nor U7792 (N_7792,N_4733,N_3642);
nand U7793 (N_7793,N_1656,N_430);
xor U7794 (N_7794,N_4716,N_1898);
or U7795 (N_7795,N_5644,N_4426);
nand U7796 (N_7796,N_57,N_4377);
xnor U7797 (N_7797,N_5114,N_5401);
and U7798 (N_7798,N_1923,N_2084);
or U7799 (N_7799,N_4842,N_4654);
nand U7800 (N_7800,N_2091,N_1312);
nand U7801 (N_7801,N_2739,N_988);
nand U7802 (N_7802,N_5134,N_3016);
or U7803 (N_7803,N_1907,N_5849);
or U7804 (N_7804,N_3302,N_3910);
and U7805 (N_7805,N_982,N_2590);
xnor U7806 (N_7806,N_971,N_3322);
xnor U7807 (N_7807,N_287,N_5526);
and U7808 (N_7808,N_2672,N_4402);
nor U7809 (N_7809,N_5412,N_1764);
and U7810 (N_7810,N_2794,N_4193);
and U7811 (N_7811,N_1598,N_5350);
and U7812 (N_7812,N_2990,N_4894);
and U7813 (N_7813,N_4926,N_3153);
nor U7814 (N_7814,N_1268,N_5338);
nand U7815 (N_7815,N_3853,N_4216);
nand U7816 (N_7816,N_1021,N_3370);
or U7817 (N_7817,N_3411,N_3375);
nor U7818 (N_7818,N_3956,N_1537);
and U7819 (N_7819,N_473,N_4186);
nor U7820 (N_7820,N_1413,N_3469);
xnor U7821 (N_7821,N_611,N_2594);
and U7822 (N_7822,N_3793,N_2274);
nor U7823 (N_7823,N_290,N_3244);
nand U7824 (N_7824,N_14,N_2178);
nor U7825 (N_7825,N_967,N_1291);
and U7826 (N_7826,N_1175,N_2900);
nor U7827 (N_7827,N_4135,N_4731);
nand U7828 (N_7828,N_2076,N_2414);
nor U7829 (N_7829,N_4735,N_5197);
or U7830 (N_7830,N_4235,N_1022);
xnor U7831 (N_7831,N_3975,N_5033);
nor U7832 (N_7832,N_2822,N_244);
and U7833 (N_7833,N_5499,N_3904);
and U7834 (N_7834,N_3103,N_3351);
or U7835 (N_7835,N_3707,N_3397);
xnor U7836 (N_7836,N_2960,N_3731);
or U7837 (N_7837,N_1657,N_4738);
nand U7838 (N_7838,N_4966,N_5931);
or U7839 (N_7839,N_2814,N_5422);
nor U7840 (N_7840,N_1755,N_5369);
or U7841 (N_7841,N_2324,N_825);
xor U7842 (N_7842,N_305,N_2584);
xnor U7843 (N_7843,N_5805,N_2395);
and U7844 (N_7844,N_1531,N_3736);
and U7845 (N_7845,N_1391,N_5408);
and U7846 (N_7846,N_560,N_4207);
xor U7847 (N_7847,N_1845,N_1055);
and U7848 (N_7848,N_2736,N_935);
and U7849 (N_7849,N_4387,N_758);
and U7850 (N_7850,N_5562,N_2664);
nand U7851 (N_7851,N_4148,N_3441);
nor U7852 (N_7852,N_1282,N_2586);
nor U7853 (N_7853,N_2697,N_3345);
nand U7854 (N_7854,N_16,N_4681);
nor U7855 (N_7855,N_112,N_5219);
nor U7856 (N_7856,N_727,N_669);
nor U7857 (N_7857,N_4722,N_79);
xnor U7858 (N_7858,N_1265,N_4528);
and U7859 (N_7859,N_3965,N_3249);
nand U7860 (N_7860,N_2448,N_765);
xor U7861 (N_7861,N_1414,N_2954);
nor U7862 (N_7862,N_2888,N_1936);
or U7863 (N_7863,N_3130,N_3864);
nand U7864 (N_7864,N_3953,N_1568);
xnor U7865 (N_7865,N_630,N_4418);
xor U7866 (N_7866,N_2442,N_2839);
nor U7867 (N_7867,N_2077,N_68);
nor U7868 (N_7868,N_1658,N_1904);
nor U7869 (N_7869,N_5225,N_5877);
nand U7870 (N_7870,N_5595,N_3640);
xnor U7871 (N_7871,N_3243,N_5837);
nand U7872 (N_7872,N_2631,N_167);
nor U7873 (N_7873,N_4625,N_4590);
nor U7874 (N_7874,N_4638,N_2957);
xnor U7875 (N_7875,N_2699,N_196);
nor U7876 (N_7876,N_4333,N_1100);
xor U7877 (N_7877,N_1921,N_3942);
nor U7878 (N_7878,N_1705,N_3718);
xnor U7879 (N_7879,N_5145,N_1726);
nand U7880 (N_7880,N_5672,N_3138);
or U7881 (N_7881,N_3278,N_297);
nor U7882 (N_7882,N_3213,N_5108);
or U7883 (N_7883,N_714,N_4309);
xor U7884 (N_7884,N_767,N_805);
nor U7885 (N_7885,N_4040,N_3267);
nand U7886 (N_7886,N_2201,N_2431);
nand U7887 (N_7887,N_705,N_3714);
nand U7888 (N_7888,N_1761,N_1236);
and U7889 (N_7889,N_3615,N_5352);
xor U7890 (N_7890,N_3090,N_396);
nor U7891 (N_7891,N_4583,N_4560);
nand U7892 (N_7892,N_3481,N_1178);
nand U7893 (N_7893,N_5669,N_4547);
nand U7894 (N_7894,N_373,N_3673);
and U7895 (N_7895,N_3977,N_884);
or U7896 (N_7896,N_1319,N_1723);
nand U7897 (N_7897,N_4736,N_2541);
and U7898 (N_7898,N_1292,N_5262);
nand U7899 (N_7899,N_4245,N_991);
and U7900 (N_7900,N_5780,N_2032);
and U7901 (N_7901,N_65,N_1730);
nor U7902 (N_7902,N_3025,N_2385);
xnor U7903 (N_7903,N_1636,N_3325);
xnor U7904 (N_7904,N_559,N_4283);
or U7905 (N_7905,N_2555,N_3547);
nor U7906 (N_7906,N_1840,N_3584);
nand U7907 (N_7907,N_4701,N_3410);
xnor U7908 (N_7908,N_1810,N_3365);
or U7909 (N_7909,N_4160,N_5885);
nor U7910 (N_7910,N_1630,N_2162);
and U7911 (N_7911,N_3199,N_2451);
or U7912 (N_7912,N_4452,N_2169);
nor U7913 (N_7913,N_5899,N_469);
nand U7914 (N_7914,N_5406,N_2136);
and U7915 (N_7915,N_5282,N_3472);
and U7916 (N_7916,N_50,N_672);
xnor U7917 (N_7917,N_1971,N_1072);
or U7918 (N_7918,N_2628,N_3759);
nand U7919 (N_7919,N_2867,N_1903);
nand U7920 (N_7920,N_752,N_3142);
nor U7921 (N_7921,N_855,N_1503);
and U7922 (N_7922,N_2591,N_676);
nor U7923 (N_7923,N_653,N_2182);
or U7924 (N_7924,N_3690,N_1608);
nand U7925 (N_7925,N_4444,N_3084);
nor U7926 (N_7926,N_764,N_4441);
xor U7927 (N_7927,N_4809,N_3654);
and U7928 (N_7928,N_5870,N_2340);
nor U7929 (N_7929,N_5253,N_1593);
nor U7930 (N_7930,N_5109,N_4499);
or U7931 (N_7931,N_5610,N_3139);
or U7932 (N_7932,N_707,N_333);
nand U7933 (N_7933,N_4634,N_4415);
xor U7934 (N_7934,N_662,N_4987);
nand U7935 (N_7935,N_2983,N_547);
nand U7936 (N_7936,N_4181,N_3430);
and U7937 (N_7937,N_3342,N_5146);
nor U7938 (N_7938,N_3336,N_5070);
and U7939 (N_7939,N_3637,N_431);
or U7940 (N_7940,N_1661,N_5153);
xor U7941 (N_7941,N_2909,N_1075);
or U7942 (N_7942,N_340,N_2578);
nor U7943 (N_7943,N_5386,N_1364);
nor U7944 (N_7944,N_5012,N_2499);
and U7945 (N_7945,N_2583,N_3927);
nor U7946 (N_7946,N_4567,N_2855);
or U7947 (N_7947,N_2202,N_5755);
nor U7948 (N_7948,N_934,N_783);
xor U7949 (N_7949,N_2072,N_2689);
nor U7950 (N_7950,N_5515,N_1041);
xor U7951 (N_7951,N_1024,N_1599);
nor U7952 (N_7952,N_2597,N_2582);
xnor U7953 (N_7953,N_4890,N_3204);
nand U7954 (N_7954,N_4321,N_3478);
or U7955 (N_7955,N_1744,N_1830);
nand U7956 (N_7956,N_2977,N_5445);
and U7957 (N_7957,N_3372,N_1204);
and U7958 (N_7958,N_1023,N_531);
nor U7959 (N_7959,N_3683,N_4082);
xnor U7960 (N_7960,N_2250,N_3840);
xnor U7961 (N_7961,N_1221,N_2777);
nand U7962 (N_7962,N_2497,N_1438);
xor U7963 (N_7963,N_1299,N_4963);
or U7964 (N_7964,N_3374,N_2986);
or U7965 (N_7965,N_3123,N_2440);
xor U7966 (N_7966,N_5173,N_656);
nor U7967 (N_7967,N_746,N_4042);
nor U7968 (N_7968,N_3307,N_2661);
nand U7969 (N_7969,N_4396,N_1009);
nand U7970 (N_7970,N_5897,N_3294);
and U7971 (N_7971,N_1406,N_3091);
nor U7972 (N_7972,N_1555,N_2844);
nor U7973 (N_7973,N_901,N_827);
and U7974 (N_7974,N_106,N_820);
xor U7975 (N_7975,N_5578,N_5936);
and U7976 (N_7976,N_1233,N_4657);
or U7977 (N_7977,N_588,N_3466);
nand U7978 (N_7978,N_275,N_2234);
nor U7979 (N_7979,N_1631,N_5287);
or U7980 (N_7980,N_578,N_3299);
xnor U7981 (N_7981,N_3112,N_466);
nand U7982 (N_7982,N_4495,N_2377);
nand U7983 (N_7983,N_2453,N_272);
xnor U7984 (N_7984,N_4695,N_749);
or U7985 (N_7985,N_3982,N_1362);
xnor U7986 (N_7986,N_4132,N_3118);
xor U7987 (N_7987,N_1026,N_2044);
nor U7988 (N_7988,N_1208,N_5704);
and U7989 (N_7989,N_3726,N_4891);
nor U7990 (N_7990,N_593,N_5009);
nand U7991 (N_7991,N_4760,N_2267);
and U7992 (N_7992,N_3766,N_2905);
or U7993 (N_7993,N_3734,N_3283);
nor U7994 (N_7994,N_3392,N_3201);
nand U7995 (N_7995,N_3337,N_4433);
or U7996 (N_7996,N_1065,N_4289);
nand U7997 (N_7997,N_2593,N_4606);
and U7998 (N_7998,N_5846,N_2502);
nand U7999 (N_7999,N_2000,N_4247);
nand U8000 (N_8000,N_3079,N_3781);
or U8001 (N_8001,N_2931,N_2788);
and U8002 (N_8002,N_3310,N_329);
nand U8003 (N_8003,N_2117,N_2813);
xnor U8004 (N_8004,N_5425,N_3567);
xor U8005 (N_8005,N_3380,N_4471);
or U8006 (N_8006,N_1339,N_2507);
and U8007 (N_8007,N_5586,N_184);
or U8008 (N_8008,N_5822,N_5732);
nand U8009 (N_8009,N_5393,N_1185);
nor U8010 (N_8010,N_5475,N_4018);
xnor U8011 (N_8011,N_5739,N_3938);
nor U8012 (N_8012,N_110,N_4691);
nand U8013 (N_8013,N_4572,N_4619);
nor U8014 (N_8014,N_3772,N_2875);
nand U8015 (N_8015,N_3191,N_2352);
xor U8016 (N_8016,N_2817,N_3099);
or U8017 (N_8017,N_2078,N_3008);
and U8018 (N_8018,N_1679,N_797);
nor U8019 (N_8019,N_2030,N_1286);
and U8020 (N_8020,N_2748,N_1681);
or U8021 (N_8021,N_3326,N_3681);
nor U8022 (N_8022,N_5530,N_5103);
xor U8023 (N_8023,N_3197,N_992);
nand U8024 (N_8024,N_5366,N_804);
xnor U8025 (N_8025,N_278,N_1866);
xor U8026 (N_8026,N_1154,N_3818);
and U8027 (N_8027,N_4331,N_5619);
xnor U8028 (N_8028,N_5062,N_129);
nor U8029 (N_8029,N_1809,N_3924);
xor U8030 (N_8030,N_222,N_5726);
and U8031 (N_8031,N_3311,N_2923);
or U8032 (N_8032,N_4997,N_4679);
and U8033 (N_8033,N_595,N_1823);
nor U8034 (N_8034,N_4389,N_4201);
and U8035 (N_8035,N_4607,N_5215);
nand U8036 (N_8036,N_911,N_3741);
or U8037 (N_8037,N_5378,N_5065);
nand U8038 (N_8038,N_3353,N_2677);
xor U8039 (N_8039,N_4218,N_1896);
xnor U8040 (N_8040,N_2911,N_5711);
nor U8041 (N_8041,N_3987,N_5453);
or U8042 (N_8042,N_3400,N_2852);
nor U8043 (N_8043,N_201,N_5293);
xnor U8044 (N_8044,N_5442,N_5841);
xor U8045 (N_8045,N_2704,N_2005);
nand U8046 (N_8046,N_5027,N_227);
and U8047 (N_8047,N_2713,N_5970);
xnor U8048 (N_8048,N_580,N_274);
and U8049 (N_8049,N_4051,N_5579);
or U8050 (N_8050,N_1772,N_4101);
nand U8051 (N_8051,N_1081,N_1699);
and U8052 (N_8052,N_4472,N_2882);
and U8053 (N_8053,N_5775,N_5567);
or U8054 (N_8054,N_1979,N_4382);
nand U8055 (N_8055,N_708,N_1104);
nor U8056 (N_8056,N_2109,N_2210);
xnor U8057 (N_8057,N_1783,N_2756);
or U8058 (N_8058,N_1359,N_4234);
nor U8059 (N_8059,N_2783,N_3504);
nand U8060 (N_8060,N_37,N_337);
nand U8061 (N_8061,N_3866,N_2214);
nand U8062 (N_8062,N_1460,N_2505);
or U8063 (N_8063,N_2551,N_5447);
xor U8064 (N_8064,N_1115,N_4932);
and U8065 (N_8065,N_3937,N_1985);
nor U8066 (N_8066,N_5481,N_266);
xor U8067 (N_8067,N_4507,N_4260);
xnor U8068 (N_8068,N_5319,N_138);
xnor U8069 (N_8069,N_5980,N_5452);
nor U8070 (N_8070,N_188,N_1335);
nand U8071 (N_8071,N_3104,N_5977);
nor U8072 (N_8072,N_5740,N_4998);
or U8073 (N_8073,N_4013,N_5086);
nand U8074 (N_8074,N_5327,N_2183);
or U8075 (N_8075,N_3164,N_1581);
nand U8076 (N_8076,N_4345,N_3241);
nor U8077 (N_8077,N_4328,N_5895);
and U8078 (N_8078,N_2918,N_2357);
xnor U8079 (N_8079,N_3111,N_1415);
xor U8080 (N_8080,N_2953,N_2843);
xor U8081 (N_8081,N_1829,N_4206);
xnor U8082 (N_8082,N_29,N_505);
or U8083 (N_8083,N_2509,N_5593);
and U8084 (N_8084,N_987,N_1053);
and U8085 (N_8085,N_3891,N_1786);
nor U8086 (N_8086,N_4298,N_3610);
or U8087 (N_8087,N_4365,N_5887);
or U8088 (N_8088,N_774,N_160);
nand U8089 (N_8089,N_849,N_2257);
and U8090 (N_8090,N_2665,N_3959);
nor U8091 (N_8091,N_817,N_3543);
or U8092 (N_8092,N_2755,N_4850);
xor U8093 (N_8093,N_2027,N_5216);
or U8094 (N_8094,N_4096,N_626);
nor U8095 (N_8095,N_4219,N_4921);
xnor U8096 (N_8096,N_223,N_4302);
or U8097 (N_8097,N_1623,N_5982);
xnor U8098 (N_8098,N_2424,N_3083);
or U8099 (N_8099,N_5078,N_5123);
and U8100 (N_8100,N_5951,N_5608);
nor U8101 (N_8101,N_485,N_1559);
nand U8102 (N_8102,N_5164,N_1616);
nand U8103 (N_8103,N_3771,N_4818);
or U8104 (N_8104,N_5606,N_2338);
xnor U8105 (N_8105,N_4597,N_4337);
xnor U8106 (N_8106,N_139,N_436);
and U8107 (N_8107,N_4802,N_2446);
nor U8108 (N_8108,N_2339,N_4734);
and U8109 (N_8109,N_5731,N_3549);
xnor U8110 (N_8110,N_544,N_3909);
xnor U8111 (N_8111,N_5705,N_5272);
and U8112 (N_8112,N_2815,N_5793);
or U8113 (N_8113,N_5973,N_3265);
or U8114 (N_8114,N_1596,N_2073);
xor U8115 (N_8115,N_2567,N_2403);
nand U8116 (N_8116,N_4955,N_2156);
or U8117 (N_8117,N_2256,N_1876);
or U8118 (N_8118,N_4088,N_2546);
nand U8119 (N_8119,N_2871,N_4074);
nand U8120 (N_8120,N_1315,N_2020);
nand U8121 (N_8121,N_5986,N_5312);
or U8122 (N_8122,N_1271,N_4420);
or U8123 (N_8123,N_5729,N_5095);
and U8124 (N_8124,N_371,N_2769);
nor U8125 (N_8125,N_3993,N_3068);
xnor U8126 (N_8126,N_88,N_3135);
or U8127 (N_8127,N_4754,N_3470);
nor U8128 (N_8128,N_4856,N_4147);
and U8129 (N_8129,N_5080,N_4978);
or U8130 (N_8130,N_4009,N_4582);
xor U8131 (N_8131,N_1571,N_3180);
nor U8132 (N_8132,N_4224,N_1566);
nor U8133 (N_8133,N_3542,N_4712);
nand U8134 (N_8134,N_3189,N_3645);
xor U8135 (N_8135,N_999,N_2487);
or U8136 (N_8136,N_5859,N_3883);
or U8137 (N_8137,N_895,N_484);
nor U8138 (N_8138,N_1013,N_5864);
or U8139 (N_8139,N_2046,N_4303);
or U8140 (N_8140,N_1138,N_1673);
xor U8141 (N_8141,N_5332,N_1877);
xnor U8142 (N_8142,N_789,N_5055);
xor U8143 (N_8143,N_440,N_1948);
xnor U8144 (N_8144,N_891,N_2645);
and U8145 (N_8145,N_1769,N_4372);
xor U8146 (N_8146,N_1384,N_293);
xnor U8147 (N_8147,N_3157,N_1813);
nand U8148 (N_8148,N_2862,N_1);
xor U8149 (N_8149,N_3019,N_2437);
or U8150 (N_8150,N_998,N_5991);
nand U8151 (N_8151,N_5820,N_3445);
and U8152 (N_8152,N_1160,N_259);
and U8153 (N_8153,N_3238,N_1121);
nor U8154 (N_8154,N_3391,N_1624);
xor U8155 (N_8155,N_4863,N_573);
xor U8156 (N_8156,N_32,N_3630);
nand U8157 (N_8157,N_3616,N_2639);
nand U8158 (N_8158,N_1721,N_5577);
nand U8159 (N_8159,N_1325,N_3192);
xnor U8160 (N_8160,N_2941,N_4469);
xnor U8161 (N_8161,N_4531,N_5167);
nand U8162 (N_8162,N_3651,N_1992);
nand U8163 (N_8163,N_2834,N_3652);
xnor U8164 (N_8164,N_841,N_426);
nor U8165 (N_8165,N_3363,N_1064);
xor U8166 (N_8166,N_4320,N_338);
and U8167 (N_8167,N_2784,N_2350);
nor U8168 (N_8168,N_1102,N_1136);
or U8169 (N_8169,N_4552,N_5853);
xor U8170 (N_8170,N_2111,N_84);
nand U8171 (N_8171,N_3425,N_2856);
nor U8172 (N_8172,N_3420,N_250);
or U8173 (N_8173,N_1038,N_2958);
and U8174 (N_8174,N_2668,N_654);
nor U8175 (N_8175,N_245,N_1905);
or U8176 (N_8176,N_2075,N_2557);
and U8177 (N_8177,N_5671,N_5534);
xnor U8178 (N_8178,N_4661,N_3609);
xnor U8179 (N_8179,N_2055,N_3580);
xor U8180 (N_8180,N_4187,N_339);
or U8181 (N_8181,N_5539,N_821);
xnor U8182 (N_8182,N_1901,N_2400);
and U8183 (N_8183,N_780,N_4740);
xor U8184 (N_8184,N_2079,N_3282);
xor U8185 (N_8185,N_745,N_1030);
and U8186 (N_8186,N_1943,N_2319);
or U8187 (N_8187,N_2420,N_3612);
and U8188 (N_8188,N_2992,N_1477);
xor U8189 (N_8189,N_1256,N_5437);
and U8190 (N_8190,N_488,N_3492);
xnor U8191 (N_8191,N_2432,N_3253);
nor U8192 (N_8192,N_4049,N_879);
nor U8193 (N_8193,N_2280,N_1880);
nand U8194 (N_8194,N_1638,N_3438);
or U8195 (N_8195,N_4637,N_734);
and U8196 (N_8196,N_3949,N_4029);
nor U8197 (N_8197,N_5006,N_1246);
xnor U8198 (N_8198,N_5646,N_2317);
nor U8199 (N_8199,N_2137,N_4546);
nand U8200 (N_8200,N_4717,N_3863);
and U8201 (N_8201,N_5209,N_614);
or U8202 (N_8202,N_5830,N_5294);
nand U8203 (N_8203,N_232,N_5624);
or U8204 (N_8204,N_4306,N_5467);
nor U8205 (N_8205,N_5411,N_1411);
or U8206 (N_8206,N_5472,N_5469);
xor U8207 (N_8207,N_1336,N_1229);
or U8208 (N_8208,N_4239,N_2939);
and U8209 (N_8209,N_202,N_5541);
nand U8210 (N_8210,N_673,N_257);
or U8211 (N_8211,N_4992,N_500);
nor U8212 (N_8212,N_4087,N_2762);
nand U8213 (N_8213,N_2724,N_3074);
nand U8214 (N_8214,N_435,N_2175);
xor U8215 (N_8215,N_1703,N_3046);
xor U8216 (N_8216,N_4803,N_5341);
or U8217 (N_8217,N_251,N_5402);
or U8218 (N_8218,N_2251,N_369);
and U8219 (N_8219,N_1860,N_2047);
nor U8220 (N_8220,N_3945,N_1101);
nand U8221 (N_8221,N_2177,N_1198);
xor U8222 (N_8222,N_5202,N_4570);
xnor U8223 (N_8223,N_2874,N_2774);
nand U8224 (N_8224,N_584,N_5687);
xor U8225 (N_8225,N_2870,N_2899);
xor U8226 (N_8226,N_1394,N_665);
nand U8227 (N_8227,N_54,N_4188);
and U8228 (N_8228,N_2213,N_3919);
xnor U8229 (N_8229,N_4144,N_447);
nor U8230 (N_8230,N_1884,N_4952);
nand U8231 (N_8231,N_591,N_5808);
and U8232 (N_8232,N_2627,N_4150);
or U8233 (N_8233,N_33,N_1123);
and U8234 (N_8234,N_1461,N_5100);
nand U8235 (N_8235,N_5655,N_4945);
nand U8236 (N_8236,N_2708,N_667);
xnor U8237 (N_8237,N_1228,N_1648);
nand U8238 (N_8238,N_3225,N_4111);
xnor U8239 (N_8239,N_2218,N_1977);
nor U8240 (N_8240,N_1388,N_2189);
and U8241 (N_8241,N_45,N_1805);
or U8242 (N_8242,N_4835,N_2293);
nand U8243 (N_8243,N_4562,N_5385);
nor U8244 (N_8244,N_4315,N_1946);
and U8245 (N_8245,N_319,N_2964);
nor U8246 (N_8246,N_5588,N_5436);
xnor U8247 (N_8247,N_1366,N_5090);
nand U8248 (N_8248,N_4557,N_312);
nor U8249 (N_8249,N_860,N_2519);
and U8250 (N_8250,N_174,N_354);
nand U8251 (N_8251,N_3171,N_5474);
xor U8252 (N_8252,N_1279,N_1640);
nand U8253 (N_8253,N_1789,N_756);
and U8254 (N_8254,N_4213,N_3092);
xnor U8255 (N_8255,N_5245,N_3918);
or U8256 (N_8256,N_898,N_5231);
xnor U8257 (N_8257,N_2980,N_1094);
nand U8258 (N_8258,N_4651,N_23);
nor U8259 (N_8259,N_4719,N_5620);
nor U8260 (N_8260,N_2103,N_938);
and U8261 (N_8261,N_2211,N_3870);
nand U8262 (N_8262,N_5941,N_5810);
and U8263 (N_8263,N_261,N_3450);
xnor U8264 (N_8264,N_4982,N_1350);
nor U8265 (N_8265,N_1025,N_5263);
and U8266 (N_8266,N_1573,N_1668);
xor U8267 (N_8267,N_5187,N_5658);
and U8268 (N_8268,N_5667,N_3205);
or U8269 (N_8269,N_585,N_2830);
nor U8270 (N_8270,N_1962,N_1617);
and U8271 (N_8271,N_4909,N_1916);
nand U8272 (N_8272,N_3166,N_1678);
nand U8273 (N_8273,N_3187,N_4970);
nor U8274 (N_8274,N_5399,N_864);
and U8275 (N_8275,N_1695,N_4112);
or U8276 (N_8276,N_1165,N_1446);
nand U8277 (N_8277,N_1820,N_5527);
xnor U8278 (N_8278,N_3885,N_1955);
xnor U8279 (N_8279,N_2003,N_114);
or U8280 (N_8280,N_2040,N_3724);
xor U8281 (N_8281,N_1435,N_5142);
xor U8282 (N_8282,N_1939,N_2207);
nand U8283 (N_8283,N_4223,N_4878);
nor U8284 (N_8284,N_978,N_330);
and U8285 (N_8285,N_1117,N_5760);
or U8286 (N_8286,N_5590,N_4820);
and U8287 (N_8287,N_513,N_4236);
xnor U8288 (N_8288,N_4329,N_3012);
nor U8289 (N_8289,N_2934,N_4461);
nor U8290 (N_8290,N_4151,N_4494);
nor U8291 (N_8291,N_1976,N_3826);
nor U8292 (N_8292,N_4769,N_3033);
xor U8293 (N_8293,N_2812,N_2743);
xor U8294 (N_8294,N_4084,N_2022);
nand U8295 (N_8295,N_1495,N_617);
nand U8296 (N_8296,N_1731,N_455);
nand U8297 (N_8297,N_574,N_5069);
and U8298 (N_8298,N_3398,N_867);
nand U8299 (N_8299,N_5129,N_1719);
or U8300 (N_8300,N_5892,N_4250);
nor U8301 (N_8301,N_1937,N_3399);
and U8302 (N_8302,N_1057,N_883);
or U8303 (N_8303,N_4801,N_1145);
nor U8304 (N_8304,N_2454,N_4270);
nor U8305 (N_8305,N_3300,N_1106);
xnor U8306 (N_8306,N_2799,N_4304);
and U8307 (N_8307,N_2759,N_5737);
xor U8308 (N_8308,N_5097,N_2796);
xor U8309 (N_8309,N_2801,N_2879);
or U8310 (N_8310,N_1869,N_2259);
and U8311 (N_8311,N_609,N_4524);
or U8312 (N_8312,N_3239,N_3281);
and U8313 (N_8313,N_3489,N_5957);
nand U8314 (N_8314,N_2333,N_4348);
nor U8315 (N_8315,N_5649,N_247);
and U8316 (N_8316,N_1459,N_2498);
nor U8317 (N_8317,N_5269,N_5816);
nor U8318 (N_8318,N_5712,N_1367);
xor U8319 (N_8319,N_285,N_1197);
or U8320 (N_8320,N_2902,N_5851);
and U8321 (N_8321,N_2685,N_5814);
nor U8322 (N_8322,N_28,N_3829);
and U8323 (N_8323,N_1892,N_359);
or U8324 (N_8324,N_3713,N_1409);
and U8325 (N_8325,N_539,N_2907);
nor U8326 (N_8326,N_1952,N_3247);
nor U8327 (N_8327,N_2529,N_2927);
or U8328 (N_8328,N_3229,N_397);
nand U8329 (N_8329,N_97,N_5302);
nand U8330 (N_8330,N_5189,N_3066);
nand U8331 (N_8331,N_1485,N_2727);
or U8332 (N_8332,N_3658,N_3525);
xnor U8333 (N_8333,N_2670,N_1601);
or U8334 (N_8334,N_2614,N_51);
and U8335 (N_8335,N_2526,N_1159);
or U8336 (N_8336,N_2252,N_877);
nand U8337 (N_8337,N_458,N_4196);
or U8338 (N_8338,N_3257,N_830);
and U8339 (N_8339,N_2846,N_1137);
or U8340 (N_8340,N_3573,N_5907);
and U8341 (N_8341,N_2539,N_3233);
or U8342 (N_8342,N_5150,N_5317);
nand U8343 (N_8343,N_3087,N_5373);
nor U8344 (N_8344,N_5322,N_3851);
or U8345 (N_8345,N_553,N_2906);
xnor U8346 (N_8346,N_3756,N_781);
xor U8347 (N_8347,N_2199,N_1712);
nor U8348 (N_8348,N_4761,N_792);
and U8349 (N_8349,N_3749,N_4322);
or U8350 (N_8350,N_3093,N_4854);
nor U8351 (N_8351,N_4035,N_957);
or U8352 (N_8352,N_2427,N_663);
or U8353 (N_8353,N_4020,N_127);
xor U8354 (N_8354,N_5771,N_4565);
xor U8355 (N_8355,N_5631,N_1970);
or U8356 (N_8356,N_5954,N_3552);
nor U8357 (N_8357,N_5226,N_3606);
nor U8358 (N_8358,N_2011,N_4650);
and U8359 (N_8359,N_1226,N_1590);
nor U8360 (N_8360,N_3429,N_2999);
or U8361 (N_8361,N_5271,N_2903);
xnor U8362 (N_8362,N_4248,N_2099);
or U8363 (N_8363,N_5559,N_3538);
nor U8364 (N_8364,N_1405,N_2971);
nor U8365 (N_8365,N_1033,N_3807);
and U8366 (N_8366,N_1402,N_4763);
xnor U8367 (N_8367,N_48,N_875);
nand U8368 (N_8368,N_5067,N_3279);
and U8369 (N_8369,N_5141,N_5570);
nor U8370 (N_8370,N_1504,N_1666);
xor U8371 (N_8371,N_5502,N_2554);
nand U8372 (N_8372,N_5641,N_5547);
xnor U8373 (N_8373,N_1849,N_1918);
xor U8374 (N_8374,N_349,N_441);
or U8375 (N_8375,N_2622,N_704);
nand U8376 (N_8376,N_3296,N_2204);
nand U8377 (N_8377,N_181,N_4758);
or U8378 (N_8378,N_1545,N_2396);
or U8379 (N_8379,N_3248,N_5845);
and U8380 (N_8380,N_5337,N_2229);
nor U8381 (N_8381,N_1139,N_1645);
nor U8382 (N_8382,N_5013,N_4064);
and U8383 (N_8383,N_5653,N_3655);
and U8384 (N_8384,N_2547,N_279);
and U8385 (N_8385,N_3126,N_4632);
xnor U8386 (N_8386,N_5343,N_1964);
or U8387 (N_8387,N_3858,N_2356);
nand U8388 (N_8388,N_575,N_4523);
or U8389 (N_8389,N_2310,N_5348);
xnor U8390 (N_8390,N_2345,N_89);
and U8391 (N_8391,N_3335,N_124);
xor U8392 (N_8392,N_4577,N_4421);
nand U8393 (N_8393,N_3809,N_1834);
and U8394 (N_8394,N_1777,N_2060);
nor U8395 (N_8395,N_1457,N_132);
nand U8396 (N_8396,N_3359,N_4106);
xnor U8397 (N_8397,N_1466,N_1954);
xor U8398 (N_8398,N_2536,N_5928);
and U8399 (N_8399,N_4514,N_376);
or U8400 (N_8400,N_4788,N_3149);
nor U8401 (N_8401,N_3386,N_85);
nor U8402 (N_8402,N_499,N_2942);
xor U8403 (N_8403,N_1051,N_1619);
xor U8404 (N_8404,N_4639,N_5330);
nand U8405 (N_8405,N_4812,N_3920);
nand U8406 (N_8406,N_4050,N_2974);
nor U8407 (N_8407,N_5903,N_2821);
nand U8408 (N_8408,N_2425,N_3728);
xnor U8409 (N_8409,N_2728,N_3708);
or U8410 (N_8410,N_1500,N_833);
nor U8411 (N_8411,N_4438,N_4475);
nor U8412 (N_8412,N_2415,N_1704);
nor U8413 (N_8413,N_1403,N_4288);
and U8414 (N_8414,N_5758,N_1527);
or U8415 (N_8415,N_2533,N_3820);
and U8416 (N_8416,N_4338,N_897);
xor U8417 (N_8417,N_699,N_25);
or U8418 (N_8418,N_4525,N_876);
or U8419 (N_8419,N_398,N_4936);
nor U8420 (N_8420,N_5435,N_1600);
xor U8421 (N_8421,N_1374,N_34);
and U8422 (N_8422,N_2173,N_709);
and U8423 (N_8423,N_5106,N_5752);
xor U8424 (N_8424,N_3415,N_2025);
nor U8425 (N_8425,N_288,N_468);
nand U8426 (N_8426,N_5345,N_5555);
and U8427 (N_8427,N_1760,N_1533);
nand U8428 (N_8428,N_2711,N_4678);
nor U8429 (N_8429,N_3692,N_5243);
nor U8430 (N_8430,N_1040,N_4267);
nand U8431 (N_8431,N_5613,N_2294);
and U8432 (N_8432,N_2543,N_5389);
nor U8433 (N_8433,N_1682,N_2258);
nor U8434 (N_8434,N_3668,N_5546);
or U8435 (N_8435,N_4559,N_4669);
nand U8436 (N_8436,N_3315,N_5428);
nor U8437 (N_8437,N_3861,N_4386);
nand U8438 (N_8438,N_1068,N_439);
and U8439 (N_8439,N_4786,N_4861);
xnor U8440 (N_8440,N_2643,N_3291);
nor U8441 (N_8441,N_1337,N_2018);
and U8442 (N_8442,N_2166,N_4817);
xor U8443 (N_8443,N_4102,N_4989);
or U8444 (N_8444,N_5769,N_4872);
or U8445 (N_8445,N_2716,N_342);
nor U8446 (N_8446,N_4628,N_5979);
and U8447 (N_8447,N_448,N_1211);
nand U8448 (N_8448,N_1430,N_3890);
nor U8449 (N_8449,N_2477,N_4375);
or U8450 (N_8450,N_5329,N_1529);
or U8451 (N_8451,N_1713,N_4214);
or U8452 (N_8452,N_5528,N_5087);
nor U8453 (N_8453,N_1259,N_4327);
or U8454 (N_8454,N_5280,N_2043);
xor U8455 (N_8455,N_5844,N_2494);
xnor U8456 (N_8456,N_3433,N_4621);
or U8457 (N_8457,N_3568,N_2608);
nor U8458 (N_8458,N_641,N_3983);
and U8459 (N_8459,N_4244,N_3867);
or U8460 (N_8460,N_5244,N_4237);
or U8461 (N_8461,N_5718,N_3096);
and U8462 (N_8462,N_2036,N_4045);
and U8463 (N_8463,N_154,N_2735);
nand U8464 (N_8464,N_1486,N_198);
or U8465 (N_8465,N_345,N_2342);
xnor U8466 (N_8466,N_1054,N_1416);
nand U8467 (N_8467,N_1118,N_2920);
nor U8468 (N_8468,N_4622,N_5905);
and U8469 (N_8469,N_819,N_3364);
nor U8470 (N_8470,N_2007,N_2522);
nand U8471 (N_8471,N_2300,N_5901);
xnor U8472 (N_8472,N_1774,N_2281);
nand U8473 (N_8473,N_1615,N_2491);
and U8474 (N_8474,N_2452,N_1194);
xnor U8475 (N_8475,N_3635,N_1873);
and U8476 (N_8476,N_845,N_2194);
or U8477 (N_8477,N_1899,N_454);
xnor U8478 (N_8478,N_4504,N_3010);
xor U8479 (N_8479,N_3907,N_386);
nand U8480 (N_8480,N_5889,N_3624);
nor U8481 (N_8481,N_695,N_2372);
nor U8482 (N_8482,N_4748,N_5256);
or U8483 (N_8483,N_1739,N_1483);
xnor U8484 (N_8484,N_331,N_2328);
nor U8485 (N_8485,N_1347,N_2123);
nand U8486 (N_8486,N_24,N_5240);
nand U8487 (N_8487,N_5234,N_70);
nand U8488 (N_8488,N_5632,N_700);
nor U8489 (N_8489,N_3020,N_572);
xnor U8490 (N_8490,N_5462,N_4700);
or U8491 (N_8491,N_2504,N_1687);
or U8492 (N_8492,N_3667,N_5423);
and U8493 (N_8493,N_1947,N_1441);
and U8494 (N_8494,N_2700,N_2479);
xnor U8495 (N_8495,N_47,N_2268);
nand U8496 (N_8496,N_5371,N_3800);
and U8497 (N_8497,N_3613,N_3050);
or U8498 (N_8498,N_5602,N_4600);
nor U8499 (N_8499,N_200,N_475);
or U8500 (N_8500,N_2048,N_1871);
xnor U8501 (N_8501,N_2087,N_568);
nand U8502 (N_8502,N_191,N_4646);
xnor U8503 (N_8503,N_3687,N_166);
or U8504 (N_8504,N_4944,N_1451);
nor U8505 (N_8505,N_1803,N_4718);
or U8506 (N_8506,N_2382,N_442);
nor U8507 (N_8507,N_2873,N_2190);
and U8508 (N_8508,N_842,N_5828);
nand U8509 (N_8509,N_1998,N_38);
nand U8510 (N_8510,N_4437,N_2969);
or U8511 (N_8511,N_4296,N_5071);
or U8512 (N_8512,N_674,N_564);
xor U8513 (N_8513,N_253,N_2709);
nand U8514 (N_8514,N_1582,N_4428);
and U8515 (N_8515,N_5850,N_4378);
xnor U8516 (N_8516,N_4286,N_2399);
or U8517 (N_8517,N_4779,N_524);
nor U8518 (N_8518,N_5860,N_3783);
xnor U8519 (N_8519,N_3561,N_811);
or U8520 (N_8520,N_5787,N_3754);
nand U8521 (N_8521,N_4208,N_3735);
and U8522 (N_8522,N_4463,N_755);
nor U8523 (N_8523,N_4450,N_1046);
nor U8524 (N_8524,N_4167,N_5756);
and U8525 (N_8525,N_2493,N_1833);
nor U8526 (N_8526,N_2749,N_2347);
nand U8527 (N_8527,N_408,N_5313);
and U8528 (N_8528,N_2303,N_472);
or U8529 (N_8529,N_284,N_3338);
nand U8530 (N_8530,N_3846,N_1864);
nand U8531 (N_8531,N_2275,N_323);
and U8532 (N_8532,N_1020,N_3044);
nor U8533 (N_8533,N_1084,N_2016);
nor U8534 (N_8534,N_254,N_1237);
xor U8535 (N_8535,N_5300,N_847);
nor U8536 (N_8536,N_1773,N_1151);
nand U8537 (N_8537,N_2144,N_169);
and U8538 (N_8538,N_3565,N_5331);
and U8539 (N_8539,N_5208,N_445);
nand U8540 (N_8540,N_3356,N_4941);
nor U8541 (N_8541,N_424,N_1882);
xnor U8542 (N_8542,N_5461,N_1707);
or U8543 (N_8543,N_2744,N_5908);
nor U8544 (N_8544,N_4374,N_5516);
and U8545 (N_8545,N_2620,N_4381);
and U8546 (N_8546,N_2816,N_5494);
nor U8547 (N_8547,N_1629,N_4133);
nor U8548 (N_8548,N_4860,N_3825);
nand U8549 (N_8549,N_5281,N_1275);
and U8550 (N_8550,N_1851,N_3158);
or U8551 (N_8551,N_2434,N_1665);
and U8552 (N_8552,N_4563,N_1795);
xnor U8553 (N_8553,N_2168,N_1484);
and U8554 (N_8554,N_5660,N_1205);
or U8555 (N_8555,N_5953,N_1857);
nor U8556 (N_8556,N_1329,N_5635);
nand U8557 (N_8557,N_941,N_2720);
or U8558 (N_8558,N_1141,N_857);
nand U8559 (N_8559,N_3216,N_1015);
and U8560 (N_8560,N_754,N_1028);
and U8561 (N_8561,N_2868,N_1610);
or U8562 (N_8562,N_2832,N_5214);
nor U8563 (N_8563,N_370,N_4311);
and U8564 (N_8564,N_983,N_5992);
xor U8565 (N_8565,N_5643,N_1525);
xnor U8566 (N_8566,N_4392,N_3794);
or U8567 (N_8567,N_3622,N_4403);
and U8568 (N_8568,N_1161,N_5532);
nand U8569 (N_8569,N_5827,N_2119);
nor U8570 (N_8570,N_3328,N_2143);
nor U8571 (N_8571,N_948,N_5952);
nand U8572 (N_8572,N_2311,N_4814);
nor U8573 (N_8573,N_393,N_4730);
and U8574 (N_8574,N_1163,N_2710);
or U8575 (N_8575,N_3048,N_4104);
or U8576 (N_8576,N_2512,N_5634);
or U8577 (N_8577,N_3184,N_1049);
and U8578 (N_8578,N_4268,N_4451);
xor U8579 (N_8579,N_2131,N_2289);
and U8580 (N_8580,N_5707,N_2707);
and U8581 (N_8581,N_252,N_3288);
or U8582 (N_8582,N_4545,N_4910);
or U8583 (N_8583,N_2998,N_873);
nor U8584 (N_8584,N_1180,N_5471);
nand U8585 (N_8585,N_3151,N_881);
xnor U8586 (N_8586,N_4983,N_5326);
xnor U8587 (N_8587,N_2206,N_1176);
or U8588 (N_8588,N_1088,N_5742);
nor U8589 (N_8589,N_5185,N_1206);
or U8590 (N_8590,N_5014,N_1867);
nor U8591 (N_8591,N_3178,N_5630);
and U8592 (N_8592,N_3933,N_2721);
nand U8593 (N_8593,N_382,N_3172);
or U8594 (N_8594,N_5854,N_3116);
and U8595 (N_8595,N_4182,N_2701);
and U8596 (N_8596,N_3627,N_5509);
nor U8597 (N_8597,N_5257,N_937);
xor U8598 (N_8598,N_2576,N_3569);
nor U8599 (N_8599,N_993,N_4109);
nand U8600 (N_8600,N_4693,N_1913);
or U8601 (N_8601,N_2089,N_3004);
nor U8602 (N_8602,N_5493,N_3503);
nand U8603 (N_8603,N_2501,N_4742);
nor U8604 (N_8604,N_5678,N_1662);
nand U8605 (N_8605,N_5395,N_1454);
nor U8606 (N_8606,N_5575,N_1222);
xor U8607 (N_8607,N_4314,N_5334);
and U8608 (N_8608,N_3773,N_1490);
or U8609 (N_8609,N_5456,N_908);
xnor U8610 (N_8610,N_3493,N_2780);
or U8611 (N_8611,N_5834,N_3086);
xor U8612 (N_8612,N_4537,N_650);
nand U8613 (N_8613,N_2550,N_1826);
or U8614 (N_8614,N_3812,N_208);
xnor U8615 (N_8615,N_3789,N_3107);
xor U8616 (N_8616,N_5975,N_4123);
or U8617 (N_8617,N_2767,N_280);
nand U8618 (N_8618,N_419,N_2948);
nand U8619 (N_8619,N_4117,N_2313);
or U8620 (N_8620,N_3434,N_4295);
or U8621 (N_8621,N_4,N_157);
xor U8622 (N_8622,N_1524,N_4424);
xnor U8623 (N_8623,N_2115,N_60);
nor U8624 (N_8624,N_4316,N_3750);
xnor U8625 (N_8625,N_1982,N_2745);
nor U8626 (N_8626,N_4030,N_3078);
nand U8627 (N_8627,N_684,N_3876);
nand U8628 (N_8628,N_2853,N_2588);
and U8629 (N_8629,N_3755,N_2388);
and U8630 (N_8630,N_2534,N_2041);
nand U8631 (N_8631,N_429,N_5640);
and U8632 (N_8632,N_4119,N_604);
and U8633 (N_8633,N_3154,N_3350);
xnor U8634 (N_8634,N_3132,N_2961);
or U8635 (N_8635,N_3507,N_83);
nor U8636 (N_8636,N_432,N_3523);
nand U8637 (N_8637,N_4620,N_3762);
and U8638 (N_8638,N_3886,N_1655);
or U8639 (N_8639,N_2604,N_423);
and U8640 (N_8640,N_2490,N_96);
or U8641 (N_8641,N_3059,N_5561);
and U8642 (N_8642,N_3984,N_2270);
xor U8643 (N_8643,N_844,N_2142);
nor U8644 (N_8644,N_379,N_2729);
xor U8645 (N_8645,N_2246,N_5981);
nor U8646 (N_8646,N_5024,N_1489);
nand U8647 (N_8647,N_3285,N_4596);
xor U8648 (N_8648,N_3703,N_1253);
xor U8649 (N_8649,N_5297,N_3897);
and U8650 (N_8650,N_19,N_966);
nand U8651 (N_8651,N_760,N_215);
nor U8652 (N_8652,N_1043,N_2126);
xor U8653 (N_8653,N_3417,N_4349);
nor U8654 (N_8654,N_437,N_3628);
nor U8655 (N_8655,N_3022,N_5314);
and U8656 (N_8656,N_2978,N_2314);
xnor U8657 (N_8657,N_277,N_2840);
and U8658 (N_8658,N_1148,N_2081);
and U8659 (N_8659,N_434,N_5673);
xnor U8660 (N_8660,N_3174,N_522);
nor U8661 (N_8661,N_2950,N_801);
and U8662 (N_8662,N_1321,N_1729);
nor U8663 (N_8663,N_4592,N_2033);
nand U8664 (N_8664,N_4721,N_2335);
and U8665 (N_8665,N_4857,N_848);
nor U8666 (N_8666,N_2596,N_3839);
xnor U8667 (N_8667,N_1073,N_1332);
xor U8668 (N_8668,N_3443,N_5473);
xor U8669 (N_8669,N_5708,N_258);
xor U8670 (N_8670,N_203,N_1034);
and U8671 (N_8671,N_856,N_4058);
or U8672 (N_8672,N_5806,N_4483);
xor U8673 (N_8673,N_3144,N_384);
and U8674 (N_8674,N_4142,N_5063);
nor U8675 (N_8675,N_4977,N_4925);
or U8676 (N_8676,N_267,N_2912);
nand U8677 (N_8677,N_3980,N_4152);
xnor U8678 (N_8678,N_554,N_1330);
and U8679 (N_8679,N_5367,N_1442);
and U8680 (N_8680,N_2753,N_2405);
xnor U8681 (N_8681,N_3544,N_4255);
nor U8682 (N_8682,N_2694,N_787);
or U8683 (N_8683,N_556,N_1281);
nor U8684 (N_8684,N_3309,N_78);
nor U8685 (N_8685,N_1887,N_2279);
xor U8686 (N_8686,N_5501,N_4939);
nand U8687 (N_8687,N_4039,N_15);
xnor U8688 (N_8688,N_3838,N_4517);
nand U8689 (N_8689,N_3346,N_4641);
nand U8690 (N_8690,N_289,N_4065);
nor U8691 (N_8691,N_1220,N_5857);
nand U8692 (N_8692,N_1469,N_204);
nand U8693 (N_8693,N_3576,N_5448);
xor U8694 (N_8694,N_5843,N_4114);
nand U8695 (N_8695,N_1888,N_5283);
and U8696 (N_8696,N_4502,N_315);
nor U8697 (N_8697,N_1642,N_3207);
or U8698 (N_8698,N_4465,N_1577);
nor U8699 (N_8699,N_4359,N_5949);
xor U8700 (N_8700,N_3031,N_304);
xnor U8701 (N_8701,N_4710,N_2215);
xnor U8702 (N_8702,N_5364,N_2031);
xor U8703 (N_8703,N_619,N_4953);
or U8704 (N_8704,N_3028,N_3183);
nor U8705 (N_8705,N_3114,N_5068);
and U8706 (N_8706,N_777,N_1396);
or U8707 (N_8707,N_961,N_4063);
nor U8708 (N_8708,N_2857,N_1135);
nor U8709 (N_8709,N_4467,N_3896);
xor U8710 (N_8710,N_3715,N_4699);
and U8711 (N_8711,N_205,N_4530);
and U8712 (N_8712,N_4703,N_5359);
nand U8713 (N_8713,N_3928,N_3698);
and U8714 (N_8714,N_5779,N_1353);
or U8715 (N_8715,N_3587,N_1968);
nand U8716 (N_8716,N_2988,N_43);
xnor U8717 (N_8717,N_3499,N_1429);
and U8718 (N_8718,N_1093,N_2039);
xor U8719 (N_8719,N_5599,N_292);
nand U8720 (N_8720,N_3110,N_5735);
and U8721 (N_8721,N_3009,N_1909);
and U8722 (N_8722,N_2803,N_5947);
xor U8723 (N_8723,N_3644,N_459);
nor U8724 (N_8724,N_2161,N_479);
xor U8725 (N_8725,N_3618,N_920);
and U8726 (N_8726,N_785,N_1431);
nand U8727 (N_8727,N_1667,N_1984);
xor U8728 (N_8728,N_3625,N_4116);
nor U8729 (N_8729,N_3252,N_3679);
and U8730 (N_8730,N_328,N_5144);
xnor U8731 (N_8731,N_1520,N_5073);
xnor U8732 (N_8732,N_5454,N_4869);
nor U8733 (N_8733,N_515,N_1996);
nor U8734 (N_8734,N_5261,N_796);
or U8735 (N_8735,N_2288,N_2277);
nor U8736 (N_8736,N_5549,N_1269);
nand U8737 (N_8737,N_4477,N_62);
nand U8738 (N_8738,N_706,N_5695);
or U8739 (N_8739,N_2845,N_121);
nand U8740 (N_8740,N_5829,N_776);
and U8741 (N_8741,N_1232,N_5295);
nand U8742 (N_8742,N_4898,N_5904);
nand U8743 (N_8743,N_4138,N_5339);
xnor U8744 (N_8744,N_3986,N_3657);
and U8745 (N_8745,N_4482,N_4489);
nor U8746 (N_8746,N_4602,N_1499);
and U8747 (N_8747,N_837,N_1131);
nor U8748 (N_8748,N_1552,N_4774);
xnor U8749 (N_8749,N_5670,N_5056);
xnor U8750 (N_8750,N_5130,N_178);
xor U8751 (N_8751,N_1250,N_2553);
nand U8752 (N_8752,N_4368,N_144);
or U8753 (N_8753,N_1142,N_4709);
xor U8754 (N_8754,N_1217,N_344);
or U8755 (N_8755,N_5023,N_907);
nor U8756 (N_8756,N_1387,N_793);
and U8757 (N_8757,N_5427,N_3227);
xor U8758 (N_8758,N_1168,N_1837);
xor U8759 (N_8759,N_806,N_4501);
and U8760 (N_8760,N_400,N_2265);
nor U8761 (N_8761,N_3957,N_3147);
and U8762 (N_8762,N_3495,N_2484);
or U8763 (N_8763,N_4897,N_3128);
or U8764 (N_8764,N_506,N_3633);
xor U8765 (N_8765,N_2476,N_5913);
nor U8766 (N_8766,N_1386,N_1798);
nand U8767 (N_8767,N_2574,N_4047);
xnor U8768 (N_8768,N_1313,N_1284);
or U8769 (N_8769,N_1832,N_2673);
xor U8770 (N_8770,N_976,N_4844);
nor U8771 (N_8771,N_5862,N_1677);
or U8772 (N_8772,N_1792,N_2220);
xor U8773 (N_8773,N_1835,N_5736);
nand U8774 (N_8774,N_5285,N_4772);
or U8775 (N_8775,N_1957,N_2093);
nand U8776 (N_8776,N_2006,N_4308);
xnor U8777 (N_8777,N_4373,N_4391);
or U8778 (N_8778,N_231,N_4675);
nand U8779 (N_8779,N_270,N_775);
and U8780 (N_8780,N_4017,N_72);
nand U8781 (N_8781,N_2650,N_5017);
or U8782 (N_8782,N_2301,N_80);
or U8783 (N_8783,N_5556,N_2531);
or U8784 (N_8784,N_5519,N_4436);
xnor U8785 (N_8785,N_5061,N_4711);
and U8786 (N_8786,N_926,N_2349);
or U8787 (N_8787,N_644,N_784);
and U8788 (N_8788,N_2290,N_2640);
and U8789 (N_8789,N_2024,N_685);
and U8790 (N_8790,N_5181,N_814);
nor U8791 (N_8791,N_740,N_5034);
xor U8792 (N_8792,N_2370,N_2842);
nand U8793 (N_8793,N_3962,N_5489);
nor U8794 (N_8794,N_4956,N_3879);
nor U8795 (N_8795,N_3943,N_3377);
xnor U8796 (N_8796,N_739,N_3770);
or U8797 (N_8797,N_3801,N_3537);
nor U8798 (N_8798,N_130,N_5201);
nand U8799 (N_8799,N_4609,N_519);
xnor U8800 (N_8800,N_729,N_69);
nand U8801 (N_8801,N_2278,N_1320);
nor U8802 (N_8802,N_5710,N_2556);
nor U8803 (N_8803,N_4916,N_3475);
or U8804 (N_8804,N_2054,N_4305);
and U8805 (N_8805,N_5925,N_3413);
nand U8806 (N_8806,N_3588,N_2601);
nand U8807 (N_8807,N_4107,N_1546);
nand U8808 (N_8808,N_3653,N_5721);
or U8809 (N_8809,N_3431,N_2825);
or U8810 (N_8810,N_2014,N_1621);
or U8811 (N_8811,N_1698,N_5790);
or U8812 (N_8812,N_2026,N_3757);
xor U8813 (N_8813,N_1449,N_4279);
xnor U8814 (N_8814,N_5548,N_3081);
and U8815 (N_8815,N_5229,N_871);
nor U8816 (N_8816,N_639,N_5972);
xnor U8817 (N_8817,N_1375,N_5200);
xnor U8818 (N_8818,N_1296,N_4713);
nor U8819 (N_8819,N_5470,N_182);
or U8820 (N_8820,N_1126,N_99);
xor U8821 (N_8821,N_3054,N_3889);
or U8822 (N_8822,N_3182,N_3934);
or U8823 (N_8823,N_5166,N_5591);
nor U8824 (N_8824,N_4508,N_452);
and U8825 (N_8825,N_1797,N_5679);
nand U8826 (N_8826,N_2922,N_1017);
and U8827 (N_8827,N_640,N_4002);
xnor U8828 (N_8828,N_450,N_433);
xnor U8829 (N_8829,N_4746,N_2468);
nand U8830 (N_8830,N_636,N_4667);
or U8831 (N_8831,N_2641,N_1836);
nand U8832 (N_8832,N_766,N_1917);
or U8833 (N_8833,N_5476,N_5296);
and U8834 (N_8834,N_1528,N_4052);
nor U8835 (N_8835,N_3527,N_990);
or U8836 (N_8836,N_1762,N_326);
xnor U8837 (N_8837,N_8,N_5563);
nand U8838 (N_8838,N_5615,N_449);
nor U8839 (N_8839,N_2195,N_4988);
nor U8840 (N_8840,N_1210,N_3585);
and U8841 (N_8841,N_2486,N_3798);
or U8842 (N_8842,N_5353,N_5520);
and U8843 (N_8843,N_1293,N_3371);
or U8844 (N_8844,N_4800,N_5507);
xor U8845 (N_8845,N_4617,N_3765);
nand U8846 (N_8846,N_5212,N_4690);
nor U8847 (N_8847,N_4929,N_1932);
and U8848 (N_8848,N_5076,N_3926);
or U8849 (N_8849,N_4141,N_4076);
and U8850 (N_8850,N_1247,N_4683);
nand U8851 (N_8851,N_5119,N_4677);
nand U8852 (N_8852,N_4579,N_5650);
nand U8853 (N_8853,N_3831,N_1243);
xnor U8854 (N_8854,N_1235,N_518);
nand U8855 (N_8855,N_91,N_5057);
nand U8856 (N_8856,N_728,N_3485);
nor U8857 (N_8857,N_4873,N_5960);
and U8858 (N_8858,N_4031,N_5553);
or U8859 (N_8859,N_5921,N_3348);
or U8860 (N_8860,N_5149,N_4831);
xor U8861 (N_8861,N_3849,N_61);
nand U8862 (N_8862,N_180,N_1008);
nand U8863 (N_8863,N_2260,N_5522);
and U8864 (N_8864,N_2771,N_5999);
or U8865 (N_8865,N_3125,N_5697);
nor U8866 (N_8866,N_3631,N_2122);
and U8867 (N_8867,N_4867,N_1672);
nand U8868 (N_8868,N_744,N_1230);
and U8869 (N_8869,N_520,N_3488);
and U8870 (N_8870,N_361,N_810);
and U8871 (N_8871,N_5848,N_5956);
or U8872 (N_8872,N_3058,N_3218);
and U8873 (N_8873,N_981,N_4307);
nor U8874 (N_8874,N_4595,N_1796);
xor U8875 (N_8875,N_1868,N_2401);
nand U8876 (N_8876,N_2355,N_1400);
nand U8877 (N_8877,N_3072,N_4125);
nand U8878 (N_8878,N_4023,N_552);
nand U8879 (N_8879,N_1540,N_1550);
nand U8880 (N_8880,N_3222,N_4947);
nand U8881 (N_8881,N_5008,N_2419);
nor U8882 (N_8882,N_576,N_4466);
xor U8883 (N_8883,N_1344,N_5093);
and U8884 (N_8884,N_1146,N_5616);
nor U8885 (N_8885,N_5211,N_1308);
nand U8886 (N_8886,N_1147,N_5432);
nor U8887 (N_8887,N_2325,N_4278);
nor U8888 (N_8888,N_3006,N_4893);
nand U8889 (N_8889,N_385,N_4462);
nor U8890 (N_8890,N_2660,N_3017);
xnor U8891 (N_8891,N_1934,N_2715);
nand U8892 (N_8892,N_3976,N_2398);
or U8893 (N_8893,N_2107,N_2894);
xor U8894 (N_8894,N_2696,N_1816);
nand U8895 (N_8895,N_5305,N_835);
nand U8896 (N_8896,N_5288,N_5565);
xor U8897 (N_8897,N_5898,N_3224);
nor U8898 (N_8898,N_3970,N_5258);
xor U8899 (N_8899,N_1521,N_822);
or U8900 (N_8900,N_4073,N_843);
and U8901 (N_8901,N_4232,N_401);
xnor U8902 (N_8902,N_2299,N_1758);
nand U8903 (N_8903,N_736,N_5663);
and U8904 (N_8904,N_813,N_2913);
xor U8905 (N_8905,N_4081,N_1263);
nor U8906 (N_8906,N_1670,N_3477);
and U8907 (N_8907,N_1945,N_52);
xnor U8908 (N_8908,N_4993,N_2973);
and U8909 (N_8909,N_4830,N_504);
nor U8910 (N_8910,N_770,N_5136);
or U8911 (N_8911,N_3264,N_4938);
nand U8912 (N_8912,N_894,N_5943);
and U8913 (N_8913,N_2651,N_5443);
and U8914 (N_8914,N_2205,N_5110);
xor U8915 (N_8915,N_2635,N_2481);
and U8916 (N_8916,N_5237,N_1953);
xnor U8917 (N_8917,N_2751,N_4341);
xnor U8918 (N_8918,N_2654,N_1358);
nand U8919 (N_8919,N_1669,N_5239);
xnor U8920 (N_8920,N_863,N_1323);
nand U8921 (N_8921,N_1195,N_5098);
and U8922 (N_8922,N_1512,N_5250);
nand U8923 (N_8923,N_394,N_5355);
nand U8924 (N_8924,N_362,N_3604);
nand U8925 (N_8925,N_3186,N_1465);
or U8926 (N_8926,N_4702,N_299);
or U8927 (N_8927,N_1379,N_1752);
or U8928 (N_8928,N_889,N_2480);
nand U8929 (N_8929,N_1042,N_523);
nand U8930 (N_8930,N_5316,N_2116);
nand U8931 (N_8931,N_5823,N_1385);
nand U8932 (N_8932,N_1346,N_286);
nand U8933 (N_8933,N_4342,N_927);
nand U8934 (N_8934,N_2524,N_3230);
nand U8935 (N_8935,N_4100,N_1548);
nor U8936 (N_8936,N_4707,N_2760);
and U8937 (N_8937,N_936,N_2824);
or U8938 (N_8938,N_659,N_4097);
nor U8939 (N_8939,N_291,N_5976);
or U8940 (N_8940,N_968,N_1886);
and U8941 (N_8941,N_4768,N_4732);
and U8942 (N_8942,N_5665,N_5838);
and U8943 (N_8943,N_3894,N_543);
nand U8944 (N_8944,N_2692,N_1365);
and U8945 (N_8945,N_914,N_4210);
nand U8946 (N_8946,N_4601,N_3917);
and U8947 (N_8947,N_666,N_1935);
or U8948 (N_8948,N_2237,N_4136);
xnor U8949 (N_8949,N_629,N_5227);
nand U8950 (N_8950,N_4439,N_2563);
nor U8951 (N_8951,N_3684,N_3057);
nor U8952 (N_8952,N_194,N_1376);
xor U8953 (N_8953,N_1633,N_751);
and U8954 (N_8954,N_5088,N_608);
nand U8955 (N_8955,N_4848,N_4986);
xnor U8956 (N_8956,N_4459,N_159);
nand U8957 (N_8957,N_3108,N_4129);
nand U8958 (N_8958,N_3188,N_3632);
xor U8959 (N_8959,N_1095,N_4380);
or U8960 (N_8960,N_1791,N_2831);
and U8961 (N_8961,N_526,N_1381);
and U8962 (N_8962,N_123,N_4485);
nand U8963 (N_8963,N_4877,N_5060);
or U8964 (N_8964,N_4197,N_5536);
or U8965 (N_8965,N_5784,N_4874);
nor U8966 (N_8966,N_4226,N_3007);
and U8967 (N_8967,N_2577,N_3516);
nand U8968 (N_8968,N_1479,N_3232);
xnor U8969 (N_8969,N_4025,N_2653);
xor U8970 (N_8970,N_995,N_5963);
nand U8971 (N_8971,N_3596,N_5937);
and U8972 (N_8972,N_3936,N_4780);
nand U8973 (N_8973,N_1432,N_5884);
xor U8974 (N_8974,N_1688,N_427);
or U8975 (N_8975,N_5238,N_3388);
xnor U8976 (N_8976,N_5965,N_4347);
xor U8977 (N_8977,N_4158,N_1660);
or U8978 (N_8978,N_5193,N_4534);
xnor U8979 (N_8979,N_5165,N_1070);
and U8980 (N_8980,N_5778,N_5446);
xnor U8981 (N_8981,N_1482,N_4843);
xor U8982 (N_8982,N_2537,N_5929);
or U8983 (N_8983,N_1354,N_4149);
nand U8984 (N_8984,N_3029,N_2936);
nand U8985 (N_8985,N_173,N_145);
xor U8986 (N_8986,N_1200,N_3739);
or U8987 (N_8987,N_1812,N_5321);
or U8988 (N_8988,N_2439,N_3560);
or U8989 (N_8989,N_925,N_4171);
or U8990 (N_8990,N_4336,N_4032);
nor U8991 (N_8991,N_5906,N_5419);
nand U8992 (N_8992,N_4093,N_872);
and U8993 (N_8993,N_4371,N_5719);
or U8994 (N_8994,N_486,N_4390);
or U8995 (N_8995,N_4604,N_5597);
nor U8996 (N_8996,N_3246,N_2058);
nor U8997 (N_8997,N_5560,N_1778);
xnor U8998 (N_8998,N_1716,N_211);
and U8999 (N_8999,N_5040,N_1802);
xnor U9000 (N_9000,N_2534,N_4855);
xnor U9001 (N_9001,N_4399,N_4273);
or U9002 (N_9002,N_1972,N_2631);
nor U9003 (N_9003,N_7,N_5794);
nand U9004 (N_9004,N_864,N_2135);
nor U9005 (N_9005,N_3222,N_2645);
nand U9006 (N_9006,N_653,N_5633);
and U9007 (N_9007,N_1962,N_5149);
nand U9008 (N_9008,N_1979,N_1335);
xnor U9009 (N_9009,N_2865,N_4643);
xnor U9010 (N_9010,N_5695,N_1490);
xnor U9011 (N_9011,N_3936,N_1996);
and U9012 (N_9012,N_3542,N_5979);
nor U9013 (N_9013,N_4964,N_5472);
or U9014 (N_9014,N_5238,N_3081);
or U9015 (N_9015,N_4472,N_1243);
or U9016 (N_9016,N_1103,N_3700);
and U9017 (N_9017,N_2424,N_5562);
nand U9018 (N_9018,N_2335,N_4424);
and U9019 (N_9019,N_4359,N_1328);
or U9020 (N_9020,N_5842,N_2184);
and U9021 (N_9021,N_3484,N_781);
nand U9022 (N_9022,N_2667,N_1234);
nor U9023 (N_9023,N_1751,N_2899);
or U9024 (N_9024,N_5499,N_2516);
xor U9025 (N_9025,N_4375,N_4952);
nand U9026 (N_9026,N_1058,N_4017);
xnor U9027 (N_9027,N_1139,N_5118);
nor U9028 (N_9028,N_4115,N_4689);
nand U9029 (N_9029,N_2800,N_1574);
xnor U9030 (N_9030,N_5462,N_2094);
or U9031 (N_9031,N_5018,N_2505);
and U9032 (N_9032,N_5093,N_1022);
xor U9033 (N_9033,N_232,N_2249);
or U9034 (N_9034,N_5450,N_4239);
nand U9035 (N_9035,N_3845,N_5299);
nor U9036 (N_9036,N_1134,N_4815);
or U9037 (N_9037,N_3184,N_3441);
nor U9038 (N_9038,N_4492,N_1892);
or U9039 (N_9039,N_3320,N_2710);
or U9040 (N_9040,N_3146,N_2665);
or U9041 (N_9041,N_505,N_5086);
and U9042 (N_9042,N_1369,N_886);
and U9043 (N_9043,N_2286,N_5342);
or U9044 (N_9044,N_5921,N_86);
nor U9045 (N_9045,N_1054,N_4628);
and U9046 (N_9046,N_5635,N_771);
nand U9047 (N_9047,N_2837,N_725);
nand U9048 (N_9048,N_787,N_2721);
nor U9049 (N_9049,N_1811,N_16);
xor U9050 (N_9050,N_5810,N_2583);
xnor U9051 (N_9051,N_3087,N_4002);
or U9052 (N_9052,N_4111,N_4009);
nand U9053 (N_9053,N_1477,N_4932);
or U9054 (N_9054,N_3036,N_2363);
and U9055 (N_9055,N_4873,N_5140);
nor U9056 (N_9056,N_5212,N_4502);
nor U9057 (N_9057,N_1243,N_5625);
or U9058 (N_9058,N_5617,N_3840);
or U9059 (N_9059,N_1005,N_345);
and U9060 (N_9060,N_2975,N_5165);
nand U9061 (N_9061,N_3374,N_3543);
nand U9062 (N_9062,N_5740,N_4815);
xor U9063 (N_9063,N_89,N_3507);
nand U9064 (N_9064,N_3435,N_5764);
xnor U9065 (N_9065,N_2590,N_667);
nor U9066 (N_9066,N_1147,N_3229);
nand U9067 (N_9067,N_4150,N_3112);
nand U9068 (N_9068,N_5154,N_4591);
or U9069 (N_9069,N_4605,N_685);
xnor U9070 (N_9070,N_3871,N_2515);
or U9071 (N_9071,N_4714,N_1093);
or U9072 (N_9072,N_4895,N_4856);
and U9073 (N_9073,N_4170,N_226);
and U9074 (N_9074,N_5498,N_4112);
xnor U9075 (N_9075,N_5828,N_5601);
nor U9076 (N_9076,N_1740,N_379);
and U9077 (N_9077,N_3533,N_1655);
and U9078 (N_9078,N_5992,N_1172);
or U9079 (N_9079,N_840,N_5834);
xor U9080 (N_9080,N_127,N_2691);
and U9081 (N_9081,N_2552,N_845);
and U9082 (N_9082,N_1309,N_926);
xnor U9083 (N_9083,N_3131,N_125);
and U9084 (N_9084,N_3573,N_4755);
nand U9085 (N_9085,N_3136,N_5144);
xor U9086 (N_9086,N_4083,N_2845);
or U9087 (N_9087,N_4044,N_174);
and U9088 (N_9088,N_608,N_4697);
and U9089 (N_9089,N_3806,N_4345);
xor U9090 (N_9090,N_5336,N_2329);
or U9091 (N_9091,N_4359,N_2120);
or U9092 (N_9092,N_4575,N_2821);
nor U9093 (N_9093,N_2592,N_5180);
and U9094 (N_9094,N_1042,N_5550);
xor U9095 (N_9095,N_2160,N_1780);
and U9096 (N_9096,N_86,N_1722);
nand U9097 (N_9097,N_5521,N_2433);
and U9098 (N_9098,N_158,N_1598);
xor U9099 (N_9099,N_325,N_3514);
and U9100 (N_9100,N_696,N_2080);
and U9101 (N_9101,N_4305,N_3636);
nor U9102 (N_9102,N_3598,N_3141);
nand U9103 (N_9103,N_1480,N_1567);
nor U9104 (N_9104,N_4707,N_5366);
nand U9105 (N_9105,N_700,N_5822);
nor U9106 (N_9106,N_2701,N_1517);
nor U9107 (N_9107,N_2199,N_4443);
nor U9108 (N_9108,N_4292,N_5533);
nor U9109 (N_9109,N_166,N_5102);
or U9110 (N_9110,N_790,N_1409);
nor U9111 (N_9111,N_422,N_5609);
or U9112 (N_9112,N_4915,N_5353);
or U9113 (N_9113,N_820,N_3485);
xnor U9114 (N_9114,N_382,N_2339);
and U9115 (N_9115,N_634,N_2868);
xor U9116 (N_9116,N_4164,N_3154);
or U9117 (N_9117,N_2838,N_790);
nor U9118 (N_9118,N_5846,N_1262);
xnor U9119 (N_9119,N_3862,N_5323);
nand U9120 (N_9120,N_3790,N_3278);
nand U9121 (N_9121,N_2768,N_783);
or U9122 (N_9122,N_5738,N_1022);
and U9123 (N_9123,N_4207,N_3405);
nand U9124 (N_9124,N_604,N_4775);
or U9125 (N_9125,N_5801,N_1712);
or U9126 (N_9126,N_2597,N_3750);
nor U9127 (N_9127,N_348,N_5120);
nor U9128 (N_9128,N_4645,N_3256);
xnor U9129 (N_9129,N_2942,N_4914);
nor U9130 (N_9130,N_2844,N_5735);
and U9131 (N_9131,N_5606,N_5162);
and U9132 (N_9132,N_2914,N_4742);
xnor U9133 (N_9133,N_5717,N_3142);
and U9134 (N_9134,N_4667,N_3794);
or U9135 (N_9135,N_4540,N_2722);
xor U9136 (N_9136,N_4219,N_5761);
or U9137 (N_9137,N_2674,N_5909);
xor U9138 (N_9138,N_1353,N_5831);
and U9139 (N_9139,N_3921,N_1312);
or U9140 (N_9140,N_2164,N_623);
and U9141 (N_9141,N_3792,N_2384);
xnor U9142 (N_9142,N_3848,N_4995);
nand U9143 (N_9143,N_2057,N_2849);
or U9144 (N_9144,N_3552,N_845);
or U9145 (N_9145,N_4187,N_5758);
nand U9146 (N_9146,N_2975,N_4921);
nor U9147 (N_9147,N_1523,N_512);
nor U9148 (N_9148,N_2743,N_1523);
and U9149 (N_9149,N_2721,N_5986);
or U9150 (N_9150,N_2659,N_3975);
or U9151 (N_9151,N_3405,N_1260);
xor U9152 (N_9152,N_5567,N_4210);
or U9153 (N_9153,N_3312,N_4693);
xor U9154 (N_9154,N_1837,N_5387);
or U9155 (N_9155,N_5216,N_5470);
nand U9156 (N_9156,N_4904,N_1022);
or U9157 (N_9157,N_3693,N_527);
xnor U9158 (N_9158,N_1849,N_587);
nand U9159 (N_9159,N_1026,N_598);
nand U9160 (N_9160,N_1440,N_756);
xnor U9161 (N_9161,N_4803,N_3582);
or U9162 (N_9162,N_3619,N_5882);
or U9163 (N_9163,N_2895,N_1841);
or U9164 (N_9164,N_5865,N_480);
xor U9165 (N_9165,N_1000,N_4145);
nand U9166 (N_9166,N_1604,N_2947);
nand U9167 (N_9167,N_447,N_4368);
nor U9168 (N_9168,N_1605,N_1133);
xor U9169 (N_9169,N_4408,N_4447);
or U9170 (N_9170,N_1374,N_3463);
and U9171 (N_9171,N_880,N_4462);
xnor U9172 (N_9172,N_535,N_1757);
xnor U9173 (N_9173,N_1131,N_111);
and U9174 (N_9174,N_3977,N_578);
nor U9175 (N_9175,N_5811,N_3999);
and U9176 (N_9176,N_2836,N_3912);
nand U9177 (N_9177,N_4280,N_1557);
nand U9178 (N_9178,N_204,N_2890);
nand U9179 (N_9179,N_5817,N_3175);
and U9180 (N_9180,N_3903,N_2811);
or U9181 (N_9181,N_2341,N_1171);
nor U9182 (N_9182,N_4556,N_2039);
or U9183 (N_9183,N_3949,N_1249);
xor U9184 (N_9184,N_5148,N_530);
or U9185 (N_9185,N_3298,N_5497);
nor U9186 (N_9186,N_3071,N_1652);
nor U9187 (N_9187,N_637,N_1994);
or U9188 (N_9188,N_4296,N_2258);
xor U9189 (N_9189,N_3033,N_492);
nand U9190 (N_9190,N_847,N_2783);
nand U9191 (N_9191,N_578,N_932);
nand U9192 (N_9192,N_5061,N_488);
xor U9193 (N_9193,N_914,N_1754);
xnor U9194 (N_9194,N_1486,N_5406);
and U9195 (N_9195,N_4221,N_503);
or U9196 (N_9196,N_3007,N_16);
and U9197 (N_9197,N_1339,N_3818);
nand U9198 (N_9198,N_1455,N_3572);
nand U9199 (N_9199,N_3681,N_2539);
nor U9200 (N_9200,N_342,N_5947);
nor U9201 (N_9201,N_1474,N_3623);
or U9202 (N_9202,N_811,N_1742);
and U9203 (N_9203,N_2843,N_3984);
nor U9204 (N_9204,N_72,N_3821);
nor U9205 (N_9205,N_5870,N_2886);
nand U9206 (N_9206,N_3828,N_3460);
and U9207 (N_9207,N_3335,N_1471);
or U9208 (N_9208,N_5983,N_5574);
and U9209 (N_9209,N_1821,N_263);
nand U9210 (N_9210,N_5461,N_2669);
nor U9211 (N_9211,N_4346,N_2959);
nand U9212 (N_9212,N_3955,N_3984);
nand U9213 (N_9213,N_1994,N_2643);
and U9214 (N_9214,N_4768,N_3105);
nand U9215 (N_9215,N_4841,N_5618);
or U9216 (N_9216,N_1155,N_596);
xnor U9217 (N_9217,N_2236,N_3416);
nor U9218 (N_9218,N_3697,N_3983);
nand U9219 (N_9219,N_5271,N_935);
nor U9220 (N_9220,N_5814,N_2647);
nand U9221 (N_9221,N_892,N_4207);
and U9222 (N_9222,N_5832,N_875);
nor U9223 (N_9223,N_1105,N_4042);
or U9224 (N_9224,N_5533,N_1914);
nand U9225 (N_9225,N_1264,N_3572);
or U9226 (N_9226,N_4432,N_1287);
nor U9227 (N_9227,N_2574,N_2384);
xnor U9228 (N_9228,N_4885,N_4473);
nor U9229 (N_9229,N_2519,N_3738);
and U9230 (N_9230,N_544,N_5342);
or U9231 (N_9231,N_1014,N_2189);
xor U9232 (N_9232,N_4664,N_2668);
and U9233 (N_9233,N_5377,N_1128);
xor U9234 (N_9234,N_5810,N_2158);
or U9235 (N_9235,N_5593,N_5335);
or U9236 (N_9236,N_4108,N_3547);
xnor U9237 (N_9237,N_4818,N_5246);
or U9238 (N_9238,N_1992,N_822);
nand U9239 (N_9239,N_1137,N_314);
or U9240 (N_9240,N_2763,N_614);
nor U9241 (N_9241,N_4469,N_2586);
or U9242 (N_9242,N_567,N_4256);
nand U9243 (N_9243,N_2699,N_2303);
nor U9244 (N_9244,N_3515,N_1534);
xor U9245 (N_9245,N_1284,N_2548);
or U9246 (N_9246,N_3149,N_2220);
xor U9247 (N_9247,N_3658,N_2953);
or U9248 (N_9248,N_3528,N_1997);
and U9249 (N_9249,N_5769,N_3124);
and U9250 (N_9250,N_5634,N_5319);
nand U9251 (N_9251,N_5848,N_33);
and U9252 (N_9252,N_426,N_4088);
or U9253 (N_9253,N_3099,N_195);
and U9254 (N_9254,N_1629,N_2686);
and U9255 (N_9255,N_3404,N_3215);
or U9256 (N_9256,N_4347,N_5647);
nand U9257 (N_9257,N_4108,N_1844);
xnor U9258 (N_9258,N_4345,N_5895);
nand U9259 (N_9259,N_4054,N_510);
or U9260 (N_9260,N_4617,N_2783);
or U9261 (N_9261,N_4374,N_1482);
nand U9262 (N_9262,N_267,N_5467);
xor U9263 (N_9263,N_289,N_339);
and U9264 (N_9264,N_1627,N_1749);
and U9265 (N_9265,N_2570,N_674);
nor U9266 (N_9266,N_4500,N_5106);
and U9267 (N_9267,N_5319,N_3113);
xnor U9268 (N_9268,N_247,N_2141);
nand U9269 (N_9269,N_3789,N_4304);
and U9270 (N_9270,N_2787,N_1588);
nor U9271 (N_9271,N_982,N_3209);
nor U9272 (N_9272,N_1753,N_49);
and U9273 (N_9273,N_3761,N_3061);
or U9274 (N_9274,N_113,N_4306);
and U9275 (N_9275,N_2103,N_4686);
nand U9276 (N_9276,N_2588,N_1900);
nor U9277 (N_9277,N_5418,N_1304);
or U9278 (N_9278,N_4217,N_5251);
nand U9279 (N_9279,N_4908,N_4326);
xor U9280 (N_9280,N_1412,N_4546);
or U9281 (N_9281,N_4339,N_3506);
nand U9282 (N_9282,N_2988,N_3521);
nand U9283 (N_9283,N_3763,N_415);
and U9284 (N_9284,N_4301,N_4917);
and U9285 (N_9285,N_5252,N_588);
and U9286 (N_9286,N_4376,N_3802);
nand U9287 (N_9287,N_1929,N_455);
nor U9288 (N_9288,N_5193,N_1425);
nand U9289 (N_9289,N_3528,N_605);
or U9290 (N_9290,N_2045,N_1079);
nand U9291 (N_9291,N_2540,N_4637);
and U9292 (N_9292,N_5994,N_4999);
and U9293 (N_9293,N_429,N_707);
xnor U9294 (N_9294,N_4755,N_856);
or U9295 (N_9295,N_4072,N_816);
and U9296 (N_9296,N_1620,N_5321);
xor U9297 (N_9297,N_5733,N_1260);
or U9298 (N_9298,N_1067,N_4099);
or U9299 (N_9299,N_3932,N_4828);
nor U9300 (N_9300,N_938,N_3887);
xor U9301 (N_9301,N_4006,N_181);
and U9302 (N_9302,N_141,N_1302);
xor U9303 (N_9303,N_5702,N_1155);
or U9304 (N_9304,N_2065,N_2872);
or U9305 (N_9305,N_2126,N_1223);
nand U9306 (N_9306,N_2699,N_547);
or U9307 (N_9307,N_2967,N_4070);
or U9308 (N_9308,N_4187,N_2914);
xnor U9309 (N_9309,N_2962,N_3489);
nor U9310 (N_9310,N_3883,N_4715);
nand U9311 (N_9311,N_808,N_719);
nand U9312 (N_9312,N_2404,N_4809);
or U9313 (N_9313,N_5680,N_4579);
and U9314 (N_9314,N_1912,N_72);
xor U9315 (N_9315,N_2479,N_2116);
nor U9316 (N_9316,N_4556,N_1832);
nor U9317 (N_9317,N_4113,N_2411);
xnor U9318 (N_9318,N_5097,N_1908);
nor U9319 (N_9319,N_2283,N_2130);
nand U9320 (N_9320,N_5084,N_1309);
nor U9321 (N_9321,N_2441,N_3016);
nand U9322 (N_9322,N_16,N_124);
nand U9323 (N_9323,N_3031,N_3350);
xnor U9324 (N_9324,N_2052,N_3417);
nand U9325 (N_9325,N_5004,N_5994);
nor U9326 (N_9326,N_2644,N_2572);
nand U9327 (N_9327,N_5682,N_5747);
nor U9328 (N_9328,N_4857,N_5787);
nor U9329 (N_9329,N_5831,N_190);
nand U9330 (N_9330,N_2248,N_2832);
xor U9331 (N_9331,N_28,N_2573);
or U9332 (N_9332,N_3216,N_1240);
nand U9333 (N_9333,N_494,N_184);
or U9334 (N_9334,N_4410,N_2434);
or U9335 (N_9335,N_718,N_268);
nor U9336 (N_9336,N_5675,N_4774);
and U9337 (N_9337,N_2515,N_1226);
and U9338 (N_9338,N_2846,N_3554);
nand U9339 (N_9339,N_5021,N_5718);
or U9340 (N_9340,N_4821,N_54);
nand U9341 (N_9341,N_2570,N_2378);
nand U9342 (N_9342,N_342,N_1577);
nand U9343 (N_9343,N_5685,N_4658);
nor U9344 (N_9344,N_757,N_5752);
or U9345 (N_9345,N_2201,N_3122);
and U9346 (N_9346,N_3064,N_2680);
and U9347 (N_9347,N_1897,N_4132);
nor U9348 (N_9348,N_1671,N_1840);
nor U9349 (N_9349,N_85,N_4652);
xor U9350 (N_9350,N_282,N_4819);
and U9351 (N_9351,N_2833,N_4819);
nor U9352 (N_9352,N_5887,N_4966);
nor U9353 (N_9353,N_3157,N_2072);
nand U9354 (N_9354,N_2593,N_1842);
nor U9355 (N_9355,N_4740,N_852);
nand U9356 (N_9356,N_4512,N_5008);
or U9357 (N_9357,N_4001,N_5872);
or U9358 (N_9358,N_2152,N_2793);
nor U9359 (N_9359,N_3552,N_5478);
and U9360 (N_9360,N_5796,N_5385);
and U9361 (N_9361,N_5904,N_5965);
xor U9362 (N_9362,N_1916,N_702);
nor U9363 (N_9363,N_201,N_3755);
xnor U9364 (N_9364,N_2495,N_2065);
nand U9365 (N_9365,N_4573,N_5949);
and U9366 (N_9366,N_5174,N_5836);
xor U9367 (N_9367,N_4448,N_2355);
nor U9368 (N_9368,N_5533,N_1611);
and U9369 (N_9369,N_493,N_2379);
and U9370 (N_9370,N_4974,N_3673);
and U9371 (N_9371,N_5087,N_3594);
or U9372 (N_9372,N_1244,N_5330);
nand U9373 (N_9373,N_3165,N_2313);
nand U9374 (N_9374,N_5378,N_547);
nand U9375 (N_9375,N_4284,N_1002);
nand U9376 (N_9376,N_3604,N_4772);
xor U9377 (N_9377,N_3458,N_5633);
or U9378 (N_9378,N_2744,N_2562);
nor U9379 (N_9379,N_5564,N_5100);
xnor U9380 (N_9380,N_4677,N_5581);
xnor U9381 (N_9381,N_3178,N_1532);
nor U9382 (N_9382,N_3642,N_2773);
nand U9383 (N_9383,N_4241,N_4421);
nor U9384 (N_9384,N_4763,N_3734);
or U9385 (N_9385,N_4122,N_3844);
xnor U9386 (N_9386,N_3405,N_1893);
or U9387 (N_9387,N_470,N_1613);
and U9388 (N_9388,N_5880,N_878);
and U9389 (N_9389,N_2863,N_1050);
or U9390 (N_9390,N_5843,N_3029);
or U9391 (N_9391,N_975,N_3973);
nor U9392 (N_9392,N_265,N_5451);
nand U9393 (N_9393,N_4540,N_803);
and U9394 (N_9394,N_4654,N_1477);
nor U9395 (N_9395,N_4247,N_2055);
nand U9396 (N_9396,N_816,N_3367);
or U9397 (N_9397,N_1383,N_5815);
and U9398 (N_9398,N_5090,N_3209);
or U9399 (N_9399,N_4328,N_2307);
xnor U9400 (N_9400,N_1161,N_2723);
nor U9401 (N_9401,N_5667,N_1749);
nand U9402 (N_9402,N_3400,N_1489);
nand U9403 (N_9403,N_2509,N_4854);
and U9404 (N_9404,N_1478,N_5743);
xnor U9405 (N_9405,N_1826,N_3182);
or U9406 (N_9406,N_2845,N_3196);
nand U9407 (N_9407,N_2535,N_4935);
or U9408 (N_9408,N_5249,N_5661);
nor U9409 (N_9409,N_3602,N_3522);
and U9410 (N_9410,N_3998,N_1924);
and U9411 (N_9411,N_844,N_4840);
or U9412 (N_9412,N_226,N_4911);
nand U9413 (N_9413,N_5659,N_2927);
xor U9414 (N_9414,N_605,N_4196);
or U9415 (N_9415,N_406,N_578);
or U9416 (N_9416,N_1231,N_372);
xnor U9417 (N_9417,N_283,N_3000);
xnor U9418 (N_9418,N_5299,N_850);
or U9419 (N_9419,N_2120,N_5842);
nand U9420 (N_9420,N_2535,N_3162);
xnor U9421 (N_9421,N_4816,N_4394);
or U9422 (N_9422,N_2342,N_3314);
xnor U9423 (N_9423,N_5052,N_1484);
and U9424 (N_9424,N_4930,N_451);
nor U9425 (N_9425,N_2248,N_676);
or U9426 (N_9426,N_552,N_3279);
nand U9427 (N_9427,N_366,N_5566);
nand U9428 (N_9428,N_1489,N_5763);
xor U9429 (N_9429,N_3073,N_3674);
nor U9430 (N_9430,N_4443,N_2423);
nor U9431 (N_9431,N_2748,N_3773);
nand U9432 (N_9432,N_1085,N_5687);
nor U9433 (N_9433,N_3342,N_359);
xnor U9434 (N_9434,N_5917,N_536);
and U9435 (N_9435,N_992,N_944);
or U9436 (N_9436,N_3772,N_945);
nor U9437 (N_9437,N_4622,N_3519);
nor U9438 (N_9438,N_5604,N_2675);
nand U9439 (N_9439,N_4806,N_4843);
nand U9440 (N_9440,N_533,N_5501);
nand U9441 (N_9441,N_717,N_3410);
and U9442 (N_9442,N_2788,N_2359);
xor U9443 (N_9443,N_2348,N_100);
and U9444 (N_9444,N_1158,N_2338);
or U9445 (N_9445,N_462,N_2356);
nor U9446 (N_9446,N_3565,N_668);
xor U9447 (N_9447,N_2117,N_137);
nand U9448 (N_9448,N_4386,N_3501);
or U9449 (N_9449,N_1287,N_3261);
xor U9450 (N_9450,N_1513,N_3410);
nand U9451 (N_9451,N_856,N_2964);
nand U9452 (N_9452,N_3292,N_4173);
xnor U9453 (N_9453,N_106,N_2233);
or U9454 (N_9454,N_1660,N_1557);
and U9455 (N_9455,N_3992,N_3614);
and U9456 (N_9456,N_3285,N_1064);
nor U9457 (N_9457,N_932,N_2507);
xor U9458 (N_9458,N_1259,N_4070);
or U9459 (N_9459,N_3184,N_3908);
and U9460 (N_9460,N_904,N_2600);
and U9461 (N_9461,N_734,N_3906);
or U9462 (N_9462,N_675,N_1713);
nor U9463 (N_9463,N_5954,N_5312);
or U9464 (N_9464,N_3022,N_5337);
or U9465 (N_9465,N_299,N_2988);
xor U9466 (N_9466,N_2407,N_69);
nand U9467 (N_9467,N_702,N_5617);
nand U9468 (N_9468,N_5797,N_1189);
nand U9469 (N_9469,N_1639,N_946);
and U9470 (N_9470,N_4217,N_4551);
nand U9471 (N_9471,N_2118,N_2559);
or U9472 (N_9472,N_2968,N_1287);
or U9473 (N_9473,N_5520,N_5335);
nor U9474 (N_9474,N_1627,N_3850);
and U9475 (N_9475,N_2526,N_1519);
or U9476 (N_9476,N_1498,N_3679);
xor U9477 (N_9477,N_3504,N_1013);
nor U9478 (N_9478,N_4189,N_602);
xnor U9479 (N_9479,N_996,N_2398);
nor U9480 (N_9480,N_3129,N_1525);
nand U9481 (N_9481,N_4985,N_4438);
and U9482 (N_9482,N_4190,N_1972);
nand U9483 (N_9483,N_5058,N_2484);
nand U9484 (N_9484,N_4118,N_2342);
nand U9485 (N_9485,N_5373,N_2377);
nand U9486 (N_9486,N_609,N_4371);
and U9487 (N_9487,N_4042,N_4857);
nor U9488 (N_9488,N_429,N_3762);
nor U9489 (N_9489,N_952,N_1635);
nand U9490 (N_9490,N_1816,N_877);
nand U9491 (N_9491,N_3644,N_2306);
xnor U9492 (N_9492,N_4564,N_3023);
nand U9493 (N_9493,N_1498,N_2310);
nand U9494 (N_9494,N_938,N_873);
nand U9495 (N_9495,N_4441,N_5813);
xor U9496 (N_9496,N_4241,N_3063);
or U9497 (N_9497,N_5486,N_4453);
nand U9498 (N_9498,N_2609,N_2266);
nor U9499 (N_9499,N_2039,N_4336);
nor U9500 (N_9500,N_624,N_4578);
xnor U9501 (N_9501,N_4330,N_2823);
xor U9502 (N_9502,N_2182,N_1201);
and U9503 (N_9503,N_4391,N_4231);
nand U9504 (N_9504,N_5558,N_2530);
nand U9505 (N_9505,N_184,N_3152);
nand U9506 (N_9506,N_3775,N_2660);
nand U9507 (N_9507,N_3100,N_5756);
xor U9508 (N_9508,N_3023,N_3192);
and U9509 (N_9509,N_2108,N_5088);
and U9510 (N_9510,N_4656,N_433);
or U9511 (N_9511,N_1835,N_5029);
nand U9512 (N_9512,N_5576,N_4545);
or U9513 (N_9513,N_5973,N_1263);
or U9514 (N_9514,N_1139,N_678);
or U9515 (N_9515,N_4496,N_703);
nand U9516 (N_9516,N_1576,N_1714);
and U9517 (N_9517,N_2602,N_3284);
nor U9518 (N_9518,N_2624,N_4453);
xnor U9519 (N_9519,N_4671,N_4842);
and U9520 (N_9520,N_2757,N_2164);
nand U9521 (N_9521,N_1312,N_3777);
xor U9522 (N_9522,N_37,N_2171);
xor U9523 (N_9523,N_4122,N_2068);
nor U9524 (N_9524,N_829,N_5213);
and U9525 (N_9525,N_1292,N_5136);
or U9526 (N_9526,N_3531,N_3296);
xnor U9527 (N_9527,N_4668,N_1141);
nand U9528 (N_9528,N_3404,N_90);
xor U9529 (N_9529,N_3167,N_3923);
and U9530 (N_9530,N_2586,N_20);
or U9531 (N_9531,N_5438,N_3386);
nand U9532 (N_9532,N_2953,N_816);
xor U9533 (N_9533,N_1467,N_639);
xnor U9534 (N_9534,N_3913,N_2536);
and U9535 (N_9535,N_345,N_779);
nand U9536 (N_9536,N_5842,N_2491);
and U9537 (N_9537,N_1142,N_2814);
or U9538 (N_9538,N_3404,N_5984);
or U9539 (N_9539,N_3345,N_3875);
nor U9540 (N_9540,N_4368,N_5331);
and U9541 (N_9541,N_5847,N_5254);
nand U9542 (N_9542,N_2191,N_5053);
or U9543 (N_9543,N_4009,N_3449);
or U9544 (N_9544,N_3078,N_3739);
xnor U9545 (N_9545,N_5514,N_5845);
nor U9546 (N_9546,N_3298,N_518);
xnor U9547 (N_9547,N_5453,N_1715);
xor U9548 (N_9548,N_2873,N_2380);
and U9549 (N_9549,N_4691,N_1463);
nand U9550 (N_9550,N_571,N_695);
nand U9551 (N_9551,N_3593,N_3972);
nand U9552 (N_9552,N_5621,N_1806);
and U9553 (N_9553,N_1440,N_2385);
xor U9554 (N_9554,N_3665,N_1818);
nor U9555 (N_9555,N_5507,N_1480);
nor U9556 (N_9556,N_5569,N_1414);
and U9557 (N_9557,N_373,N_1496);
nand U9558 (N_9558,N_4710,N_5336);
or U9559 (N_9559,N_3796,N_988);
nor U9560 (N_9560,N_4453,N_1212);
nor U9561 (N_9561,N_613,N_5937);
or U9562 (N_9562,N_4516,N_3910);
xnor U9563 (N_9563,N_2061,N_3028);
and U9564 (N_9564,N_1204,N_4853);
and U9565 (N_9565,N_132,N_4850);
or U9566 (N_9566,N_5925,N_5946);
nor U9567 (N_9567,N_1285,N_3272);
or U9568 (N_9568,N_2494,N_313);
nor U9569 (N_9569,N_4535,N_2003);
nand U9570 (N_9570,N_1512,N_1084);
nor U9571 (N_9571,N_1978,N_4842);
and U9572 (N_9572,N_3928,N_5708);
nor U9573 (N_9573,N_5858,N_5404);
xnor U9574 (N_9574,N_1173,N_4088);
xor U9575 (N_9575,N_3343,N_4440);
xor U9576 (N_9576,N_1565,N_3803);
nand U9577 (N_9577,N_1759,N_4866);
nand U9578 (N_9578,N_3648,N_3806);
xor U9579 (N_9579,N_5167,N_4912);
and U9580 (N_9580,N_2186,N_70);
and U9581 (N_9581,N_4118,N_1767);
nor U9582 (N_9582,N_1630,N_3753);
nor U9583 (N_9583,N_3083,N_2593);
nor U9584 (N_9584,N_3447,N_3280);
and U9585 (N_9585,N_3415,N_3535);
nor U9586 (N_9586,N_3794,N_5983);
nor U9587 (N_9587,N_591,N_1768);
and U9588 (N_9588,N_4215,N_3215);
xnor U9589 (N_9589,N_3181,N_3040);
nand U9590 (N_9590,N_3289,N_4169);
nor U9591 (N_9591,N_4858,N_2268);
and U9592 (N_9592,N_365,N_2722);
nor U9593 (N_9593,N_1108,N_175);
and U9594 (N_9594,N_1807,N_2088);
xnor U9595 (N_9595,N_2437,N_5151);
nor U9596 (N_9596,N_1830,N_3780);
nor U9597 (N_9597,N_4429,N_1793);
and U9598 (N_9598,N_2568,N_4955);
nand U9599 (N_9599,N_5240,N_1617);
and U9600 (N_9600,N_5164,N_3117);
xor U9601 (N_9601,N_1591,N_4314);
or U9602 (N_9602,N_4357,N_1647);
nand U9603 (N_9603,N_4833,N_2000);
nand U9604 (N_9604,N_4243,N_903);
nand U9605 (N_9605,N_5570,N_4029);
and U9606 (N_9606,N_2517,N_5181);
or U9607 (N_9607,N_2946,N_5331);
and U9608 (N_9608,N_2162,N_3811);
or U9609 (N_9609,N_4661,N_4402);
or U9610 (N_9610,N_3708,N_5479);
and U9611 (N_9611,N_4420,N_2375);
or U9612 (N_9612,N_3829,N_5098);
or U9613 (N_9613,N_238,N_1950);
and U9614 (N_9614,N_1146,N_3140);
nor U9615 (N_9615,N_5032,N_3088);
nor U9616 (N_9616,N_10,N_2914);
nand U9617 (N_9617,N_1508,N_1237);
nand U9618 (N_9618,N_2728,N_4289);
nand U9619 (N_9619,N_4952,N_3971);
nor U9620 (N_9620,N_4380,N_1271);
or U9621 (N_9621,N_1803,N_4582);
or U9622 (N_9622,N_2449,N_1174);
and U9623 (N_9623,N_3439,N_457);
nor U9624 (N_9624,N_5806,N_4200);
or U9625 (N_9625,N_2441,N_48);
nor U9626 (N_9626,N_60,N_4997);
and U9627 (N_9627,N_2606,N_3852);
and U9628 (N_9628,N_5335,N_1723);
or U9629 (N_9629,N_1589,N_870);
and U9630 (N_9630,N_1067,N_576);
or U9631 (N_9631,N_5647,N_5153);
nor U9632 (N_9632,N_5200,N_3841);
and U9633 (N_9633,N_4240,N_1513);
or U9634 (N_9634,N_5106,N_4342);
nor U9635 (N_9635,N_4415,N_291);
or U9636 (N_9636,N_58,N_128);
or U9637 (N_9637,N_2573,N_4525);
nand U9638 (N_9638,N_1476,N_1775);
and U9639 (N_9639,N_846,N_1423);
or U9640 (N_9640,N_5300,N_3001);
nand U9641 (N_9641,N_1357,N_5833);
nor U9642 (N_9642,N_3384,N_4556);
nand U9643 (N_9643,N_5269,N_5173);
nand U9644 (N_9644,N_5972,N_5238);
xnor U9645 (N_9645,N_645,N_17);
or U9646 (N_9646,N_3873,N_5990);
and U9647 (N_9647,N_752,N_2674);
nor U9648 (N_9648,N_2695,N_2290);
and U9649 (N_9649,N_735,N_3269);
nor U9650 (N_9650,N_5931,N_360);
nor U9651 (N_9651,N_2881,N_3843);
xnor U9652 (N_9652,N_5743,N_2416);
nand U9653 (N_9653,N_4086,N_926);
xnor U9654 (N_9654,N_1066,N_4386);
nand U9655 (N_9655,N_3165,N_1738);
or U9656 (N_9656,N_1242,N_1249);
xnor U9657 (N_9657,N_4535,N_3583);
or U9658 (N_9658,N_5379,N_2557);
and U9659 (N_9659,N_2051,N_2818);
nor U9660 (N_9660,N_4093,N_3418);
nand U9661 (N_9661,N_110,N_3091);
or U9662 (N_9662,N_3001,N_443);
or U9663 (N_9663,N_4785,N_3728);
nor U9664 (N_9664,N_3071,N_2893);
nor U9665 (N_9665,N_100,N_2389);
xor U9666 (N_9666,N_3678,N_2677);
or U9667 (N_9667,N_452,N_4967);
and U9668 (N_9668,N_2541,N_4432);
and U9669 (N_9669,N_5351,N_3493);
nand U9670 (N_9670,N_4217,N_4525);
or U9671 (N_9671,N_2753,N_5319);
or U9672 (N_9672,N_2929,N_5905);
nor U9673 (N_9673,N_3643,N_5724);
xnor U9674 (N_9674,N_3934,N_4885);
nor U9675 (N_9675,N_1734,N_4486);
and U9676 (N_9676,N_4932,N_4959);
and U9677 (N_9677,N_5844,N_4402);
or U9678 (N_9678,N_3398,N_5496);
and U9679 (N_9679,N_2030,N_2724);
nand U9680 (N_9680,N_5576,N_5053);
or U9681 (N_9681,N_779,N_147);
or U9682 (N_9682,N_4133,N_5846);
nand U9683 (N_9683,N_752,N_3190);
and U9684 (N_9684,N_164,N_773);
and U9685 (N_9685,N_3990,N_2986);
or U9686 (N_9686,N_2417,N_1176);
nand U9687 (N_9687,N_3667,N_3046);
and U9688 (N_9688,N_5952,N_2875);
or U9689 (N_9689,N_3884,N_1619);
xor U9690 (N_9690,N_2671,N_1564);
nor U9691 (N_9691,N_4729,N_211);
xor U9692 (N_9692,N_1055,N_1873);
or U9693 (N_9693,N_2088,N_3226);
xnor U9694 (N_9694,N_3335,N_4711);
nand U9695 (N_9695,N_1833,N_5819);
nor U9696 (N_9696,N_3780,N_287);
or U9697 (N_9697,N_5435,N_5971);
nor U9698 (N_9698,N_5225,N_1842);
xnor U9699 (N_9699,N_4843,N_1508);
xnor U9700 (N_9700,N_4925,N_3282);
nor U9701 (N_9701,N_293,N_5550);
nor U9702 (N_9702,N_4684,N_1049);
nand U9703 (N_9703,N_3114,N_5022);
nor U9704 (N_9704,N_4427,N_1035);
xnor U9705 (N_9705,N_5659,N_3452);
nor U9706 (N_9706,N_1677,N_4160);
xnor U9707 (N_9707,N_5741,N_3446);
nand U9708 (N_9708,N_2002,N_4314);
and U9709 (N_9709,N_2661,N_1725);
nor U9710 (N_9710,N_5341,N_3552);
nand U9711 (N_9711,N_4795,N_5223);
nand U9712 (N_9712,N_116,N_1171);
nor U9713 (N_9713,N_1228,N_68);
nand U9714 (N_9714,N_5392,N_2263);
and U9715 (N_9715,N_1202,N_4594);
or U9716 (N_9716,N_335,N_4065);
nor U9717 (N_9717,N_2581,N_3879);
and U9718 (N_9718,N_4887,N_5859);
and U9719 (N_9719,N_2441,N_754);
xnor U9720 (N_9720,N_5584,N_4027);
nor U9721 (N_9721,N_916,N_2875);
nor U9722 (N_9722,N_5592,N_1043);
nor U9723 (N_9723,N_3581,N_4878);
nor U9724 (N_9724,N_5590,N_2136);
or U9725 (N_9725,N_3699,N_2515);
and U9726 (N_9726,N_5094,N_5942);
and U9727 (N_9727,N_261,N_2956);
nor U9728 (N_9728,N_5923,N_4129);
or U9729 (N_9729,N_3548,N_910);
or U9730 (N_9730,N_2830,N_5749);
xor U9731 (N_9731,N_2555,N_3976);
nand U9732 (N_9732,N_4131,N_5969);
nor U9733 (N_9733,N_4852,N_4709);
nand U9734 (N_9734,N_1899,N_651);
or U9735 (N_9735,N_1206,N_3824);
nor U9736 (N_9736,N_2906,N_4972);
xor U9737 (N_9737,N_5607,N_474);
xnor U9738 (N_9738,N_616,N_4090);
or U9739 (N_9739,N_4161,N_2330);
and U9740 (N_9740,N_4650,N_4638);
or U9741 (N_9741,N_4381,N_1740);
or U9742 (N_9742,N_5935,N_279);
or U9743 (N_9743,N_1965,N_4775);
nor U9744 (N_9744,N_2885,N_5040);
nor U9745 (N_9745,N_5434,N_4519);
or U9746 (N_9746,N_4013,N_5386);
nor U9747 (N_9747,N_5811,N_1277);
xnor U9748 (N_9748,N_2293,N_5770);
nor U9749 (N_9749,N_2933,N_5100);
or U9750 (N_9750,N_5085,N_3420);
nand U9751 (N_9751,N_1666,N_760);
nor U9752 (N_9752,N_5454,N_5654);
nor U9753 (N_9753,N_3477,N_320);
or U9754 (N_9754,N_5338,N_773);
or U9755 (N_9755,N_4971,N_4441);
or U9756 (N_9756,N_4796,N_732);
xor U9757 (N_9757,N_709,N_2408);
xor U9758 (N_9758,N_1371,N_5599);
or U9759 (N_9759,N_4315,N_4666);
xnor U9760 (N_9760,N_5279,N_2280);
and U9761 (N_9761,N_3209,N_5571);
nand U9762 (N_9762,N_4023,N_2332);
nor U9763 (N_9763,N_893,N_5940);
or U9764 (N_9764,N_5688,N_3388);
or U9765 (N_9765,N_2319,N_5786);
nand U9766 (N_9766,N_4911,N_4743);
nand U9767 (N_9767,N_4984,N_3090);
and U9768 (N_9768,N_4066,N_4647);
and U9769 (N_9769,N_1244,N_913);
and U9770 (N_9770,N_3103,N_5099);
nor U9771 (N_9771,N_5305,N_1480);
xnor U9772 (N_9772,N_1056,N_3021);
xnor U9773 (N_9773,N_4935,N_5629);
and U9774 (N_9774,N_5868,N_794);
nand U9775 (N_9775,N_2452,N_5701);
xor U9776 (N_9776,N_3264,N_4907);
or U9777 (N_9777,N_5579,N_255);
nand U9778 (N_9778,N_1559,N_4662);
and U9779 (N_9779,N_5740,N_5916);
xnor U9780 (N_9780,N_2629,N_1714);
nand U9781 (N_9781,N_3806,N_2413);
and U9782 (N_9782,N_3603,N_4408);
nor U9783 (N_9783,N_5301,N_3321);
xnor U9784 (N_9784,N_5748,N_3058);
nor U9785 (N_9785,N_2978,N_387);
xnor U9786 (N_9786,N_2848,N_4921);
xor U9787 (N_9787,N_1660,N_396);
nand U9788 (N_9788,N_720,N_5566);
nor U9789 (N_9789,N_1892,N_3701);
nor U9790 (N_9790,N_930,N_2514);
and U9791 (N_9791,N_1252,N_2360);
xor U9792 (N_9792,N_1362,N_1342);
nor U9793 (N_9793,N_2567,N_3837);
nand U9794 (N_9794,N_3278,N_1130);
nand U9795 (N_9795,N_5357,N_4445);
nor U9796 (N_9796,N_2458,N_1179);
nand U9797 (N_9797,N_3256,N_1836);
and U9798 (N_9798,N_2018,N_3955);
and U9799 (N_9799,N_1555,N_2655);
and U9800 (N_9800,N_2687,N_1894);
xnor U9801 (N_9801,N_1807,N_1656);
nor U9802 (N_9802,N_3706,N_19);
nand U9803 (N_9803,N_2090,N_3465);
nand U9804 (N_9804,N_3656,N_3142);
xor U9805 (N_9805,N_374,N_885);
nand U9806 (N_9806,N_581,N_2257);
and U9807 (N_9807,N_4289,N_2965);
and U9808 (N_9808,N_3950,N_4628);
and U9809 (N_9809,N_363,N_3058);
or U9810 (N_9810,N_2225,N_4810);
nand U9811 (N_9811,N_5267,N_3719);
nand U9812 (N_9812,N_956,N_50);
or U9813 (N_9813,N_2984,N_1931);
nand U9814 (N_9814,N_4931,N_4382);
and U9815 (N_9815,N_992,N_84);
nor U9816 (N_9816,N_989,N_4838);
and U9817 (N_9817,N_4123,N_2181);
xor U9818 (N_9818,N_5214,N_2811);
or U9819 (N_9819,N_2753,N_4159);
nand U9820 (N_9820,N_5701,N_3720);
and U9821 (N_9821,N_44,N_2344);
and U9822 (N_9822,N_4629,N_1332);
nand U9823 (N_9823,N_4774,N_4265);
nand U9824 (N_9824,N_5759,N_814);
nand U9825 (N_9825,N_5897,N_3850);
nand U9826 (N_9826,N_2904,N_4700);
or U9827 (N_9827,N_4085,N_2293);
nor U9828 (N_9828,N_4870,N_306);
xor U9829 (N_9829,N_351,N_1396);
nand U9830 (N_9830,N_4395,N_4421);
nor U9831 (N_9831,N_2556,N_181);
and U9832 (N_9832,N_3674,N_2878);
or U9833 (N_9833,N_5575,N_1526);
and U9834 (N_9834,N_1063,N_2536);
and U9835 (N_9835,N_3262,N_2101);
xnor U9836 (N_9836,N_5572,N_1337);
nor U9837 (N_9837,N_3026,N_3352);
nand U9838 (N_9838,N_3610,N_4751);
or U9839 (N_9839,N_2837,N_4320);
nand U9840 (N_9840,N_5487,N_3288);
xor U9841 (N_9841,N_2734,N_3066);
nor U9842 (N_9842,N_2408,N_2104);
xnor U9843 (N_9843,N_3340,N_3835);
nor U9844 (N_9844,N_3082,N_2214);
and U9845 (N_9845,N_4897,N_3982);
nor U9846 (N_9846,N_3276,N_5499);
xnor U9847 (N_9847,N_4560,N_432);
xnor U9848 (N_9848,N_4824,N_1676);
xor U9849 (N_9849,N_4604,N_5038);
xor U9850 (N_9850,N_2275,N_254);
or U9851 (N_9851,N_1542,N_2033);
nand U9852 (N_9852,N_5629,N_4321);
nor U9853 (N_9853,N_300,N_1281);
nor U9854 (N_9854,N_2541,N_3300);
or U9855 (N_9855,N_872,N_3117);
and U9856 (N_9856,N_3223,N_1730);
xor U9857 (N_9857,N_5313,N_5452);
nand U9858 (N_9858,N_5630,N_2668);
and U9859 (N_9859,N_872,N_302);
nand U9860 (N_9860,N_3873,N_654);
nand U9861 (N_9861,N_1499,N_2421);
and U9862 (N_9862,N_4412,N_5416);
and U9863 (N_9863,N_2639,N_276);
nor U9864 (N_9864,N_5045,N_303);
nand U9865 (N_9865,N_2303,N_5198);
or U9866 (N_9866,N_4571,N_5033);
xnor U9867 (N_9867,N_136,N_5756);
or U9868 (N_9868,N_75,N_3538);
nor U9869 (N_9869,N_303,N_4288);
and U9870 (N_9870,N_3443,N_3977);
nor U9871 (N_9871,N_4932,N_4693);
and U9872 (N_9872,N_1161,N_1615);
and U9873 (N_9873,N_3428,N_105);
xor U9874 (N_9874,N_3613,N_4295);
nand U9875 (N_9875,N_3315,N_3222);
nor U9876 (N_9876,N_3419,N_4986);
nand U9877 (N_9877,N_4124,N_289);
xor U9878 (N_9878,N_1829,N_2518);
xor U9879 (N_9879,N_3931,N_2884);
xor U9880 (N_9880,N_5118,N_1098);
and U9881 (N_9881,N_3997,N_5576);
and U9882 (N_9882,N_884,N_5892);
and U9883 (N_9883,N_4605,N_3937);
or U9884 (N_9884,N_2333,N_3619);
nor U9885 (N_9885,N_85,N_4381);
nor U9886 (N_9886,N_2284,N_5248);
nor U9887 (N_9887,N_4689,N_647);
and U9888 (N_9888,N_1944,N_5027);
and U9889 (N_9889,N_3768,N_5660);
nand U9890 (N_9890,N_1829,N_4230);
nor U9891 (N_9891,N_4287,N_5922);
xnor U9892 (N_9892,N_4582,N_3511);
or U9893 (N_9893,N_1534,N_1423);
or U9894 (N_9894,N_3254,N_5641);
or U9895 (N_9895,N_4202,N_3940);
and U9896 (N_9896,N_3367,N_4180);
nor U9897 (N_9897,N_2305,N_1022);
nor U9898 (N_9898,N_1450,N_4591);
xnor U9899 (N_9899,N_3582,N_422);
nor U9900 (N_9900,N_4669,N_1636);
xor U9901 (N_9901,N_3833,N_2131);
xnor U9902 (N_9902,N_5059,N_5738);
and U9903 (N_9903,N_881,N_5041);
nor U9904 (N_9904,N_5824,N_2260);
nor U9905 (N_9905,N_3013,N_4519);
nor U9906 (N_9906,N_2947,N_1064);
or U9907 (N_9907,N_3411,N_3586);
nand U9908 (N_9908,N_846,N_4750);
nand U9909 (N_9909,N_2462,N_2568);
and U9910 (N_9910,N_2217,N_3876);
nand U9911 (N_9911,N_56,N_5689);
xor U9912 (N_9912,N_4168,N_4182);
nor U9913 (N_9913,N_5834,N_1303);
xor U9914 (N_9914,N_3739,N_2721);
nor U9915 (N_9915,N_5672,N_5101);
nor U9916 (N_9916,N_5056,N_4525);
and U9917 (N_9917,N_5577,N_5902);
or U9918 (N_9918,N_5592,N_2141);
or U9919 (N_9919,N_4002,N_991);
nor U9920 (N_9920,N_822,N_67);
nand U9921 (N_9921,N_2312,N_5124);
or U9922 (N_9922,N_3283,N_724);
nor U9923 (N_9923,N_5147,N_48);
nand U9924 (N_9924,N_5759,N_1426);
nor U9925 (N_9925,N_2274,N_1009);
xor U9926 (N_9926,N_3628,N_2393);
and U9927 (N_9927,N_2943,N_4243);
xor U9928 (N_9928,N_1927,N_1597);
nor U9929 (N_9929,N_4095,N_3855);
xor U9930 (N_9930,N_1971,N_1178);
xor U9931 (N_9931,N_4407,N_1107);
and U9932 (N_9932,N_257,N_1200);
nand U9933 (N_9933,N_3433,N_1834);
nand U9934 (N_9934,N_5670,N_5196);
xnor U9935 (N_9935,N_576,N_4804);
nor U9936 (N_9936,N_2808,N_3055);
or U9937 (N_9937,N_2412,N_3145);
nor U9938 (N_9938,N_4176,N_5671);
xnor U9939 (N_9939,N_3361,N_3088);
nor U9940 (N_9940,N_2578,N_3348);
nor U9941 (N_9941,N_5778,N_2500);
nand U9942 (N_9942,N_1147,N_3070);
nand U9943 (N_9943,N_4788,N_5682);
nor U9944 (N_9944,N_408,N_3558);
nor U9945 (N_9945,N_3928,N_2293);
or U9946 (N_9946,N_4525,N_5898);
nand U9947 (N_9947,N_1214,N_272);
nor U9948 (N_9948,N_726,N_4696);
nor U9949 (N_9949,N_5145,N_3631);
nor U9950 (N_9950,N_4302,N_290);
nor U9951 (N_9951,N_5030,N_80);
xnor U9952 (N_9952,N_5931,N_5172);
nor U9953 (N_9953,N_3197,N_3435);
or U9954 (N_9954,N_5396,N_4092);
nand U9955 (N_9955,N_1646,N_20);
or U9956 (N_9956,N_5220,N_4912);
nand U9957 (N_9957,N_433,N_1315);
nor U9958 (N_9958,N_1864,N_1673);
and U9959 (N_9959,N_5858,N_4966);
or U9960 (N_9960,N_3882,N_5430);
xor U9961 (N_9961,N_3809,N_1129);
xnor U9962 (N_9962,N_3030,N_3237);
and U9963 (N_9963,N_5131,N_1464);
and U9964 (N_9964,N_1238,N_2900);
xor U9965 (N_9965,N_4507,N_125);
or U9966 (N_9966,N_2412,N_1728);
nor U9967 (N_9967,N_5312,N_4681);
or U9968 (N_9968,N_444,N_5508);
xnor U9969 (N_9969,N_2976,N_1606);
nand U9970 (N_9970,N_3196,N_1784);
xor U9971 (N_9971,N_1104,N_436);
or U9972 (N_9972,N_351,N_609);
nand U9973 (N_9973,N_1528,N_3890);
xnor U9974 (N_9974,N_4,N_3641);
and U9975 (N_9975,N_509,N_4494);
and U9976 (N_9976,N_306,N_154);
xnor U9977 (N_9977,N_2376,N_5279);
and U9978 (N_9978,N_5682,N_4671);
or U9979 (N_9979,N_5486,N_3400);
nand U9980 (N_9980,N_736,N_1595);
or U9981 (N_9981,N_4465,N_1526);
nand U9982 (N_9982,N_1290,N_3572);
nor U9983 (N_9983,N_347,N_4991);
xor U9984 (N_9984,N_2720,N_4944);
nand U9985 (N_9985,N_613,N_320);
or U9986 (N_9986,N_4782,N_5450);
or U9987 (N_9987,N_5726,N_1386);
nor U9988 (N_9988,N_1364,N_934);
or U9989 (N_9989,N_149,N_56);
nand U9990 (N_9990,N_85,N_5760);
or U9991 (N_9991,N_5849,N_541);
nor U9992 (N_9992,N_655,N_272);
nand U9993 (N_9993,N_1140,N_5429);
and U9994 (N_9994,N_1445,N_4806);
nand U9995 (N_9995,N_5504,N_668);
nand U9996 (N_9996,N_995,N_2211);
and U9997 (N_9997,N_1428,N_3000);
and U9998 (N_9998,N_2607,N_128);
or U9999 (N_9999,N_1090,N_912);
and U10000 (N_10000,N_5238,N_4882);
nor U10001 (N_10001,N_2546,N_3556);
or U10002 (N_10002,N_5894,N_103);
nand U10003 (N_10003,N_3706,N_758);
and U10004 (N_10004,N_3958,N_2431);
nor U10005 (N_10005,N_222,N_2646);
nand U10006 (N_10006,N_2839,N_654);
xor U10007 (N_10007,N_4158,N_5125);
nand U10008 (N_10008,N_4145,N_3400);
or U10009 (N_10009,N_5828,N_4176);
and U10010 (N_10010,N_3520,N_5306);
xor U10011 (N_10011,N_3270,N_2165);
xor U10012 (N_10012,N_1172,N_5160);
or U10013 (N_10013,N_4776,N_4035);
nor U10014 (N_10014,N_1893,N_2188);
xnor U10015 (N_10015,N_2044,N_2145);
xor U10016 (N_10016,N_5182,N_542);
xor U10017 (N_10017,N_4318,N_920);
or U10018 (N_10018,N_3638,N_5497);
xor U10019 (N_10019,N_4578,N_5613);
nor U10020 (N_10020,N_1902,N_5885);
xor U10021 (N_10021,N_2932,N_1099);
or U10022 (N_10022,N_533,N_3614);
xnor U10023 (N_10023,N_833,N_2615);
and U10024 (N_10024,N_656,N_5839);
and U10025 (N_10025,N_4099,N_2699);
nor U10026 (N_10026,N_496,N_426);
nand U10027 (N_10027,N_4502,N_2479);
nand U10028 (N_10028,N_3222,N_5936);
nand U10029 (N_10029,N_5914,N_4254);
nand U10030 (N_10030,N_5022,N_4000);
or U10031 (N_10031,N_1566,N_2059);
and U10032 (N_10032,N_2807,N_5686);
xor U10033 (N_10033,N_272,N_5118);
xnor U10034 (N_10034,N_822,N_2998);
or U10035 (N_10035,N_5822,N_3459);
xor U10036 (N_10036,N_4363,N_2940);
or U10037 (N_10037,N_962,N_2362);
or U10038 (N_10038,N_4680,N_2844);
or U10039 (N_10039,N_4102,N_90);
nor U10040 (N_10040,N_2700,N_1384);
or U10041 (N_10041,N_2588,N_2736);
and U10042 (N_10042,N_4599,N_3553);
xnor U10043 (N_10043,N_5172,N_103);
and U10044 (N_10044,N_2877,N_3328);
and U10045 (N_10045,N_1316,N_3894);
nor U10046 (N_10046,N_294,N_3545);
nor U10047 (N_10047,N_1112,N_4715);
nand U10048 (N_10048,N_4765,N_4054);
or U10049 (N_10049,N_45,N_3618);
nor U10050 (N_10050,N_3773,N_2475);
and U10051 (N_10051,N_3794,N_735);
or U10052 (N_10052,N_2525,N_5664);
nand U10053 (N_10053,N_1286,N_3071);
nor U10054 (N_10054,N_4467,N_4559);
xnor U10055 (N_10055,N_3646,N_3354);
nor U10056 (N_10056,N_4936,N_718);
or U10057 (N_10057,N_1851,N_1409);
xnor U10058 (N_10058,N_1940,N_3059);
or U10059 (N_10059,N_4112,N_3332);
xnor U10060 (N_10060,N_608,N_2170);
xor U10061 (N_10061,N_3861,N_2988);
nor U10062 (N_10062,N_3488,N_671);
xnor U10063 (N_10063,N_3955,N_5486);
nor U10064 (N_10064,N_795,N_4586);
nand U10065 (N_10065,N_3446,N_4235);
and U10066 (N_10066,N_2241,N_426);
nor U10067 (N_10067,N_2690,N_4770);
nor U10068 (N_10068,N_1959,N_3990);
or U10069 (N_10069,N_1980,N_4643);
nand U10070 (N_10070,N_4030,N_1761);
xor U10071 (N_10071,N_5354,N_5231);
nand U10072 (N_10072,N_2912,N_750);
and U10073 (N_10073,N_2154,N_4098);
or U10074 (N_10074,N_3554,N_5499);
nand U10075 (N_10075,N_1010,N_5549);
nor U10076 (N_10076,N_2837,N_2956);
nor U10077 (N_10077,N_1822,N_5238);
xnor U10078 (N_10078,N_5171,N_5735);
xor U10079 (N_10079,N_3627,N_232);
and U10080 (N_10080,N_5458,N_1300);
and U10081 (N_10081,N_209,N_5189);
and U10082 (N_10082,N_3415,N_3562);
nand U10083 (N_10083,N_3465,N_458);
nand U10084 (N_10084,N_1563,N_1145);
nor U10085 (N_10085,N_1953,N_2439);
nor U10086 (N_10086,N_3777,N_3030);
or U10087 (N_10087,N_5511,N_4483);
and U10088 (N_10088,N_1920,N_547);
nor U10089 (N_10089,N_3427,N_1140);
nand U10090 (N_10090,N_1385,N_654);
xnor U10091 (N_10091,N_1459,N_4292);
xor U10092 (N_10092,N_5859,N_5171);
nand U10093 (N_10093,N_4292,N_2393);
nor U10094 (N_10094,N_4216,N_4751);
or U10095 (N_10095,N_4515,N_5621);
or U10096 (N_10096,N_1372,N_2758);
nor U10097 (N_10097,N_2319,N_3414);
nand U10098 (N_10098,N_1768,N_5657);
xnor U10099 (N_10099,N_5886,N_375);
nor U10100 (N_10100,N_3981,N_2366);
nand U10101 (N_10101,N_3022,N_2133);
or U10102 (N_10102,N_5154,N_1928);
or U10103 (N_10103,N_1064,N_3662);
nor U10104 (N_10104,N_3034,N_3387);
and U10105 (N_10105,N_5835,N_5102);
nand U10106 (N_10106,N_1696,N_3244);
xor U10107 (N_10107,N_851,N_522);
and U10108 (N_10108,N_4804,N_2353);
and U10109 (N_10109,N_2035,N_1172);
nand U10110 (N_10110,N_4345,N_870);
xor U10111 (N_10111,N_3714,N_202);
nor U10112 (N_10112,N_3823,N_4381);
or U10113 (N_10113,N_2382,N_3413);
nand U10114 (N_10114,N_3869,N_3040);
or U10115 (N_10115,N_3385,N_3433);
and U10116 (N_10116,N_2330,N_3627);
or U10117 (N_10117,N_3414,N_1108);
nor U10118 (N_10118,N_954,N_1732);
nand U10119 (N_10119,N_677,N_5246);
nor U10120 (N_10120,N_4331,N_5864);
nand U10121 (N_10121,N_772,N_2129);
or U10122 (N_10122,N_1918,N_2246);
and U10123 (N_10123,N_4181,N_1309);
xor U10124 (N_10124,N_5624,N_1334);
xor U10125 (N_10125,N_4823,N_45);
nand U10126 (N_10126,N_2935,N_1618);
and U10127 (N_10127,N_5139,N_1424);
nor U10128 (N_10128,N_4658,N_5899);
and U10129 (N_10129,N_4220,N_176);
and U10130 (N_10130,N_2780,N_2698);
or U10131 (N_10131,N_5229,N_2619);
nand U10132 (N_10132,N_4048,N_3589);
and U10133 (N_10133,N_5068,N_3084);
nand U10134 (N_10134,N_2044,N_1968);
and U10135 (N_10135,N_1824,N_1435);
nor U10136 (N_10136,N_3778,N_3877);
nand U10137 (N_10137,N_3892,N_534);
or U10138 (N_10138,N_3824,N_1035);
nand U10139 (N_10139,N_4758,N_827);
or U10140 (N_10140,N_4499,N_3163);
or U10141 (N_10141,N_200,N_656);
nand U10142 (N_10142,N_1164,N_3424);
nand U10143 (N_10143,N_5843,N_3847);
nand U10144 (N_10144,N_4934,N_1056);
xnor U10145 (N_10145,N_4324,N_3869);
xnor U10146 (N_10146,N_3302,N_817);
and U10147 (N_10147,N_789,N_3980);
nor U10148 (N_10148,N_2546,N_2848);
nor U10149 (N_10149,N_2921,N_4578);
nand U10150 (N_10150,N_1901,N_2535);
and U10151 (N_10151,N_5799,N_1647);
xor U10152 (N_10152,N_2530,N_4945);
nor U10153 (N_10153,N_830,N_5911);
and U10154 (N_10154,N_2358,N_4967);
nand U10155 (N_10155,N_5517,N_224);
xor U10156 (N_10156,N_4442,N_3888);
nand U10157 (N_10157,N_3040,N_3961);
nand U10158 (N_10158,N_56,N_2639);
and U10159 (N_10159,N_3033,N_4284);
or U10160 (N_10160,N_4547,N_2955);
and U10161 (N_10161,N_5650,N_2295);
and U10162 (N_10162,N_1114,N_3427);
or U10163 (N_10163,N_4970,N_2150);
or U10164 (N_10164,N_11,N_4455);
xor U10165 (N_10165,N_1600,N_3753);
and U10166 (N_10166,N_277,N_5374);
or U10167 (N_10167,N_129,N_548);
and U10168 (N_10168,N_165,N_1117);
nand U10169 (N_10169,N_5075,N_4571);
or U10170 (N_10170,N_5478,N_3952);
nand U10171 (N_10171,N_2098,N_1356);
nand U10172 (N_10172,N_4884,N_4943);
nand U10173 (N_10173,N_4847,N_418);
or U10174 (N_10174,N_2924,N_4680);
or U10175 (N_10175,N_5018,N_4991);
and U10176 (N_10176,N_349,N_5207);
xnor U10177 (N_10177,N_1263,N_3004);
xor U10178 (N_10178,N_32,N_2960);
nand U10179 (N_10179,N_713,N_1511);
xnor U10180 (N_10180,N_5407,N_3142);
nand U10181 (N_10181,N_4001,N_1734);
xnor U10182 (N_10182,N_1769,N_405);
nand U10183 (N_10183,N_4734,N_4119);
xnor U10184 (N_10184,N_3784,N_1612);
and U10185 (N_10185,N_1367,N_839);
or U10186 (N_10186,N_2822,N_2340);
nor U10187 (N_10187,N_2089,N_4506);
nand U10188 (N_10188,N_125,N_4720);
nand U10189 (N_10189,N_3089,N_77);
nor U10190 (N_10190,N_1041,N_986);
and U10191 (N_10191,N_5625,N_1383);
or U10192 (N_10192,N_770,N_5378);
xor U10193 (N_10193,N_1977,N_3273);
nor U10194 (N_10194,N_1506,N_5942);
nand U10195 (N_10195,N_5532,N_3923);
and U10196 (N_10196,N_2444,N_279);
nor U10197 (N_10197,N_2319,N_3257);
nand U10198 (N_10198,N_1795,N_3228);
or U10199 (N_10199,N_3906,N_2575);
nor U10200 (N_10200,N_2442,N_2330);
and U10201 (N_10201,N_379,N_2237);
xnor U10202 (N_10202,N_1136,N_1833);
xor U10203 (N_10203,N_4328,N_2381);
nand U10204 (N_10204,N_2847,N_1956);
nand U10205 (N_10205,N_281,N_809);
xnor U10206 (N_10206,N_3765,N_5056);
and U10207 (N_10207,N_5730,N_5707);
or U10208 (N_10208,N_5947,N_1161);
xor U10209 (N_10209,N_2201,N_5131);
and U10210 (N_10210,N_1397,N_2038);
and U10211 (N_10211,N_2571,N_13);
and U10212 (N_10212,N_2314,N_4556);
nand U10213 (N_10213,N_1751,N_3349);
and U10214 (N_10214,N_2237,N_4595);
xor U10215 (N_10215,N_5705,N_1273);
xor U10216 (N_10216,N_772,N_4430);
nand U10217 (N_10217,N_2650,N_1822);
or U10218 (N_10218,N_689,N_914);
nand U10219 (N_10219,N_2492,N_5673);
or U10220 (N_10220,N_5797,N_1851);
and U10221 (N_10221,N_2177,N_160);
nor U10222 (N_10222,N_764,N_2746);
or U10223 (N_10223,N_982,N_560);
and U10224 (N_10224,N_270,N_5899);
and U10225 (N_10225,N_5339,N_3917);
nor U10226 (N_10226,N_5250,N_2947);
nand U10227 (N_10227,N_1760,N_1586);
or U10228 (N_10228,N_3621,N_2092);
and U10229 (N_10229,N_1422,N_4061);
or U10230 (N_10230,N_11,N_3544);
nor U10231 (N_10231,N_5674,N_4912);
xor U10232 (N_10232,N_5897,N_3824);
xnor U10233 (N_10233,N_1003,N_4148);
nor U10234 (N_10234,N_911,N_2171);
or U10235 (N_10235,N_3470,N_5523);
xnor U10236 (N_10236,N_2377,N_890);
nor U10237 (N_10237,N_1929,N_5019);
and U10238 (N_10238,N_4081,N_5267);
nand U10239 (N_10239,N_5886,N_388);
nor U10240 (N_10240,N_3228,N_3974);
xor U10241 (N_10241,N_3289,N_1384);
nand U10242 (N_10242,N_2174,N_2655);
nand U10243 (N_10243,N_2496,N_4915);
nor U10244 (N_10244,N_5065,N_3143);
nand U10245 (N_10245,N_2423,N_2843);
and U10246 (N_10246,N_970,N_4352);
nand U10247 (N_10247,N_3341,N_5672);
or U10248 (N_10248,N_2517,N_5629);
or U10249 (N_10249,N_394,N_634);
nand U10250 (N_10250,N_3700,N_5313);
and U10251 (N_10251,N_3466,N_1192);
and U10252 (N_10252,N_1251,N_2370);
or U10253 (N_10253,N_3199,N_4110);
or U10254 (N_10254,N_2691,N_5731);
and U10255 (N_10255,N_3590,N_2188);
xor U10256 (N_10256,N_5212,N_4255);
and U10257 (N_10257,N_1302,N_3149);
and U10258 (N_10258,N_5263,N_5282);
or U10259 (N_10259,N_5773,N_4471);
or U10260 (N_10260,N_1878,N_2876);
nor U10261 (N_10261,N_1245,N_368);
nand U10262 (N_10262,N_5156,N_2141);
nor U10263 (N_10263,N_2831,N_5549);
or U10264 (N_10264,N_4906,N_1348);
or U10265 (N_10265,N_5972,N_5425);
nor U10266 (N_10266,N_3562,N_4773);
xor U10267 (N_10267,N_206,N_1916);
and U10268 (N_10268,N_3287,N_171);
xnor U10269 (N_10269,N_5663,N_5791);
or U10270 (N_10270,N_2757,N_1263);
nor U10271 (N_10271,N_2470,N_5511);
nand U10272 (N_10272,N_339,N_3659);
or U10273 (N_10273,N_4536,N_458);
and U10274 (N_10274,N_3931,N_1333);
nor U10275 (N_10275,N_527,N_1259);
or U10276 (N_10276,N_3543,N_1385);
or U10277 (N_10277,N_3423,N_2225);
xor U10278 (N_10278,N_1401,N_3716);
nor U10279 (N_10279,N_5786,N_3876);
nor U10280 (N_10280,N_5734,N_707);
xor U10281 (N_10281,N_146,N_1582);
nand U10282 (N_10282,N_311,N_4871);
nand U10283 (N_10283,N_2952,N_1015);
or U10284 (N_10284,N_3033,N_253);
nand U10285 (N_10285,N_2513,N_2379);
xnor U10286 (N_10286,N_2828,N_4215);
xnor U10287 (N_10287,N_12,N_659);
and U10288 (N_10288,N_328,N_3883);
and U10289 (N_10289,N_3797,N_3437);
xnor U10290 (N_10290,N_1466,N_2653);
or U10291 (N_10291,N_2970,N_2054);
nor U10292 (N_10292,N_2693,N_2118);
nand U10293 (N_10293,N_4348,N_4140);
xnor U10294 (N_10294,N_4370,N_2775);
or U10295 (N_10295,N_3194,N_4238);
nor U10296 (N_10296,N_3984,N_2397);
and U10297 (N_10297,N_639,N_3456);
nand U10298 (N_10298,N_3215,N_3981);
and U10299 (N_10299,N_2855,N_1899);
nor U10300 (N_10300,N_3954,N_2543);
nand U10301 (N_10301,N_3149,N_1866);
and U10302 (N_10302,N_3838,N_903);
xnor U10303 (N_10303,N_4473,N_4004);
nor U10304 (N_10304,N_3381,N_4593);
nand U10305 (N_10305,N_5408,N_3226);
nand U10306 (N_10306,N_2725,N_1336);
or U10307 (N_10307,N_1827,N_781);
nor U10308 (N_10308,N_1007,N_1473);
xor U10309 (N_10309,N_443,N_1481);
xor U10310 (N_10310,N_2269,N_770);
and U10311 (N_10311,N_5089,N_5594);
nor U10312 (N_10312,N_3291,N_3190);
nand U10313 (N_10313,N_3173,N_3316);
nand U10314 (N_10314,N_2840,N_1106);
xor U10315 (N_10315,N_1700,N_1624);
nand U10316 (N_10316,N_3601,N_122);
nand U10317 (N_10317,N_2420,N_4718);
and U10318 (N_10318,N_848,N_3759);
xor U10319 (N_10319,N_1457,N_1994);
xor U10320 (N_10320,N_3037,N_3430);
nand U10321 (N_10321,N_5794,N_763);
nand U10322 (N_10322,N_3130,N_4747);
or U10323 (N_10323,N_3068,N_4073);
or U10324 (N_10324,N_1891,N_569);
xnor U10325 (N_10325,N_1588,N_3078);
xor U10326 (N_10326,N_4865,N_1951);
or U10327 (N_10327,N_2824,N_1577);
or U10328 (N_10328,N_1899,N_4874);
nor U10329 (N_10329,N_5687,N_4584);
nand U10330 (N_10330,N_5751,N_4441);
nand U10331 (N_10331,N_4350,N_2833);
xnor U10332 (N_10332,N_5168,N_2340);
nor U10333 (N_10333,N_2913,N_3883);
xnor U10334 (N_10334,N_1110,N_1320);
and U10335 (N_10335,N_4317,N_2857);
and U10336 (N_10336,N_437,N_1452);
and U10337 (N_10337,N_2961,N_1885);
nor U10338 (N_10338,N_3954,N_2837);
xnor U10339 (N_10339,N_3915,N_2297);
nand U10340 (N_10340,N_5855,N_2679);
or U10341 (N_10341,N_3312,N_4805);
or U10342 (N_10342,N_5231,N_2365);
nor U10343 (N_10343,N_5508,N_4859);
nand U10344 (N_10344,N_175,N_3035);
xnor U10345 (N_10345,N_5424,N_2025);
and U10346 (N_10346,N_4822,N_5233);
xor U10347 (N_10347,N_5880,N_2882);
and U10348 (N_10348,N_1216,N_4834);
xor U10349 (N_10349,N_5075,N_615);
nand U10350 (N_10350,N_2391,N_4591);
nor U10351 (N_10351,N_2361,N_3842);
nand U10352 (N_10352,N_4628,N_4161);
or U10353 (N_10353,N_1547,N_4656);
and U10354 (N_10354,N_442,N_4928);
nor U10355 (N_10355,N_545,N_2002);
or U10356 (N_10356,N_3487,N_550);
nand U10357 (N_10357,N_3344,N_5965);
and U10358 (N_10358,N_2166,N_4375);
or U10359 (N_10359,N_137,N_278);
xnor U10360 (N_10360,N_5797,N_1713);
or U10361 (N_10361,N_1265,N_3634);
or U10362 (N_10362,N_4104,N_4370);
xor U10363 (N_10363,N_5841,N_1805);
and U10364 (N_10364,N_3413,N_4525);
xnor U10365 (N_10365,N_5507,N_4574);
nand U10366 (N_10366,N_5006,N_2284);
nand U10367 (N_10367,N_2607,N_5526);
xor U10368 (N_10368,N_3679,N_2420);
xor U10369 (N_10369,N_4468,N_3766);
nor U10370 (N_10370,N_1296,N_643);
nor U10371 (N_10371,N_823,N_3208);
nand U10372 (N_10372,N_3035,N_11);
xor U10373 (N_10373,N_4378,N_1939);
or U10374 (N_10374,N_565,N_394);
or U10375 (N_10375,N_3037,N_2298);
or U10376 (N_10376,N_5266,N_1526);
nand U10377 (N_10377,N_5990,N_597);
and U10378 (N_10378,N_819,N_5437);
and U10379 (N_10379,N_2761,N_5794);
nor U10380 (N_10380,N_5213,N_4530);
xor U10381 (N_10381,N_1646,N_4243);
xnor U10382 (N_10382,N_713,N_4211);
nand U10383 (N_10383,N_3401,N_2252);
nor U10384 (N_10384,N_1939,N_1433);
and U10385 (N_10385,N_3558,N_876);
nor U10386 (N_10386,N_1390,N_840);
xnor U10387 (N_10387,N_1064,N_2534);
and U10388 (N_10388,N_4447,N_3711);
xnor U10389 (N_10389,N_4413,N_3316);
or U10390 (N_10390,N_2181,N_1064);
and U10391 (N_10391,N_3894,N_739);
or U10392 (N_10392,N_2701,N_1158);
and U10393 (N_10393,N_2766,N_27);
and U10394 (N_10394,N_1773,N_401);
and U10395 (N_10395,N_534,N_5854);
or U10396 (N_10396,N_125,N_53);
xor U10397 (N_10397,N_905,N_642);
or U10398 (N_10398,N_379,N_5298);
and U10399 (N_10399,N_5805,N_758);
nand U10400 (N_10400,N_1407,N_5341);
nand U10401 (N_10401,N_1853,N_3923);
xor U10402 (N_10402,N_3828,N_5811);
or U10403 (N_10403,N_5659,N_3072);
or U10404 (N_10404,N_471,N_4321);
and U10405 (N_10405,N_1929,N_5635);
nor U10406 (N_10406,N_5779,N_3677);
nand U10407 (N_10407,N_2805,N_2883);
nor U10408 (N_10408,N_2450,N_2350);
nand U10409 (N_10409,N_3128,N_3031);
or U10410 (N_10410,N_1595,N_2303);
nor U10411 (N_10411,N_4005,N_962);
or U10412 (N_10412,N_5566,N_5288);
xnor U10413 (N_10413,N_3833,N_207);
or U10414 (N_10414,N_10,N_1288);
nand U10415 (N_10415,N_305,N_449);
nand U10416 (N_10416,N_5414,N_1468);
xnor U10417 (N_10417,N_5660,N_219);
nand U10418 (N_10418,N_577,N_2055);
xor U10419 (N_10419,N_4997,N_4781);
nand U10420 (N_10420,N_4656,N_2222);
or U10421 (N_10421,N_4797,N_1265);
xor U10422 (N_10422,N_5435,N_5251);
nor U10423 (N_10423,N_3873,N_2289);
or U10424 (N_10424,N_2540,N_5758);
or U10425 (N_10425,N_5361,N_989);
nand U10426 (N_10426,N_3045,N_4201);
nand U10427 (N_10427,N_4133,N_5433);
nor U10428 (N_10428,N_570,N_1099);
xor U10429 (N_10429,N_1281,N_4417);
or U10430 (N_10430,N_4858,N_3017);
xnor U10431 (N_10431,N_4571,N_925);
xor U10432 (N_10432,N_2062,N_4404);
and U10433 (N_10433,N_4497,N_1929);
or U10434 (N_10434,N_4545,N_1780);
xnor U10435 (N_10435,N_2454,N_5138);
nor U10436 (N_10436,N_3,N_3614);
nor U10437 (N_10437,N_4163,N_1756);
nand U10438 (N_10438,N_3602,N_12);
and U10439 (N_10439,N_729,N_3826);
or U10440 (N_10440,N_1206,N_2527);
nand U10441 (N_10441,N_2265,N_1135);
xor U10442 (N_10442,N_2537,N_2149);
or U10443 (N_10443,N_3472,N_3447);
xnor U10444 (N_10444,N_5884,N_2930);
nor U10445 (N_10445,N_2002,N_5901);
xnor U10446 (N_10446,N_2275,N_5991);
nor U10447 (N_10447,N_4340,N_188);
nand U10448 (N_10448,N_4020,N_5056);
nor U10449 (N_10449,N_1395,N_3322);
nor U10450 (N_10450,N_2959,N_5293);
xor U10451 (N_10451,N_4751,N_3092);
xor U10452 (N_10452,N_414,N_3902);
xnor U10453 (N_10453,N_1629,N_2487);
or U10454 (N_10454,N_5328,N_5258);
xor U10455 (N_10455,N_4547,N_4066);
or U10456 (N_10456,N_4171,N_820);
xor U10457 (N_10457,N_3060,N_868);
or U10458 (N_10458,N_4817,N_2745);
xnor U10459 (N_10459,N_1360,N_768);
and U10460 (N_10460,N_3103,N_5105);
nand U10461 (N_10461,N_1082,N_4233);
xnor U10462 (N_10462,N_3105,N_4951);
nor U10463 (N_10463,N_1625,N_3733);
nand U10464 (N_10464,N_2045,N_5644);
and U10465 (N_10465,N_4581,N_2050);
nand U10466 (N_10466,N_1440,N_1132);
nand U10467 (N_10467,N_5533,N_4746);
xor U10468 (N_10468,N_911,N_5271);
or U10469 (N_10469,N_423,N_2943);
or U10470 (N_10470,N_2904,N_5335);
nor U10471 (N_10471,N_3475,N_2315);
and U10472 (N_10472,N_2516,N_1945);
xnor U10473 (N_10473,N_4742,N_5940);
or U10474 (N_10474,N_91,N_4803);
nand U10475 (N_10475,N_1890,N_1070);
and U10476 (N_10476,N_5970,N_3741);
xnor U10477 (N_10477,N_3850,N_1535);
nor U10478 (N_10478,N_1166,N_3853);
nor U10479 (N_10479,N_4986,N_5228);
nor U10480 (N_10480,N_3239,N_887);
nand U10481 (N_10481,N_134,N_2301);
or U10482 (N_10482,N_4296,N_1249);
and U10483 (N_10483,N_1629,N_538);
xor U10484 (N_10484,N_5347,N_335);
nor U10485 (N_10485,N_3910,N_3397);
xor U10486 (N_10486,N_4181,N_5774);
xor U10487 (N_10487,N_1922,N_2757);
nand U10488 (N_10488,N_2401,N_3164);
xor U10489 (N_10489,N_4759,N_2782);
nor U10490 (N_10490,N_4309,N_3216);
xor U10491 (N_10491,N_3288,N_5031);
xor U10492 (N_10492,N_25,N_4641);
nand U10493 (N_10493,N_2074,N_1464);
xor U10494 (N_10494,N_1449,N_3233);
nor U10495 (N_10495,N_4450,N_4907);
or U10496 (N_10496,N_1668,N_2276);
nand U10497 (N_10497,N_3725,N_2814);
nor U10498 (N_10498,N_2474,N_313);
and U10499 (N_10499,N_1689,N_2583);
nor U10500 (N_10500,N_630,N_2488);
nand U10501 (N_10501,N_305,N_2608);
nand U10502 (N_10502,N_1356,N_4932);
and U10503 (N_10503,N_3293,N_3931);
nor U10504 (N_10504,N_2489,N_3912);
xor U10505 (N_10505,N_187,N_2982);
or U10506 (N_10506,N_96,N_3491);
or U10507 (N_10507,N_22,N_4547);
and U10508 (N_10508,N_5303,N_134);
xor U10509 (N_10509,N_583,N_2252);
nor U10510 (N_10510,N_3920,N_3454);
or U10511 (N_10511,N_1079,N_3204);
xor U10512 (N_10512,N_4254,N_2206);
or U10513 (N_10513,N_1942,N_2766);
nand U10514 (N_10514,N_1289,N_3591);
xor U10515 (N_10515,N_459,N_4207);
or U10516 (N_10516,N_5662,N_3113);
or U10517 (N_10517,N_549,N_5373);
nand U10518 (N_10518,N_5494,N_1963);
nor U10519 (N_10519,N_5636,N_4553);
xnor U10520 (N_10520,N_4417,N_3517);
nand U10521 (N_10521,N_2298,N_3699);
nor U10522 (N_10522,N_5202,N_1260);
xnor U10523 (N_10523,N_373,N_4195);
nand U10524 (N_10524,N_3909,N_3718);
xor U10525 (N_10525,N_3040,N_5963);
or U10526 (N_10526,N_3195,N_5827);
nand U10527 (N_10527,N_2930,N_5908);
xor U10528 (N_10528,N_3150,N_2181);
nor U10529 (N_10529,N_620,N_841);
nor U10530 (N_10530,N_4375,N_4732);
xor U10531 (N_10531,N_4005,N_1324);
nand U10532 (N_10532,N_1876,N_4098);
nand U10533 (N_10533,N_4009,N_819);
or U10534 (N_10534,N_751,N_4096);
nor U10535 (N_10535,N_5859,N_950);
or U10536 (N_10536,N_4129,N_2276);
nor U10537 (N_10537,N_3117,N_2231);
and U10538 (N_10538,N_5842,N_2752);
nand U10539 (N_10539,N_602,N_1200);
and U10540 (N_10540,N_5699,N_4707);
nor U10541 (N_10541,N_2283,N_4676);
nand U10542 (N_10542,N_2787,N_3715);
or U10543 (N_10543,N_1827,N_5317);
nor U10544 (N_10544,N_1536,N_1876);
nor U10545 (N_10545,N_3290,N_756);
or U10546 (N_10546,N_2836,N_3964);
and U10547 (N_10547,N_2503,N_2982);
xor U10548 (N_10548,N_4589,N_2646);
or U10549 (N_10549,N_4723,N_158);
and U10550 (N_10550,N_3506,N_4502);
nand U10551 (N_10551,N_672,N_189);
nor U10552 (N_10552,N_5653,N_3801);
and U10553 (N_10553,N_3458,N_937);
and U10554 (N_10554,N_2517,N_5508);
or U10555 (N_10555,N_2808,N_3959);
xnor U10556 (N_10556,N_4889,N_5977);
xnor U10557 (N_10557,N_5347,N_3623);
nand U10558 (N_10558,N_1109,N_5063);
and U10559 (N_10559,N_5960,N_5992);
xor U10560 (N_10560,N_555,N_5208);
nor U10561 (N_10561,N_5150,N_633);
nand U10562 (N_10562,N_1493,N_1785);
nand U10563 (N_10563,N_1844,N_65);
and U10564 (N_10564,N_1715,N_788);
and U10565 (N_10565,N_5673,N_893);
xnor U10566 (N_10566,N_5651,N_2752);
nor U10567 (N_10567,N_2594,N_4066);
and U10568 (N_10568,N_3420,N_569);
and U10569 (N_10569,N_3777,N_835);
nand U10570 (N_10570,N_2363,N_5359);
nor U10571 (N_10571,N_2334,N_2138);
nor U10572 (N_10572,N_3493,N_4076);
and U10573 (N_10573,N_1388,N_3670);
nand U10574 (N_10574,N_2532,N_2498);
nor U10575 (N_10575,N_1300,N_4376);
xor U10576 (N_10576,N_3895,N_3467);
and U10577 (N_10577,N_2451,N_3407);
nor U10578 (N_10578,N_3101,N_5446);
nand U10579 (N_10579,N_292,N_1439);
xor U10580 (N_10580,N_721,N_748);
nor U10581 (N_10581,N_1184,N_5737);
xnor U10582 (N_10582,N_4474,N_1242);
or U10583 (N_10583,N_5269,N_4722);
nor U10584 (N_10584,N_1009,N_1112);
nor U10585 (N_10585,N_4991,N_1197);
xor U10586 (N_10586,N_1715,N_2949);
and U10587 (N_10587,N_2242,N_1366);
or U10588 (N_10588,N_3810,N_1295);
nand U10589 (N_10589,N_1951,N_1786);
nand U10590 (N_10590,N_4320,N_4492);
nor U10591 (N_10591,N_1883,N_2236);
or U10592 (N_10592,N_1109,N_2487);
nor U10593 (N_10593,N_2929,N_1080);
nor U10594 (N_10594,N_5543,N_2220);
and U10595 (N_10595,N_5675,N_592);
and U10596 (N_10596,N_4159,N_4215);
nand U10597 (N_10597,N_3458,N_2299);
nand U10598 (N_10598,N_5157,N_5139);
and U10599 (N_10599,N_2761,N_5829);
xor U10600 (N_10600,N_2856,N_4394);
nand U10601 (N_10601,N_725,N_4298);
nand U10602 (N_10602,N_2328,N_2700);
or U10603 (N_10603,N_4155,N_276);
or U10604 (N_10604,N_582,N_1070);
nand U10605 (N_10605,N_2151,N_4853);
xnor U10606 (N_10606,N_2665,N_4817);
nor U10607 (N_10607,N_2192,N_118);
xor U10608 (N_10608,N_160,N_4397);
xor U10609 (N_10609,N_2914,N_2221);
and U10610 (N_10610,N_701,N_1445);
and U10611 (N_10611,N_4611,N_4174);
and U10612 (N_10612,N_1330,N_2432);
xnor U10613 (N_10613,N_2885,N_4154);
and U10614 (N_10614,N_5783,N_2899);
xnor U10615 (N_10615,N_263,N_2201);
or U10616 (N_10616,N_4852,N_5759);
and U10617 (N_10617,N_1973,N_4078);
xnor U10618 (N_10618,N_760,N_5821);
xor U10619 (N_10619,N_1488,N_1317);
or U10620 (N_10620,N_61,N_75);
xor U10621 (N_10621,N_2927,N_4799);
or U10622 (N_10622,N_1410,N_1838);
xnor U10623 (N_10623,N_3236,N_5025);
xnor U10624 (N_10624,N_4530,N_2783);
or U10625 (N_10625,N_344,N_5068);
and U10626 (N_10626,N_2377,N_2029);
xnor U10627 (N_10627,N_888,N_5111);
and U10628 (N_10628,N_1912,N_5430);
and U10629 (N_10629,N_1051,N_1317);
nand U10630 (N_10630,N_5420,N_1164);
xnor U10631 (N_10631,N_3304,N_3671);
xnor U10632 (N_10632,N_4352,N_5639);
or U10633 (N_10633,N_3511,N_1753);
xnor U10634 (N_10634,N_421,N_4165);
nor U10635 (N_10635,N_5924,N_1307);
nand U10636 (N_10636,N_859,N_343);
and U10637 (N_10637,N_353,N_2182);
or U10638 (N_10638,N_57,N_4260);
nor U10639 (N_10639,N_667,N_3841);
and U10640 (N_10640,N_3325,N_87);
or U10641 (N_10641,N_29,N_1726);
nand U10642 (N_10642,N_1855,N_5528);
or U10643 (N_10643,N_5815,N_1131);
nand U10644 (N_10644,N_2655,N_4748);
or U10645 (N_10645,N_3784,N_5560);
nand U10646 (N_10646,N_5347,N_202);
nand U10647 (N_10647,N_3225,N_3901);
nand U10648 (N_10648,N_5928,N_2330);
or U10649 (N_10649,N_5645,N_501);
xnor U10650 (N_10650,N_5365,N_2704);
and U10651 (N_10651,N_5985,N_1045);
and U10652 (N_10652,N_3429,N_304);
and U10653 (N_10653,N_2502,N_5893);
nand U10654 (N_10654,N_4250,N_2319);
nand U10655 (N_10655,N_4574,N_1038);
nor U10656 (N_10656,N_2160,N_5086);
nand U10657 (N_10657,N_4541,N_4460);
or U10658 (N_10658,N_1864,N_3182);
xor U10659 (N_10659,N_316,N_3213);
or U10660 (N_10660,N_2355,N_5666);
or U10661 (N_10661,N_3399,N_3939);
nand U10662 (N_10662,N_3079,N_2125);
and U10663 (N_10663,N_2664,N_5419);
nand U10664 (N_10664,N_5199,N_946);
nand U10665 (N_10665,N_173,N_3014);
nand U10666 (N_10666,N_1975,N_4909);
xnor U10667 (N_10667,N_1409,N_2842);
or U10668 (N_10668,N_5836,N_5564);
nand U10669 (N_10669,N_1154,N_4786);
xor U10670 (N_10670,N_1838,N_3339);
xor U10671 (N_10671,N_5684,N_5834);
or U10672 (N_10672,N_5921,N_2437);
and U10673 (N_10673,N_1954,N_2201);
nor U10674 (N_10674,N_1234,N_2495);
xor U10675 (N_10675,N_2622,N_5943);
nor U10676 (N_10676,N_3444,N_5903);
nor U10677 (N_10677,N_1042,N_5396);
nand U10678 (N_10678,N_3270,N_5122);
nor U10679 (N_10679,N_734,N_545);
and U10680 (N_10680,N_1312,N_498);
and U10681 (N_10681,N_5318,N_4915);
or U10682 (N_10682,N_2407,N_3083);
xnor U10683 (N_10683,N_3498,N_3549);
nor U10684 (N_10684,N_826,N_1054);
xnor U10685 (N_10685,N_5261,N_3653);
nor U10686 (N_10686,N_1131,N_1924);
nor U10687 (N_10687,N_4750,N_1578);
nand U10688 (N_10688,N_5070,N_5973);
or U10689 (N_10689,N_4450,N_4999);
nor U10690 (N_10690,N_4020,N_2026);
nand U10691 (N_10691,N_686,N_3069);
nand U10692 (N_10692,N_2813,N_404);
xnor U10693 (N_10693,N_3919,N_2546);
or U10694 (N_10694,N_4022,N_2113);
nand U10695 (N_10695,N_964,N_1014);
nor U10696 (N_10696,N_4412,N_2207);
or U10697 (N_10697,N_2772,N_3912);
or U10698 (N_10698,N_5921,N_3027);
xnor U10699 (N_10699,N_2786,N_5713);
xor U10700 (N_10700,N_5676,N_24);
or U10701 (N_10701,N_1757,N_5238);
and U10702 (N_10702,N_4699,N_4680);
or U10703 (N_10703,N_948,N_747);
nand U10704 (N_10704,N_4066,N_1396);
nor U10705 (N_10705,N_5461,N_50);
xnor U10706 (N_10706,N_3985,N_1364);
nand U10707 (N_10707,N_3656,N_2296);
nand U10708 (N_10708,N_5271,N_1480);
xor U10709 (N_10709,N_3151,N_5386);
nand U10710 (N_10710,N_4783,N_2012);
nor U10711 (N_10711,N_2858,N_5915);
nor U10712 (N_10712,N_702,N_3412);
and U10713 (N_10713,N_3314,N_1859);
xnor U10714 (N_10714,N_5173,N_612);
nor U10715 (N_10715,N_3106,N_4525);
nand U10716 (N_10716,N_339,N_1470);
nor U10717 (N_10717,N_2085,N_5407);
xnor U10718 (N_10718,N_230,N_1583);
nand U10719 (N_10719,N_3739,N_2999);
and U10720 (N_10720,N_4577,N_474);
nor U10721 (N_10721,N_1250,N_2284);
nor U10722 (N_10722,N_3097,N_10);
nor U10723 (N_10723,N_4027,N_2834);
or U10724 (N_10724,N_5675,N_4552);
and U10725 (N_10725,N_4102,N_1602);
nand U10726 (N_10726,N_4457,N_1334);
xnor U10727 (N_10727,N_3797,N_1734);
xnor U10728 (N_10728,N_2139,N_1531);
nor U10729 (N_10729,N_925,N_4291);
nand U10730 (N_10730,N_5609,N_116);
nor U10731 (N_10731,N_5118,N_3199);
xnor U10732 (N_10732,N_770,N_5971);
xor U10733 (N_10733,N_4435,N_2871);
xor U10734 (N_10734,N_1051,N_756);
nand U10735 (N_10735,N_757,N_1194);
and U10736 (N_10736,N_3387,N_3078);
or U10737 (N_10737,N_872,N_150);
nor U10738 (N_10738,N_3706,N_2691);
nor U10739 (N_10739,N_1455,N_344);
nor U10740 (N_10740,N_3704,N_532);
nand U10741 (N_10741,N_1288,N_5774);
nor U10742 (N_10742,N_5406,N_3905);
xor U10743 (N_10743,N_2261,N_5251);
xnor U10744 (N_10744,N_870,N_2638);
xnor U10745 (N_10745,N_1330,N_5655);
or U10746 (N_10746,N_538,N_4992);
nor U10747 (N_10747,N_3876,N_3654);
and U10748 (N_10748,N_1796,N_1698);
or U10749 (N_10749,N_5946,N_5004);
or U10750 (N_10750,N_1448,N_1925);
nor U10751 (N_10751,N_1165,N_4341);
xor U10752 (N_10752,N_282,N_4857);
xnor U10753 (N_10753,N_1287,N_5277);
and U10754 (N_10754,N_2093,N_814);
and U10755 (N_10755,N_4858,N_5745);
xnor U10756 (N_10756,N_3693,N_2293);
and U10757 (N_10757,N_1025,N_1407);
xnor U10758 (N_10758,N_2354,N_1343);
nor U10759 (N_10759,N_1751,N_990);
xor U10760 (N_10760,N_2579,N_397);
nand U10761 (N_10761,N_3514,N_5785);
xnor U10762 (N_10762,N_4933,N_2692);
and U10763 (N_10763,N_5925,N_4689);
nor U10764 (N_10764,N_1831,N_3526);
xnor U10765 (N_10765,N_2564,N_5379);
xnor U10766 (N_10766,N_2691,N_5244);
or U10767 (N_10767,N_4683,N_5763);
or U10768 (N_10768,N_3756,N_4504);
nor U10769 (N_10769,N_5856,N_3724);
xnor U10770 (N_10770,N_5495,N_5909);
and U10771 (N_10771,N_3496,N_2535);
nor U10772 (N_10772,N_3507,N_4558);
nand U10773 (N_10773,N_1322,N_674);
nor U10774 (N_10774,N_5583,N_362);
xnor U10775 (N_10775,N_3673,N_969);
or U10776 (N_10776,N_654,N_3844);
nand U10777 (N_10777,N_961,N_3220);
or U10778 (N_10778,N_5081,N_2168);
nor U10779 (N_10779,N_2935,N_973);
nand U10780 (N_10780,N_4951,N_863);
and U10781 (N_10781,N_4996,N_877);
xor U10782 (N_10782,N_4207,N_4373);
and U10783 (N_10783,N_1930,N_183);
nor U10784 (N_10784,N_5068,N_348);
or U10785 (N_10785,N_2577,N_2018);
and U10786 (N_10786,N_5729,N_408);
and U10787 (N_10787,N_5160,N_3000);
and U10788 (N_10788,N_5707,N_581);
nor U10789 (N_10789,N_3012,N_4555);
nand U10790 (N_10790,N_4614,N_2777);
and U10791 (N_10791,N_3038,N_1);
nor U10792 (N_10792,N_1523,N_5430);
or U10793 (N_10793,N_1058,N_524);
and U10794 (N_10794,N_633,N_1277);
xor U10795 (N_10795,N_2665,N_4048);
nor U10796 (N_10796,N_3203,N_113);
or U10797 (N_10797,N_3258,N_910);
and U10798 (N_10798,N_1924,N_3471);
nand U10799 (N_10799,N_1902,N_3054);
or U10800 (N_10800,N_661,N_5770);
and U10801 (N_10801,N_3176,N_4389);
xnor U10802 (N_10802,N_1178,N_1937);
xor U10803 (N_10803,N_1338,N_2147);
or U10804 (N_10804,N_459,N_1767);
or U10805 (N_10805,N_5855,N_1943);
or U10806 (N_10806,N_2052,N_1172);
or U10807 (N_10807,N_5467,N_3257);
xnor U10808 (N_10808,N_5080,N_3987);
or U10809 (N_10809,N_749,N_2402);
nand U10810 (N_10810,N_2252,N_5684);
or U10811 (N_10811,N_1166,N_3252);
nor U10812 (N_10812,N_4049,N_2477);
and U10813 (N_10813,N_2897,N_5349);
and U10814 (N_10814,N_4544,N_2391);
xor U10815 (N_10815,N_1409,N_2645);
and U10816 (N_10816,N_3065,N_513);
and U10817 (N_10817,N_599,N_2097);
or U10818 (N_10818,N_4277,N_1596);
xor U10819 (N_10819,N_463,N_1995);
xor U10820 (N_10820,N_1685,N_4400);
or U10821 (N_10821,N_1187,N_3730);
nand U10822 (N_10822,N_2639,N_3576);
nor U10823 (N_10823,N_4176,N_1170);
or U10824 (N_10824,N_4167,N_3637);
xor U10825 (N_10825,N_5255,N_5224);
and U10826 (N_10826,N_3122,N_4038);
nor U10827 (N_10827,N_5289,N_2110);
nor U10828 (N_10828,N_5871,N_5914);
or U10829 (N_10829,N_1201,N_287);
nor U10830 (N_10830,N_435,N_1899);
and U10831 (N_10831,N_3857,N_5134);
or U10832 (N_10832,N_2368,N_4402);
nand U10833 (N_10833,N_2961,N_5067);
or U10834 (N_10834,N_1286,N_5941);
nand U10835 (N_10835,N_2146,N_5641);
and U10836 (N_10836,N_616,N_2847);
or U10837 (N_10837,N_1047,N_5574);
xor U10838 (N_10838,N_4265,N_3248);
nor U10839 (N_10839,N_4210,N_4628);
nand U10840 (N_10840,N_2553,N_4007);
nor U10841 (N_10841,N_4443,N_5902);
and U10842 (N_10842,N_1011,N_4874);
or U10843 (N_10843,N_4037,N_3347);
or U10844 (N_10844,N_5957,N_1579);
nor U10845 (N_10845,N_4948,N_4677);
nand U10846 (N_10846,N_1012,N_2111);
nor U10847 (N_10847,N_1817,N_4555);
xor U10848 (N_10848,N_2941,N_4120);
xor U10849 (N_10849,N_3901,N_4214);
and U10850 (N_10850,N_3178,N_4729);
nand U10851 (N_10851,N_447,N_1218);
or U10852 (N_10852,N_3398,N_4779);
xnor U10853 (N_10853,N_4936,N_4864);
xor U10854 (N_10854,N_2198,N_3142);
xor U10855 (N_10855,N_5536,N_4744);
or U10856 (N_10856,N_5315,N_4826);
nand U10857 (N_10857,N_2257,N_5545);
nor U10858 (N_10858,N_3375,N_5028);
xor U10859 (N_10859,N_5284,N_4548);
nor U10860 (N_10860,N_1483,N_5001);
or U10861 (N_10861,N_3110,N_492);
and U10862 (N_10862,N_2786,N_2088);
and U10863 (N_10863,N_2856,N_125);
or U10864 (N_10864,N_1312,N_3568);
nand U10865 (N_10865,N_1130,N_5250);
or U10866 (N_10866,N_4521,N_5985);
and U10867 (N_10867,N_5455,N_1251);
nand U10868 (N_10868,N_2063,N_434);
and U10869 (N_10869,N_5798,N_1502);
xor U10870 (N_10870,N_562,N_5618);
and U10871 (N_10871,N_1635,N_1185);
and U10872 (N_10872,N_2932,N_5539);
or U10873 (N_10873,N_5418,N_5434);
nand U10874 (N_10874,N_4702,N_1223);
xor U10875 (N_10875,N_3654,N_1336);
nor U10876 (N_10876,N_4763,N_3544);
and U10877 (N_10877,N_4545,N_3915);
nand U10878 (N_10878,N_5678,N_4821);
xnor U10879 (N_10879,N_3931,N_3524);
and U10880 (N_10880,N_2150,N_2716);
xnor U10881 (N_10881,N_400,N_3517);
or U10882 (N_10882,N_3562,N_2430);
and U10883 (N_10883,N_2112,N_1251);
xnor U10884 (N_10884,N_2771,N_2227);
xnor U10885 (N_10885,N_3023,N_4522);
nand U10886 (N_10886,N_3505,N_2403);
and U10887 (N_10887,N_2164,N_4019);
xnor U10888 (N_10888,N_3664,N_4011);
nand U10889 (N_10889,N_141,N_3993);
and U10890 (N_10890,N_5440,N_2578);
nor U10891 (N_10891,N_3291,N_5267);
xnor U10892 (N_10892,N_5797,N_879);
nand U10893 (N_10893,N_553,N_4003);
and U10894 (N_10894,N_4922,N_2012);
nand U10895 (N_10895,N_4685,N_3790);
nor U10896 (N_10896,N_2739,N_16);
xor U10897 (N_10897,N_1848,N_5733);
xnor U10898 (N_10898,N_5203,N_3897);
or U10899 (N_10899,N_3742,N_599);
or U10900 (N_10900,N_5502,N_3601);
nor U10901 (N_10901,N_2576,N_898);
or U10902 (N_10902,N_3329,N_954);
nor U10903 (N_10903,N_5759,N_1980);
xnor U10904 (N_10904,N_3744,N_5419);
and U10905 (N_10905,N_3950,N_907);
or U10906 (N_10906,N_4419,N_5532);
nor U10907 (N_10907,N_690,N_5884);
and U10908 (N_10908,N_1238,N_3134);
nor U10909 (N_10909,N_2935,N_4687);
xnor U10910 (N_10910,N_718,N_1505);
and U10911 (N_10911,N_2433,N_4791);
xor U10912 (N_10912,N_2234,N_4190);
and U10913 (N_10913,N_2905,N_3468);
or U10914 (N_10914,N_1692,N_5750);
xor U10915 (N_10915,N_5363,N_2947);
xnor U10916 (N_10916,N_3040,N_5235);
xnor U10917 (N_10917,N_2796,N_1266);
xnor U10918 (N_10918,N_1421,N_3920);
xnor U10919 (N_10919,N_2536,N_4143);
xnor U10920 (N_10920,N_845,N_2737);
nor U10921 (N_10921,N_4860,N_363);
nand U10922 (N_10922,N_1929,N_5010);
xor U10923 (N_10923,N_3476,N_3175);
nand U10924 (N_10924,N_1634,N_952);
xnor U10925 (N_10925,N_1797,N_3940);
and U10926 (N_10926,N_4427,N_3421);
nor U10927 (N_10927,N_654,N_190);
nand U10928 (N_10928,N_1611,N_2725);
nand U10929 (N_10929,N_1415,N_2258);
nor U10930 (N_10930,N_2750,N_2729);
xor U10931 (N_10931,N_3898,N_3853);
and U10932 (N_10932,N_5578,N_938);
nand U10933 (N_10933,N_1684,N_1237);
xor U10934 (N_10934,N_3409,N_3368);
and U10935 (N_10935,N_4318,N_1300);
nor U10936 (N_10936,N_2965,N_4528);
nand U10937 (N_10937,N_1279,N_5817);
xor U10938 (N_10938,N_5300,N_3749);
xnor U10939 (N_10939,N_940,N_2427);
nand U10940 (N_10940,N_427,N_3171);
nor U10941 (N_10941,N_545,N_1384);
or U10942 (N_10942,N_2096,N_4027);
nand U10943 (N_10943,N_2992,N_3416);
xor U10944 (N_10944,N_3679,N_305);
nand U10945 (N_10945,N_5396,N_1737);
or U10946 (N_10946,N_5776,N_4316);
or U10947 (N_10947,N_1029,N_4826);
and U10948 (N_10948,N_2334,N_4535);
and U10949 (N_10949,N_3411,N_1085);
and U10950 (N_10950,N_3772,N_3052);
nor U10951 (N_10951,N_3322,N_2158);
and U10952 (N_10952,N_690,N_3176);
nor U10953 (N_10953,N_1696,N_2246);
or U10954 (N_10954,N_4135,N_2157);
nor U10955 (N_10955,N_4749,N_5392);
and U10956 (N_10956,N_5039,N_5744);
nand U10957 (N_10957,N_3916,N_231);
and U10958 (N_10958,N_3318,N_5285);
nand U10959 (N_10959,N_1690,N_5006);
xnor U10960 (N_10960,N_1489,N_787);
nand U10961 (N_10961,N_4392,N_2152);
or U10962 (N_10962,N_1291,N_387);
nor U10963 (N_10963,N_5746,N_2548);
nor U10964 (N_10964,N_1528,N_5291);
nand U10965 (N_10965,N_2403,N_2166);
and U10966 (N_10966,N_1541,N_1682);
xnor U10967 (N_10967,N_3504,N_1273);
nand U10968 (N_10968,N_5475,N_1405);
or U10969 (N_10969,N_113,N_1754);
or U10970 (N_10970,N_1854,N_4522);
nor U10971 (N_10971,N_1433,N_3600);
and U10972 (N_10972,N_326,N_1084);
or U10973 (N_10973,N_2716,N_5314);
xnor U10974 (N_10974,N_711,N_4884);
and U10975 (N_10975,N_2885,N_3853);
or U10976 (N_10976,N_2017,N_3027);
or U10977 (N_10977,N_4788,N_3412);
or U10978 (N_10978,N_1675,N_5025);
xnor U10979 (N_10979,N_3754,N_1351);
nand U10980 (N_10980,N_3642,N_233);
or U10981 (N_10981,N_4022,N_2230);
nor U10982 (N_10982,N_4175,N_249);
or U10983 (N_10983,N_283,N_1635);
xnor U10984 (N_10984,N_4002,N_4411);
or U10985 (N_10985,N_3922,N_293);
nand U10986 (N_10986,N_3816,N_5506);
and U10987 (N_10987,N_1624,N_5287);
nor U10988 (N_10988,N_530,N_487);
nor U10989 (N_10989,N_2625,N_2948);
nand U10990 (N_10990,N_3482,N_1869);
nor U10991 (N_10991,N_5600,N_4516);
nand U10992 (N_10992,N_5387,N_3295);
nand U10993 (N_10993,N_3125,N_890);
nand U10994 (N_10994,N_4896,N_1810);
xor U10995 (N_10995,N_5979,N_4682);
and U10996 (N_10996,N_127,N_992);
and U10997 (N_10997,N_1047,N_2251);
and U10998 (N_10998,N_2434,N_1616);
and U10999 (N_10999,N_2496,N_589);
and U11000 (N_11000,N_1495,N_958);
and U11001 (N_11001,N_4846,N_2658);
and U11002 (N_11002,N_1192,N_5846);
and U11003 (N_11003,N_2032,N_931);
xnor U11004 (N_11004,N_3695,N_3816);
xor U11005 (N_11005,N_4407,N_3675);
nand U11006 (N_11006,N_3697,N_2904);
nor U11007 (N_11007,N_4830,N_741);
nor U11008 (N_11008,N_710,N_3793);
nor U11009 (N_11009,N_2423,N_4018);
nand U11010 (N_11010,N_1164,N_1837);
xnor U11011 (N_11011,N_4825,N_5708);
and U11012 (N_11012,N_2907,N_4774);
nor U11013 (N_11013,N_448,N_4825);
and U11014 (N_11014,N_5481,N_726);
or U11015 (N_11015,N_633,N_757);
and U11016 (N_11016,N_1306,N_5185);
xor U11017 (N_11017,N_960,N_257);
or U11018 (N_11018,N_1798,N_5303);
and U11019 (N_11019,N_823,N_2165);
nand U11020 (N_11020,N_2692,N_2027);
and U11021 (N_11021,N_1365,N_4775);
nand U11022 (N_11022,N_1549,N_2720);
or U11023 (N_11023,N_824,N_5778);
nor U11024 (N_11024,N_5992,N_53);
xnor U11025 (N_11025,N_3513,N_4678);
nor U11026 (N_11026,N_2453,N_605);
nand U11027 (N_11027,N_438,N_2294);
or U11028 (N_11028,N_1137,N_3218);
and U11029 (N_11029,N_159,N_4737);
or U11030 (N_11030,N_4779,N_5622);
nand U11031 (N_11031,N_863,N_2455);
nor U11032 (N_11032,N_3158,N_1675);
or U11033 (N_11033,N_1435,N_4423);
and U11034 (N_11034,N_3281,N_5569);
or U11035 (N_11035,N_5826,N_5285);
nor U11036 (N_11036,N_3047,N_2547);
and U11037 (N_11037,N_5820,N_528);
nor U11038 (N_11038,N_3402,N_2046);
and U11039 (N_11039,N_2634,N_314);
or U11040 (N_11040,N_4477,N_3681);
xnor U11041 (N_11041,N_2906,N_2521);
nor U11042 (N_11042,N_3451,N_5387);
xnor U11043 (N_11043,N_5151,N_2969);
xor U11044 (N_11044,N_2285,N_276);
or U11045 (N_11045,N_235,N_1783);
and U11046 (N_11046,N_4124,N_279);
xor U11047 (N_11047,N_2855,N_1852);
or U11048 (N_11048,N_2076,N_1907);
xor U11049 (N_11049,N_1066,N_3606);
or U11050 (N_11050,N_3368,N_1024);
nor U11051 (N_11051,N_991,N_4807);
and U11052 (N_11052,N_3300,N_914);
and U11053 (N_11053,N_1820,N_5003);
xnor U11054 (N_11054,N_2642,N_2863);
and U11055 (N_11055,N_2468,N_2752);
xor U11056 (N_11056,N_2650,N_4585);
or U11057 (N_11057,N_2047,N_1100);
nand U11058 (N_11058,N_2410,N_2285);
nand U11059 (N_11059,N_5516,N_4011);
nor U11060 (N_11060,N_2491,N_2643);
or U11061 (N_11061,N_4197,N_749);
or U11062 (N_11062,N_1500,N_1600);
and U11063 (N_11063,N_4109,N_1122);
nand U11064 (N_11064,N_1174,N_2660);
xnor U11065 (N_11065,N_4997,N_780);
nand U11066 (N_11066,N_793,N_5078);
nand U11067 (N_11067,N_2929,N_604);
xor U11068 (N_11068,N_3554,N_4649);
nor U11069 (N_11069,N_4360,N_148);
nor U11070 (N_11070,N_232,N_5951);
nor U11071 (N_11071,N_4922,N_5977);
nand U11072 (N_11072,N_1080,N_2805);
or U11073 (N_11073,N_3286,N_3993);
or U11074 (N_11074,N_310,N_3690);
nor U11075 (N_11075,N_2385,N_1433);
nand U11076 (N_11076,N_5457,N_2808);
nor U11077 (N_11077,N_2659,N_3687);
and U11078 (N_11078,N_660,N_3092);
nor U11079 (N_11079,N_1961,N_2453);
and U11080 (N_11080,N_4292,N_2124);
xor U11081 (N_11081,N_4709,N_4077);
or U11082 (N_11082,N_4203,N_1994);
nor U11083 (N_11083,N_508,N_4429);
nor U11084 (N_11084,N_5685,N_4298);
and U11085 (N_11085,N_4519,N_242);
and U11086 (N_11086,N_2229,N_1503);
nand U11087 (N_11087,N_4931,N_1089);
nand U11088 (N_11088,N_3612,N_490);
xnor U11089 (N_11089,N_2164,N_2286);
or U11090 (N_11090,N_135,N_4084);
nand U11091 (N_11091,N_1466,N_406);
nor U11092 (N_11092,N_1826,N_16);
and U11093 (N_11093,N_1016,N_3230);
or U11094 (N_11094,N_677,N_4146);
and U11095 (N_11095,N_5930,N_2822);
or U11096 (N_11096,N_4804,N_1347);
xnor U11097 (N_11097,N_4211,N_1205);
nand U11098 (N_11098,N_1786,N_163);
xor U11099 (N_11099,N_758,N_2844);
or U11100 (N_11100,N_4332,N_1418);
and U11101 (N_11101,N_2052,N_850);
or U11102 (N_11102,N_194,N_1899);
nor U11103 (N_11103,N_5532,N_5620);
nand U11104 (N_11104,N_2678,N_964);
xor U11105 (N_11105,N_1693,N_3521);
and U11106 (N_11106,N_644,N_134);
nor U11107 (N_11107,N_1753,N_5721);
nor U11108 (N_11108,N_5168,N_3275);
nor U11109 (N_11109,N_2656,N_1605);
and U11110 (N_11110,N_2150,N_2893);
or U11111 (N_11111,N_3952,N_1584);
and U11112 (N_11112,N_835,N_2440);
xnor U11113 (N_11113,N_5606,N_368);
xor U11114 (N_11114,N_2782,N_1547);
xor U11115 (N_11115,N_4474,N_2084);
and U11116 (N_11116,N_3956,N_2926);
xor U11117 (N_11117,N_1975,N_3008);
and U11118 (N_11118,N_5306,N_5077);
xnor U11119 (N_11119,N_2569,N_1614);
nor U11120 (N_11120,N_5117,N_3746);
nand U11121 (N_11121,N_2904,N_4429);
nor U11122 (N_11122,N_5864,N_2000);
nand U11123 (N_11123,N_1800,N_3341);
xor U11124 (N_11124,N_5217,N_4827);
or U11125 (N_11125,N_2304,N_4420);
xnor U11126 (N_11126,N_2881,N_2641);
nor U11127 (N_11127,N_3012,N_3470);
and U11128 (N_11128,N_3136,N_638);
xor U11129 (N_11129,N_3717,N_4977);
or U11130 (N_11130,N_3674,N_1697);
and U11131 (N_11131,N_2353,N_1800);
nand U11132 (N_11132,N_2929,N_5691);
or U11133 (N_11133,N_4703,N_3082);
and U11134 (N_11134,N_4803,N_4538);
or U11135 (N_11135,N_3141,N_1157);
nor U11136 (N_11136,N_236,N_2050);
nor U11137 (N_11137,N_2287,N_4140);
or U11138 (N_11138,N_674,N_2083);
nand U11139 (N_11139,N_5237,N_2369);
nand U11140 (N_11140,N_2953,N_398);
nand U11141 (N_11141,N_5097,N_5285);
xnor U11142 (N_11142,N_2319,N_5807);
nor U11143 (N_11143,N_5000,N_2154);
nor U11144 (N_11144,N_158,N_3983);
or U11145 (N_11145,N_4595,N_2694);
nor U11146 (N_11146,N_725,N_907);
and U11147 (N_11147,N_546,N_1791);
xor U11148 (N_11148,N_5338,N_3949);
nand U11149 (N_11149,N_4328,N_317);
xor U11150 (N_11150,N_1145,N_1193);
nor U11151 (N_11151,N_3666,N_5075);
nand U11152 (N_11152,N_3023,N_249);
nand U11153 (N_11153,N_4598,N_5382);
or U11154 (N_11154,N_4570,N_4385);
nor U11155 (N_11155,N_1000,N_84);
nand U11156 (N_11156,N_4436,N_4548);
nor U11157 (N_11157,N_3505,N_1992);
nand U11158 (N_11158,N_2666,N_5308);
or U11159 (N_11159,N_5858,N_2889);
xor U11160 (N_11160,N_1410,N_1755);
and U11161 (N_11161,N_4812,N_5780);
xnor U11162 (N_11162,N_5435,N_5331);
xor U11163 (N_11163,N_5547,N_2199);
or U11164 (N_11164,N_2574,N_3114);
nor U11165 (N_11165,N_3108,N_1710);
and U11166 (N_11166,N_4873,N_119);
and U11167 (N_11167,N_484,N_4515);
nor U11168 (N_11168,N_2749,N_2058);
or U11169 (N_11169,N_5712,N_4728);
nor U11170 (N_11170,N_833,N_5222);
nor U11171 (N_11171,N_5681,N_3152);
or U11172 (N_11172,N_3774,N_4887);
nand U11173 (N_11173,N_3326,N_2937);
xor U11174 (N_11174,N_803,N_192);
xnor U11175 (N_11175,N_5135,N_1351);
and U11176 (N_11176,N_1503,N_2851);
nand U11177 (N_11177,N_5556,N_5900);
and U11178 (N_11178,N_3755,N_1535);
nand U11179 (N_11179,N_2942,N_1383);
nand U11180 (N_11180,N_4825,N_1214);
and U11181 (N_11181,N_228,N_986);
nor U11182 (N_11182,N_4348,N_3685);
and U11183 (N_11183,N_2001,N_1787);
nand U11184 (N_11184,N_5533,N_1486);
or U11185 (N_11185,N_56,N_1186);
or U11186 (N_11186,N_3358,N_903);
nor U11187 (N_11187,N_1769,N_1922);
nand U11188 (N_11188,N_39,N_5208);
and U11189 (N_11189,N_3830,N_5689);
and U11190 (N_11190,N_2215,N_950);
nor U11191 (N_11191,N_3953,N_4538);
or U11192 (N_11192,N_1254,N_1631);
xnor U11193 (N_11193,N_2939,N_2890);
and U11194 (N_11194,N_2408,N_5440);
nand U11195 (N_11195,N_4882,N_5736);
nand U11196 (N_11196,N_3415,N_1917);
nor U11197 (N_11197,N_1177,N_4584);
nand U11198 (N_11198,N_232,N_4486);
xor U11199 (N_11199,N_915,N_424);
or U11200 (N_11200,N_2788,N_4556);
or U11201 (N_11201,N_3987,N_5942);
nand U11202 (N_11202,N_3253,N_1344);
nor U11203 (N_11203,N_245,N_755);
and U11204 (N_11204,N_3376,N_5031);
nor U11205 (N_11205,N_5760,N_2730);
xnor U11206 (N_11206,N_3063,N_82);
or U11207 (N_11207,N_5892,N_5935);
nor U11208 (N_11208,N_2454,N_5927);
nor U11209 (N_11209,N_5302,N_4744);
nor U11210 (N_11210,N_5720,N_439);
and U11211 (N_11211,N_521,N_5676);
nand U11212 (N_11212,N_5632,N_4359);
xnor U11213 (N_11213,N_1283,N_5903);
xor U11214 (N_11214,N_1871,N_2244);
xor U11215 (N_11215,N_1293,N_3352);
nand U11216 (N_11216,N_5693,N_3012);
nor U11217 (N_11217,N_2471,N_4941);
nor U11218 (N_11218,N_5775,N_1324);
and U11219 (N_11219,N_3790,N_2339);
xnor U11220 (N_11220,N_2202,N_88);
or U11221 (N_11221,N_335,N_4633);
and U11222 (N_11222,N_1761,N_3103);
nand U11223 (N_11223,N_3859,N_4771);
nor U11224 (N_11224,N_500,N_3282);
xnor U11225 (N_11225,N_3712,N_4917);
xnor U11226 (N_11226,N_4372,N_936);
nor U11227 (N_11227,N_1657,N_4120);
nor U11228 (N_11228,N_3430,N_2143);
or U11229 (N_11229,N_3579,N_4898);
nand U11230 (N_11230,N_2369,N_355);
or U11231 (N_11231,N_745,N_113);
and U11232 (N_11232,N_4952,N_3983);
nand U11233 (N_11233,N_3398,N_5903);
nor U11234 (N_11234,N_4148,N_3855);
nor U11235 (N_11235,N_3300,N_2463);
and U11236 (N_11236,N_5820,N_2152);
nand U11237 (N_11237,N_2134,N_4345);
nand U11238 (N_11238,N_4071,N_4485);
nor U11239 (N_11239,N_5300,N_281);
nor U11240 (N_11240,N_3141,N_2104);
and U11241 (N_11241,N_1193,N_1314);
nand U11242 (N_11242,N_1597,N_1300);
and U11243 (N_11243,N_2113,N_4033);
nand U11244 (N_11244,N_5603,N_1346);
or U11245 (N_11245,N_919,N_4755);
or U11246 (N_11246,N_2833,N_2362);
or U11247 (N_11247,N_3985,N_1497);
xor U11248 (N_11248,N_1881,N_3214);
or U11249 (N_11249,N_3119,N_2145);
nor U11250 (N_11250,N_4861,N_4097);
and U11251 (N_11251,N_1967,N_3232);
or U11252 (N_11252,N_5531,N_4667);
nor U11253 (N_11253,N_1656,N_1256);
xor U11254 (N_11254,N_2596,N_5496);
nor U11255 (N_11255,N_3591,N_3674);
xor U11256 (N_11256,N_2106,N_5299);
nand U11257 (N_11257,N_4303,N_3075);
xnor U11258 (N_11258,N_1633,N_2707);
nor U11259 (N_11259,N_1801,N_403);
or U11260 (N_11260,N_5842,N_3291);
nand U11261 (N_11261,N_5573,N_1918);
and U11262 (N_11262,N_2224,N_3149);
nand U11263 (N_11263,N_4044,N_4629);
xor U11264 (N_11264,N_37,N_2627);
nor U11265 (N_11265,N_3120,N_159);
nor U11266 (N_11266,N_2570,N_1914);
xnor U11267 (N_11267,N_2436,N_1060);
nor U11268 (N_11268,N_1929,N_4841);
xnor U11269 (N_11269,N_131,N_4395);
and U11270 (N_11270,N_4629,N_3103);
and U11271 (N_11271,N_1796,N_2336);
and U11272 (N_11272,N_1438,N_3471);
nor U11273 (N_11273,N_2558,N_1008);
xor U11274 (N_11274,N_5145,N_3931);
nand U11275 (N_11275,N_5177,N_3525);
or U11276 (N_11276,N_1004,N_2203);
nor U11277 (N_11277,N_5265,N_3055);
nand U11278 (N_11278,N_4399,N_5914);
and U11279 (N_11279,N_1593,N_819);
xnor U11280 (N_11280,N_4623,N_5688);
nor U11281 (N_11281,N_2875,N_2994);
and U11282 (N_11282,N_4931,N_1919);
xnor U11283 (N_11283,N_3282,N_5764);
nand U11284 (N_11284,N_3043,N_3946);
nand U11285 (N_11285,N_592,N_4868);
nand U11286 (N_11286,N_3960,N_3312);
xnor U11287 (N_11287,N_2761,N_2766);
nand U11288 (N_11288,N_3799,N_4225);
and U11289 (N_11289,N_5287,N_3924);
or U11290 (N_11290,N_4714,N_724);
and U11291 (N_11291,N_5787,N_2334);
and U11292 (N_11292,N_4097,N_3332);
nor U11293 (N_11293,N_13,N_2820);
or U11294 (N_11294,N_4744,N_2703);
or U11295 (N_11295,N_3987,N_5454);
nand U11296 (N_11296,N_635,N_444);
xor U11297 (N_11297,N_2000,N_2144);
xnor U11298 (N_11298,N_4524,N_2623);
and U11299 (N_11299,N_2261,N_3381);
nand U11300 (N_11300,N_2976,N_5761);
nand U11301 (N_11301,N_721,N_5672);
xor U11302 (N_11302,N_3277,N_5413);
xnor U11303 (N_11303,N_5269,N_5195);
or U11304 (N_11304,N_5152,N_4013);
nor U11305 (N_11305,N_3307,N_2532);
nor U11306 (N_11306,N_1968,N_5690);
or U11307 (N_11307,N_2885,N_1361);
and U11308 (N_11308,N_5489,N_1142);
xor U11309 (N_11309,N_930,N_5937);
and U11310 (N_11310,N_5040,N_3975);
and U11311 (N_11311,N_2227,N_5666);
nor U11312 (N_11312,N_5045,N_5476);
and U11313 (N_11313,N_3254,N_4349);
nor U11314 (N_11314,N_172,N_3877);
and U11315 (N_11315,N_1987,N_5376);
nand U11316 (N_11316,N_1436,N_2433);
nand U11317 (N_11317,N_592,N_1889);
nor U11318 (N_11318,N_2830,N_4630);
and U11319 (N_11319,N_2526,N_3722);
nand U11320 (N_11320,N_2393,N_4727);
and U11321 (N_11321,N_704,N_5756);
or U11322 (N_11322,N_4718,N_3975);
nand U11323 (N_11323,N_699,N_2869);
xnor U11324 (N_11324,N_2134,N_4591);
or U11325 (N_11325,N_4236,N_5399);
or U11326 (N_11326,N_1630,N_3744);
or U11327 (N_11327,N_1268,N_1639);
xor U11328 (N_11328,N_2790,N_766);
or U11329 (N_11329,N_2819,N_5950);
and U11330 (N_11330,N_1200,N_3143);
nand U11331 (N_11331,N_915,N_4267);
nor U11332 (N_11332,N_5238,N_4582);
nor U11333 (N_11333,N_998,N_3054);
xnor U11334 (N_11334,N_613,N_1492);
nand U11335 (N_11335,N_2603,N_5397);
xor U11336 (N_11336,N_4143,N_3472);
nor U11337 (N_11337,N_4417,N_2978);
or U11338 (N_11338,N_3324,N_5651);
nor U11339 (N_11339,N_5436,N_624);
nand U11340 (N_11340,N_3884,N_43);
xor U11341 (N_11341,N_2357,N_3616);
nor U11342 (N_11342,N_607,N_4965);
xor U11343 (N_11343,N_4963,N_739);
xor U11344 (N_11344,N_45,N_4854);
or U11345 (N_11345,N_2448,N_2763);
xor U11346 (N_11346,N_4299,N_2389);
or U11347 (N_11347,N_4279,N_5122);
nor U11348 (N_11348,N_2671,N_1511);
xor U11349 (N_11349,N_4760,N_1437);
nand U11350 (N_11350,N_4157,N_2937);
or U11351 (N_11351,N_4494,N_3973);
nor U11352 (N_11352,N_3465,N_2983);
nor U11353 (N_11353,N_4372,N_4868);
xnor U11354 (N_11354,N_5011,N_4370);
nand U11355 (N_11355,N_3534,N_781);
or U11356 (N_11356,N_2919,N_5737);
and U11357 (N_11357,N_5579,N_534);
and U11358 (N_11358,N_2896,N_1063);
or U11359 (N_11359,N_1593,N_4976);
and U11360 (N_11360,N_2542,N_3333);
xor U11361 (N_11361,N_202,N_1869);
nand U11362 (N_11362,N_3498,N_670);
and U11363 (N_11363,N_3639,N_1339);
xor U11364 (N_11364,N_5319,N_1447);
nor U11365 (N_11365,N_4964,N_1500);
or U11366 (N_11366,N_19,N_237);
nand U11367 (N_11367,N_859,N_2789);
nor U11368 (N_11368,N_5131,N_1725);
nor U11369 (N_11369,N_2719,N_988);
or U11370 (N_11370,N_2497,N_1210);
or U11371 (N_11371,N_873,N_2274);
nor U11372 (N_11372,N_2520,N_1233);
xor U11373 (N_11373,N_4583,N_75);
or U11374 (N_11374,N_3546,N_1501);
nor U11375 (N_11375,N_4201,N_271);
nor U11376 (N_11376,N_5,N_166);
xnor U11377 (N_11377,N_822,N_815);
or U11378 (N_11378,N_3300,N_4673);
nor U11379 (N_11379,N_5038,N_20);
or U11380 (N_11380,N_634,N_4266);
or U11381 (N_11381,N_1443,N_663);
nor U11382 (N_11382,N_1006,N_1197);
nand U11383 (N_11383,N_2079,N_813);
or U11384 (N_11384,N_1043,N_1136);
nor U11385 (N_11385,N_3222,N_1201);
nand U11386 (N_11386,N_2198,N_5222);
or U11387 (N_11387,N_2090,N_2028);
or U11388 (N_11388,N_5780,N_1107);
and U11389 (N_11389,N_1783,N_4143);
and U11390 (N_11390,N_4040,N_3861);
nor U11391 (N_11391,N_4912,N_3712);
or U11392 (N_11392,N_5434,N_2517);
and U11393 (N_11393,N_1204,N_52);
nor U11394 (N_11394,N_3738,N_4341);
or U11395 (N_11395,N_1115,N_5957);
or U11396 (N_11396,N_2436,N_2688);
and U11397 (N_11397,N_3315,N_2072);
and U11398 (N_11398,N_3019,N_4779);
xnor U11399 (N_11399,N_106,N_3221);
nand U11400 (N_11400,N_4695,N_2924);
nor U11401 (N_11401,N_193,N_4960);
or U11402 (N_11402,N_4327,N_929);
nand U11403 (N_11403,N_5469,N_3677);
xor U11404 (N_11404,N_1566,N_1516);
nand U11405 (N_11405,N_2195,N_546);
nand U11406 (N_11406,N_4262,N_4119);
and U11407 (N_11407,N_5236,N_3392);
or U11408 (N_11408,N_4145,N_432);
and U11409 (N_11409,N_2139,N_3622);
xnor U11410 (N_11410,N_4233,N_722);
xnor U11411 (N_11411,N_1476,N_5608);
xnor U11412 (N_11412,N_4700,N_1666);
and U11413 (N_11413,N_727,N_2879);
or U11414 (N_11414,N_3193,N_2030);
and U11415 (N_11415,N_716,N_3045);
xnor U11416 (N_11416,N_1644,N_5172);
nand U11417 (N_11417,N_2807,N_995);
xor U11418 (N_11418,N_917,N_1486);
or U11419 (N_11419,N_4983,N_3927);
xnor U11420 (N_11420,N_4417,N_3745);
or U11421 (N_11421,N_1253,N_3474);
or U11422 (N_11422,N_5602,N_1530);
nand U11423 (N_11423,N_3560,N_5896);
nor U11424 (N_11424,N_654,N_2439);
or U11425 (N_11425,N_2187,N_5041);
nand U11426 (N_11426,N_4735,N_4891);
xor U11427 (N_11427,N_1157,N_1904);
or U11428 (N_11428,N_1745,N_4400);
nor U11429 (N_11429,N_4946,N_3998);
nor U11430 (N_11430,N_3025,N_5873);
and U11431 (N_11431,N_4704,N_2298);
nor U11432 (N_11432,N_5460,N_2429);
or U11433 (N_11433,N_5361,N_2291);
nor U11434 (N_11434,N_634,N_5075);
xor U11435 (N_11435,N_4138,N_3712);
nand U11436 (N_11436,N_1273,N_1462);
and U11437 (N_11437,N_2996,N_3031);
nand U11438 (N_11438,N_2825,N_157);
nor U11439 (N_11439,N_1118,N_929);
xnor U11440 (N_11440,N_898,N_4756);
and U11441 (N_11441,N_5596,N_5957);
nor U11442 (N_11442,N_319,N_2175);
nor U11443 (N_11443,N_4852,N_5300);
and U11444 (N_11444,N_3413,N_468);
xor U11445 (N_11445,N_293,N_223);
nor U11446 (N_11446,N_823,N_3652);
xnor U11447 (N_11447,N_5514,N_5695);
nor U11448 (N_11448,N_382,N_202);
nor U11449 (N_11449,N_4108,N_4913);
and U11450 (N_11450,N_750,N_783);
nor U11451 (N_11451,N_328,N_2718);
xnor U11452 (N_11452,N_895,N_3180);
nor U11453 (N_11453,N_5666,N_4076);
and U11454 (N_11454,N_4446,N_57);
and U11455 (N_11455,N_2611,N_5788);
and U11456 (N_11456,N_4527,N_2539);
and U11457 (N_11457,N_144,N_319);
nor U11458 (N_11458,N_1570,N_4065);
nor U11459 (N_11459,N_5149,N_5006);
xor U11460 (N_11460,N_1476,N_93);
or U11461 (N_11461,N_2199,N_268);
nor U11462 (N_11462,N_4308,N_4759);
or U11463 (N_11463,N_5598,N_1617);
nor U11464 (N_11464,N_3469,N_624);
and U11465 (N_11465,N_3879,N_2402);
nor U11466 (N_11466,N_4644,N_140);
and U11467 (N_11467,N_2501,N_4837);
nor U11468 (N_11468,N_2420,N_5062);
nand U11469 (N_11469,N_1886,N_1175);
or U11470 (N_11470,N_2843,N_5575);
nor U11471 (N_11471,N_3606,N_946);
nand U11472 (N_11472,N_3590,N_1044);
nand U11473 (N_11473,N_1835,N_5274);
and U11474 (N_11474,N_1814,N_5367);
or U11475 (N_11475,N_2057,N_3979);
and U11476 (N_11476,N_2350,N_3090);
and U11477 (N_11477,N_4872,N_1546);
nor U11478 (N_11478,N_1909,N_3575);
nand U11479 (N_11479,N_5992,N_3285);
nand U11480 (N_11480,N_905,N_975);
nand U11481 (N_11481,N_1898,N_998);
or U11482 (N_11482,N_2371,N_2224);
nand U11483 (N_11483,N_174,N_5722);
and U11484 (N_11484,N_233,N_2163);
nand U11485 (N_11485,N_4663,N_5025);
or U11486 (N_11486,N_1195,N_101);
nand U11487 (N_11487,N_2126,N_3330);
or U11488 (N_11488,N_3677,N_5930);
nand U11489 (N_11489,N_2645,N_4289);
nand U11490 (N_11490,N_1504,N_3617);
xor U11491 (N_11491,N_1773,N_1302);
or U11492 (N_11492,N_5650,N_5305);
nand U11493 (N_11493,N_2831,N_3798);
nand U11494 (N_11494,N_422,N_3741);
xnor U11495 (N_11495,N_3904,N_5877);
xor U11496 (N_11496,N_5423,N_1039);
or U11497 (N_11497,N_1887,N_4705);
or U11498 (N_11498,N_1896,N_2084);
or U11499 (N_11499,N_1051,N_3165);
nand U11500 (N_11500,N_2768,N_4864);
and U11501 (N_11501,N_1394,N_4030);
xor U11502 (N_11502,N_1846,N_442);
nor U11503 (N_11503,N_3960,N_4134);
and U11504 (N_11504,N_4338,N_1859);
or U11505 (N_11505,N_4391,N_2816);
or U11506 (N_11506,N_3371,N_3411);
or U11507 (N_11507,N_5380,N_761);
nor U11508 (N_11508,N_3731,N_910);
and U11509 (N_11509,N_5389,N_2313);
nor U11510 (N_11510,N_3975,N_1141);
nand U11511 (N_11511,N_5401,N_5690);
nand U11512 (N_11512,N_3918,N_1302);
nand U11513 (N_11513,N_2729,N_2711);
or U11514 (N_11514,N_236,N_143);
xnor U11515 (N_11515,N_4965,N_5552);
nand U11516 (N_11516,N_85,N_4322);
or U11517 (N_11517,N_4071,N_2069);
and U11518 (N_11518,N_4642,N_392);
xnor U11519 (N_11519,N_3145,N_4143);
nand U11520 (N_11520,N_4677,N_30);
or U11521 (N_11521,N_3512,N_1427);
xnor U11522 (N_11522,N_4114,N_3480);
nor U11523 (N_11523,N_4229,N_4340);
and U11524 (N_11524,N_3296,N_3406);
nor U11525 (N_11525,N_4353,N_2546);
xnor U11526 (N_11526,N_4952,N_5529);
nor U11527 (N_11527,N_2294,N_1551);
nand U11528 (N_11528,N_5274,N_3100);
and U11529 (N_11529,N_2014,N_5267);
nand U11530 (N_11530,N_956,N_727);
and U11531 (N_11531,N_2694,N_3029);
nor U11532 (N_11532,N_4168,N_5620);
or U11533 (N_11533,N_1892,N_2766);
and U11534 (N_11534,N_4011,N_4872);
or U11535 (N_11535,N_295,N_2799);
nor U11536 (N_11536,N_2797,N_780);
nand U11537 (N_11537,N_2170,N_4314);
nand U11538 (N_11538,N_4530,N_4853);
nand U11539 (N_11539,N_4983,N_514);
nand U11540 (N_11540,N_2617,N_2717);
nand U11541 (N_11541,N_1204,N_5189);
or U11542 (N_11542,N_2431,N_5085);
xor U11543 (N_11543,N_2544,N_4912);
or U11544 (N_11544,N_671,N_2338);
nand U11545 (N_11545,N_3348,N_1162);
nand U11546 (N_11546,N_2578,N_173);
nor U11547 (N_11547,N_4952,N_5097);
xnor U11548 (N_11548,N_5531,N_1336);
nand U11549 (N_11549,N_4515,N_2084);
xor U11550 (N_11550,N_1980,N_4977);
or U11551 (N_11551,N_4678,N_2828);
nor U11552 (N_11552,N_5797,N_2230);
nor U11553 (N_11553,N_1776,N_5407);
xor U11554 (N_11554,N_4121,N_377);
nor U11555 (N_11555,N_4790,N_3652);
nand U11556 (N_11556,N_671,N_5013);
xnor U11557 (N_11557,N_431,N_1294);
nor U11558 (N_11558,N_5628,N_4775);
nand U11559 (N_11559,N_2946,N_1054);
nor U11560 (N_11560,N_2907,N_4587);
nor U11561 (N_11561,N_4223,N_5585);
and U11562 (N_11562,N_4524,N_2476);
and U11563 (N_11563,N_894,N_1754);
nand U11564 (N_11564,N_4048,N_5403);
and U11565 (N_11565,N_5875,N_4774);
xor U11566 (N_11566,N_3954,N_1810);
or U11567 (N_11567,N_2787,N_1373);
nor U11568 (N_11568,N_94,N_1504);
nor U11569 (N_11569,N_2479,N_1670);
xnor U11570 (N_11570,N_1840,N_3094);
or U11571 (N_11571,N_1008,N_418);
xnor U11572 (N_11572,N_5492,N_385);
nand U11573 (N_11573,N_1179,N_4109);
or U11574 (N_11574,N_4765,N_2738);
nor U11575 (N_11575,N_2370,N_4082);
nor U11576 (N_11576,N_1869,N_2057);
nand U11577 (N_11577,N_5326,N_4805);
or U11578 (N_11578,N_2913,N_476);
and U11579 (N_11579,N_3886,N_688);
or U11580 (N_11580,N_4415,N_4876);
nand U11581 (N_11581,N_5430,N_754);
and U11582 (N_11582,N_2655,N_5629);
nor U11583 (N_11583,N_1988,N_662);
xor U11584 (N_11584,N_2456,N_3339);
nand U11585 (N_11585,N_469,N_1836);
nor U11586 (N_11586,N_3382,N_4753);
and U11587 (N_11587,N_2288,N_5701);
and U11588 (N_11588,N_283,N_2877);
nor U11589 (N_11589,N_5471,N_981);
nand U11590 (N_11590,N_266,N_3383);
nor U11591 (N_11591,N_4038,N_1813);
xnor U11592 (N_11592,N_5733,N_1602);
xnor U11593 (N_11593,N_5151,N_3829);
or U11594 (N_11594,N_842,N_3484);
nor U11595 (N_11595,N_5046,N_2015);
and U11596 (N_11596,N_5054,N_2020);
and U11597 (N_11597,N_5311,N_1560);
nor U11598 (N_11598,N_5609,N_900);
and U11599 (N_11599,N_2296,N_2068);
nor U11600 (N_11600,N_4091,N_5581);
nor U11601 (N_11601,N_2298,N_3470);
xor U11602 (N_11602,N_2742,N_5448);
xnor U11603 (N_11603,N_1426,N_339);
xnor U11604 (N_11604,N_1597,N_2793);
nor U11605 (N_11605,N_2358,N_836);
xnor U11606 (N_11606,N_5533,N_3332);
xor U11607 (N_11607,N_2409,N_5600);
or U11608 (N_11608,N_524,N_4468);
nand U11609 (N_11609,N_117,N_1091);
xor U11610 (N_11610,N_2845,N_4785);
nor U11611 (N_11611,N_317,N_5124);
nor U11612 (N_11612,N_5068,N_2271);
xor U11613 (N_11613,N_1440,N_41);
nand U11614 (N_11614,N_1910,N_4778);
or U11615 (N_11615,N_1161,N_3941);
nand U11616 (N_11616,N_3995,N_3731);
nor U11617 (N_11617,N_5464,N_5439);
nor U11618 (N_11618,N_5892,N_5718);
nor U11619 (N_11619,N_1289,N_3798);
xnor U11620 (N_11620,N_2622,N_5682);
xor U11621 (N_11621,N_558,N_5849);
and U11622 (N_11622,N_3826,N_5005);
nand U11623 (N_11623,N_333,N_717);
xor U11624 (N_11624,N_3886,N_5965);
or U11625 (N_11625,N_5479,N_2732);
and U11626 (N_11626,N_2887,N_2543);
or U11627 (N_11627,N_1270,N_3976);
nor U11628 (N_11628,N_5201,N_4696);
xor U11629 (N_11629,N_4956,N_3520);
nor U11630 (N_11630,N_5134,N_3363);
and U11631 (N_11631,N_1758,N_1992);
xnor U11632 (N_11632,N_5600,N_5487);
nor U11633 (N_11633,N_1020,N_5830);
or U11634 (N_11634,N_2554,N_3623);
or U11635 (N_11635,N_4493,N_2482);
nand U11636 (N_11636,N_5510,N_4193);
or U11637 (N_11637,N_4980,N_4433);
xor U11638 (N_11638,N_2847,N_4026);
nand U11639 (N_11639,N_5195,N_2519);
xor U11640 (N_11640,N_5860,N_4223);
nor U11641 (N_11641,N_2392,N_1855);
and U11642 (N_11642,N_3091,N_5030);
and U11643 (N_11643,N_2978,N_2042);
xnor U11644 (N_11644,N_5220,N_5370);
nor U11645 (N_11645,N_2503,N_3232);
xor U11646 (N_11646,N_1824,N_5652);
nand U11647 (N_11647,N_1491,N_3316);
nand U11648 (N_11648,N_3403,N_3589);
and U11649 (N_11649,N_5637,N_5495);
nor U11650 (N_11650,N_2779,N_4363);
nor U11651 (N_11651,N_5484,N_3029);
and U11652 (N_11652,N_524,N_2151);
nand U11653 (N_11653,N_2644,N_1090);
or U11654 (N_11654,N_3867,N_4658);
xor U11655 (N_11655,N_5951,N_2691);
and U11656 (N_11656,N_4422,N_2321);
xor U11657 (N_11657,N_5349,N_333);
and U11658 (N_11658,N_1126,N_75);
nor U11659 (N_11659,N_3075,N_1503);
nor U11660 (N_11660,N_1003,N_2020);
xnor U11661 (N_11661,N_4867,N_1992);
or U11662 (N_11662,N_1954,N_3388);
and U11663 (N_11663,N_2272,N_4009);
xnor U11664 (N_11664,N_4082,N_4112);
and U11665 (N_11665,N_5976,N_4177);
nor U11666 (N_11666,N_2666,N_621);
and U11667 (N_11667,N_1255,N_4400);
or U11668 (N_11668,N_2649,N_4851);
and U11669 (N_11669,N_5887,N_5606);
or U11670 (N_11670,N_5241,N_1772);
or U11671 (N_11671,N_3406,N_2336);
and U11672 (N_11672,N_3977,N_3573);
xnor U11673 (N_11673,N_4143,N_3504);
or U11674 (N_11674,N_3873,N_137);
nand U11675 (N_11675,N_2335,N_5892);
xor U11676 (N_11676,N_1960,N_4827);
xor U11677 (N_11677,N_5977,N_2007);
or U11678 (N_11678,N_5933,N_3591);
or U11679 (N_11679,N_4162,N_2330);
nand U11680 (N_11680,N_312,N_3397);
or U11681 (N_11681,N_4160,N_1621);
nand U11682 (N_11682,N_777,N_1989);
xnor U11683 (N_11683,N_5151,N_2966);
and U11684 (N_11684,N_3621,N_468);
and U11685 (N_11685,N_5452,N_3608);
nand U11686 (N_11686,N_5682,N_2328);
xnor U11687 (N_11687,N_2256,N_3032);
nor U11688 (N_11688,N_2534,N_1226);
and U11689 (N_11689,N_2327,N_930);
nor U11690 (N_11690,N_731,N_2592);
nor U11691 (N_11691,N_691,N_4510);
or U11692 (N_11692,N_3326,N_2035);
nand U11693 (N_11693,N_1797,N_5243);
nand U11694 (N_11694,N_3139,N_4245);
nor U11695 (N_11695,N_5107,N_2781);
and U11696 (N_11696,N_693,N_526);
nor U11697 (N_11697,N_4689,N_4022);
or U11698 (N_11698,N_3500,N_4473);
or U11699 (N_11699,N_865,N_4325);
and U11700 (N_11700,N_566,N_5841);
nand U11701 (N_11701,N_4465,N_4956);
and U11702 (N_11702,N_2415,N_892);
nand U11703 (N_11703,N_3580,N_5968);
and U11704 (N_11704,N_554,N_2845);
xor U11705 (N_11705,N_4205,N_5987);
xnor U11706 (N_11706,N_2864,N_4990);
nor U11707 (N_11707,N_4582,N_1437);
nand U11708 (N_11708,N_5930,N_3313);
nor U11709 (N_11709,N_3783,N_1089);
nor U11710 (N_11710,N_5410,N_464);
nor U11711 (N_11711,N_346,N_980);
nand U11712 (N_11712,N_1220,N_4894);
nor U11713 (N_11713,N_4057,N_5717);
nand U11714 (N_11714,N_1281,N_2798);
and U11715 (N_11715,N_4999,N_4386);
and U11716 (N_11716,N_1682,N_3642);
xor U11717 (N_11717,N_2987,N_1752);
xor U11718 (N_11718,N_560,N_5889);
nor U11719 (N_11719,N_4752,N_922);
nand U11720 (N_11720,N_3598,N_545);
and U11721 (N_11721,N_4275,N_3112);
xnor U11722 (N_11722,N_5393,N_4951);
nor U11723 (N_11723,N_1829,N_1096);
or U11724 (N_11724,N_5656,N_2974);
nor U11725 (N_11725,N_3281,N_1043);
or U11726 (N_11726,N_5707,N_3242);
and U11727 (N_11727,N_1603,N_463);
xnor U11728 (N_11728,N_2100,N_5974);
nand U11729 (N_11729,N_3946,N_2177);
or U11730 (N_11730,N_1988,N_5244);
and U11731 (N_11731,N_4505,N_626);
and U11732 (N_11732,N_1046,N_3848);
xnor U11733 (N_11733,N_5209,N_5648);
and U11734 (N_11734,N_4145,N_5288);
nor U11735 (N_11735,N_317,N_1231);
or U11736 (N_11736,N_1889,N_3971);
nand U11737 (N_11737,N_1706,N_4435);
and U11738 (N_11738,N_3439,N_5276);
and U11739 (N_11739,N_2912,N_5458);
nand U11740 (N_11740,N_4432,N_1023);
xor U11741 (N_11741,N_4114,N_2120);
or U11742 (N_11742,N_1382,N_2169);
nand U11743 (N_11743,N_5905,N_2792);
and U11744 (N_11744,N_3009,N_5827);
nor U11745 (N_11745,N_3252,N_1565);
and U11746 (N_11746,N_4081,N_5082);
or U11747 (N_11747,N_5464,N_2512);
or U11748 (N_11748,N_84,N_5632);
nor U11749 (N_11749,N_2275,N_2832);
nand U11750 (N_11750,N_1813,N_3685);
nand U11751 (N_11751,N_1053,N_1635);
nand U11752 (N_11752,N_130,N_921);
and U11753 (N_11753,N_5528,N_5688);
or U11754 (N_11754,N_532,N_1567);
nor U11755 (N_11755,N_5748,N_5495);
xor U11756 (N_11756,N_4782,N_2935);
or U11757 (N_11757,N_5188,N_2007);
and U11758 (N_11758,N_3814,N_3079);
and U11759 (N_11759,N_3941,N_4936);
or U11760 (N_11760,N_436,N_3754);
nor U11761 (N_11761,N_236,N_5117);
xnor U11762 (N_11762,N_3283,N_2013);
xnor U11763 (N_11763,N_930,N_3942);
nor U11764 (N_11764,N_3760,N_2366);
nand U11765 (N_11765,N_3955,N_116);
xor U11766 (N_11766,N_3107,N_3935);
xnor U11767 (N_11767,N_2417,N_1429);
and U11768 (N_11768,N_4852,N_607);
or U11769 (N_11769,N_2741,N_1451);
nand U11770 (N_11770,N_5746,N_3135);
nor U11771 (N_11771,N_1836,N_3178);
xor U11772 (N_11772,N_5438,N_760);
xor U11773 (N_11773,N_1466,N_3950);
nand U11774 (N_11774,N_4460,N_3747);
nor U11775 (N_11775,N_2391,N_975);
nor U11776 (N_11776,N_369,N_4684);
xor U11777 (N_11777,N_101,N_2170);
xor U11778 (N_11778,N_3798,N_195);
and U11779 (N_11779,N_4769,N_3569);
nand U11780 (N_11780,N_880,N_2472);
and U11781 (N_11781,N_806,N_3657);
or U11782 (N_11782,N_2808,N_4753);
and U11783 (N_11783,N_5883,N_5095);
xnor U11784 (N_11784,N_3907,N_5639);
xnor U11785 (N_11785,N_1524,N_1913);
nor U11786 (N_11786,N_3978,N_2885);
and U11787 (N_11787,N_128,N_4164);
nor U11788 (N_11788,N_5143,N_5409);
xor U11789 (N_11789,N_1099,N_2667);
and U11790 (N_11790,N_2670,N_2329);
nor U11791 (N_11791,N_1158,N_1045);
xor U11792 (N_11792,N_5270,N_4403);
or U11793 (N_11793,N_5809,N_4067);
xor U11794 (N_11794,N_267,N_4996);
xor U11795 (N_11795,N_1588,N_4210);
or U11796 (N_11796,N_1823,N_1828);
xor U11797 (N_11797,N_4783,N_1097);
or U11798 (N_11798,N_3345,N_2721);
or U11799 (N_11799,N_5067,N_3145);
nor U11800 (N_11800,N_176,N_5113);
or U11801 (N_11801,N_1117,N_4687);
xnor U11802 (N_11802,N_5162,N_4894);
or U11803 (N_11803,N_5253,N_4687);
nor U11804 (N_11804,N_4465,N_5073);
or U11805 (N_11805,N_3387,N_2644);
or U11806 (N_11806,N_5924,N_2756);
nand U11807 (N_11807,N_3413,N_3543);
nor U11808 (N_11808,N_732,N_3913);
xnor U11809 (N_11809,N_6,N_4620);
nor U11810 (N_11810,N_4814,N_3357);
nand U11811 (N_11811,N_1681,N_3347);
or U11812 (N_11812,N_4949,N_959);
nand U11813 (N_11813,N_4629,N_5059);
or U11814 (N_11814,N_2694,N_5204);
or U11815 (N_11815,N_2678,N_2455);
nand U11816 (N_11816,N_4687,N_2583);
xor U11817 (N_11817,N_4898,N_5760);
and U11818 (N_11818,N_3627,N_914);
and U11819 (N_11819,N_2888,N_3944);
or U11820 (N_11820,N_3188,N_5313);
xnor U11821 (N_11821,N_2281,N_182);
and U11822 (N_11822,N_4393,N_162);
xnor U11823 (N_11823,N_3598,N_135);
nor U11824 (N_11824,N_718,N_3268);
and U11825 (N_11825,N_2182,N_1141);
nand U11826 (N_11826,N_1810,N_1327);
or U11827 (N_11827,N_80,N_5683);
nand U11828 (N_11828,N_4918,N_2030);
nand U11829 (N_11829,N_5153,N_4236);
nand U11830 (N_11830,N_43,N_3035);
nand U11831 (N_11831,N_2907,N_552);
nor U11832 (N_11832,N_4528,N_5593);
or U11833 (N_11833,N_2264,N_4867);
xor U11834 (N_11834,N_2684,N_5168);
nand U11835 (N_11835,N_5386,N_241);
or U11836 (N_11836,N_4789,N_4277);
xnor U11837 (N_11837,N_120,N_1164);
nand U11838 (N_11838,N_5423,N_984);
nor U11839 (N_11839,N_406,N_1845);
nand U11840 (N_11840,N_708,N_1875);
or U11841 (N_11841,N_3975,N_1648);
nand U11842 (N_11842,N_2090,N_3208);
nand U11843 (N_11843,N_2809,N_3911);
nand U11844 (N_11844,N_1041,N_2295);
nand U11845 (N_11845,N_1779,N_5292);
xor U11846 (N_11846,N_5287,N_3051);
nor U11847 (N_11847,N_2802,N_4381);
xor U11848 (N_11848,N_5593,N_1153);
and U11849 (N_11849,N_1561,N_5187);
nor U11850 (N_11850,N_651,N_3243);
xor U11851 (N_11851,N_5618,N_4152);
nor U11852 (N_11852,N_5768,N_3038);
or U11853 (N_11853,N_3034,N_1287);
xnor U11854 (N_11854,N_1366,N_1962);
nand U11855 (N_11855,N_396,N_5746);
nor U11856 (N_11856,N_4881,N_1605);
nor U11857 (N_11857,N_1416,N_3642);
and U11858 (N_11858,N_2625,N_3288);
and U11859 (N_11859,N_2016,N_2486);
and U11860 (N_11860,N_2351,N_2839);
nand U11861 (N_11861,N_844,N_1761);
nand U11862 (N_11862,N_1886,N_3999);
and U11863 (N_11863,N_3779,N_1640);
nand U11864 (N_11864,N_5649,N_4303);
nor U11865 (N_11865,N_5214,N_2518);
nor U11866 (N_11866,N_753,N_3203);
or U11867 (N_11867,N_10,N_5837);
or U11868 (N_11868,N_5919,N_956);
or U11869 (N_11869,N_5267,N_5685);
xnor U11870 (N_11870,N_1231,N_1970);
nor U11871 (N_11871,N_2192,N_2779);
or U11872 (N_11872,N_4308,N_273);
nor U11873 (N_11873,N_4618,N_1301);
nor U11874 (N_11874,N_512,N_3142);
nor U11875 (N_11875,N_2143,N_5027);
nand U11876 (N_11876,N_2236,N_5361);
xor U11877 (N_11877,N_4254,N_2902);
and U11878 (N_11878,N_2529,N_4493);
or U11879 (N_11879,N_5012,N_3377);
nand U11880 (N_11880,N_3788,N_4040);
and U11881 (N_11881,N_388,N_4802);
nor U11882 (N_11882,N_4965,N_2297);
nor U11883 (N_11883,N_1958,N_2381);
nor U11884 (N_11884,N_4325,N_2953);
nor U11885 (N_11885,N_4785,N_5065);
nor U11886 (N_11886,N_3195,N_5464);
and U11887 (N_11887,N_2533,N_5614);
and U11888 (N_11888,N_1973,N_4709);
or U11889 (N_11889,N_2432,N_3569);
nand U11890 (N_11890,N_2928,N_5486);
nand U11891 (N_11891,N_5336,N_5854);
nor U11892 (N_11892,N_2362,N_1643);
nand U11893 (N_11893,N_2070,N_3373);
nand U11894 (N_11894,N_392,N_5073);
and U11895 (N_11895,N_3521,N_761);
or U11896 (N_11896,N_576,N_854);
and U11897 (N_11897,N_2047,N_3941);
nand U11898 (N_11898,N_5192,N_1942);
xnor U11899 (N_11899,N_305,N_1932);
nor U11900 (N_11900,N_4961,N_3250);
nand U11901 (N_11901,N_3781,N_4778);
nand U11902 (N_11902,N_1174,N_3009);
or U11903 (N_11903,N_3405,N_110);
nor U11904 (N_11904,N_3573,N_4812);
and U11905 (N_11905,N_396,N_4035);
and U11906 (N_11906,N_1212,N_5543);
nand U11907 (N_11907,N_843,N_1581);
or U11908 (N_11908,N_3465,N_461);
nand U11909 (N_11909,N_3127,N_1516);
and U11910 (N_11910,N_3726,N_1037);
and U11911 (N_11911,N_3269,N_3748);
nand U11912 (N_11912,N_669,N_975);
nor U11913 (N_11913,N_5883,N_1186);
nor U11914 (N_11914,N_3713,N_378);
or U11915 (N_11915,N_4998,N_5779);
and U11916 (N_11916,N_852,N_1032);
nor U11917 (N_11917,N_3348,N_1431);
xnor U11918 (N_11918,N_4810,N_461);
or U11919 (N_11919,N_5859,N_1075);
xnor U11920 (N_11920,N_241,N_3423);
and U11921 (N_11921,N_2805,N_3024);
and U11922 (N_11922,N_712,N_5818);
xnor U11923 (N_11923,N_670,N_2983);
xor U11924 (N_11924,N_5031,N_522);
nand U11925 (N_11925,N_3085,N_713);
nand U11926 (N_11926,N_858,N_4383);
nor U11927 (N_11927,N_51,N_1783);
or U11928 (N_11928,N_4120,N_3174);
xor U11929 (N_11929,N_378,N_5079);
xnor U11930 (N_11930,N_4601,N_4377);
or U11931 (N_11931,N_4924,N_5769);
nor U11932 (N_11932,N_4799,N_5667);
and U11933 (N_11933,N_1384,N_2725);
nand U11934 (N_11934,N_4708,N_4753);
xor U11935 (N_11935,N_2643,N_5945);
and U11936 (N_11936,N_4644,N_3524);
and U11937 (N_11937,N_1060,N_5821);
nand U11938 (N_11938,N_3930,N_135);
xnor U11939 (N_11939,N_2604,N_2437);
nor U11940 (N_11940,N_1149,N_2144);
or U11941 (N_11941,N_1109,N_1775);
xor U11942 (N_11942,N_480,N_5747);
or U11943 (N_11943,N_605,N_2138);
and U11944 (N_11944,N_5685,N_2596);
nor U11945 (N_11945,N_3874,N_129);
nor U11946 (N_11946,N_1075,N_1534);
xnor U11947 (N_11947,N_5951,N_151);
xor U11948 (N_11948,N_5391,N_351);
nor U11949 (N_11949,N_1629,N_243);
or U11950 (N_11950,N_5824,N_4384);
xnor U11951 (N_11951,N_5053,N_4715);
and U11952 (N_11952,N_2689,N_3392);
or U11953 (N_11953,N_2761,N_4290);
or U11954 (N_11954,N_5598,N_3422);
and U11955 (N_11955,N_5226,N_5074);
nand U11956 (N_11956,N_3963,N_2966);
or U11957 (N_11957,N_5881,N_4160);
or U11958 (N_11958,N_2201,N_4217);
xor U11959 (N_11959,N_2448,N_1250);
nand U11960 (N_11960,N_1703,N_112);
xnor U11961 (N_11961,N_4456,N_1030);
nor U11962 (N_11962,N_2376,N_4893);
xnor U11963 (N_11963,N_3009,N_3993);
nor U11964 (N_11964,N_1603,N_2401);
and U11965 (N_11965,N_3622,N_2454);
and U11966 (N_11966,N_1135,N_2739);
xor U11967 (N_11967,N_2116,N_4298);
and U11968 (N_11968,N_2904,N_4043);
nand U11969 (N_11969,N_3431,N_2384);
or U11970 (N_11970,N_2110,N_4113);
nor U11971 (N_11971,N_5886,N_1846);
and U11972 (N_11972,N_3415,N_5312);
xnor U11973 (N_11973,N_5620,N_2578);
nor U11974 (N_11974,N_3255,N_555);
and U11975 (N_11975,N_2108,N_640);
xnor U11976 (N_11976,N_2237,N_2091);
and U11977 (N_11977,N_4521,N_2822);
and U11978 (N_11978,N_4916,N_1951);
and U11979 (N_11979,N_1366,N_2488);
nand U11980 (N_11980,N_878,N_82);
nand U11981 (N_11981,N_4092,N_825);
nand U11982 (N_11982,N_2550,N_1299);
nand U11983 (N_11983,N_2501,N_5215);
nor U11984 (N_11984,N_329,N_923);
nand U11985 (N_11985,N_3107,N_3429);
and U11986 (N_11986,N_3529,N_5931);
and U11987 (N_11987,N_2433,N_1288);
nor U11988 (N_11988,N_4617,N_4663);
xnor U11989 (N_11989,N_372,N_4493);
nor U11990 (N_11990,N_3451,N_2169);
nor U11991 (N_11991,N_5587,N_1150);
nor U11992 (N_11992,N_4062,N_913);
and U11993 (N_11993,N_780,N_4006);
xor U11994 (N_11994,N_5677,N_164);
nand U11995 (N_11995,N_268,N_3767);
and U11996 (N_11996,N_2601,N_5046);
and U11997 (N_11997,N_1505,N_4817);
and U11998 (N_11998,N_5208,N_1429);
and U11999 (N_11999,N_2502,N_2986);
nand U12000 (N_12000,N_10789,N_11752);
and U12001 (N_12001,N_10658,N_11997);
or U12002 (N_12002,N_7206,N_8694);
xor U12003 (N_12003,N_7804,N_9310);
or U12004 (N_12004,N_7064,N_6102);
xnor U12005 (N_12005,N_9600,N_10555);
or U12006 (N_12006,N_11322,N_7481);
and U12007 (N_12007,N_9775,N_8634);
and U12008 (N_12008,N_10408,N_11349);
and U12009 (N_12009,N_10994,N_6737);
nand U12010 (N_12010,N_8548,N_10147);
nand U12011 (N_12011,N_9466,N_6209);
nand U12012 (N_12012,N_8532,N_10048);
and U12013 (N_12013,N_9887,N_8627);
xor U12014 (N_12014,N_6065,N_6949);
nand U12015 (N_12015,N_9125,N_9474);
nor U12016 (N_12016,N_6628,N_10052);
or U12017 (N_12017,N_8941,N_7374);
and U12018 (N_12018,N_9024,N_11994);
xor U12019 (N_12019,N_6201,N_9587);
nor U12020 (N_12020,N_7928,N_10380);
or U12021 (N_12021,N_11974,N_6551);
and U12022 (N_12022,N_6786,N_6269);
xnor U12023 (N_12023,N_8693,N_9961);
xnor U12024 (N_12024,N_6071,N_10350);
and U12025 (N_12025,N_6147,N_7062);
and U12026 (N_12026,N_7801,N_10566);
and U12027 (N_12027,N_11145,N_10862);
xnor U12028 (N_12028,N_11666,N_6442);
and U12029 (N_12029,N_10636,N_10691);
or U12030 (N_12030,N_6649,N_9677);
nand U12031 (N_12031,N_6886,N_10511);
xnor U12032 (N_12032,N_8144,N_8954);
nand U12033 (N_12033,N_6327,N_7993);
xnor U12034 (N_12034,N_6146,N_11754);
nor U12035 (N_12035,N_7009,N_6471);
and U12036 (N_12036,N_8538,N_6832);
xor U12037 (N_12037,N_6695,N_9098);
nor U12038 (N_12038,N_6394,N_7234);
nor U12039 (N_12039,N_8471,N_6999);
nor U12040 (N_12040,N_11118,N_11646);
and U12041 (N_12041,N_9697,N_11124);
and U12042 (N_12042,N_9872,N_7645);
nand U12043 (N_12043,N_11150,N_8417);
xnor U12044 (N_12044,N_10410,N_11230);
nor U12045 (N_12045,N_7556,N_8608);
nand U12046 (N_12046,N_7070,N_11233);
or U12047 (N_12047,N_7001,N_6054);
and U12048 (N_12048,N_11846,N_11411);
xor U12049 (N_12049,N_11595,N_8728);
and U12050 (N_12050,N_6283,N_10438);
or U12051 (N_12051,N_9852,N_10565);
xnor U12052 (N_12052,N_9649,N_10064);
or U12053 (N_12053,N_6126,N_6485);
or U12054 (N_12054,N_6780,N_6337);
nor U12055 (N_12055,N_8796,N_9810);
and U12056 (N_12056,N_9150,N_11169);
nor U12057 (N_12057,N_9953,N_9228);
and U12058 (N_12058,N_8953,N_10311);
nand U12059 (N_12059,N_10361,N_7824);
or U12060 (N_12060,N_11177,N_9154);
xor U12061 (N_12061,N_9319,N_6399);
or U12062 (N_12062,N_11389,N_7133);
nor U12063 (N_12063,N_11797,N_8340);
nor U12064 (N_12064,N_8606,N_6747);
xor U12065 (N_12065,N_10663,N_7139);
and U12066 (N_12066,N_7337,N_6069);
and U12067 (N_12067,N_6166,N_6852);
nand U12068 (N_12068,N_11221,N_10314);
or U12069 (N_12069,N_9068,N_7386);
nand U12070 (N_12070,N_11417,N_7832);
or U12071 (N_12071,N_6908,N_8576);
nor U12072 (N_12072,N_11458,N_6084);
or U12073 (N_12073,N_8907,N_7171);
xor U12074 (N_12074,N_8345,N_7840);
and U12075 (N_12075,N_8853,N_7368);
or U12076 (N_12076,N_9740,N_7291);
and U12077 (N_12077,N_7532,N_10800);
xnor U12078 (N_12078,N_10540,N_6068);
or U12079 (N_12079,N_11825,N_11686);
nand U12080 (N_12080,N_10144,N_8360);
xnor U12081 (N_12081,N_7267,N_8162);
and U12082 (N_12082,N_9511,N_7641);
xnor U12083 (N_12083,N_11794,N_7710);
nand U12084 (N_12084,N_8879,N_8258);
nor U12085 (N_12085,N_10553,N_8985);
or U12086 (N_12086,N_9389,N_10864);
or U12087 (N_12087,N_6438,N_6866);
xor U12088 (N_12088,N_7246,N_11232);
xnor U12089 (N_12089,N_9182,N_6826);
xnor U12090 (N_12090,N_9042,N_10538);
xor U12091 (N_12091,N_7297,N_9843);
nand U12092 (N_12092,N_6312,N_8450);
and U12093 (N_12093,N_10074,N_6905);
nand U12094 (N_12094,N_10488,N_9665);
and U12095 (N_12095,N_9921,N_7751);
and U12096 (N_12096,N_6221,N_11911);
or U12097 (N_12097,N_7923,N_8821);
xnor U12098 (N_12098,N_7356,N_8633);
nor U12099 (N_12099,N_9922,N_6168);
nor U12100 (N_12100,N_11796,N_10925);
nand U12101 (N_12101,N_7771,N_11048);
or U12102 (N_12102,N_7213,N_7649);
nand U12103 (N_12103,N_8234,N_11981);
and U12104 (N_12104,N_11080,N_11712);
and U12105 (N_12105,N_10459,N_7398);
nand U12106 (N_12106,N_11379,N_7612);
or U12107 (N_12107,N_7992,N_10345);
and U12108 (N_12108,N_7421,N_8556);
and U12109 (N_12109,N_9929,N_7867);
and U12110 (N_12110,N_9427,N_11845);
nand U12111 (N_12111,N_6469,N_9160);
nand U12112 (N_12112,N_6322,N_10332);
and U12113 (N_12113,N_10582,N_11348);
or U12114 (N_12114,N_11394,N_8001);
or U12115 (N_12115,N_11902,N_10460);
or U12116 (N_12116,N_6413,N_8749);
and U12117 (N_12117,N_9472,N_7781);
xnor U12118 (N_12118,N_11901,N_6087);
nor U12119 (N_12119,N_10529,N_11332);
and U12120 (N_12120,N_7554,N_10547);
and U12121 (N_12121,N_8492,N_10336);
nand U12122 (N_12122,N_6597,N_8262);
nor U12123 (N_12123,N_6308,N_9006);
and U12124 (N_12124,N_10935,N_9351);
or U12125 (N_12125,N_9036,N_6770);
xnor U12126 (N_12126,N_6278,N_9670);
nor U12127 (N_12127,N_8295,N_9373);
and U12128 (N_12128,N_10567,N_8133);
and U12129 (N_12129,N_9315,N_9714);
nor U12130 (N_12130,N_11504,N_11953);
and U12131 (N_12131,N_10161,N_6768);
xnor U12132 (N_12132,N_11689,N_9540);
xor U12133 (N_12133,N_9314,N_11571);
xor U12134 (N_12134,N_9721,N_10727);
and U12135 (N_12135,N_6742,N_6000);
or U12136 (N_12136,N_8798,N_8324);
xor U12137 (N_12137,N_8638,N_10372);
xor U12138 (N_12138,N_9103,N_8169);
nand U12139 (N_12139,N_9205,N_7869);
nand U12140 (N_12140,N_7313,N_10146);
xor U12141 (N_12141,N_6564,N_10407);
or U12142 (N_12142,N_11226,N_10014);
and U12143 (N_12143,N_7365,N_8057);
or U12144 (N_12144,N_11347,N_6321);
nor U12145 (N_12145,N_10621,N_11256);
and U12146 (N_12146,N_9440,N_11333);
nor U12147 (N_12147,N_11721,N_8085);
and U12148 (N_12148,N_6834,N_10966);
nand U12149 (N_12149,N_8692,N_10398);
and U12150 (N_12150,N_6715,N_8355);
and U12151 (N_12151,N_7559,N_9443);
or U12152 (N_12152,N_6455,N_6678);
nor U12153 (N_12153,N_10677,N_6692);
nor U12154 (N_12154,N_11579,N_11893);
xor U12155 (N_12155,N_6427,N_9486);
xor U12156 (N_12156,N_10997,N_11302);
or U12157 (N_12157,N_6009,N_9331);
nand U12158 (N_12158,N_8134,N_11019);
nand U12159 (N_12159,N_10095,N_8736);
nor U12160 (N_12160,N_8838,N_8947);
or U12161 (N_12161,N_9590,N_6237);
or U12162 (N_12162,N_8462,N_7405);
nand U12163 (N_12163,N_9952,N_10448);
nand U12164 (N_12164,N_7930,N_11661);
or U12165 (N_12165,N_10055,N_8174);
and U12166 (N_12166,N_10153,N_10525);
nor U12167 (N_12167,N_11191,N_8404);
and U12168 (N_12168,N_6589,N_11099);
and U12169 (N_12169,N_11935,N_10382);
or U12170 (N_12170,N_8385,N_11438);
or U12171 (N_12171,N_8515,N_8058);
nor U12172 (N_12172,N_9989,N_7909);
and U12173 (N_12173,N_8280,N_6723);
or U12174 (N_12174,N_6453,N_6094);
xnor U12175 (N_12175,N_6985,N_6459);
and U12176 (N_12176,N_11231,N_7491);
nor U12177 (N_12177,N_9069,N_11321);
and U12178 (N_12178,N_7021,N_11878);
nor U12179 (N_12179,N_11636,N_8398);
nand U12180 (N_12180,N_9933,N_7798);
nor U12181 (N_12181,N_8210,N_11527);
xnor U12182 (N_12182,N_10115,N_8253);
nand U12183 (N_12183,N_10212,N_8709);
nor U12184 (N_12184,N_9772,N_8686);
xor U12185 (N_12185,N_11003,N_6344);
xnor U12186 (N_12186,N_11641,N_8766);
nand U12187 (N_12187,N_11532,N_10246);
nor U12188 (N_12188,N_8122,N_11128);
xnor U12189 (N_12189,N_8211,N_8096);
or U12190 (N_12190,N_8877,N_9761);
nand U12191 (N_12191,N_6284,N_10117);
and U12192 (N_12192,N_6402,N_8380);
nand U12193 (N_12193,N_9295,N_7024);
xor U12194 (N_12194,N_11996,N_10795);
nor U12195 (N_12195,N_11551,N_7716);
nor U12196 (N_12196,N_11082,N_6355);
nor U12197 (N_12197,N_7848,N_8504);
xor U12198 (N_12198,N_9192,N_7672);
xnor U12199 (N_12199,N_7647,N_6883);
xnor U12200 (N_12200,N_9029,N_9577);
xnor U12201 (N_12201,N_9884,N_10127);
and U12202 (N_12202,N_7066,N_8804);
nand U12203 (N_12203,N_6787,N_11097);
or U12204 (N_12204,N_10722,N_9559);
nor U12205 (N_12205,N_7477,N_8035);
xnor U12206 (N_12206,N_8668,N_11060);
nor U12207 (N_12207,N_9234,N_11783);
nor U12208 (N_12208,N_7553,N_8965);
nor U12209 (N_12209,N_7677,N_6566);
nand U12210 (N_12210,N_11753,N_9751);
nor U12211 (N_12211,N_9017,N_8042);
nor U12212 (N_12212,N_9488,N_10333);
nand U12213 (N_12213,N_11471,N_8614);
nand U12214 (N_12214,N_7224,N_11208);
xnor U12215 (N_12215,N_8010,N_7745);
nor U12216 (N_12216,N_8438,N_11229);
and U12217 (N_12217,N_11516,N_11310);
xor U12218 (N_12218,N_7425,N_9461);
nor U12219 (N_12219,N_8403,N_10785);
nor U12220 (N_12220,N_11172,N_7459);
xor U12221 (N_12221,N_8151,N_11605);
or U12222 (N_12222,N_8148,N_10417);
xor U12223 (N_12223,N_9289,N_7584);
nor U12224 (N_12224,N_8795,N_7843);
and U12225 (N_12225,N_6789,N_9400);
or U12226 (N_12226,N_6488,N_9716);
nor U12227 (N_12227,N_8282,N_7921);
and U12228 (N_12228,N_10443,N_9533);
or U12229 (N_12229,N_6726,N_9951);
xnor U12230 (N_12230,N_11599,N_9354);
or U12231 (N_12231,N_10317,N_8305);
nor U12232 (N_12232,N_9517,N_9841);
nand U12233 (N_12233,N_9912,N_10360);
xnor U12234 (N_12234,N_10330,N_6019);
nor U12235 (N_12235,N_7134,N_10834);
nor U12236 (N_12236,N_7306,N_6414);
xnor U12237 (N_12237,N_8507,N_10542);
or U12238 (N_12238,N_10131,N_7176);
nor U12239 (N_12239,N_6702,N_11523);
nor U12240 (N_12240,N_8537,N_8290);
or U12241 (N_12241,N_9814,N_7568);
nor U12242 (N_12242,N_6583,N_8554);
or U12243 (N_12243,N_11803,N_10958);
xnor U12244 (N_12244,N_6819,N_10701);
nand U12245 (N_12245,N_9366,N_8664);
or U12246 (N_12246,N_11759,N_10284);
and U12247 (N_12247,N_7805,N_11422);
and U12248 (N_12248,N_7115,N_8987);
or U12249 (N_12249,N_11216,N_7172);
xnor U12250 (N_12250,N_8284,N_10008);
xor U12251 (N_12251,N_11869,N_7655);
or U12252 (N_12252,N_8126,N_11919);
nand U12253 (N_12253,N_7366,N_9689);
or U12254 (N_12254,N_9717,N_11765);
or U12255 (N_12255,N_8191,N_11555);
and U12256 (N_12256,N_11359,N_9071);
nand U12257 (N_12257,N_9546,N_7452);
and U12258 (N_12258,N_7157,N_10541);
nor U12259 (N_12259,N_8195,N_9678);
xnor U12260 (N_12260,N_10085,N_7223);
xor U12261 (N_12261,N_9504,N_6401);
and U12262 (N_12262,N_8514,N_10174);
nor U12263 (N_12263,N_6875,N_8855);
nand U12264 (N_12264,N_11076,N_11001);
xnor U12265 (N_12265,N_11009,N_9759);
nand U12266 (N_12266,N_8106,N_6396);
or U12267 (N_12267,N_9877,N_9825);
or U12268 (N_12268,N_11300,N_8753);
nor U12269 (N_12269,N_11383,N_11676);
nand U12270 (N_12270,N_10025,N_7410);
and U12271 (N_12271,N_10442,N_6127);
nand U12272 (N_12272,N_7192,N_7943);
or U12273 (N_12273,N_8744,N_8760);
or U12274 (N_12274,N_7099,N_9112);
xnor U12275 (N_12275,N_11905,N_7834);
nand U12276 (N_12276,N_7307,N_7673);
or U12277 (N_12277,N_9861,N_10742);
and U12278 (N_12278,N_11669,N_7984);
and U12279 (N_12279,N_7377,N_10044);
xor U12280 (N_12280,N_6618,N_7599);
nor U12281 (N_12281,N_10287,N_10304);
nor U12282 (N_12282,N_9875,N_8392);
xor U12283 (N_12283,N_8223,N_7401);
or U12284 (N_12284,N_8715,N_11866);
nand U12285 (N_12285,N_9332,N_6689);
xnor U12286 (N_12286,N_9538,N_7621);
nor U12287 (N_12287,N_7911,N_11610);
or U12288 (N_12288,N_8726,N_7059);
xor U12289 (N_12289,N_9403,N_6579);
or U12290 (N_12290,N_6881,N_10165);
nand U12291 (N_12291,N_8797,N_11244);
and U12292 (N_12292,N_10392,N_10856);
nor U12293 (N_12293,N_8834,N_10463);
nand U12294 (N_12294,N_11263,N_6295);
nor U12295 (N_12295,N_8991,N_9652);
xor U12296 (N_12296,N_7714,N_9597);
or U12297 (N_12297,N_6808,N_8497);
and U12298 (N_12298,N_7428,N_9679);
nand U12299 (N_12299,N_10803,N_8416);
or U12300 (N_12300,N_8182,N_6090);
nor U12301 (N_12301,N_7232,N_8321);
or U12302 (N_12302,N_6149,N_11397);
or U12303 (N_12303,N_10937,N_8865);
and U12304 (N_12304,N_11518,N_10462);
and U12305 (N_12305,N_11985,N_11014);
or U12306 (N_12306,N_11988,N_11622);
nor U12307 (N_12307,N_8542,N_10404);
nand U12308 (N_12308,N_7123,N_11780);
xnor U12309 (N_12309,N_6630,N_8669);
nor U12310 (N_12310,N_10828,N_6182);
xnor U12311 (N_12311,N_9152,N_6220);
and U12312 (N_12312,N_9076,N_6740);
nand U12313 (N_12313,N_11679,N_7169);
nand U12314 (N_12314,N_10777,N_8955);
nor U12315 (N_12315,N_10647,N_7000);
nor U12316 (N_12316,N_9102,N_6226);
nand U12317 (N_12317,N_8289,N_6123);
xnor U12318 (N_12318,N_9762,N_8571);
xor U12319 (N_12319,N_11498,N_10781);
nor U12320 (N_12320,N_10851,N_8193);
or U12321 (N_12321,N_8044,N_6021);
and U12322 (N_12322,N_9371,N_10759);
or U12323 (N_12323,N_8286,N_6178);
xor U12324 (N_12324,N_9928,N_9745);
nand U12325 (N_12325,N_9446,N_9442);
or U12326 (N_12326,N_8255,N_10486);
nor U12327 (N_12327,N_10544,N_8929);
xor U12328 (N_12328,N_8917,N_8615);
and U12329 (N_12329,N_11315,N_8406);
or U12330 (N_12330,N_8631,N_9823);
nor U12331 (N_12331,N_6945,N_8817);
nand U12332 (N_12332,N_10783,N_11465);
nor U12333 (N_12333,N_7703,N_8621);
or U12334 (N_12334,N_6807,N_7264);
or U12335 (N_12335,N_10757,N_11860);
xor U12336 (N_12336,N_9430,N_7361);
or U12337 (N_12337,N_10035,N_6075);
and U12338 (N_12338,N_9159,N_9110);
and U12339 (N_12339,N_9392,N_10194);
xnor U12340 (N_12340,N_11613,N_11822);
or U12341 (N_12341,N_10495,N_11801);
and U12342 (N_12342,N_6899,N_10293);
nor U12343 (N_12343,N_7667,N_11152);
and U12344 (N_12344,N_7855,N_8158);
or U12345 (N_12345,N_11199,N_6603);
nand U12346 (N_12346,N_11979,N_10036);
xnor U12347 (N_12347,N_8824,N_7664);
nor U12348 (N_12348,N_6530,N_9254);
nor U12349 (N_12349,N_11085,N_7773);
xor U12350 (N_12350,N_6753,N_8015);
or U12351 (N_12351,N_11002,N_11654);
or U12352 (N_12352,N_9186,N_7592);
or U12353 (N_12353,N_10340,N_9610);
nor U12354 (N_12354,N_6064,N_6380);
and U12355 (N_12355,N_10368,N_9949);
xnor U12356 (N_12356,N_6600,N_10480);
and U12357 (N_12357,N_10323,N_6943);
nand U12358 (N_12358,N_7754,N_9425);
and U12359 (N_12359,N_9022,N_7543);
and U12360 (N_12360,N_6611,N_7033);
or U12361 (N_12361,N_9657,N_6369);
nor U12362 (N_12362,N_10414,N_11173);
and U12363 (N_12363,N_7274,N_8139);
xor U12364 (N_12364,N_9360,N_7170);
or U12365 (N_12365,N_10673,N_7833);
and U12366 (N_12366,N_9776,N_8671);
or U12367 (N_12367,N_10476,N_6202);
and U12368 (N_12368,N_7625,N_7849);
xor U12369 (N_12369,N_10786,N_11714);
and U12370 (N_12370,N_6971,N_10512);
xnor U12371 (N_12371,N_11740,N_7011);
xor U12372 (N_12372,N_9352,N_11586);
xnor U12373 (N_12373,N_9777,N_6449);
and U12374 (N_12374,N_11696,N_7468);
or U12375 (N_12375,N_9247,N_9063);
xnor U12376 (N_12376,N_10349,N_6900);
nor U12377 (N_12377,N_8593,N_8039);
or U12378 (N_12378,N_8518,N_11157);
or U12379 (N_12379,N_6089,N_10867);
or U12380 (N_12380,N_10047,N_6440);
xor U12381 (N_12381,N_7931,N_6174);
nor U12382 (N_12382,N_11345,N_9363);
nand U12383 (N_12383,N_8377,N_6199);
nand U12384 (N_12384,N_11382,N_6623);
or U12385 (N_12385,N_6850,N_9215);
xor U12386 (N_12386,N_10078,N_8235);
xnor U12387 (N_12387,N_6364,N_7603);
xor U12388 (N_12388,N_9598,N_8946);
nor U12389 (N_12389,N_7802,N_11073);
and U12390 (N_12390,N_9734,N_6913);
nor U12391 (N_12391,N_7972,N_9790);
or U12392 (N_12392,N_7208,N_11473);
or U12393 (N_12393,N_9398,N_11950);
nand U12394 (N_12394,N_10390,N_11655);
xnor U12395 (N_12395,N_10659,N_11156);
nand U12396 (N_12396,N_8868,N_8016);
nor U12397 (N_12397,N_7797,N_10588);
xor U12398 (N_12398,N_7089,N_6861);
nor U12399 (N_12399,N_7014,N_7259);
or U12400 (N_12400,N_7661,N_7340);
xnor U12401 (N_12401,N_6978,N_10720);
and U12402 (N_12402,N_11312,N_11431);
and U12403 (N_12403,N_9129,N_6305);
and U12404 (N_12404,N_9082,N_8233);
nor U12405 (N_12405,N_8402,N_7389);
xnor U12406 (N_12406,N_9162,N_11200);
nor U12407 (N_12407,N_10981,N_11572);
or U12408 (N_12408,N_11298,N_9140);
or U12409 (N_12409,N_10679,N_9765);
nor U12410 (N_12410,N_6690,N_7983);
nor U12411 (N_12411,N_8499,N_6008);
and U12412 (N_12412,N_10491,N_6249);
nand U12413 (N_12413,N_11020,N_9157);
nor U12414 (N_12414,N_6426,N_8660);
nand U12415 (N_12415,N_10568,N_6470);
or U12416 (N_12416,N_6028,N_7692);
nor U12417 (N_12417,N_7535,N_11617);
and U12418 (N_12418,N_6330,N_9820);
nand U12419 (N_12419,N_6859,N_9477);
or U12420 (N_12420,N_7190,N_9555);
xnor U12421 (N_12421,N_6010,N_6655);
nand U12422 (N_12422,N_6912,N_9974);
nor U12423 (N_12423,N_6281,N_10807);
nor U12424 (N_12424,N_8143,N_10167);
nand U12425 (N_12425,N_7860,N_8906);
or U12426 (N_12426,N_11804,N_10494);
and U12427 (N_12427,N_9650,N_8069);
nor U12428 (N_12428,N_10277,N_10019);
nand U12429 (N_12429,N_11144,N_8330);
and U12430 (N_12430,N_10858,N_7498);
nand U12431 (N_12431,N_6287,N_11576);
and U12432 (N_12432,N_10703,N_9550);
or U12433 (N_12433,N_8208,N_10393);
or U12434 (N_12434,N_10973,N_8722);
nand U12435 (N_12435,N_7753,N_7686);
or U12436 (N_12436,N_7729,N_10517);
and U12437 (N_12437,N_7957,N_6975);
nor U12438 (N_12438,N_6389,N_6497);
and U12439 (N_12439,N_10394,N_7638);
xor U12440 (N_12440,N_8356,N_8800);
nand U12441 (N_12441,N_6989,N_7335);
xor U12442 (N_12442,N_7146,N_6944);
nand U12443 (N_12443,N_10501,N_8101);
nor U12444 (N_12444,N_9700,N_11251);
nor U12445 (N_12445,N_6034,N_9080);
or U12446 (N_12446,N_8653,N_9816);
nor U12447 (N_12447,N_7008,N_9576);
and U12448 (N_12448,N_10879,N_6378);
xnor U12449 (N_12449,N_6545,N_6165);
nor U12450 (N_12450,N_9703,N_9539);
and U12451 (N_12451,N_10725,N_9542);
nor U12452 (N_12452,N_8424,N_8765);
xnor U12453 (N_12453,N_10626,N_6867);
or U12454 (N_12454,N_7096,N_7036);
nor U12455 (N_12455,N_8147,N_6357);
or U12456 (N_12456,N_11027,N_9711);
or U12457 (N_12457,N_6896,N_7790);
or U12458 (N_12458,N_11006,N_10881);
and U12459 (N_12459,N_10499,N_11410);
and U12460 (N_12460,N_8752,N_6143);
or U12461 (N_12461,N_7891,N_6013);
and U12462 (N_12462,N_10746,N_8172);
nand U12463 (N_12463,N_9983,N_6769);
nor U12464 (N_12464,N_7735,N_7741);
or U12465 (N_12465,N_10887,N_7293);
nand U12466 (N_12466,N_10221,N_10401);
nor U12467 (N_12467,N_8565,N_10197);
or U12468 (N_12468,N_8129,N_8263);
xor U12469 (N_12469,N_10133,N_9224);
and U12470 (N_12470,N_10468,N_8002);
or U12471 (N_12471,N_6890,N_6940);
xnor U12472 (N_12472,N_6955,N_7912);
nand U12473 (N_12473,N_11596,N_10219);
nor U12474 (N_12474,N_7807,N_8663);
nand U12475 (N_12475,N_9072,N_10502);
nor U12476 (N_12476,N_8173,N_6779);
nand U12477 (N_12477,N_10178,N_11356);
and U12478 (N_12478,N_7292,N_7301);
xnor U12479 (N_12479,N_8103,N_10034);
xnor U12480 (N_12480,N_6889,N_11227);
or U12481 (N_12481,N_11543,N_6063);
xor U12482 (N_12482,N_11777,N_6042);
nor U12483 (N_12483,N_9758,N_11805);
and U12484 (N_12484,N_11841,N_8157);
or U12485 (N_12485,N_11848,N_7333);
xnor U12486 (N_12486,N_10860,N_10151);
and U12487 (N_12487,N_9901,N_8079);
nand U12488 (N_12488,N_10710,N_11548);
and U12489 (N_12489,N_9219,N_8501);
and U12490 (N_12490,N_8454,N_7531);
or U12491 (N_12491,N_9915,N_8754);
nor U12492 (N_12492,N_11198,N_7330);
and U12493 (N_12493,N_8183,N_7558);
nor U12494 (N_12494,N_6962,N_8276);
or U12495 (N_12495,N_6594,N_7793);
and U12496 (N_12496,N_10299,N_8118);
xor U12497 (N_12497,N_8367,N_10594);
or U12498 (N_12498,N_6309,N_7637);
or U12499 (N_12499,N_7079,N_11840);
nor U12500 (N_12500,N_6083,N_10474);
xor U12501 (N_12501,N_11282,N_11374);
and U12502 (N_12502,N_9787,N_6260);
or U12503 (N_12503,N_11398,N_8827);
xnor U12504 (N_12504,N_10906,N_10633);
nand U12505 (N_12505,N_7989,N_9936);
nor U12506 (N_12506,N_9438,N_6901);
or U12507 (N_12507,N_7818,N_6154);
nor U12508 (N_12508,N_6711,N_9632);
or U12509 (N_12509,N_8520,N_10017);
xnor U12510 (N_12510,N_11717,N_8884);
xor U12511 (N_12511,N_7354,N_11700);
nor U12512 (N_12512,N_9172,N_7392);
and U12513 (N_12513,N_7572,N_7239);
xnor U12514 (N_12514,N_11271,N_9408);
nor U12515 (N_12515,N_11880,N_11624);
and U12516 (N_12516,N_6670,N_10539);
xnor U12517 (N_12517,N_6300,N_10645);
nor U12518 (N_12518,N_10630,N_11769);
or U12519 (N_12519,N_9445,N_8783);
and U12520 (N_12520,N_6514,N_7076);
and U12521 (N_12521,N_10007,N_7888);
xor U12522 (N_12522,N_8110,N_6247);
nand U12523 (N_12523,N_7547,N_11977);
nor U12524 (N_12524,N_8325,N_9313);
xnor U12525 (N_12525,N_8241,N_10298);
and U12526 (N_12526,N_10258,N_10942);
nand U12527 (N_12527,N_6323,N_8323);
xnor U12528 (N_12528,N_6788,N_6475);
and U12529 (N_12529,N_9132,N_11888);
and U12530 (N_12530,N_9149,N_11357);
or U12531 (N_12531,N_9309,N_8994);
nor U12532 (N_12532,N_11628,N_10430);
nor U12533 (N_12533,N_7697,N_11373);
nand U12534 (N_12534,N_9984,N_6351);
or U12535 (N_12535,N_11188,N_8659);
nand U12536 (N_12536,N_6408,N_11623);
or U12537 (N_12537,N_10791,N_11699);
or U12538 (N_12538,N_9767,N_11467);
nand U12539 (N_12539,N_11580,N_9583);
nor U12540 (N_12540,N_6181,N_6446);
nor U12541 (N_12541,N_9684,N_10273);
nand U12542 (N_12542,N_9326,N_10598);
nor U12543 (N_12543,N_9568,N_10609);
or U12544 (N_12544,N_11122,N_7314);
nand U12545 (N_12545,N_9001,N_10914);
xor U12546 (N_12546,N_9712,N_10242);
nand U12547 (N_12547,N_7077,N_10387);
or U12548 (N_12548,N_8967,N_11367);
or U12549 (N_12549,N_6677,N_6976);
and U12550 (N_12550,N_9316,N_9713);
nand U12551 (N_12551,N_7345,N_9541);
nand U12552 (N_12552,N_10962,N_7737);
nor U12553 (N_12553,N_6586,N_8622);
and U12554 (N_12554,N_7479,N_6539);
or U12555 (N_12555,N_10863,N_6385);
nor U12556 (N_12556,N_9039,N_8410);
or U12557 (N_12557,N_6895,N_6317);
or U12558 (N_12558,N_6136,N_7792);
nor U12559 (N_12559,N_6011,N_8336);
nor U12560 (N_12560,N_7007,N_8541);
and U12561 (N_12561,N_10166,N_6570);
nand U12562 (N_12562,N_10081,N_9204);
nand U12563 (N_12563,N_8888,N_8384);
nor U12564 (N_12564,N_7811,N_6751);
or U12565 (N_12565,N_7632,N_11587);
nand U12566 (N_12566,N_8435,N_8575);
xor U12567 (N_12567,N_11897,N_11308);
or U12568 (N_12568,N_6984,N_10770);
xor U12569 (N_12569,N_8873,N_10040);
xor U12570 (N_12570,N_10955,N_6922);
nand U12571 (N_12571,N_11986,N_7404);
and U12572 (N_12572,N_11616,N_11541);
xnor U12573 (N_12573,N_7777,N_6014);
nor U12574 (N_12574,N_10472,N_8550);
or U12575 (N_12575,N_9947,N_9060);
xor U12576 (N_12576,N_9836,N_9201);
xor U12577 (N_12577,N_7102,N_11183);
xnor U12578 (N_12578,N_10039,N_9458);
and U12579 (N_12579,N_11695,N_11337);
and U12580 (N_12580,N_9692,N_10489);
or U12581 (N_12581,N_9556,N_6732);
and U12582 (N_12582,N_6285,N_8011);
or U12583 (N_12583,N_6142,N_10664);
and U12584 (N_12584,N_6969,N_10477);
and U12585 (N_12585,N_6452,N_11707);
xor U12586 (N_12586,N_11488,N_10080);
or U12587 (N_12587,N_10829,N_9376);
nor U12588 (N_12588,N_10778,N_7004);
xnor U12589 (N_12589,N_10919,N_10100);
nand U12590 (N_12590,N_10274,N_11035);
and U12591 (N_12591,N_8371,N_8812);
nand U12592 (N_12592,N_10849,N_8952);
xnor U12593 (N_12593,N_10079,N_10843);
xor U12594 (N_12594,N_6529,N_6637);
nand U12595 (N_12595,N_6167,N_9011);
nor U12596 (N_12596,N_7615,N_7319);
nor U12597 (N_12597,N_7295,N_8441);
xnor U12598 (N_12598,N_10953,N_7240);
nand U12599 (N_12599,N_9148,N_8525);
nor U12600 (N_12600,N_8672,N_8629);
or U12601 (N_12601,N_7764,N_6608);
xnor U12602 (N_12602,N_8818,N_7456);
nand U12603 (N_12603,N_10979,N_7039);
xor U12604 (N_12604,N_7537,N_6656);
xor U12605 (N_12605,N_7907,N_8886);
and U12606 (N_12606,N_9118,N_6782);
nor U12607 (N_12607,N_11487,N_7971);
and U12608 (N_12608,N_8860,N_10893);
xnor U12609 (N_12609,N_8981,N_7937);
or U12610 (N_12610,N_11956,N_6412);
nor U12611 (N_12611,N_7508,N_10627);
xnor U12612 (N_12612,N_11791,N_10098);
and U12613 (N_12613,N_9675,N_11225);
or U12614 (N_12614,N_11918,N_6473);
nand U12615 (N_12615,N_7328,N_8379);
and U12616 (N_12616,N_6644,N_7542);
nor U12617 (N_12617,N_11112,N_7020);
xnor U12618 (N_12618,N_9460,N_8030);
and U12619 (N_12619,N_10260,N_8100);
or U12620 (N_12620,N_10714,N_9035);
xor U12621 (N_12621,N_11049,N_8460);
xnor U12622 (N_12622,N_7412,N_6994);
or U12623 (N_12623,N_9898,N_7715);
nand U12624 (N_12624,N_11540,N_7821);
nand U12625 (N_12625,N_9604,N_8625);
nor U12626 (N_12626,N_11877,N_9340);
nor U12627 (N_12627,N_10024,N_6184);
nor U12628 (N_12628,N_9847,N_7371);
nand U12629 (N_12629,N_6721,N_9702);
and U12630 (N_12630,N_7082,N_8128);
and U12631 (N_12631,N_11106,N_6604);
nor U12632 (N_12632,N_8362,N_6610);
nor U12633 (N_12633,N_9569,N_11456);
xor U12634 (N_12634,N_6092,N_7564);
or U12635 (N_12635,N_11709,N_9292);
nor U12636 (N_12636,N_9305,N_8557);
xor U12637 (N_12637,N_9833,N_10526);
and U12638 (N_12638,N_7129,N_10190);
xor U12639 (N_12639,N_6563,N_8154);
or U12640 (N_12640,N_11800,N_8757);
nor U12641 (N_12641,N_9807,N_10030);
xor U12642 (N_12642,N_9023,N_7222);
nor U12643 (N_12643,N_10381,N_11703);
or U12644 (N_12644,N_7746,N_8521);
or U12645 (N_12645,N_11926,N_9066);
nor U12646 (N_12646,N_11187,N_6667);
nor U12647 (N_12647,N_6474,N_6502);
nor U12648 (N_12648,N_7065,N_6645);
nor U12649 (N_12649,N_8412,N_10889);
or U12650 (N_12650,N_11990,N_10083);
or U12651 (N_12651,N_11121,N_10965);
and U12652 (N_12652,N_6219,N_11266);
or U12653 (N_12653,N_7298,N_9031);
and U12654 (N_12654,N_6728,N_6239);
or U12655 (N_12655,N_10682,N_11326);
xor U12656 (N_12656,N_9012,N_9903);
or U12657 (N_12657,N_6607,N_9818);
xnor U12658 (N_12658,N_9642,N_10202);
nand U12659 (N_12659,N_11426,N_10985);
xor U12660 (N_12660,N_6734,N_8347);
and U12661 (N_12661,N_6115,N_6161);
or U12662 (N_12662,N_7488,N_9126);
nand U12663 (N_12663,N_10996,N_11578);
nor U12664 (N_12664,N_11181,N_9049);
xnor U12665 (N_12665,N_11782,N_9589);
or U12666 (N_12666,N_8474,N_6275);
nor U12667 (N_12667,N_10989,N_8993);
nand U12668 (N_12668,N_8641,N_6518);
and U12669 (N_12669,N_9307,N_9117);
nor U12670 (N_12670,N_11406,N_9770);
or U12671 (N_12671,N_9473,N_11834);
nor U12672 (N_12672,N_10076,N_6468);
and U12673 (N_12673,N_11203,N_10885);
or U12674 (N_12674,N_9164,N_10593);
nor U12675 (N_12675,N_8741,N_6370);
nand U12676 (N_12676,N_9773,N_8632);
nand U12677 (N_12677,N_7944,N_10307);
and U12678 (N_12678,N_8311,N_6045);
nand U12679 (N_12679,N_6557,N_7215);
or U12680 (N_12680,N_7590,N_6477);
xor U12681 (N_12681,N_11967,N_11484);
and U12682 (N_12682,N_9452,N_11847);
or U12683 (N_12683,N_10158,N_11638);
and U12684 (N_12684,N_10692,N_10743);
and U12685 (N_12685,N_11111,N_8856);
nand U12686 (N_12686,N_8887,N_8801);
xnor U12687 (N_12687,N_9755,N_8995);
and U12688 (N_12688,N_10043,N_11531);
nand U12689 (N_12689,N_8181,N_9333);
or U12690 (N_12690,N_7183,N_8180);
or U12691 (N_12691,N_10505,N_11909);
nand U12692 (N_12692,N_8217,N_6803);
xnor U12693 (N_12693,N_8054,N_11513);
or U12694 (N_12694,N_9211,N_8682);
nor U12695 (N_12695,N_6982,N_6335);
xnor U12696 (N_12696,N_6855,N_11391);
or U12697 (N_12697,N_6097,N_6559);
and U12698 (N_12698,N_6934,N_8020);
and U12699 (N_12699,N_7709,N_11863);
xnor U12700 (N_12700,N_7569,N_7956);
nand U12701 (N_12701,N_11884,N_6443);
nor U12702 (N_12702,N_8904,N_10113);
nor U12703 (N_12703,N_8588,N_10101);
nor U12704 (N_12704,N_9935,N_10396);
and U12705 (N_12705,N_10612,N_7496);
and U12706 (N_12706,N_7484,N_10315);
or U12707 (N_12707,N_7329,N_10600);
nand U12708 (N_12708,N_9361,N_11423);
xor U12709 (N_12709,N_10607,N_7012);
and U12710 (N_12710,N_8098,N_7154);
or U12711 (N_12711,N_11450,N_8651);
or U12712 (N_12712,N_7762,N_11723);
nor U12713 (N_12713,N_10693,N_10423);
nand U12714 (N_12714,N_9304,N_7866);
nor U12715 (N_12715,N_10852,N_11973);
and U12716 (N_12716,N_8078,N_11437);
and U12717 (N_12717,N_11432,N_7825);
nand U12718 (N_12718,N_7503,N_10504);
nor U12719 (N_12719,N_6596,N_9611);
or U12720 (N_12720,N_7669,N_7370);
nor U12721 (N_12721,N_9044,N_9216);
nand U12722 (N_12722,N_11016,N_8116);
or U12723 (N_12723,N_11671,N_6817);
xor U12724 (N_12724,N_10324,N_8595);
xnor U12725 (N_12725,N_9607,N_11983);
and U12726 (N_12726,N_10138,N_11108);
or U12727 (N_12727,N_6523,N_11132);
and U12728 (N_12728,N_10126,N_10754);
nor U12729 (N_12729,N_7679,N_10291);
or U12730 (N_12730,N_11577,N_9592);
or U12731 (N_12731,N_9557,N_11037);
and U12732 (N_12732,N_8875,N_10615);
nor U12733 (N_12733,N_7367,N_7628);
xnor U12734 (N_12734,N_9980,N_8996);
nand U12735 (N_12735,N_11447,N_6634);
nor U12736 (N_12736,N_8451,N_8568);
or U12737 (N_12737,N_10579,N_11238);
nand U12738 (N_12738,N_11311,N_8594);
nor U12739 (N_12739,N_10992,N_10253);
xor U12740 (N_12740,N_9706,N_10241);
nor U12741 (N_12741,N_10065,N_9439);
xor U12742 (N_12742,N_10911,N_11267);
and U12743 (N_12743,N_8192,N_7396);
xor U12744 (N_12744,N_8636,N_6909);
xnor U12745 (N_12745,N_8104,N_6992);
xor U12746 (N_12746,N_7995,N_8545);
or U12747 (N_12747,N_9436,N_10425);
xor U12748 (N_12748,N_9059,N_11833);
xor U12749 (N_12749,N_7022,N_9636);
nor U12750 (N_12750,N_6935,N_7251);
xnor U12751 (N_12751,N_6463,N_7271);
or U12752 (N_12752,N_8164,N_10475);
nand U12753 (N_12753,N_8177,N_10189);
xor U12754 (N_12754,N_11588,N_7439);
nand U12755 (N_12755,N_10137,N_8746);
or U12756 (N_12756,N_7597,N_10964);
xnor U12757 (N_12757,N_6560,N_9026);
nand U12758 (N_12758,N_8487,N_10343);
nand U12759 (N_12759,N_11439,N_9639);
xor U12760 (N_12760,N_8087,N_6696);
or U12761 (N_12761,N_11900,N_7813);
nor U12762 (N_12762,N_6018,N_11289);
or U12763 (N_12763,N_7052,N_7581);
nor U12764 (N_12764,N_10424,N_11309);
nor U12765 (N_12765,N_10750,N_8339);
xnor U12766 (N_12766,N_11658,N_9174);
xor U12767 (N_12767,N_11537,N_10782);
nand U12768 (N_12768,N_9385,N_8140);
nor U12769 (N_12769,N_7868,N_7967);
and U12770 (N_12770,N_6758,N_8957);
and U12771 (N_12771,N_8370,N_9151);
nor U12772 (N_12772,N_11141,N_11611);
xor U12773 (N_12773,N_11215,N_11745);
xnor U12774 (N_12774,N_8971,N_11734);
and U12775 (N_12775,N_7296,N_9725);
nand U12776 (N_12776,N_9450,N_10135);
or U12777 (N_12777,N_8244,N_9813);
and U12778 (N_12778,N_8025,N_11395);
nor U12779 (N_12779,N_11568,N_8574);
or U12780 (N_12780,N_7996,N_6286);
nand U12781 (N_12781,N_10518,N_8882);
nor U12782 (N_12782,N_9420,N_7768);
or U12783 (N_12783,N_11768,N_8207);
nor U12784 (N_12784,N_10198,N_6196);
xor U12785 (N_12785,N_11448,N_11242);
nor U12786 (N_12786,N_6495,N_8792);
xor U12787 (N_12787,N_8381,N_6486);
or U12788 (N_12788,N_6375,N_7050);
nor U12789 (N_12789,N_10186,N_10794);
xnor U12790 (N_12790,N_11861,N_7152);
or U12791 (N_12791,N_10136,N_10191);
or U12792 (N_12792,N_7565,N_8346);
nand U12793 (N_12793,N_11732,N_6384);
nor U12794 (N_12794,N_8770,N_9619);
xor U12795 (N_12795,N_10199,N_10521);
nor U12796 (N_12796,N_7261,N_8267);
xor U12797 (N_12797,N_8427,N_6892);
and U12798 (N_12798,N_9908,N_8899);
nor U12799 (N_12799,N_6521,N_6977);
nor U12800 (N_12800,N_9470,N_11408);
xor U12801 (N_12801,N_11276,N_7918);
and U12802 (N_12802,N_9617,N_8259);
or U12803 (N_12803,N_10559,N_6481);
nor U12804 (N_12804,N_6911,N_7483);
nor U12805 (N_12805,N_10531,N_7598);
nand U12806 (N_12806,N_6511,N_9729);
and U12807 (N_12807,N_6027,N_7181);
xnor U12808 (N_12808,N_7209,N_7936);
xnor U12809 (N_12809,N_6540,N_7689);
and U12810 (N_12810,N_9691,N_9737);
nor U12811 (N_12811,N_6748,N_8935);
nand U12812 (N_12812,N_11402,N_11462);
and U12813 (N_12813,N_8397,N_11615);
xnor U12814 (N_12814,N_8938,N_11891);
xor U12815 (N_12815,N_9959,N_10790);
or U12816 (N_12816,N_8500,N_9267);
and U12817 (N_12817,N_6297,N_10356);
nand U12818 (N_12818,N_8619,N_8776);
and U12819 (N_12819,N_11305,N_6537);
and U12820 (N_12820,N_7881,N_6342);
or U12821 (N_12821,N_8394,N_10634);
nand U12822 (N_12822,N_6501,N_6503);
or U12823 (N_12823,N_6499,N_9916);
xor U12824 (N_12824,N_8943,N_6821);
xor U12825 (N_12825,N_7749,N_11741);
or U12826 (N_12826,N_6081,N_11363);
xor U12827 (N_12827,N_7794,N_7433);
nor U12828 (N_12828,N_10802,N_11916);
and U12829 (N_12829,N_7595,N_7823);
and U12830 (N_12830,N_11190,N_8125);
xor U12831 (N_12831,N_9894,N_7898);
or U12832 (N_12832,N_7681,N_6580);
nor U12833 (N_12833,N_9276,N_11806);
nand U12834 (N_12834,N_8167,N_8637);
or U12835 (N_12835,N_6227,N_8053);
nand U12836 (N_12836,N_6517,N_10998);
and U12837 (N_12837,N_7149,N_9618);
nor U12838 (N_12838,N_7524,N_9213);
nand U12839 (N_12839,N_10900,N_6767);
xor U12840 (N_12840,N_6749,N_11851);
and U12841 (N_12841,N_9956,N_11667);
and U12842 (N_12842,N_8563,N_6664);
and U12843 (N_12843,N_6928,N_10051);
xor U12844 (N_12844,N_6811,N_7094);
xor U12845 (N_12845,N_6612,N_7236);
or U12846 (N_12846,N_7586,N_6428);
nor U12847 (N_12847,N_6050,N_9130);
xor U12848 (N_12848,N_9206,N_9571);
nand U12849 (N_12849,N_10589,N_11704);
nor U12850 (N_12850,N_8831,N_7364);
xnor U12851 (N_12851,N_9997,N_10355);
nand U12852 (N_12852,N_9528,N_10516);
and U12853 (N_12853,N_6114,N_9490);
nor U12854 (N_12854,N_11249,N_7475);
nor U12855 (N_12855,N_6025,N_7842);
nor U12856 (N_12856,N_9968,N_7107);
xor U12857 (N_12857,N_6411,N_11375);
or U12858 (N_12858,N_11943,N_8482);
xnor U12859 (N_12859,N_7783,N_11781);
nand U12860 (N_12860,N_11963,N_6109);
and U12861 (N_12861,N_7563,N_6450);
and U12862 (N_12862,N_10972,N_10608);
or U12863 (N_12863,N_9739,N_7245);
or U12864 (N_12864,N_6532,N_9497);
nor U12865 (N_12865,N_7892,N_10447);
or U12866 (N_12866,N_11184,N_11966);
or U12867 (N_12867,N_11303,N_10577);
or U12868 (N_12868,N_6813,N_6265);
nor U12869 (N_12869,N_7486,N_6809);
and U12870 (N_12870,N_9501,N_10395);
or U12871 (N_12871,N_9355,N_11211);
xor U12872 (N_12872,N_11131,N_8999);
nor U12873 (N_12873,N_8790,N_11631);
nor U12874 (N_12874,N_8534,N_8303);
and U12875 (N_12875,N_10551,N_10375);
nor U12876 (N_12876,N_7272,N_9527);
nand U12877 (N_12877,N_7653,N_9085);
nand U12878 (N_12878,N_6691,N_9056);
xnor U12879 (N_12879,N_6538,N_11550);
xor U12880 (N_12880,N_8490,N_9900);
nand U12881 (N_12881,N_7594,N_6512);
nor U12882 (N_12882,N_6447,N_10938);
or U12883 (N_12883,N_7268,N_7831);
xnor U12884 (N_12884,N_7789,N_11542);
or U12885 (N_12885,N_11475,N_10206);
nand U12886 (N_12886,N_7526,N_8043);
nor U12887 (N_12887,N_11729,N_7702);
or U12888 (N_12888,N_11403,N_11413);
xnor U12889 (N_12889,N_9886,N_8341);
xor U12890 (N_12890,N_7570,N_9768);
or U12891 (N_12891,N_10585,N_7375);
nand U12892 (N_12892,N_7994,N_7723);
and U12893 (N_12893,N_9522,N_11372);
xor U12894 (N_12894,N_8353,N_11069);
xor U12895 (N_12895,N_10809,N_8138);
or U12896 (N_12896,N_6764,N_9143);
or U12897 (N_12897,N_8048,N_7670);
xor U12898 (N_12898,N_7443,N_6431);
or U12899 (N_12899,N_9349,N_6192);
or U12900 (N_12900,N_7316,N_8299);
and U12901 (N_12901,N_7871,N_6920);
or U12902 (N_12902,N_6061,N_7630);
or U12903 (N_12903,N_9888,N_8005);
or U12904 (N_12904,N_11850,N_7286);
or U12905 (N_12905,N_6241,N_10105);
and U12906 (N_12906,N_7203,N_7861);
or U12907 (N_12907,N_8878,N_7463);
and U12908 (N_12908,N_9046,N_9004);
nor U12909 (N_12909,N_10201,N_7657);
nand U12910 (N_12910,N_11331,N_11143);
or U12911 (N_12911,N_7872,N_11429);
and U12912 (N_12912,N_10312,N_9448);
and U12913 (N_12913,N_9249,N_8934);
and U12914 (N_12914,N_8483,N_8200);
nor U12915 (N_12915,N_10292,N_10859);
or U12916 (N_12916,N_11036,N_6582);
nand U12917 (N_12917,N_9641,N_9502);
or U12918 (N_12918,N_10252,N_10509);
nor U12919 (N_12919,N_10846,N_9653);
nor U12920 (N_12920,N_8761,N_6960);
or U12921 (N_12921,N_10884,N_10227);
or U12922 (N_12922,N_7947,N_10091);
and U12923 (N_12923,N_8464,N_8610);
nor U12924 (N_12924,N_9284,N_7756);
xor U12925 (N_12925,N_11814,N_8612);
nand U12926 (N_12926,N_11563,N_9756);
nor U12927 (N_12927,N_7724,N_11254);
and U12928 (N_12928,N_9073,N_11436);
xnor U12929 (N_12929,N_7763,N_9645);
or U12930 (N_12930,N_11958,N_8931);
xor U12931 (N_12931,N_11463,N_8708);
nor U12932 (N_12932,N_9362,N_10811);
nor U12933 (N_12933,N_9432,N_9469);
or U12934 (N_12934,N_7582,N_6633);
nor U12935 (N_12935,N_8067,N_7403);
nand U12936 (N_12936,N_7680,N_7063);
and U12937 (N_12937,N_7257,N_11017);
nand U12938 (N_12938,N_7593,N_9671);
xnor U12939 (N_12939,N_9025,N_8012);
nor U12940 (N_12940,N_11344,N_11163);
nor U12941 (N_12941,N_8165,N_7852);
and U12942 (N_12942,N_9644,N_11174);
xor U12943 (N_12943,N_9381,N_9846);
and U12944 (N_12944,N_7362,N_6217);
xor U12945 (N_12945,N_8745,N_9454);
xor U12946 (N_12946,N_11865,N_9451);
or U12947 (N_12947,N_10968,N_9902);
nand U12948 (N_12948,N_10969,N_6484);
nor U12949 (N_12949,N_6067,N_7055);
and U12950 (N_12950,N_6948,N_9040);
xnor U12951 (N_12951,N_9880,N_10723);
xor U12952 (N_12952,N_8932,N_11358);
nor U12953 (N_12953,N_6328,N_11168);
xnor U12954 (N_12954,N_8349,N_6588);
and U12955 (N_12955,N_10247,N_8519);
and U12956 (N_12956,N_8784,N_8088);
or U12957 (N_12957,N_11307,N_11642);
nand U12958 (N_12958,N_6825,N_11399);
xnor U12959 (N_12959,N_8808,N_8539);
or U12960 (N_12960,N_6043,N_10283);
nor U12961 (N_12961,N_10915,N_10358);
nor U12962 (N_12962,N_9668,N_8359);
nor U12963 (N_12963,N_7650,N_7583);
nor U12964 (N_12964,N_10028,N_7601);
or U12965 (N_12965,N_6074,N_8781);
nor U12966 (N_12966,N_7895,N_10142);
nand U12967 (N_12967,N_11837,N_7265);
and U12968 (N_12968,N_7545,N_11207);
nand U12969 (N_12969,N_6590,N_11775);
nand U12970 (N_12970,N_6647,N_9981);
xor U12971 (N_12971,N_7720,N_11829);
and U12972 (N_12972,N_10032,N_9763);
and U12973 (N_12973,N_7474,N_10012);
nor U12974 (N_12974,N_6671,N_11835);
or U12975 (N_12975,N_9682,N_7199);
or U12976 (N_12976,N_8338,N_11167);
or U12977 (N_12977,N_9913,N_6267);
and U12978 (N_12978,N_9202,N_11932);
or U12979 (N_12979,N_8288,N_7562);
and U12980 (N_12980,N_7473,N_7447);
and U12981 (N_12981,N_10558,N_6552);
nand U12982 (N_12982,N_10507,N_7618);
nor U12983 (N_12983,N_10446,N_10503);
nand U12984 (N_12984,N_6448,N_10183);
nand U12985 (N_12985,N_8219,N_10952);
and U12986 (N_12986,N_6002,N_11644);
nor U12987 (N_12987,N_6877,N_9079);
nand U12988 (N_12988,N_7694,N_8003);
or U12989 (N_12989,N_9733,N_9905);
or U12990 (N_12990,N_9078,N_9567);
nand U12991 (N_12991,N_6107,N_11906);
nor U12992 (N_12992,N_8940,N_7504);
or U12993 (N_12993,N_8467,N_8843);
nor U12994 (N_12994,N_11361,N_11283);
xor U12995 (N_12995,N_10983,N_7144);
xor U12996 (N_12996,N_8803,N_11581);
and U12997 (N_12997,N_11602,N_6496);
nor U12998 (N_12998,N_8420,N_6232);
xnor U12999 (N_12999,N_10756,N_8335);
and U13000 (N_13000,N_8082,N_9390);
nor U13001 (N_13001,N_8391,N_8231);
xnor U13002 (N_13002,N_6250,N_10182);
or U13003 (N_13003,N_11134,N_10618);
nor U13004 (N_13004,N_10872,N_11243);
nand U13005 (N_13005,N_7053,N_11412);
or U13006 (N_13006,N_7385,N_8375);
xor U13007 (N_13007,N_6205,N_8436);
nand U13008 (N_13008,N_9727,N_11039);
nor U13009 (N_13009,N_9591,N_6675);
xor U13010 (N_13010,N_11380,N_6363);
nand U13011 (N_13011,N_7216,N_7085);
nor U13012 (N_13012,N_11813,N_10932);
or U13013 (N_13013,N_6712,N_6410);
nor U13014 (N_13014,N_7016,N_7409);
nand U13015 (N_13015,N_9296,N_11992);
nand U13016 (N_13016,N_11665,N_9456);
and U13017 (N_13017,N_11025,N_8581);
nand U13018 (N_13018,N_7506,N_10445);
nand U13019 (N_13019,N_9421,N_10006);
and U13020 (N_13020,N_8387,N_9237);
nor U13021 (N_13021,N_10428,N_7376);
or U13022 (N_13022,N_10524,N_10031);
nor U13023 (N_13023,N_9834,N_11180);
or U13024 (N_13024,N_7244,N_8056);
and U13025 (N_13025,N_7427,N_10735);
and U13026 (N_13026,N_8527,N_10439);
and U13027 (N_13027,N_9926,N_9859);
nand U13028 (N_13028,N_9280,N_11153);
nor U13029 (N_13029,N_11954,N_9519);
nor U13030 (N_13030,N_7619,N_8425);
and U13031 (N_13031,N_10850,N_8596);
nor U13032 (N_13032,N_8905,N_10054);
nand U13033 (N_13033,N_7755,N_9911);
nand U13034 (N_13034,N_7786,N_7846);
and U13035 (N_13035,N_10672,N_10591);
xor U13036 (N_13036,N_9038,N_9372);
nor U13037 (N_13037,N_9260,N_7378);
or U13038 (N_13038,N_8365,N_7431);
and U13039 (N_13039,N_8212,N_10466);
nand U13040 (N_13040,N_6991,N_11843);
nor U13041 (N_13041,N_9259,N_7683);
nor U13042 (N_13042,N_9397,N_11899);
or U13043 (N_13043,N_7164,N_10805);
or U13044 (N_13044,N_9595,N_10950);
nand U13045 (N_13045,N_8442,N_8038);
and U13046 (N_13046,N_8842,N_10765);
or U13047 (N_13047,N_11871,N_6668);
or U13048 (N_13048,N_10510,N_8062);
nor U13049 (N_13049,N_7174,N_8643);
and U13050 (N_13050,N_9545,N_10530);
and U13051 (N_13051,N_9141,N_6876);
xnor U13052 (N_13052,N_7442,N_9544);
nor U13053 (N_13053,N_6390,N_6078);
nor U13054 (N_13054,N_6766,N_7610);
or U13055 (N_13055,N_6847,N_8348);
and U13056 (N_13056,N_10797,N_9380);
nand U13057 (N_13057,N_11336,N_9909);
xnor U13058 (N_13058,N_7151,N_11064);
nand U13059 (N_13059,N_11425,N_10842);
or U13060 (N_13060,N_9812,N_10929);
nor U13061 (N_13061,N_6153,N_7613);
nor U13062 (N_13062,N_11896,N_8959);
or U13063 (N_13063,N_6930,N_6430);
xor U13064 (N_13064,N_10702,N_7916);
or U13065 (N_13065,N_8239,N_9086);
xnor U13066 (N_13066,N_6407,N_7346);
nor U13067 (N_13067,N_10669,N_10865);
nand U13068 (N_13068,N_8788,N_6291);
xor U13069 (N_13069,N_6701,N_10866);
and U13070 (N_13070,N_11949,N_7903);
nand U13071 (N_13071,N_9518,N_7238);
and U13072 (N_13072,N_9300,N_9358);
xor U13073 (N_13073,N_8681,N_11496);
or U13074 (N_13074,N_11876,N_8662);
nand U13075 (N_13075,N_10109,N_9346);
and U13076 (N_13076,N_8864,N_7381);
xor U13077 (N_13077,N_8870,N_11730);
and U13078 (N_13078,N_7812,N_7476);
nor U13079 (N_13079,N_9640,N_11650);
nand U13080 (N_13080,N_6981,N_8264);
nand U13081 (N_13081,N_8307,N_7270);
or U13082 (N_13082,N_11583,N_10458);
nand U13083 (N_13083,N_9188,N_8236);
nor U13084 (N_13084,N_6093,N_10847);
nand U13085 (N_13085,N_10419,N_11819);
nand U13086 (N_13086,N_6268,N_9020);
nand U13087 (N_13087,N_6972,N_8876);
and U13088 (N_13088,N_11535,N_6257);
xor U13089 (N_13089,N_8190,N_9185);
and U13090 (N_13090,N_7191,N_11117);
xnor U13091 (N_13091,N_6420,N_7242);
and U13092 (N_13092,N_6509,N_11341);
or U13093 (N_13093,N_8285,N_9198);
or U13094 (N_13094,N_10245,N_10734);
nand U13095 (N_13095,N_11030,N_10354);
xnor U13096 (N_13096,N_7675,N_10370);
nor U13097 (N_13097,N_7126,N_9320);
nand U13098 (N_13098,N_8652,N_10225);
nor U13099 (N_13099,N_8854,N_11396);
and U13100 (N_13100,N_8918,N_8505);
or U13101 (N_13101,N_7757,N_6683);
and U13102 (N_13102,N_8249,N_7490);
nor U13103 (N_13103,N_6739,N_7960);
xor U13104 (N_13104,N_6761,N_11685);
or U13105 (N_13105,N_8036,N_6031);
nor U13106 (N_13106,N_7395,N_7250);
or U13107 (N_13107,N_7326,N_10838);
nand U13108 (N_13108,N_7045,N_8640);
xor U13109 (N_13109,N_6658,N_8170);
and U13110 (N_13110,N_10015,N_6519);
nand U13111 (N_13111,N_10406,N_9480);
nand U13112 (N_13112,N_6553,N_6248);
xor U13113 (N_13113,N_7778,N_9096);
and U13114 (N_13114,N_10179,N_6489);
nand U13115 (N_13115,N_10467,N_6128);
nor U13116 (N_13116,N_7260,N_10342);
xnor U13117 (N_13117,N_7269,N_7981);
or U13118 (N_13118,N_9246,N_10434);
and U13119 (N_13119,N_8047,N_10764);
and U13120 (N_13120,N_11675,N_9730);
or U13121 (N_13121,N_8903,N_10341);
nor U13122 (N_13122,N_6113,N_10927);
xnor U13123 (N_13123,N_10671,N_7950);
or U13124 (N_13124,N_11858,N_11495);
xnor U13125 (N_13125,N_10170,N_6225);
nand U13126 (N_13126,N_7997,N_7550);
nand U13127 (N_13127,N_11264,N_10270);
nor U13128 (N_13128,N_11005,N_9115);
or U13129 (N_13129,N_8676,N_6795);
and U13130 (N_13130,N_7186,N_7247);
nor U13131 (N_13131,N_9274,N_6421);
and U13132 (N_13132,N_11603,N_10713);
nand U13133 (N_13133,N_9485,N_9387);
nand U13134 (N_13134,N_6814,N_10337);
xor U13135 (N_13135,N_6254,N_7616);
nor U13136 (N_13136,N_9815,N_6725);
or U13137 (N_13137,N_7782,N_6244);
nand U13138 (N_13138,N_8198,N_10799);
or U13139 (N_13139,N_11000,N_9064);
and U13140 (N_13140,N_6187,N_7974);
nor U13141 (N_13141,N_11133,N_7701);
xor U13142 (N_13142,N_10011,N_9764);
xor U13143 (N_13143,N_11553,N_10211);
and U13144 (N_13144,N_6222,N_10072);
or U13145 (N_13145,N_9867,N_10564);
and U13146 (N_13146,N_9275,N_8006);
nand U13147 (N_13147,N_11984,N_7300);
xor U13148 (N_13148,N_9742,N_10187);
or U13149 (N_13149,N_6298,N_11497);
nand U13150 (N_13150,N_10827,N_9134);
xnor U13151 (N_13151,N_7725,N_9388);
xor U13152 (N_13152,N_7419,N_8008);
xor U13153 (N_13153,N_8924,N_11776);
or U13154 (N_13154,N_11653,N_10532);
nand U13155 (N_13155,N_11659,N_7520);
and U13156 (N_13156,N_6621,N_11061);
nand U13157 (N_13157,N_6223,N_8743);
nand U13158 (N_13158,N_11802,N_9321);
nor U13159 (N_13159,N_11690,N_10934);
nor U13160 (N_13160,N_9648,N_9263);
nor U13161 (N_13161,N_10825,N_9350);
or U13162 (N_13162,N_9622,N_9356);
or U13163 (N_13163,N_6938,N_11995);
or U13164 (N_13164,N_7540,N_6765);
nand U13165 (N_13165,N_10804,N_9444);
and U13166 (N_13166,N_7158,N_6345);
nand U13167 (N_13167,N_6415,N_6973);
nand U13168 (N_13168,N_8493,N_7528);
nand U13169 (N_13169,N_7399,N_7110);
nand U13170 (N_13170,N_10945,N_6916);
or U13171 (N_13171,N_8278,N_8023);
nor U13172 (N_13172,N_9495,N_6672);
and U13173 (N_13173,N_9906,N_7678);
nor U13174 (N_13174,N_10353,N_10534);
nand U13175 (N_13175,N_7284,N_11910);
nor U13176 (N_13176,N_9531,N_11074);
or U13177 (N_13177,N_9018,N_10176);
and U13178 (N_13178,N_6640,N_8570);
xor U13179 (N_13179,N_7212,N_8530);
nor U13180 (N_13180,N_10416,N_11419);
nor U13181 (N_13181,N_7759,N_6599);
and U13182 (N_13182,N_6874,N_8846);
xor U13183 (N_13183,N_6571,N_6735);
or U13184 (N_13184,N_9231,N_9621);
nor U13185 (N_13185,N_10563,N_11409);
nor U13186 (N_13186,N_8569,N_8782);
xor U13187 (N_13187,N_7325,N_11770);
and U13188 (N_13188,N_8041,N_11371);
nand U13189 (N_13189,N_9299,N_8604);
or U13190 (N_13190,N_9088,N_8837);
nand U13191 (N_13191,N_11057,N_7589);
or U13192 (N_13192,N_11816,N_8623);
and U13193 (N_13193,N_6273,N_11757);
or U13194 (N_13194,N_8840,N_7924);
nand U13195 (N_13195,N_6015,N_9116);
or U13196 (N_13196,N_8221,N_10073);
and U13197 (N_13197,N_7938,N_8975);
or U13198 (N_13198,N_11258,N_7809);
nor U13199 (N_13199,N_11680,N_10620);
xnor U13200 (N_13200,N_11044,N_6873);
nand U13201 (N_13201,N_7391,N_9189);
and U13202 (N_13202,N_8306,N_11032);
nand U13203 (N_13203,N_6606,N_10310);
and U13204 (N_13204,N_8626,N_8408);
and U13205 (N_13205,N_11565,N_8881);
nand U13206 (N_13206,N_9757,N_7035);
nor U13207 (N_13207,N_9169,N_11245);
nand U13208 (N_13208,N_9048,N_9584);
and U13209 (N_13209,N_6392,N_10580);
or U13210 (N_13210,N_8091,N_6595);
and U13211 (N_13211,N_10450,N_8828);
nor U13212 (N_13212,N_8021,N_11625);
nand U13213 (N_13213,N_11209,N_8266);
nand U13214 (N_13214,N_9548,N_9335);
xnor U13215 (N_13215,N_7579,N_11512);
nor U13216 (N_13216,N_10845,N_7449);
xnor U13217 (N_13217,N_6398,N_6904);
nand U13218 (N_13218,N_10003,N_6416);
nand U13219 (N_13219,N_11713,N_11324);
or U13220 (N_13220,N_11784,N_7480);
nor U13221 (N_13221,N_6179,N_8992);
xor U13222 (N_13222,N_9106,N_11079);
or U13223 (N_13223,N_7317,N_11737);
xnor U13224 (N_13224,N_9285,N_6339);
xnor U13225 (N_13225,N_7985,N_10059);
and U13226 (N_13226,N_10116,N_9513);
nand U13227 (N_13227,N_11352,N_10788);
or U13228 (N_13228,N_10527,N_8222);
nand U13229 (N_13229,N_7006,N_10666);
or U13230 (N_13230,N_11360,N_7744);
nor U13231 (N_13231,N_10595,N_9269);
nand U13232 (N_13232,N_9402,N_7552);
nand U13233 (N_13233,N_6996,N_11104);
xor U13234 (N_13234,N_7998,N_10709);
or U13235 (N_13235,N_10010,N_8232);
nor U13236 (N_13236,N_7915,N_7629);
nor U13237 (N_13237,N_11601,N_6145);
or U13238 (N_13238,N_11012,N_8806);
and U13239 (N_13239,N_11923,N_9897);
nor U13240 (N_13240,N_7952,N_8510);
nand U13241 (N_13241,N_11210,N_10373);
or U13242 (N_13242,N_11657,N_7175);
nand U13243 (N_13243,N_6047,N_7687);
and U13244 (N_13244,N_10784,N_6936);
and U13245 (N_13245,N_7999,N_11071);
or U13246 (N_13246,N_7017,N_8926);
nand U13247 (N_13247,N_9221,N_6957);
xnor U13248 (N_13248,N_9008,N_11778);
nand U13249 (N_13249,N_10980,N_10088);
nor U13250 (N_13250,N_9654,N_6160);
xor U13251 (N_13251,N_8184,N_10758);
xnor U13252 (N_13252,N_10690,N_7148);
nand U13253 (N_13253,N_7511,N_11894);
nand U13254 (N_13254,N_9484,N_11955);
xor U13255 (N_13255,N_9244,N_9131);
nor U13256 (N_13256,N_8343,N_11129);
or U13257 (N_13257,N_9724,N_11376);
nand U13258 (N_13258,N_7049,N_9051);
and U13259 (N_13259,N_7060,N_11627);
xor U13260 (N_13260,N_7739,N_9178);
nand U13261 (N_13261,N_10171,N_6666);
and U13262 (N_13262,N_9710,N_11904);
xor U13263 (N_13263,N_6006,N_11115);
and U13264 (N_13264,N_11204,N_9245);
and U13265 (N_13265,N_6177,N_7155);
or U13266 (N_13266,N_6565,N_11100);
xor U13267 (N_13267,N_11787,N_9353);
or U13268 (N_13268,N_7252,N_9934);
or U13269 (N_13269,N_6476,N_7707);
nand U13270 (N_13270,N_6950,N_7662);
nor U13271 (N_13271,N_7127,N_6293);
xnor U13272 (N_13272,N_6303,N_9302);
or U13273 (N_13273,N_7121,N_11273);
and U13274 (N_13274,N_10371,N_11539);
nor U13275 (N_13275,N_11493,N_9471);
xnor U13276 (N_13276,N_9013,N_10262);
and U13277 (N_13277,N_6598,N_11094);
nor U13278 (N_13278,N_6587,N_11962);
or U13279 (N_13279,N_6842,N_11148);
and U13280 (N_13280,N_6296,N_8945);
or U13281 (N_13281,N_11123,N_8968);
nor U13282 (N_13282,N_11460,N_9464);
xnor U13283 (N_13283,N_9606,N_9434);
xnor U13284 (N_13284,N_6688,N_8066);
xnor U13285 (N_13285,N_9384,N_6235);
or U13286 (N_13286,N_8188,N_9262);
or U13287 (N_13287,N_10898,N_11961);
xnor U13288 (N_13288,N_6023,N_9599);
nor U13289 (N_13289,N_10792,N_11779);
xor U13290 (N_13290,N_9521,N_6738);
nand U13291 (N_13291,N_6206,N_7324);
xnor U13292 (N_13292,N_8666,N_11738);
nor U13293 (N_13293,N_6777,N_10616);
and U13294 (N_13294,N_8832,N_10569);
nand U13295 (N_13295,N_7432,N_10026);
nor U13296 (N_13296,N_10223,N_8224);
nand U13297 (N_13297,N_11560,N_9938);
nand U13298 (N_13298,N_11960,N_11718);
or U13299 (N_13299,N_9120,N_11991);
xnor U13300 (N_13300,N_9643,N_6533);
xor U13301 (N_13301,N_9067,N_11147);
or U13302 (N_13302,N_6360,N_7519);
nor U13303 (N_13303,N_11774,N_10286);
nor U13304 (N_13304,N_10823,N_9723);
xnor U13305 (N_13305,N_7019,N_7108);
nor U13306 (N_13306,N_9832,N_11785);
nor U13307 (N_13307,N_10652,N_9923);
and U13308 (N_13308,N_11526,N_7732);
nor U13309 (N_13309,N_9406,N_8577);
nor U13310 (N_13310,N_10321,N_8432);
or U13311 (N_13311,N_6694,N_10402);
or U13312 (N_13312,N_7857,N_10279);
and U13313 (N_13313,N_10155,N_9386);
and U13314 (N_13314,N_11166,N_6290);
or U13315 (N_13315,N_7819,N_10005);
xor U13316 (N_13316,N_11633,N_10592);
nand U13317 (N_13317,N_9858,N_7256);
xor U13318 (N_13318,N_7611,N_11218);
nand U13319 (N_13319,N_11832,N_8045);
nand U13320 (N_13320,N_7549,N_10642);
or U13321 (N_13321,N_6458,N_6137);
xnor U13322 (N_13322,N_6365,N_7128);
nor U13323 (N_13323,N_11683,N_9848);
nand U13324 (N_13324,N_6860,N_11942);
nand U13325 (N_13325,N_11815,N_9965);
xnor U13326 (N_13326,N_10899,N_10383);
nor U13327 (N_13327,N_7880,N_7770);
and U13328 (N_13328,N_8611,N_9091);
nor U13329 (N_13329,N_10533,N_6772);
nor U13330 (N_13330,N_7908,N_6004);
or U13331 (N_13331,N_6708,N_10971);
and U13332 (N_13332,N_7536,N_7742);
nand U13333 (N_13333,N_6697,N_6673);
or U13334 (N_13334,N_11951,N_7125);
or U13335 (N_13335,N_11387,N_8373);
xor U13336 (N_13336,N_9850,N_9054);
xnor U13337 (N_13337,N_6990,N_9100);
nand U13338 (N_13338,N_7901,N_7576);
and U13339 (N_13339,N_10288,N_6882);
nor U13340 (N_13340,N_6846,N_8799);
and U13341 (N_13341,N_7758,N_10637);
xor U13342 (N_13342,N_8829,N_10562);
xnor U13343 (N_13343,N_10877,N_10162);
and U13344 (N_13344,N_8491,N_9998);
xor U13345 (N_13345,N_8247,N_11142);
nand U13346 (N_13346,N_7150,N_11158);
or U13347 (N_13347,N_9525,N_6376);
or U13348 (N_13348,N_10422,N_6796);
nor U13349 (N_13349,N_8892,N_7254);
nand U13350 (N_13350,N_8458,N_10878);
and U13351 (N_13351,N_11193,N_8567);
or U13352 (N_13352,N_10075,N_7652);
or U13353 (N_13353,N_8547,N_7041);
or U13354 (N_13354,N_6352,N_8073);
xnor U13355 (N_13355,N_6246,N_8316);
nand U13356 (N_13356,N_7002,N_11314);
nor U13357 (N_13357,N_10099,N_8445);
and U13358 (N_13358,N_7202,N_11585);
and U13359 (N_13359,N_11823,N_10676);
nor U13360 (N_13360,N_9419,N_8131);
nand U13361 (N_13361,N_8055,N_7817);
and U13362 (N_13362,N_7348,N_9218);
nor U13363 (N_13363,N_6849,N_11651);
nor U13364 (N_13364,N_10921,N_7588);
or U13365 (N_13365,N_7939,N_7622);
or U13366 (N_13366,N_10560,N_9862);
or U13367 (N_13367,N_6979,N_10584);
and U13368 (N_13368,N_8413,N_10096);
or U13369 (N_13369,N_7131,N_7043);
xnor U13370 (N_13370,N_10680,N_6781);
nor U13371 (N_13371,N_10694,N_7122);
nand U13372 (N_13372,N_10421,N_11662);
xor U13373 (N_13373,N_8909,N_6213);
nand U13374 (N_13374,N_8642,N_11647);
nor U13375 (N_13375,N_7285,N_7859);
nor U13376 (N_13376,N_11809,N_6409);
nor U13377 (N_13377,N_7262,N_10455);
nor U13378 (N_13378,N_10172,N_9330);
or U13379 (N_13379,N_9345,N_9705);
nand U13380 (N_13380,N_11455,N_6148);
and U13381 (N_13381,N_7426,N_11070);
and U13382 (N_13382,N_9214,N_7422);
or U13383 (N_13383,N_9382,N_7626);
or U13384 (N_13384,N_10111,N_8819);
nand U13385 (N_13385,N_6947,N_7081);
or U13386 (N_13386,N_7897,N_9720);
nor U13387 (N_13387,N_10180,N_10871);
or U13388 (N_13388,N_8630,N_6574);
nor U13389 (N_13389,N_10653,N_8773);
nand U13390 (N_13390,N_9226,N_8973);
nand U13391 (N_13391,N_10648,N_8334);
nor U13392 (N_13392,N_11255,N_9475);
nand U13393 (N_13393,N_6176,N_10093);
and U13394 (N_13394,N_11514,N_11664);
and U13395 (N_13395,N_11464,N_6756);
nand U13396 (N_13396,N_10650,N_7357);
xor U13397 (N_13397,N_8789,N_9907);
and U13398 (N_13398,N_11928,N_8484);
or U13399 (N_13399,N_7111,N_11090);
and U13400 (N_13400,N_7114,N_10121);
and U13401 (N_13401,N_9685,N_11385);
and U13402 (N_13402,N_8976,N_11340);
nor U13403 (N_13403,N_9630,N_11536);
nor U13404 (N_13404,N_10295,N_10933);
or U13405 (N_13405,N_8841,N_6998);
and U13406 (N_13406,N_10057,N_8178);
nor U13407 (N_13407,N_9375,N_9879);
and U13408 (N_13408,N_11476,N_7253);
or U13409 (N_13409,N_7932,N_9695);
or U13410 (N_13410,N_8186,N_7177);
or U13411 (N_13411,N_8822,N_8705);
nand U13412 (N_13412,N_9236,N_11739);
nand U13413 (N_13413,N_10282,N_9753);
and U13414 (N_13414,N_10991,N_11004);
nand U13415 (N_13415,N_9301,N_8823);
and U13416 (N_13416,N_10108,N_8396);
xnor U13417 (N_13417,N_9407,N_7494);
nand U13418 (N_13418,N_6970,N_9166);
nand U13419 (N_13419,N_10038,N_8950);
or U13420 (N_13420,N_9124,N_11875);
and U13421 (N_13421,N_6891,N_8702);
nor U13422 (N_13422,N_8894,N_10651);
nand U13423 (N_13423,N_11466,N_7577);
and U13424 (N_13424,N_7027,N_6299);
xor U13425 (N_13425,N_10719,N_6830);
nor U13426 (N_13426,N_9089,N_6347);
nor U13427 (N_13427,N_7631,N_6820);
and U13428 (N_13428,N_9437,N_7061);
and U13429 (N_13429,N_11593,N_7894);
and U13430 (N_13430,N_9535,N_6049);
and U13431 (N_13431,N_10695,N_11618);
xor U13432 (N_13432,N_11883,N_9062);
and U13433 (N_13433,N_6388,N_11405);
xnor U13434 (N_13434,N_6405,N_10668);
xnor U13435 (N_13435,N_9667,N_10339);
and U13436 (N_13436,N_7492,N_10397);
nand U13437 (N_13437,N_9065,N_9719);
or U13438 (N_13438,N_8814,N_10993);
xor U13439 (N_13439,N_10978,N_9034);
xor U13440 (N_13440,N_9683,N_8573);
nand U13441 (N_13441,N_9996,N_6903);
nor U13442 (N_13442,N_8315,N_9581);
nor U13443 (N_13443,N_8587,N_6535);
xnor U13444 (N_13444,N_7440,N_8912);
or U13445 (N_13445,N_11062,N_8439);
nor U13446 (N_13446,N_9579,N_9991);
or U13447 (N_13447,N_6150,N_7747);
and U13448 (N_13448,N_9422,N_7523);
xnor U13449 (N_13449,N_7198,N_8769);
xor U13450 (N_13450,N_6816,N_8357);
xnor U13451 (N_13451,N_11214,N_11278);
nand U13452 (N_13452,N_8511,N_7600);
nor U13453 (N_13453,N_6082,N_11500);
and U13454 (N_13454,N_7363,N_6952);
and U13455 (N_13455,N_11941,N_11236);
nand U13456 (N_13456,N_10639,N_7168);
or U13457 (N_13457,N_8524,N_10334);
nor U13458 (N_13458,N_6193,N_9664);
nand U13459 (N_13459,N_9081,N_10832);
xor U13460 (N_13460,N_7889,N_10610);
or U13461 (N_13461,N_7446,N_11260);
xor U13462 (N_13462,N_9596,N_11194);
nand U13463 (N_13463,N_7935,N_10145);
xnor U13464 (N_13464,N_7691,N_7042);
and U13465 (N_13465,N_11530,N_11480);
xnor U13466 (N_13466,N_10656,N_9551);
and U13467 (N_13467,N_11938,N_10192);
and U13468 (N_13468,N_8506,N_9101);
xnor U13469 (N_13469,N_8897,N_7837);
nand U13470 (N_13470,N_10732,N_9554);
or U13471 (N_13471,N_10717,N_11138);
or U13472 (N_13472,N_8265,N_7775);
xnor U13473 (N_13473,N_8309,N_10300);
and U13474 (N_13474,N_6368,N_10160);
nand U13475 (N_13475,N_9709,N_7713);
and U13476 (N_13476,N_11175,N_7788);
and U13477 (N_13477,N_8437,N_8366);
nand U13478 (N_13478,N_10049,N_6454);
and U13479 (N_13479,N_10301,N_8522);
and U13480 (N_13480,N_9944,N_6709);
and U13481 (N_13481,N_11219,N_9468);
xnor U13482 (N_13482,N_7145,N_6674);
and U13483 (N_13483,N_9795,N_8578);
and U13484 (N_13484,N_6526,N_9789);
nor U13485 (N_13485,N_8107,N_6939);
or U13486 (N_13486,N_11722,N_7695);
nor U13487 (N_13487,N_9857,N_9687);
and U13488 (N_13488,N_6122,N_11235);
and U13489 (N_13489,N_10331,N_6907);
nand U13490 (N_13490,N_8779,N_6314);
nor U13491 (N_13491,N_11481,N_10861);
nand U13492 (N_13492,N_7966,N_11381);
nand U13493 (N_13493,N_8135,N_10338);
xor U13494 (N_13494,N_9199,N_9306);
nand U13495 (N_13495,N_9537,N_6253);
or U13496 (N_13496,N_7200,N_7970);
nor U13497 (N_13497,N_7275,N_8090);
xnor U13498 (N_13498,N_10114,N_11478);
and U13499 (N_13499,N_7914,N_8209);
and U13500 (N_13500,N_11743,N_10204);
or U13501 (N_13501,N_8889,N_7676);
or U13502 (N_13502,N_10328,N_10724);
and U13503 (N_13503,N_7334,N_7046);
nand U13504 (N_13504,N_11925,N_6125);
nor U13505 (N_13505,N_8228,N_11969);
and U13506 (N_13506,N_7359,N_9602);
nor U13507 (N_13507,N_11113,N_6332);
nand U13508 (N_13508,N_10574,N_7660);
nor U13509 (N_13509,N_8901,N_11501);
or U13510 (N_13510,N_6472,N_9179);
and U13511 (N_13511,N_11607,N_11241);
and U13512 (N_13512,N_10363,N_11534);
or U13513 (N_13513,N_9170,N_9099);
nand U13514 (N_13514,N_10261,N_9878);
nor U13515 (N_13515,N_10322,N_8628);
nand U13516 (N_13516,N_8691,N_9731);
and U13517 (N_13517,N_9158,N_6798);
xnor U13518 (N_13518,N_10599,N_10712);
or U13519 (N_13519,N_10485,N_7373);
xor U13520 (N_13520,N_6198,N_9623);
nand U13521 (N_13521,N_7227,N_9651);
and U13522 (N_13522,N_6775,N_10433);
or U13523 (N_13523,N_9465,N_9594);
nor U13524 (N_13524,N_7685,N_6258);
xor U13525 (N_13525,N_11957,N_11415);
nor U13526 (N_13526,N_7189,N_11490);
nor U13527 (N_13527,N_7904,N_6872);
and U13528 (N_13528,N_8261,N_8849);
nand U13529 (N_13529,N_7507,N_8552);
xnor U13530 (N_13530,N_11978,N_7205);
or U13531 (N_13531,N_9637,N_11879);
or U13532 (N_13532,N_6320,N_6662);
or U13533 (N_13533,N_10597,N_9348);
nand U13534 (N_13534,N_10238,N_6096);
or U13535 (N_13535,N_9726,N_6138);
xor U13536 (N_13536,N_8502,N_11018);
nor U13537 (N_13537,N_10143,N_9885);
or U13538 (N_13538,N_11098,N_7602);
nor U13539 (N_13539,N_9252,N_6718);
xnor U13540 (N_13540,N_11559,N_8735);
nand U13541 (N_13541,N_8923,N_6845);
nand U13542 (N_13542,N_11043,N_9297);
nor U13543 (N_13543,N_6870,N_11673);
and U13544 (N_13544,N_9830,N_8456);
and U13545 (N_13545,N_8202,N_8486);
nand U13546 (N_13546,N_8354,N_11839);
nand U13547 (N_13547,N_6048,N_6805);
or U13548 (N_13548,N_11136,N_9797);
nor U13549 (N_13549,N_7132,N_10269);
and U13550 (N_13550,N_9505,N_11817);
xnor U13551 (N_13551,N_7527,N_9943);
nor U13552 (N_13552,N_8670,N_10768);
nand U13553 (N_13553,N_10271,N_10070);
nor U13554 (N_13554,N_6573,N_10855);
and U13555 (N_13555,N_7380,N_11127);
nor U13556 (N_13556,N_9791,N_6231);
and U13557 (N_13557,N_10959,N_6224);
nor U13558 (N_13558,N_9405,N_7551);
nand U13559 (N_13559,N_7902,N_11296);
nand U13560 (N_13560,N_8274,N_11857);
or U13561 (N_13561,N_6632,N_11034);
or U13562 (N_13562,N_8089,N_8352);
xor U13563 (N_13563,N_9562,N_11852);
nand U13564 (N_13564,N_11140,N_9701);
or U13565 (N_13565,N_8121,N_9960);
and U13566 (N_13566,N_10209,N_11798);
nand U13567 (N_13567,N_8536,N_6432);
nand U13568 (N_13568,N_6919,N_8767);
or U13569 (N_13569,N_10793,N_9207);
nand U13570 (N_13570,N_10294,N_10755);
nand U13571 (N_13571,N_7620,N_11092);
nor U13572 (N_13572,N_6189,N_9656);
and U13573 (N_13573,N_9378,N_9137);
or U13574 (N_13574,N_6478,N_9992);
xor U13575 (N_13575,N_10205,N_8342);
nand U13576 (N_13576,N_11433,N_11663);
xnor U13577 (N_13577,N_9019,N_8785);
xnor U13578 (N_13578,N_10940,N_8279);
nand U13579 (N_13579,N_8983,N_10880);
or U13580 (N_13580,N_7417,N_7659);
nand U13581 (N_13581,N_9290,N_10548);
or U13582 (N_13582,N_10141,N_10493);
and U13583 (N_13583,N_10251,N_8962);
nor U13584 (N_13584,N_11952,N_11384);
or U13585 (N_13585,N_11288,N_8479);
nor U13586 (N_13586,N_11055,N_8956);
or U13587 (N_13587,N_10464,N_7841);
nand U13588 (N_13588,N_6554,N_10737);
nor U13589 (N_13589,N_6361,N_9057);
and U13590 (N_13590,N_11257,N_10125);
and U13591 (N_13591,N_8465,N_6080);
or U13592 (N_13592,N_8291,N_6466);
nand U13593 (N_13593,N_11890,N_6522);
and U13594 (N_13594,N_9107,N_6170);
nor U13595 (N_13595,N_6041,N_6933);
xnor U13596 (N_13596,N_6036,N_10905);
nor U13597 (N_13597,N_7718,N_9676);
xnor U13598 (N_13598,N_10470,N_7500);
and U13599 (N_13599,N_10640,N_8969);
xnor U13600 (N_13600,N_11212,N_6918);
xor U13601 (N_13601,N_8793,N_6654);
or U13602 (N_13602,N_6844,N_10278);
or U13603 (N_13603,N_10944,N_10377);
and U13604 (N_13604,N_7899,N_11971);
nor U13605 (N_13605,N_11126,N_6520);
and U13606 (N_13606,N_8893,N_6505);
xnor U13607 (N_13607,N_10046,N_7780);
nand U13608 (N_13608,N_8022,N_10982);
xnor U13609 (N_13609,N_7803,N_8468);
or U13610 (N_13610,N_11600,N_6436);
or U13611 (N_13611,N_10995,N_6024);
nor U13612 (N_13612,N_8084,N_9842);
and U13613 (N_13613,N_11517,N_8913);
or U13614 (N_13614,N_7986,N_6810);
and U13615 (N_13615,N_9416,N_6487);
and U13616 (N_13616,N_6319,N_10444);
xnor U13617 (N_13617,N_8009,N_11339);
nand U13618 (N_13618,N_6183,N_8478);
nor U13619 (N_13619,N_8916,N_8097);
and U13620 (N_13620,N_6359,N_9433);
nand U13621 (N_13621,N_7080,N_8111);
xor U13622 (N_13622,N_8925,N_9572);
xor U13623 (N_13623,N_9250,N_6577);
or U13624 (N_13624,N_8679,N_9553);
and U13625 (N_13625,N_6066,N_7838);
or U13626 (N_13626,N_6755,N_9045);
nand U13627 (N_13627,N_6967,N_11831);
nor U13628 (N_13628,N_6141,N_7858);
nor U13629 (N_13629,N_8152,N_8166);
nand U13630 (N_13630,N_8740,N_11812);
xor U13631 (N_13631,N_11924,N_8419);
xor U13632 (N_13632,N_6636,N_10685);
nand U13633 (N_13633,N_11903,N_8674);
and U13634 (N_13634,N_9659,N_7103);
and U13635 (N_13635,N_11824,N_9336);
or U13636 (N_13636,N_8858,N_10020);
nor U13637 (N_13637,N_6233,N_7740);
xnor U13638 (N_13638,N_9662,N_8687);
or U13639 (N_13639,N_8251,N_10063);
xnor U13640 (N_13640,N_11259,N_8713);
nand U13641 (N_13641,N_8748,N_9799);
or U13642 (N_13642,N_10976,N_9635);
xnor U13643 (N_13643,N_6801,N_7390);
xor U13644 (N_13644,N_10243,N_6762);
nand U13645 (N_13645,N_6030,N_8654);
and U13646 (N_13646,N_9005,N_6605);
and U13647 (N_13647,N_8509,N_11277);
nor U13648 (N_13648,N_11867,N_11907);
xor U13649 (N_13649,N_10774,N_10961);
and U13650 (N_13650,N_8885,N_8635);
and U13651 (N_13651,N_9958,N_8119);
and U13652 (N_13652,N_8920,N_11454);
and U13653 (N_13653,N_10731,N_8707);
or U13654 (N_13654,N_11697,N_7711);
xor U13655 (N_13655,N_11306,N_11873);
nor U13656 (N_13656,N_9052,N_8446);
nand U13657 (N_13657,N_11046,N_7791);
or U13658 (N_13658,N_8725,N_8826);
and U13659 (N_13659,N_9736,N_11827);
xor U13660 (N_13660,N_7814,N_7054);
nor U13661 (N_13661,N_6480,N_10817);
xor U13662 (N_13662,N_8136,N_9892);
xor U13663 (N_13663,N_9127,N_6129);
nand U13664 (N_13664,N_10500,N_11634);
nor U13665 (N_13665,N_7489,N_11711);
and U13666 (N_13666,N_10741,N_10606);
or U13667 (N_13667,N_8605,N_8755);
nor U13668 (N_13668,N_6602,N_6461);
and U13669 (N_13669,N_9871,N_8382);
or U13670 (N_13670,N_9854,N_7048);
and U13671 (N_13671,N_11728,N_7071);
nor U13672 (N_13672,N_6853,N_10457);
nor U13673 (N_13673,N_9774,N_8977);
nor U13674 (N_13674,N_10697,N_11469);
and U13675 (N_13675,N_6704,N_9851);
nor U13676 (N_13676,N_7124,N_7273);
nand U13677 (N_13677,N_8376,N_10895);
and U13678 (N_13678,N_11511,N_8308);
xor U13679 (N_13679,N_10210,N_10272);
or U13680 (N_13680,N_10762,N_11870);
or U13681 (N_13681,N_8475,N_10281);
xnor U13682 (N_13682,N_11021,N_9050);
xor U13683 (N_13683,N_7058,N_6271);
xnor U13684 (N_13684,N_11453,N_10436);
nand U13685 (N_13685,N_10218,N_7965);
xnor U13686 (N_13686,N_8225,N_7873);
nor U13687 (N_13687,N_8473,N_7413);
nor U13688 (N_13688,N_11649,N_9779);
nand U13689 (N_13689,N_11767,N_10266);
nand U13690 (N_13690,N_8583,N_7187);
xnor U13691 (N_13691,N_6843,N_6163);
nor U13692 (N_13692,N_11327,N_8895);
nor U13693 (N_13693,N_8656,N_9566);
nor U13694 (N_13694,N_8132,N_6457);
nor U13695 (N_13695,N_10986,N_6710);
nand U13696 (N_13696,N_9311,N_7827);
nor U13697 (N_13697,N_6508,N_8063);
nor U13698 (N_13698,N_6423,N_9266);
nand U13699 (N_13699,N_11087,N_7344);
nand U13700 (N_13700,N_6441,N_11993);
nand U13701 (N_13701,N_9910,N_11424);
or U13702 (N_13702,N_7226,N_6130);
or U13703 (N_13703,N_11726,N_10220);
xor U13704 (N_13704,N_9396,N_8685);
or U13705 (N_13705,N_8900,N_7567);
and U13706 (N_13706,N_6961,N_9271);
or U13707 (N_13707,N_11393,N_8815);
or U13708 (N_13708,N_11294,N_6651);
xnor U13709 (N_13709,N_7201,N_10119);
nor U13710 (N_13710,N_9945,N_7448);
nand U13711 (N_13711,N_7255,N_11976);
xor U13712 (N_13712,N_10761,N_6921);
xor U13713 (N_13713,N_11750,N_7787);
xnor U13714 (N_13714,N_7372,N_7384);
nor U13715 (N_13715,N_6100,N_9708);
nand U13716 (N_13716,N_10082,N_10773);
nand U13717 (N_13717,N_8024,N_9479);
or U13718 (N_13718,N_7382,N_8145);
and U13719 (N_13719,N_10264,N_11483);
xnor U13720 (N_13720,N_9273,N_7609);
xor U13721 (N_13721,N_9084,N_11826);
xor U13722 (N_13722,N_9673,N_10813);
nor U13723 (N_13723,N_7141,N_9491);
or U13724 (N_13724,N_10203,N_7047);
nand U13725 (N_13725,N_6055,N_10041);
nand U13726 (N_13726,N_7513,N_9530);
nand U13727 (N_13727,N_9523,N_11854);
nor U13728 (N_13728,N_7748,N_9395);
and U13729 (N_13729,N_9264,N_8095);
nor U13730 (N_13730,N_9793,N_9738);
nand U13731 (N_13731,N_11764,N_11652);
and U13732 (N_13732,N_7964,N_6614);
or U13733 (N_13733,N_8333,N_11010);
and U13734 (N_13734,N_6700,N_10787);
nand U13735 (N_13735,N_6736,N_8113);
xnor U13736 (N_13736,N_7026,N_6556);
nand U13737 (N_13737,N_8665,N_6403);
or U13738 (N_13738,N_8699,N_11047);
xnor U13739 (N_13739,N_11507,N_7922);
xnor U13740 (N_13740,N_9856,N_11746);
or U13741 (N_13741,N_10894,N_9334);
and U13742 (N_13742,N_7350,N_8982);
nor U13743 (N_13743,N_10229,N_9209);
or U13744 (N_13744,N_7185,N_11050);
xnor U13745 (N_13745,N_7233,N_10918);
xnor U13746 (N_13746,N_11786,N_9549);
xor U13747 (N_13747,N_7656,N_7905);
xor U13748 (N_13748,N_10118,N_8206);
xnor U13749 (N_13749,N_7278,N_8874);
nor U13750 (N_13750,N_7156,N_11736);
xnor U13751 (N_13751,N_8673,N_11323);
or U13752 (N_13752,N_7178,N_6354);
and U13753 (N_13753,N_9489,N_6465);
nor U13754 (N_13754,N_11239,N_7835);
and U13755 (N_13755,N_11789,N_8028);
nand U13756 (N_13756,N_9092,N_6338);
nor U13757 (N_13757,N_8857,N_7453);
nor U13758 (N_13758,N_10248,N_7514);
nor U13759 (N_13759,N_8508,N_6714);
or U13760 (N_13760,N_11472,N_8455);
or U13761 (N_13761,N_7287,N_7167);
nor U13762 (N_13762,N_6888,N_10662);
and U13763 (N_13763,N_10235,N_11279);
nand U13764 (N_13764,N_10581,N_7031);
and U13765 (N_13765,N_11246,N_8146);
and U13766 (N_13766,N_11959,N_8700);
xnor U13767 (N_13767,N_9747,N_9194);
and U13768 (N_13768,N_9139,N_6527);
nand U13769 (N_13769,N_11013,N_10496);
nand U13770 (N_13770,N_8319,N_11710);
nor U13771 (N_13771,N_8764,N_6857);
nor U13772 (N_13772,N_8272,N_7091);
xor U13773 (N_13773,N_9242,N_6880);
nor U13774 (N_13774,N_6433,N_8963);
or U13775 (N_13775,N_8650,N_11842);
xor U13776 (N_13776,N_11028,N_10700);
nand U13777 (N_13777,N_10604,N_6663);
and U13778 (N_13778,N_9616,N_6661);
and U13779 (N_13779,N_9918,N_7454);
nand U13780 (N_13780,N_6812,N_11640);
or U13781 (N_13781,N_6724,N_6575);
nand U13782 (N_13782,N_9874,N_7979);
and U13783 (N_13783,N_6393,N_11564);
or U13784 (N_13784,N_10587,N_7634);
and U13785 (N_13785,N_9957,N_6513);
or U13786 (N_13786,N_10106,N_8902);
or U13787 (N_13787,N_9780,N_7959);
nor U13788 (N_13788,N_7266,N_6741);
nand U13789 (N_13789,N_9869,N_10454);
or U13790 (N_13790,N_10359,N_10029);
nor U13791 (N_13791,N_11285,N_9904);
or U13792 (N_13792,N_6164,N_10122);
xor U13793 (N_13793,N_10175,N_6460);
nand U13794 (N_13794,N_9741,N_9977);
or U13795 (N_13795,N_9608,N_9699);
nor U13796 (N_13796,N_6642,N_8238);
and U13797 (N_13797,N_11945,N_8426);
nand U13798 (N_13798,N_7097,N_6333);
nand U13799 (N_13799,N_8980,N_7305);
nor U13800 (N_13800,N_8243,N_11771);
or U13801 (N_13801,N_8344,N_11546);
and U13802 (N_13802,N_6159,N_9409);
and U13803 (N_13803,N_6722,N_7225);
nand U13804 (N_13804,N_10686,N_6684);
or U13805 (N_13805,N_9688,N_6885);
or U13806 (N_13806,N_11849,N_6785);
xnor U13807 (N_13807,N_6665,N_9327);
xor U13808 (N_13808,N_11065,N_9155);
nand U13809 (N_13809,N_11702,N_7539);
nor U13810 (N_13810,N_9090,N_6270);
nand U13811 (N_13811,N_10469,N_7733);
nor U13812 (N_13812,N_11515,N_6827);
nand U13813 (N_13813,N_7393,N_8117);
nor U13814 (N_13814,N_6824,N_9459);
nand U13815 (N_13815,N_7025,N_10806);
xnor U13816 (N_13816,N_9303,N_7418);
nor U13817 (N_13817,N_6325,N_9097);
or U13818 (N_13818,N_7696,N_7668);
or U13819 (N_13819,N_6353,N_10820);
xor U13820 (N_13820,N_10050,N_9014);
and U13821 (N_13821,N_7571,N_10522);
and U13822 (N_13822,N_7320,N_6482);
xnor U13823 (N_13823,N_8572,N_11874);
and U13824 (N_13824,N_9626,N_8257);
or U13825 (N_13825,N_7318,N_8513);
xor U13826 (N_13826,N_6112,N_11561);
nor U13827 (N_13827,N_11040,N_7736);
xnor U13828 (N_13828,N_8802,N_7596);
nor U13829 (N_13829,N_8867,N_9890);
and U13830 (N_13830,N_10718,N_9628);
nand U13831 (N_13831,N_6185,N_10129);
or U13832 (N_13832,N_8201,N_6131);
nand U13833 (N_13833,N_8059,N_8364);
or U13834 (N_13834,N_8948,N_9418);
nand U13835 (N_13835,N_7441,N_9503);
xor U13836 (N_13836,N_10263,N_9197);
and U13837 (N_13837,N_11224,N_10655);
and U13838 (N_13838,N_8205,N_7472);
or U13839 (N_13839,N_11882,N_8727);
or U13840 (N_13840,N_10772,N_9163);
nor U13841 (N_13841,N_11528,N_6717);
nor U13842 (N_13842,N_6639,N_9680);
or U13843 (N_13843,N_6374,N_11821);
nor U13844 (N_13844,N_8489,N_8990);
and U13845 (N_13845,N_9294,N_9253);
nor U13846 (N_13846,N_10107,N_9766);
nand U13847 (N_13847,N_6456,N_10347);
xnor U13848 (N_13848,N_9404,N_6504);
xnor U13849 (N_13849,N_11416,N_9514);
nor U13850 (N_13850,N_8690,N_6914);
nand U13851 (N_13851,N_8942,N_11948);
or U13852 (N_13852,N_11914,N_10000);
xor U13853 (N_13853,N_7856,N_11748);
xnor U13854 (N_13854,N_6609,N_7093);
nor U13855 (N_13855,N_8598,N_9410);
and U13856 (N_13856,N_10831,N_10635);
xnor U13857 (N_13857,N_11701,N_8275);
and U13858 (N_13858,N_10661,N_10362);
xnor U13859 (N_13859,N_11630,N_10990);
and U13860 (N_13860,N_11684,N_7580);
xnor U13861 (N_13861,N_9547,N_7708);
xor U13862 (N_13862,N_8774,N_7878);
and U13863 (N_13863,N_6348,N_10545);
and U13864 (N_13864,N_9561,N_10596);
nor U13865 (N_13865,N_10575,N_7436);
nand U13866 (N_13866,N_6070,N_6837);
nand U13867 (N_13867,N_7138,N_8149);
nor U13868 (N_13868,N_9195,N_9661);
or U13869 (N_13869,N_9229,N_10060);
xor U13870 (N_13870,N_11041,N_9512);
nor U13871 (N_13871,N_6858,N_11101);
nand U13872 (N_13872,N_8137,N_7464);
nand U13873 (N_13873,N_8646,N_8421);
nand U13874 (N_13874,N_10901,N_6774);
xnor U13875 (N_13875,N_10711,N_7688);
nor U13876 (N_13876,N_10351,N_11930);
nand U13877 (N_13877,N_8607,N_9493);
or U13878 (N_13878,N_9819,N_11922);
and U13879 (N_13879,N_9969,N_8083);
xnor U13880 (N_13880,N_11272,N_9895);
and U13881 (N_13881,N_8701,N_9658);
nand U13882 (N_13882,N_7648,N_11619);
nand U13883 (N_13883,N_6778,N_8160);
xor U13884 (N_13884,N_8350,N_11240);
nor U13885 (N_13885,N_9690,N_7117);
and U13886 (N_13886,N_6638,N_10037);
and U13887 (N_13887,N_8648,N_7083);
nand U13888 (N_13888,N_6492,N_6869);
xor U13889 (N_13889,N_7130,N_8517);
and U13890 (N_13890,N_9899,N_10775);
or U13891 (N_13891,N_8960,N_10883);
or U13892 (N_13892,N_8014,N_11220);
and U13893 (N_13893,N_6039,N_8099);
nand U13894 (N_13894,N_11155,N_11525);
or U13895 (N_13895,N_10275,N_7029);
or U13896 (N_13896,N_9932,N_9925);
nor U13897 (N_13897,N_8127,N_9930);
and U13898 (N_13898,N_8027,N_10309);
and U13899 (N_13899,N_11404,N_7331);
or U13900 (N_13900,N_9429,N_6419);
nand U13901 (N_13901,N_6680,N_10018);
and U13902 (N_13902,N_11370,N_10267);
nand U13903 (N_13903,N_8964,N_10960);
nor U13904 (N_13904,N_6699,N_8102);
nand U13905 (N_13905,N_7705,N_8443);
nand U13906 (N_13906,N_10318,N_9190);
and U13907 (N_13907,N_7828,N_6625);
or U13908 (N_13908,N_9873,N_9037);
xnor U13909 (N_13909,N_11461,N_9796);
xnor U13910 (N_13910,N_7693,N_6218);
or U13911 (N_13911,N_10688,N_7068);
or U13912 (N_13912,N_8026,N_9529);
nor U13913 (N_13913,N_10027,N_11159);
and U13914 (N_13914,N_8283,N_10771);
or U13915 (N_13915,N_8998,N_6681);
xor U13916 (N_13916,N_7407,N_9232);
nor U13917 (N_13917,N_10745,N_8533);
nand U13918 (N_13918,N_6017,N_9855);
nor U13919 (N_13919,N_6007,N_11052);
nor U13920 (N_13920,N_7499,N_9119);
or U13921 (N_13921,N_6336,N_11088);
and U13922 (N_13922,N_7779,N_8758);
and U13923 (N_13923,N_7900,N_6056);
or U13924 (N_13924,N_9256,N_9973);
nand U13925 (N_13925,N_6173,N_8071);
and U13926 (N_13926,N_8485,N_6072);
xor U13927 (N_13927,N_7863,N_11566);
and U13928 (N_13928,N_9105,N_6062);
nand U13929 (N_13929,N_9248,N_11947);
or U13930 (N_13930,N_9669,N_6116);
nand U13931 (N_13931,N_8747,N_9286);
nand U13932 (N_13932,N_8415,N_7343);
nand U13933 (N_13933,N_11164,N_10822);
xnor U13934 (N_13934,N_6259,N_11201);
or U13935 (N_13935,N_11316,N_9161);
and U13936 (N_13936,N_11716,N_6040);
xnor U13937 (N_13937,N_9288,N_10482);
nand U13938 (N_13938,N_7289,N_10767);
nand U13939 (N_13939,N_9053,N_10366);
xor U13940 (N_13940,N_8531,N_11390);
xnor U13941 (N_13941,N_11491,N_6255);
nor U13942 (N_13942,N_6848,N_7640);
xor U13943 (N_13943,N_7119,N_7044);
and U13944 (N_13944,N_7890,N_7948);
and U13945 (N_13945,N_10519,N_7032);
or U13946 (N_13946,N_10265,N_7067);
nand U13947 (N_13947,N_6865,N_8007);
nor U13948 (N_13948,N_8401,N_11068);
or U13949 (N_13949,N_8928,N_9431);
nand U13950 (N_13950,N_6650,N_11284);
xnor U13951 (N_13951,N_8320,N_8639);
xnor U13952 (N_13952,N_9393,N_7990);
or U13953 (N_13953,N_10285,N_9184);
or U13954 (N_13954,N_7116,N_7101);
nor U13955 (N_13955,N_8052,N_7731);
nand U13956 (N_13956,N_6099,N_8644);
or U13957 (N_13957,N_7241,N_7654);
nor U13958 (N_13958,N_10483,N_8449);
or U13959 (N_13959,N_10546,N_6510);
xor U13960 (N_13960,N_11228,N_8092);
nor U13961 (N_13961,N_8312,N_8271);
and U13962 (N_13962,N_11162,N_7423);
and U13963 (N_13963,N_9752,N_11968);
nand U13964 (N_13964,N_10320,N_9534);
and U13965 (N_13965,N_6648,N_9786);
and U13966 (N_13966,N_11760,N_8961);
nor U13967 (N_13967,N_7784,N_11451);
nor U13968 (N_13968,N_9824,N_6548);
and U13969 (N_13969,N_10590,N_6279);
nor U13970 (N_13970,N_11632,N_8683);
and U13971 (N_13971,N_11470,N_7303);
nand U13972 (N_13972,N_11328,N_11621);
nand U13973 (N_13973,N_8657,N_8739);
xnor U13974 (N_13974,N_8093,N_11917);
or U13975 (N_13975,N_10403,N_11810);
or U13976 (N_13976,N_7450,N_11855);
and U13977 (N_13977,N_8771,N_9978);
xnor U13978 (N_13978,N_9783,N_6373);
xnor U13979 (N_13979,N_11913,N_11705);
and U13980 (N_13980,N_6851,N_8730);
or U13981 (N_13981,N_6576,N_10733);
nor U13982 (N_13982,N_7651,N_9999);
nor U13983 (N_13983,N_6346,N_9227);
and U13984 (N_13984,N_8459,N_8915);
xor U13985 (N_13985,N_8787,N_9552);
or U13986 (N_13986,N_7467,N_10554);
xor U13987 (N_13987,N_9483,N_10810);
and U13988 (N_13988,N_8414,N_7323);
nor U13989 (N_13989,N_9979,N_11687);
nand U13990 (N_13990,N_6720,N_11369);
or U13991 (N_13991,N_7639,N_7078);
and U13992 (N_13992,N_8496,N_11418);
and U13993 (N_13993,N_8457,N_6868);
or U13994 (N_13994,N_10506,N_6569);
and U13995 (N_13995,N_6292,N_10749);
nor U13996 (N_13996,N_7573,N_6833);
or U13997 (N_13997,N_6542,N_6215);
nand U13998 (N_13998,N_9920,N_8351);
or U13999 (N_13999,N_10892,N_7104);
xor U14000 (N_14000,N_9564,N_11089);
nor U14001 (N_14001,N_8326,N_11116);
or U14002 (N_14002,N_11582,N_7727);
nand U14003 (N_14003,N_11672,N_6863);
nor U14004 (N_14004,N_6687,N_10276);
xor U14005 (N_14005,N_6624,N_10157);
and U14006 (N_14006,N_6282,N_11795);
or U14007 (N_14007,N_6572,N_9614);
and U14008 (N_14008,N_8037,N_10427);
or U14009 (N_14009,N_7605,N_8695);
nor U14010 (N_14010,N_9413,N_8580);
xor U14011 (N_14011,N_8566,N_6003);
and U14012 (N_14012,N_11292,N_11072);
xor U14013 (N_14013,N_11749,N_8813);
nor U14014 (N_14014,N_6229,N_7864);
xnor U14015 (N_14015,N_7023,N_7608);
nand U14016 (N_14016,N_10715,N_11351);
xnor U14017 (N_14017,N_9638,N_8301);
and U14018 (N_14018,N_7438,N_7349);
xnor U14019 (N_14019,N_6155,N_10149);
xnor U14020 (N_14020,N_8986,N_7279);
nand U14021 (N_14021,N_8332,N_10641);
or U14022 (N_14022,N_6280,N_6383);
or U14023 (N_14023,N_8317,N_7098);
and U14024 (N_14024,N_7761,N_9478);
xor U14025 (N_14025,N_6171,N_10461);
nand U14026 (N_14026,N_11486,N_11042);
xnor U14027 (N_14027,N_9121,N_6616);
and U14028 (N_14028,N_6584,N_6044);
and U14029 (N_14029,N_6757,N_9338);
or U14030 (N_14030,N_8409,N_11742);
xnor U14031 (N_14031,N_9963,N_10348);
nor U14032 (N_14032,N_8481,N_10572);
nor U14033 (N_14033,N_8661,N_10479);
nand U14034 (N_14034,N_11217,N_7717);
xor U14035 (N_14035,N_11368,N_6418);
nand U14036 (N_14036,N_7147,N_9128);
or U14037 (N_14037,N_11029,N_7196);
or U14038 (N_14038,N_11549,N_7338);
nor U14039 (N_14039,N_9109,N_10987);
nand U14040 (N_14040,N_10066,N_10902);
or U14041 (N_14041,N_6245,N_9238);
and U14042 (N_14042,N_10798,N_8361);
nor U14043 (N_14043,N_10236,N_11059);
nand U14044 (N_14044,N_11026,N_7706);
or U14045 (N_14045,N_10325,N_9605);
xor U14046 (N_14046,N_11908,N_7358);
or U14047 (N_14047,N_10939,N_6467);
and U14048 (N_14048,N_9612,N_7566);
and U14049 (N_14049,N_11095,N_8189);
nand U14050 (N_14050,N_9030,N_11758);
nor U14051 (N_14051,N_6228,N_8431);
nand U14052 (N_14052,N_7961,N_11691);
and U14053 (N_14053,N_6771,N_7690);
and U14054 (N_14054,N_6358,N_7728);
xor U14055 (N_14055,N_6439,N_6371);
and U14056 (N_14056,N_9942,N_8081);
xor U14057 (N_14057,N_6743,N_7546);
and U14058 (N_14058,N_10736,N_9417);
or U14059 (N_14059,N_11430,N_9686);
or U14060 (N_14060,N_10705,N_8561);
or U14061 (N_14061,N_11887,N_10956);
or U14062 (N_14062,N_11295,N_11318);
nand U14063 (N_14063,N_8477,N_7478);
nor U14064 (N_14064,N_11982,N_7666);
nor U14065 (N_14065,N_10224,N_11269);
and U14066 (N_14066,N_7018,N_10329);
nor U14067 (N_14067,N_6301,N_10891);
nor U14068 (N_14068,N_6302,N_9829);
xor U14069 (N_14069,N_9988,N_6887);
nand U14070 (N_14070,N_9893,N_8123);
nand U14071 (N_14071,N_6026,N_11056);
xnor U14072 (N_14072,N_6406,N_6745);
and U14073 (N_14073,N_7388,N_10967);
and U14074 (N_14074,N_8237,N_8698);
xnor U14075 (N_14075,N_10103,N_7721);
or U14076 (N_14076,N_7698,N_8498);
nand U14077 (N_14077,N_10102,N_8248);
xor U14078 (N_14078,N_11677,N_7926);
xor U14079 (N_14079,N_6643,N_8281);
nor U14080 (N_14080,N_7875,N_9482);
nor U14081 (N_14081,N_10303,N_10069);
xnor U14082 (N_14082,N_10244,N_10665);
or U14083 (N_14083,N_11725,N_8717);
or U14084 (N_14084,N_8655,N_6086);
nor U14085 (N_14085,N_6500,N_11250);
xor U14086 (N_14086,N_11354,N_10744);
nand U14087 (N_14087,N_11205,N_11519);
nand U14088 (N_14088,N_6046,N_9744);
nand U14089 (N_14089,N_10452,N_6839);
or U14090 (N_14090,N_7982,N_11604);
nand U14091 (N_14091,N_6331,N_11727);
nor U14092 (N_14092,N_8386,N_7941);
or U14093 (N_14093,N_8447,N_11063);
and U14094 (N_14094,N_10215,N_10947);
or U14095 (N_14095,N_7184,N_11575);
and U14096 (N_14096,N_11420,N_10369);
or U14097 (N_14097,N_11103,N_9369);
nor U14098 (N_14098,N_6252,N_9993);
nor U14099 (N_14099,N_11562,N_11213);
nor U14100 (N_14100,N_8845,N_10316);
and U14101 (N_14101,N_10364,N_9746);
or U14102 (N_14102,N_10928,N_7844);
nand U14103 (N_14103,N_9565,N_6917);
and U14104 (N_14104,N_8503,N_6188);
nand U14105 (N_14105,N_10214,N_11744);
nor U14106 (N_14106,N_6954,N_7642);
and U14107 (N_14107,N_11388,N_10814);
nor U14108 (N_14108,N_11937,N_7015);
nor U14109 (N_14109,N_11275,N_10228);
nand U14110 (N_14110,N_8494,N_7487);
or U14111 (N_14111,N_8919,N_8559);
and U14112 (N_14112,N_6391,N_7220);
and U14113 (N_14113,N_11053,N_10670);
or U14114 (N_14114,N_6987,N_9342);
or U14115 (N_14115,N_6506,N_11335);
nor U14116 (N_14116,N_8440,N_8273);
nand U14117 (N_14117,N_7455,N_6924);
and U14118 (N_14118,N_10173,N_10931);
or U14119 (N_14119,N_6958,N_6959);
nand U14120 (N_14120,N_7315,N_8512);
and U14121 (N_14121,N_7411,N_10376);
or U14122 (N_14122,N_9970,N_6444);
nor U14123 (N_14123,N_6615,N_7962);
nand U14124 (N_14124,N_7578,N_6897);
xor U14125 (N_14125,N_10984,N_8617);
or U14126 (N_14126,N_10708,N_9176);
and U14127 (N_14127,N_9743,N_6578);
and U14128 (N_14128,N_11449,N_8017);
nand U14129 (N_14129,N_6929,N_6840);
or U14130 (N_14130,N_7587,N_11428);
nand U14131 (N_14131,N_9203,N_11386);
or U14132 (N_14132,N_6619,N_9222);
nand U14133 (N_14133,N_6434,N_9318);
and U14134 (N_14134,N_9578,N_7069);
nor U14135 (N_14135,N_7402,N_10319);
or U14136 (N_14136,N_10062,N_9508);
or U14137 (N_14137,N_11494,N_8756);
xor U14138 (N_14138,N_10840,N_6635);
xor U14139 (N_14139,N_7635,N_7460);
nor U14140 (N_14140,N_6541,N_9033);
or U14141 (N_14141,N_6234,N_9822);
nand U14142 (N_14142,N_7379,N_11110);
nor U14143 (N_14143,N_9291,N_10660);
nand U14144 (N_14144,N_6646,N_6387);
nand U14145 (N_14145,N_7005,N_9077);
and U14146 (N_14146,N_11452,N_11154);
nand U14147 (N_14147,N_11457,N_9462);
or U14148 (N_14148,N_9704,N_6657);
nor U14149 (N_14149,N_6507,N_10716);
nor U14150 (N_14150,N_8984,N_6601);
or U14151 (N_14151,N_10941,N_11965);
and U14152 (N_14152,N_11401,N_6746);
and U14153 (N_14153,N_7765,N_8216);
xor U14154 (N_14154,N_7882,N_6214);
xor U14155 (N_14155,N_10150,N_7424);
nor U14156 (N_14156,N_9344,N_8523);
nand U14157 (N_14157,N_11998,N_11570);
or U14158 (N_14158,N_8142,N_10164);
and U14159 (N_14159,N_6815,N_6549);
or U14160 (N_14160,N_6272,N_10226);
nor U14161 (N_14161,N_7826,N_9293);
and U14162 (N_14162,N_8060,N_7140);
and U14163 (N_14163,N_7548,N_10123);
and U14164 (N_14164,N_8094,N_10411);
or U14165 (N_14165,N_6053,N_8029);
xnor U14166 (N_14166,N_10543,N_6162);
or U14167 (N_14167,N_9919,N_8712);
nor U14168 (N_14168,N_8363,N_11936);
and U14169 (N_14169,N_8372,N_8908);
nor U14170 (N_14170,N_8597,N_9698);
xor U14171 (N_14171,N_11972,N_9966);
or U14172 (N_14172,N_7874,N_9235);
and U14173 (N_14173,N_9558,N_8472);
and U14174 (N_14174,N_9453,N_9575);
and U14175 (N_14175,N_9760,N_6200);
or U14176 (N_14176,N_11573,N_7829);
nor U14177 (N_14177,N_10873,N_10239);
or U14178 (N_14178,N_9827,N_8535);
xnor U14179 (N_14179,N_6417,N_11066);
xor U14180 (N_14180,N_8733,N_8226);
or U14181 (N_14181,N_9986,N_8196);
xor U14182 (N_14182,N_8310,N_6195);
and U14183 (N_14183,N_11598,N_10667);
xnor U14184 (N_14184,N_7120,N_10490);
nand U14185 (N_14185,N_8562,N_9560);
nor U14186 (N_14186,N_8331,N_9027);
and U14187 (N_14187,N_8658,N_6117);
xnor U14188 (N_14188,N_11137,N_9629);
or U14189 (N_14189,N_9261,N_10557);
or U14190 (N_14190,N_7143,N_7521);
xnor U14191 (N_14191,N_7288,N_10740);
or U14192 (N_14192,N_10230,N_10124);
nand U14193 (N_14193,N_11265,N_8618);
nand U14194 (N_14194,N_8706,N_9655);
or U14195 (N_14195,N_7614,N_10922);
xor U14196 (N_14196,N_11427,N_7434);
and U14197 (N_14197,N_11692,N_7197);
xor U14198 (N_14198,N_6400,N_10449);
nor U14199 (N_14199,N_10818,N_11763);
and U14200 (N_14200,N_8156,N_11011);
nand U14201 (N_14201,N_8337,N_10776);
nor U14202 (N_14202,N_10537,N_7712);
nand U14203 (N_14203,N_10378,N_7929);
and U14204 (N_14204,N_8109,N_6932);
and U14205 (N_14205,N_10726,N_10535);
nand U14206 (N_14206,N_8070,N_11261);
xor U14207 (N_14207,N_8429,N_9939);
xnor U14208 (N_14208,N_11584,N_6613);
nor U14209 (N_14209,N_8667,N_8033);
nand U14210 (N_14210,N_10415,N_8400);
nor U14211 (N_14211,N_9135,N_6033);
and U14212 (N_14212,N_6864,N_10839);
nand U14213 (N_14213,N_6792,N_8395);
xnor U14214 (N_14214,N_7352,N_7281);
and U14215 (N_14215,N_11179,N_6435);
xnor U14216 (N_14216,N_7682,N_7815);
xnor U14217 (N_14217,N_7851,N_9509);
and U14218 (N_14218,N_11362,N_11237);
and U14219 (N_14219,N_10975,N_8890);
xor U14220 (N_14220,N_10769,N_6925);
xnor U14221 (N_14221,N_6964,N_8939);
xor U14222 (N_14222,N_11479,N_10570);
or U14223 (N_14223,N_11165,N_8034);
and U14224 (N_14224,N_11751,N_10550);
and U14225 (N_14225,N_8734,N_8246);
nor U14226 (N_14226,N_8240,N_9940);
xnor U14227 (N_14227,N_11524,N_6862);
xnor U14228 (N_14228,N_10903,N_8296);
and U14229 (N_14229,N_10888,N_9281);
nor U14230 (N_14230,N_9693,N_6194);
or U14231 (N_14231,N_10437,N_11317);
nand U14232 (N_14232,N_10948,N_9423);
xnor U14233 (N_14233,N_9971,N_6238);
xnor U14234 (N_14234,N_10837,N_9985);
nand U14235 (N_14235,N_8049,N_11170);
nor U14236 (N_14236,N_6175,N_6956);
and U14237 (N_14237,N_11301,N_10890);
nor U14238 (N_14238,N_11274,N_7774);
nand U14239 (N_14239,N_6306,N_9817);
or U14240 (N_14240,N_8153,N_7585);
xnor U14241 (N_14241,N_6531,N_6806);
or U14242 (N_14242,N_9328,N_10625);
or U14243 (N_14243,N_9732,N_9383);
and U14244 (N_14244,N_7282,N_7230);
nor U14245 (N_14245,N_9801,N_6730);
xor U14246 (N_14246,N_10053,N_7095);
and U14247 (N_14247,N_9000,N_6274);
nor U14248 (N_14248,N_7214,N_9914);
or U14249 (N_14249,N_7946,N_6706);
or U14250 (N_14250,N_10250,N_10751);
xor U14251 (N_14251,N_11338,N_10254);
xor U14252 (N_14252,N_8852,N_6641);
and U14253 (N_14253,N_6404,N_11268);
or U14254 (N_14254,N_11964,N_7617);
nand U14255 (N_14255,N_6212,N_11083);
and U14256 (N_14256,N_10357,N_10185);
nand U14257 (N_14257,N_10678,N_10821);
and U14258 (N_14258,N_11975,N_6653);
or U14259 (N_14259,N_10738,N_6555);
or U14260 (N_14260,N_6169,N_8601);
and U14261 (N_14261,N_10022,N_6836);
xnor U14262 (N_14262,N_10646,N_7165);
or U14263 (N_14263,N_11533,N_6208);
nor U14264 (N_14264,N_10233,N_9995);
or U14265 (N_14265,N_9507,N_10603);
and U14266 (N_14266,N_10876,N_10988);
nor U14267 (N_14267,N_7118,N_8591);
xnor U14268 (N_14268,N_7607,N_8328);
nand U14269 (N_14269,N_8428,N_10868);
nor U14270 (N_14270,N_8418,N_11051);
or U14271 (N_14271,N_6316,N_7276);
nand U14272 (N_14272,N_7342,N_11146);
or U14273 (N_14273,N_6106,N_9394);
xnor U14274 (N_14274,N_7973,N_7643);
nor U14275 (N_14275,N_9146,N_8171);
and U14276 (N_14276,N_6561,N_11733);
nor U14277 (N_14277,N_11915,N_9278);
nor U14278 (N_14278,N_9074,N_7624);
xor U14279 (N_14279,N_6797,N_6593);
or U14280 (N_14280,N_9609,N_7968);
nor U14281 (N_14281,N_10826,N_7674);
and U14282 (N_14282,N_10365,N_9265);
or U14283 (N_14283,N_7075,N_6986);
xnor U14284 (N_14284,N_10573,N_8013);
and U14285 (N_14285,N_8393,N_8564);
and U14286 (N_14286,N_9696,N_11889);
or U14287 (N_14287,N_9749,N_6243);
xor U14288 (N_14288,N_7090,N_6776);
xor U14289 (N_14289,N_11828,N_10954);
and U14290 (N_14290,N_6382,N_6498);
nand U14291 (N_14291,N_10405,N_9233);
and U14292 (N_14292,N_7785,N_11435);
or U14293 (N_14293,N_7699,N_10431);
nand U14294 (N_14294,N_8820,N_7153);
or U14295 (N_14295,N_6104,N_11927);
nor U14296 (N_14296,N_7853,N_8910);
or U14297 (N_14297,N_10632,N_10134);
or U14298 (N_14298,N_6988,N_9312);
xor U14299 (N_14299,N_7051,N_11077);
nand U14300 (N_14300,N_11762,N_11081);
nor U14301 (N_14301,N_11682,N_6799);
xnor U14302 (N_14302,N_9487,N_8422);
and U14303 (N_14303,N_10441,N_10478);
or U14304 (N_14304,N_11920,N_11660);
and U14305 (N_14305,N_9588,N_10249);
nand U14306 (N_14306,N_6733,N_11544);
or U14307 (N_14307,N_9492,N_8230);
nand U14308 (N_14308,N_8068,N_8558);
xnor U14309 (N_14309,N_11818,N_7444);
nand U14310 (N_14310,N_11222,N_6001);
nor U14311 (N_14311,N_9516,N_7847);
or U14312 (N_14312,N_8871,N_7870);
and U14313 (N_14313,N_10090,N_8161);
or U14314 (N_14314,N_6620,N_10004);
xnor U14315 (N_14315,N_8444,N_10611);
or U14316 (N_14316,N_10836,N_11792);
or U14317 (N_14317,N_6942,N_6716);
or U14318 (N_14318,N_10163,N_6307);
and U14319 (N_14319,N_7515,N_7210);
nand U14320 (N_14320,N_9582,N_11521);
and U14321 (N_14321,N_11234,N_8716);
xnor U14322 (N_14322,N_7987,N_7730);
nor U14323 (N_14323,N_9785,N_7162);
and U14324 (N_14324,N_6211,N_7633);
and U14325 (N_14325,N_8389,N_7800);
or U14326 (N_14326,N_6262,N_10473);
nor U14327 (N_14327,N_11590,N_11247);
nor U14328 (N_14328,N_6902,N_6124);
nand U14329 (N_14329,N_9681,N_7913);
and U14330 (N_14330,N_8495,N_11400);
xnor U14331 (N_14331,N_10268,N_11015);
nor U14332 (N_14332,N_6111,N_7310);
xor U14333 (N_14333,N_8958,N_8187);
xnor U14334 (N_14334,N_8176,N_7429);
nor U14335 (N_14335,N_8197,N_8124);
xor U14336 (N_14336,N_8544,N_9990);
and U14337 (N_14337,N_6893,N_8729);
and U14338 (N_14338,N_7369,N_10240);
xor U14339 (N_14339,N_6134,N_9631);
xor U14340 (N_14340,N_10683,N_7283);
nand U14341 (N_14341,N_11468,N_10400);
and U14342 (N_14342,N_6763,N_9718);
or U14343 (N_14343,N_7195,N_6927);
nand U14344 (N_14344,N_6395,N_8680);
and U14345 (N_14345,N_10159,N_6029);
xor U14346 (N_14346,N_8883,N_10808);
or U14347 (N_14347,N_8074,N_10841);
and U14348 (N_14348,N_8560,N_10643);
nor U14349 (N_14349,N_10675,N_7290);
nand U14350 (N_14350,N_10308,N_7541);
or U14351 (N_14351,N_11176,N_8242);
xnor U14352 (N_14352,N_6659,N_8988);
xor U14353 (N_14353,N_11643,N_10140);
nand U14354 (N_14354,N_11023,N_8711);
xor U14355 (N_14355,N_6894,N_9424);
and U14356 (N_14356,N_7249,N_11668);
nor U14357 (N_14357,N_11989,N_10217);
nor U14358 (N_14358,N_6210,N_11626);
xor U14359 (N_14359,N_7862,N_9811);
nand U14360 (N_14360,N_10674,N_9145);
or U14361 (N_14361,N_9804,N_6906);
and U14362 (N_14362,N_7160,N_6854);
xnor U14363 (N_14363,N_10819,N_8710);
and U14364 (N_14364,N_9165,N_6120);
and U14365 (N_14365,N_7933,N_11773);
or U14366 (N_14366,N_6180,N_10549);
and U14367 (N_14367,N_10139,N_8018);
and U14368 (N_14368,N_11280,N_9243);
nor U14369 (N_14369,N_9808,N_8203);
nor U14370 (N_14370,N_11107,N_10016);
nand U14371 (N_14371,N_8287,N_7383);
nand U14372 (N_14372,N_9803,N_11719);
or U14373 (N_14373,N_8675,N_9093);
or U14374 (N_14374,N_8260,N_7072);
or U14375 (N_14375,N_9866,N_10882);
nor U14376 (N_14376,N_11365,N_6242);
xnor U14377 (N_14377,N_8390,N_11735);
xor U14378 (N_14378,N_10629,N_11656);
or U14379 (N_14379,N_7627,N_11859);
nor U14380 (N_14380,N_8830,N_11441);
or U14381 (N_14381,N_6216,N_7538);
and U14382 (N_14382,N_9032,N_10696);
or U14383 (N_14383,N_8218,N_8807);
nand U14384 (N_14384,N_10097,N_11407);
nand U14385 (N_14385,N_11346,N_11567);
and U14386 (N_14386,N_11130,N_10237);
xnor U14387 (N_14387,N_7942,N_8322);
nand U14388 (N_14388,N_8862,N_11343);
or U14389 (N_14389,N_10654,N_6534);
xnor U14390 (N_14390,N_11756,N_10957);
xnor U14391 (N_14391,N_10132,N_6923);
nor U14392 (N_14392,N_11139,N_9210);
nor U14393 (N_14393,N_10033,N_9108);
and U14394 (N_14394,N_9308,N_10779);
or U14395 (N_14395,N_8469,N_10326);
and U14396 (N_14396,N_7512,N_8433);
and U14397 (N_14397,N_9015,N_9177);
nand U14398 (N_14398,N_9778,N_8602);
nand U14399 (N_14399,N_10904,N_9268);
nor U14400 (N_14400,N_6568,N_11151);
xnor U14401 (N_14401,N_7332,N_8175);
nand U14402 (N_14402,N_7387,N_8546);
nand U14403 (N_14403,N_10657,N_8780);
nor U14404 (N_14404,N_9144,N_10886);
nor U14405 (N_14405,N_7876,N_10335);
or U14406 (N_14406,N_8204,N_9498);
nand U14407 (N_14407,N_6744,N_6547);
and U14408 (N_14408,N_6058,N_6483);
nor U14409 (N_14409,N_10681,N_6119);
nor U14410 (N_14410,N_8974,N_7530);
nor U14411 (N_14411,N_11105,N_9860);
xor U14412 (N_14412,N_8000,N_9181);
xor U14413 (N_14413,N_11830,N_8689);
or U14414 (N_14414,N_10728,N_7497);
xnor U14415 (N_14415,N_8972,N_7644);
and U14416 (N_14416,N_11192,N_8452);
and U14417 (N_14417,N_9223,N_6057);
xor U14418 (N_14418,N_9191,N_7854);
xnor U14419 (N_14419,N_9593,N_11434);
nor U14420 (N_14420,N_7294,N_6204);
nor U14421 (N_14421,N_8549,N_10128);
xnor U14422 (N_14422,N_11648,N_11609);
nand U14423 (N_14423,N_11119,N_8004);
nand U14424 (N_14424,N_6311,N_10169);
xor U14425 (N_14425,N_10484,N_10290);
or U14426 (N_14426,N_11253,N_11574);
nor U14427 (N_14427,N_11489,N_6038);
or U14428 (N_14428,N_7219,N_9982);
or U14429 (N_14429,N_6802,N_8861);
or U14430 (N_14430,N_8061,N_11939);
nand U14431 (N_14431,N_9329,N_9494);
nor U14432 (N_14432,N_7408,N_7533);
and U14433 (N_14433,N_7991,N_11620);
and U14434 (N_14434,N_9111,N_9147);
or U14435 (N_14435,N_9603,N_8304);
xor U14436 (N_14436,N_6629,N_9239);
and U14437 (N_14437,N_7885,N_7684);
nor U14438 (N_14438,N_8949,N_9574);
and U14439 (N_14439,N_9948,N_7106);
or U14440 (N_14440,N_11446,N_9347);
nor U14441 (N_14441,N_11223,N_6016);
nor U14442 (N_14442,N_6524,N_6079);
nand U14443 (N_14443,N_10824,N_6052);
nor U14444 (N_14444,N_7105,N_7623);
or U14445 (N_14445,N_9187,N_10936);
xor U14446 (N_14446,N_7179,N_7886);
xnor U14447 (N_14447,N_6794,N_6980);
and U14448 (N_14448,N_9840,N_6679);
xnor U14449 (N_14449,N_7341,N_6020);
and U14450 (N_14450,N_11698,N_7420);
or U14451 (N_14451,N_8839,N_8850);
and U14452 (N_14452,N_10084,N_6494);
xor U14453 (N_14453,N_8809,N_7034);
and U14454 (N_14454,N_7906,N_8399);
xnor U14455 (N_14455,N_6562,N_10471);
nor U14456 (N_14456,N_6838,N_9625);
xnor U14457 (N_14457,N_10086,N_9674);
xor U14458 (N_14458,N_9882,N_8914);
xor U14459 (N_14459,N_10930,N_11639);
or U14460 (N_14460,N_10451,N_7414);
nand U14461 (N_14461,N_7469,N_10848);
or U14462 (N_14462,N_11319,N_9399);
xnor U14463 (N_14463,N_9374,N_7795);
or U14464 (N_14464,N_10104,N_9515);
and U14465 (N_14465,N_11440,N_10536);
or U14466 (N_14466,N_9800,N_8329);
nor U14467 (N_14467,N_10077,N_10946);
xnor U14468 (N_14468,N_7799,N_11031);
or U14469 (N_14469,N_7509,N_8704);
xnor U14470 (N_14470,N_7243,N_6828);
nand U14471 (N_14471,N_11392,N_10346);
and U14472 (N_14472,N_11708,N_10023);
and U14473 (N_14473,N_9831,N_6822);
nand U14474 (N_14474,N_6871,N_7451);
xor U14475 (N_14475,N_8294,N_6367);
and U14476 (N_14476,N_9865,N_7109);
or U14477 (N_14477,N_10009,N_11178);
nand U14478 (N_14478,N_6133,N_11509);
xnor U14479 (N_14479,N_8696,N_7561);
and U14480 (N_14480,N_6313,N_10418);
and U14481 (N_14481,N_11898,N_11197);
nand U14482 (N_14482,N_8599,N_11474);
xor U14483 (N_14483,N_6172,N_8775);
or U14484 (N_14484,N_8866,N_10296);
and U14485 (N_14485,N_10409,N_11872);
nor U14486 (N_14486,N_7113,N_10213);
or U14487 (N_14487,N_8750,N_11793);
or U14488 (N_14488,N_7430,N_11731);
or U14489 (N_14489,N_11844,N_9251);
xor U14490 (N_14490,N_11612,N_6032);
xnor U14491 (N_14491,N_7969,N_8213);
nor U14492 (N_14492,N_8374,N_8678);
nand U14493 (N_14493,N_11637,N_11761);
or U14494 (N_14494,N_7137,N_11262);
nand U14495 (N_14495,N_11414,N_9845);
xnor U14496 (N_14496,N_10602,N_10748);
xor U14497 (N_14497,N_6157,N_10168);
or U14498 (N_14498,N_11693,N_8697);
nand U14499 (N_14499,N_8859,N_11912);
nand U14500 (N_14500,N_10833,N_7518);
and U14501 (N_14501,N_10001,N_9113);
or U14502 (N_14502,N_8155,N_10766);
and U14503 (N_14503,N_9660,N_10970);
xor U14504 (N_14504,N_9241,N_6546);
or U14505 (N_14505,N_9258,N_10752);
and U14506 (N_14506,N_9748,N_9863);
nor U14507 (N_14507,N_11807,N_7975);
nor U14508 (N_14508,N_7495,N_7057);
nor U14509 (N_14509,N_11720,N_7302);
nor U14510 (N_14510,N_10830,N_6035);
nor U14511 (N_14511,N_7796,N_6823);
nor U14512 (N_14512,N_9208,N_11589);
or U14513 (N_14513,N_7100,N_11445);
nor U14514 (N_14514,N_9377,N_9735);
nand U14515 (N_14515,N_8256,N_6139);
nor U14516 (N_14516,N_11186,N_11808);
nor U14517 (N_14517,N_6591,N_11499);
nand U14518 (N_14518,N_6263,N_10908);
xnor U14519 (N_14519,N_11606,N_6729);
nor U14520 (N_14520,N_6277,N_11329);
xor U14521 (N_14521,N_10087,N_7865);
xor U14522 (N_14522,N_6059,N_9123);
or U14523 (N_14523,N_9449,N_6951);
nand U14524 (N_14524,N_8179,N_6829);
and U14525 (N_14525,N_8966,N_8848);
nand U14526 (N_14526,N_7896,N_11248);
xor U14527 (N_14527,N_8989,N_8214);
nor U14528 (N_14528,N_10923,N_8703);
and U14529 (N_14529,N_6567,N_6585);
xnor U14530 (N_14530,N_11334,N_6544);
nand U14531 (N_14531,N_8540,N_7850);
xnor U14532 (N_14532,N_10601,N_7073);
and U14533 (N_14533,N_10619,N_9043);
or U14534 (N_14534,N_11506,N_9447);
nand U14535 (N_14535,N_7193,N_10909);
or U14536 (N_14536,N_8040,N_7752);
nand U14537 (N_14537,N_7663,N_10207);
and U14538 (N_14538,N_11444,N_7845);
nand U14539 (N_14539,N_9526,N_8772);
or U14540 (N_14540,N_7877,N_9339);
nand U14541 (N_14541,N_9021,N_6266);
xnor U14542 (N_14542,N_9476,N_7308);
nor U14543 (N_14543,N_7925,N_6132);
and U14544 (N_14544,N_7772,N_8688);
or U14545 (N_14545,N_6197,N_11135);
nor U14546 (N_14546,N_9835,N_7919);
and U14547 (N_14547,N_8076,N_6091);
nand U14548 (N_14548,N_7406,N_11160);
xor U14549 (N_14549,N_9881,N_7360);
or U14550 (N_14550,N_6310,N_11364);
nand U14551 (N_14551,N_10042,N_8292);
or U14552 (N_14552,N_10492,N_9792);
xnor U14553 (N_14553,N_7204,N_9750);
or U14554 (N_14554,N_8791,N_8019);
nor U14555 (N_14555,N_10367,N_11353);
or U14556 (N_14556,N_9196,N_7988);
or U14557 (N_14557,N_10154,N_7347);
xnor U14558 (N_14558,N_6752,N_11093);
or U14559 (N_14559,N_11502,N_9601);
nor U14560 (N_14560,N_6652,N_10907);
and U14561 (N_14561,N_6386,N_7086);
and U14562 (N_14562,N_9270,N_8150);
nor U14563 (N_14563,N_7084,N_6631);
or U14564 (N_14564,N_7836,N_9781);
and U14565 (N_14565,N_8302,N_6077);
xor U14566 (N_14566,N_8529,N_10844);
xnor U14567 (N_14567,N_8108,N_8466);
xor U14568 (N_14568,N_6261,N_10631);
xor U14569 (N_14569,N_6334,N_11557);
nor U14570 (N_14570,N_8649,N_6186);
nand U14571 (N_14571,N_6946,N_9441);
and U14572 (N_14572,N_6191,N_8252);
and U14573 (N_14573,N_7953,N_6997);
nand U14574 (N_14574,N_10605,N_11597);
or U14575 (N_14575,N_10624,N_7161);
nor U14576 (N_14576,N_10067,N_8833);
nand U14577 (N_14577,N_9889,N_9844);
nor U14578 (N_14578,N_10689,N_8072);
or U14579 (N_14579,N_9391,N_10514);
and U14580 (N_14580,N_11024,N_11999);
nand U14581 (N_14581,N_8825,N_7917);
nand U14582 (N_14582,N_11836,N_10391);
and U14583 (N_14583,N_8579,N_10780);
nand U14584 (N_14584,N_10256,N_9193);
nor U14585 (N_14585,N_7525,N_9941);
xnor U14586 (N_14586,N_6784,N_6707);
nand U14587 (N_14587,N_8719,N_6719);
xor U14588 (N_14588,N_7437,N_8358);
or U14589 (N_14589,N_11934,N_7304);
or U14590 (N_14590,N_10313,N_10638);
and U14591 (N_14591,N_7112,N_9615);
xor U14592 (N_14592,N_11766,N_11522);
and U14593 (N_14593,N_9257,N_6760);
and U14594 (N_14594,N_10920,N_8911);
xor U14595 (N_14595,N_10977,N_7237);
nor U14596 (N_14596,N_9136,N_10576);
or U14597 (N_14597,N_7400,N_6037);
or U14598 (N_14598,N_9133,N_11608);
nand U14599 (N_14599,N_7470,N_7003);
and U14600 (N_14600,N_11946,N_8937);
nand U14601 (N_14601,N_9341,N_11529);
xnor U14602 (N_14602,N_8742,N_9282);
and U14603 (N_14603,N_9142,N_8388);
and U14604 (N_14604,N_6831,N_10897);
xor U14605 (N_14605,N_6340,N_10571);
nand U14606 (N_14606,N_8844,N_7235);
and U14607 (N_14607,N_6366,N_6276);
and U14608 (N_14608,N_6022,N_7529);
xnor U14609 (N_14609,N_11706,N_7557);
nor U14610 (N_14610,N_10058,N_9839);
or U14611 (N_14611,N_10196,N_7336);
nor U14612 (N_14612,N_7726,N_6793);
and U14613 (N_14613,N_9370,N_9298);
xor U14614 (N_14614,N_11313,N_10440);
and U14615 (N_14615,N_11921,N_7510);
xnor U14616 (N_14616,N_9510,N_11320);
or U14617 (N_14617,N_8543,N_9580);
nor U14618 (N_14618,N_8229,N_11558);
and U14619 (N_14619,N_11350,N_7207);
and U14620 (N_14620,N_9769,N_9168);
nand U14621 (N_14621,N_7734,N_6879);
nand U14622 (N_14622,N_6318,N_10195);
and U14623 (N_14623,N_10528,N_9094);
xnor U14624 (N_14624,N_6528,N_10193);
nand U14625 (N_14625,N_11355,N_9964);
nand U14626 (N_14626,N_9955,N_8896);
xor U14627 (N_14627,N_10498,N_8684);
and U14628 (N_14628,N_8603,N_8721);
or U14629 (N_14629,N_6698,N_9891);
nor U14630 (N_14630,N_7028,N_7883);
xor U14631 (N_14631,N_9646,N_8250);
or U14632 (N_14632,N_8933,N_9173);
nand U14633 (N_14633,N_6963,N_9883);
nand U14634 (N_14634,N_11569,N_10426);
or U14635 (N_14635,N_10874,N_6362);
or U14636 (N_14636,N_9230,N_8731);
xor U14637 (N_14637,N_10815,N_10280);
nor U14638 (N_14638,N_7776,N_11554);
or U14639 (N_14639,N_9016,N_10374);
nand U14640 (N_14640,N_7327,N_11058);
nor U14641 (N_14641,N_6429,N_10302);
nor U14642 (N_14642,N_7435,N_8423);
or U14643 (N_14643,N_8453,N_11520);
and U14644 (N_14644,N_11503,N_9175);
nor U14645 (N_14645,N_7466,N_7808);
and U14646 (N_14646,N_8590,N_9962);
xnor U14647 (N_14647,N_8270,N_6397);
or U14648 (N_14648,N_11715,N_7951);
nor U14649 (N_14649,N_10916,N_11033);
or U14650 (N_14650,N_9010,N_7516);
nand U14651 (N_14651,N_7493,N_10729);
or U14652 (N_14652,N_11299,N_8215);
nand U14653 (N_14653,N_10487,N_11747);
xor U14654 (N_14654,N_10184,N_11552);
xor U14655 (N_14655,N_9070,N_11940);
nor U14656 (N_14656,N_8930,N_6783);
nand U14657 (N_14657,N_9950,N_8927);
xor U14658 (N_14658,N_6685,N_6703);
nand U14659 (N_14659,N_9586,N_9570);
and U14660 (N_14660,N_9722,N_11885);
nand U14661 (N_14661,N_7839,N_6993);
nor U14662 (N_14662,N_6341,N_7954);
nand U14663 (N_14663,N_8997,N_11929);
xor U14664 (N_14664,N_11084,N_6581);
or U14665 (N_14665,N_6995,N_9771);
xor U14666 (N_14666,N_6105,N_10613);
or U14667 (N_14667,N_9028,N_6898);
nor U14668 (N_14668,N_7040,N_11862);
nor U14669 (N_14669,N_10413,N_8737);
nand U14670 (N_14670,N_9853,N_6152);
nand U14671 (N_14671,N_6884,N_7229);
xor U14672 (N_14672,N_7750,N_6713);
and U14673 (N_14673,N_7415,N_9323);
nor U14674 (N_14674,N_7958,N_9520);
or U14675 (N_14675,N_8528,N_8115);
or U14676 (N_14676,N_8297,N_6515);
nand U14677 (N_14677,N_11635,N_8724);
xor U14678 (N_14678,N_10412,N_6288);
xnor U14679 (N_14679,N_8476,N_9200);
nand U14680 (N_14680,N_8816,N_9365);
or U14681 (N_14681,N_10071,N_7188);
and U14682 (N_14682,N_10753,N_7927);
nand U14683 (N_14683,N_8944,N_6236);
nand U14684 (N_14684,N_11443,N_7321);
nand U14685 (N_14685,N_9499,N_6381);
and U14686 (N_14686,N_8369,N_10216);
or U14687 (N_14687,N_6425,N_9287);
and U14688 (N_14688,N_9946,N_8835);
xnor U14689 (N_14689,N_11189,N_9058);
and U14690 (N_14690,N_9009,N_7646);
nand U14691 (N_14691,N_11045,N_10763);
nor U14692 (N_14692,N_10456,N_6759);
or U14693 (N_14693,N_8645,N_8723);
and U14694 (N_14694,N_10747,N_9864);
or U14695 (N_14695,N_8880,N_10386);
nor U14696 (N_14696,N_6151,N_11485);
and U14697 (N_14697,N_6941,N_6377);
or U14698 (N_14698,N_8922,N_9613);
and U14699 (N_14699,N_10089,N_10120);
and U14700 (N_14700,N_6256,N_9324);
and U14701 (N_14701,N_9496,N_6516);
or U14702 (N_14702,N_8112,N_9325);
nand U14703 (N_14703,N_7221,N_6804);
nand U14704 (N_14704,N_7806,N_11856);
or U14705 (N_14705,N_7502,N_7312);
or U14706 (N_14706,N_6856,N_6493);
nor U14707 (N_14707,N_8851,N_9075);
nand U14708 (N_14708,N_7665,N_6110);
xnor U14709 (N_14709,N_6379,N_6462);
nor U14710 (N_14710,N_11556,N_7879);
nand U14711 (N_14711,N_6095,N_9426);
nand U14712 (N_14712,N_8620,N_9412);
and U14713 (N_14713,N_7074,N_7397);
and U14714 (N_14714,N_8720,N_7767);
or U14715 (N_14715,N_9138,N_10796);
nand U14716 (N_14716,N_7884,N_10344);
nand U14717 (N_14717,N_9002,N_7231);
nand U14718 (N_14718,N_11772,N_10896);
or U14719 (N_14719,N_10429,N_7920);
xor U14720 (N_14720,N_10384,N_10561);
nor U14721 (N_14721,N_8624,N_10578);
and U14722 (N_14722,N_11252,N_6051);
nor U14723 (N_14723,N_6983,N_11067);
nand U14724 (N_14724,N_8254,N_6705);
and U14725 (N_14725,N_6915,N_8970);
nor U14726 (N_14726,N_10152,N_7482);
xor U14727 (N_14727,N_6088,N_7636);
nor U14728 (N_14728,N_11171,N_11592);
xnor U14729 (N_14729,N_6350,N_10289);
xnor U14730 (N_14730,N_10699,N_8300);
or U14731 (N_14731,N_7810,N_10388);
and U14732 (N_14732,N_10110,N_11330);
and U14733 (N_14733,N_9240,N_7719);
nand U14734 (N_14734,N_8836,N_9153);
xnor U14735 (N_14735,N_9055,N_10912);
or U14736 (N_14736,N_8951,N_7355);
xor U14737 (N_14737,N_9954,N_11674);
and U14738 (N_14738,N_7560,N_8516);
or U14739 (N_14739,N_9467,N_8080);
and U14740 (N_14740,N_6012,N_10917);
xnor U14741 (N_14741,N_6773,N_7671);
nor U14742 (N_14742,N_6207,N_9180);
and U14743 (N_14743,N_7822,N_8555);
nor U14744 (N_14744,N_7087,N_11790);
nand U14745 (N_14745,N_6791,N_8298);
nor U14746 (N_14746,N_10297,N_9171);
nor U14747 (N_14747,N_10949,N_7142);
and U14748 (N_14748,N_9868,N_6101);
or U14749 (N_14749,N_6464,N_8032);
xnor U14750 (N_14750,N_7458,N_7816);
nand U14751 (N_14751,N_6558,N_11281);
nand U14752 (N_14752,N_7092,N_7218);
or U14753 (N_14753,N_9379,N_8759);
nor U14754 (N_14754,N_10999,N_8794);
xor U14755 (N_14755,N_9212,N_6140);
xor U14756 (N_14756,N_11206,N_8763);
nor U14757 (N_14757,N_9826,N_10399);
and U14758 (N_14758,N_6108,N_7311);
or U14759 (N_14759,N_8141,N_9967);
nand U14760 (N_14760,N_8318,N_9167);
nor U14761 (N_14761,N_6910,N_8383);
nand U14762 (N_14762,N_8378,N_9634);
nor U14763 (N_14763,N_11688,N_6349);
xor U14764 (N_14764,N_6835,N_9620);
nand U14765 (N_14765,N_9876,N_8314);
xnor U14766 (N_14766,N_11892,N_9279);
or U14767 (N_14767,N_11287,N_8613);
xor U14768 (N_14768,N_11864,N_7194);
nand U14769 (N_14769,N_11161,N_11853);
xor U14770 (N_14770,N_11022,N_7299);
or U14771 (N_14771,N_10707,N_10305);
xnor U14772 (N_14772,N_10112,N_7517);
nor U14773 (N_14773,N_7910,N_10306);
nand U14774 (N_14774,N_6085,N_10704);
xnor U14775 (N_14775,N_10875,N_9414);
and U14776 (N_14776,N_8050,N_10389);
and U14777 (N_14777,N_9317,N_8046);
nor U14778 (N_14778,N_7445,N_11838);
or U14779 (N_14779,N_11185,N_10614);
nor U14780 (N_14780,N_7038,N_7575);
or U14781 (N_14781,N_10420,N_6790);
and U14782 (N_14782,N_6076,N_10739);
and U14783 (N_14783,N_7339,N_6190);
nand U14784 (N_14784,N_9156,N_6490);
or U14785 (N_14785,N_8979,N_9401);
xnor U14786 (N_14786,N_7182,N_11109);
nor U14787 (N_14787,N_7088,N_9694);
or U14788 (N_14788,N_11114,N_8065);
or U14789 (N_14789,N_6329,N_10508);
and U14790 (N_14790,N_7980,N_7056);
xnor U14791 (N_14791,N_6304,N_8872);
and U14792 (N_14792,N_9987,N_11694);
or U14793 (N_14793,N_8714,N_8368);
xor U14794 (N_14794,N_9931,N_8488);
nand U14795 (N_14795,N_9788,N_10177);
nor U14796 (N_14796,N_11291,N_10963);
xor U14797 (N_14797,N_7820,N_7136);
or U14798 (N_14798,N_9585,N_11421);
or U14799 (N_14799,N_8738,N_8786);
nand U14800 (N_14800,N_6158,N_6315);
and U14801 (N_14801,N_11508,N_9435);
or U14802 (N_14802,N_11820,N_10926);
nand U14803 (N_14803,N_9343,N_7462);
or U14804 (N_14804,N_9104,N_6289);
nor U14805 (N_14805,N_7351,N_7248);
or U14806 (N_14806,N_10801,N_9828);
xor U14807 (N_14807,N_10061,N_11325);
and U14808 (N_14808,N_11933,N_8114);
xnor U14809 (N_14809,N_6731,N_8245);
nor U14810 (N_14810,N_11038,N_10721);
and U14811 (N_14811,N_6669,N_6437);
nor U14812 (N_14812,N_10068,N_7461);
and U14813 (N_14813,N_10854,N_6536);
nor U14814 (N_14814,N_9061,N_7280);
nand U14815 (N_14815,N_7769,N_10232);
and U14816 (N_14816,N_9217,N_7658);
nor U14817 (N_14817,N_8159,N_7505);
or U14818 (N_14818,N_10379,N_7322);
and U14819 (N_14819,N_7180,N_9455);
xor U14820 (N_14820,N_10513,N_9003);
nor U14821 (N_14821,N_8847,N_6818);
nor U14822 (N_14822,N_7940,N_10951);
and U14823 (N_14823,N_11091,N_10913);
or U14824 (N_14824,N_8921,N_8269);
nand U14825 (N_14825,N_8647,N_7277);
and U14826 (N_14826,N_10234,N_9428);
xor U14827 (N_14827,N_6800,N_7309);
nor U14828 (N_14828,N_9255,N_9359);
and U14829 (N_14829,N_7700,N_7258);
xnor U14830 (N_14830,N_11724,N_7416);
and U14831 (N_14831,N_8768,N_7163);
xnor U14832 (N_14832,N_7394,N_9506);
nand U14833 (N_14833,N_10094,N_8811);
or U14834 (N_14834,N_11078,N_6592);
xor U14835 (N_14835,N_8293,N_7963);
or U14836 (N_14836,N_6451,N_6974);
nor U14837 (N_14837,N_9806,N_9849);
nand U14838 (N_14838,N_10385,N_9457);
or U14839 (N_14839,N_10200,N_9225);
and U14840 (N_14840,N_11538,N_11149);
or U14841 (N_14841,N_6121,N_9633);
nand U14842 (N_14842,N_8405,N_6686);
nor U14843 (N_14843,N_11378,N_8677);
or U14844 (N_14844,N_9707,N_8199);
or U14845 (N_14845,N_10853,N_9672);
nand U14846 (N_14846,N_9782,N_9927);
nor U14847 (N_14847,N_9283,N_8586);
or U14848 (N_14848,N_9532,N_9220);
nor U14849 (N_14849,N_9277,N_6424);
or U14850 (N_14850,N_7574,N_9994);
or U14851 (N_14851,N_8434,N_7501);
nand U14852 (N_14852,N_9481,N_7704);
nor U14853 (N_14853,N_10760,N_6203);
or U14854 (N_14854,N_7166,N_11931);
or U14855 (N_14855,N_6491,N_7934);
nand U14856 (N_14856,N_11510,N_9794);
nor U14857 (N_14857,N_7030,N_8936);
or U14858 (N_14858,N_10045,N_6144);
and U14859 (N_14859,N_7211,N_8526);
xnor U14860 (N_14860,N_6627,N_10222);
or U14861 (N_14861,N_7604,N_11008);
nand U14862 (N_14862,N_9937,N_11086);
and U14863 (N_14863,N_9666,N_10156);
xnor U14864 (N_14864,N_10730,N_11096);
xnor U14865 (N_14865,N_6676,N_8120);
or U14866 (N_14866,N_9007,N_11202);
or U14867 (N_14867,N_7893,N_6479);
or U14868 (N_14868,N_10869,N_8551);
nand U14869 (N_14869,N_7522,N_8584);
xnor U14870 (N_14870,N_6135,N_9821);
and U14871 (N_14871,N_8751,N_7722);
xnor U14872 (N_14872,N_9041,N_8778);
nor U14873 (N_14873,N_9463,N_10556);
nor U14874 (N_14874,N_9122,N_7945);
and U14875 (N_14875,N_10857,N_9728);
nand U14876 (N_14876,N_8313,N_10644);
nor U14877 (N_14877,N_6660,N_6626);
nor U14878 (N_14878,N_9805,N_11195);
nand U14879 (N_14879,N_9924,N_10835);
xnor U14880 (N_14880,N_8480,N_9627);
nor U14881 (N_14881,N_6445,N_10552);
or U14882 (N_14882,N_7173,N_7830);
and U14883 (N_14883,N_11881,N_9272);
or U14884 (N_14884,N_9802,N_8277);
xor U14885 (N_14885,N_11594,N_6617);
nor U14886 (N_14886,N_9047,N_7743);
nand U14887 (N_14887,N_10649,N_9411);
nor U14888 (N_14888,N_11342,N_9095);
xor U14889 (N_14889,N_11492,N_6754);
and U14890 (N_14890,N_6965,N_8585);
nor U14891 (N_14891,N_6343,N_6727);
or U14892 (N_14892,N_10432,N_9368);
xnor U14893 (N_14893,N_8869,N_10231);
nor U14894 (N_14894,N_10013,N_9798);
nor U14895 (N_14895,N_10208,N_9624);
nor U14896 (N_14896,N_10628,N_11459);
and U14897 (N_14897,N_6118,N_10706);
nor U14898 (N_14898,N_8470,N_9364);
xnor U14899 (N_14899,N_6156,N_8898);
xor U14900 (N_14900,N_10130,N_9183);
and U14901 (N_14901,N_9114,N_10617);
nand U14902 (N_14902,N_10465,N_11678);
or U14903 (N_14903,N_8411,N_11980);
nor U14904 (N_14904,N_10943,N_10974);
nand U14905 (N_14905,N_9367,N_6294);
or U14906 (N_14906,N_8600,N_10515);
nand U14907 (N_14907,N_10148,N_11811);
xor U14908 (N_14908,N_11505,N_7457);
or U14909 (N_14909,N_10352,N_11054);
and U14910 (N_14910,N_6926,N_6931);
or U14911 (N_14911,N_11970,N_7135);
and U14912 (N_14912,N_10812,N_11987);
or U14913 (N_14913,N_7760,N_7887);
nand U14914 (N_14914,N_6073,N_10687);
xnor U14915 (N_14915,N_11755,N_10698);
nor U14916 (N_14916,N_8064,N_8891);
nand U14917 (N_14917,N_10623,N_9838);
or U14918 (N_14918,N_11120,N_7010);
nor U14919 (N_14919,N_10181,N_8163);
nand U14920 (N_14920,N_8777,N_7037);
nor U14921 (N_14921,N_10481,N_11270);
nor U14922 (N_14922,N_9500,N_6937);
nand U14923 (N_14923,N_6841,N_11944);
xor U14924 (N_14924,N_10520,N_9917);
or U14925 (N_14925,N_6966,N_9715);
or U14926 (N_14926,N_10002,N_9837);
nor U14927 (N_14927,N_6543,N_6103);
or U14928 (N_14928,N_10684,N_11895);
xor U14929 (N_14929,N_7955,N_9870);
xor U14930 (N_14930,N_11293,N_8220);
or U14931 (N_14931,N_7228,N_10021);
nand U14932 (N_14932,N_10870,N_11670);
or U14933 (N_14933,N_8185,N_8077);
and U14934 (N_14934,N_8805,N_6750);
nand U14935 (N_14935,N_7949,N_9322);
xnor U14936 (N_14936,N_9337,N_9663);
xnor U14937 (N_14937,N_7013,N_11297);
xnor U14938 (N_14938,N_9976,N_11196);
and U14939 (N_14939,N_6878,N_6682);
and U14940 (N_14940,N_10435,N_10453);
nor U14941 (N_14941,N_6324,N_9415);
nor U14942 (N_14942,N_11182,N_7485);
xor U14943 (N_14943,N_11545,N_10910);
nand U14944 (N_14944,N_7555,N_11482);
nand U14945 (N_14945,N_10523,N_6060);
nand U14946 (N_14946,N_10257,N_7978);
xnor U14947 (N_14947,N_8086,N_10327);
nand U14948 (N_14948,N_6693,N_6968);
xnor U14949 (N_14949,N_9357,N_8863);
nor U14950 (N_14950,N_7591,N_9087);
nor U14951 (N_14951,N_10816,N_6953);
or U14952 (N_14952,N_11629,N_9083);
nor U14953 (N_14953,N_11799,N_6240);
nor U14954 (N_14954,N_8463,N_9524);
xor U14955 (N_14955,N_9975,N_7534);
xnor U14956 (N_14956,N_8461,N_11377);
and U14957 (N_14957,N_6251,N_7263);
nor U14958 (N_14958,N_10622,N_11007);
xor U14959 (N_14959,N_10924,N_10586);
nor U14960 (N_14960,N_7471,N_11614);
nor U14961 (N_14961,N_7766,N_7353);
xor U14962 (N_14962,N_10092,N_6356);
and U14963 (N_14963,N_7159,N_9647);
nor U14964 (N_14964,N_10056,N_11102);
and U14965 (N_14965,N_8592,N_8105);
nand U14966 (N_14966,N_11645,N_9563);
or U14967 (N_14967,N_9536,N_11868);
and U14968 (N_14968,N_8268,N_8589);
xnor U14969 (N_14969,N_11788,N_9896);
and U14970 (N_14970,N_6622,N_6550);
nor U14971 (N_14971,N_8407,N_8327);
or U14972 (N_14972,N_9573,N_9784);
and U14973 (N_14973,N_11591,N_7217);
xnor U14974 (N_14974,N_6230,N_7977);
nor U14975 (N_14975,N_11125,N_11547);
nand U14976 (N_14976,N_11286,N_8130);
and U14977 (N_14977,N_8762,N_8718);
and U14978 (N_14978,N_11290,N_7738);
xor U14979 (N_14979,N_6005,N_8430);
xor U14980 (N_14980,N_8448,N_10259);
nand U14981 (N_14981,N_9543,N_10583);
nor U14982 (N_14982,N_9972,N_11442);
or U14983 (N_14983,N_6098,N_8582);
nand U14984 (N_14984,N_6264,N_6372);
xor U14985 (N_14985,N_8978,N_8553);
and U14986 (N_14986,N_8051,N_11075);
nor U14987 (N_14987,N_10497,N_11477);
or U14988 (N_14988,N_8227,N_8075);
xor U14989 (N_14989,N_6525,N_7544);
nor U14990 (N_14990,N_10188,N_8194);
xor U14991 (N_14991,N_9754,N_7976);
xnor U14992 (N_14992,N_7465,N_11886);
nand U14993 (N_14993,N_8810,N_6326);
nor U14994 (N_14994,N_7606,N_11681);
and U14995 (N_14995,N_11366,N_9809);
or U14996 (N_14996,N_8168,N_11304);
and U14997 (N_14997,N_10255,N_8031);
nor U14998 (N_14998,N_8732,N_8616);
nor U14999 (N_14999,N_8609,N_6422);
nand U15000 (N_15000,N_8453,N_7682);
nor U15001 (N_15001,N_7600,N_8352);
nand U15002 (N_15002,N_6700,N_9750);
nand U15003 (N_15003,N_6379,N_7784);
nand U15004 (N_15004,N_7173,N_6983);
or U15005 (N_15005,N_10437,N_6149);
nand U15006 (N_15006,N_7181,N_10590);
or U15007 (N_15007,N_6192,N_6800);
nor U15008 (N_15008,N_9513,N_10386);
nand U15009 (N_15009,N_8440,N_7168);
nor U15010 (N_15010,N_11579,N_6285);
or U15011 (N_15011,N_7674,N_9668);
or U15012 (N_15012,N_10223,N_11639);
nand U15013 (N_15013,N_10347,N_11016);
and U15014 (N_15014,N_8063,N_6430);
or U15015 (N_15015,N_6703,N_8509);
and U15016 (N_15016,N_10187,N_10443);
and U15017 (N_15017,N_11304,N_7655);
nand U15018 (N_15018,N_9734,N_10262);
nand U15019 (N_15019,N_6781,N_8592);
nor U15020 (N_15020,N_10222,N_10093);
and U15021 (N_15021,N_8650,N_9893);
nor U15022 (N_15022,N_6543,N_11527);
xor U15023 (N_15023,N_6537,N_6004);
or U15024 (N_15024,N_6985,N_6496);
xor U15025 (N_15025,N_8820,N_10767);
and U15026 (N_15026,N_6445,N_8597);
nand U15027 (N_15027,N_8150,N_8156);
or U15028 (N_15028,N_7398,N_11691);
and U15029 (N_15029,N_6807,N_7964);
xor U15030 (N_15030,N_7655,N_7378);
nor U15031 (N_15031,N_11742,N_6237);
and U15032 (N_15032,N_9892,N_6058);
and U15033 (N_15033,N_8467,N_6117);
nor U15034 (N_15034,N_7331,N_10051);
nand U15035 (N_15035,N_9381,N_11034);
nor U15036 (N_15036,N_7025,N_10718);
nand U15037 (N_15037,N_8182,N_8661);
and U15038 (N_15038,N_11315,N_6232);
xor U15039 (N_15039,N_9509,N_11449);
and U15040 (N_15040,N_9808,N_7705);
nor U15041 (N_15041,N_7422,N_9410);
nor U15042 (N_15042,N_8756,N_8022);
or U15043 (N_15043,N_6881,N_7816);
and U15044 (N_15044,N_7654,N_11947);
nand U15045 (N_15045,N_11537,N_7120);
nor U15046 (N_15046,N_11232,N_6207);
xnor U15047 (N_15047,N_11500,N_10881);
nand U15048 (N_15048,N_10913,N_7568);
nor U15049 (N_15049,N_11636,N_7087);
or U15050 (N_15050,N_11261,N_11606);
and U15051 (N_15051,N_7844,N_10750);
or U15052 (N_15052,N_11422,N_8424);
or U15053 (N_15053,N_10438,N_8304);
nand U15054 (N_15054,N_11026,N_7194);
nor U15055 (N_15055,N_7415,N_7671);
xor U15056 (N_15056,N_8645,N_8474);
or U15057 (N_15057,N_10455,N_7075);
and U15058 (N_15058,N_11108,N_6687);
xor U15059 (N_15059,N_6298,N_7779);
nor U15060 (N_15060,N_9005,N_10984);
xor U15061 (N_15061,N_11379,N_6021);
and U15062 (N_15062,N_6343,N_10734);
and U15063 (N_15063,N_6418,N_7537);
and U15064 (N_15064,N_10692,N_9837);
and U15065 (N_15065,N_7449,N_7411);
or U15066 (N_15066,N_9913,N_8441);
nand U15067 (N_15067,N_9917,N_8070);
nor U15068 (N_15068,N_9382,N_9079);
xnor U15069 (N_15069,N_8270,N_7675);
nand U15070 (N_15070,N_11142,N_6364);
xor U15071 (N_15071,N_7679,N_8573);
nand U15072 (N_15072,N_9017,N_10676);
xnor U15073 (N_15073,N_9617,N_7608);
xor U15074 (N_15074,N_9224,N_9678);
or U15075 (N_15075,N_6973,N_7403);
or U15076 (N_15076,N_8397,N_11823);
and U15077 (N_15077,N_10423,N_9460);
or U15078 (N_15078,N_6287,N_10167);
and U15079 (N_15079,N_10956,N_6276);
nand U15080 (N_15080,N_11389,N_11536);
xor U15081 (N_15081,N_7245,N_9435);
xor U15082 (N_15082,N_9347,N_6998);
nor U15083 (N_15083,N_10269,N_8210);
nor U15084 (N_15084,N_7796,N_10809);
nor U15085 (N_15085,N_11952,N_9757);
nand U15086 (N_15086,N_7542,N_9333);
nand U15087 (N_15087,N_11084,N_9488);
and U15088 (N_15088,N_8289,N_7914);
nor U15089 (N_15089,N_6422,N_10163);
nor U15090 (N_15090,N_9369,N_8628);
nand U15091 (N_15091,N_9133,N_6593);
nor U15092 (N_15092,N_9426,N_6963);
xnor U15093 (N_15093,N_8485,N_6169);
xor U15094 (N_15094,N_11154,N_7246);
nor U15095 (N_15095,N_8243,N_11784);
nor U15096 (N_15096,N_9414,N_11445);
nor U15097 (N_15097,N_9436,N_8674);
nor U15098 (N_15098,N_9511,N_10808);
nand U15099 (N_15099,N_11824,N_6954);
nand U15100 (N_15100,N_8842,N_10283);
and U15101 (N_15101,N_9954,N_6176);
nand U15102 (N_15102,N_6026,N_7181);
and U15103 (N_15103,N_7192,N_7674);
nor U15104 (N_15104,N_11467,N_9031);
nor U15105 (N_15105,N_11572,N_6660);
nor U15106 (N_15106,N_10383,N_8372);
nor U15107 (N_15107,N_11552,N_9332);
or U15108 (N_15108,N_9901,N_9804);
nand U15109 (N_15109,N_7050,N_11629);
nand U15110 (N_15110,N_8316,N_9807);
nand U15111 (N_15111,N_6907,N_10657);
or U15112 (N_15112,N_7984,N_10774);
nor U15113 (N_15113,N_9342,N_6385);
or U15114 (N_15114,N_10415,N_11589);
or U15115 (N_15115,N_11826,N_7057);
nand U15116 (N_15116,N_9507,N_11534);
or U15117 (N_15117,N_9187,N_8717);
nand U15118 (N_15118,N_9212,N_7634);
xor U15119 (N_15119,N_7748,N_9400);
nand U15120 (N_15120,N_9115,N_8753);
nor U15121 (N_15121,N_8195,N_11639);
nor U15122 (N_15122,N_10563,N_9887);
and U15123 (N_15123,N_8357,N_9323);
nand U15124 (N_15124,N_9426,N_8080);
or U15125 (N_15125,N_6663,N_9678);
xor U15126 (N_15126,N_9347,N_11050);
xor U15127 (N_15127,N_9791,N_8673);
nand U15128 (N_15128,N_10042,N_10274);
and U15129 (N_15129,N_7788,N_9501);
or U15130 (N_15130,N_7283,N_9828);
nor U15131 (N_15131,N_9834,N_7344);
xor U15132 (N_15132,N_6782,N_11295);
xnor U15133 (N_15133,N_6534,N_10086);
nand U15134 (N_15134,N_8056,N_8213);
and U15135 (N_15135,N_10905,N_9095);
or U15136 (N_15136,N_11926,N_11489);
xor U15137 (N_15137,N_11789,N_7033);
and U15138 (N_15138,N_10054,N_9970);
and U15139 (N_15139,N_11572,N_7034);
or U15140 (N_15140,N_10558,N_6560);
nand U15141 (N_15141,N_10409,N_9516);
or U15142 (N_15142,N_7997,N_7394);
xor U15143 (N_15143,N_8220,N_6322);
nand U15144 (N_15144,N_7278,N_10390);
xnor U15145 (N_15145,N_7309,N_9445);
or U15146 (N_15146,N_6031,N_6231);
nand U15147 (N_15147,N_7271,N_9825);
or U15148 (N_15148,N_7348,N_8474);
or U15149 (N_15149,N_10957,N_6319);
nor U15150 (N_15150,N_10676,N_9823);
xor U15151 (N_15151,N_7145,N_6721);
or U15152 (N_15152,N_7218,N_7359);
or U15153 (N_15153,N_11506,N_6253);
and U15154 (N_15154,N_9172,N_8321);
or U15155 (N_15155,N_8645,N_7419);
xor U15156 (N_15156,N_8133,N_8417);
nand U15157 (N_15157,N_7637,N_9024);
nor U15158 (N_15158,N_9436,N_8918);
or U15159 (N_15159,N_9999,N_10200);
nor U15160 (N_15160,N_6436,N_6426);
nand U15161 (N_15161,N_6257,N_11507);
xor U15162 (N_15162,N_7987,N_10765);
or U15163 (N_15163,N_10056,N_11575);
or U15164 (N_15164,N_9213,N_6962);
and U15165 (N_15165,N_9723,N_11238);
or U15166 (N_15166,N_9975,N_11044);
and U15167 (N_15167,N_7480,N_10742);
and U15168 (N_15168,N_9581,N_8314);
and U15169 (N_15169,N_11412,N_7723);
xor U15170 (N_15170,N_6193,N_10969);
xnor U15171 (N_15171,N_11674,N_10194);
or U15172 (N_15172,N_10402,N_9172);
and U15173 (N_15173,N_7805,N_9397);
xor U15174 (N_15174,N_10241,N_11508);
nor U15175 (N_15175,N_11445,N_11121);
nand U15176 (N_15176,N_8340,N_8041);
xor U15177 (N_15177,N_7118,N_7356);
nor U15178 (N_15178,N_9241,N_10508);
nand U15179 (N_15179,N_7435,N_10045);
nand U15180 (N_15180,N_8627,N_7054);
xor U15181 (N_15181,N_11250,N_8295);
nand U15182 (N_15182,N_7550,N_10703);
xor U15183 (N_15183,N_11985,N_9602);
nand U15184 (N_15184,N_9707,N_10805);
nand U15185 (N_15185,N_9495,N_11302);
nor U15186 (N_15186,N_7228,N_11224);
and U15187 (N_15187,N_7212,N_6819);
or U15188 (N_15188,N_7842,N_9530);
or U15189 (N_15189,N_6175,N_11484);
and U15190 (N_15190,N_6923,N_6343);
and U15191 (N_15191,N_10832,N_10477);
and U15192 (N_15192,N_7865,N_11725);
nor U15193 (N_15193,N_7169,N_7506);
nor U15194 (N_15194,N_7261,N_10351);
nand U15195 (N_15195,N_11110,N_9660);
or U15196 (N_15196,N_10823,N_7174);
nor U15197 (N_15197,N_7288,N_8033);
nor U15198 (N_15198,N_10761,N_9878);
nand U15199 (N_15199,N_6661,N_11077);
xor U15200 (N_15200,N_11049,N_10400);
xnor U15201 (N_15201,N_8616,N_7647);
or U15202 (N_15202,N_10206,N_8310);
nor U15203 (N_15203,N_10499,N_8614);
nor U15204 (N_15204,N_9382,N_8552);
xnor U15205 (N_15205,N_9048,N_9852);
nor U15206 (N_15206,N_7603,N_7911);
and U15207 (N_15207,N_10022,N_11891);
and U15208 (N_15208,N_8734,N_7712);
nor U15209 (N_15209,N_6086,N_8190);
nand U15210 (N_15210,N_10685,N_10853);
or U15211 (N_15211,N_10308,N_8166);
or U15212 (N_15212,N_7690,N_11238);
and U15213 (N_15213,N_7131,N_6934);
nor U15214 (N_15214,N_10018,N_7487);
nand U15215 (N_15215,N_7634,N_6992);
xor U15216 (N_15216,N_8320,N_11047);
nand U15217 (N_15217,N_10286,N_8981);
nor U15218 (N_15218,N_8581,N_9060);
xor U15219 (N_15219,N_11517,N_8676);
nand U15220 (N_15220,N_7571,N_10515);
or U15221 (N_15221,N_6401,N_8623);
nor U15222 (N_15222,N_6285,N_7683);
nor U15223 (N_15223,N_9878,N_7291);
nand U15224 (N_15224,N_7324,N_11801);
xnor U15225 (N_15225,N_11189,N_8242);
nor U15226 (N_15226,N_6746,N_11741);
xor U15227 (N_15227,N_10111,N_8954);
nand U15228 (N_15228,N_9040,N_10207);
and U15229 (N_15229,N_11225,N_11229);
and U15230 (N_15230,N_6445,N_8426);
nand U15231 (N_15231,N_6469,N_8335);
and U15232 (N_15232,N_8060,N_9112);
xor U15233 (N_15233,N_6590,N_11378);
xor U15234 (N_15234,N_11661,N_9767);
nand U15235 (N_15235,N_8330,N_7453);
or U15236 (N_15236,N_7861,N_10275);
and U15237 (N_15237,N_7504,N_8677);
and U15238 (N_15238,N_6473,N_8867);
nor U15239 (N_15239,N_6606,N_8018);
xor U15240 (N_15240,N_10401,N_10658);
xor U15241 (N_15241,N_6197,N_11785);
nor U15242 (N_15242,N_7572,N_7536);
xnor U15243 (N_15243,N_8612,N_10448);
or U15244 (N_15244,N_11350,N_6706);
nand U15245 (N_15245,N_10183,N_10758);
or U15246 (N_15246,N_8514,N_11077);
or U15247 (N_15247,N_7525,N_9951);
xnor U15248 (N_15248,N_8628,N_7806);
or U15249 (N_15249,N_6914,N_7753);
and U15250 (N_15250,N_6618,N_11398);
or U15251 (N_15251,N_6053,N_7469);
nor U15252 (N_15252,N_6891,N_6766);
or U15253 (N_15253,N_11981,N_10945);
or U15254 (N_15254,N_9955,N_9727);
nor U15255 (N_15255,N_7333,N_9720);
nor U15256 (N_15256,N_11491,N_6561);
nor U15257 (N_15257,N_10608,N_9391);
and U15258 (N_15258,N_11016,N_11109);
nand U15259 (N_15259,N_9684,N_7628);
xnor U15260 (N_15260,N_7484,N_7805);
nand U15261 (N_15261,N_9620,N_6231);
xor U15262 (N_15262,N_8838,N_7544);
nand U15263 (N_15263,N_11693,N_7888);
and U15264 (N_15264,N_6454,N_11193);
or U15265 (N_15265,N_7045,N_10536);
nor U15266 (N_15266,N_8172,N_8184);
or U15267 (N_15267,N_10995,N_7127);
xnor U15268 (N_15268,N_10489,N_10575);
xor U15269 (N_15269,N_10640,N_10431);
xnor U15270 (N_15270,N_8420,N_9126);
nor U15271 (N_15271,N_6497,N_11368);
or U15272 (N_15272,N_10908,N_7964);
nor U15273 (N_15273,N_11604,N_6053);
nand U15274 (N_15274,N_10450,N_6939);
and U15275 (N_15275,N_8845,N_11535);
nand U15276 (N_15276,N_7133,N_11493);
and U15277 (N_15277,N_6296,N_10485);
xnor U15278 (N_15278,N_6039,N_7929);
and U15279 (N_15279,N_8230,N_8042);
nand U15280 (N_15280,N_7358,N_8302);
nand U15281 (N_15281,N_10871,N_11418);
nor U15282 (N_15282,N_8382,N_9255);
xnor U15283 (N_15283,N_11413,N_6750);
nor U15284 (N_15284,N_8793,N_7633);
or U15285 (N_15285,N_6403,N_10367);
nand U15286 (N_15286,N_7635,N_11396);
and U15287 (N_15287,N_11070,N_7825);
xor U15288 (N_15288,N_11850,N_10934);
nand U15289 (N_15289,N_11741,N_11665);
nand U15290 (N_15290,N_6261,N_8156);
nand U15291 (N_15291,N_6078,N_11500);
nor U15292 (N_15292,N_11334,N_8778);
and U15293 (N_15293,N_7031,N_6265);
nand U15294 (N_15294,N_7398,N_6640);
xor U15295 (N_15295,N_9122,N_10076);
and U15296 (N_15296,N_11426,N_6316);
and U15297 (N_15297,N_7573,N_10501);
and U15298 (N_15298,N_9511,N_8524);
or U15299 (N_15299,N_9944,N_8527);
and U15300 (N_15300,N_7538,N_9917);
or U15301 (N_15301,N_6830,N_9502);
or U15302 (N_15302,N_7779,N_6883);
nand U15303 (N_15303,N_6843,N_6237);
nor U15304 (N_15304,N_11098,N_8639);
or U15305 (N_15305,N_10741,N_11948);
nand U15306 (N_15306,N_9259,N_7847);
nand U15307 (N_15307,N_11026,N_7056);
xor U15308 (N_15308,N_10772,N_11411);
or U15309 (N_15309,N_6741,N_8960);
nor U15310 (N_15310,N_7355,N_9027);
nand U15311 (N_15311,N_11979,N_11051);
xor U15312 (N_15312,N_8419,N_7134);
and U15313 (N_15313,N_7940,N_10882);
xor U15314 (N_15314,N_10570,N_11927);
xnor U15315 (N_15315,N_9009,N_6425);
nor U15316 (N_15316,N_9578,N_7897);
and U15317 (N_15317,N_6515,N_6683);
xnor U15318 (N_15318,N_11494,N_10473);
nand U15319 (N_15319,N_6243,N_9696);
xnor U15320 (N_15320,N_10557,N_11680);
or U15321 (N_15321,N_11083,N_8753);
nor U15322 (N_15322,N_7639,N_9070);
or U15323 (N_15323,N_8577,N_7180);
nand U15324 (N_15324,N_6538,N_6759);
or U15325 (N_15325,N_11097,N_7635);
or U15326 (N_15326,N_9716,N_11760);
or U15327 (N_15327,N_9242,N_9037);
nor U15328 (N_15328,N_7445,N_11899);
xor U15329 (N_15329,N_10149,N_8164);
and U15330 (N_15330,N_11879,N_11804);
xnor U15331 (N_15331,N_10675,N_8539);
nand U15332 (N_15332,N_11635,N_8698);
nor U15333 (N_15333,N_9988,N_9021);
and U15334 (N_15334,N_9250,N_11050);
or U15335 (N_15335,N_7508,N_9770);
or U15336 (N_15336,N_6409,N_7482);
and U15337 (N_15337,N_6093,N_9824);
xor U15338 (N_15338,N_7501,N_7418);
xor U15339 (N_15339,N_8455,N_6040);
xnor U15340 (N_15340,N_11628,N_6610);
nor U15341 (N_15341,N_8077,N_11212);
or U15342 (N_15342,N_6848,N_7666);
nor U15343 (N_15343,N_8411,N_7025);
nor U15344 (N_15344,N_7066,N_6798);
or U15345 (N_15345,N_6285,N_6302);
nor U15346 (N_15346,N_8917,N_11161);
and U15347 (N_15347,N_10342,N_7365);
nand U15348 (N_15348,N_11455,N_10859);
or U15349 (N_15349,N_9393,N_11601);
and U15350 (N_15350,N_9158,N_6896);
and U15351 (N_15351,N_8124,N_6244);
or U15352 (N_15352,N_11893,N_10393);
nor U15353 (N_15353,N_10523,N_10707);
xnor U15354 (N_15354,N_10082,N_8985);
and U15355 (N_15355,N_11434,N_8644);
xnor U15356 (N_15356,N_10148,N_7837);
xor U15357 (N_15357,N_9670,N_8984);
and U15358 (N_15358,N_11656,N_9792);
or U15359 (N_15359,N_7514,N_10767);
and U15360 (N_15360,N_7297,N_11217);
xor U15361 (N_15361,N_11540,N_7381);
or U15362 (N_15362,N_11026,N_8312);
xnor U15363 (N_15363,N_11916,N_6393);
and U15364 (N_15364,N_9905,N_10117);
and U15365 (N_15365,N_10825,N_7373);
nor U15366 (N_15366,N_11940,N_7634);
nand U15367 (N_15367,N_7891,N_7902);
nor U15368 (N_15368,N_8468,N_7727);
or U15369 (N_15369,N_9131,N_8092);
or U15370 (N_15370,N_8733,N_6903);
nor U15371 (N_15371,N_9668,N_9056);
nor U15372 (N_15372,N_7666,N_11827);
nor U15373 (N_15373,N_11173,N_10251);
or U15374 (N_15374,N_8456,N_10364);
nor U15375 (N_15375,N_10474,N_7798);
or U15376 (N_15376,N_9458,N_6624);
xnor U15377 (N_15377,N_10298,N_7708);
nand U15378 (N_15378,N_8110,N_8261);
nand U15379 (N_15379,N_8460,N_7638);
nand U15380 (N_15380,N_8249,N_11576);
nor U15381 (N_15381,N_7129,N_7657);
or U15382 (N_15382,N_10767,N_10298);
nand U15383 (N_15383,N_7451,N_8019);
nand U15384 (N_15384,N_11199,N_8031);
and U15385 (N_15385,N_10645,N_9115);
and U15386 (N_15386,N_7806,N_6724);
or U15387 (N_15387,N_11936,N_8621);
and U15388 (N_15388,N_7636,N_6975);
nand U15389 (N_15389,N_6703,N_11857);
nand U15390 (N_15390,N_9064,N_10413);
xnor U15391 (N_15391,N_11546,N_8197);
nor U15392 (N_15392,N_6169,N_9459);
nand U15393 (N_15393,N_11385,N_10252);
nand U15394 (N_15394,N_7789,N_10072);
xnor U15395 (N_15395,N_9107,N_10236);
or U15396 (N_15396,N_11738,N_6483);
xor U15397 (N_15397,N_11968,N_11761);
or U15398 (N_15398,N_10138,N_10418);
nor U15399 (N_15399,N_9655,N_7200);
and U15400 (N_15400,N_11671,N_6118);
or U15401 (N_15401,N_8419,N_8742);
nand U15402 (N_15402,N_10477,N_7315);
and U15403 (N_15403,N_10453,N_9261);
nand U15404 (N_15404,N_7580,N_11463);
nor U15405 (N_15405,N_8092,N_8667);
and U15406 (N_15406,N_7094,N_7617);
and U15407 (N_15407,N_8759,N_10529);
xnor U15408 (N_15408,N_10206,N_8229);
xor U15409 (N_15409,N_11298,N_7498);
nand U15410 (N_15410,N_7896,N_9934);
or U15411 (N_15411,N_8641,N_10731);
and U15412 (N_15412,N_6936,N_9533);
or U15413 (N_15413,N_7794,N_8129);
and U15414 (N_15414,N_6976,N_7496);
and U15415 (N_15415,N_9544,N_7368);
nor U15416 (N_15416,N_11035,N_11764);
nand U15417 (N_15417,N_9700,N_6070);
nand U15418 (N_15418,N_10153,N_11602);
nand U15419 (N_15419,N_6345,N_6083);
and U15420 (N_15420,N_11331,N_10292);
nor U15421 (N_15421,N_9380,N_8222);
xor U15422 (N_15422,N_10525,N_8472);
nand U15423 (N_15423,N_7910,N_6844);
xor U15424 (N_15424,N_8420,N_8092);
or U15425 (N_15425,N_6681,N_8847);
nand U15426 (N_15426,N_9595,N_6360);
xnor U15427 (N_15427,N_8427,N_6670);
nand U15428 (N_15428,N_6919,N_7110);
and U15429 (N_15429,N_11349,N_11994);
xnor U15430 (N_15430,N_9899,N_6421);
nor U15431 (N_15431,N_8186,N_9895);
and U15432 (N_15432,N_8590,N_7097);
or U15433 (N_15433,N_11437,N_10197);
or U15434 (N_15434,N_10032,N_8634);
xnor U15435 (N_15435,N_7105,N_10028);
nand U15436 (N_15436,N_9797,N_7329);
nor U15437 (N_15437,N_10639,N_9037);
xor U15438 (N_15438,N_10174,N_11739);
or U15439 (N_15439,N_8301,N_10444);
nor U15440 (N_15440,N_11632,N_8222);
and U15441 (N_15441,N_8163,N_7227);
and U15442 (N_15442,N_11853,N_9351);
xnor U15443 (N_15443,N_8377,N_8869);
nand U15444 (N_15444,N_7882,N_11926);
xor U15445 (N_15445,N_7683,N_11683);
xnor U15446 (N_15446,N_6156,N_10204);
or U15447 (N_15447,N_7054,N_10260);
xnor U15448 (N_15448,N_9767,N_9090);
nor U15449 (N_15449,N_9961,N_10649);
nand U15450 (N_15450,N_10341,N_11465);
nand U15451 (N_15451,N_7181,N_8679);
xnor U15452 (N_15452,N_6577,N_7201);
nor U15453 (N_15453,N_10450,N_7091);
or U15454 (N_15454,N_11505,N_8101);
or U15455 (N_15455,N_11192,N_7298);
and U15456 (N_15456,N_7875,N_10766);
and U15457 (N_15457,N_11741,N_7274);
nand U15458 (N_15458,N_9928,N_9429);
and U15459 (N_15459,N_7827,N_9561);
or U15460 (N_15460,N_9904,N_10291);
nand U15461 (N_15461,N_11593,N_8965);
xor U15462 (N_15462,N_10281,N_7705);
and U15463 (N_15463,N_8099,N_11514);
nor U15464 (N_15464,N_6729,N_11699);
nor U15465 (N_15465,N_7550,N_11510);
and U15466 (N_15466,N_9563,N_10719);
nand U15467 (N_15467,N_8239,N_6379);
xnor U15468 (N_15468,N_7096,N_8733);
xnor U15469 (N_15469,N_7903,N_6884);
and U15470 (N_15470,N_7503,N_11107);
nor U15471 (N_15471,N_8752,N_8797);
and U15472 (N_15472,N_10855,N_7345);
nor U15473 (N_15473,N_7346,N_8168);
xor U15474 (N_15474,N_10262,N_7740);
and U15475 (N_15475,N_11184,N_11971);
xor U15476 (N_15476,N_11696,N_9370);
xnor U15477 (N_15477,N_6885,N_8361);
nor U15478 (N_15478,N_11074,N_11394);
nor U15479 (N_15479,N_8961,N_6867);
nor U15480 (N_15480,N_11359,N_6428);
nand U15481 (N_15481,N_6324,N_7394);
xor U15482 (N_15482,N_8264,N_10972);
xnor U15483 (N_15483,N_11111,N_6495);
nand U15484 (N_15484,N_6954,N_7956);
or U15485 (N_15485,N_8143,N_10065);
or U15486 (N_15486,N_7355,N_9174);
nor U15487 (N_15487,N_11394,N_6189);
and U15488 (N_15488,N_6094,N_6581);
xnor U15489 (N_15489,N_7615,N_6663);
or U15490 (N_15490,N_6020,N_6240);
xor U15491 (N_15491,N_9328,N_11379);
xor U15492 (N_15492,N_10565,N_10471);
and U15493 (N_15493,N_8535,N_11400);
and U15494 (N_15494,N_8761,N_11243);
xnor U15495 (N_15495,N_6380,N_9223);
nand U15496 (N_15496,N_11007,N_8729);
nand U15497 (N_15497,N_6397,N_10457);
and U15498 (N_15498,N_10492,N_11624);
nor U15499 (N_15499,N_7999,N_6022);
nor U15500 (N_15500,N_9512,N_9889);
and U15501 (N_15501,N_6116,N_7201);
or U15502 (N_15502,N_6820,N_6520);
nand U15503 (N_15503,N_7478,N_7632);
and U15504 (N_15504,N_9198,N_10419);
nor U15505 (N_15505,N_10543,N_11158);
xnor U15506 (N_15506,N_8004,N_6023);
or U15507 (N_15507,N_7490,N_6182);
or U15508 (N_15508,N_9324,N_9830);
and U15509 (N_15509,N_6342,N_6049);
xor U15510 (N_15510,N_6598,N_7084);
nand U15511 (N_15511,N_8113,N_8656);
xor U15512 (N_15512,N_11327,N_7721);
nand U15513 (N_15513,N_7111,N_7661);
or U15514 (N_15514,N_10084,N_6528);
nand U15515 (N_15515,N_8592,N_9494);
and U15516 (N_15516,N_8887,N_8396);
and U15517 (N_15517,N_8393,N_10384);
nor U15518 (N_15518,N_8418,N_10833);
or U15519 (N_15519,N_6248,N_9975);
xnor U15520 (N_15520,N_10320,N_11784);
nor U15521 (N_15521,N_9572,N_9496);
xor U15522 (N_15522,N_6180,N_10055);
xor U15523 (N_15523,N_6643,N_10134);
nand U15524 (N_15524,N_9267,N_9960);
or U15525 (N_15525,N_11100,N_8100);
or U15526 (N_15526,N_9987,N_11414);
and U15527 (N_15527,N_8797,N_11612);
nand U15528 (N_15528,N_6496,N_9114);
nor U15529 (N_15529,N_9270,N_9847);
or U15530 (N_15530,N_10840,N_11714);
xor U15531 (N_15531,N_9760,N_10144);
or U15532 (N_15532,N_10904,N_10974);
nand U15533 (N_15533,N_9867,N_7549);
or U15534 (N_15534,N_11486,N_11916);
nand U15535 (N_15535,N_8534,N_6463);
nor U15536 (N_15536,N_6395,N_10640);
nor U15537 (N_15537,N_7320,N_9135);
nand U15538 (N_15538,N_7441,N_6636);
nor U15539 (N_15539,N_8870,N_8092);
and U15540 (N_15540,N_9469,N_8850);
and U15541 (N_15541,N_11922,N_10488);
xnor U15542 (N_15542,N_10186,N_9054);
nand U15543 (N_15543,N_10737,N_10759);
nand U15544 (N_15544,N_6721,N_8939);
nand U15545 (N_15545,N_6690,N_10009);
and U15546 (N_15546,N_8028,N_9596);
nor U15547 (N_15547,N_8409,N_9763);
and U15548 (N_15548,N_11995,N_7448);
and U15549 (N_15549,N_10774,N_11984);
or U15550 (N_15550,N_6190,N_6736);
xor U15551 (N_15551,N_11750,N_8472);
nand U15552 (N_15552,N_8373,N_8706);
nand U15553 (N_15553,N_9353,N_8473);
or U15554 (N_15554,N_7565,N_11285);
xnor U15555 (N_15555,N_7070,N_11347);
and U15556 (N_15556,N_10108,N_8049);
and U15557 (N_15557,N_10086,N_8477);
nand U15558 (N_15558,N_11392,N_11619);
and U15559 (N_15559,N_7279,N_11096);
xor U15560 (N_15560,N_9213,N_8390);
nor U15561 (N_15561,N_10582,N_8829);
xnor U15562 (N_15562,N_10199,N_10357);
nor U15563 (N_15563,N_7563,N_10487);
nand U15564 (N_15564,N_6706,N_10860);
nor U15565 (N_15565,N_11703,N_7641);
xnor U15566 (N_15566,N_6881,N_10695);
nand U15567 (N_15567,N_6289,N_11274);
xnor U15568 (N_15568,N_11744,N_8014);
and U15569 (N_15569,N_9815,N_6944);
or U15570 (N_15570,N_6261,N_10918);
or U15571 (N_15571,N_10213,N_10615);
xor U15572 (N_15572,N_9583,N_6103);
nand U15573 (N_15573,N_10825,N_8896);
xnor U15574 (N_15574,N_9293,N_10196);
nor U15575 (N_15575,N_11558,N_6081);
and U15576 (N_15576,N_7837,N_11251);
nand U15577 (N_15577,N_6066,N_8934);
or U15578 (N_15578,N_7868,N_9929);
and U15579 (N_15579,N_8976,N_7672);
and U15580 (N_15580,N_10563,N_6005);
or U15581 (N_15581,N_6206,N_9230);
and U15582 (N_15582,N_8157,N_8650);
and U15583 (N_15583,N_6820,N_9726);
or U15584 (N_15584,N_11508,N_8501);
and U15585 (N_15585,N_6159,N_6487);
nand U15586 (N_15586,N_6539,N_8616);
or U15587 (N_15587,N_6921,N_6004);
or U15588 (N_15588,N_7752,N_8914);
nand U15589 (N_15589,N_7190,N_8611);
or U15590 (N_15590,N_7088,N_7707);
nor U15591 (N_15591,N_7147,N_10612);
nand U15592 (N_15592,N_11334,N_8225);
xor U15593 (N_15593,N_6840,N_9680);
xnor U15594 (N_15594,N_9251,N_8790);
and U15595 (N_15595,N_9752,N_10611);
nor U15596 (N_15596,N_10661,N_9614);
and U15597 (N_15597,N_11579,N_6015);
and U15598 (N_15598,N_6798,N_11810);
and U15599 (N_15599,N_8159,N_6372);
xor U15600 (N_15600,N_7156,N_7173);
and U15601 (N_15601,N_11398,N_8314);
xor U15602 (N_15602,N_9650,N_7372);
or U15603 (N_15603,N_6161,N_6631);
and U15604 (N_15604,N_8624,N_8017);
nor U15605 (N_15605,N_7328,N_9961);
xor U15606 (N_15606,N_8189,N_7613);
nor U15607 (N_15607,N_6555,N_8184);
xnor U15608 (N_15608,N_11300,N_8758);
nand U15609 (N_15609,N_9979,N_7278);
and U15610 (N_15610,N_11914,N_6995);
and U15611 (N_15611,N_6725,N_9323);
and U15612 (N_15612,N_8901,N_6126);
nand U15613 (N_15613,N_10595,N_8811);
or U15614 (N_15614,N_11123,N_8943);
nor U15615 (N_15615,N_8447,N_9726);
or U15616 (N_15616,N_6085,N_11417);
nand U15617 (N_15617,N_10787,N_8506);
xnor U15618 (N_15618,N_7783,N_11130);
or U15619 (N_15619,N_6878,N_10940);
nor U15620 (N_15620,N_6563,N_11096);
nand U15621 (N_15621,N_8488,N_7144);
and U15622 (N_15622,N_11454,N_9311);
nor U15623 (N_15623,N_11081,N_9927);
nand U15624 (N_15624,N_9278,N_11206);
or U15625 (N_15625,N_8572,N_11498);
and U15626 (N_15626,N_8172,N_6985);
nor U15627 (N_15627,N_11161,N_11848);
nor U15628 (N_15628,N_11312,N_8625);
nand U15629 (N_15629,N_9420,N_7510);
nand U15630 (N_15630,N_11047,N_11259);
nand U15631 (N_15631,N_10942,N_10937);
and U15632 (N_15632,N_8173,N_9699);
and U15633 (N_15633,N_10827,N_6325);
nor U15634 (N_15634,N_6702,N_6654);
nand U15635 (N_15635,N_7045,N_10973);
or U15636 (N_15636,N_11846,N_10208);
or U15637 (N_15637,N_8162,N_9331);
xnor U15638 (N_15638,N_10885,N_10654);
and U15639 (N_15639,N_10922,N_9480);
xor U15640 (N_15640,N_11777,N_9251);
nor U15641 (N_15641,N_8276,N_9391);
and U15642 (N_15642,N_9712,N_8782);
nand U15643 (N_15643,N_10398,N_7115);
and U15644 (N_15644,N_9784,N_6419);
or U15645 (N_15645,N_6893,N_6869);
or U15646 (N_15646,N_7131,N_6629);
and U15647 (N_15647,N_9260,N_6594);
xnor U15648 (N_15648,N_11793,N_9418);
and U15649 (N_15649,N_8431,N_8183);
xor U15650 (N_15650,N_11968,N_7136);
and U15651 (N_15651,N_10440,N_10325);
and U15652 (N_15652,N_6392,N_6475);
and U15653 (N_15653,N_10313,N_8319);
nor U15654 (N_15654,N_11841,N_8176);
and U15655 (N_15655,N_7377,N_10045);
nor U15656 (N_15656,N_11131,N_7269);
nor U15657 (N_15657,N_9810,N_11371);
nand U15658 (N_15658,N_9181,N_7359);
nand U15659 (N_15659,N_9834,N_10046);
or U15660 (N_15660,N_11847,N_8640);
xor U15661 (N_15661,N_9880,N_6546);
xnor U15662 (N_15662,N_9052,N_9748);
nor U15663 (N_15663,N_9359,N_7115);
xor U15664 (N_15664,N_6777,N_6669);
or U15665 (N_15665,N_6382,N_7173);
nand U15666 (N_15666,N_8805,N_11201);
nand U15667 (N_15667,N_6983,N_10002);
xor U15668 (N_15668,N_6584,N_8950);
and U15669 (N_15669,N_11657,N_7490);
xor U15670 (N_15670,N_10069,N_7899);
nor U15671 (N_15671,N_9827,N_11297);
or U15672 (N_15672,N_9555,N_6619);
xnor U15673 (N_15673,N_9653,N_7992);
and U15674 (N_15674,N_6149,N_7944);
or U15675 (N_15675,N_10028,N_10470);
nand U15676 (N_15676,N_8716,N_6087);
and U15677 (N_15677,N_11488,N_6777);
xnor U15678 (N_15678,N_6329,N_10224);
and U15679 (N_15679,N_11769,N_9987);
nand U15680 (N_15680,N_11908,N_6737);
xnor U15681 (N_15681,N_9275,N_10249);
and U15682 (N_15682,N_8465,N_8110);
nor U15683 (N_15683,N_8400,N_11616);
xor U15684 (N_15684,N_6641,N_10721);
nor U15685 (N_15685,N_11822,N_8071);
nand U15686 (N_15686,N_11508,N_8710);
or U15687 (N_15687,N_10523,N_7519);
and U15688 (N_15688,N_11492,N_8279);
nor U15689 (N_15689,N_6322,N_11270);
and U15690 (N_15690,N_9416,N_6618);
or U15691 (N_15691,N_7396,N_6493);
xnor U15692 (N_15692,N_10688,N_6672);
or U15693 (N_15693,N_11291,N_10034);
and U15694 (N_15694,N_11506,N_9997);
xor U15695 (N_15695,N_11064,N_8782);
or U15696 (N_15696,N_8422,N_7809);
nand U15697 (N_15697,N_9752,N_8000);
nor U15698 (N_15698,N_10995,N_10544);
nor U15699 (N_15699,N_7061,N_6739);
and U15700 (N_15700,N_9929,N_9705);
or U15701 (N_15701,N_7062,N_10274);
and U15702 (N_15702,N_11860,N_9744);
xnor U15703 (N_15703,N_7965,N_10934);
or U15704 (N_15704,N_9934,N_9486);
xnor U15705 (N_15705,N_9612,N_7294);
nor U15706 (N_15706,N_7044,N_11230);
or U15707 (N_15707,N_6785,N_10625);
or U15708 (N_15708,N_11525,N_11199);
and U15709 (N_15709,N_11164,N_9671);
nand U15710 (N_15710,N_11377,N_6790);
nor U15711 (N_15711,N_7389,N_10017);
or U15712 (N_15712,N_7853,N_8997);
xnor U15713 (N_15713,N_10655,N_7245);
nand U15714 (N_15714,N_9344,N_6353);
or U15715 (N_15715,N_10629,N_6286);
nor U15716 (N_15716,N_8860,N_8937);
xor U15717 (N_15717,N_8991,N_11284);
nor U15718 (N_15718,N_11989,N_10313);
nor U15719 (N_15719,N_7473,N_6495);
nor U15720 (N_15720,N_8484,N_10140);
nand U15721 (N_15721,N_10085,N_8807);
xor U15722 (N_15722,N_11057,N_11799);
xnor U15723 (N_15723,N_6711,N_9409);
xor U15724 (N_15724,N_8060,N_7562);
and U15725 (N_15725,N_6752,N_9657);
or U15726 (N_15726,N_9178,N_7825);
or U15727 (N_15727,N_10353,N_7798);
nand U15728 (N_15728,N_10637,N_9239);
xnor U15729 (N_15729,N_7682,N_8752);
or U15730 (N_15730,N_9040,N_10293);
or U15731 (N_15731,N_7658,N_9831);
or U15732 (N_15732,N_11557,N_8109);
nor U15733 (N_15733,N_6076,N_6045);
and U15734 (N_15734,N_7793,N_8971);
nor U15735 (N_15735,N_8621,N_9831);
nor U15736 (N_15736,N_8365,N_8136);
and U15737 (N_15737,N_11381,N_8480);
xnor U15738 (N_15738,N_8538,N_9765);
or U15739 (N_15739,N_11934,N_11930);
xor U15740 (N_15740,N_6885,N_11688);
nand U15741 (N_15741,N_9353,N_11575);
nor U15742 (N_15742,N_10304,N_9110);
nand U15743 (N_15743,N_10146,N_9453);
xnor U15744 (N_15744,N_10572,N_11947);
or U15745 (N_15745,N_6131,N_8928);
or U15746 (N_15746,N_10889,N_8055);
and U15747 (N_15747,N_8044,N_7674);
nor U15748 (N_15748,N_10721,N_6578);
or U15749 (N_15749,N_9380,N_6022);
nor U15750 (N_15750,N_11072,N_8508);
nand U15751 (N_15751,N_9953,N_6422);
nor U15752 (N_15752,N_9854,N_7443);
nand U15753 (N_15753,N_8694,N_7812);
or U15754 (N_15754,N_7658,N_11260);
and U15755 (N_15755,N_8323,N_8715);
or U15756 (N_15756,N_7536,N_9246);
or U15757 (N_15757,N_8744,N_7781);
or U15758 (N_15758,N_9220,N_10934);
and U15759 (N_15759,N_9012,N_9325);
xor U15760 (N_15760,N_10178,N_10091);
and U15761 (N_15761,N_8260,N_8134);
xor U15762 (N_15762,N_8666,N_9185);
xnor U15763 (N_15763,N_10118,N_10380);
nor U15764 (N_15764,N_9508,N_11741);
or U15765 (N_15765,N_11542,N_10825);
and U15766 (N_15766,N_9137,N_7625);
and U15767 (N_15767,N_7133,N_8330);
and U15768 (N_15768,N_7845,N_8673);
nand U15769 (N_15769,N_8889,N_8281);
xor U15770 (N_15770,N_7937,N_7819);
nor U15771 (N_15771,N_8075,N_10278);
xnor U15772 (N_15772,N_8388,N_8629);
nor U15773 (N_15773,N_11196,N_9099);
or U15774 (N_15774,N_6527,N_11100);
nand U15775 (N_15775,N_11250,N_6661);
or U15776 (N_15776,N_10238,N_9149);
or U15777 (N_15777,N_9674,N_11789);
nor U15778 (N_15778,N_9326,N_10029);
and U15779 (N_15779,N_11419,N_7214);
nand U15780 (N_15780,N_10059,N_10306);
xor U15781 (N_15781,N_10934,N_8388);
or U15782 (N_15782,N_6246,N_7902);
and U15783 (N_15783,N_7267,N_10531);
or U15784 (N_15784,N_6310,N_8662);
or U15785 (N_15785,N_10548,N_6269);
or U15786 (N_15786,N_10845,N_10074);
xor U15787 (N_15787,N_11404,N_7105);
and U15788 (N_15788,N_10145,N_8154);
and U15789 (N_15789,N_8157,N_11181);
nand U15790 (N_15790,N_8705,N_8423);
and U15791 (N_15791,N_8006,N_8527);
or U15792 (N_15792,N_8405,N_9153);
nand U15793 (N_15793,N_9782,N_10820);
and U15794 (N_15794,N_6560,N_6829);
and U15795 (N_15795,N_9015,N_8627);
nand U15796 (N_15796,N_6307,N_11755);
xor U15797 (N_15797,N_10175,N_9485);
xor U15798 (N_15798,N_8804,N_6836);
xor U15799 (N_15799,N_10719,N_7305);
or U15800 (N_15800,N_8076,N_9897);
nor U15801 (N_15801,N_8511,N_9516);
and U15802 (N_15802,N_11045,N_9119);
xnor U15803 (N_15803,N_7549,N_7538);
and U15804 (N_15804,N_11695,N_6055);
nand U15805 (N_15805,N_6802,N_7344);
and U15806 (N_15806,N_7234,N_7503);
nand U15807 (N_15807,N_8434,N_8943);
xor U15808 (N_15808,N_7560,N_9385);
and U15809 (N_15809,N_6726,N_9510);
and U15810 (N_15810,N_7135,N_11211);
nor U15811 (N_15811,N_6252,N_7692);
nand U15812 (N_15812,N_11174,N_8053);
xnor U15813 (N_15813,N_7482,N_6988);
nor U15814 (N_15814,N_6991,N_7485);
or U15815 (N_15815,N_7244,N_9747);
and U15816 (N_15816,N_9794,N_10570);
or U15817 (N_15817,N_10214,N_7190);
or U15818 (N_15818,N_9998,N_11739);
xnor U15819 (N_15819,N_11877,N_6008);
xor U15820 (N_15820,N_7317,N_6038);
xnor U15821 (N_15821,N_7159,N_8903);
xnor U15822 (N_15822,N_7776,N_7233);
nand U15823 (N_15823,N_7204,N_9291);
xnor U15824 (N_15824,N_6072,N_7567);
xor U15825 (N_15825,N_10627,N_7120);
nor U15826 (N_15826,N_8141,N_7179);
nor U15827 (N_15827,N_8835,N_7535);
xnor U15828 (N_15828,N_7144,N_10595);
nor U15829 (N_15829,N_6683,N_6814);
and U15830 (N_15830,N_7202,N_11436);
xor U15831 (N_15831,N_6315,N_8250);
xnor U15832 (N_15832,N_7533,N_9512);
nor U15833 (N_15833,N_10317,N_6946);
or U15834 (N_15834,N_11330,N_7819);
nor U15835 (N_15835,N_6081,N_6490);
or U15836 (N_15836,N_7508,N_11330);
and U15837 (N_15837,N_11676,N_8443);
nor U15838 (N_15838,N_10945,N_10295);
nor U15839 (N_15839,N_10420,N_6535);
xnor U15840 (N_15840,N_9583,N_9283);
xor U15841 (N_15841,N_8729,N_11627);
and U15842 (N_15842,N_9441,N_10145);
nand U15843 (N_15843,N_10399,N_10392);
and U15844 (N_15844,N_9007,N_11866);
nand U15845 (N_15845,N_7398,N_10639);
or U15846 (N_15846,N_11138,N_10634);
or U15847 (N_15847,N_8059,N_7394);
nand U15848 (N_15848,N_9314,N_8698);
nor U15849 (N_15849,N_6726,N_6576);
nor U15850 (N_15850,N_8662,N_6933);
nor U15851 (N_15851,N_11550,N_6404);
nor U15852 (N_15852,N_9130,N_11011);
and U15853 (N_15853,N_11060,N_7873);
or U15854 (N_15854,N_6802,N_6673);
or U15855 (N_15855,N_8236,N_10960);
and U15856 (N_15856,N_7573,N_9867);
and U15857 (N_15857,N_6404,N_11872);
xnor U15858 (N_15858,N_11413,N_8347);
nand U15859 (N_15859,N_10409,N_6517);
or U15860 (N_15860,N_9728,N_6621);
nor U15861 (N_15861,N_9918,N_6846);
or U15862 (N_15862,N_6341,N_10845);
nand U15863 (N_15863,N_11337,N_7125);
and U15864 (N_15864,N_11379,N_8607);
nand U15865 (N_15865,N_11712,N_9733);
and U15866 (N_15866,N_9526,N_7281);
or U15867 (N_15867,N_6217,N_9996);
or U15868 (N_15868,N_7345,N_11926);
nand U15869 (N_15869,N_8598,N_11973);
nor U15870 (N_15870,N_11223,N_9626);
and U15871 (N_15871,N_9148,N_11148);
and U15872 (N_15872,N_6936,N_7068);
xnor U15873 (N_15873,N_6204,N_6796);
or U15874 (N_15874,N_11426,N_9873);
nor U15875 (N_15875,N_7258,N_9460);
nand U15876 (N_15876,N_6273,N_10613);
nand U15877 (N_15877,N_9093,N_8239);
and U15878 (N_15878,N_10502,N_10632);
xor U15879 (N_15879,N_8467,N_7607);
nor U15880 (N_15880,N_7079,N_7747);
nand U15881 (N_15881,N_8691,N_6344);
nand U15882 (N_15882,N_8403,N_8468);
nor U15883 (N_15883,N_8761,N_9359);
or U15884 (N_15884,N_7835,N_6425);
nor U15885 (N_15885,N_7177,N_7335);
or U15886 (N_15886,N_8863,N_9444);
nor U15887 (N_15887,N_11620,N_11677);
nor U15888 (N_15888,N_10307,N_8733);
xnor U15889 (N_15889,N_6563,N_8517);
or U15890 (N_15890,N_7560,N_6359);
nor U15891 (N_15891,N_8710,N_10465);
xor U15892 (N_15892,N_10964,N_6051);
nor U15893 (N_15893,N_7339,N_6179);
xnor U15894 (N_15894,N_11264,N_9871);
nand U15895 (N_15895,N_8675,N_8249);
or U15896 (N_15896,N_6938,N_10555);
nor U15897 (N_15897,N_10625,N_6128);
or U15898 (N_15898,N_6661,N_11221);
or U15899 (N_15899,N_8900,N_9720);
and U15900 (N_15900,N_9252,N_6972);
nand U15901 (N_15901,N_6269,N_9484);
xor U15902 (N_15902,N_8103,N_11990);
and U15903 (N_15903,N_8501,N_7255);
or U15904 (N_15904,N_7135,N_10337);
nor U15905 (N_15905,N_8766,N_11785);
nor U15906 (N_15906,N_9947,N_11676);
nand U15907 (N_15907,N_7238,N_8368);
or U15908 (N_15908,N_6835,N_10007);
nor U15909 (N_15909,N_11516,N_10988);
nor U15910 (N_15910,N_10930,N_7484);
nor U15911 (N_15911,N_6846,N_8662);
and U15912 (N_15912,N_11992,N_10631);
or U15913 (N_15913,N_10760,N_6984);
nand U15914 (N_15914,N_11227,N_7794);
nand U15915 (N_15915,N_10491,N_9703);
nand U15916 (N_15916,N_7604,N_6196);
and U15917 (N_15917,N_9976,N_6246);
nor U15918 (N_15918,N_8172,N_8656);
xor U15919 (N_15919,N_6422,N_7764);
and U15920 (N_15920,N_6117,N_8318);
nand U15921 (N_15921,N_7694,N_8477);
and U15922 (N_15922,N_10369,N_6045);
xnor U15923 (N_15923,N_8388,N_7118);
nand U15924 (N_15924,N_11166,N_11942);
nand U15925 (N_15925,N_11874,N_10883);
and U15926 (N_15926,N_9330,N_9307);
and U15927 (N_15927,N_9290,N_7969);
nand U15928 (N_15928,N_6734,N_8718);
nand U15929 (N_15929,N_8554,N_8778);
nand U15930 (N_15930,N_9733,N_6353);
nand U15931 (N_15931,N_9213,N_9945);
nor U15932 (N_15932,N_8954,N_9836);
xor U15933 (N_15933,N_11551,N_10127);
and U15934 (N_15934,N_7589,N_6063);
nor U15935 (N_15935,N_6044,N_6575);
nor U15936 (N_15936,N_6221,N_7619);
nor U15937 (N_15937,N_11653,N_8656);
nand U15938 (N_15938,N_7430,N_9433);
xor U15939 (N_15939,N_8847,N_10263);
and U15940 (N_15940,N_7298,N_10265);
and U15941 (N_15941,N_8863,N_10491);
xor U15942 (N_15942,N_10565,N_8331);
and U15943 (N_15943,N_11071,N_11070);
nor U15944 (N_15944,N_10860,N_7074);
xor U15945 (N_15945,N_11409,N_6015);
xnor U15946 (N_15946,N_10744,N_11796);
nor U15947 (N_15947,N_11732,N_9864);
nor U15948 (N_15948,N_10558,N_8519);
nand U15949 (N_15949,N_7400,N_8244);
and U15950 (N_15950,N_7056,N_7136);
nor U15951 (N_15951,N_7468,N_6780);
or U15952 (N_15952,N_8869,N_8598);
nand U15953 (N_15953,N_10457,N_10531);
or U15954 (N_15954,N_8584,N_11486);
xor U15955 (N_15955,N_9537,N_9109);
or U15956 (N_15956,N_6615,N_8075);
or U15957 (N_15957,N_8251,N_6568);
xor U15958 (N_15958,N_11229,N_10918);
nor U15959 (N_15959,N_10339,N_10331);
or U15960 (N_15960,N_8627,N_6885);
and U15961 (N_15961,N_6565,N_6748);
and U15962 (N_15962,N_7343,N_11445);
nand U15963 (N_15963,N_11407,N_6494);
nand U15964 (N_15964,N_11926,N_7468);
nand U15965 (N_15965,N_11837,N_9018);
or U15966 (N_15966,N_6202,N_7468);
nand U15967 (N_15967,N_8683,N_6784);
nor U15968 (N_15968,N_11358,N_10868);
and U15969 (N_15969,N_7983,N_10818);
xnor U15970 (N_15970,N_7877,N_8558);
nand U15971 (N_15971,N_11643,N_9972);
nor U15972 (N_15972,N_6558,N_9173);
or U15973 (N_15973,N_10068,N_6316);
or U15974 (N_15974,N_10174,N_8823);
nand U15975 (N_15975,N_11876,N_11830);
nor U15976 (N_15976,N_6449,N_6524);
nand U15977 (N_15977,N_11584,N_10316);
and U15978 (N_15978,N_10030,N_6236);
xor U15979 (N_15979,N_11493,N_11596);
nand U15980 (N_15980,N_6142,N_8076);
nor U15981 (N_15981,N_7053,N_8586);
nand U15982 (N_15982,N_8407,N_8822);
nand U15983 (N_15983,N_8087,N_8795);
nand U15984 (N_15984,N_11246,N_10747);
xnor U15985 (N_15985,N_9372,N_7738);
xnor U15986 (N_15986,N_10893,N_7220);
and U15987 (N_15987,N_11273,N_10318);
xnor U15988 (N_15988,N_11996,N_8049);
and U15989 (N_15989,N_11245,N_10408);
xnor U15990 (N_15990,N_11512,N_10614);
nor U15991 (N_15991,N_9167,N_11228);
xnor U15992 (N_15992,N_10113,N_8206);
nor U15993 (N_15993,N_11675,N_8480);
and U15994 (N_15994,N_11868,N_10842);
nor U15995 (N_15995,N_9782,N_6998);
or U15996 (N_15996,N_10812,N_10603);
nand U15997 (N_15997,N_10579,N_8966);
and U15998 (N_15998,N_9512,N_10173);
and U15999 (N_15999,N_11019,N_11446);
or U16000 (N_16000,N_8097,N_11880);
or U16001 (N_16001,N_9259,N_7768);
and U16002 (N_16002,N_7307,N_8891);
and U16003 (N_16003,N_8496,N_11785);
and U16004 (N_16004,N_9306,N_7224);
and U16005 (N_16005,N_10718,N_10966);
nor U16006 (N_16006,N_9114,N_10392);
nor U16007 (N_16007,N_11581,N_8216);
xnor U16008 (N_16008,N_11363,N_11430);
nand U16009 (N_16009,N_9559,N_10793);
and U16010 (N_16010,N_6031,N_10538);
nand U16011 (N_16011,N_9511,N_11575);
or U16012 (N_16012,N_10872,N_6892);
nor U16013 (N_16013,N_9226,N_8932);
nand U16014 (N_16014,N_7993,N_10234);
nand U16015 (N_16015,N_11056,N_10148);
nand U16016 (N_16016,N_7800,N_7824);
nor U16017 (N_16017,N_7033,N_11299);
and U16018 (N_16018,N_8067,N_7000);
nand U16019 (N_16019,N_7324,N_7201);
or U16020 (N_16020,N_6165,N_10283);
nand U16021 (N_16021,N_10074,N_11280);
nand U16022 (N_16022,N_6939,N_9440);
nand U16023 (N_16023,N_10254,N_9552);
and U16024 (N_16024,N_11416,N_10708);
or U16025 (N_16025,N_9591,N_11080);
or U16026 (N_16026,N_9412,N_7231);
or U16027 (N_16027,N_9137,N_7106);
or U16028 (N_16028,N_7833,N_11479);
and U16029 (N_16029,N_10704,N_11161);
nor U16030 (N_16030,N_9824,N_10737);
xor U16031 (N_16031,N_11555,N_8048);
nor U16032 (N_16032,N_6917,N_6506);
xor U16033 (N_16033,N_9327,N_7151);
and U16034 (N_16034,N_9773,N_9895);
xor U16035 (N_16035,N_9499,N_11244);
or U16036 (N_16036,N_11513,N_8296);
and U16037 (N_16037,N_6330,N_11509);
nand U16038 (N_16038,N_11541,N_6139);
nor U16039 (N_16039,N_6790,N_6560);
nor U16040 (N_16040,N_10860,N_8052);
nor U16041 (N_16041,N_6456,N_6416);
nand U16042 (N_16042,N_11222,N_7379);
nor U16043 (N_16043,N_9092,N_7455);
or U16044 (N_16044,N_11785,N_10810);
and U16045 (N_16045,N_8536,N_11326);
and U16046 (N_16046,N_11284,N_9837);
nand U16047 (N_16047,N_6306,N_7459);
and U16048 (N_16048,N_6842,N_8200);
and U16049 (N_16049,N_10698,N_6709);
nand U16050 (N_16050,N_11501,N_8728);
or U16051 (N_16051,N_10234,N_9641);
or U16052 (N_16052,N_6847,N_10071);
nand U16053 (N_16053,N_10316,N_11862);
nand U16054 (N_16054,N_10961,N_10751);
xnor U16055 (N_16055,N_10290,N_8451);
and U16056 (N_16056,N_11899,N_6664);
xnor U16057 (N_16057,N_6784,N_8131);
nand U16058 (N_16058,N_9851,N_7562);
xor U16059 (N_16059,N_9222,N_11345);
nor U16060 (N_16060,N_10596,N_8602);
nor U16061 (N_16061,N_10466,N_9713);
nand U16062 (N_16062,N_11118,N_7857);
nor U16063 (N_16063,N_9435,N_6313);
and U16064 (N_16064,N_6759,N_9525);
nand U16065 (N_16065,N_11721,N_10748);
nor U16066 (N_16066,N_7822,N_11356);
nor U16067 (N_16067,N_7373,N_9842);
and U16068 (N_16068,N_9994,N_11531);
and U16069 (N_16069,N_10278,N_8767);
or U16070 (N_16070,N_8406,N_9889);
nand U16071 (N_16071,N_7922,N_10167);
nand U16072 (N_16072,N_11267,N_8944);
or U16073 (N_16073,N_7185,N_11492);
or U16074 (N_16074,N_9259,N_9442);
or U16075 (N_16075,N_7114,N_7101);
xor U16076 (N_16076,N_6795,N_10149);
or U16077 (N_16077,N_10271,N_11167);
xor U16078 (N_16078,N_10973,N_10327);
or U16079 (N_16079,N_10726,N_8557);
nand U16080 (N_16080,N_11442,N_7817);
or U16081 (N_16081,N_7079,N_6769);
or U16082 (N_16082,N_6335,N_10688);
nand U16083 (N_16083,N_11449,N_10624);
nor U16084 (N_16084,N_11246,N_11804);
xor U16085 (N_16085,N_10335,N_11729);
nand U16086 (N_16086,N_11388,N_10191);
nand U16087 (N_16087,N_8285,N_8594);
nor U16088 (N_16088,N_11219,N_7518);
nor U16089 (N_16089,N_6984,N_8888);
or U16090 (N_16090,N_8122,N_7210);
nand U16091 (N_16091,N_7553,N_9095);
nor U16092 (N_16092,N_7107,N_10344);
nand U16093 (N_16093,N_10861,N_10028);
or U16094 (N_16094,N_8217,N_8645);
and U16095 (N_16095,N_6909,N_8493);
and U16096 (N_16096,N_10480,N_10703);
xor U16097 (N_16097,N_7530,N_8975);
nor U16098 (N_16098,N_10320,N_11167);
nor U16099 (N_16099,N_7443,N_6543);
nand U16100 (N_16100,N_8691,N_11682);
nand U16101 (N_16101,N_10912,N_7133);
xor U16102 (N_16102,N_10838,N_6352);
or U16103 (N_16103,N_9903,N_10247);
xnor U16104 (N_16104,N_7088,N_11513);
xor U16105 (N_16105,N_7804,N_9080);
and U16106 (N_16106,N_11258,N_8448);
and U16107 (N_16107,N_10474,N_7403);
nand U16108 (N_16108,N_11836,N_6403);
or U16109 (N_16109,N_7302,N_8971);
xor U16110 (N_16110,N_6648,N_6015);
and U16111 (N_16111,N_8115,N_10391);
nor U16112 (N_16112,N_8761,N_6535);
or U16113 (N_16113,N_8751,N_10883);
nand U16114 (N_16114,N_6414,N_11994);
nand U16115 (N_16115,N_10157,N_8927);
and U16116 (N_16116,N_6992,N_8004);
xnor U16117 (N_16117,N_6091,N_6703);
or U16118 (N_16118,N_8874,N_11446);
or U16119 (N_16119,N_9058,N_10378);
or U16120 (N_16120,N_8950,N_10285);
xor U16121 (N_16121,N_6475,N_10104);
nand U16122 (N_16122,N_7528,N_11837);
nand U16123 (N_16123,N_7669,N_10505);
xnor U16124 (N_16124,N_8949,N_6747);
and U16125 (N_16125,N_10097,N_10003);
nor U16126 (N_16126,N_10562,N_10074);
and U16127 (N_16127,N_10679,N_8227);
xor U16128 (N_16128,N_11240,N_6186);
or U16129 (N_16129,N_7383,N_11514);
nand U16130 (N_16130,N_6584,N_8061);
xnor U16131 (N_16131,N_7058,N_10141);
nor U16132 (N_16132,N_10822,N_10190);
xnor U16133 (N_16133,N_11857,N_7951);
nor U16134 (N_16134,N_6794,N_6955);
and U16135 (N_16135,N_11989,N_9173);
nor U16136 (N_16136,N_9356,N_8420);
nand U16137 (N_16137,N_8766,N_11670);
nand U16138 (N_16138,N_11217,N_10873);
or U16139 (N_16139,N_6260,N_9368);
and U16140 (N_16140,N_10080,N_8751);
xnor U16141 (N_16141,N_7483,N_8658);
or U16142 (N_16142,N_8542,N_10568);
xnor U16143 (N_16143,N_7049,N_6213);
and U16144 (N_16144,N_8213,N_10678);
nand U16145 (N_16145,N_7711,N_7380);
or U16146 (N_16146,N_9002,N_6150);
nor U16147 (N_16147,N_7028,N_10778);
nand U16148 (N_16148,N_6912,N_9944);
nand U16149 (N_16149,N_6342,N_7277);
and U16150 (N_16150,N_8855,N_9033);
nand U16151 (N_16151,N_8085,N_10229);
nand U16152 (N_16152,N_7100,N_11182);
and U16153 (N_16153,N_7702,N_6185);
nand U16154 (N_16154,N_9356,N_7535);
or U16155 (N_16155,N_8425,N_6035);
and U16156 (N_16156,N_8080,N_9247);
nand U16157 (N_16157,N_10180,N_10279);
nand U16158 (N_16158,N_10435,N_11973);
and U16159 (N_16159,N_6662,N_6190);
and U16160 (N_16160,N_8240,N_7478);
nand U16161 (N_16161,N_8963,N_10769);
or U16162 (N_16162,N_7838,N_6069);
or U16163 (N_16163,N_11491,N_6553);
xor U16164 (N_16164,N_11885,N_8059);
and U16165 (N_16165,N_6076,N_9511);
or U16166 (N_16166,N_11070,N_8157);
xnor U16167 (N_16167,N_6679,N_7980);
nand U16168 (N_16168,N_8638,N_6024);
or U16169 (N_16169,N_8130,N_8508);
nand U16170 (N_16170,N_11526,N_9634);
and U16171 (N_16171,N_10288,N_9832);
nand U16172 (N_16172,N_6375,N_9837);
and U16173 (N_16173,N_7798,N_8407);
or U16174 (N_16174,N_11112,N_9556);
nand U16175 (N_16175,N_10315,N_9598);
nor U16176 (N_16176,N_6004,N_11424);
or U16177 (N_16177,N_8791,N_8420);
xor U16178 (N_16178,N_11941,N_6749);
or U16179 (N_16179,N_8132,N_7367);
and U16180 (N_16180,N_7834,N_6843);
nor U16181 (N_16181,N_9935,N_10981);
or U16182 (N_16182,N_6506,N_10364);
and U16183 (N_16183,N_9958,N_10789);
xnor U16184 (N_16184,N_7463,N_7289);
xor U16185 (N_16185,N_9727,N_11311);
xor U16186 (N_16186,N_9354,N_11565);
nand U16187 (N_16187,N_7875,N_9600);
and U16188 (N_16188,N_6216,N_11061);
nor U16189 (N_16189,N_8513,N_6090);
xnor U16190 (N_16190,N_7529,N_10163);
xor U16191 (N_16191,N_8807,N_8170);
nor U16192 (N_16192,N_7855,N_8539);
xor U16193 (N_16193,N_8242,N_9408);
or U16194 (N_16194,N_8559,N_10165);
or U16195 (N_16195,N_7357,N_8336);
nor U16196 (N_16196,N_7195,N_9001);
xor U16197 (N_16197,N_9671,N_8694);
or U16198 (N_16198,N_10542,N_6898);
xor U16199 (N_16199,N_6454,N_10715);
or U16200 (N_16200,N_9925,N_9289);
nand U16201 (N_16201,N_11171,N_7355);
or U16202 (N_16202,N_6010,N_7377);
or U16203 (N_16203,N_7846,N_7353);
nand U16204 (N_16204,N_8657,N_8590);
xnor U16205 (N_16205,N_8770,N_7001);
and U16206 (N_16206,N_7404,N_8788);
xnor U16207 (N_16207,N_8986,N_6181);
xor U16208 (N_16208,N_7285,N_9610);
nand U16209 (N_16209,N_10665,N_7112);
nand U16210 (N_16210,N_8829,N_10607);
nand U16211 (N_16211,N_11282,N_8208);
or U16212 (N_16212,N_8198,N_11443);
or U16213 (N_16213,N_8481,N_6319);
and U16214 (N_16214,N_6683,N_8173);
and U16215 (N_16215,N_6788,N_7548);
or U16216 (N_16216,N_7178,N_11028);
nand U16217 (N_16217,N_8308,N_6689);
xor U16218 (N_16218,N_10488,N_7038);
or U16219 (N_16219,N_8346,N_6491);
or U16220 (N_16220,N_8464,N_7745);
xnor U16221 (N_16221,N_6128,N_7052);
or U16222 (N_16222,N_10231,N_7964);
or U16223 (N_16223,N_11591,N_6978);
xor U16224 (N_16224,N_11858,N_8551);
or U16225 (N_16225,N_8807,N_6399);
or U16226 (N_16226,N_7564,N_9871);
nand U16227 (N_16227,N_10140,N_7540);
nor U16228 (N_16228,N_10791,N_10793);
xnor U16229 (N_16229,N_11953,N_7789);
nor U16230 (N_16230,N_7534,N_10051);
xor U16231 (N_16231,N_9994,N_10094);
xor U16232 (N_16232,N_6537,N_7138);
xor U16233 (N_16233,N_10661,N_8117);
xor U16234 (N_16234,N_7870,N_9721);
xnor U16235 (N_16235,N_9574,N_10456);
xnor U16236 (N_16236,N_6706,N_8156);
and U16237 (N_16237,N_8744,N_11524);
or U16238 (N_16238,N_10957,N_7239);
xnor U16239 (N_16239,N_10092,N_7039);
nor U16240 (N_16240,N_6439,N_7831);
and U16241 (N_16241,N_9135,N_6897);
nand U16242 (N_16242,N_8821,N_7666);
and U16243 (N_16243,N_7589,N_6393);
or U16244 (N_16244,N_9640,N_7655);
xnor U16245 (N_16245,N_10390,N_9081);
xnor U16246 (N_16246,N_10428,N_8980);
xor U16247 (N_16247,N_6439,N_11754);
nor U16248 (N_16248,N_10820,N_10750);
nand U16249 (N_16249,N_10034,N_11938);
nor U16250 (N_16250,N_10131,N_7433);
or U16251 (N_16251,N_9652,N_6500);
nor U16252 (N_16252,N_9000,N_9588);
xnor U16253 (N_16253,N_9592,N_7562);
nand U16254 (N_16254,N_6517,N_10123);
nor U16255 (N_16255,N_9151,N_11445);
nor U16256 (N_16256,N_7584,N_10911);
or U16257 (N_16257,N_6920,N_7703);
xor U16258 (N_16258,N_10663,N_10674);
nand U16259 (N_16259,N_10509,N_8644);
nor U16260 (N_16260,N_7407,N_11966);
or U16261 (N_16261,N_8405,N_7793);
nand U16262 (N_16262,N_9189,N_6034);
or U16263 (N_16263,N_7494,N_6644);
xor U16264 (N_16264,N_6457,N_10504);
nor U16265 (N_16265,N_8948,N_7959);
xnor U16266 (N_16266,N_9845,N_11605);
xor U16267 (N_16267,N_10529,N_10378);
and U16268 (N_16268,N_10890,N_8591);
and U16269 (N_16269,N_9786,N_11788);
xor U16270 (N_16270,N_8692,N_9453);
or U16271 (N_16271,N_11341,N_7593);
nand U16272 (N_16272,N_9456,N_11573);
nor U16273 (N_16273,N_9709,N_7924);
xnor U16274 (N_16274,N_6694,N_6458);
nand U16275 (N_16275,N_7140,N_8564);
and U16276 (N_16276,N_11388,N_8105);
or U16277 (N_16277,N_10000,N_6489);
and U16278 (N_16278,N_9991,N_7758);
xnor U16279 (N_16279,N_11452,N_6238);
and U16280 (N_16280,N_9019,N_11499);
nand U16281 (N_16281,N_6106,N_8464);
xnor U16282 (N_16282,N_9920,N_7646);
xor U16283 (N_16283,N_9212,N_7389);
nor U16284 (N_16284,N_7205,N_7889);
or U16285 (N_16285,N_7402,N_11026);
and U16286 (N_16286,N_10975,N_8743);
xor U16287 (N_16287,N_7927,N_11692);
xnor U16288 (N_16288,N_9226,N_9049);
and U16289 (N_16289,N_10946,N_6290);
nor U16290 (N_16290,N_9969,N_7224);
nor U16291 (N_16291,N_11047,N_11738);
nor U16292 (N_16292,N_8064,N_7975);
xor U16293 (N_16293,N_7989,N_11383);
xnor U16294 (N_16294,N_9777,N_10875);
or U16295 (N_16295,N_6019,N_6442);
nand U16296 (N_16296,N_8832,N_11762);
nor U16297 (N_16297,N_7553,N_7155);
nor U16298 (N_16298,N_6515,N_8054);
xnor U16299 (N_16299,N_8524,N_7320);
nor U16300 (N_16300,N_7978,N_11208);
xor U16301 (N_16301,N_11110,N_10351);
nor U16302 (N_16302,N_8544,N_7214);
nor U16303 (N_16303,N_7279,N_7885);
or U16304 (N_16304,N_7104,N_9196);
nor U16305 (N_16305,N_10655,N_9194);
xor U16306 (N_16306,N_7343,N_11176);
xnor U16307 (N_16307,N_11955,N_7836);
nor U16308 (N_16308,N_9288,N_9409);
nor U16309 (N_16309,N_10604,N_6124);
or U16310 (N_16310,N_11837,N_8242);
xnor U16311 (N_16311,N_7884,N_7062);
and U16312 (N_16312,N_9177,N_7173);
xnor U16313 (N_16313,N_10079,N_9220);
xor U16314 (N_16314,N_9234,N_6105);
and U16315 (N_16315,N_7801,N_11169);
and U16316 (N_16316,N_8266,N_10116);
or U16317 (N_16317,N_10486,N_8172);
xnor U16318 (N_16318,N_10368,N_8661);
and U16319 (N_16319,N_9809,N_6528);
or U16320 (N_16320,N_7739,N_10270);
nor U16321 (N_16321,N_10804,N_9008);
nor U16322 (N_16322,N_10284,N_11047);
nand U16323 (N_16323,N_11951,N_10783);
or U16324 (N_16324,N_6760,N_6155);
xor U16325 (N_16325,N_10350,N_10093);
xor U16326 (N_16326,N_6279,N_6196);
xor U16327 (N_16327,N_8423,N_7743);
xnor U16328 (N_16328,N_11504,N_7335);
nor U16329 (N_16329,N_10728,N_8666);
nand U16330 (N_16330,N_11520,N_8753);
or U16331 (N_16331,N_7653,N_9221);
and U16332 (N_16332,N_11070,N_11250);
and U16333 (N_16333,N_11451,N_11205);
and U16334 (N_16334,N_8495,N_8012);
nor U16335 (N_16335,N_10988,N_6447);
nor U16336 (N_16336,N_7063,N_7080);
and U16337 (N_16337,N_9304,N_10381);
xnor U16338 (N_16338,N_8306,N_8493);
and U16339 (N_16339,N_7605,N_11630);
nor U16340 (N_16340,N_8899,N_8664);
nand U16341 (N_16341,N_7427,N_10236);
nand U16342 (N_16342,N_11139,N_8946);
or U16343 (N_16343,N_6324,N_8248);
or U16344 (N_16344,N_8226,N_9325);
nor U16345 (N_16345,N_10290,N_7488);
and U16346 (N_16346,N_7504,N_6801);
xor U16347 (N_16347,N_9903,N_7698);
xor U16348 (N_16348,N_6798,N_6130);
nand U16349 (N_16349,N_9771,N_9416);
and U16350 (N_16350,N_6451,N_10698);
nor U16351 (N_16351,N_11152,N_10783);
and U16352 (N_16352,N_8654,N_10627);
nor U16353 (N_16353,N_11539,N_11774);
nand U16354 (N_16354,N_11760,N_11151);
xnor U16355 (N_16355,N_11883,N_11798);
nor U16356 (N_16356,N_6999,N_10855);
and U16357 (N_16357,N_7113,N_7539);
or U16358 (N_16358,N_9563,N_8013);
or U16359 (N_16359,N_7818,N_6905);
nand U16360 (N_16360,N_6674,N_6234);
xnor U16361 (N_16361,N_7225,N_7571);
nor U16362 (N_16362,N_8796,N_7533);
xor U16363 (N_16363,N_10060,N_6854);
nor U16364 (N_16364,N_11021,N_9532);
and U16365 (N_16365,N_11873,N_7305);
nor U16366 (N_16366,N_8081,N_8568);
or U16367 (N_16367,N_11717,N_7878);
and U16368 (N_16368,N_7528,N_11411);
xor U16369 (N_16369,N_9289,N_11149);
nand U16370 (N_16370,N_6894,N_6716);
nand U16371 (N_16371,N_6072,N_8755);
nor U16372 (N_16372,N_10708,N_6403);
and U16373 (N_16373,N_6055,N_9552);
nor U16374 (N_16374,N_10795,N_6308);
xnor U16375 (N_16375,N_10799,N_7075);
and U16376 (N_16376,N_9261,N_8400);
or U16377 (N_16377,N_10750,N_11710);
xnor U16378 (N_16378,N_7101,N_8179);
xnor U16379 (N_16379,N_9301,N_6942);
or U16380 (N_16380,N_11651,N_6851);
or U16381 (N_16381,N_11974,N_10583);
or U16382 (N_16382,N_6952,N_10284);
nor U16383 (N_16383,N_8194,N_11121);
nor U16384 (N_16384,N_6886,N_9915);
xor U16385 (N_16385,N_7986,N_6698);
nand U16386 (N_16386,N_6137,N_11182);
nor U16387 (N_16387,N_11810,N_8131);
and U16388 (N_16388,N_8959,N_9439);
xor U16389 (N_16389,N_10345,N_7210);
nor U16390 (N_16390,N_7671,N_9614);
xnor U16391 (N_16391,N_9997,N_8400);
xnor U16392 (N_16392,N_10651,N_9970);
nand U16393 (N_16393,N_6321,N_11960);
xnor U16394 (N_16394,N_10031,N_7337);
nor U16395 (N_16395,N_7564,N_9129);
xor U16396 (N_16396,N_11369,N_10702);
xor U16397 (N_16397,N_10325,N_11263);
xnor U16398 (N_16398,N_10034,N_6848);
nand U16399 (N_16399,N_10549,N_10864);
nor U16400 (N_16400,N_11727,N_10215);
and U16401 (N_16401,N_6289,N_9467);
nand U16402 (N_16402,N_6892,N_7656);
nor U16403 (N_16403,N_7084,N_8723);
nor U16404 (N_16404,N_11473,N_8124);
xnor U16405 (N_16405,N_6381,N_7632);
and U16406 (N_16406,N_8667,N_9379);
or U16407 (N_16407,N_11453,N_6863);
nand U16408 (N_16408,N_9301,N_8703);
nand U16409 (N_16409,N_7716,N_7308);
xor U16410 (N_16410,N_6642,N_8998);
nor U16411 (N_16411,N_10482,N_7124);
nand U16412 (N_16412,N_7557,N_6124);
or U16413 (N_16413,N_7536,N_7434);
and U16414 (N_16414,N_11324,N_10059);
or U16415 (N_16415,N_7498,N_11415);
nor U16416 (N_16416,N_11470,N_6639);
nor U16417 (N_16417,N_9633,N_6934);
nand U16418 (N_16418,N_10623,N_9992);
or U16419 (N_16419,N_10227,N_11985);
nand U16420 (N_16420,N_7996,N_6944);
or U16421 (N_16421,N_8449,N_10014);
nand U16422 (N_16422,N_11095,N_6773);
or U16423 (N_16423,N_10553,N_11577);
or U16424 (N_16424,N_9553,N_8578);
nand U16425 (N_16425,N_6853,N_7193);
xor U16426 (N_16426,N_8183,N_8534);
nor U16427 (N_16427,N_7475,N_10939);
nand U16428 (N_16428,N_11786,N_8455);
nand U16429 (N_16429,N_11702,N_10805);
nand U16430 (N_16430,N_6336,N_8488);
xnor U16431 (N_16431,N_7427,N_11986);
xor U16432 (N_16432,N_10546,N_11457);
nand U16433 (N_16433,N_10802,N_6972);
nand U16434 (N_16434,N_6771,N_9348);
nand U16435 (N_16435,N_6993,N_9349);
or U16436 (N_16436,N_10805,N_10927);
nand U16437 (N_16437,N_7116,N_10193);
xor U16438 (N_16438,N_6098,N_8014);
nand U16439 (N_16439,N_9928,N_8052);
nand U16440 (N_16440,N_11608,N_7525);
nor U16441 (N_16441,N_7946,N_8772);
xor U16442 (N_16442,N_11098,N_7679);
nand U16443 (N_16443,N_7976,N_6648);
and U16444 (N_16444,N_11802,N_6036);
xnor U16445 (N_16445,N_10864,N_8363);
and U16446 (N_16446,N_10133,N_9293);
xnor U16447 (N_16447,N_6835,N_10042);
nand U16448 (N_16448,N_10488,N_6711);
or U16449 (N_16449,N_7774,N_7876);
nand U16450 (N_16450,N_9082,N_6711);
and U16451 (N_16451,N_7461,N_6060);
xnor U16452 (N_16452,N_7212,N_10830);
nand U16453 (N_16453,N_9484,N_7427);
xor U16454 (N_16454,N_9134,N_7385);
nor U16455 (N_16455,N_6821,N_9255);
nor U16456 (N_16456,N_10240,N_11678);
and U16457 (N_16457,N_9710,N_10664);
or U16458 (N_16458,N_9656,N_7445);
nor U16459 (N_16459,N_7601,N_7337);
nand U16460 (N_16460,N_8344,N_11565);
or U16461 (N_16461,N_11050,N_9805);
nor U16462 (N_16462,N_9895,N_8048);
xor U16463 (N_16463,N_10398,N_9526);
or U16464 (N_16464,N_7612,N_6678);
nor U16465 (N_16465,N_11450,N_7007);
nand U16466 (N_16466,N_8259,N_10066);
nor U16467 (N_16467,N_7589,N_10334);
or U16468 (N_16468,N_9295,N_11625);
and U16469 (N_16469,N_9110,N_11391);
xor U16470 (N_16470,N_10887,N_7814);
or U16471 (N_16471,N_8622,N_6921);
nand U16472 (N_16472,N_6947,N_10817);
and U16473 (N_16473,N_9049,N_10834);
nor U16474 (N_16474,N_9822,N_9328);
nor U16475 (N_16475,N_8858,N_8884);
nand U16476 (N_16476,N_10384,N_7342);
xnor U16477 (N_16477,N_7820,N_8595);
xnor U16478 (N_16478,N_10211,N_9985);
nand U16479 (N_16479,N_6528,N_11843);
and U16480 (N_16480,N_6484,N_8564);
or U16481 (N_16481,N_9494,N_6704);
nand U16482 (N_16482,N_9055,N_6083);
nor U16483 (N_16483,N_7265,N_10161);
and U16484 (N_16484,N_8443,N_8044);
nand U16485 (N_16485,N_9050,N_10904);
nor U16486 (N_16486,N_10328,N_9085);
nor U16487 (N_16487,N_9191,N_11321);
and U16488 (N_16488,N_6665,N_10874);
or U16489 (N_16489,N_11969,N_9510);
or U16490 (N_16490,N_10949,N_7356);
xor U16491 (N_16491,N_6302,N_11228);
xor U16492 (N_16492,N_9340,N_8477);
nor U16493 (N_16493,N_10682,N_10825);
nand U16494 (N_16494,N_8737,N_10169);
nand U16495 (N_16495,N_11267,N_9696);
xnor U16496 (N_16496,N_7851,N_6602);
nor U16497 (N_16497,N_7201,N_8184);
and U16498 (N_16498,N_8303,N_6972);
xor U16499 (N_16499,N_11694,N_6143);
xor U16500 (N_16500,N_9411,N_7799);
xor U16501 (N_16501,N_6049,N_9972);
nand U16502 (N_16502,N_11249,N_10700);
xor U16503 (N_16503,N_7721,N_11218);
xor U16504 (N_16504,N_6572,N_11419);
or U16505 (N_16505,N_11426,N_6540);
xnor U16506 (N_16506,N_10600,N_7517);
nand U16507 (N_16507,N_7329,N_11093);
and U16508 (N_16508,N_6066,N_10173);
or U16509 (N_16509,N_7880,N_8496);
nand U16510 (N_16510,N_11550,N_9672);
nor U16511 (N_16511,N_8236,N_10658);
nand U16512 (N_16512,N_10720,N_11144);
xnor U16513 (N_16513,N_6113,N_10726);
xor U16514 (N_16514,N_7475,N_9564);
and U16515 (N_16515,N_11141,N_8607);
and U16516 (N_16516,N_9441,N_7943);
xor U16517 (N_16517,N_7741,N_10815);
or U16518 (N_16518,N_8084,N_7457);
xor U16519 (N_16519,N_8485,N_8462);
and U16520 (N_16520,N_11399,N_9072);
or U16521 (N_16521,N_6286,N_10051);
nor U16522 (N_16522,N_6282,N_11324);
nor U16523 (N_16523,N_9624,N_6825);
and U16524 (N_16524,N_9570,N_11220);
and U16525 (N_16525,N_8891,N_11945);
and U16526 (N_16526,N_11188,N_11890);
or U16527 (N_16527,N_9590,N_8189);
nand U16528 (N_16528,N_6120,N_8844);
or U16529 (N_16529,N_6067,N_7817);
xor U16530 (N_16530,N_6155,N_11725);
nand U16531 (N_16531,N_10589,N_6021);
nand U16532 (N_16532,N_6224,N_10589);
nand U16533 (N_16533,N_10098,N_11756);
nor U16534 (N_16534,N_7482,N_9376);
xor U16535 (N_16535,N_11076,N_8771);
and U16536 (N_16536,N_9699,N_6568);
xnor U16537 (N_16537,N_9785,N_8866);
xor U16538 (N_16538,N_7004,N_8413);
nor U16539 (N_16539,N_7349,N_7854);
nor U16540 (N_16540,N_6759,N_10188);
and U16541 (N_16541,N_6230,N_7650);
and U16542 (N_16542,N_10328,N_10831);
nor U16543 (N_16543,N_7309,N_8344);
nand U16544 (N_16544,N_9623,N_6769);
xnor U16545 (N_16545,N_6052,N_10003);
nand U16546 (N_16546,N_9051,N_9852);
nand U16547 (N_16547,N_8862,N_7874);
and U16548 (N_16548,N_6763,N_10922);
and U16549 (N_16549,N_6969,N_10687);
and U16550 (N_16550,N_11245,N_8595);
or U16551 (N_16551,N_9394,N_11874);
or U16552 (N_16552,N_8592,N_7312);
xnor U16553 (N_16553,N_10655,N_8765);
or U16554 (N_16554,N_7732,N_11448);
or U16555 (N_16555,N_8870,N_8351);
and U16556 (N_16556,N_7557,N_7792);
nor U16557 (N_16557,N_10645,N_9398);
xnor U16558 (N_16558,N_7833,N_10520);
xor U16559 (N_16559,N_10496,N_8909);
nor U16560 (N_16560,N_7142,N_10159);
nand U16561 (N_16561,N_11819,N_8155);
or U16562 (N_16562,N_6326,N_6047);
or U16563 (N_16563,N_7834,N_8312);
or U16564 (N_16564,N_7757,N_7972);
or U16565 (N_16565,N_10022,N_7480);
nor U16566 (N_16566,N_10273,N_6395);
xnor U16567 (N_16567,N_7631,N_9871);
nor U16568 (N_16568,N_8640,N_6918);
and U16569 (N_16569,N_6907,N_10393);
nor U16570 (N_16570,N_9073,N_9537);
nor U16571 (N_16571,N_8869,N_8510);
nand U16572 (N_16572,N_8214,N_6027);
xor U16573 (N_16573,N_11853,N_10215);
and U16574 (N_16574,N_6332,N_10293);
or U16575 (N_16575,N_10052,N_11425);
nand U16576 (N_16576,N_9734,N_9996);
nand U16577 (N_16577,N_9715,N_6984);
and U16578 (N_16578,N_8773,N_7576);
xnor U16579 (N_16579,N_8491,N_9739);
nor U16580 (N_16580,N_11368,N_7841);
and U16581 (N_16581,N_9591,N_6855);
nand U16582 (N_16582,N_9838,N_7818);
or U16583 (N_16583,N_10967,N_9702);
nand U16584 (N_16584,N_9115,N_7246);
or U16585 (N_16585,N_7182,N_10034);
nand U16586 (N_16586,N_9662,N_11718);
and U16587 (N_16587,N_9838,N_9248);
xor U16588 (N_16588,N_11174,N_6604);
xnor U16589 (N_16589,N_8542,N_6997);
and U16590 (N_16590,N_10720,N_7146);
nor U16591 (N_16591,N_8673,N_8266);
nor U16592 (N_16592,N_11593,N_8609);
and U16593 (N_16593,N_9954,N_10997);
nor U16594 (N_16594,N_11003,N_11361);
nand U16595 (N_16595,N_6033,N_11726);
xnor U16596 (N_16596,N_10924,N_11583);
and U16597 (N_16597,N_8878,N_8910);
nor U16598 (N_16598,N_6218,N_7500);
or U16599 (N_16599,N_6794,N_9046);
nor U16600 (N_16600,N_11254,N_6125);
nor U16601 (N_16601,N_9731,N_6450);
and U16602 (N_16602,N_9441,N_11858);
or U16603 (N_16603,N_7205,N_7774);
nand U16604 (N_16604,N_10075,N_6303);
or U16605 (N_16605,N_7903,N_9981);
nand U16606 (N_16606,N_7227,N_11978);
xnor U16607 (N_16607,N_7580,N_11638);
nor U16608 (N_16608,N_9764,N_11427);
nand U16609 (N_16609,N_10107,N_11501);
and U16610 (N_16610,N_10463,N_8830);
and U16611 (N_16611,N_7233,N_6251);
and U16612 (N_16612,N_11917,N_6869);
or U16613 (N_16613,N_11280,N_11458);
and U16614 (N_16614,N_8804,N_11695);
or U16615 (N_16615,N_10723,N_11127);
xnor U16616 (N_16616,N_7152,N_7069);
and U16617 (N_16617,N_11894,N_11234);
nor U16618 (N_16618,N_9645,N_8021);
or U16619 (N_16619,N_9067,N_6161);
nand U16620 (N_16620,N_10471,N_11384);
and U16621 (N_16621,N_11329,N_11261);
or U16622 (N_16622,N_9937,N_7938);
or U16623 (N_16623,N_9298,N_9954);
xor U16624 (N_16624,N_9622,N_6740);
or U16625 (N_16625,N_10118,N_9124);
or U16626 (N_16626,N_11185,N_10622);
or U16627 (N_16627,N_11540,N_11929);
and U16628 (N_16628,N_8953,N_10108);
and U16629 (N_16629,N_11347,N_9528);
nand U16630 (N_16630,N_11390,N_7914);
or U16631 (N_16631,N_10715,N_8737);
xor U16632 (N_16632,N_10936,N_9345);
nand U16633 (N_16633,N_9969,N_7173);
xor U16634 (N_16634,N_7428,N_7814);
and U16635 (N_16635,N_6727,N_9027);
nand U16636 (N_16636,N_7952,N_6748);
and U16637 (N_16637,N_6248,N_7335);
nand U16638 (N_16638,N_7117,N_8119);
xnor U16639 (N_16639,N_11147,N_9955);
nor U16640 (N_16640,N_10245,N_6260);
xnor U16641 (N_16641,N_8664,N_7136);
xnor U16642 (N_16642,N_8355,N_8242);
and U16643 (N_16643,N_7050,N_9336);
nand U16644 (N_16644,N_11273,N_6847);
nor U16645 (N_16645,N_10005,N_6370);
xor U16646 (N_16646,N_8656,N_11265);
and U16647 (N_16647,N_8292,N_11147);
nor U16648 (N_16648,N_9874,N_9626);
and U16649 (N_16649,N_7985,N_9808);
xnor U16650 (N_16650,N_11849,N_10934);
or U16651 (N_16651,N_11012,N_7055);
nor U16652 (N_16652,N_6815,N_10485);
and U16653 (N_16653,N_11318,N_6085);
nor U16654 (N_16654,N_11341,N_10573);
nor U16655 (N_16655,N_6010,N_8983);
and U16656 (N_16656,N_6922,N_10199);
and U16657 (N_16657,N_11572,N_9925);
nand U16658 (N_16658,N_7501,N_7902);
nand U16659 (N_16659,N_11059,N_9025);
or U16660 (N_16660,N_6247,N_9726);
and U16661 (N_16661,N_8990,N_7397);
nor U16662 (N_16662,N_7954,N_8391);
nand U16663 (N_16663,N_9302,N_11728);
nand U16664 (N_16664,N_6012,N_7644);
or U16665 (N_16665,N_6097,N_11983);
nand U16666 (N_16666,N_10548,N_7737);
or U16667 (N_16667,N_6340,N_10514);
nor U16668 (N_16668,N_6809,N_11248);
xnor U16669 (N_16669,N_6752,N_9960);
xor U16670 (N_16670,N_6416,N_7351);
nor U16671 (N_16671,N_10284,N_10146);
or U16672 (N_16672,N_10379,N_9979);
or U16673 (N_16673,N_6400,N_8406);
nand U16674 (N_16674,N_8921,N_9068);
nand U16675 (N_16675,N_6037,N_10979);
or U16676 (N_16676,N_10071,N_7856);
or U16677 (N_16677,N_9938,N_6713);
nor U16678 (N_16678,N_9385,N_10844);
or U16679 (N_16679,N_11112,N_11138);
xnor U16680 (N_16680,N_9281,N_6698);
or U16681 (N_16681,N_6327,N_10796);
and U16682 (N_16682,N_10577,N_8605);
nand U16683 (N_16683,N_6949,N_10446);
and U16684 (N_16684,N_10846,N_7837);
xnor U16685 (N_16685,N_8297,N_11336);
nor U16686 (N_16686,N_11914,N_11697);
nor U16687 (N_16687,N_6110,N_9023);
nor U16688 (N_16688,N_7192,N_9361);
or U16689 (N_16689,N_6623,N_6240);
and U16690 (N_16690,N_10264,N_7191);
or U16691 (N_16691,N_11875,N_8001);
and U16692 (N_16692,N_9074,N_7499);
and U16693 (N_16693,N_7987,N_7107);
and U16694 (N_16694,N_7212,N_10634);
and U16695 (N_16695,N_6166,N_8595);
and U16696 (N_16696,N_8859,N_7718);
or U16697 (N_16697,N_10068,N_9053);
nor U16698 (N_16698,N_10282,N_8351);
nor U16699 (N_16699,N_10168,N_7201);
and U16700 (N_16700,N_6856,N_11100);
xor U16701 (N_16701,N_6154,N_9508);
or U16702 (N_16702,N_11378,N_10000);
or U16703 (N_16703,N_10902,N_11144);
nand U16704 (N_16704,N_9612,N_9443);
or U16705 (N_16705,N_8045,N_11784);
or U16706 (N_16706,N_9303,N_10378);
or U16707 (N_16707,N_7180,N_10103);
and U16708 (N_16708,N_8965,N_6135);
nor U16709 (N_16709,N_6183,N_9370);
and U16710 (N_16710,N_9861,N_10431);
nor U16711 (N_16711,N_7848,N_11098);
nor U16712 (N_16712,N_8930,N_10393);
nor U16713 (N_16713,N_11782,N_6200);
and U16714 (N_16714,N_9255,N_6583);
xnor U16715 (N_16715,N_6431,N_7859);
xnor U16716 (N_16716,N_9222,N_6600);
and U16717 (N_16717,N_8158,N_8188);
and U16718 (N_16718,N_7318,N_10042);
nand U16719 (N_16719,N_7982,N_9174);
and U16720 (N_16720,N_6439,N_7402);
and U16721 (N_16721,N_11445,N_10854);
xnor U16722 (N_16722,N_7169,N_9892);
xnor U16723 (N_16723,N_11167,N_10018);
nand U16724 (N_16724,N_9583,N_8677);
and U16725 (N_16725,N_6715,N_8396);
xnor U16726 (N_16726,N_7529,N_7852);
or U16727 (N_16727,N_6634,N_8156);
nand U16728 (N_16728,N_6432,N_6972);
xor U16729 (N_16729,N_7990,N_11736);
xor U16730 (N_16730,N_9665,N_10712);
nor U16731 (N_16731,N_11503,N_7711);
xnor U16732 (N_16732,N_10943,N_11218);
and U16733 (N_16733,N_7669,N_6133);
and U16734 (N_16734,N_8094,N_10419);
nor U16735 (N_16735,N_10014,N_8464);
and U16736 (N_16736,N_6026,N_6701);
and U16737 (N_16737,N_6497,N_10325);
or U16738 (N_16738,N_8084,N_7846);
nor U16739 (N_16739,N_7584,N_9738);
and U16740 (N_16740,N_11373,N_9977);
and U16741 (N_16741,N_8270,N_10165);
xor U16742 (N_16742,N_11131,N_11818);
and U16743 (N_16743,N_10891,N_9372);
nand U16744 (N_16744,N_9951,N_10317);
and U16745 (N_16745,N_11421,N_10910);
xor U16746 (N_16746,N_6050,N_8685);
nand U16747 (N_16747,N_7356,N_9523);
or U16748 (N_16748,N_11718,N_7204);
xnor U16749 (N_16749,N_8258,N_9490);
xor U16750 (N_16750,N_10698,N_6802);
nand U16751 (N_16751,N_10791,N_6325);
nand U16752 (N_16752,N_6607,N_11682);
or U16753 (N_16753,N_10954,N_6412);
or U16754 (N_16754,N_8315,N_6286);
and U16755 (N_16755,N_8750,N_6601);
and U16756 (N_16756,N_9519,N_7482);
and U16757 (N_16757,N_10084,N_9030);
nand U16758 (N_16758,N_8429,N_10550);
and U16759 (N_16759,N_10001,N_10949);
and U16760 (N_16760,N_11088,N_11581);
nand U16761 (N_16761,N_8713,N_6790);
nand U16762 (N_16762,N_7013,N_6425);
xnor U16763 (N_16763,N_6258,N_10250);
or U16764 (N_16764,N_10290,N_8306);
or U16765 (N_16765,N_11890,N_8973);
and U16766 (N_16766,N_8056,N_9946);
nor U16767 (N_16767,N_10768,N_9916);
nor U16768 (N_16768,N_6250,N_10917);
or U16769 (N_16769,N_6785,N_8767);
nor U16770 (N_16770,N_6687,N_7829);
xor U16771 (N_16771,N_6340,N_6493);
nand U16772 (N_16772,N_6174,N_10694);
or U16773 (N_16773,N_7576,N_8841);
or U16774 (N_16774,N_6475,N_10804);
or U16775 (N_16775,N_10897,N_6902);
or U16776 (N_16776,N_10505,N_11173);
nor U16777 (N_16777,N_8670,N_8455);
or U16778 (N_16778,N_7543,N_11314);
nand U16779 (N_16779,N_6080,N_7656);
nor U16780 (N_16780,N_11640,N_7787);
and U16781 (N_16781,N_11973,N_8164);
nand U16782 (N_16782,N_9978,N_6371);
or U16783 (N_16783,N_8679,N_11656);
nor U16784 (N_16784,N_11605,N_10252);
xnor U16785 (N_16785,N_10878,N_9211);
xnor U16786 (N_16786,N_8028,N_9667);
and U16787 (N_16787,N_9496,N_11318);
nor U16788 (N_16788,N_7811,N_10601);
nand U16789 (N_16789,N_8568,N_9403);
and U16790 (N_16790,N_6104,N_8705);
nand U16791 (N_16791,N_11458,N_6202);
or U16792 (N_16792,N_7371,N_6712);
nor U16793 (N_16793,N_11913,N_10426);
and U16794 (N_16794,N_8501,N_9066);
and U16795 (N_16795,N_11775,N_6540);
nor U16796 (N_16796,N_9555,N_9086);
and U16797 (N_16797,N_7697,N_8826);
nor U16798 (N_16798,N_10026,N_6467);
nand U16799 (N_16799,N_10533,N_9224);
nand U16800 (N_16800,N_7309,N_9780);
or U16801 (N_16801,N_8123,N_10180);
or U16802 (N_16802,N_9773,N_10975);
or U16803 (N_16803,N_11421,N_9411);
or U16804 (N_16804,N_11228,N_7836);
and U16805 (N_16805,N_6099,N_10298);
and U16806 (N_16806,N_6492,N_10236);
nor U16807 (N_16807,N_10811,N_9512);
nor U16808 (N_16808,N_9206,N_11016);
nor U16809 (N_16809,N_8063,N_11984);
or U16810 (N_16810,N_6394,N_7950);
nand U16811 (N_16811,N_11792,N_7915);
nor U16812 (N_16812,N_11789,N_9441);
xor U16813 (N_16813,N_8791,N_9894);
xnor U16814 (N_16814,N_6226,N_8558);
or U16815 (N_16815,N_9372,N_11561);
or U16816 (N_16816,N_10542,N_6816);
nor U16817 (N_16817,N_7778,N_7237);
nand U16818 (N_16818,N_11432,N_11014);
and U16819 (N_16819,N_8624,N_9111);
xor U16820 (N_16820,N_11444,N_8134);
nand U16821 (N_16821,N_9171,N_10370);
and U16822 (N_16822,N_6865,N_8304);
and U16823 (N_16823,N_8010,N_10767);
or U16824 (N_16824,N_10269,N_9828);
nand U16825 (N_16825,N_6941,N_10989);
nand U16826 (N_16826,N_10824,N_8767);
or U16827 (N_16827,N_8575,N_9367);
nor U16828 (N_16828,N_7534,N_6414);
nand U16829 (N_16829,N_11155,N_8715);
and U16830 (N_16830,N_9899,N_7288);
nand U16831 (N_16831,N_6403,N_11311);
and U16832 (N_16832,N_8943,N_9912);
nand U16833 (N_16833,N_10443,N_9397);
and U16834 (N_16834,N_6205,N_6221);
xnor U16835 (N_16835,N_7689,N_9070);
and U16836 (N_16836,N_7526,N_8915);
nand U16837 (N_16837,N_10040,N_10787);
or U16838 (N_16838,N_9853,N_8336);
and U16839 (N_16839,N_8642,N_10570);
nand U16840 (N_16840,N_7242,N_6809);
nor U16841 (N_16841,N_8049,N_7750);
and U16842 (N_16842,N_7415,N_8135);
nor U16843 (N_16843,N_9165,N_10705);
xor U16844 (N_16844,N_6455,N_8800);
and U16845 (N_16845,N_11033,N_6694);
xnor U16846 (N_16846,N_8668,N_9604);
nand U16847 (N_16847,N_11908,N_9520);
nor U16848 (N_16848,N_11934,N_11308);
and U16849 (N_16849,N_8172,N_6769);
xor U16850 (N_16850,N_9451,N_6774);
xor U16851 (N_16851,N_7660,N_11320);
or U16852 (N_16852,N_7605,N_7776);
nor U16853 (N_16853,N_11547,N_6058);
and U16854 (N_16854,N_8559,N_10751);
nand U16855 (N_16855,N_11306,N_6371);
xnor U16856 (N_16856,N_6111,N_9101);
or U16857 (N_16857,N_7198,N_11838);
or U16858 (N_16858,N_8623,N_6900);
nand U16859 (N_16859,N_10876,N_7366);
and U16860 (N_16860,N_6284,N_7655);
or U16861 (N_16861,N_7823,N_11759);
xnor U16862 (N_16862,N_10321,N_8816);
xnor U16863 (N_16863,N_8329,N_6234);
nand U16864 (N_16864,N_9038,N_9416);
nand U16865 (N_16865,N_9644,N_6017);
xnor U16866 (N_16866,N_9231,N_11221);
nand U16867 (N_16867,N_7121,N_9897);
xor U16868 (N_16868,N_11495,N_8525);
nor U16869 (N_16869,N_8561,N_6178);
xor U16870 (N_16870,N_10018,N_7012);
and U16871 (N_16871,N_8029,N_6774);
nor U16872 (N_16872,N_10997,N_9904);
or U16873 (N_16873,N_9779,N_9501);
nor U16874 (N_16874,N_10347,N_11740);
and U16875 (N_16875,N_11406,N_11190);
nand U16876 (N_16876,N_9640,N_10496);
xor U16877 (N_16877,N_6963,N_9409);
nor U16878 (N_16878,N_10844,N_9815);
nand U16879 (N_16879,N_6190,N_10061);
and U16880 (N_16880,N_8576,N_6866);
nor U16881 (N_16881,N_7415,N_11188);
xor U16882 (N_16882,N_9873,N_10189);
or U16883 (N_16883,N_6750,N_6221);
xnor U16884 (N_16884,N_8488,N_11586);
nand U16885 (N_16885,N_8550,N_10085);
nor U16886 (N_16886,N_7954,N_8803);
nor U16887 (N_16887,N_8038,N_11060);
nor U16888 (N_16888,N_11961,N_9770);
or U16889 (N_16889,N_10917,N_8290);
xor U16890 (N_16890,N_6818,N_6909);
and U16891 (N_16891,N_9662,N_10585);
nand U16892 (N_16892,N_6992,N_8287);
nand U16893 (N_16893,N_11701,N_10857);
xnor U16894 (N_16894,N_7702,N_9486);
nand U16895 (N_16895,N_8362,N_8031);
xnor U16896 (N_16896,N_9445,N_8595);
xor U16897 (N_16897,N_11840,N_7064);
and U16898 (N_16898,N_9105,N_8776);
or U16899 (N_16899,N_9517,N_9994);
and U16900 (N_16900,N_8710,N_9753);
or U16901 (N_16901,N_6904,N_8441);
and U16902 (N_16902,N_8442,N_11782);
and U16903 (N_16903,N_7309,N_10100);
and U16904 (N_16904,N_7515,N_10818);
or U16905 (N_16905,N_10127,N_7186);
and U16906 (N_16906,N_7115,N_8366);
nor U16907 (N_16907,N_9244,N_9594);
nor U16908 (N_16908,N_9003,N_8671);
nor U16909 (N_16909,N_10050,N_7545);
nor U16910 (N_16910,N_8815,N_9774);
nand U16911 (N_16911,N_6236,N_7160);
or U16912 (N_16912,N_11922,N_8907);
xnor U16913 (N_16913,N_7946,N_7522);
and U16914 (N_16914,N_11162,N_9284);
and U16915 (N_16915,N_9160,N_6205);
xnor U16916 (N_16916,N_6068,N_8895);
or U16917 (N_16917,N_11778,N_7532);
or U16918 (N_16918,N_7050,N_9375);
xor U16919 (N_16919,N_8169,N_9553);
nor U16920 (N_16920,N_8672,N_6894);
nor U16921 (N_16921,N_8931,N_10499);
nor U16922 (N_16922,N_8330,N_7565);
xnor U16923 (N_16923,N_8556,N_6374);
xor U16924 (N_16924,N_11338,N_10049);
nand U16925 (N_16925,N_10347,N_9526);
xor U16926 (N_16926,N_8875,N_7200);
xnor U16927 (N_16927,N_11989,N_9298);
or U16928 (N_16928,N_8780,N_7821);
nand U16929 (N_16929,N_10854,N_6975);
nand U16930 (N_16930,N_7194,N_10177);
and U16931 (N_16931,N_8389,N_11127);
and U16932 (N_16932,N_10978,N_8115);
xor U16933 (N_16933,N_11285,N_7123);
or U16934 (N_16934,N_8576,N_9175);
xor U16935 (N_16935,N_7135,N_8193);
and U16936 (N_16936,N_8078,N_6799);
xor U16937 (N_16937,N_8563,N_8146);
nor U16938 (N_16938,N_10116,N_11873);
and U16939 (N_16939,N_6584,N_8613);
nor U16940 (N_16940,N_7417,N_9706);
nor U16941 (N_16941,N_6735,N_8137);
and U16942 (N_16942,N_6567,N_9663);
nand U16943 (N_16943,N_7084,N_9481);
xor U16944 (N_16944,N_8988,N_6806);
nor U16945 (N_16945,N_10669,N_7822);
nand U16946 (N_16946,N_10330,N_7347);
and U16947 (N_16947,N_11668,N_10014);
and U16948 (N_16948,N_7896,N_8704);
nor U16949 (N_16949,N_10174,N_7427);
nand U16950 (N_16950,N_7636,N_6979);
or U16951 (N_16951,N_9687,N_8213);
xnor U16952 (N_16952,N_8735,N_11908);
or U16953 (N_16953,N_9893,N_8292);
nor U16954 (N_16954,N_10461,N_9791);
xor U16955 (N_16955,N_7093,N_11305);
nor U16956 (N_16956,N_8160,N_8215);
or U16957 (N_16957,N_7797,N_6654);
xor U16958 (N_16958,N_10858,N_9633);
and U16959 (N_16959,N_9078,N_9432);
nand U16960 (N_16960,N_6433,N_10539);
and U16961 (N_16961,N_10838,N_10944);
xor U16962 (N_16962,N_8060,N_11942);
and U16963 (N_16963,N_11858,N_6909);
nor U16964 (N_16964,N_6169,N_7425);
nand U16965 (N_16965,N_9829,N_10035);
xor U16966 (N_16966,N_11151,N_10643);
or U16967 (N_16967,N_11661,N_6755);
nand U16968 (N_16968,N_9912,N_10055);
or U16969 (N_16969,N_7425,N_11297);
and U16970 (N_16970,N_9276,N_7927);
nand U16971 (N_16971,N_9274,N_6801);
and U16972 (N_16972,N_11629,N_6519);
xnor U16973 (N_16973,N_8163,N_7779);
xor U16974 (N_16974,N_6386,N_7460);
xnor U16975 (N_16975,N_8442,N_8395);
xnor U16976 (N_16976,N_11607,N_10204);
nand U16977 (N_16977,N_10807,N_11279);
and U16978 (N_16978,N_7731,N_10911);
nor U16979 (N_16979,N_8050,N_10514);
or U16980 (N_16980,N_10127,N_8003);
or U16981 (N_16981,N_6537,N_7258);
and U16982 (N_16982,N_10004,N_10429);
xor U16983 (N_16983,N_11532,N_7832);
nand U16984 (N_16984,N_8475,N_10441);
xor U16985 (N_16985,N_8370,N_9817);
nand U16986 (N_16986,N_8340,N_11897);
nor U16987 (N_16987,N_9620,N_8943);
and U16988 (N_16988,N_9419,N_11761);
and U16989 (N_16989,N_8594,N_10239);
nor U16990 (N_16990,N_9545,N_7041);
nand U16991 (N_16991,N_8813,N_9474);
xor U16992 (N_16992,N_6074,N_8590);
and U16993 (N_16993,N_10666,N_6458);
nand U16994 (N_16994,N_9731,N_7170);
nor U16995 (N_16995,N_11204,N_6176);
nor U16996 (N_16996,N_7675,N_6060);
and U16997 (N_16997,N_8424,N_6641);
xnor U16998 (N_16998,N_6776,N_7818);
xnor U16999 (N_16999,N_11098,N_11494);
nand U17000 (N_17000,N_6742,N_7477);
and U17001 (N_17001,N_9266,N_6990);
nand U17002 (N_17002,N_6463,N_9073);
or U17003 (N_17003,N_10037,N_9722);
nand U17004 (N_17004,N_10694,N_8951);
and U17005 (N_17005,N_10772,N_7094);
xor U17006 (N_17006,N_8531,N_11826);
xnor U17007 (N_17007,N_9390,N_6965);
nand U17008 (N_17008,N_7232,N_6016);
and U17009 (N_17009,N_10117,N_9365);
xnor U17010 (N_17010,N_11638,N_9237);
or U17011 (N_17011,N_8586,N_10543);
and U17012 (N_17012,N_9819,N_6334);
nand U17013 (N_17013,N_10416,N_10832);
nand U17014 (N_17014,N_11584,N_7203);
xor U17015 (N_17015,N_7138,N_8987);
xnor U17016 (N_17016,N_11041,N_8631);
nor U17017 (N_17017,N_8485,N_10192);
xnor U17018 (N_17018,N_10410,N_8645);
nor U17019 (N_17019,N_7961,N_11251);
nor U17020 (N_17020,N_11198,N_8689);
xor U17021 (N_17021,N_6269,N_7609);
nand U17022 (N_17022,N_8082,N_11963);
or U17023 (N_17023,N_9689,N_11670);
or U17024 (N_17024,N_10479,N_11816);
xnor U17025 (N_17025,N_9498,N_8160);
nor U17026 (N_17026,N_6893,N_7573);
and U17027 (N_17027,N_6134,N_9180);
and U17028 (N_17028,N_8647,N_8741);
and U17029 (N_17029,N_7817,N_11989);
and U17030 (N_17030,N_11243,N_6640);
and U17031 (N_17031,N_8455,N_6964);
nand U17032 (N_17032,N_10599,N_9274);
or U17033 (N_17033,N_9531,N_11582);
nor U17034 (N_17034,N_7761,N_7175);
nor U17035 (N_17035,N_6907,N_8513);
xnor U17036 (N_17036,N_10583,N_8736);
xor U17037 (N_17037,N_10546,N_10719);
nor U17038 (N_17038,N_6084,N_6192);
xor U17039 (N_17039,N_6683,N_10027);
or U17040 (N_17040,N_8548,N_9940);
nand U17041 (N_17041,N_10936,N_9342);
and U17042 (N_17042,N_6670,N_7239);
xnor U17043 (N_17043,N_8585,N_9005);
or U17044 (N_17044,N_10377,N_9406);
nor U17045 (N_17045,N_10132,N_10823);
or U17046 (N_17046,N_9336,N_8012);
nor U17047 (N_17047,N_11605,N_6447);
xnor U17048 (N_17048,N_7489,N_9730);
and U17049 (N_17049,N_7291,N_11567);
or U17050 (N_17050,N_6193,N_9452);
and U17051 (N_17051,N_10077,N_11940);
or U17052 (N_17052,N_9654,N_10428);
nor U17053 (N_17053,N_10923,N_9968);
xnor U17054 (N_17054,N_9704,N_7708);
nor U17055 (N_17055,N_9797,N_9266);
or U17056 (N_17056,N_7974,N_11200);
or U17057 (N_17057,N_7169,N_10994);
or U17058 (N_17058,N_8644,N_10824);
nand U17059 (N_17059,N_6226,N_11318);
or U17060 (N_17060,N_10205,N_11141);
nand U17061 (N_17061,N_6718,N_10589);
or U17062 (N_17062,N_6412,N_7996);
xor U17063 (N_17063,N_6828,N_11596);
nand U17064 (N_17064,N_11170,N_6728);
xor U17065 (N_17065,N_8427,N_10299);
nand U17066 (N_17066,N_11766,N_7662);
xor U17067 (N_17067,N_11275,N_6820);
nor U17068 (N_17068,N_6340,N_11536);
nand U17069 (N_17069,N_9562,N_7505);
and U17070 (N_17070,N_6532,N_6582);
nand U17071 (N_17071,N_7759,N_11616);
xor U17072 (N_17072,N_11967,N_9021);
xor U17073 (N_17073,N_8197,N_10154);
nor U17074 (N_17074,N_8150,N_7644);
and U17075 (N_17075,N_6074,N_6911);
xor U17076 (N_17076,N_9438,N_9456);
xnor U17077 (N_17077,N_7989,N_7936);
nand U17078 (N_17078,N_6394,N_7623);
nor U17079 (N_17079,N_8019,N_8245);
xor U17080 (N_17080,N_9686,N_7404);
and U17081 (N_17081,N_6271,N_6798);
and U17082 (N_17082,N_7180,N_11437);
and U17083 (N_17083,N_11250,N_8851);
nand U17084 (N_17084,N_11222,N_7521);
xnor U17085 (N_17085,N_7416,N_8763);
and U17086 (N_17086,N_8163,N_8884);
nor U17087 (N_17087,N_8155,N_11011);
or U17088 (N_17088,N_10494,N_8487);
nor U17089 (N_17089,N_8621,N_10002);
nor U17090 (N_17090,N_11221,N_7384);
or U17091 (N_17091,N_11955,N_7336);
xnor U17092 (N_17092,N_7641,N_9984);
nand U17093 (N_17093,N_7631,N_8769);
and U17094 (N_17094,N_10380,N_7473);
xnor U17095 (N_17095,N_9096,N_6612);
xor U17096 (N_17096,N_7651,N_11546);
nand U17097 (N_17097,N_8791,N_7105);
and U17098 (N_17098,N_6817,N_7446);
or U17099 (N_17099,N_10501,N_7296);
nor U17100 (N_17100,N_6476,N_6958);
nand U17101 (N_17101,N_11374,N_7768);
or U17102 (N_17102,N_7190,N_8802);
or U17103 (N_17103,N_7341,N_10285);
or U17104 (N_17104,N_6432,N_10337);
nor U17105 (N_17105,N_11677,N_7938);
xnor U17106 (N_17106,N_9692,N_8271);
nand U17107 (N_17107,N_11588,N_9551);
xnor U17108 (N_17108,N_10700,N_10954);
or U17109 (N_17109,N_7282,N_9196);
nand U17110 (N_17110,N_10412,N_7915);
and U17111 (N_17111,N_9853,N_8450);
nor U17112 (N_17112,N_7973,N_8907);
and U17113 (N_17113,N_11960,N_10012);
nor U17114 (N_17114,N_8061,N_10690);
nand U17115 (N_17115,N_9260,N_10750);
xor U17116 (N_17116,N_11353,N_8850);
nand U17117 (N_17117,N_7395,N_9217);
or U17118 (N_17118,N_10432,N_8135);
and U17119 (N_17119,N_6663,N_9588);
or U17120 (N_17120,N_8993,N_8987);
nor U17121 (N_17121,N_9781,N_9863);
and U17122 (N_17122,N_11416,N_10494);
nand U17123 (N_17123,N_11019,N_11954);
nor U17124 (N_17124,N_6432,N_11587);
nor U17125 (N_17125,N_11686,N_8871);
nand U17126 (N_17126,N_8109,N_8682);
or U17127 (N_17127,N_7908,N_7726);
nor U17128 (N_17128,N_9318,N_9026);
or U17129 (N_17129,N_7880,N_6701);
and U17130 (N_17130,N_8262,N_7195);
or U17131 (N_17131,N_8361,N_8858);
nor U17132 (N_17132,N_6918,N_8967);
nor U17133 (N_17133,N_8373,N_8022);
nand U17134 (N_17134,N_6635,N_6492);
xnor U17135 (N_17135,N_10892,N_7267);
nor U17136 (N_17136,N_11251,N_10170);
or U17137 (N_17137,N_8784,N_7420);
nor U17138 (N_17138,N_10776,N_9008);
nor U17139 (N_17139,N_9318,N_9904);
nor U17140 (N_17140,N_7124,N_8387);
and U17141 (N_17141,N_10317,N_7306);
and U17142 (N_17142,N_7157,N_10610);
nor U17143 (N_17143,N_10928,N_8035);
nand U17144 (N_17144,N_8556,N_6891);
or U17145 (N_17145,N_11248,N_7711);
xor U17146 (N_17146,N_6131,N_9053);
nand U17147 (N_17147,N_7046,N_9480);
nor U17148 (N_17148,N_7858,N_8013);
nor U17149 (N_17149,N_10950,N_11256);
nand U17150 (N_17150,N_9817,N_8225);
or U17151 (N_17151,N_9231,N_11658);
nor U17152 (N_17152,N_11520,N_8812);
xor U17153 (N_17153,N_7664,N_11761);
or U17154 (N_17154,N_9670,N_9694);
nor U17155 (N_17155,N_7112,N_8231);
nor U17156 (N_17156,N_9921,N_11820);
xor U17157 (N_17157,N_8020,N_10367);
and U17158 (N_17158,N_11775,N_9634);
or U17159 (N_17159,N_8426,N_8428);
and U17160 (N_17160,N_8164,N_6982);
nor U17161 (N_17161,N_9146,N_10395);
nand U17162 (N_17162,N_6799,N_11380);
or U17163 (N_17163,N_11570,N_11166);
nand U17164 (N_17164,N_11912,N_7764);
nor U17165 (N_17165,N_11166,N_9530);
nand U17166 (N_17166,N_7738,N_8608);
nand U17167 (N_17167,N_11228,N_7869);
and U17168 (N_17168,N_7915,N_7116);
nor U17169 (N_17169,N_11904,N_10535);
nor U17170 (N_17170,N_11871,N_8902);
nor U17171 (N_17171,N_9446,N_6508);
and U17172 (N_17172,N_9221,N_9370);
nand U17173 (N_17173,N_7832,N_10054);
nor U17174 (N_17174,N_8281,N_6852);
nor U17175 (N_17175,N_8943,N_10729);
nor U17176 (N_17176,N_10734,N_7790);
nand U17177 (N_17177,N_10144,N_10094);
and U17178 (N_17178,N_9620,N_11283);
nand U17179 (N_17179,N_6656,N_9735);
xnor U17180 (N_17180,N_10572,N_6868);
or U17181 (N_17181,N_9876,N_6960);
xnor U17182 (N_17182,N_6107,N_6515);
xnor U17183 (N_17183,N_6723,N_7045);
xnor U17184 (N_17184,N_7241,N_11079);
and U17185 (N_17185,N_9574,N_10900);
nand U17186 (N_17186,N_6358,N_10358);
nor U17187 (N_17187,N_6870,N_9972);
or U17188 (N_17188,N_10041,N_7037);
nand U17189 (N_17189,N_11670,N_8242);
and U17190 (N_17190,N_10137,N_9631);
xor U17191 (N_17191,N_9167,N_6448);
nor U17192 (N_17192,N_8389,N_9669);
nand U17193 (N_17193,N_7964,N_6283);
nand U17194 (N_17194,N_10373,N_11676);
or U17195 (N_17195,N_11316,N_9044);
nor U17196 (N_17196,N_7224,N_10607);
or U17197 (N_17197,N_6486,N_8646);
or U17198 (N_17198,N_7055,N_10971);
nor U17199 (N_17199,N_7460,N_6178);
xnor U17200 (N_17200,N_10276,N_11279);
or U17201 (N_17201,N_8341,N_10854);
and U17202 (N_17202,N_9640,N_6164);
and U17203 (N_17203,N_9287,N_7606);
and U17204 (N_17204,N_7142,N_6342);
or U17205 (N_17205,N_10808,N_7094);
nor U17206 (N_17206,N_6923,N_7559);
or U17207 (N_17207,N_9135,N_6238);
xnor U17208 (N_17208,N_8597,N_9704);
or U17209 (N_17209,N_6567,N_8581);
nand U17210 (N_17210,N_6079,N_6261);
xor U17211 (N_17211,N_8504,N_8161);
and U17212 (N_17212,N_8012,N_6387);
nand U17213 (N_17213,N_7826,N_9249);
nor U17214 (N_17214,N_6969,N_9310);
xnor U17215 (N_17215,N_9912,N_8928);
nor U17216 (N_17216,N_8534,N_9084);
and U17217 (N_17217,N_10876,N_7507);
xnor U17218 (N_17218,N_7201,N_9181);
nor U17219 (N_17219,N_6625,N_7331);
nand U17220 (N_17220,N_8986,N_7953);
and U17221 (N_17221,N_9074,N_7286);
or U17222 (N_17222,N_10595,N_11476);
or U17223 (N_17223,N_8875,N_9791);
nor U17224 (N_17224,N_6714,N_9873);
and U17225 (N_17225,N_8745,N_10360);
nor U17226 (N_17226,N_10461,N_10295);
xnor U17227 (N_17227,N_8457,N_11894);
xor U17228 (N_17228,N_10502,N_8267);
nand U17229 (N_17229,N_6237,N_10064);
or U17230 (N_17230,N_9297,N_11156);
xor U17231 (N_17231,N_10327,N_8299);
xnor U17232 (N_17232,N_8742,N_9484);
nand U17233 (N_17233,N_7800,N_9808);
nand U17234 (N_17234,N_10461,N_11385);
or U17235 (N_17235,N_7151,N_11155);
and U17236 (N_17236,N_9287,N_11276);
and U17237 (N_17237,N_8125,N_8250);
xor U17238 (N_17238,N_9817,N_10718);
xnor U17239 (N_17239,N_8230,N_11418);
nand U17240 (N_17240,N_6083,N_11814);
xnor U17241 (N_17241,N_7624,N_11570);
and U17242 (N_17242,N_6419,N_8386);
nor U17243 (N_17243,N_11657,N_9336);
nand U17244 (N_17244,N_11966,N_10546);
nor U17245 (N_17245,N_8470,N_8930);
nor U17246 (N_17246,N_11686,N_7700);
nor U17247 (N_17247,N_6653,N_10105);
xor U17248 (N_17248,N_6485,N_10292);
nand U17249 (N_17249,N_8336,N_6205);
nor U17250 (N_17250,N_8422,N_8896);
or U17251 (N_17251,N_11328,N_11971);
xnor U17252 (N_17252,N_9739,N_7620);
nor U17253 (N_17253,N_8189,N_8106);
xor U17254 (N_17254,N_10837,N_8863);
and U17255 (N_17255,N_7890,N_8776);
nand U17256 (N_17256,N_8113,N_10023);
or U17257 (N_17257,N_6484,N_9890);
or U17258 (N_17258,N_10852,N_10054);
nor U17259 (N_17259,N_6815,N_8396);
xnor U17260 (N_17260,N_6947,N_7603);
and U17261 (N_17261,N_7798,N_7241);
xor U17262 (N_17262,N_8968,N_10697);
nor U17263 (N_17263,N_11763,N_7574);
nor U17264 (N_17264,N_9290,N_6671);
xnor U17265 (N_17265,N_6904,N_6887);
nor U17266 (N_17266,N_7722,N_10665);
xnor U17267 (N_17267,N_7779,N_6728);
nor U17268 (N_17268,N_11617,N_7352);
nand U17269 (N_17269,N_8536,N_9549);
xnor U17270 (N_17270,N_8048,N_9747);
nor U17271 (N_17271,N_7355,N_10796);
and U17272 (N_17272,N_10923,N_11639);
xnor U17273 (N_17273,N_9927,N_7396);
or U17274 (N_17274,N_7296,N_10365);
xor U17275 (N_17275,N_11911,N_11820);
nand U17276 (N_17276,N_7665,N_8277);
nand U17277 (N_17277,N_10053,N_8255);
and U17278 (N_17278,N_11939,N_6801);
or U17279 (N_17279,N_7989,N_6561);
or U17280 (N_17280,N_9475,N_7366);
nand U17281 (N_17281,N_10814,N_11416);
and U17282 (N_17282,N_10589,N_7048);
or U17283 (N_17283,N_7325,N_6404);
xnor U17284 (N_17284,N_8940,N_7612);
and U17285 (N_17285,N_9895,N_9664);
and U17286 (N_17286,N_8954,N_6345);
or U17287 (N_17287,N_6183,N_10527);
nand U17288 (N_17288,N_8939,N_10467);
nor U17289 (N_17289,N_9771,N_11833);
and U17290 (N_17290,N_6426,N_11788);
xnor U17291 (N_17291,N_8076,N_8836);
or U17292 (N_17292,N_6203,N_8008);
nand U17293 (N_17293,N_8961,N_9195);
nor U17294 (N_17294,N_11774,N_7828);
xor U17295 (N_17295,N_7646,N_7286);
or U17296 (N_17296,N_11382,N_7269);
or U17297 (N_17297,N_8406,N_10233);
and U17298 (N_17298,N_8407,N_6514);
nand U17299 (N_17299,N_8521,N_9177);
nor U17300 (N_17300,N_11380,N_9323);
or U17301 (N_17301,N_7912,N_10120);
and U17302 (N_17302,N_6012,N_7940);
nand U17303 (N_17303,N_7970,N_11249);
nor U17304 (N_17304,N_8375,N_9376);
xor U17305 (N_17305,N_11393,N_6787);
or U17306 (N_17306,N_8251,N_11679);
or U17307 (N_17307,N_11645,N_11928);
nand U17308 (N_17308,N_6187,N_8879);
nor U17309 (N_17309,N_6335,N_6305);
nand U17310 (N_17310,N_9395,N_8781);
and U17311 (N_17311,N_8103,N_8570);
or U17312 (N_17312,N_9609,N_9204);
xnor U17313 (N_17313,N_10670,N_9459);
nor U17314 (N_17314,N_10558,N_10108);
and U17315 (N_17315,N_6714,N_9390);
or U17316 (N_17316,N_8028,N_10787);
nand U17317 (N_17317,N_7677,N_9570);
nor U17318 (N_17318,N_7083,N_9474);
or U17319 (N_17319,N_9974,N_6352);
xnor U17320 (N_17320,N_9146,N_6641);
and U17321 (N_17321,N_10566,N_7169);
and U17322 (N_17322,N_8016,N_7413);
nand U17323 (N_17323,N_10937,N_6633);
and U17324 (N_17324,N_10486,N_8971);
nand U17325 (N_17325,N_8362,N_8748);
or U17326 (N_17326,N_9066,N_8150);
and U17327 (N_17327,N_8577,N_6272);
and U17328 (N_17328,N_10304,N_6945);
nand U17329 (N_17329,N_7948,N_11196);
and U17330 (N_17330,N_7284,N_7568);
xor U17331 (N_17331,N_10629,N_11119);
xnor U17332 (N_17332,N_9710,N_6724);
and U17333 (N_17333,N_7427,N_8995);
nand U17334 (N_17334,N_9393,N_9448);
nor U17335 (N_17335,N_11496,N_6454);
nor U17336 (N_17336,N_9330,N_6194);
and U17337 (N_17337,N_6806,N_9687);
nor U17338 (N_17338,N_11164,N_8155);
nor U17339 (N_17339,N_8275,N_8798);
xor U17340 (N_17340,N_9928,N_11178);
nand U17341 (N_17341,N_7184,N_9849);
nor U17342 (N_17342,N_10851,N_11133);
nor U17343 (N_17343,N_11568,N_6433);
or U17344 (N_17344,N_10173,N_10828);
or U17345 (N_17345,N_7617,N_8237);
nor U17346 (N_17346,N_7601,N_7398);
nand U17347 (N_17347,N_11963,N_6723);
nor U17348 (N_17348,N_8009,N_6503);
nand U17349 (N_17349,N_6284,N_9647);
and U17350 (N_17350,N_8424,N_7478);
xor U17351 (N_17351,N_9720,N_8712);
or U17352 (N_17352,N_10622,N_8976);
xor U17353 (N_17353,N_7360,N_6865);
nand U17354 (N_17354,N_6276,N_6014);
nand U17355 (N_17355,N_6016,N_9928);
and U17356 (N_17356,N_11737,N_6886);
nand U17357 (N_17357,N_8300,N_8405);
and U17358 (N_17358,N_10640,N_9182);
nand U17359 (N_17359,N_9832,N_6261);
nor U17360 (N_17360,N_11531,N_10130);
and U17361 (N_17361,N_6259,N_9921);
or U17362 (N_17362,N_7727,N_10304);
or U17363 (N_17363,N_10553,N_7546);
nor U17364 (N_17364,N_10746,N_10762);
and U17365 (N_17365,N_11814,N_8055);
or U17366 (N_17366,N_6481,N_10181);
xor U17367 (N_17367,N_10553,N_6729);
or U17368 (N_17368,N_8907,N_10031);
nor U17369 (N_17369,N_10333,N_6328);
xnor U17370 (N_17370,N_7429,N_11339);
nand U17371 (N_17371,N_7326,N_8615);
or U17372 (N_17372,N_10131,N_9608);
or U17373 (N_17373,N_8397,N_8800);
and U17374 (N_17374,N_10479,N_11537);
or U17375 (N_17375,N_8771,N_6473);
or U17376 (N_17376,N_9004,N_8839);
nor U17377 (N_17377,N_6063,N_11359);
xor U17378 (N_17378,N_9533,N_10704);
nor U17379 (N_17379,N_7126,N_11025);
nor U17380 (N_17380,N_11094,N_6972);
xor U17381 (N_17381,N_10397,N_9538);
xor U17382 (N_17382,N_8250,N_7598);
nand U17383 (N_17383,N_10949,N_8023);
and U17384 (N_17384,N_9302,N_9582);
nor U17385 (N_17385,N_7065,N_11457);
xor U17386 (N_17386,N_11887,N_9282);
nand U17387 (N_17387,N_8328,N_8229);
and U17388 (N_17388,N_10589,N_7538);
nand U17389 (N_17389,N_6637,N_7967);
and U17390 (N_17390,N_7142,N_9737);
xor U17391 (N_17391,N_10150,N_10064);
xor U17392 (N_17392,N_9760,N_11816);
or U17393 (N_17393,N_9197,N_6665);
xnor U17394 (N_17394,N_9640,N_6823);
and U17395 (N_17395,N_9679,N_7302);
and U17396 (N_17396,N_10836,N_9542);
nor U17397 (N_17397,N_6069,N_9870);
nor U17398 (N_17398,N_7026,N_10683);
xor U17399 (N_17399,N_8878,N_8040);
nor U17400 (N_17400,N_8588,N_11193);
nand U17401 (N_17401,N_10589,N_10482);
and U17402 (N_17402,N_10962,N_6928);
xor U17403 (N_17403,N_8426,N_8688);
and U17404 (N_17404,N_8957,N_7721);
and U17405 (N_17405,N_9977,N_9016);
xor U17406 (N_17406,N_10624,N_11448);
nand U17407 (N_17407,N_7644,N_11455);
xnor U17408 (N_17408,N_9949,N_10383);
xnor U17409 (N_17409,N_7161,N_9034);
or U17410 (N_17410,N_6199,N_8551);
or U17411 (N_17411,N_11608,N_7132);
and U17412 (N_17412,N_9254,N_8354);
and U17413 (N_17413,N_7981,N_6140);
and U17414 (N_17414,N_6297,N_11228);
and U17415 (N_17415,N_6007,N_11513);
nor U17416 (N_17416,N_6990,N_6159);
and U17417 (N_17417,N_8462,N_10621);
nor U17418 (N_17418,N_9766,N_6370);
nand U17419 (N_17419,N_10139,N_9351);
or U17420 (N_17420,N_8470,N_9936);
xnor U17421 (N_17421,N_11426,N_7954);
xor U17422 (N_17422,N_10449,N_9474);
xor U17423 (N_17423,N_9228,N_11257);
nor U17424 (N_17424,N_10165,N_8926);
nand U17425 (N_17425,N_11557,N_6775);
nand U17426 (N_17426,N_6699,N_6382);
xnor U17427 (N_17427,N_7037,N_7714);
or U17428 (N_17428,N_9584,N_6831);
or U17429 (N_17429,N_6652,N_10712);
or U17430 (N_17430,N_11472,N_9589);
nor U17431 (N_17431,N_8051,N_9119);
nor U17432 (N_17432,N_10493,N_6233);
xnor U17433 (N_17433,N_8745,N_8721);
xnor U17434 (N_17434,N_8518,N_6694);
and U17435 (N_17435,N_7249,N_9375);
and U17436 (N_17436,N_11731,N_9661);
nor U17437 (N_17437,N_9298,N_11664);
or U17438 (N_17438,N_10295,N_10736);
and U17439 (N_17439,N_10326,N_10325);
or U17440 (N_17440,N_6962,N_11754);
and U17441 (N_17441,N_8027,N_10735);
or U17442 (N_17442,N_8478,N_10036);
and U17443 (N_17443,N_10911,N_11261);
nor U17444 (N_17444,N_8290,N_8080);
xor U17445 (N_17445,N_8366,N_7461);
nor U17446 (N_17446,N_8171,N_7548);
nand U17447 (N_17447,N_10700,N_9095);
nor U17448 (N_17448,N_10336,N_8687);
xnor U17449 (N_17449,N_9427,N_8814);
nor U17450 (N_17450,N_8148,N_8380);
nand U17451 (N_17451,N_10299,N_9400);
and U17452 (N_17452,N_10870,N_9437);
nor U17453 (N_17453,N_8929,N_6896);
nor U17454 (N_17454,N_11400,N_6981);
and U17455 (N_17455,N_11270,N_6165);
nor U17456 (N_17456,N_7908,N_11196);
or U17457 (N_17457,N_7447,N_10714);
nand U17458 (N_17458,N_8443,N_7539);
or U17459 (N_17459,N_11120,N_9747);
nand U17460 (N_17460,N_7974,N_11560);
nor U17461 (N_17461,N_7921,N_11878);
nor U17462 (N_17462,N_6067,N_11832);
nand U17463 (N_17463,N_9147,N_11167);
nor U17464 (N_17464,N_8964,N_10236);
nand U17465 (N_17465,N_8667,N_8029);
and U17466 (N_17466,N_6372,N_9207);
nand U17467 (N_17467,N_6695,N_7027);
nor U17468 (N_17468,N_8790,N_6772);
or U17469 (N_17469,N_6896,N_10936);
or U17470 (N_17470,N_11422,N_10488);
and U17471 (N_17471,N_8333,N_9511);
nand U17472 (N_17472,N_11511,N_6709);
nor U17473 (N_17473,N_6038,N_11279);
xor U17474 (N_17474,N_8202,N_8410);
nor U17475 (N_17475,N_10817,N_7283);
nor U17476 (N_17476,N_9245,N_8187);
xor U17477 (N_17477,N_10700,N_9220);
nand U17478 (N_17478,N_9985,N_7501);
or U17479 (N_17479,N_9444,N_10754);
xnor U17480 (N_17480,N_7398,N_11623);
nor U17481 (N_17481,N_10805,N_11648);
nand U17482 (N_17482,N_9596,N_8840);
xnor U17483 (N_17483,N_10206,N_7614);
nand U17484 (N_17484,N_6153,N_6684);
nor U17485 (N_17485,N_9563,N_9165);
xnor U17486 (N_17486,N_8348,N_6031);
or U17487 (N_17487,N_9220,N_8518);
nor U17488 (N_17488,N_6080,N_7525);
or U17489 (N_17489,N_9237,N_9801);
and U17490 (N_17490,N_11246,N_7049);
nor U17491 (N_17491,N_11170,N_9735);
nand U17492 (N_17492,N_6686,N_7281);
nor U17493 (N_17493,N_7577,N_9923);
nor U17494 (N_17494,N_6469,N_11339);
nor U17495 (N_17495,N_11600,N_10279);
and U17496 (N_17496,N_8527,N_9953);
nor U17497 (N_17497,N_9843,N_10011);
xor U17498 (N_17498,N_11263,N_6481);
and U17499 (N_17499,N_11416,N_11496);
or U17500 (N_17500,N_7498,N_11418);
nand U17501 (N_17501,N_9347,N_8828);
nor U17502 (N_17502,N_10094,N_9719);
nor U17503 (N_17503,N_10513,N_7731);
or U17504 (N_17504,N_6077,N_7319);
xnor U17505 (N_17505,N_11072,N_11600);
nand U17506 (N_17506,N_8258,N_11517);
nor U17507 (N_17507,N_9335,N_7046);
xor U17508 (N_17508,N_7083,N_10547);
xnor U17509 (N_17509,N_10769,N_11680);
or U17510 (N_17510,N_11609,N_6210);
nor U17511 (N_17511,N_7777,N_8222);
nor U17512 (N_17512,N_7187,N_11047);
or U17513 (N_17513,N_6406,N_10816);
nor U17514 (N_17514,N_6304,N_6556);
xor U17515 (N_17515,N_9839,N_8754);
or U17516 (N_17516,N_9485,N_11579);
and U17517 (N_17517,N_7967,N_8295);
and U17518 (N_17518,N_9516,N_11667);
nor U17519 (N_17519,N_8331,N_11035);
or U17520 (N_17520,N_7521,N_9434);
nor U17521 (N_17521,N_8775,N_9946);
xnor U17522 (N_17522,N_9489,N_9123);
or U17523 (N_17523,N_11157,N_11316);
nand U17524 (N_17524,N_11137,N_9409);
nor U17525 (N_17525,N_6343,N_8206);
or U17526 (N_17526,N_10344,N_8423);
and U17527 (N_17527,N_6799,N_11862);
nor U17528 (N_17528,N_7499,N_8051);
and U17529 (N_17529,N_11478,N_10992);
or U17530 (N_17530,N_6776,N_10813);
nor U17531 (N_17531,N_7862,N_7155);
nor U17532 (N_17532,N_8997,N_7747);
xnor U17533 (N_17533,N_8658,N_11321);
and U17534 (N_17534,N_7112,N_10571);
and U17535 (N_17535,N_6462,N_8356);
xnor U17536 (N_17536,N_6602,N_9767);
and U17537 (N_17537,N_11457,N_8414);
xnor U17538 (N_17538,N_6736,N_10141);
or U17539 (N_17539,N_6788,N_6289);
and U17540 (N_17540,N_7002,N_7735);
nand U17541 (N_17541,N_10916,N_8167);
xnor U17542 (N_17542,N_7642,N_9752);
or U17543 (N_17543,N_9607,N_10242);
nand U17544 (N_17544,N_7469,N_10632);
and U17545 (N_17545,N_11606,N_6397);
nor U17546 (N_17546,N_11358,N_9069);
nor U17547 (N_17547,N_9447,N_10045);
xnor U17548 (N_17548,N_7671,N_10909);
xnor U17549 (N_17549,N_11812,N_7351);
nand U17550 (N_17550,N_9814,N_10034);
and U17551 (N_17551,N_7970,N_6696);
nand U17552 (N_17552,N_7498,N_10996);
xor U17553 (N_17553,N_6094,N_7168);
xnor U17554 (N_17554,N_6751,N_11532);
and U17555 (N_17555,N_11659,N_7030);
xnor U17556 (N_17556,N_9006,N_6994);
nor U17557 (N_17557,N_10854,N_7045);
nand U17558 (N_17558,N_9657,N_8022);
nor U17559 (N_17559,N_8616,N_10788);
xnor U17560 (N_17560,N_6234,N_10728);
nor U17561 (N_17561,N_10956,N_6341);
nand U17562 (N_17562,N_6889,N_9245);
or U17563 (N_17563,N_9607,N_8686);
nand U17564 (N_17564,N_6088,N_9564);
nor U17565 (N_17565,N_11446,N_11868);
or U17566 (N_17566,N_11162,N_6069);
or U17567 (N_17567,N_9936,N_7669);
or U17568 (N_17568,N_6223,N_11405);
xnor U17569 (N_17569,N_10025,N_10748);
or U17570 (N_17570,N_11794,N_9995);
xor U17571 (N_17571,N_8126,N_11577);
or U17572 (N_17572,N_7581,N_9387);
or U17573 (N_17573,N_9504,N_8548);
xnor U17574 (N_17574,N_9461,N_9808);
and U17575 (N_17575,N_6344,N_6903);
and U17576 (N_17576,N_9292,N_10918);
nor U17577 (N_17577,N_6203,N_9933);
nor U17578 (N_17578,N_7633,N_11987);
nor U17579 (N_17579,N_6583,N_6969);
and U17580 (N_17580,N_6186,N_7124);
nand U17581 (N_17581,N_11553,N_9190);
and U17582 (N_17582,N_7096,N_7394);
and U17583 (N_17583,N_6415,N_8392);
nor U17584 (N_17584,N_6446,N_9844);
and U17585 (N_17585,N_6761,N_11673);
and U17586 (N_17586,N_8051,N_10778);
xor U17587 (N_17587,N_6907,N_6611);
or U17588 (N_17588,N_10240,N_10284);
xnor U17589 (N_17589,N_8108,N_7787);
nand U17590 (N_17590,N_11109,N_11003);
nor U17591 (N_17591,N_7135,N_8999);
or U17592 (N_17592,N_11523,N_11732);
xnor U17593 (N_17593,N_11558,N_10008);
xnor U17594 (N_17594,N_8917,N_9885);
nand U17595 (N_17595,N_7426,N_9955);
nand U17596 (N_17596,N_10610,N_7977);
or U17597 (N_17597,N_7879,N_10283);
xor U17598 (N_17598,N_7922,N_9320);
xor U17599 (N_17599,N_8023,N_7219);
nor U17600 (N_17600,N_8972,N_6467);
nand U17601 (N_17601,N_8408,N_9871);
and U17602 (N_17602,N_6381,N_6263);
and U17603 (N_17603,N_6123,N_10314);
and U17604 (N_17604,N_10104,N_8233);
nand U17605 (N_17605,N_6349,N_6433);
or U17606 (N_17606,N_11542,N_9435);
nor U17607 (N_17607,N_6449,N_6648);
or U17608 (N_17608,N_8903,N_6197);
nand U17609 (N_17609,N_8060,N_6217);
nor U17610 (N_17610,N_9510,N_10544);
xor U17611 (N_17611,N_9273,N_8740);
xnor U17612 (N_17612,N_11017,N_10648);
nor U17613 (N_17613,N_9745,N_10490);
nor U17614 (N_17614,N_6049,N_7661);
nor U17615 (N_17615,N_10896,N_11415);
nand U17616 (N_17616,N_9876,N_6028);
xor U17617 (N_17617,N_8007,N_7002);
and U17618 (N_17618,N_9646,N_6466);
and U17619 (N_17619,N_7899,N_10015);
or U17620 (N_17620,N_11768,N_8723);
xnor U17621 (N_17621,N_9288,N_10890);
nor U17622 (N_17622,N_8520,N_6333);
nor U17623 (N_17623,N_11309,N_9669);
or U17624 (N_17624,N_10051,N_11388);
xor U17625 (N_17625,N_11438,N_9998);
nand U17626 (N_17626,N_7363,N_10315);
xor U17627 (N_17627,N_7194,N_11109);
nand U17628 (N_17628,N_8096,N_11298);
nor U17629 (N_17629,N_10987,N_6625);
or U17630 (N_17630,N_10565,N_7345);
nor U17631 (N_17631,N_10152,N_10146);
nor U17632 (N_17632,N_11405,N_9007);
or U17633 (N_17633,N_10667,N_8786);
xnor U17634 (N_17634,N_7232,N_8202);
and U17635 (N_17635,N_9359,N_9044);
xor U17636 (N_17636,N_7167,N_6368);
or U17637 (N_17637,N_10260,N_8931);
xor U17638 (N_17638,N_11741,N_9803);
or U17639 (N_17639,N_11092,N_6560);
nor U17640 (N_17640,N_6889,N_10271);
and U17641 (N_17641,N_7129,N_8868);
and U17642 (N_17642,N_7812,N_11305);
or U17643 (N_17643,N_8612,N_9053);
nor U17644 (N_17644,N_11090,N_10448);
nor U17645 (N_17645,N_11543,N_11819);
and U17646 (N_17646,N_10687,N_10885);
and U17647 (N_17647,N_7294,N_11814);
nor U17648 (N_17648,N_9601,N_11204);
or U17649 (N_17649,N_7844,N_6227);
xor U17650 (N_17650,N_10738,N_10374);
or U17651 (N_17651,N_11794,N_8881);
xnor U17652 (N_17652,N_11115,N_6659);
nand U17653 (N_17653,N_8095,N_7383);
or U17654 (N_17654,N_9157,N_6219);
xnor U17655 (N_17655,N_8184,N_8900);
nand U17656 (N_17656,N_10073,N_11428);
or U17657 (N_17657,N_6094,N_9328);
xor U17658 (N_17658,N_6804,N_9036);
and U17659 (N_17659,N_6338,N_6712);
and U17660 (N_17660,N_7557,N_11785);
nor U17661 (N_17661,N_10881,N_8794);
nor U17662 (N_17662,N_9321,N_7453);
xor U17663 (N_17663,N_7546,N_11583);
xor U17664 (N_17664,N_10610,N_6606);
or U17665 (N_17665,N_9337,N_10970);
nor U17666 (N_17666,N_10798,N_7178);
or U17667 (N_17667,N_7458,N_7233);
xor U17668 (N_17668,N_8327,N_8105);
nor U17669 (N_17669,N_6563,N_10489);
xor U17670 (N_17670,N_7653,N_6031);
nor U17671 (N_17671,N_9333,N_10208);
nor U17672 (N_17672,N_11358,N_9934);
or U17673 (N_17673,N_11056,N_8113);
xnor U17674 (N_17674,N_9740,N_6328);
or U17675 (N_17675,N_9026,N_6624);
and U17676 (N_17676,N_11766,N_9661);
nor U17677 (N_17677,N_10122,N_9184);
xor U17678 (N_17678,N_8871,N_10122);
or U17679 (N_17679,N_6729,N_7190);
nand U17680 (N_17680,N_10143,N_10582);
and U17681 (N_17681,N_8088,N_11539);
and U17682 (N_17682,N_10075,N_8552);
or U17683 (N_17683,N_6793,N_7243);
xnor U17684 (N_17684,N_7280,N_10474);
nor U17685 (N_17685,N_10729,N_6998);
and U17686 (N_17686,N_8136,N_9816);
xor U17687 (N_17687,N_10301,N_8804);
nand U17688 (N_17688,N_11785,N_6053);
nor U17689 (N_17689,N_8855,N_10426);
xnor U17690 (N_17690,N_11311,N_8940);
or U17691 (N_17691,N_10648,N_10383);
and U17692 (N_17692,N_10063,N_8905);
or U17693 (N_17693,N_9215,N_8246);
xor U17694 (N_17694,N_8439,N_8341);
nor U17695 (N_17695,N_7874,N_8531);
xnor U17696 (N_17696,N_10165,N_10905);
or U17697 (N_17697,N_11318,N_10930);
nor U17698 (N_17698,N_11495,N_6686);
or U17699 (N_17699,N_7841,N_6434);
or U17700 (N_17700,N_8009,N_7897);
and U17701 (N_17701,N_6365,N_11462);
nand U17702 (N_17702,N_9498,N_11349);
and U17703 (N_17703,N_10580,N_7992);
nand U17704 (N_17704,N_7928,N_7179);
nor U17705 (N_17705,N_11126,N_11299);
nor U17706 (N_17706,N_7298,N_6937);
or U17707 (N_17707,N_7143,N_11814);
or U17708 (N_17708,N_8036,N_8463);
xor U17709 (N_17709,N_9058,N_11582);
and U17710 (N_17710,N_9710,N_6249);
and U17711 (N_17711,N_9159,N_7441);
and U17712 (N_17712,N_9281,N_6517);
nand U17713 (N_17713,N_9889,N_6774);
and U17714 (N_17714,N_7120,N_8577);
and U17715 (N_17715,N_11152,N_10256);
or U17716 (N_17716,N_8731,N_10637);
nand U17717 (N_17717,N_8463,N_11857);
nor U17718 (N_17718,N_9367,N_8649);
and U17719 (N_17719,N_11241,N_10203);
and U17720 (N_17720,N_6968,N_6173);
xor U17721 (N_17721,N_6656,N_8213);
nand U17722 (N_17722,N_6862,N_8620);
or U17723 (N_17723,N_9292,N_9399);
and U17724 (N_17724,N_11144,N_6940);
nand U17725 (N_17725,N_8193,N_10758);
xnor U17726 (N_17726,N_8006,N_7902);
nor U17727 (N_17727,N_10687,N_9046);
or U17728 (N_17728,N_10966,N_11773);
or U17729 (N_17729,N_11732,N_7285);
and U17730 (N_17730,N_11582,N_11201);
xnor U17731 (N_17731,N_7693,N_7182);
nand U17732 (N_17732,N_11806,N_6561);
and U17733 (N_17733,N_10777,N_6010);
or U17734 (N_17734,N_10176,N_11041);
and U17735 (N_17735,N_10912,N_10987);
nor U17736 (N_17736,N_6232,N_11075);
nor U17737 (N_17737,N_6597,N_9416);
nor U17738 (N_17738,N_9789,N_6988);
nand U17739 (N_17739,N_6428,N_8306);
nand U17740 (N_17740,N_9032,N_7305);
and U17741 (N_17741,N_9316,N_8634);
xnor U17742 (N_17742,N_9984,N_6524);
and U17743 (N_17743,N_8120,N_6549);
and U17744 (N_17744,N_10045,N_6660);
or U17745 (N_17745,N_11371,N_6181);
nand U17746 (N_17746,N_7117,N_8979);
nor U17747 (N_17747,N_9917,N_6720);
nor U17748 (N_17748,N_10134,N_6477);
and U17749 (N_17749,N_10861,N_6576);
xnor U17750 (N_17750,N_6427,N_7819);
xor U17751 (N_17751,N_10950,N_9658);
and U17752 (N_17752,N_6491,N_11270);
nor U17753 (N_17753,N_10520,N_6995);
nor U17754 (N_17754,N_9395,N_8116);
xnor U17755 (N_17755,N_8033,N_9898);
nor U17756 (N_17756,N_11731,N_7988);
xor U17757 (N_17757,N_11349,N_9204);
xor U17758 (N_17758,N_7655,N_10651);
or U17759 (N_17759,N_10946,N_8229);
nand U17760 (N_17760,N_9928,N_8986);
and U17761 (N_17761,N_7595,N_9581);
and U17762 (N_17762,N_10568,N_8422);
xor U17763 (N_17763,N_10652,N_6645);
or U17764 (N_17764,N_11732,N_8084);
and U17765 (N_17765,N_10967,N_8267);
and U17766 (N_17766,N_8510,N_10496);
and U17767 (N_17767,N_8771,N_10989);
nor U17768 (N_17768,N_8107,N_8776);
xor U17769 (N_17769,N_8631,N_9670);
and U17770 (N_17770,N_10306,N_6130);
nand U17771 (N_17771,N_6761,N_11627);
nor U17772 (N_17772,N_11370,N_10903);
and U17773 (N_17773,N_11559,N_11221);
nand U17774 (N_17774,N_10659,N_8920);
nand U17775 (N_17775,N_6281,N_10505);
and U17776 (N_17776,N_9741,N_7752);
nand U17777 (N_17777,N_8103,N_10031);
nand U17778 (N_17778,N_7524,N_6302);
xor U17779 (N_17779,N_6732,N_9388);
nor U17780 (N_17780,N_6488,N_8459);
or U17781 (N_17781,N_11982,N_8737);
nand U17782 (N_17782,N_8482,N_7432);
nand U17783 (N_17783,N_7927,N_7262);
and U17784 (N_17784,N_8467,N_6908);
nor U17785 (N_17785,N_9308,N_8469);
nor U17786 (N_17786,N_11155,N_7954);
xor U17787 (N_17787,N_9308,N_10094);
xnor U17788 (N_17788,N_7946,N_10733);
and U17789 (N_17789,N_11270,N_8895);
nand U17790 (N_17790,N_10189,N_7714);
nand U17791 (N_17791,N_8634,N_6112);
nand U17792 (N_17792,N_7124,N_6099);
nor U17793 (N_17793,N_6656,N_10503);
xnor U17794 (N_17794,N_9647,N_7162);
nand U17795 (N_17795,N_10701,N_6757);
xor U17796 (N_17796,N_6975,N_6863);
xnor U17797 (N_17797,N_6425,N_10430);
nor U17798 (N_17798,N_6601,N_6222);
nand U17799 (N_17799,N_9575,N_6601);
or U17800 (N_17800,N_6810,N_9026);
or U17801 (N_17801,N_8183,N_10554);
nand U17802 (N_17802,N_11548,N_10606);
or U17803 (N_17803,N_7452,N_10381);
or U17804 (N_17804,N_10936,N_11720);
xor U17805 (N_17805,N_10644,N_9145);
and U17806 (N_17806,N_8065,N_11811);
nor U17807 (N_17807,N_7151,N_10136);
xor U17808 (N_17808,N_10261,N_11026);
nand U17809 (N_17809,N_11466,N_8657);
or U17810 (N_17810,N_11879,N_8281);
or U17811 (N_17811,N_8861,N_7348);
or U17812 (N_17812,N_8081,N_8920);
nor U17813 (N_17813,N_10337,N_10320);
and U17814 (N_17814,N_8924,N_9312);
and U17815 (N_17815,N_7637,N_9691);
nand U17816 (N_17816,N_11979,N_7998);
nor U17817 (N_17817,N_7397,N_8749);
nor U17818 (N_17818,N_8559,N_6829);
or U17819 (N_17819,N_6451,N_10882);
nor U17820 (N_17820,N_8244,N_10936);
nor U17821 (N_17821,N_11851,N_6035);
xnor U17822 (N_17822,N_10768,N_10245);
or U17823 (N_17823,N_10109,N_10438);
nand U17824 (N_17824,N_10075,N_8411);
or U17825 (N_17825,N_9281,N_9966);
nand U17826 (N_17826,N_10555,N_10210);
and U17827 (N_17827,N_7165,N_10654);
and U17828 (N_17828,N_6039,N_6612);
and U17829 (N_17829,N_6585,N_8626);
nor U17830 (N_17830,N_10667,N_9293);
and U17831 (N_17831,N_11569,N_10169);
xor U17832 (N_17832,N_10613,N_8592);
or U17833 (N_17833,N_9362,N_7570);
and U17834 (N_17834,N_7123,N_7605);
nor U17835 (N_17835,N_6118,N_8698);
nand U17836 (N_17836,N_11941,N_8442);
or U17837 (N_17837,N_8789,N_10642);
xor U17838 (N_17838,N_7077,N_10971);
nand U17839 (N_17839,N_6943,N_10431);
xor U17840 (N_17840,N_9213,N_10344);
or U17841 (N_17841,N_6566,N_9406);
nor U17842 (N_17842,N_11493,N_8920);
and U17843 (N_17843,N_11672,N_6498);
nand U17844 (N_17844,N_11790,N_7420);
xnor U17845 (N_17845,N_10916,N_10364);
nor U17846 (N_17846,N_6907,N_8371);
nand U17847 (N_17847,N_9794,N_6294);
nand U17848 (N_17848,N_8624,N_6809);
nand U17849 (N_17849,N_8371,N_11122);
nor U17850 (N_17850,N_7320,N_10626);
or U17851 (N_17851,N_11338,N_6596);
or U17852 (N_17852,N_11419,N_10783);
nor U17853 (N_17853,N_9467,N_7143);
nand U17854 (N_17854,N_10791,N_8946);
xnor U17855 (N_17855,N_6625,N_8646);
nand U17856 (N_17856,N_6531,N_11971);
and U17857 (N_17857,N_11890,N_8919);
or U17858 (N_17858,N_9327,N_10208);
xnor U17859 (N_17859,N_10821,N_11223);
or U17860 (N_17860,N_8980,N_7212);
nor U17861 (N_17861,N_9194,N_8936);
xor U17862 (N_17862,N_10081,N_9604);
xor U17863 (N_17863,N_9204,N_11389);
nor U17864 (N_17864,N_11092,N_8162);
xnor U17865 (N_17865,N_6715,N_9963);
and U17866 (N_17866,N_9713,N_6531);
or U17867 (N_17867,N_11717,N_6914);
and U17868 (N_17868,N_9900,N_8719);
nor U17869 (N_17869,N_11853,N_11324);
nand U17870 (N_17870,N_6008,N_9006);
nand U17871 (N_17871,N_6750,N_9028);
nor U17872 (N_17872,N_6479,N_10023);
and U17873 (N_17873,N_8365,N_9887);
and U17874 (N_17874,N_6540,N_10255);
and U17875 (N_17875,N_6986,N_10400);
nand U17876 (N_17876,N_9572,N_10451);
xor U17877 (N_17877,N_7740,N_9745);
or U17878 (N_17878,N_10895,N_7304);
nand U17879 (N_17879,N_6365,N_10899);
nor U17880 (N_17880,N_7642,N_10954);
xor U17881 (N_17881,N_9258,N_6617);
nor U17882 (N_17882,N_9655,N_10910);
and U17883 (N_17883,N_7792,N_9685);
xor U17884 (N_17884,N_10476,N_11845);
or U17885 (N_17885,N_7679,N_6263);
and U17886 (N_17886,N_8536,N_11507);
or U17887 (N_17887,N_11233,N_7329);
nand U17888 (N_17888,N_9582,N_6529);
nor U17889 (N_17889,N_10092,N_6339);
xnor U17890 (N_17890,N_6257,N_6614);
xnor U17891 (N_17891,N_8146,N_9521);
and U17892 (N_17892,N_8033,N_7705);
xor U17893 (N_17893,N_7560,N_10748);
and U17894 (N_17894,N_6835,N_6878);
nor U17895 (N_17895,N_6641,N_7625);
xor U17896 (N_17896,N_7183,N_7130);
xnor U17897 (N_17897,N_6519,N_10938);
and U17898 (N_17898,N_8835,N_11643);
nand U17899 (N_17899,N_9015,N_11573);
nor U17900 (N_17900,N_6328,N_8063);
xnor U17901 (N_17901,N_9865,N_7273);
or U17902 (N_17902,N_7960,N_11075);
nand U17903 (N_17903,N_8054,N_10837);
or U17904 (N_17904,N_10231,N_8782);
and U17905 (N_17905,N_11644,N_7785);
or U17906 (N_17906,N_10001,N_9483);
nand U17907 (N_17907,N_8346,N_11566);
xnor U17908 (N_17908,N_10336,N_8826);
xnor U17909 (N_17909,N_11577,N_10849);
xor U17910 (N_17910,N_11217,N_10952);
and U17911 (N_17911,N_9130,N_10881);
xnor U17912 (N_17912,N_8744,N_10875);
nand U17913 (N_17913,N_10539,N_6229);
and U17914 (N_17914,N_6268,N_8944);
xor U17915 (N_17915,N_11760,N_11420);
xnor U17916 (N_17916,N_8870,N_9029);
nor U17917 (N_17917,N_6255,N_10429);
nand U17918 (N_17918,N_10404,N_11143);
nand U17919 (N_17919,N_10174,N_7109);
xnor U17920 (N_17920,N_10165,N_11920);
and U17921 (N_17921,N_11437,N_7164);
or U17922 (N_17922,N_6599,N_9391);
xor U17923 (N_17923,N_7537,N_6871);
or U17924 (N_17924,N_9255,N_11137);
or U17925 (N_17925,N_7175,N_11474);
nand U17926 (N_17926,N_10414,N_7613);
or U17927 (N_17927,N_6494,N_6966);
xnor U17928 (N_17928,N_10492,N_9969);
xnor U17929 (N_17929,N_9373,N_8268);
nand U17930 (N_17930,N_10728,N_10203);
or U17931 (N_17931,N_7995,N_10880);
nor U17932 (N_17932,N_6650,N_7954);
nand U17933 (N_17933,N_10543,N_9782);
nand U17934 (N_17934,N_8234,N_10623);
xor U17935 (N_17935,N_10189,N_8328);
or U17936 (N_17936,N_7985,N_11124);
nor U17937 (N_17937,N_9670,N_6763);
nand U17938 (N_17938,N_10584,N_8597);
or U17939 (N_17939,N_8775,N_7113);
xor U17940 (N_17940,N_10377,N_7120);
xnor U17941 (N_17941,N_7282,N_8570);
nand U17942 (N_17942,N_9346,N_9499);
or U17943 (N_17943,N_10206,N_8086);
and U17944 (N_17944,N_6037,N_7504);
nand U17945 (N_17945,N_9849,N_6012);
and U17946 (N_17946,N_11462,N_6839);
nor U17947 (N_17947,N_9168,N_7880);
nand U17948 (N_17948,N_10717,N_7624);
and U17949 (N_17949,N_9941,N_11518);
nand U17950 (N_17950,N_8055,N_8494);
xnor U17951 (N_17951,N_9959,N_8819);
or U17952 (N_17952,N_9173,N_11334);
and U17953 (N_17953,N_9075,N_7455);
nor U17954 (N_17954,N_11980,N_11102);
xnor U17955 (N_17955,N_8598,N_11528);
and U17956 (N_17956,N_10865,N_11410);
nor U17957 (N_17957,N_6938,N_9941);
or U17958 (N_17958,N_8088,N_11397);
nand U17959 (N_17959,N_11936,N_7841);
and U17960 (N_17960,N_9265,N_10931);
or U17961 (N_17961,N_10843,N_6371);
nand U17962 (N_17962,N_9500,N_10562);
xor U17963 (N_17963,N_11250,N_11574);
nand U17964 (N_17964,N_6248,N_8454);
xnor U17965 (N_17965,N_6487,N_9125);
and U17966 (N_17966,N_10149,N_7673);
xor U17967 (N_17967,N_9618,N_11038);
nor U17968 (N_17968,N_10566,N_6145);
xor U17969 (N_17969,N_7337,N_8950);
and U17970 (N_17970,N_11440,N_11680);
and U17971 (N_17971,N_9393,N_11018);
xor U17972 (N_17972,N_8855,N_8875);
or U17973 (N_17973,N_7242,N_9043);
or U17974 (N_17974,N_9032,N_10014);
or U17975 (N_17975,N_6693,N_6025);
or U17976 (N_17976,N_11062,N_8262);
nand U17977 (N_17977,N_10250,N_7944);
or U17978 (N_17978,N_11683,N_6560);
xor U17979 (N_17979,N_7776,N_7723);
nand U17980 (N_17980,N_6341,N_6703);
and U17981 (N_17981,N_10014,N_6106);
nand U17982 (N_17982,N_6224,N_7245);
xor U17983 (N_17983,N_6810,N_10958);
xor U17984 (N_17984,N_10846,N_10117);
and U17985 (N_17985,N_10944,N_9789);
nand U17986 (N_17986,N_9584,N_8847);
or U17987 (N_17987,N_7057,N_6348);
and U17988 (N_17988,N_7377,N_9732);
nand U17989 (N_17989,N_10439,N_6050);
xor U17990 (N_17990,N_6711,N_7269);
nor U17991 (N_17991,N_11094,N_10994);
nor U17992 (N_17992,N_10411,N_9935);
and U17993 (N_17993,N_11916,N_10403);
and U17994 (N_17994,N_10188,N_10142);
or U17995 (N_17995,N_9544,N_9726);
xor U17996 (N_17996,N_7206,N_10758);
or U17997 (N_17997,N_11754,N_9950);
nor U17998 (N_17998,N_10484,N_9211);
and U17999 (N_17999,N_7268,N_6540);
xnor U18000 (N_18000,N_13682,N_15673);
nand U18001 (N_18001,N_15497,N_14971);
nand U18002 (N_18002,N_14495,N_15553);
xnor U18003 (N_18003,N_12153,N_16163);
nand U18004 (N_18004,N_14638,N_13039);
and U18005 (N_18005,N_15079,N_12570);
or U18006 (N_18006,N_14582,N_12127);
nor U18007 (N_18007,N_16189,N_15718);
or U18008 (N_18008,N_12168,N_13681);
or U18009 (N_18009,N_13148,N_14944);
xnor U18010 (N_18010,N_12250,N_15552);
and U18011 (N_18011,N_17138,N_17344);
nor U18012 (N_18012,N_15484,N_12539);
xnor U18013 (N_18013,N_15751,N_13128);
nor U18014 (N_18014,N_16115,N_17008);
or U18015 (N_18015,N_12457,N_12656);
nor U18016 (N_18016,N_13136,N_15769);
nand U18017 (N_18017,N_14506,N_12590);
or U18018 (N_18018,N_16429,N_17931);
and U18019 (N_18019,N_14479,N_13757);
or U18020 (N_18020,N_13209,N_13886);
nand U18021 (N_18021,N_13871,N_15899);
xor U18022 (N_18022,N_14698,N_17258);
and U18023 (N_18023,N_15185,N_16003);
nand U18024 (N_18024,N_16892,N_12309);
nor U18025 (N_18025,N_13697,N_14326);
xor U18026 (N_18026,N_15796,N_15419);
xnor U18027 (N_18027,N_14822,N_13350);
or U18028 (N_18028,N_14268,N_17462);
nor U18029 (N_18029,N_14279,N_17019);
nor U18030 (N_18030,N_16310,N_12736);
or U18031 (N_18031,N_14264,N_14351);
or U18032 (N_18032,N_15108,N_17403);
and U18033 (N_18033,N_12100,N_13093);
nand U18034 (N_18034,N_13425,N_12244);
and U18035 (N_18035,N_15889,N_17648);
or U18036 (N_18036,N_13958,N_16778);
xor U18037 (N_18037,N_17080,N_15914);
xnor U18038 (N_18038,N_12596,N_14207);
xnor U18039 (N_18039,N_16801,N_13349);
or U18040 (N_18040,N_17074,N_13608);
and U18041 (N_18041,N_16533,N_15775);
and U18042 (N_18042,N_14448,N_16316);
nand U18043 (N_18043,N_12444,N_16386);
nor U18044 (N_18044,N_14078,N_13949);
nand U18045 (N_18045,N_12635,N_12468);
and U18046 (N_18046,N_17277,N_16265);
and U18047 (N_18047,N_16886,N_13790);
xor U18048 (N_18048,N_14601,N_13574);
xnor U18049 (N_18049,N_14300,N_16981);
nand U18050 (N_18050,N_16363,N_17967);
and U18051 (N_18051,N_16758,N_17123);
nor U18052 (N_18052,N_16447,N_16198);
or U18053 (N_18053,N_16146,N_13753);
xor U18054 (N_18054,N_16024,N_14664);
and U18055 (N_18055,N_17830,N_15839);
or U18056 (N_18056,N_15305,N_13974);
nor U18057 (N_18057,N_14146,N_13527);
or U18058 (N_18058,N_15440,N_12698);
and U18059 (N_18059,N_14567,N_17231);
xor U18060 (N_18060,N_17249,N_12239);
nor U18061 (N_18061,N_16486,N_13760);
nand U18062 (N_18062,N_12860,N_17785);
nand U18063 (N_18063,N_12864,N_15020);
and U18064 (N_18064,N_13851,N_12430);
and U18065 (N_18065,N_17101,N_16991);
xor U18066 (N_18066,N_12284,N_14017);
and U18067 (N_18067,N_15413,N_17978);
nand U18068 (N_18068,N_15625,N_16543);
xnor U18069 (N_18069,N_14870,N_16119);
xnor U18070 (N_18070,N_17065,N_13873);
xor U18071 (N_18071,N_16499,N_13567);
xnor U18072 (N_18072,N_15518,N_16093);
or U18073 (N_18073,N_12243,N_17486);
nand U18074 (N_18074,N_17173,N_16131);
xor U18075 (N_18075,N_15427,N_12876);
nand U18076 (N_18076,N_13249,N_15970);
and U18077 (N_18077,N_12392,N_15945);
nor U18078 (N_18078,N_15551,N_16688);
xor U18079 (N_18079,N_15697,N_12928);
or U18080 (N_18080,N_15711,N_17930);
xnor U18081 (N_18081,N_12565,N_17007);
and U18082 (N_18082,N_16677,N_14225);
nand U18083 (N_18083,N_15670,N_12425);
nor U18084 (N_18084,N_14115,N_15418);
and U18085 (N_18085,N_17568,N_15479);
and U18086 (N_18086,N_15187,N_17307);
or U18087 (N_18087,N_15549,N_15281);
nor U18088 (N_18088,N_15928,N_15234);
and U18089 (N_18089,N_17201,N_17832);
xor U18090 (N_18090,N_12897,N_13661);
nor U18091 (N_18091,N_16770,N_15131);
nor U18092 (N_18092,N_16451,N_14218);
xnor U18093 (N_18093,N_13602,N_16645);
or U18094 (N_18094,N_12220,N_14431);
and U18095 (N_18095,N_14366,N_14329);
nor U18096 (N_18096,N_15783,N_13151);
xor U18097 (N_18097,N_15346,N_12434);
xor U18098 (N_18098,N_14124,N_15203);
or U18099 (N_18099,N_16775,N_14782);
nor U18100 (N_18100,N_14517,N_13898);
nor U18101 (N_18101,N_17886,N_15431);
and U18102 (N_18102,N_13784,N_15962);
nand U18103 (N_18103,N_15617,N_17961);
nor U18104 (N_18104,N_13052,N_13104);
or U18105 (N_18105,N_14034,N_16640);
and U18106 (N_18106,N_13576,N_12453);
xnor U18107 (N_18107,N_16089,N_17475);
or U18108 (N_18108,N_17266,N_14070);
nand U18109 (N_18109,N_15033,N_15791);
or U18110 (N_18110,N_16592,N_14900);
nor U18111 (N_18111,N_17975,N_16492);
and U18112 (N_18112,N_13809,N_14252);
nor U18113 (N_18113,N_13872,N_13194);
xor U18114 (N_18114,N_14661,N_17021);
nor U18115 (N_18115,N_17511,N_13934);
and U18116 (N_18116,N_12569,N_15099);
or U18117 (N_18117,N_16963,N_13340);
nand U18118 (N_18118,N_16211,N_14357);
nand U18119 (N_18119,N_14219,N_16293);
nand U18120 (N_18120,N_17781,N_17126);
and U18121 (N_18121,N_15919,N_12251);
or U18122 (N_18122,N_12528,N_15955);
xnor U18123 (N_18123,N_15516,N_15843);
nand U18124 (N_18124,N_13969,N_16297);
xnor U18125 (N_18125,N_13017,N_17195);
nand U18126 (N_18126,N_15630,N_14147);
xnor U18127 (N_18127,N_17479,N_16700);
and U18128 (N_18128,N_13687,N_13018);
or U18129 (N_18129,N_16958,N_14690);
or U18130 (N_18130,N_15444,N_13843);
and U18131 (N_18131,N_15864,N_16736);
and U18132 (N_18132,N_17350,N_17049);
nor U18133 (N_18133,N_14702,N_15429);
nand U18134 (N_18134,N_13769,N_14245);
or U18135 (N_18135,N_12823,N_14989);
or U18136 (N_18136,N_16716,N_14918);
nor U18137 (N_18137,N_13620,N_15644);
or U18138 (N_18138,N_16041,N_17399);
and U18139 (N_18139,N_14312,N_17160);
xor U18140 (N_18140,N_16590,N_13038);
nor U18141 (N_18141,N_14596,N_16097);
nor U18142 (N_18142,N_14165,N_16609);
or U18143 (N_18143,N_13099,N_12353);
nand U18144 (N_18144,N_14552,N_16784);
and U18145 (N_18145,N_16002,N_17554);
nand U18146 (N_18146,N_15600,N_12573);
and U18147 (N_18147,N_17859,N_12126);
nor U18148 (N_18148,N_15909,N_17583);
nor U18149 (N_18149,N_13145,N_15814);
nor U18150 (N_18150,N_17463,N_17761);
nand U18151 (N_18151,N_14507,N_15476);
nor U18152 (N_18152,N_17692,N_15938);
and U18153 (N_18153,N_15976,N_12316);
or U18154 (N_18154,N_17082,N_13801);
xnor U18155 (N_18155,N_16122,N_17457);
nand U18156 (N_18156,N_13797,N_13802);
nor U18157 (N_18157,N_17118,N_13766);
xor U18158 (N_18158,N_17875,N_17435);
and U18159 (N_18159,N_13699,N_15638);
and U18160 (N_18160,N_16144,N_13316);
xnor U18161 (N_18161,N_17612,N_13599);
xor U18162 (N_18162,N_14851,N_13050);
nor U18163 (N_18163,N_14282,N_13207);
xor U18164 (N_18164,N_16523,N_12853);
nand U18165 (N_18165,N_12489,N_17112);
nand U18166 (N_18166,N_17974,N_17393);
xor U18167 (N_18167,N_17768,N_14770);
nor U18168 (N_18168,N_16353,N_12298);
nand U18169 (N_18169,N_14995,N_13261);
and U18170 (N_18170,N_15228,N_12686);
xor U18171 (N_18171,N_16245,N_12101);
nand U18172 (N_18172,N_17728,N_12831);
nor U18173 (N_18173,N_14413,N_16561);
and U18174 (N_18174,N_16601,N_14149);
or U18175 (N_18175,N_14217,N_17742);
and U18176 (N_18176,N_14981,N_16460);
nor U18177 (N_18177,N_17073,N_16707);
nand U18178 (N_18178,N_15038,N_14882);
nand U18179 (N_18179,N_12713,N_15143);
xor U18180 (N_18180,N_13074,N_14508);
nand U18181 (N_18181,N_14546,N_17690);
or U18182 (N_18182,N_13723,N_13816);
and U18183 (N_18183,N_16009,N_14543);
and U18184 (N_18184,N_15870,N_14815);
and U18185 (N_18185,N_15403,N_12916);
xor U18186 (N_18186,N_15577,N_13158);
xnor U18187 (N_18187,N_17217,N_14211);
nor U18188 (N_18188,N_12113,N_16955);
nand U18189 (N_18189,N_16237,N_12939);
nor U18190 (N_18190,N_17681,N_12829);
xor U18191 (N_18191,N_14297,N_17229);
nor U18192 (N_18192,N_13643,N_12557);
or U18193 (N_18193,N_17041,N_13722);
or U18194 (N_18194,N_15815,N_15822);
xnor U18195 (N_18195,N_15068,N_15107);
and U18196 (N_18196,N_15612,N_16988);
or U18197 (N_18197,N_17897,N_16067);
nand U18198 (N_18198,N_12287,N_12415);
or U18199 (N_18199,N_12895,N_12610);
nand U18200 (N_18200,N_12114,N_17800);
nor U18201 (N_18201,N_14048,N_17158);
nor U18202 (N_18202,N_12484,N_13323);
nand U18203 (N_18203,N_12073,N_14487);
nor U18204 (N_18204,N_17620,N_17539);
and U18205 (N_18205,N_12822,N_15994);
xnor U18206 (N_18206,N_14094,N_15169);
or U18207 (N_18207,N_16974,N_15681);
or U18208 (N_18208,N_13069,N_14383);
and U18209 (N_18209,N_12470,N_13839);
nor U18210 (N_18210,N_17447,N_14496);
xor U18211 (N_18211,N_15258,N_16441);
and U18212 (N_18212,N_17952,N_15098);
nand U18213 (N_18213,N_17853,N_13830);
xor U18214 (N_18214,N_17907,N_16647);
nor U18215 (N_18215,N_14714,N_13241);
xnor U18216 (N_18216,N_15027,N_16333);
nor U18217 (N_18217,N_12761,N_12027);
or U18218 (N_18218,N_13095,N_15776);
xnor U18219 (N_18219,N_14704,N_17889);
nand U18220 (N_18220,N_12029,N_12364);
or U18221 (N_18221,N_12628,N_17689);
and U18222 (N_18222,N_14750,N_17717);
xor U18223 (N_18223,N_15196,N_14370);
or U18224 (N_18224,N_15682,N_17547);
and U18225 (N_18225,N_16220,N_14043);
or U18226 (N_18226,N_16346,N_14462);
nor U18227 (N_18227,N_15318,N_16701);
nand U18228 (N_18228,N_14414,N_17998);
or U18229 (N_18229,N_14864,N_15425);
or U18230 (N_18230,N_14982,N_13692);
xor U18231 (N_18231,N_14172,N_16004);
and U18232 (N_18232,N_12799,N_13749);
or U18233 (N_18233,N_14557,N_15420);
nand U18234 (N_18234,N_14404,N_14355);
or U18235 (N_18235,N_13733,N_12174);
or U18236 (N_18236,N_13313,N_15794);
xor U18237 (N_18237,N_16855,N_17288);
or U18238 (N_18238,N_15716,N_16303);
nand U18239 (N_18239,N_13583,N_17528);
and U18240 (N_18240,N_12394,N_13512);
nand U18241 (N_18241,N_15595,N_16474);
and U18242 (N_18242,N_15650,N_17427);
xnor U18243 (N_18243,N_12796,N_13272);
nor U18244 (N_18244,N_13412,N_15987);
nand U18245 (N_18245,N_16919,N_13968);
xor U18246 (N_18246,N_12276,N_16796);
nand U18247 (N_18247,N_12901,N_16743);
nand U18248 (N_18248,N_15969,N_12151);
xor U18249 (N_18249,N_13854,N_12963);
and U18250 (N_18250,N_17760,N_14293);
xnor U18251 (N_18251,N_14899,N_16742);
xor U18252 (N_18252,N_12943,N_13308);
nand U18253 (N_18253,N_15224,N_16712);
nand U18254 (N_18254,N_17825,N_12607);
and U18255 (N_18255,N_16535,N_16473);
or U18256 (N_18256,N_12968,N_17841);
and U18257 (N_18257,N_14333,N_16488);
xnor U18258 (N_18258,N_15330,N_13948);
nand U18259 (N_18259,N_15739,N_14806);
and U18260 (N_18260,N_16532,N_13730);
and U18261 (N_18261,N_13426,N_12833);
and U18262 (N_18262,N_13546,N_13086);
xor U18263 (N_18263,N_15255,N_12070);
xor U18264 (N_18264,N_14535,N_12365);
xnor U18265 (N_18265,N_12715,N_13929);
or U18266 (N_18266,N_16449,N_15686);
nor U18267 (N_18267,N_17042,N_13744);
or U18268 (N_18268,N_15985,N_14186);
nor U18269 (N_18269,N_12280,N_12320);
xnor U18270 (N_18270,N_17521,N_13270);
or U18271 (N_18271,N_13023,N_16336);
xor U18272 (N_18272,N_17679,N_16824);
or U18273 (N_18273,N_13765,N_16766);
nand U18274 (N_18274,N_15058,N_14990);
nand U18275 (N_18275,N_17854,N_15423);
or U18276 (N_18276,N_12265,N_13078);
and U18277 (N_18277,N_16145,N_16457);
or U18278 (N_18278,N_12514,N_13568);
xor U18279 (N_18279,N_13642,N_15659);
or U18280 (N_18280,N_15911,N_12708);
and U18281 (N_18281,N_13947,N_12381);
xnor U18282 (N_18282,N_15371,N_17279);
nor U18283 (N_18283,N_14687,N_12993);
xor U18284 (N_18284,N_15599,N_17386);
and U18285 (N_18285,N_14263,N_16867);
xor U18286 (N_18286,N_16270,N_14859);
xnor U18287 (N_18287,N_15387,N_12477);
xnor U18288 (N_18288,N_17204,N_17437);
xnor U18289 (N_18289,N_12268,N_17418);
xor U18290 (N_18290,N_14608,N_13778);
and U18291 (N_18291,N_17341,N_13072);
or U18292 (N_18292,N_13719,N_14046);
xor U18293 (N_18293,N_13075,N_15626);
or U18294 (N_18294,N_17358,N_13237);
nor U18295 (N_18295,N_12196,N_14522);
and U18296 (N_18296,N_17563,N_15462);
xnor U18297 (N_18297,N_12001,N_14424);
nand U18298 (N_18298,N_13509,N_13247);
or U18299 (N_18299,N_12850,N_15661);
nor U18300 (N_18300,N_14948,N_17223);
and U18301 (N_18301,N_15740,N_13795);
xnor U18302 (N_18302,N_16977,N_13991);
xor U18303 (N_18303,N_12751,N_12877);
nand U18304 (N_18304,N_16608,N_12915);
and U18305 (N_18305,N_14038,N_14620);
or U18306 (N_18306,N_12687,N_12111);
xnor U18307 (N_18307,N_15583,N_14532);
xor U18308 (N_18308,N_14937,N_15102);
xnor U18309 (N_18309,N_16513,N_15047);
xnor U18310 (N_18310,N_16327,N_17735);
and U18311 (N_18311,N_16788,N_13331);
and U18312 (N_18312,N_12124,N_13764);
xnor U18313 (N_18313,N_12272,N_15023);
nor U18314 (N_18314,N_17412,N_14785);
or U18315 (N_18315,N_14723,N_14602);
or U18316 (N_18316,N_12206,N_15593);
nor U18317 (N_18317,N_16182,N_13963);
nand U18318 (N_18318,N_17855,N_17608);
nand U18319 (N_18319,N_13665,N_17860);
and U18320 (N_18320,N_13876,N_13793);
nor U18321 (N_18321,N_14660,N_16498);
nand U18322 (N_18322,N_12116,N_16774);
nor U18323 (N_18323,N_16510,N_15627);
nand U18324 (N_18324,N_13694,N_15326);
nor U18325 (N_18325,N_14468,N_12966);
nor U18326 (N_18326,N_17794,N_16943);
xnor U18327 (N_18327,N_13625,N_13381);
nor U18328 (N_18328,N_12150,N_17647);
or U18329 (N_18329,N_17848,N_12544);
nand U18330 (N_18330,N_17845,N_12676);
nand U18331 (N_18331,N_17782,N_15035);
and U18332 (N_18332,N_15441,N_14276);
and U18333 (N_18333,N_16816,N_16044);
nand U18334 (N_18334,N_12112,N_13214);
nor U18335 (N_18335,N_13456,N_13782);
nor U18336 (N_18336,N_12002,N_14190);
and U18337 (N_18337,N_12741,N_14184);
nand U18338 (N_18338,N_15110,N_13179);
and U18339 (N_18339,N_13912,N_17614);
nand U18340 (N_18340,N_17045,N_17169);
or U18341 (N_18341,N_15542,N_15194);
nand U18342 (N_18342,N_12862,N_13515);
xor U18343 (N_18343,N_13796,N_16483);
or U18344 (N_18344,N_15894,N_15189);
nand U18345 (N_18345,N_17092,N_17194);
nor U18346 (N_18346,N_13337,N_16411);
nor U18347 (N_18347,N_15589,N_16560);
and U18348 (N_18348,N_14463,N_15188);
nor U18349 (N_18349,N_12214,N_17773);
or U18350 (N_18350,N_17550,N_13475);
or U18351 (N_18351,N_15931,N_13591);
nand U18352 (N_18352,N_16016,N_15292);
and U18353 (N_18353,N_15550,N_16582);
or U18354 (N_18354,N_17410,N_13362);
xor U18355 (N_18355,N_17044,N_17895);
xor U18356 (N_18356,N_17110,N_12630);
xor U18357 (N_18357,N_15932,N_12804);
or U18358 (N_18358,N_17569,N_13980);
nand U18359 (N_18359,N_17164,N_16376);
xor U18360 (N_18360,N_12140,N_12617);
nor U18361 (N_18361,N_15746,N_12671);
and U18362 (N_18362,N_16407,N_16833);
nor U18363 (N_18363,N_12807,N_16908);
nor U18364 (N_18364,N_15057,N_16020);
nand U18365 (N_18365,N_14030,N_17365);
or U18366 (N_18366,N_15037,N_15119);
or U18367 (N_18367,N_13021,N_17771);
xor U18368 (N_18368,N_12899,N_12917);
and U18369 (N_18369,N_15588,N_16347);
nor U18370 (N_18370,N_17879,N_14974);
or U18371 (N_18371,N_12692,N_14340);
nand U18372 (N_18372,N_14833,N_12185);
or U18373 (N_18373,N_15773,N_13924);
or U18374 (N_18374,N_13965,N_12060);
nor U18375 (N_18375,N_17091,N_12670);
or U18376 (N_18376,N_17817,N_17216);
xor U18377 (N_18377,N_15111,N_13484);
xor U18378 (N_18378,N_13492,N_15685);
nand U18379 (N_18379,N_16884,N_16406);
and U18380 (N_18380,N_12718,N_13696);
nand U18381 (N_18381,N_15745,N_12324);
or U18382 (N_18382,N_15755,N_15443);
nand U18383 (N_18383,N_16162,N_17718);
and U18384 (N_18384,N_13227,N_17373);
or U18385 (N_18385,N_16719,N_15301);
nand U18386 (N_18386,N_13079,N_17107);
xor U18387 (N_18387,N_17413,N_15486);
nor U18388 (N_18388,N_17762,N_12691);
nand U18389 (N_18389,N_16841,N_12305);
and U18390 (N_18390,N_13926,N_17150);
xnor U18391 (N_18391,N_16373,N_13286);
nand U18392 (N_18392,N_17987,N_16383);
and U18393 (N_18393,N_17752,N_12158);
nor U18394 (N_18394,N_14636,N_14604);
or U18395 (N_18395,N_12537,N_16665);
or U18396 (N_18396,N_17208,N_13800);
or U18397 (N_18397,N_16082,N_15930);
nor U18398 (N_18398,N_17565,N_14528);
nor U18399 (N_18399,N_15042,N_17751);
nand U18400 (N_18400,N_12660,N_13650);
nor U18401 (N_18401,N_13728,N_14461);
and U18402 (N_18402,N_12615,N_16466);
or U18403 (N_18403,N_15095,N_13312);
xor U18404 (N_18404,N_13742,N_17347);
or U18405 (N_18405,N_15948,N_14629);
nand U18406 (N_18406,N_13850,N_16141);
and U18407 (N_18407,N_12984,N_13666);
nand U18408 (N_18408,N_13216,N_12995);
nor U18409 (N_18409,N_15777,N_17495);
xnor U18410 (N_18410,N_13283,N_13551);
nand U18411 (N_18411,N_15980,N_16231);
xnor U18412 (N_18412,N_15083,N_14827);
nor U18413 (N_18413,N_14547,N_13131);
nand U18414 (N_18414,N_14967,N_16858);
and U18415 (N_18415,N_13265,N_16199);
and U18416 (N_18416,N_16204,N_17221);
or U18417 (N_18417,N_17453,N_16922);
or U18418 (N_18418,N_15322,N_17601);
and U18419 (N_18419,N_17948,N_17954);
and U18420 (N_18420,N_12212,N_16390);
xnor U18421 (N_18421,N_17245,N_16127);
and U18422 (N_18422,N_13825,N_13314);
xor U18423 (N_18423,N_12896,N_13009);
xnor U18424 (N_18424,N_12293,N_14823);
and U18425 (N_18425,N_15536,N_12962);
and U18426 (N_18426,N_15295,N_15736);
nor U18427 (N_18427,N_14761,N_13906);
nand U18428 (N_18428,N_14783,N_14485);
or U18429 (N_18429,N_12375,N_17929);
xnor U18430 (N_18430,N_17693,N_12322);
nand U18431 (N_18431,N_17669,N_13834);
and U18432 (N_18432,N_15276,N_12157);
nor U18433 (N_18433,N_17787,N_15863);
nand U18434 (N_18434,N_17582,N_16495);
nor U18435 (N_18435,N_15106,N_12357);
xor U18436 (N_18436,N_17891,N_14458);
and U18437 (N_18437,N_15400,N_14656);
and U18438 (N_18438,N_13068,N_14984);
nor U18439 (N_18439,N_14028,N_16720);
nand U18440 (N_18440,N_14369,N_16754);
xnor U18441 (N_18441,N_14179,N_12504);
xnor U18442 (N_18442,N_16143,N_15679);
or U18443 (N_18443,N_14405,N_13669);
or U18444 (N_18444,N_17856,N_16682);
nand U18445 (N_18445,N_12495,N_16021);
xnor U18446 (N_18446,N_12765,N_16875);
xnor U18447 (N_18447,N_15758,N_14708);
or U18448 (N_18448,N_16140,N_16167);
and U18449 (N_18449,N_15983,N_14756);
xnor U18450 (N_18450,N_16197,N_15528);
nor U18451 (N_18451,N_14983,N_14811);
nand U18452 (N_18452,N_17087,N_12410);
nand U18453 (N_18453,N_17602,N_17309);
xor U18454 (N_18454,N_15494,N_14755);
or U18455 (N_18455,N_17411,N_16803);
and U18456 (N_18456,N_13732,N_15202);
nand U18457 (N_18457,N_14232,N_14086);
nor U18458 (N_18458,N_15103,N_12530);
nor U18459 (N_18459,N_12256,N_13914);
and U18460 (N_18460,N_14001,N_14313);
and U18461 (N_18461,N_15272,N_12122);
nor U18462 (N_18462,N_13799,N_15459);
or U18463 (N_18463,N_13154,N_16377);
nor U18464 (N_18464,N_15967,N_17115);
and U18465 (N_18465,N_13907,N_16087);
nand U18466 (N_18466,N_12082,N_15250);
nor U18467 (N_18467,N_15376,N_17869);
xnor U18468 (N_18468,N_17814,N_13613);
and U18469 (N_18469,N_12420,N_17490);
or U18470 (N_18470,N_14876,N_12198);
xnor U18471 (N_18471,N_12568,N_16201);
or U18472 (N_18472,N_15069,N_15927);
xnor U18473 (N_18473,N_14465,N_14084);
xnor U18474 (N_18474,N_13667,N_16520);
nand U18475 (N_18475,N_12437,N_15534);
xor U18476 (N_18476,N_16030,N_13186);
xor U18477 (N_18477,N_14634,N_13204);
nand U18478 (N_18478,N_17757,N_17624);
nor U18479 (N_18479,N_13459,N_12689);
or U18480 (N_18480,N_12732,N_17094);
or U18481 (N_18481,N_12325,N_16555);
or U18482 (N_18482,N_15508,N_12460);
xor U18483 (N_18483,N_15460,N_17989);
or U18484 (N_18484,N_13427,N_12471);
nor U18485 (N_18485,N_17604,N_17270);
or U18486 (N_18486,N_17591,N_17077);
or U18487 (N_18487,N_14008,N_17459);
and U18488 (N_18488,N_12839,N_12575);
nand U18489 (N_18489,N_12851,N_17441);
and U18490 (N_18490,N_15873,N_15956);
nand U18491 (N_18491,N_12428,N_17900);
xor U18492 (N_18492,N_12631,N_16863);
nand U18493 (N_18493,N_16038,N_15537);
xnor U18494 (N_18494,N_12584,N_16502);
or U18495 (N_18495,N_17178,N_16638);
and U18496 (N_18496,N_13045,N_14749);
and U18497 (N_18497,N_13975,N_15744);
or U18498 (N_18498,N_14097,N_12503);
nor U18499 (N_18499,N_17755,N_14940);
nand U18500 (N_18500,N_15025,N_12932);
nand U18501 (N_18501,N_13223,N_17766);
xnor U18502 (N_18502,N_13960,N_16945);
nand U18503 (N_18503,N_13915,N_16990);
xnor U18504 (N_18504,N_13371,N_14652);
and U18505 (N_18505,N_17982,N_17375);
xnor U18506 (N_18506,N_13556,N_16056);
nand U18507 (N_18507,N_12781,N_12066);
nor U18508 (N_18508,N_16033,N_15026);
nor U18509 (N_18509,N_17285,N_15286);
xor U18510 (N_18510,N_13918,N_14069);
and U18511 (N_18511,N_14807,N_13443);
and U18512 (N_18512,N_13363,N_13610);
xnor U18513 (N_18513,N_17202,N_15003);
and U18514 (N_18514,N_12216,N_14996);
or U18515 (N_18515,N_13082,N_15858);
nand U18516 (N_18516,N_14534,N_12764);
nand U18517 (N_18517,N_17981,N_12663);
nor U18518 (N_18518,N_13811,N_17536);
and U18519 (N_18519,N_17053,N_17289);
nor U18520 (N_18520,N_13675,N_14295);
nand U18521 (N_18521,N_15097,N_14878);
xor U18522 (N_18522,N_16463,N_12934);
nand U18523 (N_18523,N_17426,N_13863);
nand U18524 (N_18524,N_17449,N_15653);
nand U18525 (N_18525,N_13382,N_15748);
xnor U18526 (N_18526,N_13521,N_14997);
nor U18527 (N_18527,N_15906,N_14685);
or U18528 (N_18528,N_14377,N_15901);
or U18529 (N_18529,N_13455,N_15687);
and U18530 (N_18530,N_12775,N_17708);
nand U18531 (N_18531,N_14352,N_14515);
or U18532 (N_18532,N_12595,N_17744);
nor U18533 (N_18533,N_16574,N_13702);
nor U18534 (N_18534,N_12821,N_15018);
nor U18535 (N_18535,N_17917,N_14800);
nand U18536 (N_18536,N_14427,N_12292);
and U18537 (N_18537,N_12929,N_12762);
and U18538 (N_18538,N_15446,N_13133);
xor U18539 (N_18539,N_13940,N_12819);
nand U18540 (N_18540,N_16046,N_13259);
nor U18541 (N_18541,N_14025,N_13152);
and U18542 (N_18542,N_17084,N_14382);
and U18543 (N_18543,N_17192,N_15565);
or U18544 (N_18544,N_17772,N_17137);
or U18545 (N_18545,N_15408,N_15380);
nand U18546 (N_18546,N_12709,N_14646);
nor U18547 (N_18547,N_16355,N_12258);
and U18548 (N_18548,N_12559,N_13306);
and U18549 (N_18549,N_16010,N_13496);
or U18550 (N_18550,N_16280,N_15317);
or U18551 (N_18551,N_12363,N_13225);
nand U18552 (N_18552,N_14315,N_15892);
or U18553 (N_18553,N_15261,N_13434);
xnor U18554 (N_18554,N_17968,N_12389);
and U18555 (N_18555,N_14445,N_16802);
or U18556 (N_18556,N_16099,N_15929);
nor U18557 (N_18557,N_13932,N_14917);
nand U18558 (N_18558,N_14849,N_14055);
nor U18559 (N_18559,N_16356,N_13451);
or U18560 (N_18560,N_17335,N_13184);
nand U18561 (N_18561,N_14693,N_13277);
or U18562 (N_18562,N_14011,N_13255);
nand U18563 (N_18563,N_13366,N_13070);
nand U18564 (N_18564,N_13046,N_16173);
xnor U18565 (N_18565,N_12106,N_16966);
xnor U18566 (N_18566,N_17481,N_12578);
or U18567 (N_18567,N_12767,N_12529);
nor U18568 (N_18568,N_12228,N_15029);
nor U18569 (N_18569,N_12626,N_13325);
xor U18570 (N_18570,N_14188,N_15364);
nor U18571 (N_18571,N_16586,N_12380);
or U18572 (N_18572,N_16320,N_15857);
nor U18573 (N_18573,N_16838,N_16018);
nand U18574 (N_18574,N_15604,N_12221);
or U18575 (N_18575,N_17622,N_16181);
xnor U18576 (N_18576,N_13715,N_13541);
nor U18577 (N_18577,N_14240,N_13806);
nand U18578 (N_18578,N_13821,N_17362);
or U18579 (N_18579,N_16900,N_15200);
nand U18580 (N_18580,N_15061,N_16480);
nand U18581 (N_18581,N_13105,N_16428);
and U18582 (N_18582,N_13619,N_14667);
nand U18583 (N_18583,N_15172,N_14116);
and U18584 (N_18584,N_15040,N_13930);
nor U18585 (N_18585,N_15067,N_12427);
and U18586 (N_18586,N_13467,N_17054);
and U18587 (N_18587,N_12562,N_14922);
or U18588 (N_18588,N_14033,N_12040);
xnor U18589 (N_18589,N_15012,N_12035);
xor U18590 (N_18590,N_16779,N_13494);
nor U18591 (N_18591,N_14406,N_16302);
nor U18592 (N_18592,N_14887,N_17581);
and U18593 (N_18593,N_13649,N_14901);
nor U18594 (N_18594,N_16408,N_17318);
nor U18595 (N_18595,N_13976,N_13112);
nand U18596 (N_18596,N_13822,N_15306);
nor U18597 (N_18597,N_15296,N_12857);
or U18598 (N_18598,N_16092,N_17348);
or U18599 (N_18599,N_14277,N_16274);
nand U18600 (N_18600,N_16953,N_17576);
or U18601 (N_18601,N_15559,N_12875);
and U18602 (N_18602,N_16216,N_14666);
nor U18603 (N_18603,N_13919,N_16137);
xor U18604 (N_18604,N_16672,N_17100);
nand U18605 (N_18605,N_14450,N_16098);
and U18606 (N_18606,N_12612,N_15205);
nor U18607 (N_18607,N_12348,N_14139);
or U18608 (N_18608,N_13327,N_16073);
nand U18609 (N_18609,N_12662,N_13770);
nor U18610 (N_18610,N_14627,N_17764);
nand U18611 (N_18611,N_16959,N_12036);
and U18612 (N_18612,N_13543,N_17846);
or U18613 (N_18613,N_14612,N_13985);
xor U18614 (N_18614,N_16080,N_17531);
nand U18615 (N_18615,N_12231,N_12217);
nand U18616 (N_18616,N_14679,N_17136);
and U18617 (N_18617,N_15946,N_17714);
and U18618 (N_18618,N_15451,N_13904);
nor U18619 (N_18619,N_13413,N_13200);
xnor U18620 (N_18620,N_17505,N_12605);
or U18621 (N_18621,N_14503,N_15044);
nor U18622 (N_18622,N_15424,N_13664);
nor U18623 (N_18623,N_12177,N_15381);
or U18624 (N_18624,N_13993,N_12386);
nor U18625 (N_18625,N_16865,N_13920);
nand U18626 (N_18626,N_16291,N_14863);
xnor U18627 (N_18627,N_17600,N_16589);
xnor U18628 (N_18628,N_13368,N_17154);
xor U18629 (N_18629,N_16685,N_15327);
nor U18630 (N_18630,N_13626,N_15504);
xor U18631 (N_18631,N_12694,N_13091);
nor U18632 (N_18632,N_12515,N_14428);
and U18633 (N_18633,N_14578,N_14100);
or U18634 (N_18634,N_15651,N_13833);
nor U18635 (N_18635,N_12401,N_16104);
and U18636 (N_18636,N_17246,N_12043);
and U18637 (N_18637,N_16583,N_16168);
and U18638 (N_18638,N_12508,N_12015);
xnor U18639 (N_18639,N_13693,N_17088);
and U18640 (N_18640,N_15757,N_12519);
or U18641 (N_18641,N_15760,N_13003);
nor U18642 (N_18642,N_15471,N_12200);
or U18643 (N_18643,N_15865,N_15692);
and U18644 (N_18644,N_15880,N_12638);
or U18645 (N_18645,N_16597,N_16554);
nand U18646 (N_18646,N_12990,N_13376);
xnor U18647 (N_18647,N_17488,N_17310);
or U18648 (N_18648,N_15806,N_13606);
and U18649 (N_18649,N_17610,N_15860);
nor U18650 (N_18650,N_15869,N_15329);
nor U18651 (N_18651,N_17725,N_13013);
nand U18652 (N_18652,N_17852,N_15468);
nand U18653 (N_18653,N_13239,N_17237);
or U18654 (N_18654,N_16744,N_15960);
nor U18655 (N_18655,N_12951,N_12290);
and U18656 (N_18656,N_17176,N_13804);
or U18657 (N_18657,N_16613,N_14751);
nor U18658 (N_18658,N_13561,N_16230);
nand U18659 (N_18659,N_16292,N_15084);
and U18660 (N_18660,N_14549,N_16595);
and U18661 (N_18661,N_12024,N_13335);
or U18662 (N_18662,N_17440,N_17432);
nor U18663 (N_18663,N_17469,N_17370);
xor U18664 (N_18664,N_15359,N_12756);
nor U18665 (N_18665,N_16911,N_12237);
or U18666 (N_18666,N_14840,N_13288);
nor U18667 (N_18667,N_12026,N_15293);
and U18668 (N_18668,N_14059,N_15952);
nor U18669 (N_18669,N_17619,N_14183);
nor U18670 (N_18670,N_12296,N_13100);
nor U18671 (N_18671,N_15936,N_17361);
nor U18672 (N_18672,N_14928,N_12855);
or U18673 (N_18673,N_12306,N_12782);
or U18674 (N_18674,N_12843,N_14935);
and U18675 (N_18675,N_13309,N_17177);
and U18676 (N_18676,N_12922,N_15134);
nand U18677 (N_18677,N_12885,N_12142);
and U18678 (N_18678,N_15470,N_12563);
and U18679 (N_18679,N_15513,N_14654);
xor U18680 (N_18680,N_14469,N_14668);
and U18681 (N_18681,N_17522,N_13466);
nor U18682 (N_18682,N_15637,N_13373);
and U18683 (N_18683,N_12545,N_17039);
xnor U18684 (N_18684,N_15949,N_13526);
xor U18685 (N_18685,N_15629,N_13534);
or U18686 (N_18686,N_13653,N_16323);
or U18687 (N_18687,N_15940,N_14275);
nor U18688 (N_18688,N_16263,N_15309);
and U18689 (N_18689,N_12820,N_15498);
nor U18690 (N_18690,N_16813,N_13185);
nand U18691 (N_18691,N_16961,N_14700);
xnor U18692 (N_18692,N_12814,N_17997);
nand U18693 (N_18693,N_16248,N_14364);
xnor U18694 (N_18694,N_14308,N_13064);
nor U18695 (N_18695,N_14019,N_15951);
nand U18696 (N_18696,N_15544,N_16806);
nor U18697 (N_18697,N_16371,N_16951);
nor U18698 (N_18698,N_17503,N_16023);
nand U18699 (N_18699,N_16795,N_17443);
and U18700 (N_18700,N_16112,N_17663);
or U18701 (N_18701,N_16702,N_17838);
and U18702 (N_18702,N_12771,N_15005);
nor U18703 (N_18703,N_13637,N_17902);
and U18704 (N_18704,N_12128,N_14730);
and U18705 (N_18705,N_17259,N_17242);
nor U18706 (N_18706,N_17458,N_15587);
xor U18707 (N_18707,N_15677,N_12770);
nand U18708 (N_18708,N_15126,N_14266);
and U18709 (N_18709,N_16063,N_13129);
nor U18710 (N_18710,N_17777,N_12703);
or U18711 (N_18711,N_17227,N_16299);
or U18712 (N_18712,N_16036,N_15885);
xor U18713 (N_18713,N_15959,N_14888);
nor U18714 (N_18714,N_17661,N_12661);
xnor U18715 (N_18715,N_16026,N_14169);
and U18716 (N_18716,N_17269,N_12131);
or U18717 (N_18717,N_14689,N_12411);
nand U18718 (N_18718,N_12824,N_13959);
and U18719 (N_18719,N_17685,N_13585);
xnor U18720 (N_18720,N_12666,N_14570);
or U18721 (N_18721,N_17061,N_12706);
nand U18722 (N_18722,N_14455,N_13228);
and U18723 (N_18723,N_16129,N_15915);
nand U18724 (N_18724,N_16239,N_15132);
nor U18725 (N_18725,N_16587,N_17342);
and U18726 (N_18726,N_12918,N_14720);
or U18727 (N_18727,N_13529,N_13059);
and U18728 (N_18728,N_14026,N_12838);
or U18729 (N_18729,N_14360,N_14215);
nand U18730 (N_18730,N_17867,N_13213);
nor U18731 (N_18731,N_13103,N_14764);
nor U18732 (N_18732,N_13724,N_17184);
or U18733 (N_18733,N_14344,N_13780);
nand U18734 (N_18734,N_15941,N_15704);
or U18735 (N_18735,N_12688,N_12218);
and U18736 (N_18736,N_12743,N_14694);
nor U18737 (N_18737,N_13739,N_12006);
nand U18738 (N_18738,N_17791,N_12952);
nor U18739 (N_18739,N_16068,N_17686);
or U18740 (N_18740,N_16440,N_13848);
nand U18741 (N_18741,N_13967,N_14007);
nand U18742 (N_18742,N_15231,N_14719);
and U18743 (N_18743,N_14104,N_17416);
nand U18744 (N_18744,N_16591,N_12488);
xnor U18745 (N_18745,N_17325,N_12505);
and U18746 (N_18746,N_17696,N_16894);
or U18747 (N_18747,N_16123,N_12555);
and U18748 (N_18748,N_16281,N_12926);
nand U18749 (N_18749,N_12476,N_13005);
xnor U18750 (N_18750,N_14301,N_16968);
nor U18751 (N_18751,N_17476,N_15100);
xnor U18752 (N_18752,N_12500,N_16037);
nand U18753 (N_18753,N_12658,N_14272);
xnor U18754 (N_18754,N_14538,N_12009);
and U18755 (N_18755,N_16739,N_16435);
nor U18756 (N_18756,N_15094,N_15574);
xor U18757 (N_18757,N_14705,N_16653);
nor U18758 (N_18758,N_12310,N_12391);
or U18759 (N_18759,N_13379,N_17816);
or U18760 (N_18760,N_12780,N_12739);
and U18761 (N_18761,N_16848,N_12891);
nor U18762 (N_18762,N_13051,N_17527);
and U18763 (N_18763,N_17585,N_13645);
and U18764 (N_18764,N_15648,N_14681);
xor U18765 (N_18765,N_15953,N_12093);
nor U18766 (N_18766,N_13172,N_15086);
and U18767 (N_18767,N_14002,N_14904);
or U18768 (N_18768,N_15798,N_14611);
and U18769 (N_18769,N_13471,N_13336);
nor U18770 (N_18770,N_14391,N_15167);
nor U18771 (N_18771,N_17460,N_14903);
and U18772 (N_18772,N_14595,N_12271);
or U18773 (N_18773,N_16630,N_12913);
or U18774 (N_18774,N_15974,N_12248);
nand U18775 (N_18775,N_17134,N_12129);
or U18776 (N_18776,N_17944,N_15137);
nand U18777 (N_18777,N_13849,N_14564);
and U18778 (N_18778,N_15140,N_17894);
xnor U18779 (N_18779,N_15456,N_13096);
and U18780 (N_18780,N_15836,N_14839);
nand U18781 (N_18781,N_13221,N_14288);
nor U18782 (N_18782,N_14621,N_14205);
nand U18783 (N_18783,N_13215,N_17085);
and U18784 (N_18784,N_13973,N_13604);
nor U18785 (N_18785,N_16670,N_17759);
and U18786 (N_18786,N_14566,N_16161);
xnor U18787 (N_18787,N_17064,N_13955);
nor U18788 (N_18788,N_16529,N_17155);
or U18789 (N_18789,N_12974,N_12961);
nor U18790 (N_18790,N_17519,N_16102);
or U18791 (N_18791,N_16730,N_15605);
or U18792 (N_18792,N_14717,N_17618);
nand U18793 (N_18793,N_17850,N_17038);
nor U18794 (N_18794,N_13590,N_15664);
xor U18795 (N_18795,N_14828,N_17501);
xnor U18796 (N_18796,N_13041,N_15581);
xnor U18797 (N_18797,N_15555,N_16581);
xnor U18798 (N_18798,N_13440,N_13431);
xnor U18799 (N_18799,N_16714,N_14177);
nand U18800 (N_18800,N_16748,N_14743);
nor U18801 (N_18801,N_13882,N_13437);
xnor U18802 (N_18802,N_14056,N_16012);
nand U18803 (N_18803,N_17356,N_17908);
or U18804 (N_18804,N_12577,N_12524);
nand U18805 (N_18805,N_16360,N_15835);
nand U18806 (N_18806,N_17477,N_14881);
and U18807 (N_18807,N_15576,N_17297);
and U18808 (N_18808,N_17677,N_16866);
nand U18809 (N_18809,N_14453,N_16183);
xnor U18810 (N_18810,N_17298,N_14441);
nor U18811 (N_18811,N_15000,N_15789);
or U18812 (N_18812,N_16147,N_15358);
or U18813 (N_18813,N_12187,N_14735);
or U18814 (N_18814,N_12672,N_12076);
nor U18815 (N_18815,N_16124,N_13385);
or U18816 (N_18816,N_12145,N_13089);
nand U18817 (N_18817,N_14339,N_12016);
nor U18818 (N_18818,N_15934,N_15240);
and U18819 (N_18819,N_12283,N_16438);
nor U18820 (N_18820,N_14440,N_12640);
or U18821 (N_18821,N_17431,N_14797);
and U18822 (N_18822,N_17970,N_15719);
nor U18823 (N_18823,N_14052,N_17515);
xnor U18824 (N_18824,N_13773,N_16880);
nand U18825 (N_18825,N_17301,N_16234);
xor U18826 (N_18826,N_12600,N_14473);
nor U18827 (N_18827,N_13468,N_13372);
nand U18828 (N_18828,N_13077,N_14518);
or U18829 (N_18829,N_15421,N_14415);
nor U18830 (N_18830,N_14492,N_15325);
xnor U18831 (N_18831,N_14867,N_15561);
xor U18832 (N_18832,N_12955,N_12792);
or U18833 (N_18833,N_15332,N_15607);
nor U18834 (N_18834,N_15239,N_14227);
and U18835 (N_18835,N_12979,N_15168);
and U18836 (N_18836,N_17187,N_17367);
or U18837 (N_18837,N_14747,N_13598);
xnor U18838 (N_18838,N_13476,N_16564);
or U18839 (N_18839,N_17198,N_14083);
or U18840 (N_18840,N_16873,N_16433);
nand U18841 (N_18841,N_16361,N_17993);
nand U18842 (N_18842,N_15762,N_15208);
nor U18843 (N_18843,N_14247,N_15877);
and U18844 (N_18844,N_15699,N_16957);
xnor U18845 (N_18845,N_17542,N_15232);
nand U18846 (N_18846,N_16276,N_13163);
and U18847 (N_18847,N_15321,N_16315);
and U18848 (N_18848,N_14623,N_12785);
nor U18849 (N_18849,N_15756,N_16521);
xor U18850 (N_18850,N_17928,N_15384);
or U18851 (N_18851,N_15572,N_14163);
xnor U18852 (N_18852,N_12004,N_16541);
nor U18853 (N_18853,N_17887,N_16049);
or U18854 (N_18854,N_14790,N_12911);
and U18855 (N_18855,N_13002,N_13140);
xor U18856 (N_18856,N_15824,N_12475);
xnor U18857 (N_18857,N_12651,N_17197);
nor U18858 (N_18858,N_13705,N_15563);
and U18859 (N_18859,N_14187,N_12361);
nand U18860 (N_18860,N_16585,N_17387);
or U18861 (N_18861,N_13260,N_15527);
xnor U18862 (N_18862,N_14449,N_16525);
nor U18863 (N_18863,N_16108,N_13549);
nand U18864 (N_18864,N_12621,N_12034);
nor U18865 (N_18865,N_15817,N_16427);
xnor U18866 (N_18866,N_15201,N_12439);
and U18867 (N_18867,N_12472,N_16646);
nand U18868 (N_18868,N_16404,N_16296);
or U18869 (N_18869,N_12190,N_17036);
nor U18870 (N_18870,N_12802,N_14796);
and U18871 (N_18871,N_14718,N_15557);
nor U18872 (N_18872,N_13473,N_15900);
nor U18873 (N_18873,N_13305,N_14330);
and U18874 (N_18874,N_14640,N_12343);
and U18875 (N_18875,N_16626,N_15362);
nor U18876 (N_18876,N_13520,N_17424);
or U18877 (N_18877,N_14140,N_13141);
xor U18878 (N_18878,N_15219,N_13088);
and U18879 (N_18879,N_12372,N_14726);
xnor U18880 (N_18880,N_16169,N_12749);
nor U18881 (N_18881,N_14649,N_14058);
and U18882 (N_18882,N_17081,N_17711);
or U18883 (N_18883,N_15640,N_14579);
or U18884 (N_18884,N_13655,N_15569);
or U18885 (N_18885,N_15535,N_15585);
xnor U18886 (N_18886,N_14143,N_17214);
nand U18887 (N_18887,N_16807,N_16015);
nand U18888 (N_18888,N_12003,N_16667);
and U18889 (N_18889,N_12096,N_15186);
nand U18890 (N_18890,N_16178,N_12267);
xnor U18891 (N_18891,N_14234,N_14421);
xnor U18892 (N_18892,N_12556,N_12087);
or U18893 (N_18893,N_12399,N_14774);
nor U18894 (N_18894,N_13944,N_15336);
nor U18895 (N_18895,N_16725,N_14788);
xor U18896 (N_18896,N_14057,N_17935);
xnor U18897 (N_18897,N_16054,N_15643);
nand U18898 (N_18898,N_13375,N_15343);
xor U18899 (N_18899,N_13365,N_16970);
nand U18900 (N_18900,N_13071,N_16074);
xnor U18901 (N_18901,N_13166,N_12902);
and U18902 (N_18902,N_15071,N_13243);
nor U18903 (N_18903,N_16088,N_12146);
nand U18904 (N_18904,N_15039,N_15717);
and U18905 (N_18905,N_13049,N_17023);
nand U18906 (N_18906,N_17995,N_14283);
xnor U18907 (N_18907,N_13772,N_15818);
xor U18908 (N_18908,N_17621,N_14302);
or U18909 (N_18909,N_14909,N_16690);
and U18910 (N_18910,N_13798,N_15856);
nand U18911 (N_18911,N_14214,N_12977);
nand U18912 (N_18912,N_15529,N_15006);
and U18913 (N_18913,N_16191,N_13652);
or U18914 (N_18914,N_13121,N_13754);
or U18915 (N_18915,N_13460,N_16611);
or U18916 (N_18916,N_15998,N_16271);
or U18917 (N_18917,N_15348,N_17843);
and U18918 (N_18918,N_16750,N_12205);
and U18919 (N_18919,N_16139,N_13605);
or U18920 (N_18920,N_16412,N_14290);
xor U18921 (N_18921,N_13852,N_12407);
xor U18922 (N_18922,N_16747,N_13393);
xnor U18923 (N_18923,N_14223,N_13609);
nor U18924 (N_18924,N_15354,N_12970);
nand U18925 (N_18925,N_17938,N_13125);
or U18926 (N_18926,N_17797,N_16051);
and U18927 (N_18927,N_14505,N_17286);
or U18928 (N_18928,N_13818,N_13188);
nand U18929 (N_18929,N_12699,N_17480);
nor U18930 (N_18930,N_16757,N_12627);
xor U18931 (N_18931,N_13755,N_17884);
and U18932 (N_18932,N_17813,N_17419);
nand U18933 (N_18933,N_15850,N_17175);
xor U18934 (N_18934,N_16418,N_16117);
nand U18935 (N_18935,N_16872,N_17487);
or U18936 (N_18936,N_16625,N_13866);
xor U18937 (N_18937,N_14703,N_14307);
and U18938 (N_18938,N_17986,N_17865);
xnor U18939 (N_18939,N_12641,N_14299);
and U18940 (N_18940,N_12645,N_13193);
and U18941 (N_18941,N_17901,N_13449);
or U18942 (N_18942,N_15093,N_14934);
nand U18943 (N_18943,N_14821,N_12281);
nor U18944 (N_18944,N_14961,N_14408);
nand U18945 (N_18945,N_14318,N_15345);
or U18946 (N_18946,N_17129,N_14423);
nand U18947 (N_18947,N_13846,N_14483);
and U18948 (N_18948,N_16294,N_13159);
or U18949 (N_18949,N_17371,N_16741);
xor U18950 (N_18950,N_12067,N_15436);
nand U18951 (N_18951,N_13180,N_16138);
and U18952 (N_18952,N_15623,N_13311);
nor U18953 (N_18953,N_17343,N_12675);
and U18954 (N_18954,N_15197,N_15658);
or U18955 (N_18955,N_12286,N_15793);
nand U18956 (N_18956,N_13597,N_14337);
nor U18957 (N_18957,N_15392,N_16527);
xnor U18958 (N_18958,N_16477,N_17434);
nand U18959 (N_18959,N_15242,N_13407);
xnor U18960 (N_18960,N_14773,N_15675);
and U18961 (N_18961,N_14641,N_14925);
and U18962 (N_18962,N_15049,N_16444);
nand U18963 (N_18963,N_15961,N_15011);
or U18964 (N_18964,N_13292,N_16511);
nand U18965 (N_18965,N_15539,N_12852);
and U18966 (N_18966,N_15743,N_15377);
xor U18967 (N_18967,N_15248,N_12517);
nor U18968 (N_18968,N_17116,N_12880);
or U18969 (N_18969,N_12582,N_12176);
and U18970 (N_18970,N_17658,N_16338);
nand U18971 (N_18971,N_14545,N_17271);
xnor U18972 (N_18972,N_12253,N_16641);
and U18973 (N_18973,N_12117,N_13761);
nor U18974 (N_18974,N_17529,N_15920);
nand U18975 (N_18975,N_13578,N_15233);
nand U18976 (N_18976,N_17206,N_15442);
and U18977 (N_18977,N_13890,N_12866);
or U18978 (N_18978,N_15267,N_14632);
xor U18979 (N_18979,N_15828,N_17264);
and U18980 (N_18980,N_17133,N_15603);
and U18981 (N_18981,N_12704,N_17337);
and U18982 (N_18982,N_17001,N_15430);
xnor U18983 (N_18983,N_12815,N_12368);
nand U18984 (N_18984,N_17122,N_14494);
xor U18985 (N_18985,N_17220,N_16478);
nor U18986 (N_18986,N_13395,N_12774);
xnor U18987 (N_18987,N_13630,N_14341);
nor U18988 (N_18988,N_12816,N_15511);
or U18989 (N_18989,N_13470,N_17429);
nor U18990 (N_18990,N_17636,N_15116);
and U18991 (N_18991,N_16551,N_14153);
and U18992 (N_18992,N_12720,N_16703);
and U18993 (N_18993,N_13408,N_15917);
nor U18994 (N_18994,N_14906,N_12921);
nor U18995 (N_18995,N_16496,N_15161);
nor U18996 (N_18996,N_16313,N_16516);
nor U18997 (N_18997,N_13295,N_14511);
nand U18998 (N_18998,N_17376,N_17646);
or U18999 (N_18999,N_17250,N_14865);
or U19000 (N_19000,N_13785,N_16737);
nand U19001 (N_19001,N_16733,N_17530);
xnor U19002 (N_19002,N_14409,N_15790);
xor U19003 (N_19003,N_13905,N_13008);
nor U19004 (N_19004,N_13428,N_14004);
nand U19005 (N_19005,N_13224,N_17445);
or U19006 (N_19006,N_14577,N_14943);
xor U19007 (N_19007,N_15721,N_12423);
nand U19008 (N_19008,N_12849,N_17723);
or U19009 (N_19009,N_15338,N_14931);
nand U19010 (N_19010,N_12812,N_12031);
nor U19011 (N_19011,N_14643,N_16090);
or U19012 (N_19012,N_17822,N_13555);
nor U19013 (N_19013,N_14651,N_16217);
nor U19014 (N_19014,N_13352,N_17218);
nor U19015 (N_19015,N_17035,N_17546);
or U19016 (N_19016,N_14875,N_15320);
nand U19017 (N_19017,N_14072,N_12259);
xnor U19018 (N_19018,N_14616,N_14655);
nand U19019 (N_19019,N_12199,N_17267);
and U19020 (N_19020,N_12078,N_13518);
nand U19021 (N_19021,N_15397,N_17538);
xnor U19022 (N_19022,N_16709,N_15398);
nand U19023 (N_19023,N_15922,N_14310);
nand U19024 (N_19024,N_12997,N_15316);
or U19025 (N_19025,N_17595,N_13252);
or U19026 (N_19026,N_14617,N_15252);
nor U19027 (N_19027,N_17651,N_13826);
xor U19028 (N_19028,N_14748,N_15649);
or U19029 (N_19029,N_17037,N_13615);
or U19030 (N_19030,N_14707,N_14243);
and U19031 (N_19031,N_12465,N_13341);
nand U19032 (N_19032,N_14475,N_16228);
nor U19033 (N_19033,N_14258,N_15059);
or U19034 (N_19034,N_13533,N_13575);
and U19035 (N_19035,N_16790,N_17211);
nor U19036 (N_19036,N_17504,N_12904);
xnor U19037 (N_19037,N_13324,N_14599);
nand U19038 (N_19038,N_12240,N_16394);
xor U19039 (N_19039,N_14433,N_15433);
nor U19040 (N_19040,N_17306,N_14908);
nand U19041 (N_19041,N_13403,N_16983);
nand U19042 (N_19042,N_16534,N_16399);
and U19043 (N_19043,N_15337,N_13823);
nor U19044 (N_19044,N_13808,N_15547);
nor U19045 (N_19045,N_17737,N_16649);
xor U19046 (N_19046,N_15405,N_12697);
nand U19047 (N_19047,N_16930,N_14491);
nor U19048 (N_19048,N_17425,N_12059);
nor U19049 (N_19049,N_16258,N_17668);
and U19050 (N_19050,N_13545,N_16596);
xor U19051 (N_19051,N_15001,N_16780);
and U19052 (N_19052,N_12601,N_15448);
nor U19053 (N_19053,N_16728,N_16059);
or U19054 (N_19054,N_12154,N_12037);
and U19055 (N_19055,N_14562,N_14945);
nand U19056 (N_19056,N_16125,N_16836);
or U19057 (N_19057,N_14886,N_14711);
and U19058 (N_19058,N_16135,N_13531);
nor U19059 (N_19059,N_15515,N_17130);
nand U19060 (N_19060,N_16022,N_14500);
xnor U19061 (N_19061,N_17012,N_14678);
nand U19062 (N_19062,N_14968,N_17616);
and U19063 (N_19063,N_15680,N_16650);
xor U19064 (N_19064,N_12763,N_16614);
nand U19065 (N_19065,N_17372,N_17507);
nand U19066 (N_19066,N_17700,N_13027);
nand U19067 (N_19067,N_15750,N_15241);
and U19068 (N_19068,N_16687,N_16257);
xor U19069 (N_19069,N_15302,N_12546);
nand U19070 (N_19070,N_14343,N_15779);
and U19071 (N_19071,N_15153,N_17096);
or U19072 (N_19072,N_14189,N_13572);
and U19073 (N_19073,N_14674,N_17145);
or U19074 (N_19074,N_17758,N_16772);
nor U19075 (N_19075,N_12512,N_13383);
nand U19076 (N_19076,N_14154,N_14837);
nand U19077 (N_19077,N_13402,N_15474);
or U19078 (N_19078,N_13894,N_12451);
xnor U19079 (N_19079,N_15160,N_17163);
nor U19080 (N_19080,N_16075,N_15827);
xnor U19081 (N_19081,N_12940,N_12793);
or U19082 (N_19082,N_16556,N_12710);
or U19083 (N_19083,N_12074,N_14320);
nor U19084 (N_19084,N_17821,N_13627);
xor U19085 (N_19085,N_14972,N_13040);
nor U19086 (N_19086,N_16782,N_12312);
or U19087 (N_19087,N_12525,N_16954);
xnor U19088 (N_19088,N_14529,N_16882);
and U19089 (N_19089,N_15616,N_17525);
nor U19090 (N_19090,N_17783,N_15875);
xor U19091 (N_19091,N_14789,N_13210);
nor U19092 (N_19092,N_16542,N_17637);
and U19093 (N_19093,N_12455,N_12356);
xor U19094 (N_19094,N_13548,N_12321);
or U19095 (N_19095,N_14388,N_13617);
and U19096 (N_19096,N_17956,N_12738);
and U19097 (N_19097,N_16572,N_14480);
and U19098 (N_19098,N_16870,N_15512);
or U19099 (N_19099,N_14619,N_15493);
nor U19100 (N_19100,N_17165,N_13995);
nand U19101 (N_19101,N_13758,N_12105);
xor U19102 (N_19102,N_16013,N_14117);
nor U19103 (N_19103,N_15073,N_15091);
or U19104 (N_19104,N_13720,N_13631);
xnor U19105 (N_19105,N_15117,N_17363);
nor U19106 (N_19106,N_17029,N_14523);
xnor U19107 (N_19107,N_15733,N_12338);
or U19108 (N_19108,N_12273,N_13322);
nor U19109 (N_19109,N_17873,N_14037);
and U19110 (N_19110,N_15414,N_14884);
nand U19111 (N_19111,N_13339,N_16846);
nand U19112 (N_19112,N_12098,N_17626);
or U19113 (N_19113,N_13477,N_12712);
nand U19114 (N_19114,N_12552,N_16934);
or U19115 (N_19115,N_14613,N_13701);
nor U19116 (N_19116,N_16065,N_12048);
and U19117 (N_19117,N_17790,N_15933);
nor U19118 (N_19118,N_12813,N_17255);
or U19119 (N_19119,N_15412,N_17719);
nor U19120 (N_19120,N_12887,N_16793);
nor U19121 (N_19121,N_13714,N_16721);
and U19122 (N_19122,N_14265,N_14260);
nand U19123 (N_19123,N_13536,N_14986);
nand U19124 (N_19124,N_13144,N_12443);
xnor U19125 (N_19125,N_17026,N_16949);
nor U19126 (N_19126,N_17324,N_14885);
and U19127 (N_19127,N_14706,N_17936);
and U19128 (N_19128,N_13596,N_12247);
and U19129 (N_19129,N_17506,N_17167);
nor U19130 (N_19130,N_14919,N_14435);
xnor U19131 (N_19131,N_17840,N_12667);
nand U19132 (N_19132,N_12723,N_13982);
nor U19133 (N_19133,N_17170,N_12390);
nor U19134 (N_19134,N_17028,N_12125);
and U19135 (N_19135,N_14447,N_12827);
or U19136 (N_19136,N_13409,N_13174);
nand U19137 (N_19137,N_13195,N_15268);
or U19138 (N_19138,N_12266,N_15584);
nand U19139 (N_19139,N_17113,N_17157);
xnor U19140 (N_19140,N_16184,N_17716);
or U19141 (N_19141,N_15204,N_17423);
or U19142 (N_19142,N_12300,N_15646);
nor U19143 (N_19143,N_16799,N_13579);
xor U19144 (N_19144,N_15394,N_12674);
xnor U19145 (N_19145,N_12086,N_14390);
and U19146 (N_19146,N_14765,N_15310);
xnor U19147 (N_19147,N_16000,N_13423);
nand U19148 (N_19148,N_15771,N_17659);
and U19149 (N_19149,N_16996,N_13789);
nor U19150 (N_19150,N_12417,N_12914);
xor U19151 (N_19151,N_15191,N_17912);
nand U19152 (N_19152,N_14049,N_14999);
or U19153 (N_19153,N_17687,N_17179);
or U19154 (N_19154,N_12421,N_13624);
nor U19155 (N_19155,N_12362,N_14970);
and U19156 (N_19156,N_17837,N_16705);
or U19157 (N_19157,N_15958,N_13592);
or U19158 (N_19158,N_13347,N_15797);
nor U19159 (N_19159,N_15105,N_15916);
xnor U19160 (N_19160,N_17397,N_14650);
or U19161 (N_19161,N_16989,N_15669);
xnor U19162 (N_19162,N_16380,N_15409);
nand U19163 (N_19163,N_14402,N_16151);
nand U19164 (N_19164,N_16322,N_13570);
nand U19165 (N_19165,N_16318,N_14289);
or U19166 (N_19166,N_12791,N_15165);
or U19167 (N_19167,N_15782,N_16506);
xor U19168 (N_19168,N_16912,N_13562);
and U19169 (N_19169,N_14574,N_16531);
xnor U19170 (N_19170,N_16573,N_17420);
xor U19171 (N_19171,N_17071,N_16545);
nor U19172 (N_19172,N_15297,N_17117);
and U19173 (N_19173,N_14820,N_15155);
nand U19174 (N_19174,N_12186,N_14362);
nor U19175 (N_19175,N_14734,N_14464);
nand U19176 (N_19176,N_17051,N_13491);
or U19177 (N_19177,N_13767,N_12986);
nand U19178 (N_19178,N_12382,N_12204);
and U19179 (N_19179,N_15846,N_13123);
xor U19180 (N_19180,N_16992,N_15586);
xor U19181 (N_19181,N_12611,N_12183);
nor U19182 (N_19182,N_14235,N_16365);
or U19183 (N_19183,N_12242,N_13805);
and U19184 (N_19184,N_17349,N_14824);
nor U19185 (N_19185,N_17144,N_16909);
xnor U19186 (N_19186,N_17580,N_16273);
xnor U19187 (N_19187,N_14257,N_17067);
nand U19188 (N_19188,N_12017,N_14896);
nor U19189 (N_19189,N_15904,N_14525);
xnor U19190 (N_19190,N_17575,N_14573);
nor U19191 (N_19191,N_14794,N_12486);
or U19192 (N_19192,N_13633,N_17345);
or U19193 (N_19193,N_17428,N_13101);
xor U19194 (N_19194,N_14436,N_12314);
nand U19195 (N_19195,N_16238,N_16861);
nand U19196 (N_19196,N_17864,N_17055);
or U19197 (N_19197,N_15837,N_17139);
nor U19198 (N_19198,N_14537,N_17260);
nor U19199 (N_19199,N_16910,N_13662);
xnor U19200 (N_19200,N_13729,N_16448);
xor U19201 (N_19201,N_13462,N_16325);
xnor U19202 (N_19202,N_12564,N_13560);
nand U19203 (N_19203,N_16654,N_16244);
and U19204 (N_19204,N_13302,N_16368);
or U19205 (N_19205,N_16103,N_12442);
and U19206 (N_19206,N_14161,N_15973);
or U19207 (N_19207,N_12028,N_16771);
nor U19208 (N_19208,N_15883,N_13155);
xnor U19209 (N_19209,N_16752,N_12207);
or U19210 (N_19210,N_15714,N_14195);
xnor U19211 (N_19211,N_17934,N_15363);
nor U19212 (N_19212,N_17357,N_13589);
nor U19213 (N_19213,N_14624,N_15524);
and U19214 (N_19214,N_15968,N_13025);
or U19215 (N_19215,N_14763,N_17649);
and U19216 (N_19216,N_13752,N_15114);
or U19217 (N_19217,N_13565,N_12933);
nand U19218 (N_19218,N_16329,N_13291);
nand U19219 (N_19219,N_13119,N_16634);
nor U19220 (N_19220,N_16105,N_12433);
nand U19221 (N_19221,N_15613,N_13741);
nand U19222 (N_19222,N_14662,N_16116);
nand U19223 (N_19223,N_12182,N_15768);
xnor U19224 (N_19224,N_17317,N_15887);
xnor U19225 (N_19225,N_14880,N_12107);
or U19226 (N_19226,N_15881,N_12099);
nand U19227 (N_19227,N_16717,N_12130);
nand U19228 (N_19228,N_15556,N_17566);
nor U19229 (N_19229,N_17905,N_14843);
nand U19230 (N_19230,N_17631,N_12033);
and U19231 (N_19231,N_13686,N_14762);
or U19232 (N_19232,N_13880,N_17911);
or U19233 (N_19233,N_16612,N_13250);
and U19234 (N_19234,N_13231,N_17512);
nor U19235 (N_19235,N_14933,N_14814);
or U19236 (N_19236,N_17190,N_17359);
and U19237 (N_19237,N_15399,N_16328);
xor U19238 (N_19238,N_14891,N_16019);
nor U19239 (N_19239,N_13464,N_16121);
xor U19240 (N_19240,N_15939,N_13020);
nor U19241 (N_19241,N_16240,N_15543);
or U19242 (N_19242,N_16695,N_12227);
nor U19243 (N_19243,N_12958,N_17075);
and U19244 (N_19244,N_12238,N_15439);
or U19245 (N_19245,N_13775,N_15813);
or U19246 (N_19246,N_13057,N_17253);
nand U19247 (N_19247,N_17407,N_16819);
nor U19248 (N_19248,N_15080,N_14791);
xnor U19249 (N_19249,N_12493,N_13083);
nor U19250 (N_19250,N_14378,N_17535);
and U19251 (N_19251,N_15375,N_12175);
nand U19252 (N_19252,N_12378,N_12592);
nor U19253 (N_19253,N_17111,N_12996);
and U19254 (N_19254,N_14697,N_17366);
nor U19255 (N_19255,N_17180,N_13097);
and U19256 (N_19256,N_12510,N_13783);
nor U19257 (N_19257,N_12526,N_14724);
nand U19258 (N_19258,N_13024,N_17018);
xor U19259 (N_19259,N_17212,N_12737);
or U19260 (N_19260,N_14499,N_15988);
nand U19261 (N_19261,N_13814,N_15123);
or U19262 (N_19262,N_15609,N_17143);
nor U19263 (N_19263,N_16885,N_16241);
nor U19264 (N_19264,N_16839,N_17513);
xor U19265 (N_19265,N_14677,N_14335);
nor U19266 (N_19266,N_17980,N_15212);
nand U19267 (N_19267,N_12482,N_17667);
or U19268 (N_19268,N_16927,N_12121);
and U19269 (N_19269,N_14803,N_17556);
or U19270 (N_19270,N_16829,N_12733);
xor U19271 (N_19271,N_16070,N_14319);
nor U19272 (N_19272,N_13378,N_16006);
or U19273 (N_19273,N_13691,N_13810);
or U19274 (N_19274,N_17265,N_12301);
xor U19275 (N_19275,N_17820,N_16462);
xor U19276 (N_19276,N_14191,N_13683);
xor U19277 (N_19277,N_15801,N_12754);
nand U19278 (N_19278,N_16339,N_12599);
xor U19279 (N_19279,N_16617,N_17025);
or U19280 (N_19280,N_17593,N_12777);
nor U19281 (N_19281,N_15876,N_12936);
and U19282 (N_19282,N_17715,N_14929);
nor U19283 (N_19283,N_15844,N_15825);
nand U19284 (N_19284,N_16937,N_13359);
xnor U19285 (N_19285,N_17655,N_15121);
nand U19286 (N_19286,N_13344,N_14085);
and U19287 (N_19287,N_17652,N_17352);
xnor U19288 (N_19288,N_13678,N_16393);
and U19289 (N_19289,N_12077,N_15656);
nor U19290 (N_19290,N_17965,N_14198);
and U19291 (N_19291,N_15823,N_12553);
xnor U19292 (N_19292,N_16205,N_13330);
xor U19293 (N_19293,N_13168,N_17430);
or U19294 (N_19294,N_12892,N_15738);
or U19295 (N_19295,N_13146,N_15608);
and U19296 (N_19296,N_14553,N_13945);
xnor U19297 (N_19297,N_15918,N_13236);
xor U19298 (N_19298,N_13348,N_16643);
and U19299 (N_19299,N_12690,N_12166);
nor U19300 (N_19300,N_14597,N_15464);
and U19301 (N_19301,N_16540,N_16536);
nand U19302 (N_19302,N_12714,N_12797);
nand U19303 (N_19303,N_12854,N_14568);
or U19304 (N_19304,N_13029,N_17181);
or U19305 (N_19305,N_16290,N_16481);
nand U19306 (N_19306,N_16632,N_16896);
nand U19307 (N_19307,N_17340,N_13829);
and U19308 (N_19308,N_16563,N_17446);
nor U19309 (N_19309,N_12978,N_14199);
and U19310 (N_19310,N_14285,N_14965);
and U19311 (N_19311,N_14905,N_12057);
nor U19312 (N_19312,N_16374,N_15386);
or U19313 (N_19313,N_16604,N_12345);
or U19314 (N_19314,N_12397,N_14539);
xnor U19315 (N_19315,N_14145,N_16175);
or U19316 (N_19316,N_16312,N_15833);
nor U19317 (N_19317,N_12180,N_13067);
nand U19318 (N_19318,N_14838,N_16998);
nand U19319 (N_19319,N_16094,N_12701);
nand U19320 (N_19320,N_17609,N_13511);
xor U19321 (N_19321,N_17455,N_16490);
xor U19322 (N_19322,N_12264,N_12441);
nor U19323 (N_19323,N_13011,N_14363);
and U19324 (N_19324,N_15164,N_13153);
and U19325 (N_19325,N_16950,N_12908);
nand U19326 (N_19326,N_12745,N_15729);
nand U19327 (N_19327,N_15192,N_15963);
or U19328 (N_19328,N_14563,N_16948);
xor U19329 (N_19329,N_13505,N_15606);
nor U19330 (N_19330,N_15554,N_16759);
nand U19331 (N_19331,N_17451,N_16491);
xnor U19332 (N_19332,N_14292,N_16710);
nand U19333 (N_19333,N_13726,N_12795);
or U19334 (N_19334,N_15636,N_15975);
xor U19335 (N_19335,N_12336,N_14410);
xor U19336 (N_19336,N_17866,N_12211);
or U19337 (N_19337,N_17960,N_15360);
nor U19338 (N_19338,N_15218,N_16761);
xor U19339 (N_19339,N_12163,N_16043);
xor U19340 (N_19340,N_16432,N_17584);
nor U19341 (N_19341,N_12729,N_16843);
or U19342 (N_19342,N_13552,N_14066);
nand U19343 (N_19343,N_13503,N_12481);
xor U19344 (N_19344,N_14897,N_16620);
and U19345 (N_19345,N_16662,N_17793);
xnor U19346 (N_19346,N_16308,N_15162);
xnor U19347 (N_19347,N_13006,N_15349);
nand U19348 (N_19348,N_15280,N_14739);
nand U19349 (N_19349,N_14498,N_13853);
or U19350 (N_19350,N_14873,N_12013);
nor U19351 (N_19351,N_14399,N_16691);
or U19352 (N_19352,N_15571,N_14963);
nor U19353 (N_19353,N_13446,N_14594);
or U19354 (N_19354,N_13925,N_15816);
xnor U19355 (N_19355,N_15832,N_17736);
xor U19356 (N_19356,N_12352,N_12055);
and U19357 (N_19357,N_15820,N_17355);
nor U19358 (N_19358,N_14672,N_14854);
nor U19359 (N_19359,N_14280,N_16235);
nand U19360 (N_19360,N_14132,N_16446);
nand U19361 (N_19361,N_13418,N_17872);
nand U19362 (N_19362,N_16187,N_12935);
or U19363 (N_19363,N_17109,N_16773);
nor U19364 (N_19364,N_13736,N_15180);
xor U19365 (N_19365,N_15490,N_17971);
nor U19366 (N_19366,N_16337,N_12828);
xor U19367 (N_19367,N_14422,N_14210);
nand U19368 (N_19368,N_12625,N_13053);
nor U19369 (N_19369,N_15992,N_15016);
nand U19370 (N_19370,N_13218,N_15713);
or U19371 (N_19371,N_12806,N_15036);
nor U19372 (N_19372,N_17382,N_14196);
nor U19373 (N_19373,N_16849,N_12859);
nand U19374 (N_19374,N_12463,N_15357);
xnor U19375 (N_19375,N_16425,N_13935);
or U19376 (N_19376,N_13177,N_16785);
or U19377 (N_19377,N_15179,N_14555);
nand U19378 (N_19378,N_14385,N_13499);
xnor U19379 (N_19379,N_12506,N_13334);
or U19380 (N_19380,N_14152,N_15452);
nand U19381 (N_19381,N_17645,N_14799);
and U19382 (N_19382,N_17819,N_15434);
xnor U19383 (N_19383,N_15195,N_14394);
and U19384 (N_19384,N_13315,N_15142);
nor U19385 (N_19385,N_12097,N_17230);
xnor U19386 (N_19386,N_13355,N_17189);
xor U19387 (N_19387,N_12467,N_15030);
nand U19388 (N_19388,N_17239,N_14778);
xor U19389 (N_19389,N_16837,N_17215);
xnor U19390 (N_19390,N_13257,N_14178);
and U19391 (N_19391,N_15764,N_16698);
nor U19392 (N_19392,N_12492,N_13868);
and U19393 (N_19393,N_12919,N_12079);
xnor U19394 (N_19394,N_12927,N_14023);
nand U19395 (N_19395,N_15601,N_13289);
nand U19396 (N_19396,N_17775,N_13763);
xnor U19397 (N_19397,N_12554,N_14669);
or U19398 (N_19398,N_16366,N_17336);
nand U19399 (N_19399,N_15088,N_15652);
xnor U19400 (N_19400,N_15428,N_16984);
nor U19401 (N_19401,N_12772,N_15538);
and U19402 (N_19402,N_16252,N_13030);
xnor U19403 (N_19403,N_17056,N_14920);
nor U19404 (N_19404,N_17746,N_12440);
nand U19405 (N_19405,N_15435,N_14536);
and U19406 (N_19406,N_12541,N_13614);
nand U19407 (N_19407,N_13582,N_15416);
and U19408 (N_19408,N_15056,N_16616);
and U19409 (N_19409,N_17786,N_12527);
and U19410 (N_19410,N_14973,N_12724);
nor U19411 (N_19411,N_16476,N_15220);
nor U19412 (N_19412,N_16422,N_16111);
nor U19413 (N_19413,N_16295,N_14979);
and U19414 (N_19414,N_17323,N_16602);
or U19415 (N_19415,N_16424,N_14281);
or U19416 (N_19416,N_17570,N_15727);
or U19417 (N_19417,N_12836,N_14345);
xnor U19418 (N_19418,N_14204,N_15668);
or U19419 (N_19419,N_12985,N_16369);
nor U19420 (N_19420,N_15991,N_14045);
xor U19421 (N_19421,N_12719,N_16713);
and U19422 (N_19422,N_12234,N_17332);
or U19423 (N_19423,N_14176,N_12809);
xnor U19424 (N_19424,N_12054,N_13254);
nor U19425 (N_19425,N_12566,N_17161);
or U19426 (N_19426,N_12637,N_14956);
nor U19427 (N_19427,N_14593,N_16227);
or U19428 (N_19428,N_15298,N_13126);
nand U19429 (N_19429,N_13299,N_14291);
nor U19430 (N_19430,N_17605,N_14831);
nor U19431 (N_19431,N_12095,N_17877);
nand U19432 (N_19432,N_14271,N_15795);
nand U19433 (N_19433,N_17290,N_16172);
nor U19434 (N_19434,N_15903,N_12889);
xor U19435 (N_19435,N_16781,N_13495);
and U19436 (N_19436,N_15315,N_17398);
and U19437 (N_19437,N_14951,N_15395);
or U19438 (N_19438,N_17034,N_16150);
nor U19439 (N_19439,N_12883,N_12606);
xnor U19440 (N_19440,N_16976,N_13285);
xnor U19441 (N_19441,N_13577,N_16465);
and U19442 (N_19442,N_13397,N_13881);
or U19443 (N_19443,N_15666,N_12395);
and U19444 (N_19444,N_16933,N_14015);
nor U19445 (N_19445,N_16631,N_15225);
and U19446 (N_19446,N_12695,N_12167);
xor U19447 (N_19447,N_15072,N_16944);
nor U19448 (N_19448,N_17494,N_12075);
nand U19449 (N_19449,N_14856,N_15999);
xnor U19450 (N_19450,N_17839,N_12181);
nand U19451 (N_19451,N_13012,N_16155);
xnor U19452 (N_19452,N_14346,N_13328);
nor U19453 (N_19453,N_12586,N_14779);
and U19454 (N_19454,N_16436,N_17014);
nand U19455 (N_19455,N_15570,N_13745);
nor U19456 (N_19456,N_16729,N_12583);
nand U19457 (N_19457,N_12534,N_12721);
nand U19458 (N_19458,N_14671,N_12647);
nor U19459 (N_19459,N_14715,N_14110);
nor U19460 (N_19460,N_17209,N_15671);
or U19461 (N_19461,N_14395,N_16426);
nor U19462 (N_19462,N_12379,N_13164);
nor U19463 (N_19463,N_15009,N_17226);
xor U19464 (N_19464,N_16745,N_15564);
xnor U19465 (N_19465,N_14114,N_16528);
nor U19466 (N_19466,N_16575,N_15678);
and U19467 (N_19467,N_12905,N_16735);
nand U19468 (N_19468,N_16349,N_14349);
nand U19469 (N_19469,N_16853,N_12753);
nor U19470 (N_19470,N_14696,N_15965);
xor U19471 (N_19471,N_16860,N_17321);
nand U19472 (N_19472,N_13278,N_13913);
nand U19473 (N_19473,N_14874,N_12371);
or U19474 (N_19474,N_12051,N_15347);
nor U19475 (N_19475,N_15174,N_16214);
nand U19476 (N_19476,N_12705,N_14278);
or U19477 (N_19477,N_14509,N_13684);
and U19478 (N_19478,N_14373,N_13102);
nor U19479 (N_19479,N_17656,N_16859);
xor U19480 (N_19480,N_12619,N_15361);
or U19481 (N_19481,N_13056,N_13862);
and U19482 (N_19482,N_12614,N_15251);
nand U19483 (N_19483,N_16915,N_14105);
nor U19484 (N_19484,N_16423,N_12065);
nor U19485 (N_19485,N_12090,N_16815);
nand U19486 (N_19486,N_14975,N_14569);
and U19487 (N_19487,N_16567,N_15211);
nand U19488 (N_19488,N_13329,N_12094);
and U19489 (N_19489,N_16403,N_14630);
or U19490 (N_19490,N_14752,N_17549);
and U19491 (N_19491,N_16856,N_15223);
nand U19492 (N_19492,N_14332,N_14834);
or U19493 (N_19493,N_12108,N_12903);
and U19494 (N_19494,N_15597,N_13160);
xnor U19495 (N_19495,N_12551,N_12169);
or U19496 (N_19496,N_13864,N_13127);
xor U19497 (N_19497,N_14141,N_17408);
or U19498 (N_19498,N_13992,N_16600);
nor U19499 (N_19499,N_14472,N_13986);
nand U19500 (N_19500,N_12328,N_15008);
xor U19501 (N_19501,N_15540,N_12702);
or U19502 (N_19502,N_12585,N_16128);
nor U19503 (N_19503,N_16878,N_17274);
xor U19504 (N_19504,N_12373,N_12047);
nor U19505 (N_19505,N_14439,N_12912);
nor U19506 (N_19506,N_16469,N_16400);
nand U19507 (N_19507,N_17188,N_17910);
nand U19508 (N_19508,N_17921,N_12744);
or U19509 (N_19509,N_12776,N_13634);
xnor U19510 (N_19510,N_15082,N_14845);
xor U19511 (N_19511,N_15019,N_16935);
and U19512 (N_19512,N_14572,N_16285);
xor U19513 (N_19513,N_14665,N_16906);
or U19514 (N_19514,N_17171,N_14589);
and U19515 (N_19515,N_15206,N_12178);
and U19516 (N_19516,N_15130,N_17950);
nand U19517 (N_19517,N_14801,N_15385);
or U19518 (N_19518,N_15157,N_13353);
xor U19519 (N_19519,N_12032,N_17422);
or U19520 (N_19520,N_15138,N_14581);
xnor U19521 (N_19521,N_13656,N_17594);
nor U19522 (N_19522,N_15710,N_12277);
nor U19523 (N_19523,N_16558,N_16678);
and U19524 (N_19524,N_16267,N_12413);
nor U19525 (N_19525,N_17383,N_16648);
or U19526 (N_19526,N_14741,N_16210);
nor U19527 (N_19527,N_17417,N_16221);
nor U19528 (N_19528,N_15496,N_15667);
nand U19529 (N_19529,N_14924,N_17847);
nand U19530 (N_19530,N_12319,N_12334);
nand U19531 (N_19531,N_12161,N_13498);
nand U19532 (N_19532,N_12768,N_13273);
nor U19533 (N_19533,N_16809,N_13756);
nor U19534 (N_19534,N_14262,N_16553);
and U19535 (N_19535,N_16133,N_17093);
xor U19536 (N_19536,N_13688,N_17776);
nand U19537 (N_19537,N_16453,N_15693);
nor U19538 (N_19538,N_15532,N_15720);
nor U19539 (N_19539,N_16660,N_15896);
xnor U19540 (N_19540,N_13107,N_16580);
and U19541 (N_19541,N_15388,N_13276);
xor U19542 (N_19542,N_17868,N_13869);
and U19543 (N_19543,N_12646,N_14393);
xnor U19544 (N_19544,N_14802,N_15522);
nor U19545 (N_19545,N_13594,N_17172);
nor U19546 (N_19546,N_15314,N_13149);
nand U19547 (N_19547,N_13388,N_14089);
or U19548 (N_19548,N_13034,N_15957);
xnor U19549 (N_19549,N_17069,N_14095);
or U19550 (N_19550,N_15924,N_17207);
and U19551 (N_19551,N_16967,N_17015);
and U19552 (N_19552,N_13092,N_14321);
xor U19553 (N_19553,N_12022,N_13663);
nand U19554 (N_19554,N_14311,N_16445);
xnor U19555 (N_19555,N_17598,N_14826);
and U19556 (N_19556,N_13436,N_15120);
and U19557 (N_19557,N_12890,N_14712);
nand U19558 (N_19558,N_15159,N_15766);
xor U19559 (N_19559,N_16298,N_13891);
nand U19560 (N_19560,N_14663,N_12536);
nand U19561 (N_19561,N_17009,N_17017);
xor U19562 (N_19562,N_17240,N_13392);
and U19563 (N_19563,N_16154,N_13815);
xnor U19564 (N_19564,N_12673,N_16464);
nand U19565 (N_19565,N_12311,N_16651);
nand U19566 (N_19566,N_15007,N_13855);
and U19567 (N_19567,N_13718,N_16956);
nor U19568 (N_19568,N_12302,N_16925);
nand U19569 (N_19569,N_12869,N_17162);
nand U19570 (N_19570,N_15182,N_14401);
nor U19571 (N_19571,N_13298,N_16862);
nand U19572 (N_19572,N_15819,N_16897);
xnor U19573 (N_19573,N_17579,N_12152);
nand U19574 (N_19574,N_12456,N_17103);
nor U19575 (N_19575,N_16077,N_14159);
nor U19576 (N_19576,N_14162,N_14603);
or U19577 (N_19577,N_16208,N_15492);
or U19578 (N_19578,N_17369,N_16225);
and U19579 (N_19579,N_15575,N_17127);
nand U19580 (N_19580,N_13607,N_15696);
or U19581 (N_19581,N_13970,N_13421);
nor U19582 (N_19582,N_16823,N_15034);
and U19583 (N_19583,N_17660,N_16594);
nand U19584 (N_19584,N_15765,N_14194);
and U19585 (N_19585,N_17106,N_12848);
and U19586 (N_19586,N_13461,N_12679);
nor U19587 (N_19587,N_15070,N_17806);
xor U19588 (N_19588,N_14063,N_14091);
or U19589 (N_19589,N_15096,N_17683);
nor U19590 (N_19590,N_14338,N_13803);
xor U19591 (N_19591,N_13938,N_13502);
nand U19592 (N_19592,N_15523,N_16835);
or U19593 (N_19593,N_15647,N_14497);
and U19594 (N_19594,N_15500,N_16618);
nand U19595 (N_19595,N_14150,N_15489);
and U19596 (N_19596,N_15175,N_13781);
or U19597 (N_19597,N_13084,N_12682);
and U19598 (N_19598,N_17022,N_14164);
or U19599 (N_19599,N_15373,N_16566);
or U19600 (N_19600,N_12778,N_17984);
nand U19601 (N_19601,N_16031,N_17147);
nand U19602 (N_19602,N_16693,N_13708);
nand U19603 (N_19603,N_16565,N_17829);
and U19604 (N_19604,N_14484,N_17951);
or U19605 (N_19605,N_13896,N_13047);
xnor U19606 (N_19606,N_14993,N_17470);
nand U19607 (N_19607,N_17142,N_13621);
nor U19608 (N_19608,N_12757,N_12409);
nand U19609 (N_19609,N_14812,N_14626);
xor U19610 (N_19610,N_15144,N_16971);
xnor U19611 (N_19611,N_13844,N_15438);
nand U19612 (N_19612,N_17384,N_13672);
xor U19613 (N_19613,N_16283,N_14871);
nand U19614 (N_19614,N_12225,N_14478);
xnor U19615 (N_19615,N_14456,N_16229);
nor U19616 (N_19616,N_16375,N_14201);
and U19617 (N_19617,N_15810,N_13874);
or U19618 (N_19618,N_16034,N_15215);
xnor U19619 (N_19619,N_14817,N_14502);
xnor U19620 (N_19620,N_17541,N_14426);
and U19621 (N_19621,N_16039,N_17228);
nor U19622 (N_19622,N_13922,N_12818);
nand U19623 (N_19623,N_16907,N_14957);
and U19624 (N_19624,N_12422,N_15229);
or U19625 (N_19625,N_17125,N_15112);
nand U19626 (N_19626,N_17151,N_12335);
nand U19627 (N_19627,N_14157,N_12624);
xnor U19628 (N_19628,N_15558,N_14296);
or U19629 (N_19629,N_14250,N_17684);
nor U19630 (N_19630,N_14206,N_14107);
or U19631 (N_19631,N_16764,N_16633);
and U19632 (N_19632,N_17724,N_17964);
and U19633 (N_19633,N_15582,N_16623);
nand U19634 (N_19634,N_13448,N_16007);
nor U19635 (N_19635,N_14978,N_15289);
and U19636 (N_19636,N_14653,N_13507);
and U19637 (N_19637,N_14106,N_15989);
xor U19638 (N_19638,N_14786,N_15324);
and U19639 (N_19639,N_17628,N_16903);
nand U19640 (N_19640,N_12783,N_12257);
nand U19641 (N_19641,N_13824,N_14442);
or U19642 (N_19642,N_16941,N_16149);
and U19643 (N_19643,N_15311,N_14927);
nor U19644 (N_19644,N_16522,N_17966);
xnor U19645 (N_19645,N_14728,N_17320);
xor U19646 (N_19646,N_15907,N_14548);
or U19647 (N_19647,N_17642,N_14368);
nor U19648 (N_19648,N_12872,N_13048);
nand U19649 (N_19649,N_14598,N_17774);
xnor U19650 (N_19650,N_16253,N_16675);
xnor U19651 (N_19651,N_16518,N_13841);
and U19652 (N_19652,N_15333,N_13130);
nand U19653 (N_19653,N_16079,N_17493);
xnor U19654 (N_19654,N_13603,N_15115);
nor U19655 (N_19655,N_12110,N_16840);
nand U19656 (N_19656,N_14527,N_16442);
xor U19657 (N_19657,N_15312,N_16250);
or U19658 (N_19658,N_17284,N_14417);
and U19659 (N_19659,N_16040,N_15300);
xnor U19660 (N_19660,N_13996,N_13861);
nor U19661 (N_19661,N_17739,N_12359);
and U19662 (N_19662,N_12408,N_13061);
xnor U19663 (N_19663,N_14798,N_13558);
nor U19664 (N_19664,N_17809,N_12740);
or U19665 (N_19665,N_14682,N_14889);
nand U19666 (N_19666,N_16185,N_13226);
or U19667 (N_19667,N_15749,N_16917);
or U19668 (N_19668,N_17497,N_13978);
nor U19669 (N_19669,N_14514,N_17640);
nand U19670 (N_19670,N_12414,N_13199);
nand U19671 (N_19671,N_17959,N_14027);
nand U19672 (N_19672,N_13709,N_16603);
xor U19673 (N_19673,N_17379,N_17499);
nand U19674 (N_19674,N_14571,N_16898);
nand U19675 (N_19675,N_14460,N_17523);
or U19676 (N_19676,N_15520,N_12571);
and U19677 (N_19677,N_17962,N_13326);
nand U19678 (N_19678,N_13161,N_13169);
or U19679 (N_19679,N_12490,N_12307);
nor U19680 (N_19680,N_13819,N_14113);
or U19681 (N_19681,N_16689,N_17607);
and U19682 (N_19682,N_14087,N_16621);
or U19683 (N_19683,N_14160,N_15283);
nand U19684 (N_19684,N_12604,N_17390);
or U19685 (N_19685,N_12135,N_17874);
and U19686 (N_19686,N_17234,N_12870);
xor U19687 (N_19687,N_17880,N_17857);
nand U19688 (N_19688,N_16415,N_16673);
or U19689 (N_19689,N_15473,N_17812);
nor U19690 (N_19690,N_12748,N_13441);
nand U19691 (N_19691,N_17128,N_14416);
nand U19692 (N_19692,N_14322,N_17070);
xnor U19693 (N_19693,N_13233,N_14284);
xor U19694 (N_19694,N_16724,N_15128);
or U19695 (N_19695,N_12260,N_16156);
nor U19696 (N_19696,N_17156,N_13998);
nand U19697 (N_19697,N_13338,N_17999);
nand U19698 (N_19698,N_12387,N_16979);
nand U19699 (N_19699,N_15912,N_12418);
or U19700 (N_19700,N_15808,N_17878);
xor U19701 (N_19701,N_13192,N_16929);
nand U19702 (N_19702,N_14530,N_13026);
nand U19703 (N_19703,N_17862,N_13390);
nor U19704 (N_19704,N_12118,N_16791);
and U19705 (N_19705,N_12226,N_15639);
or U19706 (N_19706,N_17406,N_12574);
xnor U19707 (N_19707,N_16636,N_17489);
xnor U19708 (N_19708,N_16852,N_15087);
xnor U19709 (N_19709,N_15382,N_15450);
xnor U19710 (N_19710,N_15090,N_16808);
and U19711 (N_19711,N_12998,N_17913);
nand U19712 (N_19712,N_15178,N_14174);
nor U19713 (N_19713,N_17729,N_15707);
xnor U19714 (N_19714,N_12801,N_17276);
xor U19715 (N_19715,N_17979,N_14606);
xor U19716 (N_19716,N_17508,N_13087);
nand U19717 (N_19717,N_16272,N_14261);
and U19718 (N_19718,N_17072,N_13647);
and U19719 (N_19719,N_15050,N_12920);
or U19720 (N_19720,N_12727,N_17168);
nor U19721 (N_19721,N_12332,N_17104);
xnor U19722 (N_19722,N_14003,N_14883);
nor U19723 (N_19723,N_15747,N_13892);
nor U19724 (N_19724,N_14809,N_13883);
nand U19725 (N_19725,N_16776,N_16025);
xor U19726 (N_19726,N_12261,N_15238);
and U19727 (N_19727,N_17763,N_13911);
and U19728 (N_19728,N_13445,N_13135);
xor U19729 (N_19729,N_13138,N_14861);
and U19730 (N_19730,N_17904,N_16136);
nor U19731 (N_19731,N_14142,N_12452);
and U19732 (N_19732,N_12937,N_12092);
nand U19733 (N_19733,N_17300,N_14403);
or U19734 (N_19734,N_12957,N_14760);
nand U19735 (N_19735,N_13820,N_17353);
and U19736 (N_19736,N_17551,N_16249);
and U19737 (N_19737,N_16195,N_14942);
nand U19738 (N_19738,N_14998,N_14926);
nand U19739 (N_19739,N_16190,N_15902);
and U19740 (N_19740,N_15458,N_12023);
nand U19741 (N_19741,N_12007,N_15879);
xor U19742 (N_19742,N_12197,N_13611);
xnor U19743 (N_19743,N_17316,N_16765);
or U19744 (N_19744,N_14583,N_16497);
and U19745 (N_19745,N_15545,N_13836);
nor U19746 (N_19746,N_17564,N_15742);
nor U19747 (N_19747,N_14476,N_16027);
or U19748 (N_19748,N_16084,N_15893);
and U19749 (N_19749,N_15703,N_14158);
nand U19750 (N_19750,N_16501,N_15149);
xnor U19751 (N_19751,N_13304,N_14112);
nand U19752 (N_19752,N_17254,N_14716);
nor U19753 (N_19753,N_13658,N_13695);
nand U19754 (N_19754,N_12788,N_17990);
and U19755 (N_19755,N_17442,N_15127);
nand U19756 (N_19756,N_16726,N_16755);
nand U19757 (N_19757,N_16060,N_16202);
or U19758 (N_19758,N_12700,N_16507);
nor U19759 (N_19759,N_17888,N_17043);
xor U19760 (N_19760,N_17388,N_14857);
or U19761 (N_19761,N_12561,N_17701);
xnor U19762 (N_19762,N_13933,N_12466);
xnor U19763 (N_19763,N_17333,N_17313);
nor U19764 (N_19764,N_13957,N_15243);
xor U19765 (N_19765,N_16157,N_17559);
and U19766 (N_19766,N_15285,N_14200);
nand U19767 (N_19767,N_15199,N_12487);
xnor U19768 (N_19768,N_14550,N_15618);
nand U19769 (N_19769,N_14012,N_12102);
or U19770 (N_19770,N_12229,N_17263);
nor U19771 (N_19771,N_12138,N_17454);
nand U19772 (N_19772,N_15950,N_13979);
xor U19773 (N_19773,N_17040,N_12245);
and U19774 (N_19774,N_16057,N_12591);
nand U19775 (N_19775,N_15614,N_14103);
nor U19776 (N_19776,N_16343,N_14044);
nand U19777 (N_19777,N_12841,N_12722);
nand U19778 (N_19778,N_12549,N_17500);
xor U19779 (N_19779,N_13690,N_17743);
nand U19780 (N_19780,N_16877,N_14138);
or U19781 (N_19781,N_16972,N_13928);
nor U19782 (N_19782,N_14365,N_15402);
nor U19783 (N_19783,N_15454,N_13768);
nor U19784 (N_19784,N_13189,N_17704);
nand U19785 (N_19785,N_12270,N_14893);
or U19786 (N_19786,N_16402,N_13563);
nand U19787 (N_19787,N_13364,N_12072);
or U19788 (N_19788,N_14542,N_12837);
nor U19789 (N_19789,N_12730,N_14151);
or U19790 (N_19790,N_16072,N_14228);
and U19791 (N_19791,N_17404,N_17484);
nand U19792 (N_19792,N_12947,N_13196);
nor U19793 (N_19793,N_15076,N_13717);
and U19794 (N_19794,N_15712,N_13544);
or U19795 (N_19795,N_12629,N_17526);
xor U19796 (N_19796,N_13660,N_12279);
nand U19797 (N_19797,N_16975,N_13506);
nor U19798 (N_19798,N_17058,N_15514);
and U19799 (N_19799,N_15624,N_12878);
nor U19800 (N_19800,N_15031,N_15177);
or U19801 (N_19801,N_12462,N_17734);
and U19802 (N_19802,N_17592,N_16834);
xor U19803 (N_19803,N_16871,N_13707);
and U19804 (N_19804,N_12289,N_17364);
nor U19805 (N_19805,N_12518,N_16756);
nor U19806 (N_19806,N_14988,N_12104);
or U19807 (N_19807,N_12580,N_14111);
xor U19808 (N_19808,N_16668,N_15594);
and U19809 (N_19809,N_13676,N_16456);
nor U19810 (N_19810,N_12404,N_17149);
nand U19811 (N_19811,N_17275,N_15852);
or U19812 (N_19812,N_13983,N_16397);
nand U19813 (N_19813,N_15217,N_12542);
xor U19814 (N_19814,N_12734,N_17796);
nor U19815 (N_19815,N_14013,N_12976);
xnor U19816 (N_19816,N_17244,N_12832);
and U19817 (N_19817,N_15284,N_16331);
xnor U19818 (N_19818,N_12008,N_14810);
and U19819 (N_19819,N_14584,N_14987);
or U19820 (N_19820,N_15845,N_13977);
nand U19821 (N_19821,N_14531,N_14098);
nor U19822 (N_19822,N_17827,N_13990);
xor U19823 (N_19823,N_13245,N_17132);
nand U19824 (N_19824,N_12360,N_13564);
xor U19825 (N_19825,N_12025,N_17046);
xor U19826 (N_19826,N_13406,N_15075);
or U19827 (N_19827,N_15051,N_15226);
nor U19828 (N_19828,N_17611,N_17464);
nor U19829 (N_19829,N_17257,N_14216);
nand U19830 (N_19830,N_17589,N_14102);
and U19831 (N_19831,N_13424,N_12587);
and U19832 (N_19832,N_14064,N_16850);
nand U19833 (N_19833,N_16749,N_14644);
or U19834 (N_19834,N_14912,N_16277);
nor U19835 (N_19835,N_13671,N_16552);
and U19836 (N_19836,N_13190,N_12454);
and U19837 (N_19837,N_16995,N_17119);
or U19838 (N_19838,N_15465,N_14510);
nor U19839 (N_19839,N_16324,N_14036);
or U19840 (N_19840,N_14016,N_13670);
nor U19841 (N_19841,N_14932,N_12779);
nand U19842 (N_19842,N_12123,N_16340);
xnor U19843 (N_19843,N_15984,N_16194);
and U19844 (N_19844,N_14135,N_15139);
or U19845 (N_19845,N_17048,N_17792);
nor U19846 (N_19846,N_17705,N_13411);
or U19847 (N_19847,N_15722,N_16576);
and U19848 (N_19848,N_14119,N_16081);
xor U19849 (N_19849,N_17219,N_12021);
or U19850 (N_19850,N_17146,N_16787);
xnor U19851 (N_19851,N_14792,N_12171);
and U19852 (N_19852,N_17392,N_15726);
nor U19853 (N_19853,N_12502,N_12046);
or U19854 (N_19854,N_17871,N_15807);
nor U19855 (N_19855,N_17665,N_13165);
and U19856 (N_19856,N_13015,N_13346);
xor U19857 (N_19857,N_15905,N_13307);
xor U19858 (N_19858,N_17326,N_16264);
nor U19859 (N_19859,N_13535,N_14121);
xnor U19860 (N_19860,N_14222,N_12071);
or U19861 (N_19861,N_14590,N_15081);
xnor U19862 (N_19862,N_13367,N_17893);
or U19863 (N_19863,N_14852,N_16357);
nor U19864 (N_19864,N_15800,N_14220);
xor U19865 (N_19865,N_13310,N_13832);
xor U19866 (N_19866,N_17988,N_12044);
nor U19867 (N_19867,N_15908,N_15319);
nor U19868 (N_19868,N_17828,N_17741);
nor U19869 (N_19869,N_16683,N_17765);
nor U19870 (N_19870,N_15525,N_16635);
and U19871 (N_19871,N_13644,N_12080);
nor U19872 (N_19872,N_15986,N_17906);
or U19873 (N_19873,N_15472,N_17833);
and U19874 (N_19874,N_17294,N_13429);
nand U19875 (N_19875,N_12350,N_12331);
or U19876 (N_19876,N_14591,N_17671);
and U19877 (N_19877,N_17063,N_17916);
xor U19878 (N_19878,N_12956,N_15274);
or U19879 (N_19879,N_15052,N_12548);
nand U19880 (N_19880,N_13946,N_17557);
nand U19881 (N_19881,N_17485,N_12540);
nor U19882 (N_19882,N_12766,N_13875);
xnor U19883 (N_19883,N_17924,N_17745);
nand U19884 (N_19884,N_14249,N_17516);
or U19885 (N_19885,N_13007,N_16017);
and U19886 (N_19886,N_12449,N_17826);
nor U19887 (N_19887,N_14808,N_16921);
xnor U19888 (N_19888,N_13414,N_13281);
xor U19889 (N_19889,N_12039,N_12683);
and U19890 (N_19890,N_17945,N_17712);
xor U19891 (N_19891,N_13386,N_16420);
nand U19892 (N_19892,N_15829,N_13486);
nand U19893 (N_19893,N_13525,N_15415);
and U19894 (N_19894,N_13942,N_14432);
nand U19895 (N_19895,N_14746,N_15642);
nand U19896 (N_19896,N_12479,N_14742);
or U19897 (N_19897,N_13113,N_13037);
and U19898 (N_19898,N_15503,N_17016);
nor U19899 (N_19899,N_17969,N_16334);
and U19900 (N_19900,N_13747,N_16658);
nand U19901 (N_19901,N_15259,N_16413);
xor U19902 (N_19902,N_17958,N_17823);
nand U19903 (N_19903,N_12684,N_17377);
xnor U19904 (N_19904,N_14658,N_12755);
and U19905 (N_19905,N_14923,N_12195);
or U19906 (N_19906,N_17801,N_15568);
nor U19907 (N_19907,N_12275,N_16546);
xnor U19908 (N_19908,N_17779,N_13036);
or U19909 (N_19909,N_12909,N_16045);
or U19910 (N_19910,N_12907,N_13208);
and U19911 (N_19911,N_16686,N_16114);
and U19912 (N_19912,N_13659,N_17066);
nand U19913 (N_19913,N_16384,N_12374);
nor U19914 (N_19914,N_14212,N_16732);
nand U19915 (N_19915,N_16421,N_13094);
and U19916 (N_19916,N_12370,N_14766);
and U19917 (N_19917,N_17334,N_14173);
and U19918 (N_19918,N_15411,N_13219);
xnor U19919 (N_19919,N_16484,N_17955);
nand U19920 (N_19920,N_12179,N_13251);
or U19921 (N_19921,N_14955,N_13420);
nand U19922 (N_19922,N_16475,N_16110);
or U19923 (N_19923,N_15694,N_14793);
and U19924 (N_19924,N_14354,N_15078);
and U19925 (N_19925,N_13035,N_14331);
or U19926 (N_19926,N_13167,N_15331);
or U19927 (N_19927,N_15447,N_16165);
xnor U19928 (N_19928,N_13939,N_16174);
xor U19929 (N_19929,N_16918,N_12355);
and U19930 (N_19930,N_13004,N_15173);
nand U19931 (N_19931,N_17272,N_16419);
nand U19932 (N_19932,N_14625,N_14438);
and U19933 (N_19933,N_17558,N_14855);
nand U19934 (N_19934,N_17560,N_17328);
nor U19935 (N_19935,N_16468,N_15735);
and U19936 (N_19936,N_17492,N_16610);
xnor U19937 (N_19937,N_16266,N_14444);
and U19938 (N_19938,N_13238,N_12983);
nand U19939 (N_19939,N_17909,N_16544);
or U19940 (N_19940,N_17561,N_13847);
and U19941 (N_19941,N_14118,N_14642);
or U19942 (N_19942,N_17243,N_15654);
or U19943 (N_19943,N_13677,N_12354);
and U19944 (N_19944,N_12416,N_17076);
and U19945 (N_19945,N_16987,N_17293);
nor U19946 (N_19946,N_14588,N_14858);
nand U19947 (N_19947,N_14434,N_17078);
nor U19948 (N_19948,N_16416,N_17385);
nor U19949 (N_19949,N_13351,N_12317);
nor U19950 (N_19950,N_17727,N_15148);
nor U19951 (N_19951,N_14358,N_13230);
and U19952 (N_19952,N_12164,N_16166);
nand U19953 (N_19953,N_15591,N_14913);
or U19954 (N_19954,N_12346,N_13680);
nand U19955 (N_19955,N_13950,N_16904);
xor U19956 (N_19956,N_15853,N_15787);
nand U19957 (N_19957,N_17510,N_14729);
and U19958 (N_19958,N_13244,N_16179);
or U19959 (N_19959,N_14185,N_16171);
nand U19960 (N_19960,N_16096,N_14000);
nand U19961 (N_19961,N_12707,N_13916);
nor U19962 (N_19962,N_16381,N_15483);
nand U19963 (N_19963,N_15966,N_14137);
or U19964 (N_19964,N_13399,N_14067);
nor U19965 (N_19965,N_16512,N_15222);
or U19966 (N_19966,N_13867,N_17491);
nand U19967 (N_19967,N_17627,N_14246);
xor U19968 (N_19968,N_16118,N_17205);
nor U19969 (N_19969,N_16370,N_13356);
or U19970 (N_19970,N_13137,N_13931);
and U19971 (N_19971,N_15113,N_16450);
and U19972 (N_19972,N_12041,N_15313);
nand U19973 (N_19973,N_16920,N_14736);
and U19974 (N_19974,N_17638,N_17466);
nand U19975 (N_19975,N_15133,N_14088);
and U19976 (N_19976,N_14551,N_12252);
xnor U19977 (N_19977,N_12726,N_17680);
and U19978 (N_19978,N_13073,N_17520);
nand U19979 (N_19979,N_17941,N_15867);
or U19980 (N_19980,N_15621,N_17824);
or U19981 (N_19981,N_15566,N_14136);
nor U19982 (N_19982,N_15684,N_15700);
or U19983 (N_19983,N_16261,N_12139);
nand U19984 (N_19984,N_13812,N_14396);
and U19985 (N_19985,N_17032,N_15665);
xnor U19986 (N_19986,N_17327,N_16409);
xnor U19987 (N_19987,N_17803,N_17807);
nand U19988 (N_19988,N_17641,N_17517);
nor U19989 (N_19989,N_12967,N_16639);
and U19990 (N_19990,N_16854,N_14600);
nor U19991 (N_19991,N_12136,N_16434);
and U19992 (N_19992,N_16851,N_13043);
or U19993 (N_19993,N_14949,N_13547);
nand U19994 (N_19994,N_16344,N_15979);
and U19995 (N_19995,N_12230,N_15834);
nand U19996 (N_19996,N_15690,N_15695);
nor U19997 (N_19997,N_15578,N_17933);
or U19998 (N_19998,N_13725,N_13550);
xnor U19999 (N_19999,N_12064,N_13458);
or U20000 (N_20000,N_12172,N_16879);
xor U20001 (N_20001,N_12014,N_15379);
or U20002 (N_20002,N_12473,N_12081);
nand U20003 (N_20003,N_12303,N_17555);
nand U20004 (N_20004,N_12288,N_15278);
nor U20005 (N_20005,N_16076,N_13539);
xnor U20006 (N_20006,N_16304,N_14474);
and U20007 (N_20007,N_14607,N_16053);
nand U20008 (N_20008,N_13422,N_17740);
and U20009 (N_20009,N_13234,N_14359);
and U20010 (N_20010,N_17972,N_13727);
xnor U20011 (N_20011,N_12973,N_14692);
and U20012 (N_20012,N_17433,N_14512);
nand U20013 (N_20013,N_13966,N_14985);
xor U20014 (N_20014,N_12632,N_16538);
xor U20015 (N_20015,N_17834,N_14371);
xnor U20016 (N_20016,N_16246,N_17183);
xnor U20017 (N_20017,N_14053,N_13435);
nand U20018 (N_20018,N_16827,N_13751);
and U20019 (N_20019,N_16269,N_16676);
xor U20020 (N_20020,N_13463,N_15709);
nand U20021 (N_20021,N_16509,N_13674);
or U20022 (N_20022,N_16152,N_15481);
xnor U20023 (N_20023,N_17380,N_14872);
and U20024 (N_20024,N_12366,N_12285);
or U20025 (N_20025,N_12084,N_13398);
nor U20026 (N_20026,N_13828,N_16697);
xnor U20027 (N_20027,N_16286,N_13903);
or U20028 (N_20028,N_14869,N_12329);
xor U20029 (N_20029,N_15227,N_13280);
nand U20030 (N_20030,N_13638,N_17473);
xnor U20031 (N_20031,N_13114,N_16794);
nand U20032 (N_20032,N_12982,N_16874);
or U20033 (N_20033,N_14122,N_14236);
and U20034 (N_20034,N_14192,N_17024);
and U20035 (N_20035,N_14202,N_13794);
or U20036 (N_20036,N_12810,N_16939);
nor U20037 (N_20037,N_13354,N_12535);
and U20038 (N_20038,N_17844,N_17709);
xnor U20039 (N_20039,N_15022,N_13178);
nand U20040 (N_20040,N_14060,N_16734);
or U20041 (N_20041,N_17983,N_16385);
and U20042 (N_20042,N_13487,N_14504);
nand U20043 (N_20043,N_14126,N_15437);
and U20044 (N_20044,N_15821,N_15509);
and U20045 (N_20045,N_14079,N_16845);
or U20046 (N_20046,N_13275,N_12249);
and U20047 (N_20047,N_14050,N_15874);
nor U20048 (N_20048,N_15691,N_13333);
or U20049 (N_20049,N_12861,N_14921);
nor U20050 (N_20050,N_12330,N_17973);
xnor U20051 (N_20051,N_13877,N_17378);
nand U20052 (N_20052,N_16159,N_16515);
or U20053 (N_20053,N_17892,N_17731);
nand U20054 (N_20054,N_15831,N_16664);
and U20055 (N_20055,N_16926,N_14129);
nor U20056 (N_20056,N_17287,N_16367);
nor U20057 (N_20057,N_16341,N_17694);
or U20058 (N_20058,N_17676,N_13899);
xnor U20059 (N_20059,N_13994,N_15266);
nor U20060 (N_20060,N_15246,N_17394);
and U20061 (N_20061,N_13954,N_12262);
and U20062 (N_20062,N_14721,N_17625);
nor U20063 (N_20063,N_16663,N_14323);
nand U20064 (N_20064,N_14911,N_17199);
xor U20065 (N_20065,N_15404,N_17863);
or U20066 (N_20066,N_16969,N_12222);
xnor U20067 (N_20067,N_17391,N_17252);
or U20068 (N_20068,N_16605,N_16568);
xnor U20069 (N_20069,N_13318,N_13404);
xnor U20070 (N_20070,N_17811,N_17120);
nor U20071 (N_20071,N_12835,N_17518);
nand U20072 (N_20072,N_13290,N_14635);
nor U20073 (N_20073,N_17268,N_13612);
xor U20074 (N_20074,N_14907,N_15124);
nor U20075 (N_20075,N_13116,N_16769);
or U20076 (N_20076,N_13481,N_12192);
or U20077 (N_20077,N_12438,N_15277);
xor U20078 (N_20078,N_14488,N_15921);
and U20079 (N_20079,N_12622,N_16694);
and U20080 (N_20080,N_13762,N_13698);
xnor U20081 (N_20081,N_13791,N_14737);
nor U20082 (N_20082,N_17678,N_13117);
nand U20083 (N_20083,N_13032,N_13542);
nor U20084 (N_20084,N_13740,N_13173);
xnor U20085 (N_20085,N_17182,N_14753);
nor U20086 (N_20086,N_13716,N_17697);
nor U20087 (N_20087,N_13465,N_17247);
xnor U20088 (N_20088,N_14061,N_14701);
or U20089 (N_20089,N_13641,N_16176);
nand U20090 (N_20090,N_15176,N_15151);
xor U20091 (N_20091,N_17932,N_17577);
nand U20092 (N_20092,N_14695,N_14868);
or U20093 (N_20093,N_13584,N_13917);
and U20094 (N_20094,N_12491,N_17262);
or U20095 (N_20095,N_17849,N_17885);
xor U20096 (N_20096,N_14541,N_15417);
xor U20097 (N_20097,N_15480,N_14231);
nor U20098 (N_20098,N_12263,N_14732);
nand U20099 (N_20099,N_15104,N_14039);
nand U20100 (N_20100,N_13108,N_12485);
and U20101 (N_20101,N_13971,N_13317);
or U20102 (N_20102,N_12061,N_12388);
nor U20103 (N_20103,N_15294,N_16767);
xnor U20104 (N_20104,N_15043,N_16158);
and U20105 (N_20105,N_12208,N_16607);
nor U20106 (N_20106,N_15590,N_16405);
or U20107 (N_20107,N_16042,N_16786);
xnor U20108 (N_20108,N_17815,N_16913);
xnor U20109 (N_20109,N_12790,N_14622);
and U20110 (N_20110,N_16431,N_14819);
nor U20111 (N_20111,N_15249,N_13743);
nand U20112 (N_20112,N_16723,N_12202);
xnor U20113 (N_20113,N_14556,N_12209);
xnor U20114 (N_20114,N_13171,N_16458);
xnor U20115 (N_20115,N_12063,N_17251);
and U20116 (N_20116,N_15141,N_14389);
xor U20117 (N_20117,N_15944,N_13493);
nand U20118 (N_20118,N_14520,N_13921);
xnor U20119 (N_20119,N_17261,N_15840);
and U20120 (N_20120,N_12115,N_15851);
nor U20121 (N_20121,N_12089,N_17213);
nor U20122 (N_20122,N_14397,N_15763);
or U20123 (N_20123,N_15213,N_17329);
xnor U20124 (N_20124,N_12241,N_13831);
xor U20125 (N_20125,N_15015,N_12494);
nor U20126 (N_20126,N_12450,N_16301);
xnor U20127 (N_20127,N_13923,N_16083);
nor U20128 (N_20128,N_17027,N_15171);
and U20129 (N_20129,N_13953,N_16001);
nor U20130 (N_20130,N_14144,N_13019);
nand U20131 (N_20131,N_17943,N_15995);
and U20132 (N_20132,N_16461,N_15368);
nand U20133 (N_20133,N_12946,N_13293);
and U20134 (N_20134,N_14076,N_14559);
and U20135 (N_20135,N_15754,N_12784);
or U20136 (N_20136,N_14454,N_13629);
or U20137 (N_20137,N_13842,N_13396);
or U20138 (N_20138,N_15978,N_14519);
and U20139 (N_20139,N_14816,N_15032);
and U20140 (N_20140,N_15021,N_16524);
nor U20141 (N_20141,N_17224,N_16711);
nor U20142 (N_20142,N_14767,N_16482);
nor U20143 (N_20143,N_13268,N_15872);
and U20144 (N_20144,N_13343,N_17721);
xor U20145 (N_20145,N_13710,N_14648);
nor U20146 (N_20146,N_12567,N_14051);
and U20147 (N_20147,N_17623,N_12844);
nor U20148 (N_20148,N_15092,N_17732);
nor U20149 (N_20149,N_17389,N_14862);
and U20150 (N_20150,N_14605,N_14101);
xor U20151 (N_20151,N_13943,N_13734);
xor U20152 (N_20152,N_12213,N_17153);
or U20153 (N_20153,N_12634,N_14580);
and U20154 (N_20154,N_16345,N_13559);
nand U20155 (N_20155,N_12235,N_13962);
or U20156 (N_20156,N_13063,N_15971);
xor U20157 (N_20157,N_15734,N_17553);
xnor U20158 (N_20158,N_13838,N_15045);
or U20159 (N_20159,N_15737,N_15805);
nor U20160 (N_20160,N_16066,N_16430);
nand U20161 (N_20161,N_17381,N_12725);
nand U20162 (N_20162,N_15510,N_17303);
nand U20163 (N_20163,N_15365,N_15705);
nor U20164 (N_20164,N_15010,N_17802);
or U20165 (N_20165,N_13369,N_13410);
and U20166 (N_20166,N_15256,N_16132);
nor U20167 (N_20167,N_16530,N_12746);
nor U20168 (N_20168,N_17540,N_17699);
xnor U20169 (N_20169,N_16186,N_17052);
or U20170 (N_20170,N_14877,N_17804);
or U20171 (N_20171,N_14670,N_12980);
xnor U20172 (N_20172,N_15546,N_13220);
xnor U20173 (N_20173,N_14647,N_14123);
or U20174 (N_20174,N_16193,N_17571);
xor U20175 (N_20175,N_15046,N_17597);
nand U20176 (N_20176,N_17196,N_17000);
and U20177 (N_20177,N_13893,N_15401);
xnor U20178 (N_20178,N_16762,N_14306);
nand U20179 (N_20179,N_17472,N_17011);
and U20180 (N_20180,N_16417,N_15732);
or U20181 (N_20181,N_15125,N_14980);
or U20182 (N_20182,N_16307,N_17114);
nor U20183 (N_20183,N_13157,N_12648);
and U20184 (N_20184,N_15635,N_13028);
xor U20185 (N_20185,N_12393,N_15871);
nand U20186 (N_20186,N_12805,N_16443);
or U20187 (N_20187,N_12201,N_14353);
and U20188 (N_20188,N_15445,N_14916);
nor U20189 (N_20189,N_16895,N_12347);
nor U20190 (N_20190,N_14042,N_17068);
or U20191 (N_20191,N_13401,N_12149);
nor U20192 (N_20192,N_15676,N_15449);
nand U20193 (N_20193,N_15291,N_15759);
xor U20194 (N_20194,N_17726,N_15628);
and U20195 (N_20195,N_16508,N_13703);
xor U20196 (N_20196,N_15060,N_17368);
or U20197 (N_20197,N_16078,N_16107);
and U20198 (N_20198,N_17461,N_13500);
or U20199 (N_20199,N_17836,N_14244);
xnor U20200 (N_20200,N_13432,N_14470);
and U20201 (N_20201,N_17915,N_13022);
nand U20202 (N_20202,N_12533,N_13377);
and U20203 (N_20203,N_13908,N_16615);
nor U20204 (N_20204,N_13109,N_13430);
nor U20205 (N_20205,N_15055,N_17644);
xor U20206 (N_20206,N_16284,N_12184);
nor U20207 (N_20207,N_15526,N_14374);
nand U20208 (N_20208,N_15487,N_17703);
nand U20209 (N_20209,N_12881,N_12091);
or U20210 (N_20210,N_15531,N_15560);
nor U20211 (N_20211,N_13972,N_12817);
or U20212 (N_20212,N_12162,N_14197);
xor U20213 (N_20213,N_13787,N_15260);
nand U20214 (N_20214,N_13706,N_14342);
xnor U20215 (N_20215,N_12429,N_14379);
xnor U20216 (N_20216,N_12735,N_14938);
xnor U20217 (N_20217,N_17675,N_14071);
nor U20218 (N_20218,N_12988,N_15785);
and U20219 (N_20219,N_12432,N_13419);
or U20220 (N_20220,N_13845,N_15158);
and U20221 (N_20221,N_13081,N_13587);
xnor U20222 (N_20222,N_12522,N_17673);
nand U20223 (N_20223,N_13616,N_14787);
and U20224 (N_20224,N_12333,N_15378);
and U20225 (N_20225,N_13080,N_15466);
or U20226 (N_20226,N_16452,N_15146);
and U20227 (N_20227,N_12137,N_12898);
nor U20228 (N_20228,N_12669,N_15422);
nor U20229 (N_20229,N_17031,N_12255);
nor U20230 (N_20230,N_16657,N_13183);
or U20231 (N_20231,N_13514,N_12950);
xor U20232 (N_20232,N_16569,N_16305);
or U20233 (N_20233,N_15341,N_13066);
nand U20234 (N_20234,N_13150,N_13593);
nand U20235 (N_20235,N_12579,N_14251);
nor U20236 (N_20236,N_16681,N_15723);
or U20237 (N_20237,N_16817,N_13654);
nand U20238 (N_20238,N_16622,N_17401);
and U20239 (N_20239,N_13294,N_12447);
or U20240 (N_20240,N_16940,N_12461);
nor U20241 (N_20241,N_15477,N_16679);
nand U20242 (N_20242,N_14309,N_13374);
and U20243 (N_20243,N_16706,N_17939);
xnor U20244 (N_20244,N_15517,N_17898);
or U20245 (N_20245,N_14452,N_17003);
nand U20246 (N_20246,N_14501,N_13110);
nor U20247 (N_20247,N_14127,N_13198);
xor U20248 (N_20248,N_16627,N_12846);
and U20249 (N_20249,N_16789,N_14725);
nand U20250 (N_20250,N_14361,N_17033);
nor U20251 (N_20251,N_14759,N_16177);
and U20252 (N_20252,N_12062,N_17351);
nor U20253 (N_20253,N_13405,N_14738);
and U20254 (N_20254,N_16652,N_16454);
nor U20255 (N_20255,N_14575,N_15156);
nand U20256 (N_20256,N_14237,N_12464);
xnor U20257 (N_20257,N_17108,N_15407);
nand U20258 (N_20258,N_17421,N_12377);
xnor U20259 (N_20259,N_13668,N_13952);
nand U20260 (N_20260,N_14047,N_17590);
or U20261 (N_20261,N_13523,N_12254);
nor U20262 (N_20262,N_15752,N_15024);
nor U20263 (N_20263,N_12948,N_12189);
nor U20264 (N_20264,N_15533,N_16275);
nor U20265 (N_20265,N_12304,N_17105);
xnor U20266 (N_20266,N_15334,N_13888);
nand U20267 (N_20267,N_13750,N_17282);
and U20268 (N_20268,N_14254,N_17089);
or U20269 (N_20269,N_12758,N_12516);
or U20270 (N_20270,N_13636,N_14657);
or U20271 (N_20271,N_14683,N_13387);
or U20272 (N_20272,N_16014,N_17976);
or U20273 (N_20273,N_13357,N_17296);
nand U20274 (N_20274,N_16811,N_13287);
or U20275 (N_20275,N_17992,N_17903);
nand U20276 (N_20276,N_17248,N_12608);
or U20277 (N_20277,N_16109,N_12308);
nor U20278 (N_20278,N_14771,N_13122);
xnor U20279 (N_20279,N_16485,N_12019);
nor U20280 (N_20280,N_16887,N_15632);
nor U20281 (N_20281,N_14991,N_14615);
and U20282 (N_20282,N_16655,N_14560);
and U20283 (N_20283,N_16153,N_14068);
xor U20284 (N_20284,N_16389,N_13319);
nand U20285 (N_20285,N_16262,N_15689);
nor U20286 (N_20286,N_16120,N_16222);
nand U20287 (N_20287,N_17799,N_12603);
xnor U20288 (N_20288,N_13452,N_16962);
and U20289 (N_20289,N_14936,N_16207);
and U20290 (N_20290,N_17396,N_12000);
or U20291 (N_20291,N_12224,N_12448);
and U20292 (N_20292,N_15530,N_15622);
xor U20293 (N_20293,N_17292,N_12873);
nor U20294 (N_20294,N_16914,N_16637);
xnor U20295 (N_20295,N_17062,N_13999);
nor U20296 (N_20296,N_13483,N_12653);
and U20297 (N_20297,N_16980,N_13442);
xor U20298 (N_20298,N_14156,N_15118);
nand U20299 (N_20299,N_14209,N_15841);
and U20300 (N_20300,N_16378,N_12215);
nand U20301 (N_20301,N_14009,N_16644);
and U20302 (N_20302,N_14969,N_15184);
nor U20303 (N_20303,N_12383,N_17047);
and U20304 (N_20304,N_16106,N_15273);
or U20305 (N_20305,N_16946,N_17985);
or U20306 (N_20306,N_17672,N_17405);
nand U20307 (N_20307,N_12616,N_15662);
xor U20308 (N_20308,N_13748,N_15269);
or U20309 (N_20309,N_13016,N_15868);
and U20310 (N_20310,N_13901,N_13600);
nor U20311 (N_20311,N_12133,N_14411);
nor U20312 (N_20312,N_15236,N_14006);
nor U20313 (N_20313,N_14895,N_17346);
or U20314 (N_20314,N_17599,N_16148);
nor U20315 (N_20315,N_12318,N_13321);
nand U20316 (N_20316,N_13738,N_17544);
nor U20317 (N_20317,N_16902,N_17587);
nand U20318 (N_20318,N_12643,N_16810);
nand U20319 (N_20319,N_12405,N_17914);
nor U20320 (N_20320,N_14035,N_13737);
and U20321 (N_20321,N_14772,N_15041);
or U20322 (N_20322,N_15383,N_14467);
nor U20323 (N_20323,N_13482,N_17578);
or U20324 (N_20324,N_12794,N_17842);
or U20325 (N_20325,N_14684,N_12678);
xnor U20326 (N_20326,N_12558,N_14267);
nor U20327 (N_20327,N_17653,N_17141);
xor U20328 (N_20328,N_13651,N_17942);
nand U20329 (N_20329,N_13792,N_17953);
or U20330 (N_20330,N_12981,N_12965);
and U20331 (N_20331,N_15937,N_17720);
or U20332 (N_20332,N_16048,N_16606);
nand U20333 (N_20333,N_14032,N_17185);
and U20334 (N_20334,N_16215,N_15610);
or U20335 (N_20335,N_12680,N_12924);
or U20336 (N_20336,N_16768,N_12170);
or U20337 (N_20337,N_15660,N_15467);
and U20338 (N_20338,N_15335,N_12949);
nand U20339 (N_20339,N_12103,N_14093);
nand U20340 (N_20340,N_14941,N_13859);
or U20341 (N_20341,N_13235,N_14784);
nand U20342 (N_20342,N_17004,N_13646);
nand U20343 (N_20343,N_17509,N_17030);
nand U20344 (N_20344,N_14894,N_12572);
nand U20345 (N_20345,N_16062,N_13508);
nor U20346 (N_20346,N_14521,N_17483);
nand U20347 (N_20347,N_14108,N_15002);
nand U20348 (N_20348,N_14675,N_16661);
or U20349 (N_20349,N_14255,N_17870);
or U20350 (N_20350,N_12384,N_17574);
and U20351 (N_20351,N_14585,N_13835);
or U20352 (N_20352,N_15715,N_17632);
or U20353 (N_20353,N_15253,N_15708);
xor U20354 (N_20354,N_16656,N_13635);
and U20355 (N_20355,N_15109,N_14544);
nand U20356 (N_20356,N_12020,N_13746);
and U20357 (N_20357,N_17186,N_12143);
nand U20358 (N_20358,N_15501,N_17937);
or U20359 (N_20359,N_14134,N_16550);
nor U20360 (N_20360,N_15943,N_17890);
xor U20361 (N_20361,N_14994,N_16008);
nor U20362 (N_20362,N_14238,N_17005);
xor U20363 (N_20363,N_14699,N_13279);
xnor U20364 (N_20364,N_16459,N_16830);
xor U20365 (N_20365,N_15802,N_17747);
and U20366 (N_20366,N_14631,N_16278);
and U20367 (N_20367,N_16814,N_12148);
nand U20368 (N_20368,N_14540,N_12618);
nand U20369 (N_20369,N_13033,N_17468);
and U20370 (N_20370,N_13469,N_12501);
and U20371 (N_20371,N_12942,N_14780);
xnor U20372 (N_20372,N_17534,N_14776);
nand U20373 (N_20373,N_13885,N_12842);
xor U20374 (N_20374,N_15830,N_17835);
nor U20375 (N_20375,N_12058,N_16259);
or U20376 (N_20376,N_16388,N_16317);
xnor U20377 (N_20377,N_17949,N_13519);
xor U20378 (N_20378,N_13076,N_16330);
xor U20379 (N_20379,N_17278,N_15741);
nor U20380 (N_20380,N_15247,N_14221);
or U20381 (N_20381,N_16410,N_15898);
xor U20382 (N_20382,N_15406,N_13176);
nand U20383 (N_20383,N_16126,N_15340);
nand U20384 (N_20384,N_12884,N_14848);
nor U20385 (N_20385,N_13139,N_17977);
nor U20386 (N_20386,N_13689,N_14080);
nand U20387 (N_20387,N_16753,N_16113);
and U20388 (N_20388,N_15244,N_13358);
xor U20389 (N_20389,N_14954,N_17281);
nor U20390 (N_20390,N_17496,N_16517);
and U20391 (N_20391,N_16800,N_14850);
and U20392 (N_20392,N_13370,N_14493);
nor U20393 (N_20393,N_14673,N_12620);
and U20394 (N_20394,N_12056,N_14898);
and U20395 (N_20395,N_17354,N_17302);
nor U20396 (N_20396,N_16058,N_14298);
nor U20397 (N_20397,N_12830,N_15287);
nand U20398 (N_20398,N_12773,N_15154);
or U20399 (N_20399,N_17330,N_14731);
xor U20400 (N_20400,N_13197,N_14303);
xnor U20401 (N_20401,N_17400,N_17409);
nor U20402 (N_20402,N_13807,N_15101);
xor U20403 (N_20403,N_13156,N_13910);
nand U20404 (N_20404,N_15631,N_15181);
xor U20405 (N_20405,N_16256,N_13622);
xnor U20406 (N_20406,N_12436,N_14412);
and U20407 (N_20407,N_16359,N_14167);
nand U20408 (N_20408,N_15981,N_17899);
xor U20409 (N_20409,N_15457,N_14171);
and U20410 (N_20410,N_14964,N_12581);
nor U20411 (N_20411,N_14830,N_15351);
or U20412 (N_20412,N_14148,N_14733);
nor U20413 (N_20413,N_16101,N_12419);
and U20414 (N_20414,N_13263,N_17010);
nor U20415 (N_20415,N_14274,N_15147);
and U20416 (N_20416,N_15923,N_12521);
and U20417 (N_20417,N_13472,N_13417);
nand U20418 (N_20418,N_17666,N_12233);
and U20419 (N_20419,N_13776,N_16395);
nand U20420 (N_20420,N_16881,N_16864);
nand U20421 (N_20421,N_14419,N_17121);
or U20422 (N_20422,N_12236,N_17465);
xor U20423 (N_20423,N_13517,N_15878);
nand U20424 (N_20424,N_15135,N_13700);
or U20425 (N_20425,N_15350,N_14099);
nor U20426 (N_20426,N_17083,N_17805);
nor U20427 (N_20427,N_14407,N_12431);
and U20428 (N_20428,N_12269,N_15548);
and U20429 (N_20429,N_12639,N_16889);
xor U20430 (N_20430,N_12141,N_14316);
nor U20431 (N_20431,N_14375,N_15389);
nor U20432 (N_20432,N_12385,N_17291);
or U20433 (N_20433,N_15913,N_12693);
or U20434 (N_20434,N_13106,N_12787);
nor U20435 (N_20435,N_14336,N_13817);
xor U20436 (N_20436,N_12867,N_15838);
and U20437 (N_20437,N_15263,N_13222);
nand U20438 (N_20438,N_15028,N_12728);
xor U20439 (N_20439,N_16362,N_16519);
or U20440 (N_20440,N_15166,N_14637);
xor U20441 (N_20441,N_17996,N_14526);
nand U20442 (N_20442,N_15214,N_14392);
and U20443 (N_20443,N_13118,N_15767);
nor U20444 (N_20444,N_14757,N_13711);
nor U20445 (N_20445,N_15725,N_14367);
or U20446 (N_20446,N_13332,N_14074);
and U20447 (N_20447,N_13501,N_17707);
nor U20448 (N_20448,N_12406,N_12650);
or U20449 (N_20449,N_17013,N_12808);
nand U20450 (N_20450,N_14633,N_14804);
and U20451 (N_20451,N_15619,N_14558);
nand U20452 (N_20452,N_13648,N_14860);
or U20453 (N_20453,N_16061,N_14304);
nor U20454 (N_20454,N_12369,N_14618);
xnor U20455 (N_20455,N_16584,N_12633);
or U20456 (N_20456,N_16993,N_13628);
nor U20457 (N_20457,N_17586,N_14029);
and U20458 (N_20458,N_16692,N_16642);
nor U20459 (N_20459,N_17635,N_13837);
xor U20460 (N_20460,N_13062,N_16287);
nor U20461 (N_20461,N_17688,N_15190);
and U20462 (N_20462,N_13142,N_17478);
or U20463 (N_20463,N_12478,N_17572);
and U20464 (N_20464,N_12589,N_15282);
and U20465 (N_20465,N_14645,N_14740);
nor U20466 (N_20466,N_14958,N_15390);
or U20467 (N_20467,N_16069,N_16825);
xor U20468 (N_20468,N_12941,N_17238);
or U20469 (N_20469,N_15935,N_12845);
nand U20470 (N_20470,N_13927,N_16254);
xnor U20471 (N_20471,N_14586,N_14892);
xnor U20472 (N_20472,N_12654,N_13217);
and U20473 (N_20473,N_14813,N_14946);
nor U20474 (N_20474,N_13524,N_13111);
or U20475 (N_20475,N_12341,N_12964);
or U20476 (N_20476,N_14805,N_16134);
and U20477 (N_20477,N_15478,N_17920);
nor U20478 (N_20478,N_14902,N_17548);
and U20479 (N_20479,N_12011,N_16055);
xnor U20480 (N_20480,N_13415,N_12953);
nor U20481 (N_20481,N_12613,N_14680);
nor U20482 (N_20482,N_17532,N_17191);
nand U20483 (N_20483,N_17706,N_17851);
nand U20484 (N_20484,N_13857,N_15264);
nor U20485 (N_20485,N_17713,N_16537);
nand U20486 (N_20486,N_15065,N_15826);
nand U20487 (N_20487,N_13360,N_13870);
xnor U20488 (N_20488,N_15862,N_14287);
and U20489 (N_20489,N_16251,N_16047);
and U20490 (N_20490,N_14193,N_17818);
nand U20491 (N_20491,N_15672,N_16905);
nand U20492 (N_20492,N_17808,N_15308);
nor U20493 (N_20493,N_17918,N_16598);
or U20494 (N_20494,N_15270,N_16978);
xor U20495 (N_20495,N_15772,N_16489);
nor U20496 (N_20496,N_12210,N_15393);
xor U20497 (N_20497,N_14398,N_13391);
nor U20498 (N_20498,N_17861,N_12109);
and U20499 (N_20499,N_15455,N_15683);
xor U20500 (N_20500,N_17159,N_12752);
or U20501 (N_20501,N_16188,N_13297);
nor U20502 (N_20502,N_16994,N_17533);
nand U20503 (N_20503,N_13961,N_13632);
or U20504 (N_20504,N_13187,N_13595);
and U20505 (N_20505,N_12085,N_14754);
nor U20506 (N_20506,N_12340,N_15633);
nor U20507 (N_20507,N_13001,N_13573);
and U20508 (N_20508,N_16219,N_14915);
nand U20509 (N_20509,N_17314,N_12938);
and U20510 (N_20510,N_14065,N_13447);
xnor U20511 (N_20511,N_17524,N_16899);
and U20512 (N_20512,N_15602,N_17926);
nor U20513 (N_20513,N_12886,N_15702);
nand U20514 (N_20514,N_15884,N_14182);
and U20515 (N_20515,N_17006,N_12858);
nand U20516 (N_20516,N_16321,N_17436);
and U20517 (N_20517,N_14836,N_12987);
nand U20518 (N_20518,N_13779,N_16751);
or U20519 (N_20519,N_15063,N_12147);
and U20520 (N_20520,N_17338,N_15339);
nand U20521 (N_20521,N_15897,N_12826);
nor U20522 (N_20522,N_14175,N_17881);
nor U20523 (N_20523,N_14253,N_16722);
or U20524 (N_20524,N_17135,N_16050);
nor U20525 (N_20525,N_17273,N_14947);
nand U20526 (N_20526,N_12282,N_12278);
nand U20527 (N_20527,N_16562,N_14208);
nand U20528 (N_20528,N_13438,N_14489);
nor U20529 (N_20529,N_13704,N_13580);
and U20530 (N_20530,N_13444,N_12246);
and U20531 (N_20531,N_13640,N_15849);
xor U20532 (N_20532,N_12030,N_13262);
or U20533 (N_20533,N_16965,N_14092);
nand U20534 (N_20534,N_16247,N_16212);
nor U20535 (N_20535,N_14829,N_15925);
and U20536 (N_20536,N_14131,N_13480);
or U20537 (N_20537,N_15074,N_12644);
xor U20538 (N_20538,N_17050,N_12543);
xor U20539 (N_20539,N_15342,N_16666);
nor U20540 (N_20540,N_12717,N_13510);
or U20541 (N_20541,N_12358,N_16577);
nor U20542 (N_20542,N_16100,N_12868);
xor U20543 (N_20543,N_16342,N_16401);
or U20544 (N_20544,N_15066,N_12344);
or U20545 (N_20545,N_12403,N_13997);
xnor U20546 (N_20546,N_14203,N_15842);
and U20547 (N_20547,N_14587,N_17174);
nand U20548 (N_20548,N_17710,N_15786);
and U20549 (N_20549,N_12513,N_12173);
nand U20550 (N_20550,N_13936,N_12291);
or U20551 (N_20551,N_16335,N_14420);
nor U20552 (N_20552,N_14910,N_13981);
xnor U20553 (N_20553,N_12696,N_12991);
xor U20554 (N_20554,N_12944,N_12523);
nand U20555 (N_20555,N_13300,N_14241);
or U20556 (N_20556,N_14168,N_12800);
or U20557 (N_20557,N_15804,N_16715);
xor U20558 (N_20558,N_13044,N_14328);
xnor U20559 (N_20559,N_14376,N_17319);
and U20560 (N_20560,N_16332,N_16674);
xnor U20561 (N_20561,N_17543,N_12299);
nand U20562 (N_20562,N_16624,N_17770);
and U20563 (N_20563,N_12598,N_17283);
nor U20564 (N_20564,N_14890,N_17654);
and U20565 (N_20565,N_17097,N_12742);
or U20566 (N_20566,N_16997,N_14021);
xor U20567 (N_20567,N_17991,N_13206);
nand U20568 (N_20568,N_16526,N_16289);
or U20569 (N_20569,N_15620,N_17166);
and U20570 (N_20570,N_15150,N_16472);
nor U20571 (N_20571,N_14481,N_15366);
or U20572 (N_20572,N_15657,N_13147);
nor U20573 (N_20573,N_13513,N_14325);
xnor U20574 (N_20574,N_14777,N_15706);
or U20575 (N_20575,N_12906,N_14639);
nor U20576 (N_20576,N_15505,N_17573);
xor U20577 (N_20577,N_16932,N_16396);
nand U20578 (N_20578,N_12445,N_16479);
xor U20579 (N_20579,N_13897,N_12893);
nor U20580 (N_20580,N_15495,N_14437);
xor U20581 (N_20581,N_15367,N_12458);
xnor U20582 (N_20582,N_17002,N_12274);
nand U20583 (N_20583,N_12509,N_17148);
xor U20584 (N_20584,N_14844,N_17753);
nor U20585 (N_20585,N_13713,N_13586);
and U20586 (N_20586,N_12376,N_16578);
nand U20587 (N_20587,N_15910,N_13301);
and U20588 (N_20588,N_12657,N_12049);
and U20589 (N_20589,N_17498,N_12750);
or U20590 (N_20590,N_17730,N_12469);
and U20591 (N_20591,N_16282,N_13042);
or U20592 (N_20592,N_16699,N_12349);
and U20593 (N_20593,N_13528,N_12847);
and U20594 (N_20594,N_12930,N_12888);
nor U20595 (N_20595,N_13941,N_15370);
nand U20596 (N_20596,N_12342,N_14350);
and U20597 (N_20597,N_16309,N_16973);
nor U20598 (N_20598,N_14096,N_14482);
and U20599 (N_20599,N_12803,N_15426);
and U20600 (N_20600,N_16314,N_16999);
or U20601 (N_20601,N_15254,N_15303);
nor U20602 (N_20602,N_13303,N_16470);
and U20603 (N_20603,N_16792,N_12018);
nor U20604 (N_20604,N_13439,N_16209);
nand U20605 (N_20605,N_16559,N_13673);
xor U20606 (N_20606,N_13457,N_16547);
nand U20607 (N_20607,N_13014,N_13865);
or U20608 (N_20608,N_12038,N_14533);
nand U20609 (N_20609,N_15198,N_15170);
and U20610 (N_20610,N_13900,N_13361);
nor U20611 (N_20611,N_17322,N_12435);
or U20612 (N_20612,N_16233,N_13735);
nor U20613 (N_20613,N_14305,N_12731);
and U20614 (N_20614,N_16931,N_14125);
or U20615 (N_20615,N_14710,N_16085);
nor U20616 (N_20616,N_16487,N_15499);
and U20617 (N_20617,N_14952,N_15210);
xor U20618 (N_20618,N_16842,N_16391);
and U20619 (N_20619,N_13454,N_15353);
nand U20620 (N_20620,N_16821,N_13266);
or U20621 (N_20621,N_15136,N_13090);
nand U20622 (N_20622,N_13889,N_15886);
xnor U20623 (N_20623,N_12520,N_14966);
nor U20624 (N_20624,N_14744,N_17923);
nor U20625 (N_20625,N_12894,N_14524);
nor U20626 (N_20626,N_15271,N_12367);
and U20627 (N_20627,N_14041,N_15048);
xnor U20628 (N_20628,N_14294,N_13987);
nor U20629 (N_20629,N_12160,N_17798);
nor U20630 (N_20630,N_17502,N_14879);
xnor U20631 (N_20631,N_17225,N_12954);
nand U20632 (N_20632,N_13258,N_14372);
and U20633 (N_20633,N_17963,N_16255);
or U20634 (N_20634,N_16064,N_14082);
or U20635 (N_20635,N_12120,N_13453);
nor U20636 (N_20636,N_12193,N_15369);
nor U20637 (N_20637,N_15947,N_14181);
and U20638 (N_20638,N_13416,N_14486);
xor U20639 (N_20639,N_15866,N_12188);
or U20640 (N_20640,N_17402,N_13532);
nand U20641 (N_20641,N_17617,N_15770);
or U20642 (N_20642,N_16130,N_16890);
xnor U20643 (N_20643,N_16588,N_14430);
nand U20644 (N_20644,N_16684,N_13937);
xor U20645 (N_20645,N_14120,N_13554);
nand U20646 (N_20646,N_13813,N_16696);
and U20647 (N_20647,N_15861,N_17876);
nand U20648 (N_20648,N_17643,N_14381);
nor U20649 (N_20649,N_16095,N_15077);
nor U20650 (N_20650,N_17615,N_15129);
nor U20651 (N_20651,N_17312,N_14425);
nor U20652 (N_20652,N_15688,N_15304);
xor U20653 (N_20653,N_16226,N_17545);
xnor U20654 (N_20654,N_16539,N_15781);
nand U20655 (N_20655,N_14166,N_17331);
and U20656 (N_20656,N_16218,N_15847);
nand U20657 (N_20657,N_16268,N_12834);
or U20658 (N_20658,N_17749,N_13774);
and U20659 (N_20659,N_14459,N_16804);
xor U20660 (N_20660,N_14018,N_12396);
or U20661 (N_20661,N_14713,N_12083);
nor U20662 (N_20662,N_16514,N_14451);
or U20663 (N_20663,N_12191,N_16669);
and U20664 (N_20664,N_16243,N_17634);
and U20665 (N_20665,N_16471,N_17994);
nor U20666 (N_20666,N_12576,N_17695);
xnor U20667 (N_20667,N_15262,N_14628);
xnor U20668 (N_20668,N_12925,N_16805);
and U20669 (N_20669,N_15997,N_13777);
nor U20670 (N_20670,N_12623,N_14090);
nor U20671 (N_20671,N_16869,N_12194);
and U20672 (N_20672,N_15089,N_12840);
nand U20673 (N_20673,N_16868,N_16822);
and U20674 (N_20674,N_13342,N_16828);
nor U20675 (N_20675,N_17438,N_12119);
or U20676 (N_20676,N_14334,N_14380);
xor U20677 (N_20677,N_12900,N_15230);
and U20678 (N_20678,N_14062,N_15356);
xnor U20679 (N_20679,N_17280,N_15778);
or U20680 (N_20680,N_12931,N_14841);
xor U20681 (N_20681,N_13143,N_16467);
nand U20682 (N_20682,N_12498,N_12865);
and U20683 (N_20683,N_17603,N_14960);
nor U20684 (N_20684,N_15982,N_15882);
or U20685 (N_20685,N_12975,N_17662);
nor U20686 (N_20686,N_13242,N_14347);
or U20687 (N_20687,N_14758,N_13516);
xor U20688 (N_20688,N_12923,N_16326);
xor U20689 (N_20689,N_15372,N_17922);
and U20690 (N_20690,N_14256,N_16628);
or U20691 (N_20691,N_17789,N_16260);
nand U20692 (N_20692,N_16071,N_17414);
nand U20693 (N_20693,N_14565,N_12459);
nand U20694 (N_20694,N_13909,N_17308);
or U20695 (N_20695,N_12716,N_15663);
and U20696 (N_20696,N_16311,N_16826);
nor U20697 (N_20697,N_15145,N_17769);
and U20698 (N_20698,N_14576,N_14609);
and U20699 (N_20699,N_14825,N_17831);
nor U20700 (N_20700,N_13490,N_12747);
nor U20701 (N_20701,N_15634,N_12685);
xor U20702 (N_20702,N_17754,N_12480);
and U20703 (N_20703,N_15152,N_17474);
nand U20704 (N_20704,N_13010,N_12426);
xor U20705 (N_20705,N_15013,N_16192);
xor U20706 (N_20706,N_13557,N_12398);
xor U20707 (N_20707,N_13248,N_16005);
and U20708 (N_20708,N_16936,N_12655);
or U20709 (N_20709,N_13474,N_16731);
and U20710 (N_20710,N_16032,N_17882);
nor U20711 (N_20711,N_17305,N_13055);
and U20712 (N_20712,N_14109,N_15859);
or U20713 (N_20713,N_13685,N_12295);
nor U20714 (N_20714,N_12400,N_17810);
nand U20715 (N_20715,N_15641,N_15307);
xnor U20716 (N_20716,N_14745,N_13284);
and U20717 (N_20717,N_13191,N_17079);
and U20718 (N_20718,N_12219,N_15237);
nor U20719 (N_20719,N_12969,N_15774);
and U20720 (N_20720,N_15792,N_13054);
nand U20721 (N_20721,N_12511,N_17057);
nand U20722 (N_20722,N_14073,N_16035);
and U20723 (N_20723,N_16797,N_13569);
and U20724 (N_20724,N_13553,N_15017);
nor U20725 (N_20725,N_16387,N_17095);
nor U20726 (N_20726,N_17748,N_12424);
nor U20727 (N_20727,N_14387,N_13282);
and U20728 (N_20728,N_12313,N_16232);
nand U20729 (N_20729,N_12203,N_12825);
and U20730 (N_20730,N_17858,N_16680);
or U20731 (N_20731,N_14081,N_15788);
or U20732 (N_20732,N_13759,N_13956);
nand U20733 (N_20733,N_14930,N_14457);
nor U20734 (N_20734,N_12474,N_13878);
xnor U20735 (N_20735,N_17456,N_13731);
or U20736 (N_20736,N_16224,N_16818);
nand U20737 (N_20737,N_14768,N_16348);
or U20738 (N_20738,N_14795,N_15521);
nand U20739 (N_20739,N_17925,N_13433);
or U20740 (N_20740,N_17090,N_13902);
or U20741 (N_20741,N_16382,N_12339);
or U20742 (N_20742,N_17152,N_14686);
and U20743 (N_20743,N_12010,N_17099);
and U20744 (N_20744,N_16548,N_17467);
nor U20745 (N_20745,N_15461,N_15488);
xnor U20746 (N_20746,N_16952,N_15926);
or U20747 (N_20747,N_16820,N_16777);
xnor U20748 (N_20748,N_17629,N_17606);
or U20749 (N_20749,N_17222,N_16300);
xor U20750 (N_20750,N_14832,N_14224);
xnor U20751 (N_20751,N_13170,N_16557);
or U20752 (N_20752,N_14054,N_16170);
nor U20753 (N_20753,N_16372,N_12668);
xor U20754 (N_20754,N_17722,N_16727);
nand U20755 (N_20755,N_12882,N_13246);
xnor U20756 (N_20756,N_17940,N_14031);
nor U20757 (N_20757,N_14248,N_16964);
and U20758 (N_20758,N_15964,N_15507);
nor U20759 (N_20759,N_17767,N_15519);
nand U20760 (N_20760,N_12560,N_16746);
nor U20761 (N_20761,N_15396,N_17756);
nor U20762 (N_20762,N_12496,N_12531);
xor U20763 (N_20763,N_17304,N_15954);
xnor U20764 (N_20764,N_17059,N_12550);
nand U20765 (N_20765,N_17927,N_15275);
or U20766 (N_20766,N_13212,N_17315);
and U20767 (N_20767,N_15491,N_17439);
and U20768 (N_20768,N_17674,N_15753);
or U20769 (N_20769,N_16960,N_13296);
nand U20770 (N_20770,N_14259,N_12232);
nand U20771 (N_20771,N_17537,N_16704);
or U20772 (N_20772,N_15265,N_14592);
and U20773 (N_20773,N_13618,N_15855);
nand U20774 (N_20774,N_16011,N_16916);
or U20775 (N_20775,N_14213,N_16494);
xor U20776 (N_20776,N_13132,N_12050);
xor U20777 (N_20777,N_17374,N_13202);
or U20778 (N_20778,N_15977,N_14953);
or U20779 (N_20779,N_15482,N_12005);
xor U20780 (N_20780,N_12652,N_13400);
nand U20781 (N_20781,N_15355,N_14075);
nor U20782 (N_20782,N_12134,N_14914);
xor U20783 (N_20783,N_15502,N_14180);
or U20784 (N_20784,N_16364,N_16242);
and U20785 (N_20785,N_13478,N_12879);
xnor U20786 (N_20786,N_15391,N_16847);
or U20787 (N_20787,N_13182,N_13267);
xnor U20788 (N_20788,N_15701,N_13639);
and U20789 (N_20789,N_17256,N_16319);
and U20790 (N_20790,N_17020,N_17193);
or U20791 (N_20791,N_16358,N_16659);
nor U20792 (N_20792,N_13211,N_16893);
nand U20793 (N_20793,N_12588,N_15888);
xnor U20794 (N_20794,N_17795,N_12856);
nor U20795 (N_20795,N_17471,N_13488);
and U20796 (N_20796,N_14769,N_16570);
nor U20797 (N_20797,N_15290,N_13879);
nor U20798 (N_20798,N_13264,N_17124);
nand U20799 (N_20799,N_12483,N_17780);
and U20800 (N_20800,N_14676,N_14688);
nand U20801 (N_20801,N_17778,N_17733);
nand U20802 (N_20802,N_17919,N_13181);
or U20803 (N_20803,N_13098,N_15580);
and U20804 (N_20804,N_13712,N_15288);
xor U20805 (N_20805,N_17691,N_14477);
nor U20806 (N_20806,N_17200,N_13504);
or U20807 (N_20807,N_15323,N_16279);
nor U20808 (N_20808,N_14324,N_17738);
xor U20809 (N_20809,N_17946,N_15453);
nor U20810 (N_20810,N_14847,N_16832);
nor U20811 (N_20811,N_12759,N_17650);
and U20812 (N_20812,N_15328,N_14317);
nand U20813 (N_20813,N_17360,N_12053);
xnor U20814 (N_20814,N_12786,N_15848);
nand U20815 (N_20815,N_14269,N_12446);
xor U20816 (N_20816,N_16571,N_15592);
nor U20817 (N_20817,N_16629,N_13497);
and U20818 (N_20818,N_12538,N_12959);
nand U20819 (N_20819,N_12649,N_12972);
nor U20820 (N_20820,N_13085,N_14040);
nand U20821 (N_20821,N_17339,N_15062);
xor U20822 (N_20822,N_16763,N_14230);
nand U20823 (N_20823,N_15730,N_12681);
and U20824 (N_20824,N_14722,N_14005);
or U20825 (N_20825,N_16938,N_12642);
nand U20826 (N_20826,N_16593,N_12863);
and U20827 (N_20827,N_12677,N_12507);
and U20828 (N_20828,N_15344,N_16379);
nor U20829 (N_20829,N_12499,N_13530);
nor U20830 (N_20830,N_14835,N_16883);
xnor U20831 (N_20831,N_15299,N_15645);
and U20832 (N_20832,N_16986,N_13989);
nand U20833 (N_20833,N_16857,N_17232);
nor U20834 (N_20834,N_17452,N_14962);
xnor U20835 (N_20835,N_17482,N_15611);
xnor U20836 (N_20836,N_14513,N_12402);
nand U20837 (N_20837,N_14959,N_17241);
and U20838 (N_20838,N_13253,N_13380);
xnor U20839 (N_20839,N_15257,N_15596);
nor U20840 (N_20840,N_14327,N_15053);
or U20841 (N_20841,N_14939,N_12315);
nor U20842 (N_20842,N_13000,N_16783);
or U20843 (N_20843,N_12597,N_16437);
xor U20844 (N_20844,N_15674,N_15698);
and U20845 (N_20845,N_14233,N_12012);
nand U20846 (N_20846,N_15761,N_12636);
and U20847 (N_20847,N_14554,N_15993);
nand U20848 (N_20848,N_12760,N_13571);
xor U20849 (N_20849,N_14014,N_17060);
or U20850 (N_20850,N_12351,N_13271);
xnor U20851 (N_20851,N_17947,N_13538);
nor U20852 (N_20852,N_14273,N_15475);
nand U20853 (N_20853,N_15193,N_17395);
nor U20854 (N_20854,N_17639,N_12144);
xor U20855 (N_20855,N_16947,N_16503);
xor U20856 (N_20856,N_12223,N_12711);
nand U20857 (N_20857,N_14384,N_16928);
nor U20858 (N_20858,N_15410,N_17883);
or U20859 (N_20859,N_15485,N_12068);
xnor U20860 (N_20860,N_16439,N_16352);
and U20861 (N_20861,N_16740,N_14992);
and U20862 (N_20862,N_15209,N_17596);
and U20863 (N_20863,N_17233,N_17235);
or U20864 (N_20864,N_17567,N_12323);
xnor U20865 (N_20865,N_16718,N_15972);
nand U20866 (N_20866,N_15352,N_12156);
or U20867 (N_20867,N_12609,N_15780);
or U20868 (N_20868,N_14130,N_17311);
xnor U20869 (N_20869,N_12665,N_15122);
nor U20870 (N_20870,N_16500,N_14781);
or U20871 (N_20871,N_12945,N_16923);
xor U20872 (N_20872,N_16350,N_14446);
or U20873 (N_20873,N_13657,N_15728);
xnor U20874 (N_20874,N_13951,N_16831);
xor U20875 (N_20875,N_15216,N_12960);
nor U20876 (N_20876,N_12155,N_15996);
nor U20877 (N_20877,N_14846,N_14418);
nor U20878 (N_20878,N_15615,N_12337);
xor U20879 (N_20879,N_16901,N_12042);
xor U20880 (N_20880,N_12088,N_14400);
and U20881 (N_20881,N_16180,N_17630);
nand U20882 (N_20882,N_13389,N_14239);
or U20883 (N_20883,N_15799,N_17299);
xnor U20884 (N_20884,N_13858,N_12165);
and U20885 (N_20885,N_15245,N_13120);
and U20886 (N_20886,N_14490,N_17788);
and U20887 (N_20887,N_13274,N_16671);
and U20888 (N_20888,N_13124,N_16203);
and U20889 (N_20889,N_14818,N_14386);
xor U20890 (N_20890,N_17613,N_15811);
and U20891 (N_20891,N_15724,N_12664);
nand U20892 (N_20892,N_12910,N_13060);
or U20893 (N_20893,N_12326,N_17295);
nand U20894 (N_20894,N_14270,N_15432);
nor U20895 (N_20895,N_15463,N_12159);
and U20896 (N_20896,N_14242,N_16029);
xnor U20897 (N_20897,N_12659,N_16223);
xnor U20898 (N_20898,N_13856,N_15374);
and U20899 (N_20899,N_17896,N_16505);
nor U20900 (N_20900,N_13964,N_13240);
and U20901 (N_20901,N_12594,N_13581);
xnor U20902 (N_20902,N_16888,N_13394);
and U20903 (N_20903,N_12602,N_14022);
xor U20904 (N_20904,N_12412,N_15784);
and U20905 (N_20905,N_15573,N_14128);
xor U20906 (N_20906,N_16028,N_16549);
and U20907 (N_20907,N_12045,N_13884);
nor U20908 (N_20908,N_16985,N_15895);
nor U20909 (N_20909,N_14155,N_12992);
nor U20910 (N_20910,N_12593,N_12874);
xnor U20911 (N_20911,N_14286,N_13984);
and U20912 (N_20912,N_15163,N_17657);
xor U20913 (N_20913,N_13566,N_17140);
nor U20914 (N_20914,N_13489,N_16392);
and U20915 (N_20915,N_16844,N_16164);
nand U20916 (N_20916,N_15541,N_17784);
nor U20917 (N_20917,N_16599,N_13115);
and U20918 (N_20918,N_17588,N_13450);
and U20919 (N_20919,N_16812,N_15567);
xnor U20920 (N_20920,N_13065,N_14314);
xnor U20921 (N_20921,N_13134,N_15562);
and U20922 (N_20922,N_14866,N_15235);
or U20923 (N_20923,N_13479,N_16579);
or U20924 (N_20924,N_14853,N_12994);
nor U20925 (N_20925,N_13232,N_13840);
or U20926 (N_20926,N_16160,N_13522);
xnor U20927 (N_20927,N_16398,N_12069);
or U20928 (N_20928,N_15054,N_12971);
or U20929 (N_20929,N_13345,N_13256);
xor U20930 (N_20930,N_15279,N_14691);
xnor U20931 (N_20931,N_12811,N_12294);
nand U20932 (N_20932,N_12327,N_16455);
and U20933 (N_20933,N_17415,N_17102);
nand U20934 (N_20934,N_16924,N_14429);
nor U20935 (N_20935,N_13601,N_16236);
xor U20936 (N_20936,N_12497,N_13540);
nand U20937 (N_20937,N_14976,N_17682);
or U20938 (N_20938,N_15469,N_15064);
xor U20939 (N_20939,N_13887,N_17236);
or U20940 (N_20940,N_13229,N_14610);
xnor U20941 (N_20941,N_13788,N_16504);
nand U20942 (N_20942,N_16619,N_17086);
nand U20943 (N_20943,N_14561,N_15731);
xnor U20944 (N_20944,N_17670,N_12871);
or U20945 (N_20945,N_16351,N_12132);
nand U20946 (N_20946,N_17957,N_14709);
or U20947 (N_20947,N_15207,N_16306);
and U20948 (N_20948,N_14977,N_17562);
nand U20949 (N_20949,N_13269,N_16798);
nor U20950 (N_20950,N_17210,N_14226);
xor U20951 (N_20951,N_17203,N_12532);
or U20952 (N_20952,N_13771,N_14775);
nand U20953 (N_20953,N_15598,N_14020);
or U20954 (N_20954,N_15183,N_17664);
xnor U20955 (N_20955,N_14356,N_12798);
and U20956 (N_20956,N_14950,N_14614);
and U20957 (N_20957,N_13895,N_13588);
xor U20958 (N_20958,N_12989,N_17098);
nand U20959 (N_20959,N_16200,N_16091);
and U20960 (N_20960,N_13320,N_13988);
nand U20961 (N_20961,N_17450,N_16708);
and U20962 (N_20962,N_17552,N_15506);
nand U20963 (N_20963,N_16196,N_15004);
and U20964 (N_20964,N_13058,N_14659);
xor U20965 (N_20965,N_13162,N_16760);
and U20966 (N_20966,N_13537,N_13485);
or U20967 (N_20967,N_13786,N_16206);
or U20968 (N_20968,N_14010,N_13203);
xnor U20969 (N_20969,N_15579,N_17698);
nand U20970 (N_20970,N_14727,N_15890);
xor U20971 (N_20971,N_17750,N_15014);
nor U20972 (N_20972,N_15812,N_12297);
xor U20973 (N_20973,N_13860,N_17131);
and U20974 (N_20974,N_13827,N_13201);
nor U20975 (N_20975,N_15891,N_13679);
xor U20976 (N_20976,N_14229,N_15085);
or U20977 (N_20977,N_13205,N_16876);
xnor U20978 (N_20978,N_12052,N_15803);
nand U20979 (N_20979,N_16288,N_13175);
xor U20980 (N_20980,N_13384,N_12547);
xnor U20981 (N_20981,N_17633,N_15942);
or U20982 (N_20982,N_14170,N_14516);
xnor U20983 (N_20983,N_17702,N_16354);
or U20984 (N_20984,N_12769,N_15655);
nor U20985 (N_20985,N_14133,N_16738);
xnor U20986 (N_20986,N_14466,N_16414);
nor U20987 (N_20987,N_14443,N_16891);
xor U20988 (N_20988,N_15854,N_15809);
xor U20989 (N_20989,N_14348,N_13623);
xnor U20990 (N_20990,N_17448,N_15221);
or U20991 (N_20991,N_14471,N_17514);
and U20992 (N_20992,N_16086,N_16942);
nand U20993 (N_20993,N_13031,N_14077);
nand U20994 (N_20994,N_16052,N_16142);
nand U20995 (N_20995,N_15990,N_12789);
or U20996 (N_20996,N_14842,N_16982);
nor U20997 (N_20997,N_17444,N_16493);
or U20998 (N_20998,N_12999,N_14024);
and U20999 (N_20999,N_16213,N_13721);
or U21000 (N_21000,N_14674,N_12196);
nor U21001 (N_21001,N_14892,N_14375);
nand U21002 (N_21002,N_14020,N_15124);
and U21003 (N_21003,N_17869,N_16987);
and U21004 (N_21004,N_13811,N_13162);
or U21005 (N_21005,N_15770,N_17312);
nor U21006 (N_21006,N_14986,N_13973);
nor U21007 (N_21007,N_14530,N_16719);
nor U21008 (N_21008,N_14870,N_15668);
and U21009 (N_21009,N_16492,N_15066);
nor U21010 (N_21010,N_16657,N_13212);
nor U21011 (N_21011,N_17313,N_15662);
nand U21012 (N_21012,N_15072,N_13947);
and U21013 (N_21013,N_16005,N_16555);
or U21014 (N_21014,N_17320,N_13932);
xnor U21015 (N_21015,N_14379,N_16174);
and U21016 (N_21016,N_17547,N_15966);
nor U21017 (N_21017,N_15193,N_13158);
or U21018 (N_21018,N_13185,N_17462);
xnor U21019 (N_21019,N_13062,N_15134);
nor U21020 (N_21020,N_17771,N_16253);
nor U21021 (N_21021,N_16142,N_17940);
nor U21022 (N_21022,N_16454,N_13188);
and U21023 (N_21023,N_14345,N_13045);
nor U21024 (N_21024,N_15785,N_12731);
or U21025 (N_21025,N_12943,N_13266);
xor U21026 (N_21026,N_17805,N_12882);
nor U21027 (N_21027,N_16126,N_17973);
and U21028 (N_21028,N_14378,N_15169);
xnor U21029 (N_21029,N_12095,N_13977);
and U21030 (N_21030,N_12007,N_17822);
or U21031 (N_21031,N_12047,N_17408);
and U21032 (N_21032,N_17315,N_16837);
or U21033 (N_21033,N_15123,N_12859);
or U21034 (N_21034,N_14981,N_13804);
and U21035 (N_21035,N_12849,N_17072);
and U21036 (N_21036,N_13896,N_16263);
xor U21037 (N_21037,N_16815,N_16674);
or U21038 (N_21038,N_17302,N_13857);
xnor U21039 (N_21039,N_15043,N_16764);
and U21040 (N_21040,N_12913,N_12626);
nor U21041 (N_21041,N_16077,N_17914);
xnor U21042 (N_21042,N_14623,N_14854);
or U21043 (N_21043,N_12378,N_17271);
nand U21044 (N_21044,N_17854,N_15256);
nor U21045 (N_21045,N_14142,N_15718);
nand U21046 (N_21046,N_12332,N_15935);
nor U21047 (N_21047,N_16949,N_15702);
xnor U21048 (N_21048,N_17959,N_13912);
nor U21049 (N_21049,N_17246,N_17397);
nor U21050 (N_21050,N_17582,N_14454);
xor U21051 (N_21051,N_15701,N_16726);
or U21052 (N_21052,N_16154,N_15262);
and U21053 (N_21053,N_17217,N_16453);
nor U21054 (N_21054,N_12187,N_16969);
nor U21055 (N_21055,N_12348,N_13900);
xnor U21056 (N_21056,N_13146,N_12234);
nor U21057 (N_21057,N_13767,N_16142);
xor U21058 (N_21058,N_12805,N_13870);
nor U21059 (N_21059,N_13706,N_16967);
nand U21060 (N_21060,N_17761,N_14057);
xnor U21061 (N_21061,N_14451,N_17456);
or U21062 (N_21062,N_16236,N_15384);
nor U21063 (N_21063,N_15441,N_17117);
and U21064 (N_21064,N_12801,N_12138);
nor U21065 (N_21065,N_13398,N_13795);
nand U21066 (N_21066,N_13002,N_17472);
xor U21067 (N_21067,N_12005,N_17621);
and U21068 (N_21068,N_13880,N_13198);
and U21069 (N_21069,N_13911,N_17561);
or U21070 (N_21070,N_17874,N_16968);
nand U21071 (N_21071,N_16644,N_17062);
nand U21072 (N_21072,N_12168,N_16680);
nor U21073 (N_21073,N_15075,N_15095);
nand U21074 (N_21074,N_16177,N_14828);
nand U21075 (N_21075,N_13097,N_16785);
and U21076 (N_21076,N_12222,N_15997);
xnor U21077 (N_21077,N_14702,N_13976);
xor U21078 (N_21078,N_13490,N_13895);
xor U21079 (N_21079,N_16247,N_16248);
xor U21080 (N_21080,N_14608,N_16949);
xor U21081 (N_21081,N_13417,N_16250);
xnor U21082 (N_21082,N_15877,N_17647);
and U21083 (N_21083,N_16083,N_12914);
or U21084 (N_21084,N_12148,N_17910);
nand U21085 (N_21085,N_12288,N_12677);
and U21086 (N_21086,N_12290,N_12297);
xnor U21087 (N_21087,N_17127,N_12169);
nor U21088 (N_21088,N_17277,N_14242);
xnor U21089 (N_21089,N_12520,N_17971);
and U21090 (N_21090,N_12250,N_13259);
nor U21091 (N_21091,N_17292,N_16274);
nand U21092 (N_21092,N_14142,N_17924);
xor U21093 (N_21093,N_13323,N_13494);
nor U21094 (N_21094,N_14449,N_16046);
or U21095 (N_21095,N_16960,N_13928);
nor U21096 (N_21096,N_12475,N_15030);
xnor U21097 (N_21097,N_14697,N_16533);
or U21098 (N_21098,N_16902,N_16907);
and U21099 (N_21099,N_15785,N_15568);
nor U21100 (N_21100,N_13919,N_15004);
xnor U21101 (N_21101,N_15324,N_14672);
and U21102 (N_21102,N_14779,N_15745);
nor U21103 (N_21103,N_12101,N_17852);
and U21104 (N_21104,N_15623,N_13863);
nor U21105 (N_21105,N_16703,N_15385);
or U21106 (N_21106,N_16157,N_12166);
nand U21107 (N_21107,N_14926,N_14291);
and U21108 (N_21108,N_15167,N_15523);
nor U21109 (N_21109,N_13902,N_15466);
nand U21110 (N_21110,N_16240,N_17202);
nand U21111 (N_21111,N_14279,N_15422);
and U21112 (N_21112,N_12060,N_17545);
nor U21113 (N_21113,N_16132,N_13703);
and U21114 (N_21114,N_16988,N_15681);
and U21115 (N_21115,N_12671,N_13081);
or U21116 (N_21116,N_14570,N_16307);
nand U21117 (N_21117,N_16244,N_12482);
or U21118 (N_21118,N_16550,N_17233);
or U21119 (N_21119,N_16652,N_16433);
nor U21120 (N_21120,N_13378,N_16660);
xnor U21121 (N_21121,N_13764,N_15289);
and U21122 (N_21122,N_13118,N_14153);
or U21123 (N_21123,N_13482,N_16263);
nand U21124 (N_21124,N_13781,N_15987);
nand U21125 (N_21125,N_17732,N_13635);
xnor U21126 (N_21126,N_15435,N_15951);
xnor U21127 (N_21127,N_14681,N_14789);
nand U21128 (N_21128,N_16960,N_16443);
and U21129 (N_21129,N_15195,N_15976);
nor U21130 (N_21130,N_16975,N_17828);
xor U21131 (N_21131,N_13521,N_15442);
nand U21132 (N_21132,N_17406,N_15592);
nor U21133 (N_21133,N_14940,N_17308);
and U21134 (N_21134,N_17675,N_17997);
and U21135 (N_21135,N_16730,N_14589);
nor U21136 (N_21136,N_16257,N_14068);
xnor U21137 (N_21137,N_16443,N_17953);
nor U21138 (N_21138,N_12705,N_16896);
and U21139 (N_21139,N_14128,N_14017);
or U21140 (N_21140,N_17181,N_17099);
and U21141 (N_21141,N_16099,N_13875);
or U21142 (N_21142,N_15518,N_14884);
or U21143 (N_21143,N_15089,N_17433);
nor U21144 (N_21144,N_13991,N_14167);
nand U21145 (N_21145,N_17745,N_13122);
nand U21146 (N_21146,N_13381,N_13939);
and U21147 (N_21147,N_14478,N_16719);
and U21148 (N_21148,N_15670,N_17694);
nand U21149 (N_21149,N_14344,N_13844);
and U21150 (N_21150,N_12660,N_15526);
and U21151 (N_21151,N_15504,N_14779);
and U21152 (N_21152,N_17475,N_17529);
nor U21153 (N_21153,N_14469,N_15718);
and U21154 (N_21154,N_15490,N_12092);
nor U21155 (N_21155,N_13681,N_14019);
xor U21156 (N_21156,N_15341,N_17712);
xnor U21157 (N_21157,N_14393,N_17139);
nor U21158 (N_21158,N_14440,N_12617);
nand U21159 (N_21159,N_15450,N_12517);
and U21160 (N_21160,N_16812,N_15721);
nand U21161 (N_21161,N_14633,N_16379);
or U21162 (N_21162,N_16244,N_15269);
nor U21163 (N_21163,N_15098,N_12733);
or U21164 (N_21164,N_12987,N_17573);
xor U21165 (N_21165,N_13564,N_15425);
xnor U21166 (N_21166,N_17539,N_15193);
nor U21167 (N_21167,N_12804,N_15056);
and U21168 (N_21168,N_12581,N_15382);
xnor U21169 (N_21169,N_17598,N_14599);
and U21170 (N_21170,N_15517,N_13159);
nand U21171 (N_21171,N_17051,N_15924);
or U21172 (N_21172,N_13737,N_16810);
nand U21173 (N_21173,N_13095,N_15786);
nand U21174 (N_21174,N_15163,N_12066);
nor U21175 (N_21175,N_15238,N_13749);
and U21176 (N_21176,N_17904,N_17155);
nor U21177 (N_21177,N_13935,N_12915);
xor U21178 (N_21178,N_12024,N_15796);
nand U21179 (N_21179,N_13192,N_15253);
or U21180 (N_21180,N_15449,N_15484);
or U21181 (N_21181,N_14706,N_15107);
xnor U21182 (N_21182,N_13991,N_16558);
nor U21183 (N_21183,N_14786,N_17976);
and U21184 (N_21184,N_13710,N_14944);
xor U21185 (N_21185,N_15083,N_12130);
xnor U21186 (N_21186,N_17521,N_13016);
or U21187 (N_21187,N_15744,N_12564);
or U21188 (N_21188,N_17931,N_12068);
xnor U21189 (N_21189,N_14820,N_14680);
and U21190 (N_21190,N_14504,N_17955);
or U21191 (N_21191,N_12878,N_16755);
or U21192 (N_21192,N_14992,N_12036);
and U21193 (N_21193,N_12155,N_17591);
nand U21194 (N_21194,N_14971,N_13906);
nand U21195 (N_21195,N_15347,N_14149);
and U21196 (N_21196,N_12670,N_12135);
nand U21197 (N_21197,N_14646,N_17057);
nand U21198 (N_21198,N_13119,N_13047);
nor U21199 (N_21199,N_12551,N_13569);
nand U21200 (N_21200,N_15055,N_12039);
nor U21201 (N_21201,N_14902,N_16442);
and U21202 (N_21202,N_13159,N_17524);
nor U21203 (N_21203,N_16005,N_15758);
nor U21204 (N_21204,N_13408,N_17691);
and U21205 (N_21205,N_16056,N_16686);
nand U21206 (N_21206,N_15257,N_13374);
or U21207 (N_21207,N_15669,N_14103);
and U21208 (N_21208,N_15195,N_14574);
xor U21209 (N_21209,N_17210,N_12559);
and U21210 (N_21210,N_13972,N_13888);
nand U21211 (N_21211,N_12795,N_14789);
nor U21212 (N_21212,N_15976,N_16627);
xor U21213 (N_21213,N_17137,N_12983);
or U21214 (N_21214,N_12872,N_14556);
and U21215 (N_21215,N_15073,N_16296);
nor U21216 (N_21216,N_12784,N_14252);
or U21217 (N_21217,N_17077,N_12947);
xor U21218 (N_21218,N_14949,N_13581);
nor U21219 (N_21219,N_14197,N_13166);
nand U21220 (N_21220,N_15586,N_15543);
or U21221 (N_21221,N_14242,N_13904);
and U21222 (N_21222,N_13335,N_14244);
nand U21223 (N_21223,N_16571,N_15597);
nor U21224 (N_21224,N_13799,N_16959);
or U21225 (N_21225,N_15375,N_15924);
nor U21226 (N_21226,N_14897,N_14997);
or U21227 (N_21227,N_15399,N_13509);
nand U21228 (N_21228,N_15386,N_14777);
or U21229 (N_21229,N_17832,N_16225);
nor U21230 (N_21230,N_14490,N_16177);
or U21231 (N_21231,N_17341,N_15919);
or U21232 (N_21232,N_13380,N_17986);
or U21233 (N_21233,N_17569,N_12780);
nor U21234 (N_21234,N_13031,N_15327);
and U21235 (N_21235,N_12589,N_13165);
nor U21236 (N_21236,N_14161,N_13347);
xnor U21237 (N_21237,N_16540,N_13426);
or U21238 (N_21238,N_17149,N_14864);
or U21239 (N_21239,N_15814,N_16340);
xor U21240 (N_21240,N_14936,N_17778);
nand U21241 (N_21241,N_14322,N_13167);
nand U21242 (N_21242,N_14699,N_16627);
xor U21243 (N_21243,N_17396,N_14375);
xnor U21244 (N_21244,N_15197,N_15106);
nand U21245 (N_21245,N_17958,N_16666);
and U21246 (N_21246,N_17893,N_17678);
nor U21247 (N_21247,N_14935,N_17165);
nor U21248 (N_21248,N_15723,N_12845);
or U21249 (N_21249,N_14847,N_15979);
nor U21250 (N_21250,N_15477,N_12347);
nand U21251 (N_21251,N_12283,N_15136);
nand U21252 (N_21252,N_17374,N_12362);
or U21253 (N_21253,N_16790,N_14772);
nor U21254 (N_21254,N_14505,N_15421);
xnor U21255 (N_21255,N_14721,N_17574);
and U21256 (N_21256,N_15257,N_14445);
or U21257 (N_21257,N_14208,N_15404);
nand U21258 (N_21258,N_14885,N_12438);
xor U21259 (N_21259,N_12145,N_15937);
xor U21260 (N_21260,N_15801,N_14165);
or U21261 (N_21261,N_13985,N_13962);
nor U21262 (N_21262,N_12741,N_14370);
nand U21263 (N_21263,N_16853,N_16199);
nor U21264 (N_21264,N_17587,N_15234);
and U21265 (N_21265,N_17962,N_16960);
or U21266 (N_21266,N_16145,N_14554);
and U21267 (N_21267,N_17778,N_14481);
nand U21268 (N_21268,N_14382,N_16570);
xor U21269 (N_21269,N_14869,N_12232);
xor U21270 (N_21270,N_17321,N_17827);
and U21271 (N_21271,N_16122,N_16081);
nor U21272 (N_21272,N_14946,N_12402);
xor U21273 (N_21273,N_14740,N_12686);
nor U21274 (N_21274,N_12696,N_14310);
or U21275 (N_21275,N_17945,N_16289);
nand U21276 (N_21276,N_13479,N_13030);
nand U21277 (N_21277,N_12244,N_13001);
nor U21278 (N_21278,N_13404,N_17862);
xor U21279 (N_21279,N_14958,N_16470);
or U21280 (N_21280,N_13121,N_16510);
and U21281 (N_21281,N_16307,N_12532);
xor U21282 (N_21282,N_16922,N_16492);
nor U21283 (N_21283,N_15414,N_13920);
nand U21284 (N_21284,N_16604,N_15826);
and U21285 (N_21285,N_13583,N_16551);
nand U21286 (N_21286,N_15264,N_17329);
nand U21287 (N_21287,N_16797,N_13716);
nor U21288 (N_21288,N_15322,N_13271);
nor U21289 (N_21289,N_14472,N_14452);
xnor U21290 (N_21290,N_13076,N_17282);
or U21291 (N_21291,N_16652,N_16359);
nand U21292 (N_21292,N_12703,N_15290);
nand U21293 (N_21293,N_15976,N_17984);
xnor U21294 (N_21294,N_13399,N_17459);
xor U21295 (N_21295,N_14474,N_16808);
nor U21296 (N_21296,N_12362,N_16570);
and U21297 (N_21297,N_13252,N_13557);
nand U21298 (N_21298,N_15249,N_16083);
xor U21299 (N_21299,N_13100,N_15521);
nand U21300 (N_21300,N_17535,N_13579);
or U21301 (N_21301,N_14696,N_12930);
and U21302 (N_21302,N_16962,N_15696);
xor U21303 (N_21303,N_16762,N_13873);
or U21304 (N_21304,N_16709,N_12364);
and U21305 (N_21305,N_15809,N_12209);
and U21306 (N_21306,N_17668,N_14816);
nand U21307 (N_21307,N_17567,N_17191);
or U21308 (N_21308,N_13720,N_12679);
nand U21309 (N_21309,N_13081,N_13844);
nand U21310 (N_21310,N_14462,N_16142);
nand U21311 (N_21311,N_13978,N_17211);
nor U21312 (N_21312,N_12413,N_15807);
xor U21313 (N_21313,N_12926,N_15420);
and U21314 (N_21314,N_15629,N_14641);
xnor U21315 (N_21315,N_16141,N_15698);
and U21316 (N_21316,N_13947,N_13769);
nor U21317 (N_21317,N_14518,N_13691);
nand U21318 (N_21318,N_13336,N_14988);
or U21319 (N_21319,N_15205,N_13421);
xor U21320 (N_21320,N_13176,N_12665);
nor U21321 (N_21321,N_16875,N_16358);
xnor U21322 (N_21322,N_14325,N_15226);
xnor U21323 (N_21323,N_15544,N_16233);
or U21324 (N_21324,N_14488,N_17314);
and U21325 (N_21325,N_12914,N_15242);
nand U21326 (N_21326,N_12836,N_17034);
nand U21327 (N_21327,N_14035,N_14693);
nor U21328 (N_21328,N_13188,N_17626);
or U21329 (N_21329,N_16697,N_12283);
or U21330 (N_21330,N_12189,N_14601);
and U21331 (N_21331,N_15482,N_17224);
or U21332 (N_21332,N_17592,N_15990);
or U21333 (N_21333,N_17305,N_17721);
nor U21334 (N_21334,N_16138,N_16972);
and U21335 (N_21335,N_14317,N_16759);
and U21336 (N_21336,N_14067,N_17732);
nor U21337 (N_21337,N_13097,N_16830);
nor U21338 (N_21338,N_17746,N_13693);
or U21339 (N_21339,N_12631,N_14435);
xnor U21340 (N_21340,N_15415,N_16493);
or U21341 (N_21341,N_13724,N_17253);
xnor U21342 (N_21342,N_16715,N_17878);
nand U21343 (N_21343,N_15761,N_14658);
nor U21344 (N_21344,N_17740,N_14396);
xor U21345 (N_21345,N_13042,N_15728);
nor U21346 (N_21346,N_14323,N_16372);
and U21347 (N_21347,N_17831,N_17850);
and U21348 (N_21348,N_15733,N_14077);
nor U21349 (N_21349,N_15087,N_13081);
xor U21350 (N_21350,N_12011,N_12648);
and U21351 (N_21351,N_13010,N_13911);
or U21352 (N_21352,N_12911,N_16680);
nor U21353 (N_21353,N_17411,N_12498);
xor U21354 (N_21354,N_17612,N_17502);
xnor U21355 (N_21355,N_14468,N_17471);
xor U21356 (N_21356,N_15297,N_13399);
nor U21357 (N_21357,N_17258,N_17412);
xor U21358 (N_21358,N_13104,N_12152);
xnor U21359 (N_21359,N_14928,N_14281);
nand U21360 (N_21360,N_16001,N_17321);
nor U21361 (N_21361,N_14266,N_13759);
nand U21362 (N_21362,N_14347,N_13591);
or U21363 (N_21363,N_15458,N_15374);
xnor U21364 (N_21364,N_12374,N_15563);
nor U21365 (N_21365,N_12994,N_12517);
and U21366 (N_21366,N_14141,N_16622);
nand U21367 (N_21367,N_17480,N_12649);
or U21368 (N_21368,N_15197,N_13767);
and U21369 (N_21369,N_12052,N_12829);
xnor U21370 (N_21370,N_17258,N_13352);
or U21371 (N_21371,N_16715,N_12340);
xnor U21372 (N_21372,N_15200,N_14498);
xor U21373 (N_21373,N_17480,N_12029);
nor U21374 (N_21374,N_12467,N_16933);
and U21375 (N_21375,N_12793,N_12554);
nand U21376 (N_21376,N_13918,N_16861);
xnor U21377 (N_21377,N_16924,N_13539);
nand U21378 (N_21378,N_17995,N_16873);
and U21379 (N_21379,N_17813,N_15052);
and U21380 (N_21380,N_13724,N_14765);
xor U21381 (N_21381,N_15671,N_14102);
xor U21382 (N_21382,N_15342,N_15744);
or U21383 (N_21383,N_15779,N_16662);
and U21384 (N_21384,N_13191,N_13092);
xnor U21385 (N_21385,N_16738,N_15302);
xor U21386 (N_21386,N_16805,N_17982);
or U21387 (N_21387,N_16846,N_15469);
xor U21388 (N_21388,N_16443,N_12237);
or U21389 (N_21389,N_16164,N_16647);
or U21390 (N_21390,N_12824,N_16487);
and U21391 (N_21391,N_14843,N_16417);
or U21392 (N_21392,N_17485,N_14682);
nor U21393 (N_21393,N_16920,N_13214);
xor U21394 (N_21394,N_13572,N_13302);
nand U21395 (N_21395,N_15966,N_14245);
and U21396 (N_21396,N_12380,N_12762);
xor U21397 (N_21397,N_16746,N_13604);
nor U21398 (N_21398,N_17990,N_17839);
nand U21399 (N_21399,N_16911,N_16487);
xor U21400 (N_21400,N_17253,N_13472);
and U21401 (N_21401,N_16412,N_14213);
and U21402 (N_21402,N_14955,N_16383);
and U21403 (N_21403,N_12498,N_16537);
or U21404 (N_21404,N_15630,N_13191);
nor U21405 (N_21405,N_15876,N_16570);
nand U21406 (N_21406,N_13753,N_13669);
or U21407 (N_21407,N_12254,N_16349);
nor U21408 (N_21408,N_17013,N_17168);
xor U21409 (N_21409,N_12598,N_16042);
nor U21410 (N_21410,N_12684,N_15790);
nor U21411 (N_21411,N_15482,N_17430);
or U21412 (N_21412,N_12024,N_17430);
or U21413 (N_21413,N_17425,N_15786);
nor U21414 (N_21414,N_13181,N_13595);
or U21415 (N_21415,N_14804,N_13450);
nor U21416 (N_21416,N_12780,N_16685);
or U21417 (N_21417,N_16346,N_13620);
xnor U21418 (N_21418,N_12686,N_17851);
or U21419 (N_21419,N_14292,N_12096);
nor U21420 (N_21420,N_15231,N_15252);
xnor U21421 (N_21421,N_13036,N_13251);
xor U21422 (N_21422,N_14815,N_14574);
or U21423 (N_21423,N_15406,N_16929);
xor U21424 (N_21424,N_14155,N_15043);
and U21425 (N_21425,N_12162,N_12882);
or U21426 (N_21426,N_17753,N_16713);
or U21427 (N_21427,N_17524,N_17415);
xnor U21428 (N_21428,N_17757,N_16399);
or U21429 (N_21429,N_13357,N_15261);
nand U21430 (N_21430,N_16724,N_14869);
or U21431 (N_21431,N_15053,N_12521);
or U21432 (N_21432,N_12828,N_13017);
nand U21433 (N_21433,N_17116,N_13301);
nand U21434 (N_21434,N_17041,N_16456);
xnor U21435 (N_21435,N_16575,N_16900);
and U21436 (N_21436,N_12749,N_17007);
or U21437 (N_21437,N_12221,N_16141);
nor U21438 (N_21438,N_15922,N_17963);
nor U21439 (N_21439,N_12662,N_12417);
nand U21440 (N_21440,N_13003,N_14869);
xnor U21441 (N_21441,N_13374,N_12005);
xnor U21442 (N_21442,N_12051,N_16692);
nor U21443 (N_21443,N_12510,N_17822);
or U21444 (N_21444,N_12919,N_13258);
xnor U21445 (N_21445,N_12347,N_13770);
or U21446 (N_21446,N_12796,N_15697);
or U21447 (N_21447,N_14425,N_13993);
and U21448 (N_21448,N_12006,N_15082);
nand U21449 (N_21449,N_15487,N_13913);
nand U21450 (N_21450,N_17171,N_12909);
nand U21451 (N_21451,N_17515,N_12960);
or U21452 (N_21452,N_17723,N_13465);
xor U21453 (N_21453,N_16526,N_16907);
nor U21454 (N_21454,N_14759,N_15425);
and U21455 (N_21455,N_12081,N_14035);
or U21456 (N_21456,N_16853,N_15062);
xnor U21457 (N_21457,N_14157,N_14439);
or U21458 (N_21458,N_14078,N_17607);
and U21459 (N_21459,N_16080,N_14041);
nor U21460 (N_21460,N_14891,N_13740);
and U21461 (N_21461,N_14962,N_12950);
or U21462 (N_21462,N_14721,N_16258);
or U21463 (N_21463,N_16295,N_15371);
and U21464 (N_21464,N_13479,N_12430);
xor U21465 (N_21465,N_14936,N_14850);
nand U21466 (N_21466,N_14717,N_15107);
nand U21467 (N_21467,N_16470,N_15574);
nand U21468 (N_21468,N_16568,N_12829);
and U21469 (N_21469,N_15582,N_17355);
and U21470 (N_21470,N_14631,N_13901);
xnor U21471 (N_21471,N_15570,N_15280);
nand U21472 (N_21472,N_14240,N_17137);
nand U21473 (N_21473,N_14030,N_15064);
and U21474 (N_21474,N_12353,N_14661);
xnor U21475 (N_21475,N_13899,N_14697);
xnor U21476 (N_21476,N_17191,N_12688);
or U21477 (N_21477,N_15425,N_13674);
xnor U21478 (N_21478,N_15004,N_16800);
xnor U21479 (N_21479,N_13008,N_17748);
nand U21480 (N_21480,N_17285,N_15172);
xnor U21481 (N_21481,N_13435,N_17276);
xnor U21482 (N_21482,N_13344,N_12096);
and U21483 (N_21483,N_15223,N_14318);
xor U21484 (N_21484,N_14909,N_12001);
xor U21485 (N_21485,N_13806,N_16997);
or U21486 (N_21486,N_17259,N_15684);
xor U21487 (N_21487,N_13594,N_13821);
nand U21488 (N_21488,N_16631,N_13548);
or U21489 (N_21489,N_17948,N_17557);
and U21490 (N_21490,N_12726,N_15528);
xnor U21491 (N_21491,N_14634,N_12224);
nor U21492 (N_21492,N_12628,N_14429);
nor U21493 (N_21493,N_15938,N_13174);
or U21494 (N_21494,N_13759,N_13536);
or U21495 (N_21495,N_14763,N_12213);
or U21496 (N_21496,N_17579,N_13188);
nor U21497 (N_21497,N_13337,N_16739);
nor U21498 (N_21498,N_14664,N_16014);
xor U21499 (N_21499,N_12506,N_16968);
or U21500 (N_21500,N_12961,N_12945);
nor U21501 (N_21501,N_17316,N_14160);
nor U21502 (N_21502,N_13315,N_15220);
nor U21503 (N_21503,N_13422,N_15950);
nand U21504 (N_21504,N_15325,N_15985);
nor U21505 (N_21505,N_12418,N_16142);
xor U21506 (N_21506,N_13900,N_13058);
xor U21507 (N_21507,N_17977,N_17888);
and U21508 (N_21508,N_13388,N_17455);
nand U21509 (N_21509,N_14947,N_14294);
nand U21510 (N_21510,N_17898,N_13714);
xnor U21511 (N_21511,N_12795,N_16172);
and U21512 (N_21512,N_16427,N_14318);
and U21513 (N_21513,N_17405,N_16433);
nand U21514 (N_21514,N_17056,N_12537);
and U21515 (N_21515,N_16201,N_17660);
or U21516 (N_21516,N_13521,N_17132);
or U21517 (N_21517,N_17724,N_15781);
xor U21518 (N_21518,N_15216,N_16830);
xnor U21519 (N_21519,N_17243,N_17249);
or U21520 (N_21520,N_16007,N_14483);
nand U21521 (N_21521,N_16495,N_12483);
and U21522 (N_21522,N_13130,N_15309);
or U21523 (N_21523,N_13589,N_16694);
xor U21524 (N_21524,N_16858,N_15008);
and U21525 (N_21525,N_17105,N_14543);
or U21526 (N_21526,N_12875,N_15775);
or U21527 (N_21527,N_15946,N_13189);
nor U21528 (N_21528,N_14098,N_12923);
nor U21529 (N_21529,N_16576,N_16337);
xor U21530 (N_21530,N_14739,N_13974);
nand U21531 (N_21531,N_17229,N_14836);
and U21532 (N_21532,N_15402,N_14454);
nor U21533 (N_21533,N_14892,N_16013);
or U21534 (N_21534,N_15002,N_16429);
nand U21535 (N_21535,N_16978,N_13012);
xnor U21536 (N_21536,N_14383,N_12409);
nand U21537 (N_21537,N_12738,N_12529);
or U21538 (N_21538,N_15117,N_16063);
xor U21539 (N_21539,N_12387,N_15249);
and U21540 (N_21540,N_15424,N_17886);
and U21541 (N_21541,N_13426,N_12585);
xnor U21542 (N_21542,N_16805,N_12608);
or U21543 (N_21543,N_14231,N_14793);
and U21544 (N_21544,N_15154,N_12503);
nand U21545 (N_21545,N_15642,N_15374);
and U21546 (N_21546,N_15458,N_15101);
or U21547 (N_21547,N_15604,N_15802);
or U21548 (N_21548,N_12932,N_17339);
and U21549 (N_21549,N_17554,N_17733);
and U21550 (N_21550,N_12383,N_14104);
nor U21551 (N_21551,N_13218,N_12640);
and U21552 (N_21552,N_13833,N_17202);
or U21553 (N_21553,N_15219,N_13895);
xor U21554 (N_21554,N_12779,N_16384);
nand U21555 (N_21555,N_14907,N_17054);
nand U21556 (N_21556,N_14675,N_16113);
nand U21557 (N_21557,N_13282,N_14924);
and U21558 (N_21558,N_12385,N_17604);
xnor U21559 (N_21559,N_14020,N_17639);
and U21560 (N_21560,N_17598,N_16821);
nor U21561 (N_21561,N_16634,N_16400);
nand U21562 (N_21562,N_14554,N_14153);
nand U21563 (N_21563,N_17686,N_15318);
nor U21564 (N_21564,N_12399,N_13405);
and U21565 (N_21565,N_13488,N_15004);
or U21566 (N_21566,N_17664,N_12110);
xnor U21567 (N_21567,N_15706,N_13611);
nand U21568 (N_21568,N_12140,N_14043);
and U21569 (N_21569,N_13784,N_13989);
nor U21570 (N_21570,N_14394,N_13920);
nor U21571 (N_21571,N_15506,N_14703);
xnor U21572 (N_21572,N_17523,N_12515);
nor U21573 (N_21573,N_16334,N_17131);
or U21574 (N_21574,N_12203,N_12131);
xnor U21575 (N_21575,N_14291,N_15021);
xnor U21576 (N_21576,N_16592,N_14954);
and U21577 (N_21577,N_15871,N_17746);
nand U21578 (N_21578,N_13000,N_16443);
or U21579 (N_21579,N_12745,N_15652);
and U21580 (N_21580,N_13371,N_15758);
nand U21581 (N_21581,N_16478,N_14313);
xnor U21582 (N_21582,N_17328,N_13072);
and U21583 (N_21583,N_17177,N_17724);
and U21584 (N_21584,N_16639,N_17971);
nor U21585 (N_21585,N_12091,N_15344);
nand U21586 (N_21586,N_13630,N_16781);
xor U21587 (N_21587,N_16455,N_17361);
xor U21588 (N_21588,N_17433,N_17882);
nand U21589 (N_21589,N_14541,N_16539);
xor U21590 (N_21590,N_12070,N_12389);
xor U21591 (N_21591,N_13015,N_15522);
or U21592 (N_21592,N_16370,N_15431);
nor U21593 (N_21593,N_12015,N_13035);
or U21594 (N_21594,N_12602,N_13645);
and U21595 (N_21595,N_14266,N_12210);
nor U21596 (N_21596,N_15222,N_15354);
nand U21597 (N_21597,N_16321,N_15369);
xor U21598 (N_21598,N_13690,N_17187);
nor U21599 (N_21599,N_12562,N_17497);
nand U21600 (N_21600,N_16133,N_12019);
or U21601 (N_21601,N_16917,N_17711);
and U21602 (N_21602,N_13187,N_15497);
nor U21603 (N_21603,N_16986,N_13591);
and U21604 (N_21604,N_17643,N_15145);
or U21605 (N_21605,N_16200,N_13160);
nand U21606 (N_21606,N_17956,N_14838);
nand U21607 (N_21607,N_14759,N_17879);
or U21608 (N_21608,N_12882,N_16803);
nand U21609 (N_21609,N_16080,N_15173);
nor U21610 (N_21610,N_17107,N_13216);
nor U21611 (N_21611,N_12044,N_13238);
nor U21612 (N_21612,N_17971,N_12991);
and U21613 (N_21613,N_16451,N_16883);
nand U21614 (N_21614,N_12158,N_17148);
nand U21615 (N_21615,N_12075,N_13404);
xnor U21616 (N_21616,N_14221,N_14241);
or U21617 (N_21617,N_14100,N_13779);
nor U21618 (N_21618,N_16104,N_12180);
xor U21619 (N_21619,N_16326,N_16148);
xnor U21620 (N_21620,N_15665,N_15431);
xnor U21621 (N_21621,N_17455,N_14583);
nor U21622 (N_21622,N_14182,N_14285);
xnor U21623 (N_21623,N_13179,N_12066);
nand U21624 (N_21624,N_12568,N_14707);
or U21625 (N_21625,N_17592,N_15822);
and U21626 (N_21626,N_16599,N_16071);
or U21627 (N_21627,N_12713,N_16860);
nand U21628 (N_21628,N_14960,N_12304);
and U21629 (N_21629,N_17543,N_12624);
nand U21630 (N_21630,N_15345,N_12703);
or U21631 (N_21631,N_14019,N_16681);
nand U21632 (N_21632,N_13448,N_13180);
nand U21633 (N_21633,N_16270,N_17311);
or U21634 (N_21634,N_15661,N_14312);
or U21635 (N_21635,N_15843,N_13479);
and U21636 (N_21636,N_16814,N_17690);
or U21637 (N_21637,N_15616,N_16303);
or U21638 (N_21638,N_17322,N_17563);
and U21639 (N_21639,N_15987,N_16134);
nor U21640 (N_21640,N_16765,N_14272);
nor U21641 (N_21641,N_14587,N_16663);
nand U21642 (N_21642,N_17174,N_14338);
nand U21643 (N_21643,N_16513,N_13700);
or U21644 (N_21644,N_17406,N_15151);
nand U21645 (N_21645,N_16367,N_16350);
and U21646 (N_21646,N_14439,N_12935);
nor U21647 (N_21647,N_17211,N_12934);
or U21648 (N_21648,N_16282,N_16891);
nand U21649 (N_21649,N_15501,N_15194);
nand U21650 (N_21650,N_16343,N_16915);
and U21651 (N_21651,N_14896,N_14961);
and U21652 (N_21652,N_13586,N_15923);
nand U21653 (N_21653,N_15833,N_16732);
and U21654 (N_21654,N_13596,N_15659);
nor U21655 (N_21655,N_14621,N_12806);
and U21656 (N_21656,N_17868,N_17788);
xor U21657 (N_21657,N_17579,N_13969);
or U21658 (N_21658,N_15165,N_13672);
nand U21659 (N_21659,N_16536,N_16288);
xor U21660 (N_21660,N_16087,N_12790);
and U21661 (N_21661,N_13015,N_13617);
nand U21662 (N_21662,N_14055,N_17821);
nand U21663 (N_21663,N_16068,N_16763);
and U21664 (N_21664,N_14078,N_13113);
nor U21665 (N_21665,N_17485,N_15555);
nand U21666 (N_21666,N_14014,N_17991);
and U21667 (N_21667,N_14740,N_16450);
nor U21668 (N_21668,N_13711,N_17749);
and U21669 (N_21669,N_13360,N_13070);
xor U21670 (N_21670,N_16142,N_16411);
xor U21671 (N_21671,N_13745,N_13434);
and U21672 (N_21672,N_16509,N_16753);
and U21673 (N_21673,N_13324,N_12631);
nand U21674 (N_21674,N_17120,N_12558);
xnor U21675 (N_21675,N_16638,N_16260);
and U21676 (N_21676,N_12748,N_16454);
xor U21677 (N_21677,N_13573,N_13134);
nand U21678 (N_21678,N_14548,N_13916);
xor U21679 (N_21679,N_17669,N_14977);
and U21680 (N_21680,N_13775,N_14034);
xor U21681 (N_21681,N_13347,N_12966);
nor U21682 (N_21682,N_13340,N_16683);
and U21683 (N_21683,N_16028,N_16902);
nor U21684 (N_21684,N_13972,N_17850);
and U21685 (N_21685,N_12786,N_12985);
nand U21686 (N_21686,N_17138,N_14084);
nor U21687 (N_21687,N_13480,N_17127);
nand U21688 (N_21688,N_17559,N_15339);
nor U21689 (N_21689,N_14012,N_14073);
nand U21690 (N_21690,N_14570,N_13616);
or U21691 (N_21691,N_15235,N_15906);
or U21692 (N_21692,N_17263,N_12354);
xnor U21693 (N_21693,N_13455,N_14422);
or U21694 (N_21694,N_15412,N_15159);
or U21695 (N_21695,N_14055,N_15882);
nand U21696 (N_21696,N_13265,N_15703);
or U21697 (N_21697,N_16384,N_14735);
xor U21698 (N_21698,N_16449,N_14178);
and U21699 (N_21699,N_16269,N_15560);
and U21700 (N_21700,N_15069,N_17791);
or U21701 (N_21701,N_13031,N_14364);
nor U21702 (N_21702,N_15391,N_14369);
or U21703 (N_21703,N_15526,N_16105);
nor U21704 (N_21704,N_15959,N_17914);
nor U21705 (N_21705,N_13902,N_15387);
nand U21706 (N_21706,N_13532,N_15405);
xor U21707 (N_21707,N_14252,N_15189);
or U21708 (N_21708,N_16268,N_12281);
or U21709 (N_21709,N_16388,N_17258);
xor U21710 (N_21710,N_16484,N_15800);
nand U21711 (N_21711,N_16174,N_13821);
xor U21712 (N_21712,N_12105,N_13765);
nand U21713 (N_21713,N_12418,N_17297);
or U21714 (N_21714,N_12210,N_17661);
xor U21715 (N_21715,N_13665,N_12219);
and U21716 (N_21716,N_15333,N_15181);
or U21717 (N_21717,N_15731,N_14795);
or U21718 (N_21718,N_13284,N_17406);
or U21719 (N_21719,N_12940,N_14535);
or U21720 (N_21720,N_13542,N_17826);
and U21721 (N_21721,N_13834,N_16816);
nor U21722 (N_21722,N_12219,N_15478);
nor U21723 (N_21723,N_12261,N_13981);
or U21724 (N_21724,N_15439,N_13253);
nand U21725 (N_21725,N_13859,N_17117);
or U21726 (N_21726,N_16841,N_15771);
or U21727 (N_21727,N_12554,N_15981);
nor U21728 (N_21728,N_12863,N_17211);
xor U21729 (N_21729,N_15895,N_13525);
or U21730 (N_21730,N_14937,N_13036);
nor U21731 (N_21731,N_16087,N_13487);
nand U21732 (N_21732,N_14179,N_17384);
nand U21733 (N_21733,N_14591,N_16145);
nor U21734 (N_21734,N_14776,N_12244);
and U21735 (N_21735,N_17367,N_16618);
or U21736 (N_21736,N_13676,N_16018);
or U21737 (N_21737,N_14355,N_14407);
xor U21738 (N_21738,N_13457,N_14697);
and U21739 (N_21739,N_14506,N_17717);
xnor U21740 (N_21740,N_15285,N_15669);
nor U21741 (N_21741,N_16994,N_14088);
nand U21742 (N_21742,N_15965,N_17746);
nand U21743 (N_21743,N_13906,N_16749);
and U21744 (N_21744,N_15076,N_13467);
and U21745 (N_21745,N_16600,N_13292);
nand U21746 (N_21746,N_12482,N_15799);
xnor U21747 (N_21747,N_14461,N_15437);
nand U21748 (N_21748,N_14150,N_17951);
nand U21749 (N_21749,N_17206,N_14309);
nor U21750 (N_21750,N_16448,N_13441);
xor U21751 (N_21751,N_13530,N_13379);
nand U21752 (N_21752,N_14307,N_13342);
nand U21753 (N_21753,N_16954,N_14798);
or U21754 (N_21754,N_16711,N_12063);
xor U21755 (N_21755,N_17074,N_14689);
xnor U21756 (N_21756,N_13571,N_15394);
and U21757 (N_21757,N_15544,N_14490);
xnor U21758 (N_21758,N_12057,N_15482);
nand U21759 (N_21759,N_15033,N_15274);
xor U21760 (N_21760,N_13281,N_16349);
xor U21761 (N_21761,N_17753,N_12331);
nor U21762 (N_21762,N_15277,N_12979);
nand U21763 (N_21763,N_17353,N_17853);
xor U21764 (N_21764,N_12842,N_12158);
or U21765 (N_21765,N_13597,N_16399);
and U21766 (N_21766,N_13242,N_12273);
nand U21767 (N_21767,N_15181,N_17405);
nand U21768 (N_21768,N_14035,N_17940);
and U21769 (N_21769,N_15546,N_17203);
nor U21770 (N_21770,N_13289,N_14234);
xnor U21771 (N_21771,N_14471,N_13333);
nor U21772 (N_21772,N_16455,N_12838);
or U21773 (N_21773,N_13600,N_12575);
nor U21774 (N_21774,N_16585,N_17546);
xnor U21775 (N_21775,N_12321,N_13884);
and U21776 (N_21776,N_15996,N_14579);
nand U21777 (N_21777,N_14094,N_14250);
xnor U21778 (N_21778,N_15098,N_16099);
nand U21779 (N_21779,N_17721,N_13240);
and U21780 (N_21780,N_14742,N_13942);
nor U21781 (N_21781,N_12183,N_13869);
nor U21782 (N_21782,N_13082,N_16631);
and U21783 (N_21783,N_14061,N_13110);
nand U21784 (N_21784,N_13476,N_16343);
nor U21785 (N_21785,N_14843,N_12729);
and U21786 (N_21786,N_15789,N_12504);
nor U21787 (N_21787,N_17527,N_14277);
nand U21788 (N_21788,N_17850,N_12966);
and U21789 (N_21789,N_15280,N_16121);
nor U21790 (N_21790,N_16741,N_15470);
nand U21791 (N_21791,N_15461,N_15042);
or U21792 (N_21792,N_13868,N_14898);
xor U21793 (N_21793,N_12378,N_13120);
nand U21794 (N_21794,N_16405,N_17114);
nand U21795 (N_21795,N_17656,N_15252);
nor U21796 (N_21796,N_13817,N_12697);
or U21797 (N_21797,N_13233,N_12861);
and U21798 (N_21798,N_17519,N_13235);
or U21799 (N_21799,N_12166,N_15486);
or U21800 (N_21800,N_13373,N_16841);
and U21801 (N_21801,N_14634,N_15769);
xnor U21802 (N_21802,N_15827,N_12415);
nand U21803 (N_21803,N_14324,N_17573);
xnor U21804 (N_21804,N_16054,N_13187);
nand U21805 (N_21805,N_13393,N_17620);
xor U21806 (N_21806,N_13017,N_15569);
xnor U21807 (N_21807,N_15872,N_17495);
nor U21808 (N_21808,N_14185,N_13163);
nand U21809 (N_21809,N_17388,N_17069);
and U21810 (N_21810,N_17460,N_16346);
nor U21811 (N_21811,N_13365,N_15284);
or U21812 (N_21812,N_17316,N_14686);
or U21813 (N_21813,N_13118,N_16033);
nor U21814 (N_21814,N_15447,N_12527);
nand U21815 (N_21815,N_16879,N_12798);
and U21816 (N_21816,N_14042,N_14018);
nor U21817 (N_21817,N_15153,N_17250);
and U21818 (N_21818,N_16150,N_16607);
or U21819 (N_21819,N_14115,N_14672);
nor U21820 (N_21820,N_12573,N_15129);
or U21821 (N_21821,N_12118,N_14248);
and U21822 (N_21822,N_13421,N_15400);
nand U21823 (N_21823,N_17135,N_12169);
nand U21824 (N_21824,N_12468,N_15395);
or U21825 (N_21825,N_15621,N_13385);
and U21826 (N_21826,N_16490,N_14476);
nor U21827 (N_21827,N_15078,N_17600);
nor U21828 (N_21828,N_13138,N_14671);
xnor U21829 (N_21829,N_12675,N_15212);
and U21830 (N_21830,N_16510,N_16042);
or U21831 (N_21831,N_17664,N_16375);
nor U21832 (N_21832,N_17435,N_12376);
nor U21833 (N_21833,N_14602,N_14951);
or U21834 (N_21834,N_17205,N_16407);
nor U21835 (N_21835,N_12330,N_16853);
nand U21836 (N_21836,N_13219,N_17889);
xor U21837 (N_21837,N_13505,N_14870);
and U21838 (N_21838,N_14560,N_12538);
xnor U21839 (N_21839,N_12868,N_16029);
xor U21840 (N_21840,N_13624,N_12073);
nor U21841 (N_21841,N_13963,N_16943);
xnor U21842 (N_21842,N_14894,N_17627);
nor U21843 (N_21843,N_15345,N_12484);
and U21844 (N_21844,N_16560,N_14405);
and U21845 (N_21845,N_17694,N_13783);
xnor U21846 (N_21846,N_15192,N_15472);
xor U21847 (N_21847,N_17023,N_13695);
nand U21848 (N_21848,N_13656,N_13878);
or U21849 (N_21849,N_12956,N_12785);
or U21850 (N_21850,N_13924,N_17445);
or U21851 (N_21851,N_15491,N_16337);
xnor U21852 (N_21852,N_16070,N_17554);
nand U21853 (N_21853,N_16815,N_12191);
or U21854 (N_21854,N_16907,N_14642);
xor U21855 (N_21855,N_13630,N_12427);
xor U21856 (N_21856,N_14578,N_14927);
or U21857 (N_21857,N_15848,N_14504);
and U21858 (N_21858,N_14548,N_15023);
xnor U21859 (N_21859,N_12962,N_17922);
or U21860 (N_21860,N_15582,N_16670);
or U21861 (N_21861,N_13744,N_12492);
nand U21862 (N_21862,N_14375,N_17428);
and U21863 (N_21863,N_15661,N_12163);
nand U21864 (N_21864,N_15367,N_17952);
nor U21865 (N_21865,N_15814,N_15705);
nor U21866 (N_21866,N_13649,N_13330);
nor U21867 (N_21867,N_14857,N_12207);
nand U21868 (N_21868,N_14639,N_14005);
nor U21869 (N_21869,N_13107,N_13354);
xor U21870 (N_21870,N_14414,N_16331);
nand U21871 (N_21871,N_17961,N_16532);
xnor U21872 (N_21872,N_16096,N_17798);
and U21873 (N_21873,N_15060,N_17428);
or U21874 (N_21874,N_14603,N_16824);
or U21875 (N_21875,N_14357,N_17610);
nor U21876 (N_21876,N_12847,N_14765);
or U21877 (N_21877,N_12992,N_15715);
nand U21878 (N_21878,N_14504,N_12085);
xor U21879 (N_21879,N_13213,N_14391);
or U21880 (N_21880,N_17433,N_14656);
or U21881 (N_21881,N_16091,N_14569);
or U21882 (N_21882,N_12475,N_13012);
or U21883 (N_21883,N_16529,N_17819);
and U21884 (N_21884,N_16481,N_12314);
or U21885 (N_21885,N_14221,N_14542);
and U21886 (N_21886,N_15390,N_15086);
or U21887 (N_21887,N_14324,N_14442);
xnor U21888 (N_21888,N_17743,N_15199);
or U21889 (N_21889,N_12777,N_13315);
nor U21890 (N_21890,N_14624,N_17894);
nor U21891 (N_21891,N_15652,N_12977);
nand U21892 (N_21892,N_14342,N_15039);
nand U21893 (N_21893,N_16242,N_15883);
nand U21894 (N_21894,N_16970,N_14097);
nand U21895 (N_21895,N_13973,N_14584);
and U21896 (N_21896,N_14471,N_14523);
and U21897 (N_21897,N_15538,N_13481);
xnor U21898 (N_21898,N_12734,N_16357);
and U21899 (N_21899,N_16368,N_14008);
or U21900 (N_21900,N_13720,N_14154);
nand U21901 (N_21901,N_16100,N_17712);
xnor U21902 (N_21902,N_15998,N_14927);
and U21903 (N_21903,N_16876,N_17704);
nor U21904 (N_21904,N_17636,N_16200);
nor U21905 (N_21905,N_16257,N_16306);
nor U21906 (N_21906,N_13450,N_13456);
and U21907 (N_21907,N_17801,N_14225);
nor U21908 (N_21908,N_12557,N_14262);
nand U21909 (N_21909,N_12857,N_14109);
nor U21910 (N_21910,N_17470,N_16698);
or U21911 (N_21911,N_13425,N_17153);
xnor U21912 (N_21912,N_13188,N_12169);
or U21913 (N_21913,N_15616,N_16687);
xor U21914 (N_21914,N_13161,N_17424);
or U21915 (N_21915,N_12966,N_12154);
xnor U21916 (N_21916,N_12769,N_13409);
nand U21917 (N_21917,N_15210,N_12523);
and U21918 (N_21918,N_15604,N_12500);
xor U21919 (N_21919,N_13035,N_14905);
or U21920 (N_21920,N_16279,N_13922);
nand U21921 (N_21921,N_12233,N_15858);
and U21922 (N_21922,N_13457,N_15244);
or U21923 (N_21923,N_17463,N_16755);
xor U21924 (N_21924,N_17030,N_17929);
xor U21925 (N_21925,N_13699,N_12341);
xor U21926 (N_21926,N_13377,N_17513);
xnor U21927 (N_21927,N_15875,N_13316);
nand U21928 (N_21928,N_16298,N_16075);
and U21929 (N_21929,N_17011,N_12075);
and U21930 (N_21930,N_17316,N_17537);
nand U21931 (N_21931,N_16139,N_15107);
or U21932 (N_21932,N_14359,N_15471);
and U21933 (N_21933,N_17942,N_14494);
and U21934 (N_21934,N_15031,N_13839);
nand U21935 (N_21935,N_15808,N_16094);
nor U21936 (N_21936,N_12487,N_12491);
or U21937 (N_21937,N_12906,N_16035);
xnor U21938 (N_21938,N_16819,N_16253);
xor U21939 (N_21939,N_14813,N_15409);
and U21940 (N_21940,N_14290,N_13940);
xnor U21941 (N_21941,N_14265,N_16903);
or U21942 (N_21942,N_13615,N_14898);
nand U21943 (N_21943,N_13987,N_15914);
xor U21944 (N_21944,N_16752,N_15558);
and U21945 (N_21945,N_13413,N_12431);
xnor U21946 (N_21946,N_12648,N_15594);
xor U21947 (N_21947,N_17093,N_16169);
or U21948 (N_21948,N_12271,N_16559);
nand U21949 (N_21949,N_17816,N_16348);
and U21950 (N_21950,N_13168,N_17612);
and U21951 (N_21951,N_12444,N_14525);
nand U21952 (N_21952,N_15111,N_14610);
nand U21953 (N_21953,N_12991,N_14242);
or U21954 (N_21954,N_13935,N_12833);
xnor U21955 (N_21955,N_13277,N_13196);
xor U21956 (N_21956,N_16753,N_17519);
xor U21957 (N_21957,N_16595,N_15746);
nand U21958 (N_21958,N_14756,N_13019);
xor U21959 (N_21959,N_12993,N_12249);
nor U21960 (N_21960,N_13382,N_12474);
nor U21961 (N_21961,N_17964,N_17946);
xor U21962 (N_21962,N_13524,N_12680);
xor U21963 (N_21963,N_13584,N_14144);
xnor U21964 (N_21964,N_14375,N_13665);
or U21965 (N_21965,N_14295,N_13038);
and U21966 (N_21966,N_12763,N_12630);
nor U21967 (N_21967,N_16192,N_12569);
nor U21968 (N_21968,N_16388,N_12286);
or U21969 (N_21969,N_17062,N_14421);
nor U21970 (N_21970,N_17195,N_12919);
nand U21971 (N_21971,N_16610,N_14939);
xnor U21972 (N_21972,N_13139,N_14161);
and U21973 (N_21973,N_15829,N_15251);
or U21974 (N_21974,N_14529,N_14730);
nand U21975 (N_21975,N_14664,N_15919);
or U21976 (N_21976,N_13551,N_12250);
nor U21977 (N_21977,N_13141,N_13711);
nor U21978 (N_21978,N_16252,N_16566);
and U21979 (N_21979,N_14953,N_16535);
nor U21980 (N_21980,N_16419,N_16223);
nand U21981 (N_21981,N_16144,N_15139);
and U21982 (N_21982,N_13109,N_15479);
or U21983 (N_21983,N_15980,N_16021);
or U21984 (N_21984,N_16280,N_14942);
nor U21985 (N_21985,N_15370,N_13683);
or U21986 (N_21986,N_16149,N_15718);
xor U21987 (N_21987,N_13085,N_14583);
or U21988 (N_21988,N_12465,N_13357);
and U21989 (N_21989,N_14705,N_17569);
and U21990 (N_21990,N_16497,N_15111);
or U21991 (N_21991,N_13925,N_12728);
or U21992 (N_21992,N_12430,N_12093);
xnor U21993 (N_21993,N_12595,N_16569);
nor U21994 (N_21994,N_12883,N_13114);
xor U21995 (N_21995,N_17645,N_12522);
or U21996 (N_21996,N_12489,N_14075);
nand U21997 (N_21997,N_14789,N_15719);
and U21998 (N_21998,N_14883,N_13695);
or U21999 (N_21999,N_15579,N_16234);
nor U22000 (N_22000,N_16409,N_17059);
xnor U22001 (N_22001,N_15420,N_14266);
nand U22002 (N_22002,N_12326,N_16672);
and U22003 (N_22003,N_17348,N_14198);
or U22004 (N_22004,N_16598,N_13203);
nor U22005 (N_22005,N_14727,N_17170);
xnor U22006 (N_22006,N_15502,N_14612);
and U22007 (N_22007,N_13736,N_12873);
or U22008 (N_22008,N_13006,N_15228);
or U22009 (N_22009,N_13875,N_13107);
xnor U22010 (N_22010,N_14708,N_12635);
nand U22011 (N_22011,N_14829,N_15280);
or U22012 (N_22012,N_14966,N_17725);
or U22013 (N_22013,N_13902,N_14825);
or U22014 (N_22014,N_17134,N_12240);
xor U22015 (N_22015,N_17007,N_13802);
nand U22016 (N_22016,N_13679,N_15454);
nor U22017 (N_22017,N_15044,N_16888);
or U22018 (N_22018,N_15276,N_14962);
nand U22019 (N_22019,N_13739,N_17202);
nor U22020 (N_22020,N_12508,N_17898);
or U22021 (N_22021,N_12952,N_12947);
nand U22022 (N_22022,N_15063,N_15818);
nor U22023 (N_22023,N_16102,N_13870);
nor U22024 (N_22024,N_16859,N_12422);
xor U22025 (N_22025,N_12356,N_14901);
xnor U22026 (N_22026,N_14684,N_15555);
xor U22027 (N_22027,N_16141,N_12762);
nand U22028 (N_22028,N_12073,N_15468);
or U22029 (N_22029,N_15705,N_16769);
or U22030 (N_22030,N_14251,N_17942);
nand U22031 (N_22031,N_14067,N_17028);
or U22032 (N_22032,N_12452,N_17823);
nor U22033 (N_22033,N_12865,N_12060);
xor U22034 (N_22034,N_12093,N_17840);
xor U22035 (N_22035,N_15466,N_12302);
or U22036 (N_22036,N_12229,N_12564);
xor U22037 (N_22037,N_13105,N_15454);
or U22038 (N_22038,N_14284,N_17985);
or U22039 (N_22039,N_12262,N_14745);
xor U22040 (N_22040,N_13275,N_14714);
and U22041 (N_22041,N_13252,N_14398);
nand U22042 (N_22042,N_14687,N_16521);
nand U22043 (N_22043,N_14580,N_12459);
nand U22044 (N_22044,N_16922,N_15455);
and U22045 (N_22045,N_17881,N_16280);
and U22046 (N_22046,N_17234,N_13379);
nand U22047 (N_22047,N_17185,N_13441);
xnor U22048 (N_22048,N_17651,N_13794);
and U22049 (N_22049,N_13486,N_16088);
nand U22050 (N_22050,N_12957,N_17558);
nand U22051 (N_22051,N_14453,N_16784);
or U22052 (N_22052,N_16720,N_16991);
nand U22053 (N_22053,N_13365,N_15855);
or U22054 (N_22054,N_13200,N_12144);
and U22055 (N_22055,N_15102,N_12709);
xnor U22056 (N_22056,N_17140,N_17603);
xor U22057 (N_22057,N_13678,N_16366);
nand U22058 (N_22058,N_12431,N_13739);
xnor U22059 (N_22059,N_14875,N_16127);
nand U22060 (N_22060,N_13511,N_17807);
and U22061 (N_22061,N_16366,N_16706);
nor U22062 (N_22062,N_13380,N_17299);
and U22063 (N_22063,N_12905,N_14375);
nand U22064 (N_22064,N_15281,N_17575);
and U22065 (N_22065,N_15520,N_12779);
and U22066 (N_22066,N_17117,N_17199);
xnor U22067 (N_22067,N_12070,N_17912);
nor U22068 (N_22068,N_15393,N_13428);
nor U22069 (N_22069,N_15815,N_12148);
xnor U22070 (N_22070,N_15601,N_12237);
nor U22071 (N_22071,N_17946,N_12218);
nand U22072 (N_22072,N_17528,N_14571);
nor U22073 (N_22073,N_16158,N_15342);
or U22074 (N_22074,N_15734,N_16876);
nand U22075 (N_22075,N_12982,N_16825);
xnor U22076 (N_22076,N_12278,N_13683);
xor U22077 (N_22077,N_12373,N_16553);
or U22078 (N_22078,N_17111,N_13655);
nand U22079 (N_22079,N_12394,N_12553);
nand U22080 (N_22080,N_13910,N_16902);
nor U22081 (N_22081,N_14558,N_16902);
or U22082 (N_22082,N_16838,N_13187);
and U22083 (N_22083,N_13917,N_17944);
nand U22084 (N_22084,N_17826,N_14842);
and U22085 (N_22085,N_17929,N_12040);
xor U22086 (N_22086,N_17351,N_13769);
nand U22087 (N_22087,N_12702,N_17634);
xor U22088 (N_22088,N_16400,N_17078);
and U22089 (N_22089,N_16710,N_12550);
nand U22090 (N_22090,N_16916,N_12351);
nand U22091 (N_22091,N_16384,N_15548);
and U22092 (N_22092,N_16542,N_16122);
and U22093 (N_22093,N_17879,N_13941);
or U22094 (N_22094,N_15881,N_16930);
nand U22095 (N_22095,N_16362,N_14863);
nor U22096 (N_22096,N_16081,N_16075);
and U22097 (N_22097,N_17185,N_16576);
xnor U22098 (N_22098,N_16517,N_13401);
or U22099 (N_22099,N_13216,N_17555);
or U22100 (N_22100,N_17076,N_16556);
or U22101 (N_22101,N_12825,N_12016);
nor U22102 (N_22102,N_15514,N_12049);
or U22103 (N_22103,N_13648,N_14809);
nor U22104 (N_22104,N_16853,N_14621);
nor U22105 (N_22105,N_16735,N_12311);
xnor U22106 (N_22106,N_14244,N_16987);
xor U22107 (N_22107,N_14941,N_15284);
nor U22108 (N_22108,N_14991,N_12453);
xnor U22109 (N_22109,N_15029,N_15943);
or U22110 (N_22110,N_16307,N_16718);
nor U22111 (N_22111,N_14257,N_17164);
xor U22112 (N_22112,N_12619,N_12395);
nor U22113 (N_22113,N_15309,N_15542);
xor U22114 (N_22114,N_13751,N_12117);
and U22115 (N_22115,N_13367,N_16560);
and U22116 (N_22116,N_12035,N_13414);
nor U22117 (N_22117,N_15434,N_13151);
or U22118 (N_22118,N_16660,N_16178);
nand U22119 (N_22119,N_13811,N_17103);
xnor U22120 (N_22120,N_15678,N_17930);
and U22121 (N_22121,N_16707,N_15030);
nand U22122 (N_22122,N_12790,N_14455);
xor U22123 (N_22123,N_16847,N_16515);
nor U22124 (N_22124,N_12733,N_17889);
nand U22125 (N_22125,N_13601,N_13443);
nand U22126 (N_22126,N_13835,N_12412);
nor U22127 (N_22127,N_16983,N_12623);
nand U22128 (N_22128,N_14210,N_13768);
nor U22129 (N_22129,N_14547,N_14416);
or U22130 (N_22130,N_12053,N_17989);
nand U22131 (N_22131,N_13384,N_13738);
or U22132 (N_22132,N_16640,N_15472);
xnor U22133 (N_22133,N_15118,N_12244);
and U22134 (N_22134,N_15790,N_16543);
nand U22135 (N_22135,N_12665,N_14059);
nand U22136 (N_22136,N_12986,N_12571);
nor U22137 (N_22137,N_17408,N_17877);
or U22138 (N_22138,N_14491,N_17273);
or U22139 (N_22139,N_12315,N_12328);
nor U22140 (N_22140,N_12734,N_12867);
or U22141 (N_22141,N_14154,N_12327);
xor U22142 (N_22142,N_14964,N_17706);
or U22143 (N_22143,N_17194,N_15367);
xnor U22144 (N_22144,N_14059,N_16578);
or U22145 (N_22145,N_17583,N_17699);
and U22146 (N_22146,N_17360,N_17262);
nor U22147 (N_22147,N_16014,N_13273);
xnor U22148 (N_22148,N_15578,N_12974);
nand U22149 (N_22149,N_17840,N_16258);
or U22150 (N_22150,N_14391,N_17958);
nor U22151 (N_22151,N_12549,N_14222);
xnor U22152 (N_22152,N_13366,N_15052);
xor U22153 (N_22153,N_15965,N_15430);
nor U22154 (N_22154,N_13249,N_15199);
xor U22155 (N_22155,N_12450,N_13635);
and U22156 (N_22156,N_16433,N_14307);
xor U22157 (N_22157,N_15733,N_12126);
nor U22158 (N_22158,N_12886,N_12345);
nand U22159 (N_22159,N_13343,N_14780);
nand U22160 (N_22160,N_12667,N_12747);
nand U22161 (N_22161,N_14804,N_17839);
xor U22162 (N_22162,N_14782,N_16225);
xor U22163 (N_22163,N_13716,N_12331);
nand U22164 (N_22164,N_16830,N_13727);
nor U22165 (N_22165,N_13646,N_13740);
nor U22166 (N_22166,N_12362,N_14047);
nor U22167 (N_22167,N_15196,N_12487);
xor U22168 (N_22168,N_15883,N_13520);
or U22169 (N_22169,N_15663,N_16601);
xor U22170 (N_22170,N_17251,N_17120);
nor U22171 (N_22171,N_14093,N_13106);
nand U22172 (N_22172,N_15625,N_15783);
xnor U22173 (N_22173,N_12252,N_14809);
and U22174 (N_22174,N_15645,N_12261);
nand U22175 (N_22175,N_12599,N_17575);
or U22176 (N_22176,N_13775,N_17216);
and U22177 (N_22177,N_14206,N_17549);
xnor U22178 (N_22178,N_16260,N_17076);
xnor U22179 (N_22179,N_16214,N_12946);
and U22180 (N_22180,N_17264,N_17626);
nand U22181 (N_22181,N_14053,N_12424);
nor U22182 (N_22182,N_17824,N_16412);
or U22183 (N_22183,N_12151,N_17402);
nand U22184 (N_22184,N_15207,N_13829);
nand U22185 (N_22185,N_15857,N_14401);
nor U22186 (N_22186,N_15044,N_17681);
nand U22187 (N_22187,N_17092,N_16979);
and U22188 (N_22188,N_13123,N_15370);
or U22189 (N_22189,N_13979,N_14315);
nand U22190 (N_22190,N_14177,N_16476);
nand U22191 (N_22191,N_16764,N_15538);
nor U22192 (N_22192,N_17059,N_12844);
nand U22193 (N_22193,N_15359,N_12307);
nand U22194 (N_22194,N_16829,N_17384);
and U22195 (N_22195,N_17356,N_12208);
or U22196 (N_22196,N_17253,N_13599);
or U22197 (N_22197,N_12571,N_12059);
nor U22198 (N_22198,N_16651,N_12213);
nand U22199 (N_22199,N_15524,N_17294);
and U22200 (N_22200,N_13847,N_14316);
or U22201 (N_22201,N_15724,N_14909);
or U22202 (N_22202,N_14912,N_15338);
or U22203 (N_22203,N_13381,N_16822);
or U22204 (N_22204,N_16975,N_14737);
xor U22205 (N_22205,N_14730,N_13823);
xor U22206 (N_22206,N_17520,N_16485);
and U22207 (N_22207,N_16440,N_16216);
nor U22208 (N_22208,N_12489,N_17414);
xor U22209 (N_22209,N_12546,N_13553);
xor U22210 (N_22210,N_12097,N_14482);
xnor U22211 (N_22211,N_17123,N_12019);
xor U22212 (N_22212,N_14830,N_14871);
xor U22213 (N_22213,N_15622,N_16096);
or U22214 (N_22214,N_16601,N_16129);
xor U22215 (N_22215,N_13819,N_14434);
or U22216 (N_22216,N_17415,N_12681);
or U22217 (N_22217,N_16367,N_14355);
and U22218 (N_22218,N_16694,N_14955);
nor U22219 (N_22219,N_16826,N_16397);
or U22220 (N_22220,N_12571,N_15962);
nor U22221 (N_22221,N_14796,N_14772);
xor U22222 (N_22222,N_15601,N_17873);
xor U22223 (N_22223,N_16616,N_13799);
and U22224 (N_22224,N_13740,N_16821);
nor U22225 (N_22225,N_12466,N_15096);
nand U22226 (N_22226,N_14030,N_13003);
or U22227 (N_22227,N_16267,N_14390);
nor U22228 (N_22228,N_15989,N_17070);
xnor U22229 (N_22229,N_12413,N_15490);
and U22230 (N_22230,N_14556,N_17956);
xnor U22231 (N_22231,N_12317,N_12762);
or U22232 (N_22232,N_15158,N_17493);
or U22233 (N_22233,N_16573,N_16504);
nor U22234 (N_22234,N_17186,N_12825);
and U22235 (N_22235,N_15392,N_13952);
or U22236 (N_22236,N_12928,N_15104);
nor U22237 (N_22237,N_14185,N_15373);
xor U22238 (N_22238,N_16287,N_13836);
nand U22239 (N_22239,N_12261,N_14513);
or U22240 (N_22240,N_12795,N_15395);
nand U22241 (N_22241,N_13051,N_12411);
xnor U22242 (N_22242,N_14006,N_12505);
or U22243 (N_22243,N_16991,N_13857);
or U22244 (N_22244,N_13420,N_16796);
nand U22245 (N_22245,N_12224,N_12160);
or U22246 (N_22246,N_12917,N_12276);
nor U22247 (N_22247,N_14703,N_13056);
nor U22248 (N_22248,N_16229,N_14987);
and U22249 (N_22249,N_17818,N_12457);
nor U22250 (N_22250,N_17594,N_15577);
and U22251 (N_22251,N_16081,N_13507);
and U22252 (N_22252,N_15333,N_14901);
nor U22253 (N_22253,N_14808,N_15807);
nand U22254 (N_22254,N_14574,N_16435);
xnor U22255 (N_22255,N_17331,N_15510);
or U22256 (N_22256,N_12247,N_12458);
xnor U22257 (N_22257,N_13988,N_17424);
or U22258 (N_22258,N_15205,N_13606);
nand U22259 (N_22259,N_13598,N_12738);
xnor U22260 (N_22260,N_17521,N_12342);
nor U22261 (N_22261,N_16809,N_15291);
xor U22262 (N_22262,N_14313,N_12121);
nand U22263 (N_22263,N_12131,N_15726);
or U22264 (N_22264,N_16867,N_12097);
and U22265 (N_22265,N_12970,N_17874);
nor U22266 (N_22266,N_16888,N_15482);
and U22267 (N_22267,N_13934,N_15326);
nor U22268 (N_22268,N_16544,N_12586);
nand U22269 (N_22269,N_17232,N_15839);
nor U22270 (N_22270,N_17571,N_13158);
nor U22271 (N_22271,N_17912,N_15276);
nor U22272 (N_22272,N_16184,N_12427);
xor U22273 (N_22273,N_14059,N_16667);
xnor U22274 (N_22274,N_12732,N_14733);
and U22275 (N_22275,N_16293,N_17513);
nor U22276 (N_22276,N_17418,N_14764);
nor U22277 (N_22277,N_15221,N_13649);
or U22278 (N_22278,N_16217,N_17414);
nor U22279 (N_22279,N_12730,N_16811);
and U22280 (N_22280,N_15566,N_17786);
or U22281 (N_22281,N_13505,N_15559);
nor U22282 (N_22282,N_17419,N_16627);
and U22283 (N_22283,N_16154,N_17339);
and U22284 (N_22284,N_15762,N_17578);
nand U22285 (N_22285,N_16092,N_14450);
xnor U22286 (N_22286,N_14974,N_15530);
xnor U22287 (N_22287,N_16645,N_12913);
nand U22288 (N_22288,N_17747,N_12746);
and U22289 (N_22289,N_17252,N_13596);
and U22290 (N_22290,N_16814,N_14498);
xnor U22291 (N_22291,N_13276,N_13105);
xnor U22292 (N_22292,N_15866,N_15666);
or U22293 (N_22293,N_17257,N_15296);
or U22294 (N_22294,N_17954,N_12305);
xor U22295 (N_22295,N_15603,N_16580);
nor U22296 (N_22296,N_15019,N_15858);
xnor U22297 (N_22297,N_12158,N_12424);
and U22298 (N_22298,N_12256,N_14484);
nor U22299 (N_22299,N_14187,N_16759);
nand U22300 (N_22300,N_12509,N_15222);
nor U22301 (N_22301,N_14208,N_13180);
and U22302 (N_22302,N_15826,N_14924);
and U22303 (N_22303,N_15102,N_13374);
or U22304 (N_22304,N_13079,N_16985);
or U22305 (N_22305,N_15933,N_15960);
or U22306 (N_22306,N_15107,N_13014);
xor U22307 (N_22307,N_17498,N_14529);
and U22308 (N_22308,N_16049,N_15642);
nor U22309 (N_22309,N_13421,N_14638);
nand U22310 (N_22310,N_15076,N_15784);
nor U22311 (N_22311,N_14183,N_16931);
xor U22312 (N_22312,N_16574,N_16278);
xnor U22313 (N_22313,N_14331,N_13652);
nor U22314 (N_22314,N_15747,N_14864);
nand U22315 (N_22315,N_13092,N_13113);
xnor U22316 (N_22316,N_14206,N_16577);
nand U22317 (N_22317,N_15630,N_12429);
and U22318 (N_22318,N_12253,N_13784);
nor U22319 (N_22319,N_14603,N_14752);
nor U22320 (N_22320,N_13269,N_14551);
and U22321 (N_22321,N_12527,N_13014);
nor U22322 (N_22322,N_16692,N_17172);
xnor U22323 (N_22323,N_14571,N_14919);
and U22324 (N_22324,N_15088,N_17388);
nor U22325 (N_22325,N_16952,N_16991);
and U22326 (N_22326,N_16300,N_17064);
nand U22327 (N_22327,N_17936,N_16087);
or U22328 (N_22328,N_15355,N_12224);
or U22329 (N_22329,N_12531,N_13649);
and U22330 (N_22330,N_17685,N_13207);
nand U22331 (N_22331,N_17069,N_17107);
and U22332 (N_22332,N_16165,N_14450);
xor U22333 (N_22333,N_15935,N_16811);
xor U22334 (N_22334,N_17863,N_12080);
xnor U22335 (N_22335,N_16222,N_14566);
nand U22336 (N_22336,N_15763,N_17794);
xor U22337 (N_22337,N_16254,N_12253);
xnor U22338 (N_22338,N_17097,N_17214);
and U22339 (N_22339,N_17359,N_14548);
nor U22340 (N_22340,N_16145,N_12074);
nand U22341 (N_22341,N_14012,N_15526);
nand U22342 (N_22342,N_12534,N_12873);
nand U22343 (N_22343,N_15056,N_16070);
nor U22344 (N_22344,N_14396,N_15723);
nor U22345 (N_22345,N_12719,N_17768);
or U22346 (N_22346,N_13076,N_12999);
nor U22347 (N_22347,N_17207,N_17130);
and U22348 (N_22348,N_14030,N_17628);
nor U22349 (N_22349,N_16368,N_14662);
xnor U22350 (N_22350,N_13736,N_14849);
or U22351 (N_22351,N_14695,N_14080);
and U22352 (N_22352,N_14656,N_13018);
or U22353 (N_22353,N_14751,N_16067);
nand U22354 (N_22354,N_16800,N_12910);
or U22355 (N_22355,N_16604,N_13891);
and U22356 (N_22356,N_15145,N_17039);
nor U22357 (N_22357,N_13739,N_15521);
or U22358 (N_22358,N_13753,N_12812);
nor U22359 (N_22359,N_17990,N_17482);
nor U22360 (N_22360,N_14207,N_16955);
or U22361 (N_22361,N_15118,N_16870);
or U22362 (N_22362,N_16407,N_13860);
xor U22363 (N_22363,N_17887,N_13995);
nand U22364 (N_22364,N_14287,N_15387);
or U22365 (N_22365,N_12392,N_15601);
and U22366 (N_22366,N_13264,N_13197);
or U22367 (N_22367,N_17339,N_16626);
xnor U22368 (N_22368,N_15491,N_16234);
and U22369 (N_22369,N_16767,N_13483);
nand U22370 (N_22370,N_15812,N_12643);
and U22371 (N_22371,N_17049,N_16155);
nand U22372 (N_22372,N_15618,N_15490);
nor U22373 (N_22373,N_16008,N_17805);
nor U22374 (N_22374,N_12543,N_15805);
nor U22375 (N_22375,N_17833,N_14765);
or U22376 (N_22376,N_15013,N_14325);
and U22377 (N_22377,N_15982,N_15110);
and U22378 (N_22378,N_14763,N_16177);
or U22379 (N_22379,N_12344,N_16581);
or U22380 (N_22380,N_17536,N_12808);
or U22381 (N_22381,N_13477,N_17094);
xnor U22382 (N_22382,N_16996,N_16354);
and U22383 (N_22383,N_13748,N_14258);
nor U22384 (N_22384,N_17745,N_15299);
nand U22385 (N_22385,N_16869,N_13623);
nand U22386 (N_22386,N_12958,N_15280);
nand U22387 (N_22387,N_15347,N_12861);
xnor U22388 (N_22388,N_14309,N_14302);
nand U22389 (N_22389,N_12257,N_17669);
xor U22390 (N_22390,N_16504,N_14628);
or U22391 (N_22391,N_13413,N_12812);
or U22392 (N_22392,N_16340,N_13154);
and U22393 (N_22393,N_13309,N_15273);
xor U22394 (N_22394,N_17316,N_17313);
nor U22395 (N_22395,N_14291,N_12315);
xnor U22396 (N_22396,N_13278,N_15805);
and U22397 (N_22397,N_16782,N_14180);
or U22398 (N_22398,N_15887,N_16242);
or U22399 (N_22399,N_16905,N_17170);
or U22400 (N_22400,N_17394,N_12361);
nand U22401 (N_22401,N_13200,N_15970);
xor U22402 (N_22402,N_16515,N_13089);
nor U22403 (N_22403,N_13129,N_13412);
nor U22404 (N_22404,N_17886,N_16283);
xnor U22405 (N_22405,N_13831,N_14042);
xnor U22406 (N_22406,N_12676,N_15204);
or U22407 (N_22407,N_14675,N_15077);
nand U22408 (N_22408,N_17964,N_14728);
nor U22409 (N_22409,N_15204,N_14234);
nand U22410 (N_22410,N_15027,N_12391);
and U22411 (N_22411,N_17096,N_16836);
nand U22412 (N_22412,N_14338,N_17566);
nor U22413 (N_22413,N_17966,N_15130);
or U22414 (N_22414,N_13487,N_12885);
nand U22415 (N_22415,N_15375,N_17885);
nand U22416 (N_22416,N_12954,N_15965);
nor U22417 (N_22417,N_16079,N_14555);
or U22418 (N_22418,N_15435,N_13329);
and U22419 (N_22419,N_14140,N_15295);
nor U22420 (N_22420,N_13330,N_16107);
nand U22421 (N_22421,N_13670,N_16914);
nand U22422 (N_22422,N_17596,N_14211);
nand U22423 (N_22423,N_17584,N_15849);
or U22424 (N_22424,N_14372,N_13209);
nand U22425 (N_22425,N_17231,N_17249);
or U22426 (N_22426,N_15423,N_15909);
xnor U22427 (N_22427,N_13151,N_17676);
nor U22428 (N_22428,N_15644,N_17860);
nand U22429 (N_22429,N_15871,N_14827);
nand U22430 (N_22430,N_12952,N_14083);
xor U22431 (N_22431,N_15474,N_17734);
nand U22432 (N_22432,N_15068,N_17013);
xnor U22433 (N_22433,N_16214,N_12034);
xor U22434 (N_22434,N_15959,N_13634);
xnor U22435 (N_22435,N_13235,N_14474);
nand U22436 (N_22436,N_15241,N_13001);
nand U22437 (N_22437,N_15770,N_16167);
nor U22438 (N_22438,N_14618,N_17792);
nor U22439 (N_22439,N_15520,N_16855);
and U22440 (N_22440,N_12201,N_15870);
nand U22441 (N_22441,N_14405,N_14721);
nand U22442 (N_22442,N_12337,N_17299);
xor U22443 (N_22443,N_17844,N_13136);
nand U22444 (N_22444,N_16677,N_16418);
xor U22445 (N_22445,N_15566,N_16410);
nand U22446 (N_22446,N_14208,N_16698);
or U22447 (N_22447,N_15302,N_15888);
nand U22448 (N_22448,N_14160,N_14277);
or U22449 (N_22449,N_12451,N_15871);
or U22450 (N_22450,N_16806,N_15405);
nor U22451 (N_22451,N_15840,N_15749);
nor U22452 (N_22452,N_14637,N_17004);
or U22453 (N_22453,N_16890,N_17893);
xnor U22454 (N_22454,N_16848,N_16262);
or U22455 (N_22455,N_14470,N_14514);
xor U22456 (N_22456,N_15746,N_16779);
xor U22457 (N_22457,N_12505,N_17038);
nand U22458 (N_22458,N_12502,N_16141);
xnor U22459 (N_22459,N_17875,N_14984);
and U22460 (N_22460,N_12667,N_16255);
and U22461 (N_22461,N_16853,N_15050);
xor U22462 (N_22462,N_13348,N_17788);
or U22463 (N_22463,N_15153,N_17921);
nor U22464 (N_22464,N_16536,N_14384);
and U22465 (N_22465,N_17962,N_16243);
and U22466 (N_22466,N_12316,N_14079);
or U22467 (N_22467,N_16574,N_16453);
nand U22468 (N_22468,N_16326,N_12259);
nor U22469 (N_22469,N_13852,N_12321);
and U22470 (N_22470,N_14286,N_14110);
nor U22471 (N_22471,N_16819,N_12222);
xnor U22472 (N_22472,N_15464,N_12578);
nor U22473 (N_22473,N_15499,N_12036);
xor U22474 (N_22474,N_13586,N_15557);
nand U22475 (N_22475,N_14138,N_14528);
nand U22476 (N_22476,N_12045,N_12900);
or U22477 (N_22477,N_16332,N_17200);
or U22478 (N_22478,N_15905,N_14412);
xor U22479 (N_22479,N_12716,N_12469);
and U22480 (N_22480,N_14257,N_14303);
xnor U22481 (N_22481,N_13024,N_16118);
xor U22482 (N_22482,N_13563,N_14930);
nand U22483 (N_22483,N_17672,N_12710);
nand U22484 (N_22484,N_17032,N_13512);
xnor U22485 (N_22485,N_16833,N_12946);
nand U22486 (N_22486,N_17556,N_17066);
and U22487 (N_22487,N_16057,N_14150);
and U22488 (N_22488,N_15077,N_16554);
nor U22489 (N_22489,N_17562,N_15951);
nand U22490 (N_22490,N_17247,N_13464);
nor U22491 (N_22491,N_17588,N_15898);
nor U22492 (N_22492,N_16942,N_17397);
or U22493 (N_22493,N_13186,N_15811);
and U22494 (N_22494,N_12339,N_17339);
or U22495 (N_22495,N_14731,N_13147);
nand U22496 (N_22496,N_14983,N_13846);
xor U22497 (N_22497,N_13242,N_16471);
nand U22498 (N_22498,N_15540,N_17069);
nor U22499 (N_22499,N_12225,N_12339);
nand U22500 (N_22500,N_14565,N_13547);
and U22501 (N_22501,N_16224,N_17911);
nand U22502 (N_22502,N_15871,N_14816);
and U22503 (N_22503,N_16715,N_15978);
and U22504 (N_22504,N_14215,N_13929);
nand U22505 (N_22505,N_12666,N_13476);
or U22506 (N_22506,N_15735,N_14112);
xor U22507 (N_22507,N_17976,N_14873);
or U22508 (N_22508,N_16058,N_17488);
nor U22509 (N_22509,N_15905,N_16837);
and U22510 (N_22510,N_15581,N_15234);
nor U22511 (N_22511,N_17298,N_12414);
xor U22512 (N_22512,N_16816,N_12091);
nand U22513 (N_22513,N_17782,N_15093);
or U22514 (N_22514,N_13133,N_17030);
nand U22515 (N_22515,N_12282,N_12227);
nor U22516 (N_22516,N_15377,N_12237);
nor U22517 (N_22517,N_15049,N_14704);
or U22518 (N_22518,N_14980,N_13975);
nand U22519 (N_22519,N_16666,N_12618);
xor U22520 (N_22520,N_12966,N_14539);
and U22521 (N_22521,N_15572,N_14431);
nand U22522 (N_22522,N_15869,N_14563);
xnor U22523 (N_22523,N_15197,N_13432);
xnor U22524 (N_22524,N_16019,N_15951);
nor U22525 (N_22525,N_17201,N_13850);
xnor U22526 (N_22526,N_17208,N_15608);
xor U22527 (N_22527,N_16417,N_17192);
or U22528 (N_22528,N_12015,N_15188);
and U22529 (N_22529,N_12958,N_14376);
or U22530 (N_22530,N_17759,N_14500);
and U22531 (N_22531,N_15228,N_15358);
nor U22532 (N_22532,N_16996,N_17499);
nand U22533 (N_22533,N_15290,N_17206);
and U22534 (N_22534,N_16531,N_13813);
nor U22535 (N_22535,N_13833,N_17428);
xnor U22536 (N_22536,N_16536,N_13019);
and U22537 (N_22537,N_14439,N_13406);
nor U22538 (N_22538,N_16228,N_16520);
nand U22539 (N_22539,N_17302,N_15299);
nor U22540 (N_22540,N_13656,N_15974);
or U22541 (N_22541,N_16462,N_14870);
nand U22542 (N_22542,N_14499,N_14376);
nand U22543 (N_22543,N_15085,N_17829);
xor U22544 (N_22544,N_17985,N_17152);
nor U22545 (N_22545,N_15569,N_17670);
and U22546 (N_22546,N_12412,N_13140);
nor U22547 (N_22547,N_14425,N_16934);
and U22548 (N_22548,N_14709,N_14078);
nand U22549 (N_22549,N_12800,N_13404);
nor U22550 (N_22550,N_14969,N_12236);
xor U22551 (N_22551,N_12098,N_14735);
nand U22552 (N_22552,N_13493,N_16987);
nor U22553 (N_22553,N_17398,N_13898);
nand U22554 (N_22554,N_16335,N_17279);
nor U22555 (N_22555,N_16793,N_16804);
or U22556 (N_22556,N_12517,N_16048);
or U22557 (N_22557,N_17204,N_15712);
or U22558 (N_22558,N_12663,N_16266);
and U22559 (N_22559,N_15834,N_15580);
or U22560 (N_22560,N_12358,N_12874);
xnor U22561 (N_22561,N_12551,N_12160);
and U22562 (N_22562,N_13474,N_17069);
or U22563 (N_22563,N_14276,N_12841);
nand U22564 (N_22564,N_15459,N_14560);
or U22565 (N_22565,N_14012,N_16176);
nor U22566 (N_22566,N_14194,N_15878);
xnor U22567 (N_22567,N_17601,N_16020);
or U22568 (N_22568,N_15776,N_14654);
nand U22569 (N_22569,N_12549,N_15430);
or U22570 (N_22570,N_12928,N_16020);
nor U22571 (N_22571,N_14393,N_15543);
xor U22572 (N_22572,N_17812,N_17395);
and U22573 (N_22573,N_14787,N_12409);
nand U22574 (N_22574,N_17651,N_14575);
and U22575 (N_22575,N_12667,N_13308);
nand U22576 (N_22576,N_14916,N_16225);
or U22577 (N_22577,N_14146,N_15876);
nor U22578 (N_22578,N_15411,N_14717);
xnor U22579 (N_22579,N_13766,N_17831);
nand U22580 (N_22580,N_13094,N_12845);
and U22581 (N_22581,N_15776,N_16397);
nand U22582 (N_22582,N_17485,N_14214);
and U22583 (N_22583,N_12195,N_15508);
nor U22584 (N_22584,N_15618,N_17008);
nand U22585 (N_22585,N_13736,N_15091);
or U22586 (N_22586,N_17820,N_13279);
nor U22587 (N_22587,N_13773,N_15396);
nand U22588 (N_22588,N_17313,N_13881);
nand U22589 (N_22589,N_14647,N_12077);
xor U22590 (N_22590,N_14404,N_16871);
and U22591 (N_22591,N_12549,N_15553);
xnor U22592 (N_22592,N_12280,N_12863);
or U22593 (N_22593,N_15660,N_13405);
nand U22594 (N_22594,N_15750,N_14526);
xnor U22595 (N_22595,N_14854,N_17042);
and U22596 (N_22596,N_15690,N_14903);
nor U22597 (N_22597,N_15034,N_15230);
and U22598 (N_22598,N_14909,N_13523);
or U22599 (N_22599,N_15603,N_13610);
and U22600 (N_22600,N_14156,N_16087);
nand U22601 (N_22601,N_14328,N_15781);
or U22602 (N_22602,N_15902,N_17703);
nor U22603 (N_22603,N_15325,N_13341);
or U22604 (N_22604,N_13079,N_17599);
nor U22605 (N_22605,N_17670,N_16261);
nor U22606 (N_22606,N_15411,N_14292);
nand U22607 (N_22607,N_16892,N_17603);
nor U22608 (N_22608,N_15573,N_12261);
nor U22609 (N_22609,N_15288,N_13220);
nor U22610 (N_22610,N_12484,N_16080);
nand U22611 (N_22611,N_14367,N_17474);
xor U22612 (N_22612,N_17063,N_13484);
or U22613 (N_22613,N_15840,N_17953);
or U22614 (N_22614,N_14410,N_15949);
nand U22615 (N_22615,N_17502,N_17572);
and U22616 (N_22616,N_12176,N_16494);
nor U22617 (N_22617,N_17834,N_12981);
nand U22618 (N_22618,N_15390,N_13633);
nand U22619 (N_22619,N_14604,N_16833);
or U22620 (N_22620,N_14999,N_14390);
or U22621 (N_22621,N_16242,N_17986);
nor U22622 (N_22622,N_12710,N_12074);
xor U22623 (N_22623,N_15529,N_12901);
nor U22624 (N_22624,N_12452,N_13753);
nor U22625 (N_22625,N_14438,N_16066);
nor U22626 (N_22626,N_16271,N_12306);
and U22627 (N_22627,N_17450,N_14272);
or U22628 (N_22628,N_12312,N_13293);
or U22629 (N_22629,N_14359,N_17002);
nand U22630 (N_22630,N_12449,N_14181);
nor U22631 (N_22631,N_15483,N_13757);
nor U22632 (N_22632,N_12961,N_13852);
and U22633 (N_22633,N_13146,N_17789);
or U22634 (N_22634,N_17562,N_16970);
nor U22635 (N_22635,N_16551,N_12180);
or U22636 (N_22636,N_15293,N_13216);
xnor U22637 (N_22637,N_15025,N_14797);
nand U22638 (N_22638,N_13815,N_15414);
or U22639 (N_22639,N_14387,N_13786);
or U22640 (N_22640,N_13718,N_17082);
and U22641 (N_22641,N_15575,N_16425);
and U22642 (N_22642,N_15189,N_15872);
nor U22643 (N_22643,N_15472,N_17510);
or U22644 (N_22644,N_12213,N_16634);
nand U22645 (N_22645,N_14100,N_16553);
xor U22646 (N_22646,N_12514,N_17521);
nand U22647 (N_22647,N_12944,N_17327);
and U22648 (N_22648,N_15581,N_16439);
xnor U22649 (N_22649,N_14434,N_15064);
xnor U22650 (N_22650,N_15896,N_16849);
xnor U22651 (N_22651,N_13327,N_14680);
or U22652 (N_22652,N_16313,N_16357);
or U22653 (N_22653,N_13156,N_12635);
or U22654 (N_22654,N_12833,N_16235);
or U22655 (N_22655,N_17180,N_14393);
or U22656 (N_22656,N_17515,N_15009);
nand U22657 (N_22657,N_16327,N_12990);
nand U22658 (N_22658,N_17378,N_16254);
and U22659 (N_22659,N_14324,N_15807);
nor U22660 (N_22660,N_16066,N_13588);
nor U22661 (N_22661,N_15264,N_15875);
nor U22662 (N_22662,N_17099,N_12188);
nand U22663 (N_22663,N_17930,N_16956);
nor U22664 (N_22664,N_17062,N_14228);
nand U22665 (N_22665,N_14042,N_16736);
and U22666 (N_22666,N_16043,N_16032);
nand U22667 (N_22667,N_14536,N_15210);
xnor U22668 (N_22668,N_13978,N_17847);
or U22669 (N_22669,N_13190,N_12913);
nor U22670 (N_22670,N_16903,N_13347);
nor U22671 (N_22671,N_14297,N_16054);
and U22672 (N_22672,N_15416,N_16123);
or U22673 (N_22673,N_17889,N_16478);
nor U22674 (N_22674,N_16500,N_15656);
xor U22675 (N_22675,N_16558,N_17770);
xnor U22676 (N_22676,N_17537,N_17086);
nand U22677 (N_22677,N_16346,N_16731);
xnor U22678 (N_22678,N_16983,N_12824);
and U22679 (N_22679,N_13029,N_14089);
xnor U22680 (N_22680,N_12114,N_15618);
or U22681 (N_22681,N_12688,N_12829);
nand U22682 (N_22682,N_14638,N_14595);
or U22683 (N_22683,N_12537,N_17248);
and U22684 (N_22684,N_16595,N_15539);
nor U22685 (N_22685,N_13706,N_16691);
and U22686 (N_22686,N_13524,N_13889);
xor U22687 (N_22687,N_12135,N_13580);
xnor U22688 (N_22688,N_17674,N_13686);
nor U22689 (N_22689,N_17540,N_16896);
xnor U22690 (N_22690,N_12887,N_17125);
and U22691 (N_22691,N_12038,N_17127);
and U22692 (N_22692,N_15170,N_17517);
nor U22693 (N_22693,N_17301,N_13701);
or U22694 (N_22694,N_17175,N_14612);
nor U22695 (N_22695,N_16777,N_14930);
nor U22696 (N_22696,N_15647,N_13205);
or U22697 (N_22697,N_13206,N_14321);
nand U22698 (N_22698,N_16374,N_16458);
nor U22699 (N_22699,N_16385,N_16377);
or U22700 (N_22700,N_17510,N_16339);
and U22701 (N_22701,N_14632,N_14188);
and U22702 (N_22702,N_16091,N_14140);
and U22703 (N_22703,N_17363,N_13192);
or U22704 (N_22704,N_16782,N_15033);
nand U22705 (N_22705,N_14536,N_13906);
and U22706 (N_22706,N_13475,N_12836);
and U22707 (N_22707,N_17745,N_14686);
nor U22708 (N_22708,N_16710,N_14095);
and U22709 (N_22709,N_14432,N_13398);
and U22710 (N_22710,N_15587,N_17392);
nor U22711 (N_22711,N_14134,N_15922);
and U22712 (N_22712,N_14913,N_16038);
and U22713 (N_22713,N_16958,N_14031);
nor U22714 (N_22714,N_13695,N_13512);
nor U22715 (N_22715,N_16695,N_15775);
xor U22716 (N_22716,N_16487,N_16244);
and U22717 (N_22717,N_17265,N_14547);
xnor U22718 (N_22718,N_16845,N_17639);
nor U22719 (N_22719,N_14452,N_14308);
nand U22720 (N_22720,N_16931,N_13950);
nor U22721 (N_22721,N_15818,N_12750);
or U22722 (N_22722,N_16139,N_15521);
nand U22723 (N_22723,N_14375,N_16684);
nand U22724 (N_22724,N_17055,N_17418);
nand U22725 (N_22725,N_14551,N_12365);
nand U22726 (N_22726,N_13218,N_15121);
or U22727 (N_22727,N_14902,N_16698);
or U22728 (N_22728,N_17881,N_13240);
xnor U22729 (N_22729,N_15449,N_15210);
or U22730 (N_22730,N_13556,N_14169);
and U22731 (N_22731,N_13709,N_13319);
and U22732 (N_22732,N_13775,N_14617);
xnor U22733 (N_22733,N_12697,N_15187);
and U22734 (N_22734,N_16626,N_12209);
and U22735 (N_22735,N_16981,N_14780);
xor U22736 (N_22736,N_13076,N_12682);
xnor U22737 (N_22737,N_13497,N_15678);
or U22738 (N_22738,N_12401,N_15105);
xor U22739 (N_22739,N_14146,N_17145);
and U22740 (N_22740,N_15329,N_16855);
nor U22741 (N_22741,N_13269,N_15538);
nand U22742 (N_22742,N_14706,N_12870);
and U22743 (N_22743,N_16222,N_12696);
and U22744 (N_22744,N_17259,N_17307);
nand U22745 (N_22745,N_13763,N_15879);
xor U22746 (N_22746,N_15400,N_15302);
xnor U22747 (N_22747,N_12323,N_14358);
or U22748 (N_22748,N_12582,N_12477);
nand U22749 (N_22749,N_12768,N_16672);
and U22750 (N_22750,N_17458,N_13941);
or U22751 (N_22751,N_16855,N_12035);
nor U22752 (N_22752,N_15322,N_17117);
xor U22753 (N_22753,N_12409,N_12528);
xor U22754 (N_22754,N_17696,N_15150);
nand U22755 (N_22755,N_13911,N_13612);
or U22756 (N_22756,N_15584,N_15185);
nand U22757 (N_22757,N_16708,N_12460);
nor U22758 (N_22758,N_14346,N_13504);
nand U22759 (N_22759,N_13135,N_13872);
or U22760 (N_22760,N_14953,N_17123);
and U22761 (N_22761,N_16460,N_14753);
or U22762 (N_22762,N_15447,N_16263);
and U22763 (N_22763,N_16887,N_15929);
nand U22764 (N_22764,N_13282,N_12774);
and U22765 (N_22765,N_12074,N_17366);
or U22766 (N_22766,N_14070,N_13013);
or U22767 (N_22767,N_14567,N_15489);
or U22768 (N_22768,N_13241,N_13708);
and U22769 (N_22769,N_13768,N_17267);
or U22770 (N_22770,N_13203,N_13916);
nor U22771 (N_22771,N_15036,N_17890);
nor U22772 (N_22772,N_15095,N_15891);
nor U22773 (N_22773,N_12279,N_12867);
and U22774 (N_22774,N_16424,N_12660);
nor U22775 (N_22775,N_17400,N_16097);
or U22776 (N_22776,N_17652,N_16029);
and U22777 (N_22777,N_17515,N_13672);
nor U22778 (N_22778,N_17312,N_13083);
xor U22779 (N_22779,N_15354,N_13112);
or U22780 (N_22780,N_13669,N_16098);
and U22781 (N_22781,N_15156,N_14221);
nor U22782 (N_22782,N_12232,N_17270);
nor U22783 (N_22783,N_12886,N_13069);
nand U22784 (N_22784,N_12582,N_14929);
and U22785 (N_22785,N_16101,N_13493);
nor U22786 (N_22786,N_15421,N_13205);
nor U22787 (N_22787,N_14824,N_14923);
and U22788 (N_22788,N_12560,N_12440);
or U22789 (N_22789,N_15038,N_14085);
or U22790 (N_22790,N_16177,N_13618);
and U22791 (N_22791,N_12525,N_14006);
nor U22792 (N_22792,N_13153,N_12608);
nand U22793 (N_22793,N_13417,N_14465);
nand U22794 (N_22794,N_13369,N_16477);
and U22795 (N_22795,N_15168,N_15482);
or U22796 (N_22796,N_16865,N_13130);
nor U22797 (N_22797,N_17457,N_15571);
nor U22798 (N_22798,N_14707,N_14957);
or U22799 (N_22799,N_14812,N_12733);
nand U22800 (N_22800,N_13381,N_15860);
xor U22801 (N_22801,N_12339,N_14561);
and U22802 (N_22802,N_16798,N_16423);
or U22803 (N_22803,N_15893,N_13642);
nor U22804 (N_22804,N_16551,N_13619);
xor U22805 (N_22805,N_17205,N_14376);
nor U22806 (N_22806,N_15181,N_12727);
nor U22807 (N_22807,N_13651,N_12293);
nor U22808 (N_22808,N_12289,N_13196);
nor U22809 (N_22809,N_13780,N_12047);
nand U22810 (N_22810,N_12950,N_12114);
nor U22811 (N_22811,N_17531,N_15952);
and U22812 (N_22812,N_15079,N_15017);
and U22813 (N_22813,N_15856,N_14198);
or U22814 (N_22814,N_16083,N_15290);
and U22815 (N_22815,N_15548,N_13846);
nand U22816 (N_22816,N_13685,N_13139);
nor U22817 (N_22817,N_13435,N_17997);
nand U22818 (N_22818,N_14187,N_16822);
nor U22819 (N_22819,N_14588,N_13278);
nor U22820 (N_22820,N_12042,N_17700);
nand U22821 (N_22821,N_15892,N_12602);
nor U22822 (N_22822,N_17281,N_16247);
and U22823 (N_22823,N_13026,N_16036);
nor U22824 (N_22824,N_17287,N_13810);
nand U22825 (N_22825,N_12562,N_15397);
and U22826 (N_22826,N_17815,N_17536);
and U22827 (N_22827,N_13817,N_16169);
nor U22828 (N_22828,N_16518,N_16567);
nor U22829 (N_22829,N_13751,N_14730);
nor U22830 (N_22830,N_17572,N_15678);
and U22831 (N_22831,N_12900,N_17589);
nor U22832 (N_22832,N_12869,N_14738);
xor U22833 (N_22833,N_16995,N_16404);
xnor U22834 (N_22834,N_15591,N_16916);
nor U22835 (N_22835,N_17822,N_14801);
nor U22836 (N_22836,N_14070,N_16876);
nor U22837 (N_22837,N_13654,N_14932);
or U22838 (N_22838,N_12743,N_16694);
and U22839 (N_22839,N_16134,N_12604);
xor U22840 (N_22840,N_15005,N_14083);
and U22841 (N_22841,N_17980,N_15073);
xor U22842 (N_22842,N_17136,N_15439);
and U22843 (N_22843,N_17111,N_12530);
nand U22844 (N_22844,N_14906,N_16337);
or U22845 (N_22845,N_13421,N_16037);
nand U22846 (N_22846,N_13141,N_15466);
nor U22847 (N_22847,N_12365,N_16370);
and U22848 (N_22848,N_12555,N_14767);
and U22849 (N_22849,N_12621,N_12216);
or U22850 (N_22850,N_17626,N_12207);
and U22851 (N_22851,N_12165,N_16500);
xor U22852 (N_22852,N_14598,N_16634);
nor U22853 (N_22853,N_13754,N_13148);
and U22854 (N_22854,N_13827,N_13611);
nor U22855 (N_22855,N_13818,N_17795);
xnor U22856 (N_22856,N_13280,N_14751);
or U22857 (N_22857,N_15029,N_13653);
xor U22858 (N_22858,N_16973,N_13203);
or U22859 (N_22859,N_12620,N_15285);
xnor U22860 (N_22860,N_13835,N_16043);
and U22861 (N_22861,N_13820,N_13576);
and U22862 (N_22862,N_12029,N_14463);
xor U22863 (N_22863,N_17330,N_17724);
or U22864 (N_22864,N_12493,N_14539);
or U22865 (N_22865,N_17972,N_12466);
nor U22866 (N_22866,N_17989,N_13749);
nor U22867 (N_22867,N_12457,N_15712);
xnor U22868 (N_22868,N_16988,N_14220);
xnor U22869 (N_22869,N_12068,N_16640);
xnor U22870 (N_22870,N_12813,N_17294);
nor U22871 (N_22871,N_15641,N_17336);
xor U22872 (N_22872,N_13181,N_14214);
nor U22873 (N_22873,N_14827,N_16564);
and U22874 (N_22874,N_14896,N_16591);
nand U22875 (N_22875,N_14090,N_17436);
or U22876 (N_22876,N_17572,N_16163);
xnor U22877 (N_22877,N_15851,N_16378);
xnor U22878 (N_22878,N_13793,N_12385);
and U22879 (N_22879,N_12649,N_16421);
and U22880 (N_22880,N_13694,N_15275);
nor U22881 (N_22881,N_12686,N_12158);
xnor U22882 (N_22882,N_15559,N_14401);
nor U22883 (N_22883,N_17661,N_14634);
and U22884 (N_22884,N_13395,N_16241);
nor U22885 (N_22885,N_12555,N_14226);
nand U22886 (N_22886,N_17674,N_16232);
and U22887 (N_22887,N_16162,N_12531);
and U22888 (N_22888,N_14002,N_16236);
nand U22889 (N_22889,N_14043,N_13868);
and U22890 (N_22890,N_13557,N_14402);
or U22891 (N_22891,N_15672,N_17305);
and U22892 (N_22892,N_16799,N_15763);
nor U22893 (N_22893,N_16111,N_16530);
or U22894 (N_22894,N_13704,N_14030);
nand U22895 (N_22895,N_14997,N_12019);
xor U22896 (N_22896,N_17164,N_15184);
xnor U22897 (N_22897,N_16416,N_13982);
nand U22898 (N_22898,N_13529,N_13275);
nor U22899 (N_22899,N_14817,N_13085);
and U22900 (N_22900,N_15075,N_16161);
xor U22901 (N_22901,N_14344,N_16808);
or U22902 (N_22902,N_12228,N_12242);
or U22903 (N_22903,N_15213,N_17118);
nor U22904 (N_22904,N_13513,N_15093);
or U22905 (N_22905,N_14092,N_12177);
or U22906 (N_22906,N_14636,N_15651);
or U22907 (N_22907,N_13074,N_15208);
nor U22908 (N_22908,N_15257,N_12100);
nand U22909 (N_22909,N_14661,N_12485);
or U22910 (N_22910,N_17777,N_12582);
nor U22911 (N_22911,N_12923,N_12771);
xnor U22912 (N_22912,N_14919,N_13493);
or U22913 (N_22913,N_15119,N_16216);
nor U22914 (N_22914,N_17303,N_13097);
nand U22915 (N_22915,N_14713,N_13150);
xnor U22916 (N_22916,N_14747,N_12696);
and U22917 (N_22917,N_16638,N_15078);
nor U22918 (N_22918,N_12714,N_14503);
and U22919 (N_22919,N_15677,N_15436);
xor U22920 (N_22920,N_13197,N_12211);
or U22921 (N_22921,N_12986,N_13504);
nand U22922 (N_22922,N_17795,N_16845);
xnor U22923 (N_22923,N_12763,N_17184);
nor U22924 (N_22924,N_15768,N_15034);
nor U22925 (N_22925,N_16079,N_17473);
and U22926 (N_22926,N_17407,N_13705);
nand U22927 (N_22927,N_14019,N_12354);
and U22928 (N_22928,N_15185,N_15191);
nor U22929 (N_22929,N_16249,N_12694);
nor U22930 (N_22930,N_15763,N_12179);
nor U22931 (N_22931,N_15250,N_17827);
or U22932 (N_22932,N_12035,N_12134);
or U22933 (N_22933,N_12667,N_17491);
nand U22934 (N_22934,N_14006,N_17894);
xor U22935 (N_22935,N_16863,N_14261);
or U22936 (N_22936,N_15337,N_16292);
nand U22937 (N_22937,N_13061,N_13278);
or U22938 (N_22938,N_15072,N_12543);
xnor U22939 (N_22939,N_12254,N_12830);
nor U22940 (N_22940,N_12517,N_13665);
and U22941 (N_22941,N_17828,N_13716);
nand U22942 (N_22942,N_16989,N_12605);
or U22943 (N_22943,N_12709,N_16290);
and U22944 (N_22944,N_12734,N_17020);
or U22945 (N_22945,N_13397,N_12170);
and U22946 (N_22946,N_17638,N_12859);
xnor U22947 (N_22947,N_16227,N_17781);
or U22948 (N_22948,N_12680,N_15389);
nor U22949 (N_22949,N_14156,N_16498);
and U22950 (N_22950,N_13058,N_17220);
xnor U22951 (N_22951,N_13296,N_12617);
or U22952 (N_22952,N_12825,N_14137);
or U22953 (N_22953,N_16387,N_13300);
nor U22954 (N_22954,N_15123,N_17431);
and U22955 (N_22955,N_17655,N_16534);
xnor U22956 (N_22956,N_13373,N_14749);
xnor U22957 (N_22957,N_14600,N_15326);
or U22958 (N_22958,N_17911,N_15410);
or U22959 (N_22959,N_17188,N_15031);
or U22960 (N_22960,N_17838,N_12688);
nand U22961 (N_22961,N_12513,N_15436);
and U22962 (N_22962,N_17540,N_17515);
xor U22963 (N_22963,N_17706,N_12931);
nand U22964 (N_22964,N_14992,N_13508);
nor U22965 (N_22965,N_15798,N_17167);
nor U22966 (N_22966,N_13314,N_17045);
and U22967 (N_22967,N_12215,N_14518);
and U22968 (N_22968,N_15367,N_12984);
xnor U22969 (N_22969,N_12592,N_12133);
and U22970 (N_22970,N_12636,N_14510);
xnor U22971 (N_22971,N_15938,N_15975);
or U22972 (N_22972,N_16333,N_16632);
nor U22973 (N_22973,N_15046,N_12273);
nor U22974 (N_22974,N_12161,N_17603);
nor U22975 (N_22975,N_17644,N_14541);
nand U22976 (N_22976,N_16583,N_16486);
or U22977 (N_22977,N_17778,N_15504);
or U22978 (N_22978,N_17032,N_12936);
nor U22979 (N_22979,N_17532,N_13138);
or U22980 (N_22980,N_16589,N_14851);
xor U22981 (N_22981,N_14566,N_17200);
and U22982 (N_22982,N_13860,N_12555);
and U22983 (N_22983,N_16529,N_14840);
nor U22984 (N_22984,N_15996,N_16876);
xor U22985 (N_22985,N_17202,N_16356);
and U22986 (N_22986,N_14903,N_16019);
xnor U22987 (N_22987,N_17945,N_17224);
and U22988 (N_22988,N_14515,N_13102);
or U22989 (N_22989,N_12493,N_15755);
and U22990 (N_22990,N_14203,N_15167);
and U22991 (N_22991,N_14960,N_12386);
nand U22992 (N_22992,N_14416,N_12511);
or U22993 (N_22993,N_16910,N_16943);
nor U22994 (N_22994,N_17396,N_17359);
nand U22995 (N_22995,N_15708,N_16881);
or U22996 (N_22996,N_14450,N_16296);
nand U22997 (N_22997,N_15457,N_17115);
xnor U22998 (N_22998,N_15086,N_13069);
and U22999 (N_22999,N_15588,N_16369);
and U23000 (N_23000,N_17470,N_14524);
xor U23001 (N_23001,N_13763,N_14913);
and U23002 (N_23002,N_12260,N_14121);
nand U23003 (N_23003,N_12957,N_17292);
or U23004 (N_23004,N_15875,N_12380);
and U23005 (N_23005,N_16714,N_16663);
and U23006 (N_23006,N_14005,N_12770);
xnor U23007 (N_23007,N_14428,N_16007);
nor U23008 (N_23008,N_17950,N_13467);
nor U23009 (N_23009,N_12600,N_12965);
xnor U23010 (N_23010,N_14586,N_15225);
or U23011 (N_23011,N_12432,N_14501);
and U23012 (N_23012,N_15204,N_14662);
nor U23013 (N_23013,N_12387,N_17486);
and U23014 (N_23014,N_13429,N_15577);
xor U23015 (N_23015,N_12646,N_13136);
and U23016 (N_23016,N_12017,N_17407);
xor U23017 (N_23017,N_12047,N_15676);
nand U23018 (N_23018,N_12285,N_12378);
nand U23019 (N_23019,N_12139,N_14494);
xnor U23020 (N_23020,N_15641,N_17132);
and U23021 (N_23021,N_16314,N_15468);
nand U23022 (N_23022,N_15357,N_14467);
nand U23023 (N_23023,N_15027,N_17784);
and U23024 (N_23024,N_15196,N_16236);
or U23025 (N_23025,N_15242,N_14703);
and U23026 (N_23026,N_14429,N_12642);
nor U23027 (N_23027,N_13127,N_16622);
and U23028 (N_23028,N_15218,N_17430);
and U23029 (N_23029,N_13958,N_13935);
and U23030 (N_23030,N_12180,N_13950);
and U23031 (N_23031,N_17202,N_16199);
xor U23032 (N_23032,N_14253,N_13269);
and U23033 (N_23033,N_15471,N_15231);
nand U23034 (N_23034,N_15547,N_13660);
xnor U23035 (N_23035,N_15809,N_14279);
xnor U23036 (N_23036,N_13963,N_14096);
nor U23037 (N_23037,N_15167,N_16020);
xor U23038 (N_23038,N_13113,N_15259);
nor U23039 (N_23039,N_17599,N_13701);
or U23040 (N_23040,N_15486,N_12885);
nor U23041 (N_23041,N_13968,N_16724);
or U23042 (N_23042,N_14727,N_17649);
or U23043 (N_23043,N_12521,N_14697);
or U23044 (N_23044,N_17799,N_16615);
or U23045 (N_23045,N_17204,N_15386);
xor U23046 (N_23046,N_16814,N_14471);
or U23047 (N_23047,N_15624,N_12664);
xnor U23048 (N_23048,N_15904,N_13425);
nand U23049 (N_23049,N_17878,N_16920);
nand U23050 (N_23050,N_17661,N_17531);
or U23051 (N_23051,N_13007,N_13583);
and U23052 (N_23052,N_17651,N_12607);
xor U23053 (N_23053,N_12226,N_16479);
and U23054 (N_23054,N_12151,N_16406);
nand U23055 (N_23055,N_12478,N_17035);
nand U23056 (N_23056,N_12529,N_15648);
nor U23057 (N_23057,N_12191,N_16515);
nor U23058 (N_23058,N_13760,N_16645);
xor U23059 (N_23059,N_17591,N_17398);
nor U23060 (N_23060,N_13512,N_16536);
xor U23061 (N_23061,N_12257,N_13254);
nand U23062 (N_23062,N_14144,N_12592);
nand U23063 (N_23063,N_13289,N_14223);
and U23064 (N_23064,N_15620,N_17904);
nand U23065 (N_23065,N_12635,N_13948);
and U23066 (N_23066,N_17056,N_12251);
nand U23067 (N_23067,N_16078,N_14841);
xnor U23068 (N_23068,N_16270,N_16828);
or U23069 (N_23069,N_16498,N_16785);
and U23070 (N_23070,N_17730,N_14473);
and U23071 (N_23071,N_12836,N_15494);
xnor U23072 (N_23072,N_16434,N_16089);
xor U23073 (N_23073,N_12038,N_17133);
nand U23074 (N_23074,N_16216,N_14391);
or U23075 (N_23075,N_12999,N_14698);
or U23076 (N_23076,N_14585,N_17871);
or U23077 (N_23077,N_14886,N_16921);
or U23078 (N_23078,N_13358,N_14180);
xor U23079 (N_23079,N_17194,N_13271);
or U23080 (N_23080,N_17905,N_12509);
nor U23081 (N_23081,N_14610,N_14627);
nor U23082 (N_23082,N_13793,N_15470);
and U23083 (N_23083,N_16769,N_15474);
xnor U23084 (N_23084,N_15139,N_15928);
or U23085 (N_23085,N_13593,N_12657);
nand U23086 (N_23086,N_14595,N_16521);
nand U23087 (N_23087,N_12271,N_17376);
and U23088 (N_23088,N_15352,N_14365);
and U23089 (N_23089,N_13945,N_13153);
or U23090 (N_23090,N_13707,N_16171);
or U23091 (N_23091,N_14587,N_14517);
or U23092 (N_23092,N_12705,N_16240);
or U23093 (N_23093,N_16409,N_17184);
nand U23094 (N_23094,N_16992,N_14012);
xnor U23095 (N_23095,N_13917,N_13796);
xnor U23096 (N_23096,N_12419,N_13609);
nand U23097 (N_23097,N_15743,N_12933);
and U23098 (N_23098,N_16925,N_17406);
nand U23099 (N_23099,N_15695,N_13113);
nor U23100 (N_23100,N_13270,N_15039);
nor U23101 (N_23101,N_12040,N_17168);
and U23102 (N_23102,N_14128,N_13435);
or U23103 (N_23103,N_15575,N_12330);
and U23104 (N_23104,N_16676,N_12073);
nor U23105 (N_23105,N_15086,N_15917);
xor U23106 (N_23106,N_15852,N_13681);
nor U23107 (N_23107,N_13181,N_13306);
nor U23108 (N_23108,N_16331,N_12022);
and U23109 (N_23109,N_16454,N_14660);
or U23110 (N_23110,N_16749,N_12171);
or U23111 (N_23111,N_16835,N_14559);
or U23112 (N_23112,N_16180,N_16535);
nor U23113 (N_23113,N_15036,N_17487);
xor U23114 (N_23114,N_12272,N_12933);
xnor U23115 (N_23115,N_16705,N_13998);
nor U23116 (N_23116,N_13616,N_12179);
or U23117 (N_23117,N_17466,N_17602);
and U23118 (N_23118,N_17419,N_14050);
nor U23119 (N_23119,N_13867,N_14342);
nor U23120 (N_23120,N_16494,N_12071);
nor U23121 (N_23121,N_13685,N_17652);
xor U23122 (N_23122,N_13727,N_16337);
nand U23123 (N_23123,N_13146,N_17370);
nor U23124 (N_23124,N_12053,N_13826);
or U23125 (N_23125,N_13405,N_12663);
and U23126 (N_23126,N_16049,N_13653);
nand U23127 (N_23127,N_17556,N_14949);
and U23128 (N_23128,N_15582,N_15244);
nand U23129 (N_23129,N_14101,N_17388);
or U23130 (N_23130,N_16840,N_17729);
xor U23131 (N_23131,N_14422,N_12970);
and U23132 (N_23132,N_15752,N_13623);
xnor U23133 (N_23133,N_15105,N_13595);
nor U23134 (N_23134,N_14824,N_13363);
and U23135 (N_23135,N_15973,N_15142);
nor U23136 (N_23136,N_15638,N_15283);
nor U23137 (N_23137,N_16602,N_15118);
nor U23138 (N_23138,N_14006,N_17652);
nand U23139 (N_23139,N_16750,N_13524);
nor U23140 (N_23140,N_15243,N_14165);
or U23141 (N_23141,N_17903,N_17279);
and U23142 (N_23142,N_12643,N_13284);
nand U23143 (N_23143,N_13745,N_15844);
and U23144 (N_23144,N_14645,N_15728);
nand U23145 (N_23145,N_14020,N_12280);
nand U23146 (N_23146,N_16106,N_17615);
and U23147 (N_23147,N_13474,N_12134);
or U23148 (N_23148,N_14169,N_15017);
or U23149 (N_23149,N_15317,N_12082);
nor U23150 (N_23150,N_17751,N_14554);
xor U23151 (N_23151,N_14465,N_14848);
or U23152 (N_23152,N_17155,N_13004);
nor U23153 (N_23153,N_12946,N_13035);
nand U23154 (N_23154,N_16455,N_14205);
nor U23155 (N_23155,N_15129,N_13594);
nor U23156 (N_23156,N_13666,N_17973);
and U23157 (N_23157,N_16556,N_16742);
and U23158 (N_23158,N_17031,N_17241);
nor U23159 (N_23159,N_16392,N_13386);
and U23160 (N_23160,N_12104,N_15421);
or U23161 (N_23161,N_15951,N_14122);
nor U23162 (N_23162,N_14408,N_14538);
and U23163 (N_23163,N_17415,N_17203);
or U23164 (N_23164,N_13212,N_12788);
nor U23165 (N_23165,N_15737,N_14448);
nor U23166 (N_23166,N_14092,N_12237);
xnor U23167 (N_23167,N_15563,N_17716);
nand U23168 (N_23168,N_16237,N_13036);
or U23169 (N_23169,N_16811,N_15789);
xnor U23170 (N_23170,N_12911,N_12793);
nand U23171 (N_23171,N_13151,N_13888);
or U23172 (N_23172,N_15754,N_17026);
nand U23173 (N_23173,N_13858,N_12859);
xnor U23174 (N_23174,N_14709,N_13253);
nand U23175 (N_23175,N_12869,N_17942);
xor U23176 (N_23176,N_16463,N_15718);
nor U23177 (N_23177,N_13557,N_13318);
nand U23178 (N_23178,N_16678,N_16905);
and U23179 (N_23179,N_12328,N_16359);
nand U23180 (N_23180,N_14527,N_15209);
nor U23181 (N_23181,N_15542,N_17276);
xnor U23182 (N_23182,N_16536,N_12772);
xor U23183 (N_23183,N_13502,N_16746);
or U23184 (N_23184,N_14622,N_14625);
nand U23185 (N_23185,N_15840,N_15234);
nor U23186 (N_23186,N_17970,N_12649);
and U23187 (N_23187,N_15475,N_13867);
and U23188 (N_23188,N_12700,N_13871);
or U23189 (N_23189,N_16886,N_17653);
nand U23190 (N_23190,N_16776,N_16191);
xnor U23191 (N_23191,N_15963,N_16461);
nand U23192 (N_23192,N_12936,N_13580);
nor U23193 (N_23193,N_17619,N_14740);
and U23194 (N_23194,N_15324,N_14032);
or U23195 (N_23195,N_15501,N_13795);
and U23196 (N_23196,N_16429,N_12339);
nand U23197 (N_23197,N_14570,N_16800);
and U23198 (N_23198,N_14448,N_15120);
nor U23199 (N_23199,N_14217,N_12933);
nor U23200 (N_23200,N_16208,N_12283);
or U23201 (N_23201,N_13748,N_16961);
and U23202 (N_23202,N_14330,N_14010);
or U23203 (N_23203,N_13760,N_15726);
or U23204 (N_23204,N_16026,N_12836);
nor U23205 (N_23205,N_17971,N_12283);
xor U23206 (N_23206,N_13432,N_15725);
or U23207 (N_23207,N_16925,N_12280);
nand U23208 (N_23208,N_17008,N_12619);
xor U23209 (N_23209,N_16639,N_12560);
and U23210 (N_23210,N_15883,N_13921);
nor U23211 (N_23211,N_17193,N_14612);
or U23212 (N_23212,N_16065,N_12041);
and U23213 (N_23213,N_17267,N_14307);
and U23214 (N_23214,N_17458,N_14094);
nor U23215 (N_23215,N_13561,N_16488);
nand U23216 (N_23216,N_13927,N_12603);
and U23217 (N_23217,N_15359,N_13584);
nand U23218 (N_23218,N_14527,N_17865);
and U23219 (N_23219,N_15092,N_17753);
xnor U23220 (N_23220,N_13042,N_12276);
or U23221 (N_23221,N_15582,N_15070);
or U23222 (N_23222,N_15397,N_14771);
nand U23223 (N_23223,N_17283,N_12690);
nand U23224 (N_23224,N_12462,N_14724);
and U23225 (N_23225,N_13309,N_13578);
xor U23226 (N_23226,N_16854,N_12675);
and U23227 (N_23227,N_15855,N_15752);
and U23228 (N_23228,N_16478,N_15160);
nand U23229 (N_23229,N_15405,N_13090);
and U23230 (N_23230,N_14436,N_12375);
and U23231 (N_23231,N_16325,N_14119);
and U23232 (N_23232,N_15985,N_12658);
xnor U23233 (N_23233,N_14659,N_12555);
and U23234 (N_23234,N_13631,N_14343);
or U23235 (N_23235,N_15579,N_14815);
or U23236 (N_23236,N_12040,N_14415);
and U23237 (N_23237,N_16787,N_15093);
nor U23238 (N_23238,N_12910,N_13704);
or U23239 (N_23239,N_16179,N_13619);
nor U23240 (N_23240,N_14173,N_12476);
or U23241 (N_23241,N_14699,N_13944);
and U23242 (N_23242,N_15922,N_15619);
or U23243 (N_23243,N_14670,N_14525);
and U23244 (N_23244,N_14651,N_17059);
and U23245 (N_23245,N_15091,N_17343);
or U23246 (N_23246,N_15577,N_16636);
xor U23247 (N_23247,N_13480,N_15767);
and U23248 (N_23248,N_17784,N_15404);
nand U23249 (N_23249,N_12868,N_15436);
xnor U23250 (N_23250,N_14695,N_13760);
or U23251 (N_23251,N_17744,N_14322);
xnor U23252 (N_23252,N_15230,N_17085);
xnor U23253 (N_23253,N_15370,N_16986);
and U23254 (N_23254,N_15037,N_13417);
or U23255 (N_23255,N_17732,N_15598);
and U23256 (N_23256,N_12057,N_15636);
nor U23257 (N_23257,N_13295,N_15692);
xnor U23258 (N_23258,N_12869,N_13125);
nand U23259 (N_23259,N_17729,N_14518);
or U23260 (N_23260,N_13256,N_13790);
or U23261 (N_23261,N_12194,N_13753);
or U23262 (N_23262,N_15559,N_17806);
and U23263 (N_23263,N_16768,N_12952);
xor U23264 (N_23264,N_16519,N_15602);
nor U23265 (N_23265,N_13874,N_14769);
or U23266 (N_23266,N_16926,N_17305);
xnor U23267 (N_23267,N_17967,N_17939);
xnor U23268 (N_23268,N_12118,N_16330);
or U23269 (N_23269,N_14016,N_15082);
nand U23270 (N_23270,N_15754,N_16304);
or U23271 (N_23271,N_12800,N_17693);
nor U23272 (N_23272,N_13309,N_12282);
or U23273 (N_23273,N_15940,N_16922);
and U23274 (N_23274,N_15268,N_13322);
nor U23275 (N_23275,N_12447,N_14401);
xnor U23276 (N_23276,N_16846,N_13573);
nor U23277 (N_23277,N_12606,N_13390);
nand U23278 (N_23278,N_16661,N_14646);
xnor U23279 (N_23279,N_12452,N_12162);
and U23280 (N_23280,N_14902,N_14641);
nor U23281 (N_23281,N_15100,N_13373);
and U23282 (N_23282,N_12512,N_13452);
nand U23283 (N_23283,N_14064,N_12020);
nor U23284 (N_23284,N_16082,N_17832);
or U23285 (N_23285,N_13507,N_16874);
or U23286 (N_23286,N_17309,N_14414);
nor U23287 (N_23287,N_17044,N_14623);
nor U23288 (N_23288,N_14588,N_14327);
xnor U23289 (N_23289,N_17822,N_17903);
nor U23290 (N_23290,N_15740,N_17129);
and U23291 (N_23291,N_15948,N_17121);
nor U23292 (N_23292,N_17148,N_16560);
and U23293 (N_23293,N_17233,N_13733);
xor U23294 (N_23294,N_14375,N_14855);
nand U23295 (N_23295,N_12072,N_16848);
nand U23296 (N_23296,N_14502,N_13382);
nor U23297 (N_23297,N_14588,N_15351);
xnor U23298 (N_23298,N_14868,N_12954);
nand U23299 (N_23299,N_12881,N_12636);
nor U23300 (N_23300,N_16660,N_15050);
xor U23301 (N_23301,N_13624,N_14653);
nor U23302 (N_23302,N_12144,N_16573);
or U23303 (N_23303,N_15256,N_14500);
and U23304 (N_23304,N_16424,N_13922);
or U23305 (N_23305,N_13931,N_15756);
nor U23306 (N_23306,N_12061,N_14865);
and U23307 (N_23307,N_13487,N_12314);
nor U23308 (N_23308,N_12144,N_15537);
xnor U23309 (N_23309,N_12605,N_12091);
xnor U23310 (N_23310,N_16965,N_17566);
nand U23311 (N_23311,N_17729,N_12117);
nand U23312 (N_23312,N_14086,N_15868);
xor U23313 (N_23313,N_14377,N_12202);
or U23314 (N_23314,N_15902,N_15461);
and U23315 (N_23315,N_14664,N_15230);
xnor U23316 (N_23316,N_13734,N_13074);
or U23317 (N_23317,N_17914,N_15712);
xnor U23318 (N_23318,N_16540,N_17670);
nor U23319 (N_23319,N_12005,N_13708);
and U23320 (N_23320,N_15666,N_13350);
or U23321 (N_23321,N_17235,N_13370);
or U23322 (N_23322,N_13129,N_13155);
or U23323 (N_23323,N_14419,N_12790);
nor U23324 (N_23324,N_16007,N_13620);
nor U23325 (N_23325,N_17363,N_12529);
xor U23326 (N_23326,N_17670,N_16631);
or U23327 (N_23327,N_15924,N_16360);
nand U23328 (N_23328,N_15280,N_15184);
xor U23329 (N_23329,N_17138,N_17337);
nand U23330 (N_23330,N_14450,N_12637);
and U23331 (N_23331,N_14406,N_16107);
and U23332 (N_23332,N_16770,N_12950);
and U23333 (N_23333,N_17266,N_15842);
xor U23334 (N_23334,N_16396,N_17170);
nor U23335 (N_23335,N_15856,N_13076);
nand U23336 (N_23336,N_16224,N_15671);
or U23337 (N_23337,N_12007,N_12332);
and U23338 (N_23338,N_12310,N_13344);
nor U23339 (N_23339,N_15978,N_15689);
nor U23340 (N_23340,N_17589,N_14170);
or U23341 (N_23341,N_14840,N_13462);
xnor U23342 (N_23342,N_16333,N_15173);
nor U23343 (N_23343,N_17940,N_17353);
or U23344 (N_23344,N_15208,N_13578);
xor U23345 (N_23345,N_17763,N_15505);
nor U23346 (N_23346,N_17289,N_17308);
and U23347 (N_23347,N_14905,N_12108);
nor U23348 (N_23348,N_14511,N_14010);
and U23349 (N_23349,N_12121,N_13766);
xor U23350 (N_23350,N_16415,N_16867);
xnor U23351 (N_23351,N_16339,N_15107);
nor U23352 (N_23352,N_13622,N_12509);
nand U23353 (N_23353,N_17921,N_12650);
xnor U23354 (N_23354,N_14478,N_12251);
or U23355 (N_23355,N_14879,N_13730);
nand U23356 (N_23356,N_12377,N_16918);
and U23357 (N_23357,N_16386,N_16816);
nor U23358 (N_23358,N_15401,N_17966);
xor U23359 (N_23359,N_12944,N_14048);
and U23360 (N_23360,N_13899,N_17814);
nor U23361 (N_23361,N_17196,N_17065);
nand U23362 (N_23362,N_14180,N_14708);
and U23363 (N_23363,N_16127,N_12340);
and U23364 (N_23364,N_15384,N_16389);
or U23365 (N_23365,N_13118,N_12876);
and U23366 (N_23366,N_14990,N_17474);
nand U23367 (N_23367,N_16158,N_15739);
or U23368 (N_23368,N_17108,N_14145);
and U23369 (N_23369,N_17927,N_12337);
xor U23370 (N_23370,N_17422,N_12678);
or U23371 (N_23371,N_13417,N_15146);
nor U23372 (N_23372,N_16012,N_14907);
or U23373 (N_23373,N_13854,N_12690);
nand U23374 (N_23374,N_12968,N_16482);
or U23375 (N_23375,N_16937,N_14064);
or U23376 (N_23376,N_15949,N_13071);
xor U23377 (N_23377,N_15778,N_12331);
xor U23378 (N_23378,N_15353,N_12831);
nand U23379 (N_23379,N_16760,N_16381);
nor U23380 (N_23380,N_12946,N_17446);
nand U23381 (N_23381,N_16224,N_17743);
nand U23382 (N_23382,N_15959,N_17770);
or U23383 (N_23383,N_16492,N_13755);
nor U23384 (N_23384,N_16049,N_16765);
nor U23385 (N_23385,N_13225,N_12622);
nor U23386 (N_23386,N_15940,N_12732);
nor U23387 (N_23387,N_16249,N_14709);
nand U23388 (N_23388,N_12516,N_13490);
and U23389 (N_23389,N_16784,N_13690);
and U23390 (N_23390,N_13580,N_12719);
xor U23391 (N_23391,N_17904,N_14266);
nand U23392 (N_23392,N_14897,N_15030);
xor U23393 (N_23393,N_13451,N_14276);
or U23394 (N_23394,N_12546,N_17699);
or U23395 (N_23395,N_14890,N_17107);
xor U23396 (N_23396,N_15364,N_16260);
or U23397 (N_23397,N_15174,N_12722);
nand U23398 (N_23398,N_14772,N_12415);
xor U23399 (N_23399,N_15931,N_12455);
nor U23400 (N_23400,N_16238,N_15511);
xor U23401 (N_23401,N_15900,N_15080);
or U23402 (N_23402,N_12739,N_14123);
and U23403 (N_23403,N_15165,N_16600);
and U23404 (N_23404,N_15077,N_13087);
and U23405 (N_23405,N_12816,N_13952);
xor U23406 (N_23406,N_14560,N_17629);
nand U23407 (N_23407,N_14027,N_14383);
and U23408 (N_23408,N_13240,N_15128);
xnor U23409 (N_23409,N_12690,N_15473);
and U23410 (N_23410,N_17579,N_14675);
and U23411 (N_23411,N_12403,N_17408);
or U23412 (N_23412,N_15422,N_16322);
nand U23413 (N_23413,N_13047,N_14430);
nand U23414 (N_23414,N_16958,N_15847);
and U23415 (N_23415,N_13188,N_14577);
and U23416 (N_23416,N_13993,N_15084);
nand U23417 (N_23417,N_17514,N_12338);
nor U23418 (N_23418,N_15162,N_17437);
and U23419 (N_23419,N_17458,N_14652);
nand U23420 (N_23420,N_15962,N_15922);
and U23421 (N_23421,N_13012,N_12268);
nor U23422 (N_23422,N_16266,N_13836);
xnor U23423 (N_23423,N_17971,N_17565);
or U23424 (N_23424,N_13861,N_16554);
or U23425 (N_23425,N_13996,N_12392);
or U23426 (N_23426,N_14948,N_13773);
or U23427 (N_23427,N_15703,N_13949);
nand U23428 (N_23428,N_16277,N_13613);
xnor U23429 (N_23429,N_15706,N_14310);
xor U23430 (N_23430,N_17152,N_16033);
nand U23431 (N_23431,N_15012,N_16007);
or U23432 (N_23432,N_12073,N_14570);
xor U23433 (N_23433,N_13762,N_12016);
nand U23434 (N_23434,N_16162,N_17734);
xor U23435 (N_23435,N_12660,N_14802);
and U23436 (N_23436,N_16273,N_13902);
or U23437 (N_23437,N_13906,N_16076);
xor U23438 (N_23438,N_13204,N_17826);
nand U23439 (N_23439,N_14847,N_17394);
or U23440 (N_23440,N_14854,N_13001);
nor U23441 (N_23441,N_14048,N_12218);
xnor U23442 (N_23442,N_14132,N_16550);
or U23443 (N_23443,N_15693,N_17432);
nor U23444 (N_23444,N_12011,N_13387);
nor U23445 (N_23445,N_15762,N_17751);
xnor U23446 (N_23446,N_12646,N_13673);
xor U23447 (N_23447,N_16833,N_12841);
or U23448 (N_23448,N_12776,N_17237);
and U23449 (N_23449,N_12134,N_13730);
nand U23450 (N_23450,N_17832,N_14418);
and U23451 (N_23451,N_13199,N_16646);
nand U23452 (N_23452,N_15401,N_13027);
nand U23453 (N_23453,N_15504,N_16616);
nor U23454 (N_23454,N_16693,N_13879);
nor U23455 (N_23455,N_12143,N_17890);
and U23456 (N_23456,N_14094,N_15068);
nand U23457 (N_23457,N_16756,N_12407);
nor U23458 (N_23458,N_15971,N_15399);
or U23459 (N_23459,N_13371,N_12460);
xnor U23460 (N_23460,N_13544,N_16798);
nor U23461 (N_23461,N_17310,N_16463);
or U23462 (N_23462,N_16069,N_17267);
nor U23463 (N_23463,N_12724,N_14765);
and U23464 (N_23464,N_13400,N_17849);
or U23465 (N_23465,N_13489,N_16794);
and U23466 (N_23466,N_14360,N_17808);
nor U23467 (N_23467,N_13020,N_16706);
nand U23468 (N_23468,N_13381,N_17527);
nor U23469 (N_23469,N_16841,N_17003);
or U23470 (N_23470,N_14885,N_16911);
or U23471 (N_23471,N_17397,N_13286);
and U23472 (N_23472,N_12673,N_14348);
nand U23473 (N_23473,N_14326,N_15782);
nor U23474 (N_23474,N_14549,N_13462);
nor U23475 (N_23475,N_16483,N_14701);
xor U23476 (N_23476,N_14319,N_14953);
xor U23477 (N_23477,N_15362,N_15603);
nor U23478 (N_23478,N_13256,N_15956);
nor U23479 (N_23479,N_12058,N_13403);
nor U23480 (N_23480,N_15613,N_14171);
nor U23481 (N_23481,N_13801,N_15060);
nor U23482 (N_23482,N_17615,N_17229);
nand U23483 (N_23483,N_14995,N_16777);
xor U23484 (N_23484,N_14972,N_13933);
nor U23485 (N_23485,N_15466,N_17811);
or U23486 (N_23486,N_13428,N_17167);
or U23487 (N_23487,N_14869,N_12959);
and U23488 (N_23488,N_16708,N_15218);
xnor U23489 (N_23489,N_15258,N_17853);
or U23490 (N_23490,N_15216,N_12804);
or U23491 (N_23491,N_17492,N_13938);
or U23492 (N_23492,N_16738,N_12020);
nand U23493 (N_23493,N_12526,N_17774);
nor U23494 (N_23494,N_12023,N_12131);
and U23495 (N_23495,N_17052,N_12569);
or U23496 (N_23496,N_13501,N_17201);
nor U23497 (N_23497,N_13375,N_15127);
or U23498 (N_23498,N_17783,N_15271);
and U23499 (N_23499,N_12304,N_12567);
xor U23500 (N_23500,N_17893,N_16318);
nand U23501 (N_23501,N_12650,N_12768);
xor U23502 (N_23502,N_15898,N_13109);
nor U23503 (N_23503,N_12039,N_12817);
and U23504 (N_23504,N_16756,N_14908);
or U23505 (N_23505,N_15227,N_17231);
and U23506 (N_23506,N_12565,N_14489);
or U23507 (N_23507,N_13745,N_12794);
or U23508 (N_23508,N_14999,N_12592);
xor U23509 (N_23509,N_16770,N_14155);
nand U23510 (N_23510,N_13637,N_12040);
nor U23511 (N_23511,N_13999,N_15775);
nor U23512 (N_23512,N_14215,N_17965);
and U23513 (N_23513,N_13754,N_16626);
nand U23514 (N_23514,N_17809,N_12244);
and U23515 (N_23515,N_17105,N_13766);
or U23516 (N_23516,N_15609,N_17898);
nor U23517 (N_23517,N_16556,N_13649);
nor U23518 (N_23518,N_13261,N_13247);
and U23519 (N_23519,N_13359,N_17056);
xor U23520 (N_23520,N_12932,N_15890);
and U23521 (N_23521,N_13633,N_17857);
nor U23522 (N_23522,N_16852,N_12511);
and U23523 (N_23523,N_17707,N_13287);
and U23524 (N_23524,N_13878,N_13187);
nand U23525 (N_23525,N_15361,N_12795);
xnor U23526 (N_23526,N_16218,N_13900);
and U23527 (N_23527,N_15257,N_13448);
xor U23528 (N_23528,N_15548,N_12025);
and U23529 (N_23529,N_12827,N_12987);
nand U23530 (N_23530,N_13495,N_12410);
nor U23531 (N_23531,N_17357,N_13357);
xor U23532 (N_23532,N_12272,N_16690);
or U23533 (N_23533,N_16695,N_14191);
or U23534 (N_23534,N_12088,N_13973);
or U23535 (N_23535,N_16400,N_14801);
xor U23536 (N_23536,N_13796,N_12504);
nor U23537 (N_23537,N_16202,N_13495);
nor U23538 (N_23538,N_17380,N_14994);
xnor U23539 (N_23539,N_12237,N_17019);
nand U23540 (N_23540,N_15409,N_15774);
xnor U23541 (N_23541,N_17052,N_13652);
or U23542 (N_23542,N_12084,N_16989);
nand U23543 (N_23543,N_14395,N_13031);
xnor U23544 (N_23544,N_12451,N_17041);
or U23545 (N_23545,N_15696,N_12989);
nor U23546 (N_23546,N_15797,N_15390);
xnor U23547 (N_23547,N_17442,N_13045);
nand U23548 (N_23548,N_16744,N_17200);
xor U23549 (N_23549,N_14629,N_16182);
or U23550 (N_23550,N_13034,N_16673);
nand U23551 (N_23551,N_14023,N_13571);
or U23552 (N_23552,N_17524,N_12559);
nor U23553 (N_23553,N_17817,N_16653);
or U23554 (N_23554,N_15631,N_14511);
nand U23555 (N_23555,N_15449,N_16447);
and U23556 (N_23556,N_17222,N_13520);
xnor U23557 (N_23557,N_12046,N_14725);
or U23558 (N_23558,N_16896,N_12798);
or U23559 (N_23559,N_12429,N_14485);
or U23560 (N_23560,N_17814,N_15927);
xnor U23561 (N_23561,N_17728,N_14677);
and U23562 (N_23562,N_16913,N_12818);
xor U23563 (N_23563,N_14700,N_14453);
nor U23564 (N_23564,N_14091,N_15586);
and U23565 (N_23565,N_16168,N_14402);
or U23566 (N_23566,N_17366,N_15232);
nor U23567 (N_23567,N_14038,N_16622);
nand U23568 (N_23568,N_12092,N_12326);
xnor U23569 (N_23569,N_13230,N_14511);
or U23570 (N_23570,N_17275,N_13369);
xor U23571 (N_23571,N_13589,N_16392);
or U23572 (N_23572,N_12827,N_17287);
and U23573 (N_23573,N_14663,N_16158);
nor U23574 (N_23574,N_16829,N_16873);
xnor U23575 (N_23575,N_17897,N_16657);
nor U23576 (N_23576,N_13687,N_13866);
nor U23577 (N_23577,N_15660,N_14225);
nand U23578 (N_23578,N_13873,N_13770);
and U23579 (N_23579,N_16529,N_14636);
or U23580 (N_23580,N_13606,N_13533);
xor U23581 (N_23581,N_12996,N_15466);
nand U23582 (N_23582,N_14933,N_15878);
nor U23583 (N_23583,N_14860,N_15437);
nand U23584 (N_23584,N_14064,N_14083);
xnor U23585 (N_23585,N_12521,N_17056);
nand U23586 (N_23586,N_14340,N_15213);
or U23587 (N_23587,N_14144,N_14605);
nor U23588 (N_23588,N_12523,N_16035);
xnor U23589 (N_23589,N_13107,N_13885);
nor U23590 (N_23590,N_17745,N_13496);
nand U23591 (N_23591,N_13097,N_13092);
nor U23592 (N_23592,N_12447,N_17886);
and U23593 (N_23593,N_14451,N_12675);
xnor U23594 (N_23594,N_16098,N_15835);
and U23595 (N_23595,N_13753,N_12817);
or U23596 (N_23596,N_17962,N_15631);
and U23597 (N_23597,N_12516,N_17777);
nor U23598 (N_23598,N_16014,N_12199);
or U23599 (N_23599,N_15280,N_12721);
nor U23600 (N_23600,N_13427,N_12829);
nand U23601 (N_23601,N_17478,N_17003);
nor U23602 (N_23602,N_12336,N_14748);
nand U23603 (N_23603,N_17026,N_15579);
or U23604 (N_23604,N_12843,N_13118);
and U23605 (N_23605,N_17112,N_12815);
or U23606 (N_23606,N_12155,N_13470);
nand U23607 (N_23607,N_15940,N_13037);
nor U23608 (N_23608,N_13094,N_15908);
nand U23609 (N_23609,N_12337,N_17897);
nor U23610 (N_23610,N_15821,N_14111);
and U23611 (N_23611,N_15891,N_16841);
nand U23612 (N_23612,N_13626,N_15077);
or U23613 (N_23613,N_16092,N_17621);
xor U23614 (N_23614,N_16540,N_17214);
nor U23615 (N_23615,N_16782,N_13059);
nand U23616 (N_23616,N_15570,N_17785);
and U23617 (N_23617,N_17240,N_15086);
nand U23618 (N_23618,N_13793,N_14269);
xor U23619 (N_23619,N_16493,N_12510);
nand U23620 (N_23620,N_12710,N_15141);
or U23621 (N_23621,N_14312,N_17332);
xnor U23622 (N_23622,N_12342,N_12053);
nor U23623 (N_23623,N_17179,N_15021);
nand U23624 (N_23624,N_12661,N_14852);
nor U23625 (N_23625,N_16813,N_12546);
and U23626 (N_23626,N_13120,N_13675);
nor U23627 (N_23627,N_16529,N_12887);
nand U23628 (N_23628,N_15769,N_17706);
and U23629 (N_23629,N_15575,N_17544);
or U23630 (N_23630,N_17075,N_15939);
nor U23631 (N_23631,N_15525,N_17929);
nor U23632 (N_23632,N_15531,N_12627);
xnor U23633 (N_23633,N_17577,N_14670);
and U23634 (N_23634,N_12040,N_13833);
xor U23635 (N_23635,N_16080,N_14022);
xor U23636 (N_23636,N_14787,N_17345);
and U23637 (N_23637,N_13128,N_14514);
and U23638 (N_23638,N_14876,N_16387);
nand U23639 (N_23639,N_17884,N_16495);
or U23640 (N_23640,N_12275,N_17905);
and U23641 (N_23641,N_17109,N_16552);
or U23642 (N_23642,N_14018,N_15332);
xor U23643 (N_23643,N_15658,N_12401);
nor U23644 (N_23644,N_16928,N_12195);
nand U23645 (N_23645,N_13520,N_12502);
nor U23646 (N_23646,N_17254,N_16654);
xor U23647 (N_23647,N_15899,N_12509);
or U23648 (N_23648,N_13691,N_16533);
or U23649 (N_23649,N_15932,N_12979);
nor U23650 (N_23650,N_15061,N_15317);
or U23651 (N_23651,N_16194,N_12468);
and U23652 (N_23652,N_14729,N_14567);
xnor U23653 (N_23653,N_13479,N_14621);
nand U23654 (N_23654,N_15814,N_12946);
nor U23655 (N_23655,N_16927,N_17764);
or U23656 (N_23656,N_12458,N_16612);
nand U23657 (N_23657,N_13061,N_17578);
nor U23658 (N_23658,N_13485,N_14357);
xnor U23659 (N_23659,N_16449,N_14696);
nand U23660 (N_23660,N_12504,N_14772);
and U23661 (N_23661,N_17468,N_17330);
and U23662 (N_23662,N_14741,N_15044);
or U23663 (N_23663,N_14013,N_15014);
or U23664 (N_23664,N_17110,N_14435);
nor U23665 (N_23665,N_14350,N_16224);
nand U23666 (N_23666,N_12482,N_16194);
and U23667 (N_23667,N_12275,N_14725);
or U23668 (N_23668,N_16288,N_17125);
and U23669 (N_23669,N_13811,N_13775);
nor U23670 (N_23670,N_12830,N_16719);
xor U23671 (N_23671,N_16916,N_12965);
or U23672 (N_23672,N_13157,N_14430);
or U23673 (N_23673,N_16778,N_15896);
nor U23674 (N_23674,N_16585,N_14755);
or U23675 (N_23675,N_17555,N_12792);
and U23676 (N_23676,N_16970,N_15920);
and U23677 (N_23677,N_16902,N_17837);
and U23678 (N_23678,N_12868,N_12776);
nor U23679 (N_23679,N_17780,N_15279);
xnor U23680 (N_23680,N_14653,N_15844);
xnor U23681 (N_23681,N_14845,N_15022);
xnor U23682 (N_23682,N_17738,N_13383);
xnor U23683 (N_23683,N_14163,N_12189);
and U23684 (N_23684,N_17459,N_17938);
xnor U23685 (N_23685,N_16465,N_14637);
nor U23686 (N_23686,N_16080,N_15378);
and U23687 (N_23687,N_14681,N_16035);
xnor U23688 (N_23688,N_13400,N_12257);
xnor U23689 (N_23689,N_14888,N_15524);
or U23690 (N_23690,N_13417,N_14931);
or U23691 (N_23691,N_12016,N_14586);
nand U23692 (N_23692,N_12917,N_16690);
or U23693 (N_23693,N_14471,N_14587);
or U23694 (N_23694,N_15425,N_13595);
xnor U23695 (N_23695,N_16134,N_12239);
and U23696 (N_23696,N_15645,N_16601);
xnor U23697 (N_23697,N_12965,N_15834);
nand U23698 (N_23698,N_15105,N_12169);
xor U23699 (N_23699,N_15870,N_15610);
and U23700 (N_23700,N_13129,N_14533);
nor U23701 (N_23701,N_13116,N_17200);
and U23702 (N_23702,N_14470,N_13396);
nand U23703 (N_23703,N_16674,N_17986);
and U23704 (N_23704,N_12074,N_12601);
and U23705 (N_23705,N_14907,N_15583);
nand U23706 (N_23706,N_16951,N_16235);
nand U23707 (N_23707,N_15220,N_15300);
nor U23708 (N_23708,N_15412,N_16674);
and U23709 (N_23709,N_13337,N_17274);
nor U23710 (N_23710,N_16551,N_15928);
or U23711 (N_23711,N_15210,N_12045);
and U23712 (N_23712,N_17099,N_12145);
or U23713 (N_23713,N_16752,N_12601);
xnor U23714 (N_23714,N_14309,N_16946);
nor U23715 (N_23715,N_13528,N_14955);
nand U23716 (N_23716,N_17407,N_17004);
nand U23717 (N_23717,N_14454,N_12525);
or U23718 (N_23718,N_16291,N_16726);
xnor U23719 (N_23719,N_16817,N_15666);
nor U23720 (N_23720,N_12943,N_17919);
xnor U23721 (N_23721,N_17657,N_12369);
nand U23722 (N_23722,N_16269,N_16291);
nand U23723 (N_23723,N_13219,N_14542);
and U23724 (N_23724,N_17942,N_15937);
and U23725 (N_23725,N_14261,N_15354);
nand U23726 (N_23726,N_14121,N_17229);
nor U23727 (N_23727,N_12572,N_14502);
and U23728 (N_23728,N_15797,N_17664);
xnor U23729 (N_23729,N_15705,N_15367);
nand U23730 (N_23730,N_13426,N_13660);
xor U23731 (N_23731,N_14634,N_14317);
xnor U23732 (N_23732,N_15585,N_14511);
xor U23733 (N_23733,N_12378,N_12092);
nand U23734 (N_23734,N_14861,N_17257);
nand U23735 (N_23735,N_15293,N_13315);
or U23736 (N_23736,N_16940,N_14417);
or U23737 (N_23737,N_14193,N_13130);
and U23738 (N_23738,N_13266,N_15037);
nor U23739 (N_23739,N_15126,N_14054);
or U23740 (N_23740,N_12710,N_12809);
xor U23741 (N_23741,N_16820,N_15148);
xnor U23742 (N_23742,N_15335,N_16042);
nor U23743 (N_23743,N_13809,N_13023);
nand U23744 (N_23744,N_12438,N_14257);
xnor U23745 (N_23745,N_12817,N_15305);
or U23746 (N_23746,N_16609,N_17634);
nor U23747 (N_23747,N_16140,N_13943);
or U23748 (N_23748,N_12504,N_14937);
or U23749 (N_23749,N_17865,N_13469);
and U23750 (N_23750,N_14097,N_15822);
nor U23751 (N_23751,N_12894,N_14479);
and U23752 (N_23752,N_17496,N_15817);
or U23753 (N_23753,N_17236,N_15752);
and U23754 (N_23754,N_12320,N_16499);
or U23755 (N_23755,N_16204,N_13075);
nand U23756 (N_23756,N_14679,N_17531);
nand U23757 (N_23757,N_17897,N_15268);
or U23758 (N_23758,N_13499,N_15114);
nand U23759 (N_23759,N_13324,N_13243);
or U23760 (N_23760,N_15418,N_17716);
nand U23761 (N_23761,N_15409,N_17899);
and U23762 (N_23762,N_17956,N_14142);
nor U23763 (N_23763,N_12316,N_13979);
nor U23764 (N_23764,N_15313,N_16167);
and U23765 (N_23765,N_16030,N_17665);
nand U23766 (N_23766,N_12566,N_15020);
and U23767 (N_23767,N_17041,N_14694);
nor U23768 (N_23768,N_14733,N_14011);
or U23769 (N_23769,N_14116,N_16534);
and U23770 (N_23770,N_12893,N_14469);
nor U23771 (N_23771,N_17455,N_13677);
xnor U23772 (N_23772,N_17401,N_15870);
nor U23773 (N_23773,N_17481,N_14729);
or U23774 (N_23774,N_13424,N_15517);
xnor U23775 (N_23775,N_15529,N_12242);
nor U23776 (N_23776,N_17145,N_13366);
and U23777 (N_23777,N_15823,N_16241);
nor U23778 (N_23778,N_14699,N_16183);
and U23779 (N_23779,N_12268,N_12426);
and U23780 (N_23780,N_13501,N_16553);
nand U23781 (N_23781,N_15239,N_15846);
nor U23782 (N_23782,N_12432,N_16045);
nor U23783 (N_23783,N_13935,N_14000);
or U23784 (N_23784,N_17023,N_14845);
or U23785 (N_23785,N_17310,N_15706);
or U23786 (N_23786,N_15806,N_15513);
nor U23787 (N_23787,N_14753,N_15278);
nand U23788 (N_23788,N_13597,N_17238);
and U23789 (N_23789,N_13228,N_12236);
nand U23790 (N_23790,N_15349,N_14254);
or U23791 (N_23791,N_16156,N_13476);
xnor U23792 (N_23792,N_16252,N_17289);
nor U23793 (N_23793,N_14078,N_13971);
or U23794 (N_23794,N_17397,N_13981);
xor U23795 (N_23795,N_16273,N_15811);
or U23796 (N_23796,N_12941,N_12898);
xor U23797 (N_23797,N_17950,N_15599);
or U23798 (N_23798,N_15996,N_17963);
nor U23799 (N_23799,N_15134,N_13679);
and U23800 (N_23800,N_16801,N_13871);
and U23801 (N_23801,N_13380,N_16347);
xnor U23802 (N_23802,N_17753,N_12109);
nand U23803 (N_23803,N_13316,N_14574);
or U23804 (N_23804,N_12785,N_16109);
and U23805 (N_23805,N_16359,N_13332);
or U23806 (N_23806,N_13750,N_12100);
and U23807 (N_23807,N_16215,N_12042);
nor U23808 (N_23808,N_17907,N_15961);
nor U23809 (N_23809,N_12469,N_16948);
or U23810 (N_23810,N_12276,N_12114);
nor U23811 (N_23811,N_17953,N_15729);
and U23812 (N_23812,N_13086,N_12296);
and U23813 (N_23813,N_15519,N_15039);
nand U23814 (N_23814,N_16436,N_17176);
and U23815 (N_23815,N_14140,N_13442);
xor U23816 (N_23816,N_14069,N_17345);
nor U23817 (N_23817,N_17215,N_15156);
and U23818 (N_23818,N_13989,N_17104);
or U23819 (N_23819,N_13653,N_13697);
or U23820 (N_23820,N_14857,N_17247);
xnor U23821 (N_23821,N_12550,N_17098);
xor U23822 (N_23822,N_16179,N_15718);
and U23823 (N_23823,N_14668,N_16345);
nor U23824 (N_23824,N_15704,N_13177);
nand U23825 (N_23825,N_17530,N_13912);
nand U23826 (N_23826,N_17988,N_12115);
xnor U23827 (N_23827,N_17157,N_13408);
nor U23828 (N_23828,N_17787,N_15627);
nor U23829 (N_23829,N_17810,N_12719);
nand U23830 (N_23830,N_14903,N_17671);
nor U23831 (N_23831,N_12903,N_15584);
nand U23832 (N_23832,N_17654,N_17463);
or U23833 (N_23833,N_14624,N_15108);
and U23834 (N_23834,N_14449,N_16359);
and U23835 (N_23835,N_15793,N_12059);
xor U23836 (N_23836,N_12687,N_17138);
nand U23837 (N_23837,N_16426,N_16765);
and U23838 (N_23838,N_15148,N_17813);
nor U23839 (N_23839,N_14103,N_17094);
xnor U23840 (N_23840,N_17606,N_14670);
or U23841 (N_23841,N_16475,N_13267);
or U23842 (N_23842,N_14503,N_16136);
or U23843 (N_23843,N_14744,N_12254);
xor U23844 (N_23844,N_16982,N_17730);
nor U23845 (N_23845,N_17076,N_13801);
nand U23846 (N_23846,N_14674,N_15680);
and U23847 (N_23847,N_14658,N_17460);
or U23848 (N_23848,N_12984,N_17353);
xor U23849 (N_23849,N_15767,N_13882);
xnor U23850 (N_23850,N_17261,N_16393);
xor U23851 (N_23851,N_15181,N_12414);
nor U23852 (N_23852,N_16756,N_16341);
and U23853 (N_23853,N_17277,N_15495);
xor U23854 (N_23854,N_14532,N_14422);
or U23855 (N_23855,N_13396,N_16506);
nor U23856 (N_23856,N_12812,N_13719);
or U23857 (N_23857,N_14881,N_15392);
nor U23858 (N_23858,N_13180,N_13893);
and U23859 (N_23859,N_14037,N_16012);
or U23860 (N_23860,N_16057,N_17252);
nor U23861 (N_23861,N_15810,N_14613);
nor U23862 (N_23862,N_17801,N_13968);
xor U23863 (N_23863,N_15287,N_16211);
nor U23864 (N_23864,N_14328,N_14165);
and U23865 (N_23865,N_16245,N_13019);
or U23866 (N_23866,N_17782,N_15807);
xor U23867 (N_23867,N_12932,N_16080);
or U23868 (N_23868,N_15486,N_15452);
and U23869 (N_23869,N_15885,N_17431);
nor U23870 (N_23870,N_14258,N_14605);
and U23871 (N_23871,N_14431,N_15943);
nor U23872 (N_23872,N_17467,N_13050);
nand U23873 (N_23873,N_14015,N_15883);
nand U23874 (N_23874,N_16636,N_14632);
nand U23875 (N_23875,N_17688,N_15592);
nor U23876 (N_23876,N_13674,N_16750);
or U23877 (N_23877,N_17920,N_15278);
nor U23878 (N_23878,N_13687,N_16376);
nand U23879 (N_23879,N_12766,N_13784);
xor U23880 (N_23880,N_16914,N_17689);
xnor U23881 (N_23881,N_16222,N_16374);
and U23882 (N_23882,N_13655,N_14809);
nand U23883 (N_23883,N_17607,N_12154);
or U23884 (N_23884,N_15503,N_14820);
and U23885 (N_23885,N_16587,N_17106);
nor U23886 (N_23886,N_12232,N_17662);
and U23887 (N_23887,N_13111,N_12555);
and U23888 (N_23888,N_13129,N_16549);
or U23889 (N_23889,N_17294,N_17924);
and U23890 (N_23890,N_12843,N_12218);
nor U23891 (N_23891,N_13006,N_17035);
or U23892 (N_23892,N_14165,N_14383);
and U23893 (N_23893,N_14834,N_12903);
nand U23894 (N_23894,N_12772,N_12197);
and U23895 (N_23895,N_15012,N_15912);
xor U23896 (N_23896,N_16334,N_15904);
and U23897 (N_23897,N_15441,N_13718);
or U23898 (N_23898,N_16136,N_14816);
nand U23899 (N_23899,N_14713,N_17213);
nand U23900 (N_23900,N_15538,N_13195);
and U23901 (N_23901,N_16342,N_16649);
and U23902 (N_23902,N_16488,N_17413);
nor U23903 (N_23903,N_12606,N_15673);
nor U23904 (N_23904,N_15393,N_13309);
and U23905 (N_23905,N_14586,N_17670);
or U23906 (N_23906,N_15418,N_14452);
nand U23907 (N_23907,N_15080,N_15436);
nand U23908 (N_23908,N_16633,N_16691);
xnor U23909 (N_23909,N_15970,N_17191);
nand U23910 (N_23910,N_12572,N_13375);
xnor U23911 (N_23911,N_13885,N_12926);
or U23912 (N_23912,N_12790,N_15039);
nand U23913 (N_23913,N_12590,N_14672);
xor U23914 (N_23914,N_13276,N_12040);
nand U23915 (N_23915,N_17208,N_14004);
nor U23916 (N_23916,N_14247,N_13049);
or U23917 (N_23917,N_16351,N_16779);
or U23918 (N_23918,N_13906,N_16638);
and U23919 (N_23919,N_16488,N_14815);
or U23920 (N_23920,N_15755,N_15713);
or U23921 (N_23921,N_12223,N_17733);
xnor U23922 (N_23922,N_12793,N_14331);
or U23923 (N_23923,N_15814,N_15397);
nor U23924 (N_23924,N_16146,N_13491);
and U23925 (N_23925,N_16474,N_16490);
xor U23926 (N_23926,N_14147,N_15755);
or U23927 (N_23927,N_14508,N_15904);
xor U23928 (N_23928,N_14807,N_15368);
nand U23929 (N_23929,N_17706,N_14458);
or U23930 (N_23930,N_17605,N_13051);
xnor U23931 (N_23931,N_17273,N_12725);
nand U23932 (N_23932,N_16486,N_12698);
or U23933 (N_23933,N_13592,N_15483);
or U23934 (N_23934,N_13808,N_14178);
nand U23935 (N_23935,N_13508,N_13127);
xor U23936 (N_23936,N_16713,N_14782);
xor U23937 (N_23937,N_17437,N_15831);
or U23938 (N_23938,N_17243,N_16586);
and U23939 (N_23939,N_17263,N_15003);
nand U23940 (N_23940,N_14376,N_13923);
xnor U23941 (N_23941,N_15515,N_16658);
xnor U23942 (N_23942,N_16081,N_14667);
nor U23943 (N_23943,N_16602,N_14830);
xnor U23944 (N_23944,N_17360,N_14590);
or U23945 (N_23945,N_12209,N_16722);
or U23946 (N_23946,N_17593,N_14472);
xnor U23947 (N_23947,N_14895,N_15801);
xor U23948 (N_23948,N_15110,N_14461);
and U23949 (N_23949,N_15057,N_17003);
and U23950 (N_23950,N_17375,N_15889);
or U23951 (N_23951,N_15272,N_13044);
or U23952 (N_23952,N_12960,N_16401);
nor U23953 (N_23953,N_12773,N_13506);
xor U23954 (N_23954,N_17722,N_15244);
nor U23955 (N_23955,N_14954,N_13889);
or U23956 (N_23956,N_17543,N_15692);
or U23957 (N_23957,N_16792,N_17236);
xor U23958 (N_23958,N_17666,N_12275);
or U23959 (N_23959,N_14589,N_13877);
nor U23960 (N_23960,N_17121,N_12639);
nor U23961 (N_23961,N_17590,N_14892);
nor U23962 (N_23962,N_15262,N_14453);
or U23963 (N_23963,N_15160,N_17684);
and U23964 (N_23964,N_16735,N_12696);
and U23965 (N_23965,N_14378,N_16127);
and U23966 (N_23966,N_12978,N_12599);
xor U23967 (N_23967,N_15891,N_13972);
or U23968 (N_23968,N_12406,N_17573);
or U23969 (N_23969,N_12386,N_12074);
and U23970 (N_23970,N_12837,N_15704);
nor U23971 (N_23971,N_17029,N_14823);
nand U23972 (N_23972,N_16360,N_12922);
xor U23973 (N_23973,N_13997,N_16713);
nand U23974 (N_23974,N_17192,N_13834);
xnor U23975 (N_23975,N_14357,N_16404);
or U23976 (N_23976,N_15761,N_15830);
nor U23977 (N_23977,N_13928,N_17868);
or U23978 (N_23978,N_12266,N_13199);
nand U23979 (N_23979,N_12269,N_13765);
nand U23980 (N_23980,N_17290,N_15644);
nand U23981 (N_23981,N_17143,N_17136);
xor U23982 (N_23982,N_14327,N_12917);
nand U23983 (N_23983,N_17755,N_12031);
nor U23984 (N_23984,N_16899,N_17915);
xnor U23985 (N_23985,N_12607,N_13709);
nand U23986 (N_23986,N_15214,N_12457);
nand U23987 (N_23987,N_13434,N_12022);
and U23988 (N_23988,N_13093,N_15742);
or U23989 (N_23989,N_17715,N_14560);
xor U23990 (N_23990,N_12558,N_14293);
nand U23991 (N_23991,N_15709,N_17986);
and U23992 (N_23992,N_17212,N_14658);
nand U23993 (N_23993,N_15907,N_16163);
nor U23994 (N_23994,N_17860,N_16234);
or U23995 (N_23995,N_16090,N_12343);
nand U23996 (N_23996,N_16275,N_12307);
xor U23997 (N_23997,N_14716,N_15310);
and U23998 (N_23998,N_14477,N_16190);
or U23999 (N_23999,N_14737,N_17999);
xor U24000 (N_24000,N_18731,N_19833);
and U24001 (N_24001,N_22594,N_23077);
and U24002 (N_24002,N_18978,N_22628);
nor U24003 (N_24003,N_22929,N_22902);
or U24004 (N_24004,N_20415,N_21841);
or U24005 (N_24005,N_22647,N_18326);
nor U24006 (N_24006,N_21181,N_18093);
and U24007 (N_24007,N_22466,N_23487);
nand U24008 (N_24008,N_19824,N_18290);
xor U24009 (N_24009,N_22931,N_22437);
nor U24010 (N_24010,N_22955,N_21222);
xnor U24011 (N_24011,N_18234,N_19009);
or U24012 (N_24012,N_23766,N_21720);
nand U24013 (N_24013,N_18128,N_18944);
xnor U24014 (N_24014,N_18140,N_23179);
nand U24015 (N_24015,N_18425,N_22361);
and U24016 (N_24016,N_18231,N_20658);
and U24017 (N_24017,N_19523,N_21646);
xor U24018 (N_24018,N_20717,N_20984);
nor U24019 (N_24019,N_20331,N_23217);
nor U24020 (N_24020,N_22606,N_18984);
and U24021 (N_24021,N_18262,N_22401);
xor U24022 (N_24022,N_21159,N_21191);
or U24023 (N_24023,N_20412,N_23801);
nand U24024 (N_24024,N_22014,N_20048);
and U24025 (N_24025,N_19881,N_18903);
nand U24026 (N_24026,N_18412,N_21826);
xor U24027 (N_24027,N_19567,N_21232);
nand U24028 (N_24028,N_19400,N_22362);
nand U24029 (N_24029,N_22152,N_18213);
nand U24030 (N_24030,N_19304,N_20535);
or U24031 (N_24031,N_19301,N_20038);
nor U24032 (N_24032,N_20343,N_19158);
xor U24033 (N_24033,N_22516,N_21060);
nand U24034 (N_24034,N_20792,N_23853);
nand U24035 (N_24035,N_23352,N_22118);
xor U24036 (N_24036,N_19163,N_18301);
or U24037 (N_24037,N_18765,N_18468);
nor U24038 (N_24038,N_18586,N_23159);
or U24039 (N_24039,N_20114,N_21581);
or U24040 (N_24040,N_22618,N_20126);
or U24041 (N_24041,N_23274,N_18693);
nand U24042 (N_24042,N_23640,N_23484);
nand U24043 (N_24043,N_19593,N_22589);
or U24044 (N_24044,N_19219,N_22866);
nand U24045 (N_24045,N_18293,N_19021);
xnor U24046 (N_24046,N_20312,N_23943);
nand U24047 (N_24047,N_18806,N_20565);
nand U24048 (N_24048,N_21196,N_19760);
nand U24049 (N_24049,N_19726,N_18799);
and U24050 (N_24050,N_21344,N_21270);
nor U24051 (N_24051,N_22002,N_19141);
nand U24052 (N_24052,N_22204,N_23239);
nor U24053 (N_24053,N_19595,N_18993);
or U24054 (N_24054,N_23224,N_19637);
nand U24055 (N_24055,N_22764,N_21388);
and U24056 (N_24056,N_22781,N_18171);
nand U24057 (N_24057,N_22649,N_20944);
or U24058 (N_24058,N_22693,N_20327);
xor U24059 (N_24059,N_21948,N_21884);
and U24060 (N_24060,N_18461,N_18168);
nand U24061 (N_24061,N_21278,N_22735);
nand U24062 (N_24062,N_19641,N_21850);
xnor U24063 (N_24063,N_19214,N_18871);
xnor U24064 (N_24064,N_22135,N_20386);
nand U24065 (N_24065,N_23592,N_18682);
xnor U24066 (N_24066,N_18013,N_20716);
or U24067 (N_24067,N_19585,N_23229);
or U24068 (N_24068,N_18417,N_22938);
nor U24069 (N_24069,N_22733,N_23886);
nand U24070 (N_24070,N_20437,N_18732);
xnor U24071 (N_24071,N_21048,N_18325);
nor U24072 (N_24072,N_22293,N_22311);
and U24073 (N_24073,N_19771,N_20270);
nor U24074 (N_24074,N_20684,N_22245);
and U24075 (N_24075,N_21978,N_18440);
xnor U24076 (N_24076,N_20598,N_23090);
xnor U24077 (N_24077,N_23845,N_21102);
or U24078 (N_24078,N_21992,N_23339);
nor U24079 (N_24079,N_19081,N_22302);
and U24080 (N_24080,N_21951,N_20674);
nand U24081 (N_24081,N_23325,N_22831);
or U24082 (N_24082,N_21925,N_23702);
nor U24083 (N_24083,N_18380,N_20215);
and U24084 (N_24084,N_20006,N_19413);
or U24085 (N_24085,N_23662,N_23779);
nand U24086 (N_24086,N_18343,N_20457);
xor U24087 (N_24087,N_18888,N_18609);
xnor U24088 (N_24088,N_19457,N_21307);
or U24089 (N_24089,N_19763,N_19189);
or U24090 (N_24090,N_23740,N_18037);
and U24091 (N_24091,N_22111,N_23467);
xor U24092 (N_24092,N_22000,N_19484);
or U24093 (N_24093,N_18347,N_18579);
or U24094 (N_24094,N_19607,N_21084);
or U24095 (N_24095,N_18865,N_21195);
and U24096 (N_24096,N_20683,N_18083);
and U24097 (N_24097,N_19472,N_23656);
nand U24098 (N_24098,N_20851,N_21299);
or U24099 (N_24099,N_18740,N_19737);
or U24100 (N_24100,N_21888,N_19370);
xnor U24101 (N_24101,N_18349,N_19900);
or U24102 (N_24102,N_21397,N_22853);
xnor U24103 (N_24103,N_23628,N_19330);
or U24104 (N_24104,N_21249,N_18334);
xor U24105 (N_24105,N_19112,N_21557);
and U24106 (N_24106,N_21027,N_18738);
nor U24107 (N_24107,N_20118,N_21979);
and U24108 (N_24108,N_22230,N_20795);
and U24109 (N_24109,N_19405,N_23583);
nor U24110 (N_24110,N_19530,N_18775);
and U24111 (N_24111,N_20209,N_19804);
xor U24112 (N_24112,N_19398,N_20157);
and U24113 (N_24113,N_21303,N_23660);
nand U24114 (N_24114,N_18381,N_23303);
nor U24115 (N_24115,N_19409,N_21173);
nor U24116 (N_24116,N_18906,N_18991);
or U24117 (N_24117,N_20772,N_22464);
or U24118 (N_24118,N_21106,N_19799);
nor U24119 (N_24119,N_23675,N_19871);
or U24120 (N_24120,N_18717,N_20849);
xnor U24121 (N_24121,N_21927,N_22462);
nor U24122 (N_24122,N_22829,N_20340);
nor U24123 (N_24123,N_18031,N_19351);
nor U24124 (N_24124,N_21785,N_20621);
or U24125 (N_24125,N_22818,N_19019);
xor U24126 (N_24126,N_22729,N_20862);
nand U24127 (N_24127,N_20787,N_19912);
nor U24128 (N_24128,N_23896,N_19551);
xor U24129 (N_24129,N_22890,N_22834);
xor U24130 (N_24130,N_18627,N_23335);
nor U24131 (N_24131,N_18421,N_23361);
or U24132 (N_24132,N_23389,N_23259);
xor U24133 (N_24133,N_18721,N_23541);
and U24134 (N_24134,N_20810,N_19806);
nor U24135 (N_24135,N_21513,N_22832);
nor U24136 (N_24136,N_21440,N_19849);
nand U24137 (N_24137,N_18921,N_23122);
xnor U24138 (N_24138,N_18813,N_21832);
nor U24139 (N_24139,N_20866,N_19324);
xor U24140 (N_24140,N_21748,N_23499);
nand U24141 (N_24141,N_18176,N_23071);
xnor U24142 (N_24142,N_22080,N_22292);
and U24143 (N_24143,N_23643,N_21004);
or U24144 (N_24144,N_20274,N_18265);
nor U24145 (N_24145,N_19436,N_20328);
xnor U24146 (N_24146,N_22461,N_21620);
and U24147 (N_24147,N_19942,N_20891);
nor U24148 (N_24148,N_22752,N_23986);
or U24149 (N_24149,N_22428,N_21330);
nand U24150 (N_24150,N_19181,N_23859);
nor U24151 (N_24151,N_21914,N_23203);
nor U24152 (N_24152,N_21063,N_18306);
xor U24153 (N_24153,N_22430,N_20617);
nor U24154 (N_24154,N_22574,N_23852);
or U24155 (N_24155,N_19596,N_22003);
nand U24156 (N_24156,N_22656,N_19521);
xor U24157 (N_24157,N_19820,N_19783);
and U24158 (N_24158,N_21648,N_18597);
and U24159 (N_24159,N_18174,N_20148);
xor U24160 (N_24160,N_23510,N_19801);
and U24161 (N_24161,N_19227,N_21714);
or U24162 (N_24162,N_22728,N_22793);
or U24163 (N_24163,N_18870,N_18324);
and U24164 (N_24164,N_18418,N_21057);
xnor U24165 (N_24165,N_19561,N_18822);
and U24166 (N_24166,N_23447,N_19813);
nand U24167 (N_24167,N_22185,N_22256);
nor U24168 (N_24168,N_20175,N_18605);
nor U24169 (N_24169,N_18848,N_19188);
nand U24170 (N_24170,N_22774,N_23584);
nand U24171 (N_24171,N_20171,N_23772);
or U24172 (N_24172,N_18021,N_21120);
and U24173 (N_24173,N_23863,N_23915);
xnor U24174 (N_24174,N_19240,N_19468);
xor U24175 (N_24175,N_21685,N_23210);
or U24176 (N_24176,N_23815,N_20162);
nor U24177 (N_24177,N_23514,N_22335);
nor U24178 (N_24178,N_22605,N_23644);
and U24179 (N_24179,N_20623,N_18785);
nand U24180 (N_24180,N_21917,N_22154);
nor U24181 (N_24181,N_18518,N_23212);
or U24182 (N_24182,N_23101,N_18669);
xnor U24183 (N_24183,N_22388,N_21010);
and U24184 (N_24184,N_19314,N_21151);
xnor U24185 (N_24185,N_21877,N_21259);
xor U24186 (N_24186,N_22346,N_23348);
and U24187 (N_24187,N_18164,N_19842);
xnor U24188 (N_24188,N_19583,N_18635);
or U24189 (N_24189,N_21313,N_23561);
nand U24190 (N_24190,N_23028,N_19446);
nand U24191 (N_24191,N_21852,N_20149);
and U24192 (N_24192,N_23918,N_20092);
or U24193 (N_24193,N_19213,N_19111);
nand U24194 (N_24194,N_23084,N_23106);
nand U24195 (N_24195,N_23835,N_21198);
nand U24196 (N_24196,N_21326,N_22508);
nand U24197 (N_24197,N_21081,N_20050);
xor U24198 (N_24198,N_20473,N_23051);
nor U24199 (N_24199,N_18291,N_21954);
xor U24200 (N_24200,N_18153,N_21752);
nand U24201 (N_24201,N_18481,N_22963);
or U24202 (N_24202,N_20797,N_23301);
xnor U24203 (N_24203,N_23578,N_18216);
and U24204 (N_24204,N_21290,N_23385);
and U24205 (N_24205,N_22059,N_23962);
or U24206 (N_24206,N_23802,N_20714);
nand U24207 (N_24207,N_22526,N_21491);
xor U24208 (N_24208,N_23354,N_19401);
xnor U24209 (N_24209,N_19461,N_18986);
nand U24210 (N_24210,N_20534,N_18695);
nor U24211 (N_24211,N_19016,N_23668);
or U24212 (N_24212,N_22912,N_20697);
nor U24213 (N_24213,N_23572,N_18646);
nor U24214 (N_24214,N_23450,N_23518);
or U24215 (N_24215,N_20817,N_20715);
or U24216 (N_24216,N_20291,N_20545);
xor U24217 (N_24217,N_20301,N_22104);
nor U24218 (N_24218,N_22144,N_21035);
nand U24219 (N_24219,N_19389,N_23594);
or U24220 (N_24220,N_18444,N_23092);
xor U24221 (N_24221,N_20221,N_18295);
nand U24222 (N_24222,N_19495,N_20601);
xor U24223 (N_24223,N_22398,N_21508);
xnor U24224 (N_24224,N_21835,N_19078);
nand U24225 (N_24225,N_23520,N_18655);
and U24226 (N_24226,N_18115,N_19095);
xnor U24227 (N_24227,N_19230,N_21241);
nand U24228 (N_24228,N_18482,N_23650);
or U24229 (N_24229,N_22253,N_18555);
or U24230 (N_24230,N_21506,N_22572);
or U24231 (N_24231,N_19173,N_21127);
and U24232 (N_24232,N_21972,N_18100);
xnor U24233 (N_24233,N_18413,N_18471);
xnor U24234 (N_24234,N_21940,N_19253);
or U24235 (N_24235,N_20916,N_23190);
nand U24236 (N_24236,N_23688,N_23708);
or U24237 (N_24237,N_20678,N_21495);
nor U24238 (N_24238,N_21148,N_18652);
nand U24239 (N_24239,N_19149,N_19030);
and U24240 (N_24240,N_21235,N_20699);
or U24241 (N_24241,N_19348,N_19500);
nand U24242 (N_24242,N_22157,N_20177);
nand U24243 (N_24243,N_21336,N_20094);
xnor U24244 (N_24244,N_21580,N_20831);
nor U24245 (N_24245,N_21309,N_18948);
and U24246 (N_24246,N_21398,N_18263);
and U24247 (N_24247,N_18648,N_21369);
nor U24248 (N_24248,N_20317,N_21414);
and U24249 (N_24249,N_20285,N_22262);
and U24250 (N_24250,N_23933,N_19805);
nor U24251 (N_24251,N_18369,N_20346);
and U24252 (N_24252,N_22261,N_23832);
xnor U24253 (N_24253,N_19283,N_23817);
xnor U24254 (N_24254,N_23654,N_20250);
or U24255 (N_24255,N_19822,N_20021);
and U24256 (N_24256,N_23007,N_21983);
xnor U24257 (N_24257,N_19717,N_20139);
nand U24258 (N_24258,N_19200,N_20975);
or U24259 (N_24259,N_20144,N_23938);
and U24260 (N_24260,N_21759,N_20252);
xnor U24261 (N_24261,N_22962,N_22721);
or U24262 (N_24262,N_18243,N_18708);
xor U24263 (N_24263,N_22331,N_21026);
xor U24264 (N_24264,N_22786,N_23983);
nor U24265 (N_24265,N_22778,N_21650);
and U24266 (N_24266,N_22484,N_21087);
and U24267 (N_24267,N_22994,N_22737);
nor U24268 (N_24268,N_19210,N_20937);
or U24269 (N_24269,N_22524,N_18182);
and U24270 (N_24270,N_20142,N_22825);
xor U24271 (N_24271,N_23439,N_23011);
nand U24272 (N_24272,N_22474,N_18284);
and U24273 (N_24273,N_20326,N_19483);
nand U24274 (N_24274,N_18667,N_19302);
nor U24275 (N_24275,N_22493,N_19627);
and U24276 (N_24276,N_21923,N_23449);
nand U24277 (N_24277,N_21565,N_22378);
nand U24278 (N_24278,N_23907,N_22250);
xor U24279 (N_24279,N_19733,N_21392);
or U24280 (N_24280,N_18055,N_18023);
nor U24281 (N_24281,N_23649,N_19925);
nor U24282 (N_24282,N_23707,N_23037);
or U24283 (N_24283,N_22838,N_21510);
xnor U24284 (N_24284,N_20962,N_19543);
xor U24285 (N_24285,N_20485,N_20593);
xor U24286 (N_24286,N_22951,N_19242);
and U24287 (N_24287,N_20650,N_23277);
xnor U24288 (N_24288,N_20664,N_22323);
nand U24289 (N_24289,N_20675,N_22556);
xor U24290 (N_24290,N_23889,N_23836);
xor U24291 (N_24291,N_20219,N_23999);
and U24292 (N_24292,N_22449,N_20248);
xor U24293 (N_24293,N_19212,N_21422);
and U24294 (N_24294,N_19557,N_21089);
nand U24295 (N_24295,N_19877,N_21962);
xor U24296 (N_24296,N_23704,N_20348);
and U24297 (N_24297,N_21533,N_19671);
nor U24298 (N_24298,N_18286,N_23284);
or U24299 (N_24299,N_19698,N_23042);
nor U24300 (N_24300,N_22149,N_18416);
nor U24301 (N_24301,N_19266,N_21047);
and U24302 (N_24302,N_18882,N_21994);
or U24303 (N_24303,N_22222,N_19318);
nor U24304 (N_24304,N_19657,N_19037);
and U24305 (N_24305,N_19613,N_20635);
xnor U24306 (N_24306,N_23305,N_22661);
xnor U24307 (N_24307,N_23838,N_23356);
or U24308 (N_24308,N_20324,N_20434);
and U24309 (N_24309,N_20035,N_19829);
nor U24310 (N_24310,N_23368,N_21690);
or U24311 (N_24311,N_23876,N_22382);
xor U24312 (N_24312,N_19375,N_22209);
and U24313 (N_24313,N_20280,N_23590);
or U24314 (N_24314,N_19152,N_20199);
nor U24315 (N_24315,N_18762,N_22117);
and U24316 (N_24316,N_20237,N_21211);
or U24317 (N_24317,N_20395,N_23266);
nand U24318 (N_24318,N_21781,N_22132);
nor U24319 (N_24319,N_22566,N_21499);
nor U24320 (N_24320,N_20741,N_23940);
and U24321 (N_24321,N_19395,N_22455);
and U24322 (N_24322,N_23846,N_22543);
nand U24323 (N_24323,N_20159,N_18119);
or U24324 (N_24324,N_22568,N_20080);
xnor U24325 (N_24325,N_23534,N_18887);
nor U24326 (N_24326,N_18159,N_20709);
nor U24327 (N_24327,N_23196,N_23908);
nor U24328 (N_24328,N_21522,N_23755);
xnor U24329 (N_24329,N_22620,N_18607);
nand U24330 (N_24330,N_20712,N_23519);
xor U24331 (N_24331,N_23105,N_20099);
nand U24332 (N_24332,N_23235,N_23782);
and U24333 (N_24333,N_23155,N_18001);
xor U24334 (N_24334,N_23652,N_21054);
or U24335 (N_24335,N_20030,N_22699);
and U24336 (N_24336,N_18217,N_19990);
and U24337 (N_24337,N_21790,N_23016);
or U24338 (N_24338,N_19605,N_21480);
nor U24339 (N_24339,N_18285,N_20400);
or U24340 (N_24340,N_21283,N_20201);
and U24341 (N_24341,N_19216,N_18446);
nor U24342 (N_24342,N_21163,N_22360);
nor U24343 (N_24343,N_23147,N_19044);
xnor U24344 (N_24344,N_18668,N_21433);
nor U24345 (N_24345,N_18014,N_22792);
xnor U24346 (N_24346,N_20961,N_23981);
or U24347 (N_24347,N_19207,N_19178);
nand U24348 (N_24348,N_20034,N_22928);
nand U24349 (N_24349,N_22894,N_22557);
nand U24350 (N_24350,N_23809,N_21217);
or U24351 (N_24351,N_18151,N_18149);
xnor U24352 (N_24352,N_22026,N_18508);
nor U24353 (N_24353,N_23552,N_22807);
nor U24354 (N_24354,N_19006,N_20785);
and U24355 (N_24355,N_18707,N_22217);
nand U24356 (N_24356,N_19451,N_20638);
xor U24357 (N_24357,N_23685,N_18485);
and U24358 (N_24358,N_20679,N_19083);
xor U24359 (N_24359,N_19133,N_21100);
xnor U24360 (N_24360,N_21920,N_19703);
and U24361 (N_24361,N_23635,N_18756);
nand U24362 (N_24362,N_20003,N_18229);
nand U24363 (N_24363,N_21965,N_23083);
nor U24364 (N_24364,N_18615,N_18420);
or U24365 (N_24365,N_22776,N_21518);
or U24366 (N_24366,N_20549,N_20055);
nand U24367 (N_24367,N_18340,N_21589);
xnor U24368 (N_24368,N_23880,N_18356);
or U24369 (N_24369,N_21571,N_19930);
and U24370 (N_24370,N_18506,N_23930);
nor U24371 (N_24371,N_23360,N_21399);
or U24372 (N_24372,N_23837,N_20934);
or U24373 (N_24373,N_21042,N_23587);
or U24374 (N_24374,N_20041,N_23373);
and U24375 (N_24375,N_18666,N_22748);
xnor U24376 (N_24376,N_23285,N_23489);
nor U24377 (N_24377,N_20686,N_20311);
nand U24378 (N_24378,N_20592,N_22422);
and U24379 (N_24379,N_18104,N_18179);
and U24380 (N_24380,N_18298,N_20668);
nand U24381 (N_24381,N_20408,N_19843);
nand U24382 (N_24382,N_21188,N_19923);
xnor U24383 (N_24383,N_19626,N_22800);
xnor U24384 (N_24384,N_22314,N_19208);
nand U24385 (N_24385,N_23425,N_18138);
nand U24386 (N_24386,N_20193,N_18706);
and U24387 (N_24387,N_20267,N_19864);
xnor U24388 (N_24388,N_22050,N_20421);
nand U24389 (N_24389,N_23371,N_21966);
xnor U24390 (N_24390,N_19780,N_22861);
or U24391 (N_24391,N_20854,N_22827);
or U24392 (N_24392,N_21825,N_20472);
nor U24393 (N_24393,N_18452,N_20941);
nor U24394 (N_24394,N_22723,N_21612);
or U24395 (N_24395,N_22761,N_22489);
nor U24396 (N_24396,N_22053,N_19121);
or U24397 (N_24397,N_23351,N_19299);
and U24398 (N_24398,N_21012,N_19182);
and U24399 (N_24399,N_22719,N_18114);
nand U24400 (N_24400,N_22141,N_19416);
nand U24401 (N_24401,N_21238,N_21809);
nand U24402 (N_24402,N_21347,N_22796);
and U24403 (N_24403,N_21981,N_19385);
or U24404 (N_24404,N_22101,N_23446);
xor U24405 (N_24405,N_20737,N_22054);
xor U24406 (N_24406,N_23563,N_23430);
xnor U24407 (N_24407,N_23270,N_23298);
or U24408 (N_24408,N_22582,N_20186);
nand U24409 (N_24409,N_22201,N_22874);
xnor U24410 (N_24410,N_23062,N_23513);
and U24411 (N_24411,N_22034,N_21197);
nor U24412 (N_24412,N_23233,N_23067);
xor U24413 (N_24413,N_18089,N_21097);
nor U24414 (N_24414,N_18257,N_18724);
nand U24415 (N_24415,N_23666,N_23453);
or U24416 (N_24416,N_23040,N_18893);
nand U24417 (N_24417,N_18391,N_18971);
and U24418 (N_24418,N_20163,N_23942);
and U24419 (N_24419,N_23673,N_18253);
nor U24420 (N_24420,N_22757,N_19172);
and U24421 (N_24421,N_19339,N_19345);
nor U24422 (N_24422,N_23615,N_20560);
nor U24423 (N_24423,N_20316,N_20014);
xnor U24424 (N_24424,N_22056,N_19466);
nor U24425 (N_24425,N_19393,N_18337);
nand U24426 (N_24426,N_20747,N_23992);
or U24427 (N_24427,N_22531,N_23681);
or U24428 (N_24428,N_18733,N_23140);
nand U24429 (N_24429,N_18059,N_19408);
and U24430 (N_24430,N_22773,N_22358);
nor U24431 (N_24431,N_19866,N_19480);
and U24432 (N_24432,N_21767,N_19778);
and U24433 (N_24433,N_20085,N_18519);
xor U24434 (N_24434,N_21154,N_20834);
nor U24435 (N_24435,N_19835,N_22751);
or U24436 (N_24436,N_21803,N_18955);
or U24437 (N_24437,N_22161,N_19767);
or U24438 (N_24438,N_20389,N_21339);
nor U24439 (N_24439,N_22944,N_18117);
nand U24440 (N_24440,N_23299,N_22456);
nor U24441 (N_24441,N_22978,N_21267);
nor U24442 (N_24442,N_18538,N_19144);
nor U24443 (N_24443,N_20833,N_23820);
nand U24444 (N_24444,N_19916,N_21955);
or U24445 (N_24445,N_20983,N_18504);
nor U24446 (N_24446,N_18945,N_22642);
nor U24447 (N_24447,N_21432,N_19373);
or U24448 (N_24448,N_23205,N_20302);
or U24449 (N_24449,N_21555,N_21654);
and U24450 (N_24450,N_18010,N_20548);
and U24451 (N_24451,N_23283,N_21056);
nor U24452 (N_24452,N_21618,N_20289);
nor U24453 (N_24453,N_18543,N_22479);
nor U24454 (N_24454,N_22240,N_18297);
xnor U24455 (N_24455,N_22279,N_21221);
xor U24456 (N_24456,N_18791,N_22224);
nand U24457 (N_24457,N_18233,N_20583);
nor U24458 (N_24458,N_21219,N_20122);
xnor U24459 (N_24459,N_18201,N_20543);
nor U24460 (N_24460,N_21740,N_20970);
or U24461 (N_24461,N_22425,N_19546);
nor U24462 (N_24462,N_20682,N_18235);
nor U24463 (N_24463,N_19784,N_23240);
nor U24464 (N_24464,N_19024,N_22775);
and U24465 (N_24465,N_23279,N_22846);
nor U24466 (N_24466,N_20294,N_19802);
nor U24467 (N_24467,N_21611,N_19825);
or U24468 (N_24468,N_23181,N_19071);
nor U24469 (N_24469,N_19744,N_23134);
or U24470 (N_24470,N_22328,N_19659);
and U24471 (N_24471,N_18226,N_23693);
nand U24472 (N_24472,N_18372,N_21601);
nor U24473 (N_24473,N_20380,N_20631);
or U24474 (N_24474,N_18946,N_18102);
or U24475 (N_24475,N_21916,N_21390);
xor U24476 (N_24476,N_23100,N_22913);
xnor U24477 (N_24477,N_18219,N_22924);
nand U24478 (N_24478,N_20812,N_18890);
and U24479 (N_24479,N_21817,N_22885);
and U24480 (N_24480,N_23516,N_23340);
and U24481 (N_24481,N_19211,N_22068);
nor U24482 (N_24482,N_21293,N_19809);
xor U24483 (N_24483,N_18805,N_20403);
xnor U24484 (N_24484,N_19287,N_18645);
or U24485 (N_24485,N_22867,N_21607);
or U24486 (N_24486,N_19128,N_23378);
nand U24487 (N_24487,N_22213,N_22452);
xnor U24488 (N_24488,N_23984,N_19797);
and U24489 (N_24489,N_19988,N_19278);
or U24490 (N_24490,N_22958,N_23794);
nand U24491 (N_24491,N_18815,N_18747);
xnor U24492 (N_24492,N_22547,N_21323);
or U24493 (N_24493,N_22961,N_22105);
nand U24494 (N_24494,N_18981,N_23332);
nor U24495 (N_24495,N_20360,N_19166);
xor U24496 (N_24496,N_21667,N_22463);
nand U24497 (N_24497,N_23202,N_23714);
xnor U24498 (N_24498,N_20663,N_18886);
and U24499 (N_24499,N_23952,N_22264);
nand U24500 (N_24500,N_20208,N_20746);
nand U24501 (N_24501,N_23829,N_23133);
and U24502 (N_24502,N_18510,N_23479);
or U24503 (N_24503,N_20512,N_23677);
nor U24504 (N_24504,N_22259,N_20824);
xnor U24505 (N_24505,N_23504,N_21813);
nor U24506 (N_24506,N_21861,N_23557);
or U24507 (N_24507,N_23443,N_18766);
or U24508 (N_24508,N_21530,N_19445);
and U24509 (N_24509,N_18432,N_23819);
and U24510 (N_24510,N_21507,N_23207);
and U24511 (N_24511,N_18047,N_21797);
nor U24512 (N_24512,N_21367,N_19839);
or U24513 (N_24513,N_22387,N_22943);
nand U24514 (N_24514,N_21125,N_18969);
nand U24515 (N_24515,N_19334,N_22207);
and U24516 (N_24516,N_23760,N_21967);
or U24517 (N_24517,N_22614,N_19929);
nor U24518 (N_24518,N_21157,N_22465);
xor U24519 (N_24519,N_22453,N_20432);
and U24520 (N_24520,N_22438,N_19258);
nand U24521 (N_24521,N_20732,N_21572);
or U24522 (N_24522,N_20758,N_19903);
or U24523 (N_24523,N_20517,N_20275);
nor U24524 (N_24524,N_19552,N_23475);
or U24525 (N_24525,N_20856,N_21335);
nor U24526 (N_24526,N_19708,N_22754);
nor U24527 (N_24527,N_23599,N_19740);
nand U24528 (N_24528,N_19217,N_20224);
and U24529 (N_24529,N_21800,N_19701);
xnor U24530 (N_24530,N_21678,N_20843);
or U24531 (N_24531,N_22629,N_20268);
nor U24532 (N_24532,N_18261,N_20132);
xnor U24533 (N_24533,N_18925,N_23927);
and U24534 (N_24534,N_18036,N_20197);
nand U24535 (N_24535,N_20460,N_22870);
or U24536 (N_24536,N_22544,N_21280);
nor U24537 (N_24537,N_19146,N_18483);
nand U24538 (N_24538,N_23193,N_22784);
and U24539 (N_24539,N_22036,N_20019);
and U24540 (N_24540,N_23642,N_21535);
nand U24541 (N_24541,N_21673,N_22597);
and U24542 (N_24542,N_20662,N_22654);
and U24543 (N_24543,N_22511,N_18474);
xor U24544 (N_24544,N_21041,N_21713);
and U24545 (N_24545,N_22932,N_20243);
or U24546 (N_24546,N_22007,N_23657);
nand U24547 (N_24547,N_23429,N_22653);
or U24548 (N_24548,N_18215,N_19067);
nand U24549 (N_24549,N_18212,N_22083);
xor U24550 (N_24550,N_22226,N_22860);
or U24551 (N_24551,N_23795,N_18591);
and U24552 (N_24552,N_19218,N_19147);
or U24553 (N_24553,N_23956,N_22692);
and U24554 (N_24554,N_21577,N_23018);
nand U24555 (N_24555,N_18469,N_19588);
or U24556 (N_24556,N_21466,N_22095);
xor U24557 (N_24557,N_18647,N_23920);
nand U24558 (N_24558,N_21664,N_20639);
nor U24559 (N_24559,N_22970,N_20943);
xor U24560 (N_24560,N_20829,N_22148);
and U24561 (N_24561,N_19664,N_18786);
xnor U24562 (N_24562,N_23579,N_19406);
nand U24563 (N_24563,N_19841,N_22040);
nor U24564 (N_24564,N_19893,N_22167);
xnor U24565 (N_24565,N_20606,N_18629);
xnor U24566 (N_24566,N_19417,N_18237);
nor U24567 (N_24567,N_22227,N_18496);
and U24568 (N_24568,N_20337,N_19538);
xor U24569 (N_24569,N_21333,N_23793);
xnor U24570 (N_24570,N_20618,N_22016);
xnor U24571 (N_24571,N_20059,N_20037);
and U24572 (N_24572,N_18379,N_22413);
or U24573 (N_24573,N_21421,N_22330);
and U24574 (N_24574,N_21791,N_23086);
nor U24575 (N_24575,N_19886,N_21402);
and U24576 (N_24576,N_20054,N_21327);
and U24577 (N_24577,N_20959,N_19225);
and U24578 (N_24578,N_19658,N_22959);
or U24579 (N_24579,N_21281,N_20012);
and U24580 (N_24580,N_23913,N_19704);
nand U24581 (N_24581,N_19116,N_21452);
nand U24582 (N_24582,N_22948,N_22174);
nor U24583 (N_24583,N_22659,N_21670);
nor U24584 (N_24584,N_20367,N_20546);
xnor U24585 (N_24585,N_23003,N_22713);
or U24586 (N_24586,N_21961,N_22492);
and U24587 (N_24587,N_23576,N_21101);
xnor U24588 (N_24588,N_21123,N_22389);
or U24589 (N_24589,N_23039,N_20755);
and U24590 (N_24590,N_23941,N_18323);
xnor U24591 (N_24591,N_22797,N_20176);
xnor U24592 (N_24592,N_23728,N_19646);
or U24593 (N_24593,N_20731,N_22234);
and U24594 (N_24594,N_20942,N_22611);
or U24595 (N_24595,N_18088,N_20440);
nand U24596 (N_24596,N_20835,N_19844);
or U24597 (N_24597,N_23393,N_18982);
xor U24598 (N_24598,N_22192,N_22027);
xnor U24599 (N_24599,N_22880,N_23286);
or U24600 (N_24600,N_19562,N_20043);
xor U24601 (N_24601,N_19296,N_22646);
and U24602 (N_24602,N_23789,N_22716);
nor U24603 (N_24603,N_21512,N_21150);
nor U24604 (N_24604,N_19108,N_20932);
xnor U24605 (N_24605,N_21723,N_19630);
nor U24606 (N_24606,N_19870,N_22790);
nor U24607 (N_24607,N_23517,N_19404);
nor U24608 (N_24608,N_20123,N_21700);
nand U24609 (N_24609,N_23197,N_18292);
nor U24610 (N_24610,N_18409,N_21420);
nand U24611 (N_24611,N_22889,N_22717);
nand U24612 (N_24612,N_20116,N_21822);
nor U24613 (N_24613,N_23870,N_18875);
nand U24614 (N_24614,N_19196,N_20161);
or U24615 (N_24615,N_19695,N_19911);
xor U24616 (N_24616,N_23770,N_21078);
nor U24617 (N_24617,N_22617,N_23209);
xor U24618 (N_24618,N_23168,N_18502);
xor U24619 (N_24619,N_19859,N_23616);
and U24620 (N_24620,N_22475,N_23738);
nand U24621 (N_24621,N_20134,N_20595);
nand U24622 (N_24622,N_19510,N_20318);
and U24623 (N_24623,N_19553,N_21540);
or U24624 (N_24624,N_22496,N_23231);
nor U24625 (N_24625,N_19969,N_20053);
or U24626 (N_24626,N_21756,N_21735);
nand U24627 (N_24627,N_18384,N_21856);
and U24628 (N_24628,N_19935,N_21444);
and U24629 (N_24629,N_18961,N_21069);
nand U24630 (N_24630,N_23024,N_23383);
nor U24631 (N_24631,N_19335,N_23626);
xnor U24632 (N_24632,N_21739,N_22412);
or U24633 (N_24633,N_18807,N_18715);
nor U24634 (N_24634,N_21694,N_19117);
and U24635 (N_24635,N_23464,N_19966);
and U24636 (N_24636,N_21090,N_20910);
xor U24637 (N_24637,N_21243,N_21400);
nor U24638 (N_24638,N_18689,N_21609);
or U24639 (N_24639,N_22780,N_23800);
or U24640 (N_24640,N_20304,N_20351);
nand U24641 (N_24641,N_22417,N_18095);
xor U24642 (N_24642,N_20153,N_22655);
nor U24643 (N_24643,N_20445,N_21586);
and U24644 (N_24644,N_22826,N_22359);
xnor U24645 (N_24645,N_20469,N_18889);
xor U24646 (N_24646,N_18388,N_19080);
nor U24647 (N_24647,N_23163,N_21606);
nand U24648 (N_24648,N_18433,N_19366);
nand U24649 (N_24649,N_18039,N_23522);
or U24650 (N_24650,N_20661,N_19180);
nor U24651 (N_24651,N_19379,N_18795);
nor U24652 (N_24652,N_20098,N_21705);
nand U24653 (N_24653,N_18983,N_18335);
xor U24654 (N_24654,N_23618,N_22355);
and U24655 (N_24655,N_19968,N_20373);
or U24656 (N_24656,N_22200,N_20488);
xnor U24657 (N_24657,N_23512,N_23630);
or U24658 (N_24658,N_23515,N_19018);
xor U24659 (N_24659,N_21682,N_21155);
nand U24660 (N_24660,N_21551,N_18523);
xnor U24661 (N_24661,N_21292,N_23581);
nand U24662 (N_24662,N_18636,N_21496);
nor U24663 (N_24663,N_21941,N_19901);
and U24664 (N_24664,N_19656,N_23554);
xor U24665 (N_24665,N_19458,N_22501);
and U24666 (N_24666,N_18784,N_18147);
or U24667 (N_24667,N_19363,N_19331);
nor U24668 (N_24668,N_19176,N_22952);
nand U24669 (N_24669,N_18087,N_19647);
nor U24670 (N_24670,N_19440,N_21317);
and U24671 (N_24671,N_21391,N_23866);
or U24672 (N_24672,N_22123,N_19392);
nor U24673 (N_24673,N_20898,N_19983);
nand U24674 (N_24674,N_23690,N_21409);
and U24675 (N_24675,N_23937,N_18407);
and U24676 (N_24676,N_20751,N_23065);
xor U24677 (N_24677,N_22709,N_20049);
or U24678 (N_24678,N_22865,N_20587);
xnor U24679 (N_24679,N_18252,N_19066);
or U24680 (N_24680,N_18414,N_23979);
or U24681 (N_24681,N_20046,N_23509);
nand U24682 (N_24682,N_22383,N_19110);
nand U24683 (N_24683,N_20702,N_23638);
or U24684 (N_24684,N_22186,N_20945);
or U24685 (N_24685,N_20001,N_22202);
nand U24686 (N_24686,N_19683,N_23349);
and U24687 (N_24687,N_20837,N_18282);
nor U24688 (N_24688,N_18022,N_18737);
xnor U24689 (N_24689,N_18312,N_21038);
or U24690 (N_24690,N_23763,N_20152);
or U24691 (N_24691,N_18304,N_18866);
xor U24692 (N_24692,N_23906,N_20227);
or U24693 (N_24693,N_18368,N_21470);
and U24694 (N_24694,N_20451,N_20615);
nor U24695 (N_24695,N_18054,N_22879);
and U24696 (N_24696,N_21271,N_19234);
or U24697 (N_24697,N_20620,N_21153);
nor U24698 (N_24698,N_18818,N_22872);
or U24699 (N_24699,N_18068,N_23603);
nand U24700 (N_24700,N_20936,N_23392);
nand U24701 (N_24701,N_21692,N_20950);
xnor U24702 (N_24702,N_23735,N_18074);
nand U24703 (N_24703,N_22384,N_20399);
or U24704 (N_24704,N_22339,N_19816);
and U24705 (N_24705,N_18402,N_21576);
xnor U24706 (N_24706,N_23494,N_20591);
nand U24707 (N_24707,N_18736,N_20708);
nand U24708 (N_24708,N_22238,N_19976);
or U24709 (N_24709,N_23893,N_23035);
and U24710 (N_24710,N_21025,N_18012);
or U24711 (N_24711,N_19010,N_19862);
or U24712 (N_24712,N_19539,N_22678);
nand U24713 (N_24713,N_18441,N_22715);
nand U24714 (N_24714,N_18331,N_19097);
or U24715 (N_24715,N_18926,N_18264);
nor U24716 (N_24716,N_18267,N_18107);
or U24717 (N_24717,N_19410,N_22812);
and U24718 (N_24718,N_19524,N_18517);
and U24719 (N_24719,N_18949,N_22940);
xor U24720 (N_24720,N_21461,N_18614);
xor U24721 (N_24721,N_23264,N_22927);
and U24722 (N_24722,N_23379,N_20551);
or U24723 (N_24723,N_22510,N_19376);
nor U24724 (N_24724,N_19791,N_22988);
nor U24725 (N_24725,N_20156,N_20586);
nand U24726 (N_24726,N_21177,N_23624);
xnor U24727 (N_24727,N_21865,N_18396);
nand U24728 (N_24728,N_19086,N_19892);
or U24729 (N_24729,N_22783,N_18530);
nand U24730 (N_24730,N_19713,N_23068);
nand U24731 (N_24731,N_23397,N_20504);
nand U24732 (N_24732,N_23875,N_18662);
or U24733 (N_24733,N_21132,N_22067);
and U24734 (N_24734,N_19965,N_22112);
and U24735 (N_24735,N_22512,N_21517);
nand U24736 (N_24736,N_23785,N_22497);
or U24737 (N_24737,N_21144,N_18514);
and U24738 (N_24738,N_20588,N_20334);
xnor U24739 (N_24739,N_22469,N_20476);
and U24740 (N_24740,N_21710,N_18802);
nand U24741 (N_24741,N_23536,N_22163);
and U24742 (N_24742,N_20698,N_19624);
or U24743 (N_24743,N_22416,N_22142);
and U24744 (N_24744,N_20920,N_22899);
nor U24745 (N_24745,N_20428,N_19049);
xor U24746 (N_24746,N_21531,N_18977);
xor U24747 (N_24747,N_18521,N_18397);
nor U24748 (N_24748,N_21384,N_22917);
nand U24749 (N_24749,N_19634,N_19955);
or U24750 (N_24750,N_20801,N_20721);
xnor U24751 (N_24751,N_19810,N_21039);
or U24752 (N_24752,N_18678,N_23495);
xor U24753 (N_24753,N_19945,N_20557);
nor U24754 (N_24754,N_18162,N_23890);
or U24755 (N_24755,N_21866,N_21130);
and U24756 (N_24756,N_22273,N_20695);
and U24757 (N_24757,N_18399,N_19764);
xnor U24758 (N_24758,N_23483,N_23410);
nor U24759 (N_24759,N_23508,N_19633);
and U24760 (N_24760,N_18734,N_19272);
and U24761 (N_24761,N_18589,N_20909);
nand U24762 (N_24762,N_23448,N_21113);
and U24763 (N_24763,N_21820,N_21624);
xor U24764 (N_24764,N_23715,N_20840);
nor U24765 (N_24765,N_23107,N_20225);
or U24766 (N_24766,N_20022,N_19918);
xnor U24767 (N_24767,N_20232,N_23366);
or U24768 (N_24768,N_18208,N_19327);
or U24769 (N_24769,N_18842,N_20977);
xnor U24770 (N_24770,N_20191,N_19621);
and U24771 (N_24771,N_22420,N_18363);
nor U24772 (N_24772,N_20515,N_21903);
and U24773 (N_24773,N_21778,N_21152);
nor U24774 (N_24774,N_22631,N_23502);
xnor U24775 (N_24775,N_21165,N_22058);
or U24776 (N_24776,N_21233,N_21683);
nand U24777 (N_24777,N_21112,N_23713);
and U24778 (N_24778,N_22005,N_19773);
nor U24779 (N_24779,N_21831,N_19710);
nor U24780 (N_24780,N_20418,N_18250);
and U24781 (N_24781,N_22682,N_23204);
or U24782 (N_24782,N_21076,N_20939);
nor U24783 (N_24783,N_19300,N_23444);
nor U24784 (N_24784,N_18844,N_18281);
or U24785 (N_24785,N_22808,N_21647);
or U24786 (N_24786,N_22981,N_21524);
xnor U24787 (N_24787,N_20808,N_18700);
nand U24788 (N_24788,N_18351,N_21891);
xnor U24789 (N_24789,N_18673,N_23469);
nor U24790 (N_24790,N_19992,N_23574);
and U24791 (N_24791,N_19126,N_22408);
nor U24792 (N_24792,N_21110,N_23712);
or U24793 (N_24793,N_23249,N_23121);
nor U24794 (N_24794,N_23069,N_18193);
xnor U24795 (N_24795,N_22559,N_23547);
nand U24796 (N_24796,N_23953,N_21469);
nor U24797 (N_24797,N_21652,N_19443);
or U24798 (N_24798,N_19391,N_22357);
or U24799 (N_24799,N_21200,N_22158);
xor U24800 (N_24800,N_20181,N_19123);
nor U24801 (N_24801,N_18513,N_22785);
xor U24802 (N_24802,N_18714,N_19738);
or U24803 (N_24803,N_20366,N_18624);
nand U24804 (N_24804,N_20002,N_21649);
or U24805 (N_24805,N_22257,N_23271);
and U24806 (N_24806,N_18537,N_23973);
and U24807 (N_24807,N_22334,N_22502);
nand U24808 (N_24808,N_23525,N_21793);
xor U24809 (N_24809,N_20529,N_23546);
or U24810 (N_24810,N_20754,N_21385);
xor U24811 (N_24811,N_19948,N_18760);
xor U24812 (N_24812,N_23309,N_21003);
nor U24813 (N_24813,N_23296,N_21699);
and U24814 (N_24814,N_21590,N_19469);
and U24815 (N_24815,N_21834,N_21406);
xor U24816 (N_24816,N_22613,N_22685);
or U24817 (N_24817,N_18808,N_18225);
and U24818 (N_24818,N_18310,N_20264);
or U24819 (N_24819,N_21288,N_22436);
and U24820 (N_24820,N_19175,N_23314);
nand U24821 (N_24821,N_22191,N_19932);
nand U24822 (N_24822,N_18135,N_21990);
xor U24823 (N_24823,N_19115,N_20521);
nand U24824 (N_24824,N_18392,N_21031);
or U24825 (N_24825,N_20846,N_19691);
nand U24826 (N_24826,N_21924,N_20329);
or U24827 (N_24827,N_23355,N_22710);
or U24828 (N_24828,N_19554,N_20816);
and U24829 (N_24829,N_21184,N_18727);
or U24830 (N_24830,N_18670,N_21253);
and U24831 (N_24831,N_20901,N_22766);
xnor U24832 (N_24832,N_20989,N_21828);
xnor U24833 (N_24833,N_20218,N_19244);
or U24834 (N_24834,N_19623,N_22377);
or U24835 (N_24835,N_20349,N_18692);
nand U24836 (N_24836,N_22042,N_22621);
or U24837 (N_24837,N_18854,N_19026);
nand U24838 (N_24838,N_22326,N_21977);
nand U24839 (N_24839,N_20492,N_23535);
and U24840 (N_24840,N_18400,N_19507);
nor U24841 (N_24841,N_18723,N_20759);
or U24842 (N_24842,N_21529,N_23593);
or U24843 (N_24843,N_21872,N_18338);
or U24844 (N_24844,N_22364,N_20396);
nor U24845 (N_24845,N_19411,N_18899);
nor U24846 (N_24846,N_23316,N_22409);
xnor U24847 (N_24847,N_18393,N_23384);
xor U24848 (N_24848,N_21337,N_21744);
and U24849 (N_24849,N_18341,N_19956);
xor U24850 (N_24850,N_18473,N_23622);
or U24851 (N_24851,N_20112,N_22386);
and U24852 (N_24852,N_21009,N_20015);
xor U24853 (N_24853,N_19350,N_19533);
nor U24854 (N_24854,N_20981,N_18053);
and U24855 (N_24855,N_21519,N_18319);
or U24856 (N_24856,N_22632,N_21462);
or U24857 (N_24857,N_19853,N_18828);
nor U24858 (N_24858,N_21279,N_22035);
nor U24859 (N_24859,N_20889,N_21525);
or U24860 (N_24860,N_22064,N_18959);
nand U24861 (N_24861,N_23604,N_20969);
nand U24862 (N_24862,N_23849,N_18148);
or U24863 (N_24863,N_21294,N_23609);
or U24864 (N_24864,N_20867,N_20985);
nor U24865 (N_24865,N_23230,N_21185);
and U24866 (N_24866,N_19506,N_20217);
nor U24867 (N_24867,N_21212,N_20844);
nor U24868 (N_24868,N_19256,N_18480);
xnor U24869 (N_24869,N_18099,N_22004);
xor U24870 (N_24870,N_18686,N_18540);
xor U24871 (N_24871,N_19888,N_21446);
and U24872 (N_24872,N_21645,N_23651);
and U24873 (N_24873,N_23423,N_21411);
or U24874 (N_24874,N_18545,N_18487);
nor U24875 (N_24875,N_23967,N_22183);
or U24876 (N_24876,N_19706,N_20235);
nor U24877 (N_24877,N_20173,N_21228);
xnor U24878 (N_24878,N_22546,N_18145);
xnor U24879 (N_24879,N_19959,N_19645);
or U24880 (N_24880,N_19481,N_20377);
nor U24881 (N_24881,N_19320,N_22237);
nand U24882 (N_24882,N_21383,N_19157);
and U24883 (N_24883,N_23720,N_21273);
xor U24884 (N_24884,N_23804,N_18869);
and U24885 (N_24885,N_18972,N_23914);
and U24886 (N_24886,N_20443,N_22418);
and U24887 (N_24887,N_20701,N_19537);
and U24888 (N_24888,N_21715,N_19346);
xnor U24889 (N_24889,N_21787,N_20155);
and U24890 (N_24890,N_20150,N_22558);
xor U24891 (N_24891,N_23046,N_19622);
or U24892 (N_24892,N_21215,N_18631);
xor U24893 (N_24893,N_21812,N_18565);
and U24894 (N_24894,N_20370,N_21248);
nor U24895 (N_24895,N_23369,N_19952);
nor U24896 (N_24896,N_22208,N_23187);
nand U24897 (N_24897,N_21868,N_21192);
xnor U24898 (N_24898,N_22933,N_23434);
nand U24899 (N_24899,N_22269,N_23637);
or U24900 (N_24900,N_18309,N_18781);
xnor U24901 (N_24901,N_22426,N_21769);
nor U24902 (N_24902,N_19798,N_22972);
xor U24903 (N_24903,N_22537,N_20414);
nor U24904 (N_24904,N_18562,N_22906);
nor U24905 (N_24905,N_23313,N_20480);
nand U24906 (N_24906,N_21560,N_22674);
and U24907 (N_24907,N_18038,N_21023);
and U24908 (N_24908,N_21592,N_23784);
nor U24909 (N_24909,N_23588,N_23294);
or U24910 (N_24910,N_21362,N_21805);
or U24911 (N_24911,N_18069,N_19631);
and U24912 (N_24912,N_23252,N_18139);
nor U24913 (N_24913,N_18429,N_18641);
nand U24914 (N_24914,N_22451,N_20857);
or U24915 (N_24915,N_20244,N_18794);
or U24916 (N_24916,N_19919,N_20929);
and U24917 (N_24917,N_23734,N_20086);
nand U24918 (N_24918,N_19017,N_21050);
and U24919 (N_24919,N_20522,N_18160);
xor U24920 (N_24920,N_20454,N_23073);
xnor U24921 (N_24921,N_20826,N_21651);
and U24922 (N_24922,N_19290,N_20713);
and U24923 (N_24923,N_19674,N_23273);
or U24924 (N_24924,N_18950,N_22247);
nor U24925 (N_24925,N_22243,N_23826);
nor U24926 (N_24926,N_22098,N_20687);
xor U24927 (N_24927,N_18923,N_20863);
and U24928 (N_24928,N_22025,N_21908);
nor U24929 (N_24929,N_23362,N_19137);
nor U24930 (N_24930,N_18025,N_19322);
or U24931 (N_24931,N_21762,N_22600);
and U24932 (N_24932,N_19653,N_23898);
or U24933 (N_24933,N_19516,N_20079);
nand U24934 (N_24934,N_18167,N_19846);
and U24935 (N_24935,N_22769,N_21407);
nor U24936 (N_24936,N_18405,N_22268);
nor U24937 (N_24937,N_20076,N_18531);
xor U24938 (N_24938,N_23120,N_23756);
nand U24939 (N_24939,N_20527,N_22284);
nor U24940 (N_24940,N_18470,N_21108);
and U24941 (N_24941,N_18920,N_18867);
nor U24942 (N_24942,N_21665,N_22725);
nor U24943 (N_24943,N_18774,N_19023);
xnor U24944 (N_24944,N_20371,N_22814);
and U24945 (N_24945,N_18333,N_19699);
xor U24946 (N_24946,N_18080,N_19534);
nor U24947 (N_24947,N_20506,N_21239);
nor U24948 (N_24948,N_20249,N_23745);
nor U24949 (N_24949,N_23894,N_19697);
and U24950 (N_24950,N_20212,N_21505);
nand U24951 (N_24951,N_23009,N_20158);
or U24952 (N_24952,N_22322,N_19970);
and U24953 (N_24953,N_18048,N_22714);
nand U24954 (N_24954,N_23928,N_23684);
nand U24955 (N_24955,N_18595,N_19615);
or U24956 (N_24956,N_20198,N_23087);
nand U24957 (N_24957,N_18078,N_23506);
and U24958 (N_24958,N_23432,N_19310);
or U24959 (N_24959,N_19241,N_23811);
nor U24960 (N_24960,N_22150,N_18507);
xor U24961 (N_24961,N_20693,N_22173);
xnor U24962 (N_24962,N_22841,N_20052);
nor U24963 (N_24963,N_22973,N_21029);
nor U24964 (N_24964,N_20023,N_21541);
nor U24965 (N_24965,N_21901,N_19758);
and U24966 (N_24966,N_22127,N_21542);
or U24967 (N_24967,N_19984,N_23004);
xor U24968 (N_24968,N_22011,N_20166);
xnor U24969 (N_24969,N_20335,N_23545);
nand U24970 (N_24970,N_23996,N_20827);
or U24971 (N_24971,N_23839,N_19861);
nand U24972 (N_24972,N_19609,N_23272);
nand U24973 (N_24973,N_20231,N_19399);
xor U24974 (N_24974,N_20778,N_18927);
nor U24975 (N_24975,N_19103,N_21013);
nor U24976 (N_24976,N_19487,N_18255);
nand U24977 (N_24977,N_20140,N_23641);
and U24978 (N_24978,N_20718,N_22231);
or U24979 (N_24979,N_21942,N_20542);
nor U24980 (N_24980,N_21912,N_23295);
or U24981 (N_24981,N_19160,N_18105);
xnor U24982 (N_24982,N_20890,N_18224);
nor U24983 (N_24983,N_19761,N_18464);
nor U24984 (N_24984,N_23869,N_22286);
and U24985 (N_24985,N_19281,N_22277);
nor U24986 (N_24986,N_19786,N_19882);
nand U24987 (N_24987,N_20354,N_19341);
and U24988 (N_24988,N_22816,N_20530);
nand U24989 (N_24989,N_20105,N_18045);
and U24990 (N_24990,N_19709,N_18750);
nand U24991 (N_24991,N_22266,N_22433);
xnor U24992 (N_24992,N_21729,N_20628);
nor U24993 (N_24993,N_22576,N_18663);
nor U24994 (N_24994,N_18051,N_18588);
nand U24995 (N_24995,N_23059,N_22126);
nor U24996 (N_24996,N_23421,N_22223);
nand U24997 (N_24997,N_23363,N_18316);
or U24998 (N_24998,N_21230,N_19449);
nor U24999 (N_24999,N_20066,N_19197);
nand U25000 (N_25000,N_18063,N_21236);
nor U25001 (N_25001,N_18832,N_23897);
xor U25002 (N_25002,N_23931,N_22491);
xnor U25003 (N_25003,N_18364,N_20455);
nand U25004 (N_25004,N_20069,N_23474);
and U25005 (N_25005,N_19342,N_23873);
nand U25006 (N_25006,N_19077,N_23226);
or U25007 (N_25007,N_22634,N_18783);
nand U25008 (N_25008,N_18796,N_22995);
xor U25009 (N_25009,N_20828,N_18868);
and U25010 (N_25010,N_20852,N_21457);
xnor U25011 (N_25011,N_18841,N_22008);
nand U25012 (N_25012,N_21706,N_22049);
or U25013 (N_25013,N_23132,N_22974);
or U25014 (N_25014,N_21881,N_18735);
xnor U25015 (N_25015,N_18956,N_21324);
nor U25016 (N_25016,N_19374,N_19425);
xor U25017 (N_25017,N_22313,N_21074);
nand U25018 (N_25018,N_23376,N_21681);
nand U25019 (N_25019,N_22195,N_21939);
or U25020 (N_25020,N_22315,N_18770);
or U25021 (N_25021,N_21911,N_22110);
nor U25022 (N_25022,N_22957,N_22645);
nand U25023 (N_25023,N_19274,N_19192);
nand U25024 (N_25024,N_22478,N_18902);
and U25025 (N_25025,N_22069,N_18650);
or U25026 (N_25026,N_19519,N_20536);
nand U25027 (N_25027,N_20940,N_21958);
xnor U25028 (N_25028,N_21503,N_20507);
nand U25029 (N_25029,N_19140,N_21252);
or U25030 (N_25030,N_20120,N_22084);
nor U25031 (N_25031,N_18551,N_19328);
nor U25032 (N_25032,N_21088,N_20058);
nand U25033 (N_25033,N_19675,N_23929);
nor U25034 (N_25034,N_20466,N_19043);
or U25035 (N_25035,N_18124,N_22092);
nor U25036 (N_25036,N_22666,N_22505);
nand U25037 (N_25037,N_23719,N_23023);
and U25038 (N_25038,N_19245,N_22130);
nand U25039 (N_25039,N_23135,N_20309);
xnor U25040 (N_25040,N_22177,N_22536);
xnor U25041 (N_25041,N_23097,N_20385);
nor U25042 (N_25042,N_20988,N_19085);
and U25043 (N_25043,N_23950,N_21575);
and U25044 (N_25044,N_20992,N_22616);
nand U25045 (N_25045,N_21905,N_23548);
nand U25046 (N_25046,N_19815,N_19426);
and U25047 (N_25047,N_18705,N_20470);
and U25048 (N_25048,N_18314,N_19672);
xor U25049 (N_25049,N_20673,N_19365);
nand U25050 (N_25050,N_19511,N_18894);
nand U25051 (N_25051,N_18940,N_18064);
or U25052 (N_25052,N_21666,N_19476);
nand U25053 (N_25053,N_20074,N_20921);
and U25054 (N_25054,N_20948,N_23833);
nand U25055 (N_25055,N_21174,N_22176);
nand U25056 (N_25056,N_20930,N_18449);
nor U25057 (N_25057,N_20907,N_19313);
and U25058 (N_25058,N_23398,N_22345);
nor U25059 (N_25059,N_19323,N_22909);
nand U25060 (N_25060,N_18685,N_18988);
nor U25061 (N_25061,N_20845,N_20045);
or U25062 (N_25062,N_23968,N_22063);
or U25063 (N_25063,N_18814,N_23786);
or U25064 (N_25064,N_22583,N_18488);
nand U25065 (N_25065,N_18273,N_20660);
nor U25066 (N_25066,N_22180,N_22998);
nand U25067 (N_25067,N_18610,N_19676);
and U25068 (N_25068,N_21109,N_23173);
xnor U25069 (N_25069,N_21436,N_18827);
nand U25070 (N_25070,N_18568,N_18509);
nand U25071 (N_25071,N_20478,N_18761);
and U25072 (N_25072,N_20995,N_18448);
nand U25073 (N_25073,N_18938,N_21332);
nor U25074 (N_25074,N_22303,N_21770);
and U25075 (N_25075,N_19574,N_22473);
nor U25076 (N_25076,N_21860,N_23165);
nand U25077 (N_25077,N_18511,N_18157);
nand U25078 (N_25078,N_21932,N_22477);
xor U25079 (N_25079,N_21583,N_22525);
xor U25080 (N_25080,N_21599,N_18498);
xor U25081 (N_25081,N_23386,N_22637);
nand U25082 (N_25082,N_18897,N_21935);
or U25083 (N_25083,N_20036,N_19800);
xnor U25084 (N_25084,N_19294,N_19994);
nor U25085 (N_25085,N_19384,N_23387);
or U25086 (N_25086,N_22684,N_18017);
nor U25087 (N_25087,N_19332,N_18367);
nand U25088 (N_25088,N_23032,N_22579);
or U25089 (N_25089,N_18456,N_20903);
or U25090 (N_25090,N_19803,N_21376);
or U25091 (N_25091,N_20009,N_19985);
xnor U25092 (N_25092,N_21987,N_21305);
nor U25093 (N_25093,N_23900,N_23566);
nor U25094 (N_25094,N_19759,N_20135);
nand U25095 (N_25095,N_18376,N_18857);
or U25096 (N_25096,N_21458,N_19584);
nand U25097 (N_25097,N_19828,N_18460);
nor U25098 (N_25098,N_23238,N_19573);
and U25099 (N_25099,N_19665,N_19191);
nand U25100 (N_25100,N_23206,N_23595);
xnor U25101 (N_25101,N_18375,N_21286);
and U25102 (N_25102,N_21423,N_22133);
xor U25103 (N_25103,N_21450,N_20781);
nor U25104 (N_25104,N_22338,N_23406);
and U25105 (N_25105,N_21558,N_18419);
nor U25106 (N_25106,N_19702,N_18266);
or U25107 (N_25107,N_19151,N_22839);
and U25108 (N_25108,N_23300,N_20063);
and U25109 (N_25109,N_21237,N_22533);
or U25110 (N_25110,N_19246,N_23511);
nand U25111 (N_25111,N_18081,N_20878);
xnor U25112 (N_25112,N_19670,N_18541);
or U25113 (N_25113,N_19262,N_21206);
nor U25114 (N_25114,N_22843,N_23645);
or U25115 (N_25115,N_19479,N_20576);
nor U25116 (N_25116,N_19243,N_23008);
or U25117 (N_25117,N_20487,N_19421);
and U25118 (N_25118,N_19662,N_22830);
or U25119 (N_25119,N_20994,N_21523);
nor U25120 (N_25120,N_21062,N_23413);
nand U25121 (N_25121,N_18445,N_21479);
or U25122 (N_25122,N_20641,N_19441);
and U25123 (N_25123,N_20409,N_20786);
nand U25124 (N_25124,N_21882,N_23631);
xor U25125 (N_25125,N_20999,N_20509);
or U25126 (N_25126,N_18759,N_22667);
or U25127 (N_25127,N_23427,N_23810);
xor U25128 (N_25128,N_22569,N_21443);
and U25129 (N_25129,N_19034,N_20067);
nor U25130 (N_25130,N_18209,N_23861);
and U25131 (N_25131,N_22607,N_20392);
xor U25132 (N_25132,N_23317,N_19439);
nor U25133 (N_25133,N_23458,N_21350);
nand U25134 (N_25134,N_23851,N_22017);
and U25135 (N_25135,N_22487,N_20338);
nand U25136 (N_25136,N_22937,N_23823);
nand U25137 (N_25137,N_19655,N_21680);
xor U25138 (N_25138,N_23706,N_21262);
nand U25139 (N_25139,N_21117,N_21956);
nor U25140 (N_25140,N_23606,N_21372);
or U25141 (N_25141,N_23551,N_22001);
or U25142 (N_25142,N_19909,N_23454);
xor U25143 (N_25143,N_21363,N_20207);
or U25144 (N_25144,N_21573,N_18953);
or U25145 (N_25145,N_19390,N_22532);
xnor U25146 (N_25146,N_22038,N_21131);
xor U25147 (N_25147,N_18205,N_22571);
or U25148 (N_25148,N_21274,N_23268);
nand U25149 (N_25149,N_22400,N_21049);
and U25150 (N_25150,N_20908,N_19680);
nand U25151 (N_25151,N_19667,N_21118);
xnor U25152 (N_25152,N_18979,N_23328);
and U25153 (N_25153,N_20575,N_22856);
and U25154 (N_25154,N_20347,N_21814);
nor U25155 (N_25155,N_20951,N_20511);
xor U25156 (N_25156,N_18251,N_22404);
nor U25157 (N_25157,N_23969,N_21310);
nand U25158 (N_25158,N_20514,N_20911);
xnor U25159 (N_25159,N_21640,N_19865);
and U25160 (N_25160,N_23597,N_21055);
nor U25161 (N_25161,N_22787,N_20375);
nor U25162 (N_25162,N_18353,N_22235);
or U25163 (N_25163,N_20743,N_20734);
nand U25164 (N_25164,N_23891,N_21162);
or U25165 (N_25165,N_21774,N_22267);
and U25166 (N_25166,N_20025,N_18896);
nor U25167 (N_25167,N_20416,N_21570);
or U25168 (N_25168,N_18370,N_18438);
xor U25169 (N_25169,N_18744,N_22795);
nand U25170 (N_25170,N_23420,N_22651);
nand U25171 (N_25171,N_23537,N_18122);
or U25172 (N_25172,N_20770,N_18008);
nor U25173 (N_25173,N_18158,N_21361);
xnor U25174 (N_25174,N_19700,N_19353);
or U25175 (N_25175,N_21613,N_18125);
xor U25176 (N_25176,N_22380,N_21946);
nor U25177 (N_25177,N_18939,N_21208);
or U25178 (N_25178,N_23758,N_18230);
and U25179 (N_25179,N_23753,N_19794);
xor U25180 (N_25180,N_21082,N_23409);
and U25181 (N_25181,N_20143,N_22254);
nand U25182 (N_25182,N_21138,N_23211);
xnor U25183 (N_25183,N_20029,N_20154);
xnor U25184 (N_25184,N_22876,N_18121);
xnor U25185 (N_25185,N_19060,N_22702);
xnor U25186 (N_25186,N_23951,N_20957);
nor U25187 (N_25187,N_19722,N_22971);
nor U25188 (N_25188,N_18362,N_21285);
or U25189 (N_25189,N_22242,N_20057);
nor U25190 (N_25190,N_19982,N_19419);
nand U25191 (N_25191,N_22285,N_18611);
nor U25192 (N_25192,N_20609,N_18960);
and U25193 (N_25193,N_22051,N_20883);
and U25194 (N_25194,N_22619,N_22519);
xnor U25195 (N_25195,N_22969,N_21913);
or U25196 (N_25196,N_19231,N_22304);
or U25197 (N_25197,N_22424,N_19490);
xor U25198 (N_25198,N_22746,N_18150);
or U25199 (N_25199,N_18272,N_20008);
or U25200 (N_25200,N_19632,N_20580);
nand U25201 (N_25201,N_18112,N_22037);
xnor U25202 (N_25202,N_20384,N_22316);
nor U25203 (N_25203,N_21464,N_23263);
nand U25204 (N_25204,N_23175,N_22405);
xnor U25205 (N_25205,N_20426,N_22106);
xor U25206 (N_25206,N_22143,N_20502);
nor U25207 (N_25207,N_18476,N_21091);
nand U25208 (N_25208,N_21115,N_22138);
or U25209 (N_25209,N_23341,N_20872);
nand U25210 (N_25210,N_20865,N_19728);
xor U25211 (N_25211,N_23658,N_23730);
nand U25212 (N_25212,N_18970,N_19986);
or U25213 (N_25213,N_22145,N_22393);
nor U25214 (N_25214,N_18559,N_18757);
and U25215 (N_25215,N_22833,N_18183);
nor U25216 (N_25216,N_19369,N_18679);
xor U25217 (N_25217,N_18691,N_18245);
nand U25218 (N_25218,N_20355,N_19750);
nor U25219 (N_25219,N_21937,N_23885);
or U25220 (N_25220,N_18567,N_23236);
and U25221 (N_25221,N_21104,N_23333);
nand U25222 (N_25222,N_23318,N_22196);
nand U25223 (N_25223,N_19271,N_18475);
nand U25224 (N_25224,N_23172,N_21947);
and U25225 (N_25225,N_21161,N_18524);
nand U25226 (N_25226,N_19666,N_19132);
and U25227 (N_25227,N_23468,N_18644);
nand U25228 (N_25228,N_20468,N_23026);
nor U25229 (N_25229,N_18677,N_19308);
xnor U25230 (N_25230,N_19032,N_21585);
and U25231 (N_25231,N_18912,N_21857);
and U25232 (N_25232,N_22467,N_21980);
nand U25233 (N_25233,N_18303,N_21593);
and U25234 (N_25234,N_23189,N_21716);
or U25235 (N_25235,N_19378,N_20255);
nand U25236 (N_25236,N_23698,N_22356);
and U25237 (N_25237,N_21094,N_18625);
xnor U25238 (N_25238,N_23364,N_18103);
xnor U25239 (N_25239,N_21695,N_23130);
nor U25240 (N_25240,N_22029,N_23103);
and U25241 (N_25241,N_19280,N_19450);
nand U25242 (N_25242,N_22099,N_18443);
and U25243 (N_25243,N_23401,N_23460);
and U25244 (N_25244,N_23043,N_19355);
nor U25245 (N_25245,N_23353,N_18999);
nand U25246 (N_25246,N_22472,N_18554);
nand U25247 (N_25247,N_20442,N_19890);
nor U25248 (N_25248,N_19513,N_18722);
and U25249 (N_25249,N_21053,N_22498);
nor U25250 (N_25250,N_19792,N_19229);
or U25251 (N_25251,N_19494,N_20240);
nand U25252 (N_25252,N_21945,N_20727);
and U25253 (N_25253,N_22441,N_18930);
xnor U25254 (N_25254,N_21321,N_23808);
nor U25255 (N_25255,N_21642,N_23019);
xor U25256 (N_25256,N_21095,N_19442);
xnor U25257 (N_25257,N_19719,N_20438);
xnor U25258 (N_25258,N_23402,N_22402);
nor U25259 (N_25259,N_21657,N_22018);
xnor U25260 (N_25260,N_22915,N_22082);
xnor U25261 (N_25261,N_23456,N_22371);
nor U25262 (N_25262,N_20788,N_22499);
or U25263 (N_25263,N_19154,N_22435);
nand U25264 (N_25264,N_23711,N_22128);
or U25265 (N_25265,N_19340,N_19635);
or U25266 (N_25266,N_22694,N_18451);
or U25267 (N_25267,N_18260,N_23222);
or U25268 (N_25268,N_21471,N_18491);
xnor U25269 (N_25269,N_21594,N_21494);
xnor U25270 (N_25270,N_18289,N_20216);
nor U25271 (N_25271,N_19381,N_19669);
or U25272 (N_25272,N_20125,N_18661);
nand U25273 (N_25273,N_23375,N_18330);
and U25274 (N_25274,N_20669,N_20526);
or U25275 (N_25275,N_22798,N_20953);
nor U25276 (N_25276,N_19088,N_21209);
or U25277 (N_25277,N_18877,N_21349);
nand U25278 (N_25278,N_19852,N_21482);
and U25279 (N_25279,N_19493,N_18703);
and U25280 (N_25280,N_21405,N_22139);
nand U25281 (N_25281,N_21633,N_22859);
and U25282 (N_25282,N_20290,N_20256);
or U25283 (N_25283,N_22503,N_18825);
or U25284 (N_25284,N_23195,N_20777);
or U25285 (N_25285,N_20325,N_20971);
xnor U25286 (N_25286,N_21855,N_22575);
xor U25287 (N_25287,N_22297,N_22060);
or U25288 (N_25288,N_23762,N_23052);
and U25289 (N_25289,N_22012,N_20774);
xor U25290 (N_25290,N_20491,N_22976);
or U25291 (N_25291,N_20005,N_20692);
nand U25292 (N_25292,N_23381,N_18185);
or U25293 (N_25293,N_21511,N_20077);
nor U25294 (N_25294,N_18816,N_20211);
nor U25295 (N_25295,N_20558,N_19592);
nor U25296 (N_25296,N_21070,N_19755);
nor U25297 (N_25297,N_23946,N_23461);
nand U25298 (N_25298,N_20703,N_23776);
and U25299 (N_25299,N_22763,N_20924);
nor U25300 (N_25300,N_21435,N_18154);
or U25301 (N_25301,N_23710,N_20189);
nand U25302 (N_25302,N_23408,N_18357);
nor U25303 (N_25303,N_22837,N_22310);
and U25304 (N_25304,N_19040,N_22641);
xor U25305 (N_25305,N_21364,N_20246);
and U25306 (N_25306,N_18430,N_19896);
nand U25307 (N_25307,N_21068,N_19317);
nor U25308 (N_25308,N_20811,N_19620);
xor U25309 (N_25309,N_22854,N_23424);
xor U25310 (N_25310,N_18322,N_21621);
nand U25311 (N_25311,N_22595,N_19560);
and U25312 (N_25312,N_20228,N_19193);
nor U25313 (N_25313,N_19387,N_23292);
nor U25314 (N_25314,N_19412,N_19462);
nand U25315 (N_25315,N_21455,N_19169);
or U25316 (N_25316,N_18874,N_19074);
or U25317 (N_25317,N_18681,N_19498);
nor U25318 (N_25318,N_19383,N_18075);
nand U25319 (N_25319,N_18980,N_21895);
nand U25320 (N_25320,N_21226,N_20071);
or U25321 (N_25321,N_19102,N_23248);
xor U25322 (N_25322,N_22028,N_20406);
nand U25323 (N_25323,N_19811,N_21234);
nand U25324 (N_25324,N_22031,N_23255);
and U25325 (N_25325,N_18120,N_22283);
and U25326 (N_25326,N_22299,N_19107);
nor U25327 (N_25327,N_19860,N_18500);
nand U25328 (N_25328,N_20564,N_23213);
and U25329 (N_25329,N_22187,N_20559);
nor U25330 (N_25330,N_23828,N_21894);
xor U25331 (N_25331,N_20720,N_18287);
or U25332 (N_25332,N_21373,N_21022);
nor U25333 (N_25333,N_23747,N_18690);
nor U25334 (N_25334,N_19768,N_22538);
or U25335 (N_25335,N_21839,N_23462);
or U25336 (N_25336,N_19259,N_21801);
xor U25337 (N_25337,N_22294,N_22440);
nor U25338 (N_25338,N_20516,N_18073);
nor U25339 (N_25339,N_19928,N_23882);
xnor U25340 (N_25340,N_19687,N_18726);
or U25341 (N_25341,N_22910,N_21568);
nand U25342 (N_25342,N_21742,N_19059);
xnor U25343 (N_25343,N_23764,N_23276);
and U25344 (N_25344,N_19471,N_18294);
or U25345 (N_25345,N_23470,N_19962);
nand U25346 (N_25346,N_22585,N_21660);
and U25347 (N_25347,N_23403,N_22762);
nor U25348 (N_25348,N_19045,N_21147);
xor U25349 (N_25349,N_18581,N_23687);
xnor U25350 (N_25350,N_21024,N_20707);
xnor U25351 (N_25351,N_20722,N_23334);
or U25352 (N_25352,N_19319,N_20281);
and U25353 (N_25353,N_23119,N_21741);
or U25354 (N_25354,N_23006,N_19960);
or U25355 (N_25355,N_23778,N_22696);
nand U25356 (N_25356,N_19122,N_19582);
and U25357 (N_25357,N_19195,N_22065);
nor U25358 (N_25358,N_20821,N_19424);
nor U25359 (N_25359,N_22347,N_19818);
or U25360 (N_25360,N_19558,N_19777);
nor U25361 (N_25361,N_19025,N_19179);
nor U25362 (N_25362,N_21105,N_19291);
nand U25363 (N_25363,N_22193,N_21546);
nand U25364 (N_25364,N_19951,N_23227);
and U25365 (N_25365,N_18501,N_21354);
nor U25366 (N_25366,N_22669,N_21697);
xnor U25367 (N_25367,N_21869,N_19485);
and U25368 (N_25368,N_18041,N_21921);
xnor U25369 (N_25369,N_22251,N_22587);
and U25370 (N_25370,N_21799,N_18918);
xor U25371 (N_25371,N_23899,N_20195);
and U25372 (N_25372,N_19575,N_21342);
and U25373 (N_25373,N_18582,N_22707);
nand U25374 (N_25374,N_21485,N_23768);
nand U25375 (N_25375,N_22119,N_18242);
nand U25376 (N_25376,N_23257,N_23064);
or U25377 (N_25377,N_19987,N_20251);
nand U25378 (N_25378,N_18665,N_21562);
or U25379 (N_25379,N_23457,N_20894);
or U25380 (N_25380,N_23796,N_23058);
or U25381 (N_25381,N_22239,N_20608);
and U25382 (N_25382,N_20952,N_19600);
nand U25383 (N_25383,N_20407,N_19577);
or U25384 (N_25384,N_21871,N_22560);
or U25385 (N_25385,N_18454,N_19288);
or U25386 (N_25386,N_20665,N_21698);
nand U25387 (N_25387,N_18829,N_21260);
xnor U25388 (N_25388,N_19284,N_20807);
nand U25389 (N_25389,N_20928,N_22156);
and U25390 (N_25390,N_20544,N_21504);
nor U25391 (N_25391,N_22336,N_23418);
or U25392 (N_25392,N_19867,N_23220);
and U25393 (N_25393,N_18900,N_20160);
nand U25394 (N_25394,N_22964,N_23939);
xnor U25395 (N_25395,N_18850,N_18401);
xor U25396 (N_25396,N_19854,N_19765);
xor U25397 (N_25397,N_21481,N_23633);
and U25398 (N_25398,N_20310,N_18797);
and U25399 (N_25399,N_23047,N_20818);
nor U25400 (N_25400,N_19268,N_20425);
or U25401 (N_25401,N_19514,N_19922);
nand U25402 (N_25402,N_22312,N_18194);
and U25403 (N_25403,N_18049,N_22047);
nor U25404 (N_25404,N_21930,N_19171);
nor U25405 (N_25405,N_19431,N_21122);
nand U25406 (N_25406,N_20900,N_20750);
nand U25407 (N_25407,N_20167,N_20966);
xnor U25408 (N_25408,N_20885,N_19520);
xor U25409 (N_25409,N_22802,N_19131);
nor U25410 (N_25410,N_20913,N_23428);
and U25411 (N_25411,N_18108,N_18746);
nor U25412 (N_25412,N_21674,N_20762);
nor U25413 (N_25413,N_20490,N_19295);
nand U25414 (N_25414,N_20876,N_21845);
and U25415 (N_25415,N_18751,N_19452);
xor U25416 (N_25416,N_19958,N_22896);
nand U25417 (N_25417,N_18793,N_19237);
or U25418 (N_25418,N_23577,N_23072);
nand U25419 (N_25419,N_18884,N_20017);
nand U25420 (N_25420,N_18674,N_20624);
or U25421 (N_25421,N_18329,N_20634);
nor U25422 (N_25422,N_18811,N_20738);
nand U25423 (N_25423,N_21460,N_19046);
and U25424 (N_25424,N_18709,N_18339);
nor U25425 (N_25425,N_18742,N_22370);
or U25426 (N_25426,N_18550,N_21447);
and U25427 (N_25427,N_18928,N_23347);
or U25428 (N_25428,N_18598,N_23827);
and U25429 (N_25429,N_18600,N_18004);
xor U25430 (N_25430,N_18009,N_20004);
and U25431 (N_25431,N_23944,N_19766);
or U25432 (N_25432,N_20633,N_22431);
nor U25433 (N_25433,N_22087,N_21141);
xor U25434 (N_25434,N_23049,N_19943);
or U25435 (N_25435,N_21623,N_19875);
and U25436 (N_25436,N_18915,N_19447);
xnor U25437 (N_25437,N_22708,N_23112);
and U25438 (N_25438,N_22021,N_18527);
or U25439 (N_25439,N_19528,N_18366);
or U25440 (N_25440,N_21944,N_22015);
nor U25441 (N_25441,N_21688,N_22949);
and U25442 (N_25442,N_23718,N_19608);
or U25443 (N_25443,N_19145,N_23610);
or U25444 (N_25444,N_18878,N_22374);
nor U25445 (N_25445,N_19429,N_20424);
nand U25446 (N_25446,N_19337,N_23336);
xnor U25447 (N_25447,N_20330,N_20303);
and U25448 (N_25448,N_23623,N_18618);
xor U25449 (N_25449,N_18584,N_19532);
nand U25450 (N_25450,N_22657,N_20704);
nand U25451 (N_25451,N_19587,N_23166);
nor U25452 (N_25452,N_19474,N_23312);
nor U25453 (N_25453,N_22043,N_23396);
nand U25454 (N_25454,N_19578,N_23902);
xnor U25455 (N_25455,N_23840,N_22348);
xnor U25456 (N_25456,N_19357,N_20146);
nand U25457 (N_25457,N_19012,N_18275);
nor U25458 (N_25458,N_22791,N_21798);
xnor U25459 (N_25459,N_19084,N_19950);
nor U25460 (N_25460,N_18697,N_23975);
nor U25461 (N_25461,N_19312,N_20295);
xor U25462 (N_25462,N_21415,N_19731);
and U25463 (N_25463,N_21287,N_22367);
nor U25464 (N_25464,N_21549,N_18643);
and U25465 (N_25465,N_18106,N_20358);
xor U25466 (N_25466,N_23818,N_20204);
nand U25467 (N_25467,N_18532,N_19906);
xor U25468 (N_25468,N_18493,N_21319);
nor U25469 (N_25469,N_20525,N_20474);
nor U25470 (N_25470,N_23523,N_20103);
and U25471 (N_25471,N_18553,N_20642);
and U25472 (N_25472,N_18028,N_21514);
nand U25473 (N_25473,N_19590,N_19382);
or U25474 (N_25474,N_23151,N_18315);
nand U25475 (N_25475,N_21302,N_21371);
or U25476 (N_25476,N_22891,N_22935);
xnor U25477 (N_25477,N_20090,N_22296);
nor U25478 (N_25478,N_23542,N_22947);
and U25479 (N_25479,N_22379,N_18881);
and U25480 (N_25480,N_22668,N_21598);
nand U25481 (N_25481,N_18018,N_23390);
nand U25482 (N_25482,N_21600,N_18497);
xor U25483 (N_25483,N_18029,N_23478);
and U25484 (N_25484,N_23031,N_21949);
or U25485 (N_25485,N_18539,N_20666);
xor U25486 (N_25486,N_20192,N_18382);
nand U25487 (N_25487,N_21205,N_21722);
nand U25488 (N_25488,N_18861,N_19995);
or U25489 (N_25489,N_18007,N_23307);
nor U25490 (N_25490,N_20706,N_23797);
nor U25491 (N_25491,N_19606,N_18197);
or U25492 (N_25492,N_18490,N_23716);
xor U25493 (N_25493,N_18833,N_23167);
nand U25494 (N_25494,N_23030,N_22701);
or U25495 (N_25495,N_23754,N_23966);
or U25496 (N_25496,N_22439,N_22460);
or U25497 (N_25497,N_22965,N_22591);
xnor U25498 (N_25498,N_19403,N_23883);
nor U25499 (N_25499,N_18308,N_22365);
xor U25500 (N_25500,N_23582,N_23670);
xnor U25501 (N_25501,N_19475,N_23726);
nor U25502 (N_25502,N_21794,N_19070);
nand U25503 (N_25503,N_22916,N_22652);
nor U25504 (N_25504,N_23338,N_23445);
and U25505 (N_25505,N_23225,N_18424);
nand U25506 (N_25506,N_18776,N_20926);
or U25507 (N_25507,N_21064,N_23076);
or U25508 (N_25508,N_21092,N_20261);
and U25509 (N_25509,N_20960,N_23002);
xnor U25510 (N_25510,N_20109,N_20178);
and U25511 (N_25511,N_23857,N_23680);
and U25512 (N_25512,N_18427,N_22022);
and U25513 (N_25513,N_21873,N_23503);
xnor U25514 (N_25514,N_20973,N_18863);
nor U25515 (N_25515,N_23750,N_21497);
and U25516 (N_25516,N_22580,N_23777);
or U25517 (N_25517,N_22504,N_18729);
nand U25518 (N_25518,N_23160,N_20405);
and U25519 (N_25519,N_18423,N_22246);
nand U25520 (N_25520,N_22993,N_20382);
and U25521 (N_25521,N_19725,N_18913);
and U25522 (N_25522,N_23477,N_23174);
nor U25523 (N_25523,N_21737,N_22045);
xor U25524 (N_25524,N_20286,N_18574);
xnor U25525 (N_25525,N_20368,N_23663);
xnor U25526 (N_25526,N_20283,N_23847);
nand U25527 (N_25527,N_18113,N_18876);
nand U25528 (N_25528,N_23759,N_20585);
and U25529 (N_25529,N_19597,N_19913);
xor U25530 (N_25530,N_21795,N_19614);
nand U25531 (N_25531,N_23669,N_23977);
xnor U25532 (N_25532,N_22070,N_20263);
nor U25533 (N_25533,N_22921,N_22615);
and U25534 (N_25534,N_18091,N_23034);
nand U25535 (N_25535,N_20336,N_20825);
xnor U25536 (N_25536,N_23602,N_21996);
nand U25537 (N_25537,N_20705,N_18719);
nand U25538 (N_25538,N_20239,N_18831);
xor U25539 (N_25539,N_23412,N_20496);
xor U25540 (N_25540,N_23293,N_19252);
nor U25541 (N_25541,N_21107,N_23729);
xnor U25542 (N_25542,N_20258,N_20110);
nor U25543 (N_25543,N_20356,N_21077);
nand U25544 (N_25544,N_21434,N_22622);
and U25545 (N_25545,N_18911,N_20726);
nand U25546 (N_25546,N_22904,N_21677);
or U25547 (N_25547,N_19418,N_20372);
nand U25548 (N_25548,N_21454,N_23442);
and U25549 (N_25549,N_20376,N_23182);
or U25550 (N_25550,N_18809,N_20520);
nand U25551 (N_25551,N_20446,N_23558);
nor U25552 (N_25552,N_19000,N_19690);
or U25553 (N_25553,N_22010,N_21067);
nand U25554 (N_25554,N_19265,N_19056);
nor U25555 (N_25555,N_22590,N_22041);
xnor U25556 (N_25556,N_22454,N_23543);
or U25557 (N_25557,N_22181,N_22100);
or U25558 (N_25558,N_20579,N_23380);
nor U25559 (N_25559,N_19752,N_21072);
nor U25560 (N_25560,N_23586,N_22055);
xor U25561 (N_25561,N_22395,N_21712);
nand U25562 (N_25562,N_22549,N_21158);
and U25563 (N_25563,N_23887,N_18020);
nand U25564 (N_25564,N_20262,N_19753);
nor U25565 (N_25565,N_22551,N_23123);
xnor U25566 (N_25566,N_22160,N_21277);
nor U25567 (N_25567,N_18684,N_21528);
nand U25568 (N_25568,N_20626,N_18355);
or U25569 (N_25569,N_20582,N_21782);
or U25570 (N_25570,N_19029,N_21103);
nand U25571 (N_25571,N_22633,N_21893);
nand U25572 (N_25572,N_20033,N_23001);
nor U25573 (N_25573,N_22643,N_19576);
or U25574 (N_25574,N_21240,N_18111);
nor U25575 (N_25575,N_23530,N_18556);
or U25576 (N_25576,N_23253,N_21015);
xnor U25577 (N_25577,N_19678,N_21203);
xor U25578 (N_25578,N_22136,N_23830);
or U25579 (N_25579,N_22228,N_22020);
xor U25580 (N_25580,N_19604,N_23437);
xnor U25581 (N_25581,N_20381,N_20974);
nor U25582 (N_25582,N_18092,N_20127);
nor U25583 (N_25583,N_22248,N_18557);
or U25584 (N_25584,N_22066,N_18634);
and U25585 (N_25585,N_20539,N_21375);
and U25586 (N_25586,N_20918,N_21412);
or U25587 (N_25587,N_23154,N_18603);
and U25588 (N_25588,N_23287,N_22983);
nor U25589 (N_25589,N_18390,N_23909);
nor U25590 (N_25590,N_22914,N_22809);
xnor U25591 (N_25591,N_20996,N_21245);
nor U25592 (N_25592,N_23116,N_21672);
nand U25593 (N_25593,N_23145,N_20700);
nor U25594 (N_25594,N_23526,N_18987);
nor U25595 (N_25595,N_18864,N_20987);
nor U25596 (N_25596,N_22317,N_22108);
nor U25597 (N_25597,N_22697,N_22679);
or U25598 (N_25598,N_21658,N_20805);
nand U25599 (N_25599,N_18002,N_19872);
nor U25600 (N_25600,N_19648,N_20065);
nand U25601 (N_25601,N_18056,N_23185);
nand U25602 (N_25602,N_19961,N_20131);
and U25603 (N_25603,N_18593,N_19423);
xor U25604 (N_25604,N_23057,N_18860);
or U25605 (N_25605,N_22561,N_18317);
xor U25606 (N_25606,N_19402,N_21201);
or U25607 (N_25607,N_22768,N_19505);
and U25608 (N_25608,N_20622,N_22146);
or U25609 (N_25609,N_19226,N_22680);
nor U25610 (N_25610,N_22903,N_18142);
nand U25611 (N_25611,N_21114,N_22731);
nand U25612 (N_25612,N_20070,N_23613);
xor U25613 (N_25613,N_18467,N_20649);
nor U25614 (N_25614,N_22506,N_23463);
or U25615 (N_25615,N_23216,N_19138);
and U25616 (N_25616,N_19186,N_22024);
and U25617 (N_25617,N_21544,N_20848);
and U25618 (N_25618,N_18097,N_21352);
nand U25619 (N_25619,N_18753,N_23722);
and U25620 (N_25620,N_22521,N_20503);
nand U25621 (N_25621,N_22023,N_20119);
xor U25622 (N_25622,N_23585,N_23925);
xnor U25623 (N_25623,N_23343,N_20899);
xor U25624 (N_25624,N_22073,N_20498);
xor U25625 (N_25625,N_22090,N_19993);
nand U25626 (N_25626,N_23320,N_22749);
nor U25627 (N_25627,N_22252,N_19309);
or U25628 (N_25628,N_18767,N_21509);
and U25629 (N_25629,N_23061,N_23141);
nand U25630 (N_25630,N_18654,N_22500);
nor U25631 (N_25631,N_22683,N_20879);
nor U25632 (N_25632,N_23136,N_23790);
xor U25633 (N_25633,N_21521,N_20581);
and U25634 (N_25634,N_23813,N_21255);
or U25635 (N_25635,N_22664,N_21365);
xnor U25636 (N_25636,N_18570,N_19286);
nor U25637 (N_25637,N_18155,N_23053);
or U25638 (N_25638,N_18664,N_20972);
xor U25639 (N_25639,N_18688,N_22162);
xor U25640 (N_25640,N_18371,N_23302);
and U25641 (N_25641,N_20956,N_21430);
nor U25642 (N_25642,N_21093,N_19949);
nand U25643 (N_25643,N_20528,N_18962);
nor U25644 (N_25644,N_18327,N_18386);
nand U25645 (N_25645,N_18395,N_20724);
nor U25646 (N_25646,N_21356,N_19433);
and U25647 (N_25647,N_23600,N_23157);
nand U25648 (N_25648,N_19174,N_22578);
nand U25649 (N_25649,N_19610,N_19836);
nor U25650 (N_25650,N_22344,N_19826);
or U25651 (N_25651,N_21351,N_21548);
nor U25652 (N_25652,N_21394,N_23858);
and U25653 (N_25653,N_20205,N_21653);
or U25654 (N_25654,N_20648,N_21761);
nand U25655 (N_25655,N_23831,N_19711);
nand U25656 (N_25656,N_23686,N_18254);
xor U25657 (N_25657,N_20815,N_18873);
xor U25658 (N_25658,N_22563,N_23659);
nand U25659 (N_25659,N_21538,N_23374);
xor U25660 (N_25660,N_18572,N_18852);
xnor U25661 (N_25661,N_21156,N_20282);
nor U25662 (N_25662,N_21536,N_22429);
nand U25663 (N_25663,N_19688,N_23689);
or U25664 (N_25664,N_22623,N_21296);
and U25665 (N_25665,N_19343,N_22703);
or U25666 (N_25666,N_21328,N_18564);
nand U25667 (N_25667,N_22676,N_20602);
or U25668 (N_25668,N_22771,N_20637);
and U25669 (N_25669,N_22309,N_22900);
or U25670 (N_25670,N_21247,N_19535);
nor U25671 (N_25671,N_23872,N_20739);
nand U25672 (N_25672,N_22442,N_20032);
nand U25673 (N_25673,N_18687,N_19769);
nor U25674 (N_25674,N_18085,N_20482);
or U25675 (N_25675,N_20729,N_23773);
or U25676 (N_25676,N_23391,N_18533);
nor U25677 (N_25677,N_21772,N_23324);
and U25678 (N_25678,N_21885,N_19570);
and U25679 (N_25679,N_23556,N_21559);
xnor U25680 (N_25680,N_18973,N_18466);
nor U25681 (N_25681,N_19684,N_23965);
xor U25682 (N_25682,N_23114,N_20172);
xnor U25683 (N_25683,N_20691,N_19856);
or U25684 (N_25684,N_19707,N_20026);
nor U25685 (N_25685,N_20806,N_20869);
nand U25686 (N_25686,N_21892,N_19201);
nand U25687 (N_25687,N_18773,N_19098);
nor U25688 (N_25688,N_22534,N_20596);
and U25689 (N_25689,N_20383,N_23260);
and U25690 (N_25690,N_23171,N_20607);
xor U25691 (N_25691,N_19090,N_21838);
nor U25692 (N_25692,N_22329,N_23089);
nor U25693 (N_25693,N_23612,N_19650);
xnor U25694 (N_25694,N_20341,N_23289);
nand U25695 (N_25695,N_20711,N_20954);
or U25696 (N_25696,N_19770,N_20978);
xor U25697 (N_25697,N_22290,N_21308);
xor U25698 (N_25698,N_19364,N_21734);
and U25699 (N_25699,N_20611,N_19106);
nor U25700 (N_25700,N_19549,N_18365);
and U25701 (N_25701,N_20864,N_19795);
xnor U25702 (N_25702,N_23571,N_18123);
nor U25703 (N_25703,N_19721,N_19526);
and U25704 (N_25704,N_22255,N_19124);
nand U25705 (N_25705,N_22844,N_23721);
xnor U25706 (N_25706,N_21539,N_22923);
and U25707 (N_25707,N_18583,N_22953);
or U25708 (N_25708,N_21659,N_19198);
xor U25709 (N_25709,N_18835,N_18716);
xnor U25710 (N_25710,N_20266,N_19954);
nor U25711 (N_25711,N_18947,N_19202);
nand U25712 (N_25712,N_22332,N_19898);
xnor U25713 (N_25713,N_22089,N_19858);
or U25714 (N_25714,N_21066,N_22403);
or U25715 (N_25715,N_19581,N_22691);
nand U25716 (N_25716,N_21040,N_23848);
and U25717 (N_25717,N_21413,N_19663);
and U25718 (N_25718,N_21816,N_19094);
xor U25719 (N_25719,N_20423,N_21875);
and U25720 (N_25720,N_19022,N_19910);
and U25721 (N_25721,N_22057,N_22934);
or U25722 (N_25722,N_18090,N_21655);
or U25723 (N_25723,N_20236,N_18764);
nand U25724 (N_25724,N_18373,N_21065);
xor U25725 (N_25725,N_20257,N_18060);
xnor U25726 (N_25726,N_21906,N_23559);
xor U25727 (N_25727,N_19847,N_22857);
xor U25728 (N_25728,N_20187,N_18810);
nand U25729 (N_25729,N_19156,N_20458);
or U25730 (N_25730,N_21187,N_20319);
or U25731 (N_25731,N_18184,N_22221);
nand U25732 (N_25732,N_22061,N_22258);
nor U25733 (N_25733,N_22599,N_19880);
or U25734 (N_25734,N_20020,N_21493);
nor U25735 (N_25735,N_23490,N_22280);
or U25736 (N_25736,N_22319,N_19790);
or U25737 (N_25737,N_23881,N_20494);
nor U25738 (N_25738,N_18082,N_22555);
nor U25739 (N_25739,N_23737,N_20430);
nand U25740 (N_25740,N_20214,N_23919);
or U25741 (N_25741,N_22772,N_22828);
nand U25742 (N_25742,N_18146,N_22210);
or U25743 (N_25743,N_18223,N_23005);
nor U25744 (N_25744,N_20632,N_19727);
or U25745 (N_25745,N_18079,N_18596);
or U25746 (N_25746,N_20500,N_22232);
xor U25747 (N_25747,N_23564,N_22071);
nor U25748 (N_25748,N_19448,N_19837);
nor U25749 (N_25749,N_21696,N_20234);
and U25750 (N_25750,N_18907,N_20419);
xor U25751 (N_25751,N_22881,N_22114);
or U25752 (N_25752,N_22373,N_22581);
nor U25753 (N_25753,N_18035,N_19052);
or U25754 (N_25754,N_19277,N_20276);
or U25755 (N_25755,N_20401,N_23310);
and U25756 (N_25756,N_18131,N_19661);
nor U25757 (N_25757,N_21224,N_18134);
nor U25758 (N_25758,N_18300,N_21395);
nor U25759 (N_25759,N_23085,N_19082);
and U25760 (N_25760,N_22835,N_23108);
nand U25761 (N_25761,N_19787,N_20133);
nor U25762 (N_25762,N_21880,N_23555);
or U25763 (N_25763,N_18768,N_21417);
and U25764 (N_25764,N_23824,N_20841);
nand U25765 (N_25765,N_18494,N_19338);
xnor U25766 (N_25766,N_23036,N_21751);
nand U25767 (N_25767,N_20073,N_19644);
and U25768 (N_25768,N_21419,N_20450);
and U25769 (N_25769,N_19586,N_19772);
xnor U25770 (N_25770,N_19155,N_20655);
xor U25771 (N_25771,N_20809,N_21033);
xor U25772 (N_25772,N_19008,N_21970);
nand U25773 (N_25773,N_23709,N_22815);
xor U25774 (N_25774,N_21904,N_19908);
and U25775 (N_25775,N_18576,N_20087);
or U25776 (N_25776,N_23705,N_22427);
nand U25777 (N_25777,N_19883,N_23304);
xnor U25778 (N_25778,N_22190,N_21346);
nand U25779 (N_25779,N_23321,N_20461);
and U25780 (N_25780,N_18642,N_23812);
and U25781 (N_25781,N_21345,N_18463);
or U25782 (N_25782,N_22410,N_20321);
nand U25783 (N_25783,N_19967,N_18613);
and U25784 (N_25784,N_18166,N_21316);
or U25785 (N_25785,N_23575,N_18777);
nand U25786 (N_25786,N_20313,N_23544);
xor U25787 (N_25787,N_22085,N_19432);
or U25788 (N_25788,N_22385,N_22665);
nand U25789 (N_25789,N_23288,N_23993);
or U25790 (N_25790,N_18136,N_20183);
or U25791 (N_25791,N_18271,N_19499);
nor U25792 (N_25792,N_22274,N_23524);
nand U25793 (N_25793,N_19428,N_23632);
or U25794 (N_25794,N_23048,N_20391);
and U25795 (N_25795,N_21989,N_21474);
xnor U25796 (N_25796,N_22539,N_23480);
and U25797 (N_25797,N_19739,N_19508);
nor U25798 (N_25798,N_22608,N_18305);
nor U25799 (N_25799,N_21408,N_21755);
and U25800 (N_25800,N_20489,N_23214);
nor U25801 (N_25801,N_19061,N_22626);
and U25802 (N_25802,N_20394,N_18222);
or U25803 (N_25803,N_22570,N_21687);
nand U25804 (N_25804,N_23247,N_18752);
nor U25805 (N_25805,N_20344,N_19209);
nor U25806 (N_25806,N_21636,N_22911);
or U25807 (N_25807,N_23878,N_18211);
and U25808 (N_25808,N_21368,N_18499);
or U25809 (N_25809,N_20823,N_19689);
xor U25810 (N_25810,N_21867,N_20010);
or U25811 (N_25811,N_19307,N_19823);
or U25812 (N_25812,N_23743,N_20456);
and U25813 (N_25813,N_20031,N_20555);
xor U25814 (N_25814,N_18426,N_23308);
nand U25815 (N_25815,N_22887,N_19536);
nor U25816 (N_25816,N_20273,N_21034);
xnor U25817 (N_25817,N_22343,N_23749);
or U25818 (N_25818,N_22091,N_18246);
nand U25819 (N_25819,N_21124,N_21478);
and U25820 (N_25820,N_19705,N_23115);
and U25821 (N_25821,N_22907,N_20388);
xnor U25822 (N_25822,N_20101,N_20393);
and U25823 (N_25823,N_20568,N_19555);
or U25824 (N_25824,N_19885,N_22321);
and U25825 (N_25825,N_21135,N_20681);
xor U25826 (N_25826,N_20685,N_18258);
or U25827 (N_25827,N_22794,N_23792);
or U25828 (N_25828,N_23044,N_23476);
and U25829 (N_25829,N_22662,N_21833);
nand U25830 (N_25830,N_19311,N_21145);
or U25831 (N_25831,N_20735,N_20730);
nand U25832 (N_25832,N_19001,N_21359);
or U25833 (N_25833,N_19832,N_19515);
nor U25834 (N_25834,N_18755,N_22514);
or U25835 (N_25835,N_21707,N_19270);
or U25836 (N_25836,N_22840,N_20571);
nand U25837 (N_25837,N_18268,N_18442);
nor U25838 (N_25838,N_22046,N_21807);
xor U25839 (N_25839,N_18387,N_20935);
and U25840 (N_25840,N_18782,N_19735);
or U25841 (N_25841,N_21445,N_19142);
xor U25842 (N_25842,N_20567,N_22205);
nand U25843 (N_25843,N_20614,N_19233);
and U25844 (N_25844,N_21315,N_19559);
and U25845 (N_25845,N_19602,N_19518);
and U25846 (N_25846,N_22997,N_20688);
or U25847 (N_25847,N_18116,N_20292);
or U25848 (N_25848,N_23290,N_21726);
and U25849 (N_25849,N_20117,N_21900);
or U25850 (N_25850,N_20893,N_21139);
nor U25851 (N_25851,N_21425,N_21806);
nand U25852 (N_25852,N_18276,N_20333);
and U25853 (N_25853,N_23256,N_18279);
nor U25854 (N_25854,N_18170,N_19746);
or U25855 (N_25855,N_19638,N_23949);
or U25856 (N_25856,N_21250,N_21547);
xor U25857 (N_25857,N_20630,N_20771);
or U25858 (N_25858,N_21584,N_21644);
nand U25859 (N_25859,N_20084,N_21468);
nand U25860 (N_25860,N_19285,N_19113);
and U25861 (N_25861,N_18922,N_19069);
xnor U25862 (N_25862,N_20763,N_22817);
xor U25863 (N_25863,N_23000,N_20007);
or U25864 (N_25864,N_18710,N_23291);
xnor U25865 (N_25865,N_20378,N_20300);
nor U25866 (N_25866,N_21379,N_20299);
xnor U25867 (N_25867,N_19566,N_20210);
xnor U25868 (N_25868,N_22353,N_23415);
and U25869 (N_25869,N_19224,N_21675);
xnor U25870 (N_25870,N_22908,N_22308);
or U25871 (N_25871,N_21061,N_22298);
and U25872 (N_25872,N_19789,N_22718);
nor U25873 (N_25873,N_22922,N_20271);
nor U25874 (N_25874,N_21837,N_18859);
and U25875 (N_25875,N_20107,N_23126);
and U25876 (N_25876,N_19781,N_23625);
nor U25877 (N_25877,N_20448,N_22756);
and U25878 (N_25878,N_20253,N_18302);
xor U25879 (N_25879,N_21561,N_18580);
nand U25880 (N_25880,N_20091,N_20769);
xor U25881 (N_25881,N_19686,N_18566);
nand U25882 (N_25882,N_20130,N_20636);
or U25883 (N_25883,N_20510,N_22747);
nor U25884 (N_25884,N_23269,N_22170);
and U25885 (N_25885,N_19589,N_19628);
xnor U25886 (N_25886,N_20444,N_23850);
nand U25887 (N_25887,N_23807,N_19352);
and U25888 (N_25888,N_20452,N_21897);
or U25889 (N_25889,N_22324,N_23653);
nand U25890 (N_25890,N_23395,N_19238);
nor U25891 (N_25891,N_19047,N_20484);
xor U25892 (N_25892,N_21574,N_21724);
xor U25893 (N_25893,N_22086,N_19522);
nor U25894 (N_25894,N_18891,N_18015);
nand U25895 (N_25895,N_23345,N_18130);
and U25896 (N_25896,N_20947,N_21017);
nand U25897 (N_25897,N_23787,N_22340);
or U25898 (N_25898,N_22636,N_21170);
xor U25899 (N_25899,N_18758,N_21229);
or U25900 (N_25900,N_18227,N_20868);
nor U25901 (N_25901,N_18214,N_19580);
nor U25902 (N_25902,N_21227,N_18249);
or U25903 (N_25903,N_23075,N_18606);
nand U25904 (N_25904,N_18819,N_22287);
nand U25905 (N_25905,N_19297,N_23219);
xnor U25906 (N_25906,N_23727,N_19931);
or U25907 (N_25907,N_20141,N_19114);
xnor U25908 (N_25908,N_21631,N_22480);
nor U25909 (N_25909,N_22823,N_18711);
xor U25910 (N_25910,N_21849,N_23856);
xor U25911 (N_25911,N_21701,N_18772);
or U25912 (N_25912,N_23647,N_19396);
or U25913 (N_25913,N_21747,N_18342);
or U25914 (N_25914,N_18479,N_23098);
or U25915 (N_25915,N_22077,N_19978);
nand U25916 (N_25916,N_20505,N_18076);
and U25917 (N_25917,N_20387,N_19397);
nand U25918 (N_25918,N_20241,N_22120);
nand U25919 (N_25919,N_22188,N_20108);
nand U25920 (N_25920,N_22320,N_18528);
xor U25921 (N_25921,N_18459,N_19333);
and U25922 (N_25922,N_22753,N_18431);
nor U25923 (N_25923,N_18277,N_20188);
nor U25924 (N_25924,N_22241,N_18307);
and U25925 (N_25925,N_19463,N_18910);
and U25926 (N_25926,N_20931,N_21629);
and U25927 (N_25927,N_21300,N_21428);
nand U25928 (N_25928,N_21486,N_19251);
and U25929 (N_25929,N_23275,N_20991);
or U25930 (N_25930,N_18798,N_23199);
or U25931 (N_25931,N_18997,N_23791);
nor U25932 (N_25932,N_22411,N_23433);
and U25933 (N_25933,N_23822,N_22712);
xor U25934 (N_25934,N_19129,N_23221);
nor U25935 (N_25935,N_23497,N_21830);
nor U25936 (N_25936,N_20072,N_21441);
xnor U25937 (N_25937,N_23761,N_20501);
xor U25938 (N_25938,N_22663,N_20284);
nor U25939 (N_25939,N_23357,N_19039);
xnor U25940 (N_25940,N_19529,N_21532);
and U25941 (N_25941,N_23932,N_22198);
xnor U25942 (N_25942,N_19730,N_18964);
and U25943 (N_25943,N_18571,N_18361);
xor U25944 (N_25944,N_21193,N_20552);
and U25945 (N_25945,N_21121,N_20306);
nor U25946 (N_25946,N_22318,N_21266);
nand U25947 (N_25947,N_22967,N_20915);
nor U25948 (N_25948,N_21591,N_19749);
nand U25949 (N_25949,N_20860,N_23529);
xnor U25950 (N_25950,N_21876,N_20222);
and U25951 (N_25951,N_19668,N_20129);
or U25952 (N_25952,N_19564,N_21276);
nand U25953 (N_25953,N_18071,N_20145);
and U25954 (N_25954,N_21804,N_21043);
xor U25955 (N_25955,N_20659,N_22520);
and U25956 (N_25956,N_19015,N_20136);
and U25957 (N_25957,N_23237,N_19276);
nand U25958 (N_25958,N_20804,N_18694);
and U25959 (N_25959,N_18846,N_20315);
nor U25960 (N_25960,N_22494,N_23528);
nor U25961 (N_25961,N_19934,N_23862);
nand U25962 (N_25962,N_18622,N_21008);
and U25963 (N_25963,N_20464,N_22006);
nor U25964 (N_25964,N_18458,N_23404);
xor U25965 (N_25965,N_18065,N_21265);
or U25966 (N_25966,N_20884,N_23533);
and U25967 (N_25967,N_22720,N_19685);
xnor U25968 (N_25968,N_19143,N_20039);
nand U25969 (N_25969,N_22468,N_23634);
nor U25970 (N_25970,N_21037,N_23431);
nand U25971 (N_25971,N_22168,N_19957);
and U25972 (N_25972,N_19235,N_23124);
or U25973 (N_25973,N_20838,N_22936);
nor U25974 (N_25974,N_22509,N_18406);
nand U25975 (N_25975,N_18623,N_22598);
nor U25976 (N_25976,N_20345,N_23580);
nor U25977 (N_25977,N_19643,N_21475);
nand U25978 (N_25978,N_20213,N_23491);
nand U25979 (N_25979,N_23280,N_23947);
or U25980 (N_25980,N_21556,N_19422);
nand U25981 (N_25981,N_20779,N_18098);
or U25982 (N_25982,N_18455,N_22851);
or U25983 (N_25983,N_20570,N_22596);
and U25984 (N_25984,N_23080,N_23183);
or U25985 (N_25985,N_19640,N_18404);
nand U25986 (N_25986,N_21896,N_21304);
or U25987 (N_25987,N_22877,N_22991);
or U25988 (N_25988,N_21183,N_18515);
and U25989 (N_25989,N_23377,N_22421);
or U25990 (N_25990,N_22724,N_19273);
nand U25991 (N_25991,N_20725,N_20279);
and U25992 (N_25992,N_19517,N_18651);
nor U25993 (N_25993,N_19924,N_23903);
nor U25994 (N_25994,N_18200,N_18792);
or U25995 (N_25995,N_23012,N_21973);
nor U25996 (N_25996,N_21059,N_19547);
nand U25997 (N_25997,N_21777,N_18963);
xnor U25998 (N_25998,N_23063,N_20508);
nand U25999 (N_25999,N_20680,N_18909);
and U26000 (N_26000,N_19279,N_23591);
and U26001 (N_26001,N_19972,N_22996);
nor U26002 (N_26002,N_21738,N_19895);
nor U26003 (N_26003,N_18328,N_19367);
xor U26004 (N_26004,N_22689,N_18288);
nor U26005 (N_26005,N_23228,N_18975);
or U26006 (N_26006,N_23982,N_21732);
nand U26007 (N_26007,N_22446,N_20922);
nand U26008 (N_26008,N_22577,N_19062);
and U26009 (N_26009,N_18998,N_22982);
and U26010 (N_26010,N_21314,N_22806);
or U26011 (N_26011,N_18210,N_20397);
or U26012 (N_26012,N_21827,N_22515);
nor U26013 (N_26013,N_20042,N_23074);
xnor U26014 (N_26014,N_19048,N_22448);
and U26015 (N_26015,N_19840,N_21743);
xnor U26016 (N_26016,N_21702,N_18587);
or U26017 (N_26017,N_22895,N_23164);
nand U26018 (N_26018,N_21718,N_21686);
nand U26019 (N_26019,N_21907,N_19120);
and U26020 (N_26020,N_18658,N_21587);
nor U26021 (N_26021,N_23865,N_19512);
xnor U26022 (N_26022,N_23608,N_23621);
xor U26023 (N_26023,N_18858,N_20742);
and U26024 (N_26024,N_20589,N_23118);
and U26025 (N_26025,N_23879,N_21216);
nand U26026 (N_26026,N_18512,N_20892);
and U26027 (N_26027,N_20499,N_20923);
nand U26028 (N_26028,N_21019,N_20439);
or U26029 (N_26029,N_22366,N_21382);
xor U26030 (N_26030,N_20082,N_21502);
xnor U26031 (N_26031,N_22179,N_22624);
and U26032 (N_26032,N_18026,N_20610);
nand U26033 (N_26033,N_20646,N_19263);
nor U26034 (N_26034,N_21016,N_22381);
or U26035 (N_26035,N_20562,N_18280);
nor U26036 (N_26036,N_23331,N_18608);
and U26037 (N_26037,N_19361,N_18638);
xor U26038 (N_26038,N_19497,N_22052);
nor U26039 (N_26039,N_21424,N_20798);
and U26040 (N_26040,N_23976,N_18005);
nand U26041 (N_26041,N_23201,N_22153);
nand U26042 (N_26042,N_18935,N_18919);
nand U26043 (N_26043,N_21291,N_21619);
nor U26044 (N_26044,N_23245,N_18763);
nor U26045 (N_26045,N_19775,N_18633);
nand U26046 (N_26046,N_18769,N_23957);
or U26047 (N_26047,N_22945,N_21488);
xor U26048 (N_26048,N_23573,N_23746);
and U26049 (N_26049,N_19556,N_21588);
or U26050 (N_26050,N_23884,N_22233);
nor U26051 (N_26051,N_21933,N_19185);
nor U26052 (N_26052,N_19162,N_22288);
nor U26053 (N_26053,N_23987,N_21403);
xor U26054 (N_26054,N_19254,N_20640);
xnor U26055 (N_26055,N_22804,N_23033);
and U26056 (N_26056,N_20556,N_21886);
xnor U26057 (N_26057,N_21032,N_20993);
and U26058 (N_26058,N_20245,N_19531);
xnor U26059 (N_26059,N_23095,N_23306);
xor U26060 (N_26060,N_23570,N_18415);
and U26061 (N_26061,N_22276,N_23451);
nand U26062 (N_26062,N_19362,N_23960);
or U26063 (N_26063,N_20060,N_22272);
nand U26064 (N_26064,N_21899,N_22788);
nand U26065 (N_26065,N_23752,N_18837);
nor U26066 (N_26066,N_21357,N_20690);
xor U26067 (N_26067,N_21853,N_19855);
or U26068 (N_26068,N_19745,N_23311);
nand U26069 (N_26069,N_19055,N_23841);
nor U26070 (N_26070,N_22893,N_21998);
nor U26071 (N_26071,N_20554,N_21879);
and U26072 (N_26072,N_18966,N_22397);
nor U26073 (N_26073,N_19239,N_18995);
nor U26074 (N_26074,N_23901,N_19444);
nand U26075 (N_26075,N_19827,N_21137);
nand U26076 (N_26076,N_20097,N_20272);
xnor U26077 (N_26077,N_21360,N_22586);
or U26078 (N_26078,N_21451,N_21169);
and U26079 (N_26079,N_19359,N_21142);
or U26080 (N_26080,N_19148,N_22740);
xnor U26081 (N_26081,N_20320,N_21044);
xnor U26082 (N_26082,N_19220,N_23521);
nor U26083 (N_26083,N_21864,N_18332);
nand U26084 (N_26084,N_21982,N_20566);
or U26085 (N_26085,N_23691,N_20475);
nand U26086 (N_26086,N_23493,N_23496);
or U26087 (N_26087,N_21802,N_23013);
nor U26088 (N_26088,N_18640,N_23091);
nor U26089 (N_26089,N_22419,N_22432);
xor U26090 (N_26090,N_22878,N_22905);
and U26091 (N_26091,N_22169,N_23683);
nand U26092 (N_26092,N_19894,N_21656);
and U26093 (N_26093,N_22044,N_21453);
and U26094 (N_26094,N_20352,N_19100);
nand U26095 (N_26095,N_18383,N_18560);
xor U26096 (N_26096,N_22609,N_21244);
or U26097 (N_26097,N_21563,N_19161);
nand U26098 (N_26098,N_23695,N_20550);
and U26099 (N_26099,N_21136,N_23170);
and U26100 (N_26100,N_18851,N_22869);
and U26101 (N_26101,N_22888,N_21207);
nor U26102 (N_26102,N_19887,N_23974);
or U26103 (N_26103,N_23188,N_20062);
nor U26104 (N_26104,N_20796,N_20671);
and U26105 (N_26105,N_19716,N_23646);
and U26106 (N_26106,N_21725,N_18712);
nor U26107 (N_26107,N_23549,N_19946);
xnor U26108 (N_26108,N_20018,N_19977);
nor U26109 (N_26109,N_20075,N_22677);
nand U26110 (N_26110,N_18061,N_22076);
and U26111 (N_26111,N_22550,N_19915);
or U26112 (N_26112,N_20051,N_21353);
or U26113 (N_26113,N_19344,N_23639);
or U26114 (N_26114,N_19150,N_23924);
nor U26115 (N_26115,N_23617,N_19467);
xor U26116 (N_26116,N_21489,N_18704);
and U26117 (N_26117,N_21058,N_22507);
and U26118 (N_26118,N_21964,N_21870);
xnor U26119 (N_26119,N_18992,N_21028);
nand U26120 (N_26120,N_22767,N_18590);
xor U26121 (N_26121,N_18616,N_18558);
xor U26122 (N_26122,N_23945,N_19031);
nor U26123 (N_26123,N_22390,N_19796);
or U26124 (N_26124,N_22736,N_20963);
xnor U26125 (N_26125,N_18743,N_23055);
nand U26126 (N_26126,N_18601,N_20839);
nand U26127 (N_26127,N_20749,N_23094);
xor U26128 (N_26128,N_21988,N_23733);
nand U26129 (N_26129,N_23910,N_23598);
and U26130 (N_26130,N_22072,N_22372);
or U26131 (N_26131,N_21604,N_23921);
xor U26132 (N_26132,N_19257,N_19618);
nand U26133 (N_26133,N_18141,N_22535);
nor U26134 (N_26134,N_19989,N_20728);
and U26135 (N_26135,N_22414,N_21679);
nand U26136 (N_26136,N_21487,N_19941);
and U26137 (N_26137,N_21214,N_19407);
xor U26138 (N_26138,N_20656,N_21483);
nor U26139 (N_26139,N_18617,N_23081);
or U26140 (N_26140,N_23892,N_23664);
xor U26141 (N_26141,N_21079,N_18186);
nand U26142 (N_26142,N_20185,N_21639);
nand U26143 (N_26143,N_22423,N_19550);
and U26144 (N_26144,N_22819,N_21637);
and U26145 (N_26145,N_20113,N_21632);
and U26146 (N_26146,N_21520,N_23242);
or U26147 (N_26147,N_22635,N_19380);
nor U26148 (N_26148,N_19681,N_22822);
nand U26149 (N_26149,N_22075,N_23131);
nor U26150 (N_26150,N_20537,N_21898);
or U26151 (N_26151,N_23742,N_21527);
and U26152 (N_26152,N_20229,N_21366);
and U26153 (N_26153,N_18748,N_20047);
or U26154 (N_26154,N_23877,N_21306);
or U26155 (N_26155,N_20733,N_19255);
or U26156 (N_26156,N_20182,N_23176);
and U26157 (N_26157,N_19041,N_19459);
nor U26158 (N_26158,N_23775,N_22470);
nor U26159 (N_26159,N_23964,N_20651);
nor U26160 (N_26160,N_19134,N_22081);
nor U26161 (N_26161,N_19057,N_18024);
or U26162 (N_26162,N_23117,N_18787);
or U26163 (N_26163,N_21331,N_23125);
nand U26164 (N_26164,N_18843,N_22805);
nand U26165 (N_26165,N_23278,N_22883);
xnor U26166 (N_26166,N_20398,N_20179);
nand U26167 (N_26167,N_19568,N_22977);
and U26168 (N_26168,N_18594,N_22755);
and U26169 (N_26169,N_19347,N_20223);
or U26170 (N_26170,N_21704,N_22140);
xnor U26171 (N_26171,N_20873,N_21552);
nor U26172 (N_26172,N_21874,N_23128);
nor U26173 (N_26173,N_21284,N_23803);
or U26174 (N_26174,N_23821,N_18885);
xor U26175 (N_26175,N_23056,N_19206);
nor U26176 (N_26176,N_20736,N_20880);
or U26177 (N_26177,N_22742,N_19305);
nor U26178 (N_26178,N_19127,N_21746);
nor U26179 (N_26179,N_20799,N_18360);
xor U26180 (N_26180,N_23459,N_23329);
xnor U26181 (N_26181,N_18350,N_18996);
and U26182 (N_26182,N_21641,N_18630);
or U26183 (N_26183,N_23382,N_23388);
nor U26184 (N_26184,N_19293,N_22490);
nor U26185 (N_26185,N_22225,N_18296);
nand U26186 (N_26186,N_21498,N_22705);
nor U26187 (N_26187,N_22864,N_23372);
nand U26188 (N_26188,N_19187,N_23717);
or U26189 (N_26189,N_21377,N_20653);
nor U26190 (N_26190,N_23436,N_22444);
and U26191 (N_26191,N_19068,N_21773);
nand U26192 (N_26192,N_23844,N_18779);
xnor U26193 (N_26193,N_20563,N_20902);
and U26194 (N_26194,N_21431,N_23916);
nor U26195 (N_26195,N_20447,N_23041);
or U26196 (N_26196,N_23079,N_20647);
or U26197 (N_26197,N_20121,N_18529);
xor U26198 (N_26198,N_18632,N_21289);
or U26199 (N_26199,N_19248,N_18133);
xor U26200 (N_26200,N_19869,N_20577);
or U26201 (N_26201,N_21928,N_23078);
xor U26202 (N_26202,N_18132,N_19540);
and U26203 (N_26203,N_22573,N_19594);
nor U26204 (N_26204,N_18247,N_18656);
nor U26205 (N_26205,N_20061,N_20495);
xor U26206 (N_26206,N_22604,N_18465);
and U26207 (N_26207,N_23322,N_20784);
nand U26208 (N_26208,N_20979,N_22074);
or U26209 (N_26209,N_21387,N_18283);
or U26210 (N_26210,N_23358,N_19473);
nand U26211 (N_26211,N_22687,N_21991);
nor U26212 (N_26212,N_23926,N_20206);
nand U26213 (N_26213,N_18932,N_19504);
nand U26214 (N_26214,N_19503,N_22351);
nor U26215 (N_26215,N_19492,N_22175);
xor U26216 (N_26216,N_20190,N_20569);
nor U26217 (N_26217,N_21887,N_23326);
nand U26218 (N_26218,N_23015,N_23250);
xor U26219 (N_26219,N_19964,N_18954);
or U26220 (N_26220,N_23568,N_21764);
nor U26221 (N_26221,N_22249,N_23991);
or U26222 (N_26222,N_21566,N_19571);
and U26223 (N_26223,N_18192,N_21709);
and U26224 (N_26224,N_20677,N_18019);
and U26225 (N_26225,N_20858,N_18311);
xor U26226 (N_26226,N_19430,N_18957);
or U26227 (N_26227,N_20104,N_19649);
nand U26228 (N_26228,N_20194,N_23153);
nand U26229 (N_26229,N_22166,N_20265);
xnor U26230 (N_26230,N_21936,N_23601);
xor U26231 (N_26231,N_21727,N_19205);
nor U26232 (N_26232,N_21765,N_21578);
xor U26233 (N_26233,N_21844,N_20756);
xnor U26234 (N_26234,N_18542,N_19269);
nand U26235 (N_26235,N_19679,N_23994);
or U26236 (N_26236,N_21919,N_21676);
xor U26237 (N_26237,N_20723,N_20540);
xnor U26238 (N_26238,N_22376,N_19694);
nor U26239 (N_26239,N_23027,N_20308);
xor U26240 (N_26240,N_18985,N_20369);
and U26241 (N_26241,N_22528,N_21763);
xnor U26242 (N_26242,N_18336,N_23636);
or U26243 (N_26243,N_19636,N_19501);
xnor U26244 (N_26244,N_18320,N_22396);
and U26245 (N_26245,N_23605,N_22103);
nor U26246 (N_26246,N_20657,N_23367);
xnor U26247 (N_26247,N_21661,N_20486);
or U26248 (N_26248,N_23254,N_20761);
xnor U26249 (N_26249,N_23997,N_23104);
nand U26250 (N_26250,N_23319,N_21140);
xnor U26251 (N_26251,N_22548,N_18203);
nor U26252 (N_26252,N_23667,N_22670);
and U26253 (N_26253,N_21199,N_20881);
and U26254 (N_26254,N_23178,N_22946);
xor U26255 (N_26255,N_20613,N_20493);
or U26256 (N_26256,N_18126,N_23414);
and U26257 (N_26257,N_18790,N_21858);
and U26258 (N_26258,N_22706,N_20998);
or U26259 (N_26259,N_19072,N_20362);
nor U26260 (N_26260,N_22124,N_22131);
and U26261 (N_26261,N_23482,N_22529);
nor U26262 (N_26262,N_19692,N_22734);
nand U26263 (N_26263,N_20748,N_20938);
nand U26264 (N_26264,N_20332,N_19036);
or U26265 (N_26265,N_20672,N_21975);
or U26266 (N_26266,N_23111,N_19747);
nor U26267 (N_26267,N_18967,N_23569);
or U26268 (N_26268,N_20906,N_18046);
nor U26269 (N_26269,N_20305,N_20773);
or U26270 (N_26270,N_23038,N_18549);
or U26271 (N_26271,N_20603,N_19599);
nor U26272 (N_26272,N_23342,N_22375);
or U26273 (N_26273,N_22992,N_18621);
or U26274 (N_26274,N_22275,N_19491);
xnor U26275 (N_26275,N_23565,N_23465);
or U26276 (N_26276,N_18495,N_19232);
and U26277 (N_26277,N_22471,N_19222);
nor U26278 (N_26278,N_22886,N_19812);
or U26279 (N_26279,N_23099,N_21459);
xnor U26280 (N_26280,N_21343,N_21526);
xnor U26281 (N_26281,N_20100,N_18803);
nor U26282 (N_26282,N_21821,N_20719);
nand U26283 (N_26283,N_20242,N_18974);
nand U26284 (N_26284,N_20497,N_21515);
or U26285 (N_26285,N_20980,N_19165);
and U26286 (N_26286,N_23696,N_19455);
and U26287 (N_26287,N_20949,N_18239);
nand U26288 (N_26288,N_22137,N_21223);
and U26289 (N_26289,N_21175,N_21760);
and U26290 (N_26290,N_22415,N_23531);
xnor U26291 (N_26291,N_22968,N_21634);
nand U26292 (N_26292,N_21176,N_20689);
and U26293 (N_26293,N_18378,N_19002);
and U26294 (N_26294,N_19857,N_23732);
nand U26295 (N_26295,N_20578,N_19734);
and U26296 (N_26296,N_23935,N_20803);
nand U26297 (N_26297,N_23798,N_22602);
or U26298 (N_26298,N_21608,N_19963);
nand U26299 (N_26299,N_19130,N_18933);
nand U26300 (N_26300,N_22744,N_19748);
nand U26301 (N_26301,N_23682,N_19496);
and U26302 (N_26302,N_19569,N_21001);
nor U26303 (N_26303,N_20233,N_19488);
nor U26304 (N_26304,N_18552,N_21976);
and U26305 (N_26305,N_18525,N_19776);
nand U26306 (N_26306,N_20976,N_21143);
nand U26307 (N_26307,N_18161,N_22950);
nand U26308 (N_26308,N_18898,N_21579);
xnor U26309 (N_26309,N_20802,N_23265);
xnor U26310 (N_26310,N_20106,N_19014);
and U26311 (N_26311,N_21605,N_21616);
nor U26312 (N_26312,N_23904,N_20676);
and U26313 (N_26313,N_23359,N_23678);
or U26314 (N_26314,N_18659,N_20404);
nand U26315 (N_26315,N_21210,N_22695);
xnor U26316 (N_26316,N_20594,N_20259);
nand U26317 (N_26317,N_19033,N_21036);
xor U26318 (N_26318,N_18181,N_22182);
xnor U26319 (N_26319,N_21358,N_23452);
nor U26320 (N_26320,N_19817,N_21014);
and U26321 (N_26321,N_19603,N_22545);
and U26322 (N_26322,N_18410,N_23970);
or U26323 (N_26323,N_22333,N_19616);
or U26324 (N_26324,N_22214,N_19028);
or U26325 (N_26325,N_19168,N_18492);
or U26326 (N_26326,N_18094,N_19891);
or U26327 (N_26327,N_21166,N_18033);
nand U26328 (N_26328,N_19548,N_23679);
or U26329 (N_26329,N_22960,N_18745);
or U26330 (N_26330,N_18671,N_19715);
xnor U26331 (N_26331,N_21126,N_22918);
or U26332 (N_26332,N_22109,N_21918);
nor U26333 (N_26333,N_22765,N_22627);
and U26334 (N_26334,N_18931,N_18771);
or U26335 (N_26335,N_19619,N_20364);
xor U26336 (N_26336,N_21922,N_23692);
or U26337 (N_26337,N_23805,N_23158);
or U26338 (N_26338,N_21329,N_23560);
or U26339 (N_26339,N_18849,N_20184);
and U26340 (N_26340,N_18163,N_22873);
nor U26341 (N_26341,N_18976,N_18437);
and U26342 (N_26342,N_19742,N_23816);
xor U26343 (N_26343,N_21257,N_22686);
xor U26344 (N_26344,N_22836,N_20068);
and U26345 (N_26345,N_21374,N_23774);
nand U26346 (N_26346,N_18248,N_21968);
nor U26347 (N_26347,N_18830,N_22013);
nand U26348 (N_26348,N_19087,N_23337);
or U26349 (N_26349,N_21766,N_18152);
xnor U26350 (N_26350,N_21736,N_22097);
and U26351 (N_26351,N_22553,N_21129);
xor U26352 (N_26352,N_18472,N_22445);
nand U26353 (N_26353,N_21194,N_20350);
xnor U26354 (N_26354,N_22941,N_18352);
and U26355 (N_26355,N_23985,N_19927);
xnor U26356 (N_26356,N_19236,N_23532);
or U26357 (N_26357,N_23344,N_20410);
xor U26358 (N_26358,N_21338,N_20477);
nor U26359 (N_26359,N_18698,N_22030);
xnor U26360 (N_26360,N_22688,N_18345);
nor U26361 (N_26361,N_19464,N_18236);
xnor U26362 (N_26362,N_22700,N_20652);
nand U26363 (N_26363,N_22481,N_18526);
nor U26364 (N_26364,N_19093,N_20604);
nand U26365 (N_26365,N_22630,N_18118);
xnor U26366 (N_26366,N_19876,N_22681);
xnor U26367 (N_26367,N_22567,N_23251);
nand U26368 (N_26368,N_19926,N_22770);
nand U26369 (N_26369,N_18892,N_21442);
xnor U26370 (N_26370,N_20925,N_18259);
and U26371 (N_26371,N_19905,N_18188);
nand U26372 (N_26372,N_19199,N_19435);
or U26373 (N_26373,N_20895,N_18195);
nor U26374 (N_26374,N_22926,N_20277);
nand U26375 (N_26375,N_21789,N_22942);
or U26376 (N_26376,N_22758,N_18880);
nand U26377 (N_26377,N_18994,N_21878);
and U26378 (N_26378,N_22354,N_21931);
and U26379 (N_26379,N_23017,N_18066);
and U26380 (N_26380,N_22975,N_20170);
nand U26381 (N_26381,N_21189,N_19917);
and U26382 (N_26382,N_22956,N_22842);
nor U26383 (N_26383,N_21997,N_22265);
xor U26384 (N_26384,N_18812,N_22517);
nand U26385 (N_26385,N_21295,N_19598);
or U26386 (N_26386,N_19177,N_19975);
nor U26387 (N_26387,N_23241,N_21851);
nand U26388 (N_26388,N_20820,N_22939);
and U26389 (N_26389,N_20411,N_21883);
xor U26390 (N_26390,N_18032,N_22610);
or U26391 (N_26391,N_21603,N_18238);
nand U26392 (N_26392,N_20174,N_23150);
xnor U26393 (N_26393,N_22151,N_22121);
or U26394 (N_26394,N_19164,N_19696);
nor U26395 (N_26395,N_18862,N_19118);
nand U26396 (N_26396,N_18408,N_20102);
or U26397 (N_26397,N_23486,N_23177);
and U26398 (N_26398,N_22824,N_19054);
and U26399 (N_26399,N_18845,N_18232);
nand U26400 (N_26400,N_22459,N_19303);
nor U26401 (N_26401,N_22399,N_21030);
xnor U26402 (N_26402,N_21476,N_23400);
nor U26403 (N_26403,N_18478,N_23671);
or U26404 (N_26404,N_21902,N_20760);
nand U26405 (N_26405,N_22062,N_20093);
xor U26406 (N_26406,N_18683,N_18516);
and U26407 (N_26407,N_19058,N_23066);
nor U26408 (N_26408,N_21717,N_19831);
and U26409 (N_26409,N_23405,N_18847);
xnor U26410 (N_26410,N_19005,N_18274);
nand U26411 (N_26411,N_22892,N_22820);
nand U26412 (N_26412,N_19326,N_23701);
or U26413 (N_26413,N_20870,N_19354);
nand U26414 (N_26414,N_20361,N_18718);
xor U26415 (N_26415,N_18354,N_19011);
or U26416 (N_26416,N_21768,N_19541);
nor U26417 (N_26417,N_18578,N_21477);
and U26418 (N_26418,N_18701,N_22039);
nor U26419 (N_26419,N_22270,N_18637);
and U26420 (N_26420,N_19275,N_18626);
and U26421 (N_26421,N_23980,N_22088);
or U26422 (N_26422,N_23655,N_22306);
nand U26423 (N_26423,N_23146,N_21164);
and U26424 (N_26424,N_18522,N_18942);
and U26425 (N_26425,N_20541,N_22673);
xor U26426 (N_26426,N_18270,N_23143);
or U26427 (N_26427,N_21182,N_22094);
and U26428 (N_26428,N_23736,N_23699);
or U26429 (N_26429,N_23110,N_20000);
xnor U26430 (N_26430,N_21180,N_20427);
xnor U26431 (N_26431,N_18072,N_22488);
nor U26432 (N_26432,N_21808,N_21610);
xor U26433 (N_26433,N_21779,N_21071);
and U26434 (N_26434,N_23911,N_18477);
and U26435 (N_26435,N_21098,N_22019);
nor U26436 (N_26436,N_21730,N_19261);
or U26437 (N_26437,N_23438,N_18191);
xor U26438 (N_26438,N_18220,N_19625);
or U26439 (N_26439,N_21815,N_18535);
xnor U26440 (N_26440,N_21969,N_21146);
or U26441 (N_26441,N_19563,N_20379);
nand U26442 (N_26442,N_21251,N_19007);
or U26443 (N_26443,N_21534,N_22782);
and U26444 (N_26444,N_23161,N_23050);
nand U26445 (N_26445,N_23814,N_23665);
or U26446 (N_26446,N_19377,N_18937);
nand U26447 (N_26447,N_20481,N_21272);
and U26448 (N_26448,N_21426,N_18422);
and U26449 (N_26449,N_22189,N_18968);
and U26450 (N_26450,N_20877,N_21627);
and U26451 (N_26451,N_18042,N_20363);
or U26452 (N_26452,N_20453,N_21703);
nor U26453 (N_26453,N_18207,N_22644);
xor U26454 (N_26454,N_19762,N_20783);
xor U26455 (N_26455,N_23093,N_19720);
nand U26456 (N_26456,N_20629,N_21753);
nand U26457 (N_26457,N_20429,N_19470);
and U26458 (N_26458,N_19360,N_18908);
nor U26459 (N_26459,N_20402,N_23144);
and U26460 (N_26460,N_21775,N_18318);
xor U26461 (N_26461,N_20547,N_21389);
nand U26462 (N_26462,N_18749,N_18696);
and U26463 (N_26463,N_21439,N_21086);
and U26464 (N_26464,N_23152,N_20220);
or U26465 (N_26465,N_19617,N_18044);
or U26466 (N_26466,N_19712,N_23948);
nor U26467 (N_26467,N_20946,N_18620);
nand U26468 (N_26468,N_18003,N_18905);
or U26469 (N_26469,N_22648,N_18180);
and U26470 (N_26470,N_18096,N_18872);
xnor U26471 (N_26471,N_23109,N_18278);
nor U26472 (N_26472,N_18269,N_21448);
and U26473 (N_26473,N_18720,N_22341);
and U26474 (N_26474,N_21863,N_21348);
nor U26475 (N_26475,N_22450,N_19050);
xnor U26476 (N_26476,N_21745,N_22349);
or U26477 (N_26477,N_20024,N_18741);
or U26478 (N_26478,N_21275,N_19454);
and U26479 (N_26479,N_18206,N_20605);
nor U26480 (N_26480,N_21128,N_18929);
xnor U26481 (N_26481,N_20766,N_18062);
xor U26482 (N_26482,N_20967,N_19944);
nand U26483 (N_26483,N_18439,N_23180);
nand U26484 (N_26484,N_20814,N_23054);
nor U26485 (N_26485,N_23488,N_20757);
nand U26486 (N_26486,N_23922,N_22527);
and U26487 (N_26487,N_19756,N_22260);
nand U26488 (N_26488,N_21792,N_22675);
xnor U26489 (N_26489,N_23961,N_20365);
nor U26490 (N_26490,N_23998,N_23481);
or U26491 (N_26491,N_21393,N_21796);
nand U26492 (N_26492,N_19845,N_23029);
nand U26493 (N_26493,N_21213,N_22650);
xor U26494 (N_26494,N_19939,N_19356);
nand U26495 (N_26495,N_23350,N_18628);
xnor U26496 (N_26496,N_21757,N_19427);
xnor U26497 (N_26497,N_19874,N_21083);
xor U26498 (N_26498,N_23672,N_20089);
or U26499 (N_26499,N_23169,N_19096);
or U26500 (N_26500,N_19316,N_18129);
or U26501 (N_26501,N_23113,N_21960);
and U26502 (N_26502,N_23959,N_23958);
nand U26503 (N_26503,N_23540,N_21134);
or U26504 (N_26504,N_21957,N_19153);
and U26505 (N_26505,N_22178,N_19572);
or U26506 (N_26506,N_19486,N_20441);
and U26507 (N_26507,N_22989,N_23860);
nand U26508 (N_26508,N_19204,N_19868);
nand U26509 (N_26509,N_23088,N_18034);
xnor U26510 (N_26510,N_20990,N_19907);
nand U26511 (N_26511,N_19830,N_22552);
nor U26512 (N_26512,N_18403,N_22979);
nor U26513 (N_26513,N_19673,N_20357);
nand U26514 (N_26514,N_23629,N_21179);
nor U26515 (N_26515,N_18256,N_19063);
nand U26516 (N_26516,N_23370,N_21218);
nor U26517 (N_26517,N_23741,N_21501);
or U26518 (N_26518,N_18569,N_18101);
nor U26519 (N_26519,N_22406,N_20744);
or U26520 (N_26520,N_20417,N_20600);
and U26521 (N_26521,N_22102,N_21264);
nand U26522 (N_26522,N_22801,N_22999);
or U26523 (N_26523,N_22392,N_23267);
or U26524 (N_26524,N_21045,N_18853);
xor U26525 (N_26525,N_19741,N_21622);
xor U26526 (N_26526,N_18725,N_19073);
xor U26527 (N_26527,N_19509,N_21202);
xor U26528 (N_26528,N_23022,N_21595);
nand U26529 (N_26529,N_20269,N_23315);
xnor U26530 (N_26530,N_22919,N_22639);
and U26531 (N_26531,N_19751,N_22483);
nand U26532 (N_26532,N_21258,N_23739);
nand U26533 (N_26533,N_23139,N_19013);
and U26534 (N_26534,N_19223,N_21325);
or U26535 (N_26535,N_20088,N_22855);
xor U26536 (N_26536,N_18486,N_19850);
and U26537 (N_26537,N_21671,N_21020);
or U26538 (N_26538,N_20483,N_18165);
or U26539 (N_26539,N_23021,N_23567);
xor U26540 (N_26540,N_23855,N_22482);
or U26541 (N_26541,N_19947,N_23455);
or U26542 (N_26542,N_21602,N_21824);
nand U26543 (N_26543,N_18000,N_22847);
or U26544 (N_26544,N_20616,N_22485);
or U26545 (N_26545,N_21297,N_19079);
or U26546 (N_26546,N_20670,N_23194);
nand U26547 (N_26547,N_22897,N_23703);
nand U26548 (N_26548,N_20524,N_18299);
and U26549 (N_26549,N_19099,N_22486);
and U26550 (N_26550,N_21052,N_18680);
nor U26551 (N_26551,N_21075,N_21617);
and U26552 (N_26552,N_22518,N_19502);
and U26553 (N_26553,N_19542,N_20933);
xor U26554 (N_26554,N_22147,N_18879);
xnor U26555 (N_26555,N_23912,N_18058);
nor U26556 (N_26556,N_21758,N_20875);
nor U26557 (N_26557,N_20745,N_21490);
and U26558 (N_26558,N_21771,N_20390);
nand U26559 (N_26559,N_18447,N_22184);
nor U26560 (N_26560,N_22194,N_22779);
and U26561 (N_26561,N_23281,N_22789);
xnor U26562 (N_26562,N_20919,N_23435);
or U26563 (N_26563,N_19884,N_21635);
nor U26564 (N_26564,N_20790,N_19035);
nor U26565 (N_26565,N_20342,N_18043);
or U26566 (N_26566,N_20644,N_21691);
nor U26567 (N_26567,N_19267,N_18434);
nand U26568 (N_26568,N_23466,N_23874);
and U26569 (N_26569,N_22698,N_23539);
nand U26570 (N_26570,N_19437,N_20654);
nand U26571 (N_26571,N_18917,N_20830);
xor U26572 (N_26572,N_23989,N_18202);
nand U26573 (N_26573,N_21995,N_18836);
or U26574 (N_26574,N_20768,N_18840);
xor U26575 (N_26575,N_21537,N_21986);
and U26576 (N_26576,N_23936,N_20599);
xor U26577 (N_26577,N_20203,N_19076);
or U26578 (N_26578,N_21628,N_18389);
xnor U26579 (N_26579,N_22588,N_19834);
and U26580 (N_26580,N_18109,N_19456);
nor U26581 (N_26581,N_22236,N_23407);
nand U26582 (N_26582,N_18052,N_21719);
and U26583 (N_26583,N_22301,N_18639);
or U26584 (N_26584,N_18653,N_22920);
nor U26585 (N_26585,N_22852,N_18672);
nor U26586 (N_26586,N_18649,N_18901);
nor U26587 (N_26587,N_22218,N_21263);
or U26588 (N_26588,N_19394,N_19996);
or U26589 (N_26589,N_18070,N_19438);
nor U26590 (N_26590,N_20882,N_21909);
or U26591 (N_26591,N_20561,N_22672);
nand U26592 (N_26592,N_22862,N_22671);
xor U26593 (N_26593,N_21953,N_19897);
xor U26594 (N_26594,N_23799,N_23538);
nand U26595 (N_26595,N_21225,N_23215);
and U26596 (N_26596,N_20111,N_19349);
xor U26597 (N_26597,N_22750,N_20986);
nor U26598 (N_26598,N_19184,N_21085);
or U26599 (N_26599,N_21006,N_21320);
or U26600 (N_26600,N_22032,N_20064);
and U26601 (N_26601,N_19065,N_20847);
nor U26602 (N_26602,N_20196,N_18221);
nand U26603 (N_26603,N_20782,N_19902);
nor U26604 (N_26604,N_21380,N_22327);
and U26605 (N_26605,N_22530,N_23825);
or U26606 (N_26606,N_21269,N_21859);
nor U26607 (N_26607,N_20422,N_22199);
nor U26608 (N_26608,N_21318,N_18359);
nand U26609 (N_26609,N_22565,N_21750);
nor U26610 (N_26610,N_20200,N_19652);
nand U26611 (N_26611,N_22799,N_20128);
nand U26612 (N_26612,N_18592,N_18989);
xnor U26613 (N_26613,N_21111,N_22848);
nand U26614 (N_26614,N_20413,N_19075);
nand U26615 (N_26615,N_19289,N_19642);
or U26616 (N_26616,N_18713,N_21172);
xnor U26617 (N_26617,N_22165,N_23864);
or U26618 (N_26618,N_22863,N_21021);
xnor U26619 (N_26619,N_18754,N_23323);
nor U26620 (N_26620,N_20016,N_22868);
xor U26621 (N_26621,N_23138,N_23218);
or U26622 (N_26622,N_18398,N_21463);
xnor U26623 (N_26623,N_21543,N_21334);
nand U26624 (N_26624,N_18943,N_20147);
nor U26625 (N_26625,N_18778,N_22305);
xor U26626 (N_26626,N_23767,N_18462);
nand U26627 (N_26627,N_20584,N_21862);
nand U26628 (N_26628,N_21569,N_22352);
and U26629 (N_26629,N_23441,N_23674);
or U26630 (N_26630,N_22727,N_19482);
xor U26631 (N_26631,N_19170,N_21890);
nor U26632 (N_26632,N_19579,N_20997);
xor U26633 (N_26633,N_23471,N_22542);
nand U26634 (N_26634,N_20169,N_22850);
nor U26635 (N_26635,N_21668,N_20625);
and U26636 (N_26636,N_23411,N_20513);
nor U26637 (N_26637,N_20471,N_20164);
xor U26638 (N_26638,N_20436,N_20519);
xor U26639 (N_26639,N_18739,N_23868);
nand U26640 (N_26640,N_22134,N_22107);
nor U26641 (N_26641,N_20226,N_21080);
and U26642 (N_26642,N_21168,N_22096);
xnor U26643 (N_26643,N_21254,N_20793);
or U26644 (N_26644,N_21840,N_20287);
or U26645 (N_26645,N_20293,N_23905);
or U26646 (N_26646,N_23096,N_19991);
nor U26647 (N_26647,N_18958,N_21818);
nor U26648 (N_26648,N_20297,N_18453);
or U26649 (N_26649,N_21943,N_20574);
or U26650 (N_26650,N_19292,N_21733);
xor U26651 (N_26651,N_21149,N_21754);
nor U26652 (N_26652,N_18934,N_18240);
nand U26653 (N_26653,N_18728,N_20776);
or U26654 (N_26654,N_20968,N_21938);
nor U26655 (N_26655,N_21246,N_20056);
nand U26656 (N_26656,N_23676,N_20696);
and U26657 (N_26657,N_20278,N_19105);
or U26658 (N_26658,N_22197,N_18110);
nand U26659 (N_26659,N_22513,N_19863);
or U26660 (N_26660,N_21829,N_18505);
or U26661 (N_26661,N_23697,N_21662);
nand U26662 (N_26662,N_23589,N_18199);
nor U26663 (N_26663,N_22845,N_21934);
xnor U26664 (N_26664,N_20912,N_19109);
or U26665 (N_26665,N_21516,N_21971);
and U26666 (N_26666,N_22300,N_21915);
xnor U26667 (N_26667,N_21018,N_23244);
nand U26668 (N_26668,N_21985,N_23148);
or U26669 (N_26669,N_21811,N_19336);
and U26670 (N_26670,N_20307,N_19591);
nand U26671 (N_26671,N_22495,N_19660);
nand U26672 (N_26672,N_23500,N_22093);
nor U26673 (N_26673,N_22821,N_19135);
nand U26674 (N_26674,N_18951,N_18675);
nand U26675 (N_26675,N_18990,N_21711);
or U26676 (N_26676,N_20800,N_20151);
nor U26677 (N_26677,N_23045,N_23744);
and U26678 (N_26678,N_19848,N_19119);
nor U26679 (N_26679,N_22159,N_20011);
or U26680 (N_26680,N_21910,N_22215);
nand U26681 (N_26681,N_19973,N_19793);
or U26682 (N_26682,N_19899,N_22592);
or U26683 (N_26683,N_21322,N_18489);
nor U26684 (N_26684,N_23806,N_22363);
nor U26685 (N_26685,N_22206,N_23417);
nor U26686 (N_26686,N_20775,N_23020);
xnor U26687 (N_26687,N_23070,N_18077);
and U26688 (N_26688,N_20165,N_22282);
nor U26689 (N_26689,N_19329,N_20083);
or U26690 (N_26690,N_20819,N_18175);
nand U26691 (N_26691,N_21007,N_19807);
nand U26692 (N_26692,N_18660,N_21370);
and U26693 (N_26693,N_22690,N_22337);
nor U26694 (N_26694,N_18086,N_20433);
nand U26695 (N_26695,N_19682,N_18936);
xnor U26696 (N_26696,N_20359,N_20765);
xor U26697 (N_26697,N_18198,N_22898);
xnor U26698 (N_26698,N_19092,N_21749);
xnor U26699 (N_26699,N_20288,N_21492);
nand U26700 (N_26700,N_21073,N_22625);
nand U26701 (N_26701,N_20314,N_21597);
nand U26702 (N_26702,N_21449,N_18358);
nor U26703 (N_26703,N_23262,N_22291);
nand U26704 (N_26704,N_18702,N_23010);
or U26705 (N_26705,N_21564,N_23757);
and U26706 (N_26706,N_19489,N_19612);
xor U26707 (N_26707,N_21401,N_22171);
nand U26708 (N_26708,N_21626,N_22562);
or U26709 (N_26709,N_21731,N_19420);
nor U26710 (N_26710,N_18855,N_22244);
and U26711 (N_26711,N_21708,N_21550);
or U26712 (N_26712,N_21984,N_23297);
or U26713 (N_26713,N_20855,N_19136);
nor U26714 (N_26714,N_23507,N_21404);
and U26715 (N_26715,N_19190,N_20238);
or U26716 (N_26716,N_22369,N_22954);
xnor U26717 (N_26717,N_22875,N_21231);
nand U26718 (N_26718,N_18377,N_20619);
nor U26719 (N_26719,N_22554,N_20861);
xor U26720 (N_26720,N_23723,N_22033);
xnor U26721 (N_26721,N_19003,N_22871);
xnor U26722 (N_26722,N_19478,N_19677);
and U26723 (N_26723,N_21396,N_18914);
xnor U26724 (N_26724,N_18244,N_18204);
or U26725 (N_26725,N_20138,N_20168);
xor U26726 (N_26726,N_23917,N_23346);
nor U26727 (N_26727,N_18006,N_22760);
and U26728 (N_26728,N_21614,N_23440);
nor U26729 (N_26729,N_21000,N_18824);
nand U26730 (N_26730,N_19851,N_22116);
nand U26731 (N_26731,N_22984,N_23399);
and U26732 (N_26732,N_19757,N_19782);
or U26733 (N_26733,N_21256,N_19999);
nor U26734 (N_26734,N_20965,N_21186);
xor U26735 (N_26735,N_20040,N_19042);
xnor U26736 (N_26736,N_23156,N_21046);
xnor U26737 (N_26737,N_23895,N_20791);
xor U26738 (N_26738,N_20353,N_22858);
xnor U26739 (N_26739,N_21116,N_20078);
nand U26740 (N_26740,N_20853,N_23192);
nor U26741 (N_26741,N_19779,N_22115);
nor U26742 (N_26742,N_18428,N_20573);
nor U26743 (N_26743,N_22443,N_19004);
or U26744 (N_26744,N_19386,N_23955);
and U26745 (N_26745,N_21836,N_20914);
xor U26746 (N_26746,N_23191,N_21465);
xnor U26747 (N_26747,N_22777,N_18169);
xnor U26748 (N_26748,N_23854,N_18127);
xnor U26749 (N_26749,N_19921,N_23751);
nand U26750 (N_26750,N_20115,N_18040);
nand U26751 (N_26751,N_18561,N_23834);
or U26752 (N_26752,N_18838,N_19525);
and U26753 (N_26753,N_21784,N_19937);
xnor U26754 (N_26754,N_19249,N_22447);
nand U26755 (N_26755,N_22540,N_19139);
nor U26756 (N_26756,N_22278,N_18834);
or U26757 (N_26757,N_21842,N_22342);
xnor U26758 (N_26758,N_21473,N_20836);
and U26759 (N_26759,N_19998,N_22391);
or U26760 (N_26760,N_23550,N_23149);
or U26761 (N_26761,N_21854,N_18156);
and U26762 (N_26762,N_23990,N_20137);
nand U26763 (N_26763,N_18143,N_20794);
nor U26764 (N_26764,N_18573,N_23473);
nor U26765 (N_26765,N_21643,N_21410);
xnor U26766 (N_26766,N_20298,N_19089);
or U26767 (N_26767,N_21950,N_23184);
nand U26768 (N_26768,N_19714,N_20927);
nor U26769 (N_26769,N_23783,N_23258);
or U26770 (N_26770,N_23365,N_19260);
or U26771 (N_26771,N_19940,N_21625);
nor U26772 (N_26772,N_20822,N_20740);
or U26773 (N_26773,N_20096,N_19639);
and U26774 (N_26774,N_19980,N_19247);
nor U26775 (N_26775,N_18619,N_23223);
or U26776 (N_26776,N_18904,N_20202);
or U26777 (N_26777,N_19953,N_21437);
or U26778 (N_26778,N_19091,N_20322);
and U26779 (N_26779,N_22732,N_22350);
xor U26780 (N_26780,N_20871,N_23781);
nand U26781 (N_26781,N_21728,N_18057);
xnor U26782 (N_26782,N_21204,N_20449);
and U26783 (N_26783,N_18575,N_23327);
xor U26784 (N_26784,N_18027,N_19545);
xor U26785 (N_26785,N_22281,N_21567);
nor U26786 (N_26786,N_20532,N_23243);
nor U26787 (N_26787,N_18177,N_20459);
xor U26788 (N_26788,N_19104,N_18190);
or U26789 (N_26789,N_22884,N_23419);
nand U26790 (N_26790,N_21484,N_19053);
nand U26791 (N_26791,N_18536,N_21783);
and U26792 (N_26792,N_21011,N_23082);
nor U26793 (N_26793,N_21171,N_22541);
and U26794 (N_26794,N_23978,N_19838);
and U26795 (N_26795,N_23614,N_19565);
or U26796 (N_26796,N_21721,N_18547);
nand U26797 (N_26797,N_22930,N_18952);
nor U26798 (N_26798,N_18883,N_20533);
xor U26799 (N_26799,N_22048,N_23842);
nand U26800 (N_26800,N_18801,N_21926);
nand U26801 (N_26801,N_22811,N_21340);
nand U26802 (N_26802,N_18313,N_21355);
and U26803 (N_26803,N_19601,N_23596);
xnor U26804 (N_26804,N_18657,N_21381);
nor U26805 (N_26805,N_23694,N_18503);
xor U26806 (N_26806,N_23867,N_20752);
nand U26807 (N_26807,N_20467,N_23934);
or U26808 (N_26808,N_18839,N_18030);
nand U26809 (N_26809,N_18577,N_19453);
nand U26810 (N_26810,N_18374,N_20572);
or U26811 (N_26811,N_18321,N_19038);
or U26812 (N_26812,N_22640,N_21638);
or U26813 (N_26813,N_22113,N_19788);
nand U26814 (N_26814,N_23661,N_19325);
xnor U26815 (N_26815,N_21615,N_21002);
nand U26816 (N_26816,N_18789,N_22155);
and U26817 (N_26817,N_23724,N_21282);
nor U26818 (N_26818,N_20813,N_18800);
nand U26819 (N_26819,N_22122,N_20180);
or U26820 (N_26820,N_18394,N_22434);
nand U26821 (N_26821,N_20028,N_21472);
and U26822 (N_26822,N_20694,N_21843);
and U26823 (N_26823,N_23780,N_18546);
nor U26824 (N_26824,N_22212,N_23871);
nand U26825 (N_26825,N_18602,N_19873);
nand U26826 (N_26826,N_20850,N_19629);
nor U26827 (N_26827,N_18820,N_23137);
or U26828 (N_26828,N_21500,N_21553);
or U26829 (N_26829,N_21929,N_18450);
nand U26830 (N_26830,N_20904,N_21596);
nor U26831 (N_26831,N_18823,N_19938);
xnor U26832 (N_26832,N_20518,N_20339);
nand U26833 (N_26833,N_20254,N_22743);
nand U26834 (N_26834,N_18137,N_22216);
nor U26835 (N_26835,N_22638,N_22307);
nand U26836 (N_26836,N_19611,N_23527);
xor U26837 (N_26837,N_19974,N_23888);
nand U26838 (N_26838,N_23025,N_23505);
or U26839 (N_26839,N_22078,N_21889);
nor U26840 (N_26840,N_21780,N_19785);
nor U26841 (N_26841,N_20767,N_19814);
or U26842 (N_26842,N_19368,N_19250);
and U26843 (N_26843,N_18821,N_20897);
xor U26844 (N_26844,N_19221,N_23162);
nor U26845 (N_26845,N_20888,N_19228);
and U26846 (N_26846,N_18436,N_20896);
nand U26847 (N_26847,N_23282,N_23142);
or U26848 (N_26848,N_20780,N_23963);
nand U26849 (N_26849,N_18241,N_20435);
and U26850 (N_26850,N_20627,N_23700);
xor U26851 (N_26851,N_20842,N_22660);
xor U26852 (N_26852,N_21846,N_22289);
nor U26853 (N_26853,N_19101,N_19933);
and U26854 (N_26854,N_23988,N_18178);
xor U26855 (N_26855,N_18699,N_20247);
xnor U26856 (N_26856,N_18520,N_22125);
nand U26857 (N_26857,N_22966,N_22658);
and U26858 (N_26858,N_22987,N_23627);
nor U26859 (N_26859,N_23198,N_19315);
and U26860 (N_26860,N_23485,N_22741);
and U26861 (N_26861,N_18228,N_20296);
nand U26862 (N_26862,N_21427,N_22603);
nand U26863 (N_26863,N_19693,N_20832);
nand U26864 (N_26864,N_20789,N_21663);
xnor U26865 (N_26865,N_18050,N_23620);
or U26866 (N_26866,N_23995,N_22522);
nor U26867 (N_26867,N_19460,N_19981);
nor U26868 (N_26868,N_20260,N_18344);
or U26869 (N_26869,N_19415,N_19718);
or U26870 (N_26870,N_20538,N_20463);
nor U26871 (N_26871,N_20553,N_23843);
nor U26872 (N_26872,N_22612,N_19527);
nor U26873 (N_26873,N_21298,N_22164);
and U26874 (N_26874,N_20465,N_20982);
or U26875 (N_26875,N_23765,N_22220);
xnor U26876 (N_26876,N_18187,N_22263);
xnor U26877 (N_26877,N_23607,N_19167);
xor U26878 (N_26878,N_19194,N_21848);
nand U26879 (N_26879,N_21630,N_20643);
and U26880 (N_26880,N_21096,N_18457);
nor U26881 (N_26881,N_18346,N_18548);
and U26882 (N_26882,N_21312,N_21810);
or U26883 (N_26883,N_22394,N_19654);
xor U26884 (N_26884,N_19774,N_20905);
nand U26885 (N_26885,N_18788,N_22803);
or U26886 (N_26886,N_22986,N_21974);
nor U26887 (N_26887,N_23769,N_21669);
or U26888 (N_26888,N_22129,N_21311);
and U26889 (N_26889,N_19821,N_18173);
nor U26890 (N_26890,N_22271,N_23619);
nand U26891 (N_26891,N_19878,N_21819);
nand U26892 (N_26892,N_22990,N_22476);
nor U26893 (N_26893,N_21689,N_19159);
or U26894 (N_26894,N_21220,N_22172);
and U26895 (N_26895,N_20590,N_22722);
and U26896 (N_26896,N_23562,N_23748);
xnor U26897 (N_26897,N_19215,N_18172);
nor U26898 (N_26898,N_20753,N_18916);
xor U26899 (N_26899,N_21051,N_21160);
or U26900 (N_26900,N_21133,N_21418);
or U26901 (N_26901,N_22901,N_20964);
and U26902 (N_26902,N_22584,N_18563);
and U26903 (N_26903,N_23725,N_18924);
xnor U26904 (N_26904,N_18895,N_19414);
xor U26905 (N_26905,N_21005,N_19321);
nor U26906 (N_26906,N_18196,N_19808);
and U26907 (N_26907,N_20764,N_18385);
nand U26908 (N_26908,N_23731,N_22325);
nand U26909 (N_26909,N_23501,N_19203);
nand U26910 (N_26910,N_22704,N_18965);
nand U26911 (N_26911,N_19914,N_23186);
nor U26912 (N_26912,N_18604,N_21119);
and U26913 (N_26913,N_20859,N_18676);
xnor U26914 (N_26914,N_23498,N_23954);
nand U26915 (N_26915,N_18348,N_20230);
nand U26916 (N_26916,N_21416,N_23416);
nand U26917 (N_26917,N_23014,N_19819);
and U26918 (N_26918,N_18941,N_21959);
xnor U26919 (N_26919,N_23234,N_22211);
or U26920 (N_26920,N_22564,N_19282);
or U26921 (N_26921,N_19889,N_19298);
and U26922 (N_26922,N_22368,N_22882);
and U26923 (N_26923,N_22980,N_19051);
nand U26924 (N_26924,N_23972,N_23422);
xnor U26925 (N_26925,N_19979,N_20955);
nand U26926 (N_26926,N_19651,N_22849);
nor U26927 (N_26927,N_21554,N_22925);
and U26928 (N_26928,N_19183,N_18730);
nand U26929 (N_26929,N_18585,N_21823);
nor U26930 (N_26930,N_19743,N_18435);
xor U26931 (N_26931,N_18826,N_20323);
xnor U26932 (N_26932,N_18534,N_19372);
and U26933 (N_26933,N_23200,N_22985);
nand U26934 (N_26934,N_22711,N_23648);
nand U26935 (N_26935,N_23553,N_22407);
xor U26936 (N_26936,N_18856,N_22730);
xnor U26937 (N_26937,N_18011,N_23771);
xnor U26938 (N_26938,N_20667,N_21456);
or U26939 (N_26939,N_19306,N_21467);
or U26940 (N_26940,N_23971,N_19736);
xnor U26941 (N_26941,N_19465,N_21582);
nor U26942 (N_26942,N_19358,N_19920);
and U26943 (N_26943,N_22295,N_21693);
xor U26944 (N_26944,N_19879,N_22229);
xor U26945 (N_26945,N_18817,N_22726);
nor U26946 (N_26946,N_18016,N_20044);
nor U26947 (N_26947,N_19020,N_21993);
or U26948 (N_26948,N_22810,N_20420);
and U26949 (N_26949,N_22759,N_19936);
and U26950 (N_26950,N_21684,N_20874);
nor U26951 (N_26951,N_19724,N_20597);
or U26952 (N_26952,N_21847,N_23492);
nor U26953 (N_26953,N_19971,N_19064);
nand U26954 (N_26954,N_20531,N_18067);
xnor U26955 (N_26955,N_19388,N_22079);
or U26956 (N_26956,N_23330,N_18804);
xor U26957 (N_26957,N_19027,N_19544);
xor U26958 (N_26958,N_21776,N_20886);
xnor U26959 (N_26959,N_21301,N_21963);
or U26960 (N_26960,N_23472,N_21378);
nor U26961 (N_26961,N_23923,N_20027);
nor U26962 (N_26962,N_19125,N_18144);
nor U26963 (N_26963,N_21786,N_23394);
nor U26964 (N_26964,N_22601,N_22203);
nor U26965 (N_26965,N_18780,N_22738);
or U26966 (N_26966,N_23232,N_18084);
or U26967 (N_26967,N_21167,N_18189);
xnor U26968 (N_26968,N_18599,N_23611);
xor U26969 (N_26969,N_23426,N_19264);
nor U26970 (N_26970,N_20081,N_20095);
and U26971 (N_26971,N_20523,N_21178);
xnor U26972 (N_26972,N_20645,N_18612);
or U26973 (N_26973,N_22745,N_20431);
nand U26974 (N_26974,N_23129,N_23246);
and U26975 (N_26975,N_20124,N_21099);
or U26976 (N_26976,N_23261,N_22813);
xnor U26977 (N_26977,N_21952,N_19434);
nand U26978 (N_26978,N_19754,N_23208);
xor U26979 (N_26979,N_18218,N_21341);
nand U26980 (N_26980,N_22739,N_20374);
nand U26981 (N_26981,N_21788,N_23127);
or U26982 (N_26982,N_21429,N_22523);
and U26983 (N_26983,N_18544,N_22458);
and U26984 (N_26984,N_18411,N_22457);
nand U26985 (N_26985,N_21268,N_20710);
nand U26986 (N_26986,N_19732,N_19904);
xnor U26987 (N_26987,N_20013,N_19477);
nand U26988 (N_26988,N_19723,N_20887);
nand U26989 (N_26989,N_18484,N_23102);
xnor U26990 (N_26990,N_19997,N_19729);
nor U26991 (N_26991,N_19371,N_20462);
xor U26992 (N_26992,N_23060,N_21261);
nand U26993 (N_26993,N_22009,N_20958);
xnor U26994 (N_26994,N_21242,N_21386);
xnor U26995 (N_26995,N_22219,N_21438);
nor U26996 (N_26996,N_21190,N_23788);
xnor U26997 (N_26997,N_20917,N_22593);
nand U26998 (N_26998,N_20612,N_21545);
nor U26999 (N_26999,N_20479,N_21999);
xnor U27000 (N_27000,N_20276,N_21753);
nand U27001 (N_27001,N_21274,N_19511);
nor U27002 (N_27002,N_23149,N_21384);
nand U27003 (N_27003,N_22936,N_23204);
and U27004 (N_27004,N_21382,N_18087);
nor U27005 (N_27005,N_18511,N_22524);
xor U27006 (N_27006,N_21985,N_22938);
and U27007 (N_27007,N_19630,N_18253);
nand U27008 (N_27008,N_21840,N_18095);
xnor U27009 (N_27009,N_19200,N_19887);
nor U27010 (N_27010,N_20910,N_21759);
nor U27011 (N_27011,N_23847,N_21063);
xor U27012 (N_27012,N_23538,N_21830);
xnor U27013 (N_27013,N_18190,N_18436);
or U27014 (N_27014,N_19515,N_22078);
xor U27015 (N_27015,N_22737,N_18013);
or U27016 (N_27016,N_19396,N_22441);
and U27017 (N_27017,N_23328,N_19852);
and U27018 (N_27018,N_18290,N_23942);
nand U27019 (N_27019,N_22516,N_19637);
xnor U27020 (N_27020,N_22924,N_20047);
nand U27021 (N_27021,N_20565,N_21464);
or U27022 (N_27022,N_20198,N_20615);
or U27023 (N_27023,N_18061,N_18259);
nor U27024 (N_27024,N_22227,N_23612);
nand U27025 (N_27025,N_23705,N_20678);
nor U27026 (N_27026,N_18725,N_22679);
and U27027 (N_27027,N_19100,N_20882);
xnor U27028 (N_27028,N_18143,N_23904);
or U27029 (N_27029,N_19695,N_18949);
xnor U27030 (N_27030,N_18187,N_18957);
xnor U27031 (N_27031,N_23993,N_18693);
nand U27032 (N_27032,N_20859,N_23692);
xor U27033 (N_27033,N_20020,N_22247);
nor U27034 (N_27034,N_20347,N_20176);
and U27035 (N_27035,N_22366,N_20739);
nor U27036 (N_27036,N_22845,N_19531);
xnor U27037 (N_27037,N_21886,N_23892);
and U27038 (N_27038,N_19818,N_18802);
or U27039 (N_27039,N_21508,N_18607);
xnor U27040 (N_27040,N_19412,N_23886);
xnor U27041 (N_27041,N_20325,N_20323);
xnor U27042 (N_27042,N_21766,N_23900);
nor U27043 (N_27043,N_18919,N_23716);
nor U27044 (N_27044,N_19676,N_20299);
nor U27045 (N_27045,N_21450,N_21451);
and U27046 (N_27046,N_19408,N_23004);
or U27047 (N_27047,N_18973,N_19826);
or U27048 (N_27048,N_18011,N_20362);
and U27049 (N_27049,N_19695,N_23558);
or U27050 (N_27050,N_20267,N_23091);
nor U27051 (N_27051,N_19146,N_21234);
and U27052 (N_27052,N_21785,N_21960);
nand U27053 (N_27053,N_19108,N_21731);
or U27054 (N_27054,N_19429,N_18437);
and U27055 (N_27055,N_21906,N_22011);
nor U27056 (N_27056,N_21430,N_22880);
xnor U27057 (N_27057,N_21023,N_18229);
and U27058 (N_27058,N_18383,N_22638);
or U27059 (N_27059,N_20988,N_21333);
xnor U27060 (N_27060,N_20748,N_19186);
and U27061 (N_27061,N_21931,N_22993);
xor U27062 (N_27062,N_23868,N_20578);
nor U27063 (N_27063,N_21527,N_20775);
or U27064 (N_27064,N_20872,N_22911);
nor U27065 (N_27065,N_20897,N_20983);
xor U27066 (N_27066,N_23019,N_19526);
or U27067 (N_27067,N_23359,N_18727);
and U27068 (N_27068,N_22443,N_23077);
and U27069 (N_27069,N_20756,N_22274);
xor U27070 (N_27070,N_19825,N_20154);
xnor U27071 (N_27071,N_19536,N_18341);
or U27072 (N_27072,N_20655,N_22854);
or U27073 (N_27073,N_20672,N_18626);
nor U27074 (N_27074,N_19925,N_23883);
and U27075 (N_27075,N_20435,N_20580);
or U27076 (N_27076,N_20416,N_23402);
nand U27077 (N_27077,N_20274,N_20768);
or U27078 (N_27078,N_23535,N_22334);
nor U27079 (N_27079,N_20189,N_20950);
or U27080 (N_27080,N_21739,N_18520);
nand U27081 (N_27081,N_22986,N_23353);
nand U27082 (N_27082,N_23826,N_18032);
and U27083 (N_27083,N_23329,N_23128);
nand U27084 (N_27084,N_23930,N_20189);
xor U27085 (N_27085,N_23369,N_20435);
or U27086 (N_27086,N_21334,N_23982);
or U27087 (N_27087,N_23265,N_22586);
or U27088 (N_27088,N_21525,N_21541);
and U27089 (N_27089,N_19543,N_23283);
nor U27090 (N_27090,N_18811,N_18847);
nand U27091 (N_27091,N_19112,N_23097);
and U27092 (N_27092,N_20591,N_19293);
xnor U27093 (N_27093,N_23824,N_23734);
and U27094 (N_27094,N_21671,N_20835);
xnor U27095 (N_27095,N_18976,N_21629);
and U27096 (N_27096,N_23532,N_18204);
and U27097 (N_27097,N_18792,N_20096);
nor U27098 (N_27098,N_18514,N_23065);
nor U27099 (N_27099,N_19218,N_18567);
nand U27100 (N_27100,N_19908,N_23582);
nand U27101 (N_27101,N_22816,N_19606);
nor U27102 (N_27102,N_21363,N_19030);
nand U27103 (N_27103,N_21125,N_18819);
nand U27104 (N_27104,N_23259,N_18343);
and U27105 (N_27105,N_22672,N_19719);
nor U27106 (N_27106,N_22345,N_21656);
nand U27107 (N_27107,N_18822,N_19635);
xnor U27108 (N_27108,N_21140,N_21792);
xnor U27109 (N_27109,N_19962,N_23993);
or U27110 (N_27110,N_19215,N_22374);
nand U27111 (N_27111,N_19446,N_20648);
or U27112 (N_27112,N_18123,N_18781);
or U27113 (N_27113,N_19232,N_20734);
xor U27114 (N_27114,N_22638,N_19138);
nor U27115 (N_27115,N_18742,N_21597);
nor U27116 (N_27116,N_18294,N_20664);
xnor U27117 (N_27117,N_19277,N_21872);
xnor U27118 (N_27118,N_23479,N_23176);
and U27119 (N_27119,N_20147,N_23187);
nor U27120 (N_27120,N_20041,N_22731);
nand U27121 (N_27121,N_20106,N_19762);
nor U27122 (N_27122,N_18719,N_19990);
nand U27123 (N_27123,N_19709,N_20855);
or U27124 (N_27124,N_22651,N_21646);
nor U27125 (N_27125,N_19476,N_23482);
or U27126 (N_27126,N_20033,N_23026);
nor U27127 (N_27127,N_19404,N_22204);
and U27128 (N_27128,N_21271,N_20824);
or U27129 (N_27129,N_18076,N_19761);
or U27130 (N_27130,N_18873,N_22554);
nand U27131 (N_27131,N_19812,N_23038);
and U27132 (N_27132,N_20923,N_23819);
nor U27133 (N_27133,N_18431,N_22861);
or U27134 (N_27134,N_20055,N_21964);
and U27135 (N_27135,N_23980,N_23693);
nand U27136 (N_27136,N_23208,N_23160);
xor U27137 (N_27137,N_22716,N_19837);
nand U27138 (N_27138,N_21764,N_19696);
nand U27139 (N_27139,N_20909,N_23787);
nor U27140 (N_27140,N_19981,N_21203);
nor U27141 (N_27141,N_19105,N_21273);
xnor U27142 (N_27142,N_18744,N_21446);
nand U27143 (N_27143,N_21358,N_22456);
xor U27144 (N_27144,N_20559,N_18034);
nand U27145 (N_27145,N_23284,N_18439);
or U27146 (N_27146,N_23816,N_18819);
xor U27147 (N_27147,N_19727,N_23498);
xor U27148 (N_27148,N_18844,N_20133);
or U27149 (N_27149,N_20869,N_21146);
nand U27150 (N_27150,N_23691,N_20511);
nor U27151 (N_27151,N_22432,N_18414);
and U27152 (N_27152,N_19884,N_22569);
nand U27153 (N_27153,N_19743,N_21287);
nand U27154 (N_27154,N_22799,N_23516);
nand U27155 (N_27155,N_23033,N_19302);
xnor U27156 (N_27156,N_18054,N_22100);
nand U27157 (N_27157,N_19907,N_23587);
nand U27158 (N_27158,N_18069,N_20165);
nand U27159 (N_27159,N_22373,N_21453);
or U27160 (N_27160,N_19881,N_20842);
nand U27161 (N_27161,N_18503,N_18486);
and U27162 (N_27162,N_22555,N_20144);
nor U27163 (N_27163,N_18421,N_21355);
xnor U27164 (N_27164,N_21015,N_22317);
and U27165 (N_27165,N_21169,N_22104);
or U27166 (N_27166,N_19421,N_21300);
xnor U27167 (N_27167,N_20252,N_21124);
nand U27168 (N_27168,N_23158,N_23604);
nand U27169 (N_27169,N_18859,N_21679);
and U27170 (N_27170,N_23875,N_20430);
and U27171 (N_27171,N_19863,N_22043);
and U27172 (N_27172,N_23939,N_20932);
nor U27173 (N_27173,N_18661,N_20433);
nand U27174 (N_27174,N_23256,N_22249);
xnor U27175 (N_27175,N_20634,N_22744);
or U27176 (N_27176,N_20126,N_21542);
and U27177 (N_27177,N_22677,N_19450);
nor U27178 (N_27178,N_18262,N_18560);
or U27179 (N_27179,N_18136,N_21989);
and U27180 (N_27180,N_18620,N_23273);
nor U27181 (N_27181,N_21043,N_23431);
nand U27182 (N_27182,N_21013,N_19601);
or U27183 (N_27183,N_22422,N_21469);
or U27184 (N_27184,N_19062,N_22156);
nor U27185 (N_27185,N_20877,N_23447);
or U27186 (N_27186,N_22955,N_18530);
or U27187 (N_27187,N_23210,N_21653);
or U27188 (N_27188,N_20061,N_22118);
nand U27189 (N_27189,N_22201,N_23108);
nor U27190 (N_27190,N_20260,N_21869);
nor U27191 (N_27191,N_21201,N_19119);
xor U27192 (N_27192,N_19815,N_18165);
nand U27193 (N_27193,N_23717,N_23195);
nor U27194 (N_27194,N_23969,N_23078);
xor U27195 (N_27195,N_19905,N_23380);
or U27196 (N_27196,N_23183,N_22601);
or U27197 (N_27197,N_22633,N_18434);
and U27198 (N_27198,N_23286,N_18854);
and U27199 (N_27199,N_23585,N_20619);
nand U27200 (N_27200,N_23280,N_21577);
nand U27201 (N_27201,N_22031,N_22521);
nor U27202 (N_27202,N_22593,N_23633);
xnor U27203 (N_27203,N_23057,N_18403);
nand U27204 (N_27204,N_23608,N_21189);
xnor U27205 (N_27205,N_22157,N_23385);
xnor U27206 (N_27206,N_18260,N_20175);
and U27207 (N_27207,N_20662,N_21387);
and U27208 (N_27208,N_21122,N_22407);
nor U27209 (N_27209,N_18937,N_23109);
xor U27210 (N_27210,N_20564,N_21829);
and U27211 (N_27211,N_22100,N_23678);
xnor U27212 (N_27212,N_18757,N_21752);
nor U27213 (N_27213,N_21933,N_18155);
xnor U27214 (N_27214,N_22830,N_18042);
nor U27215 (N_27215,N_20516,N_23455);
xor U27216 (N_27216,N_18197,N_20963);
and U27217 (N_27217,N_18916,N_19963);
nand U27218 (N_27218,N_20767,N_23487);
and U27219 (N_27219,N_18315,N_20383);
nor U27220 (N_27220,N_23630,N_19014);
nand U27221 (N_27221,N_20642,N_21983);
xor U27222 (N_27222,N_23217,N_19458);
nand U27223 (N_27223,N_21422,N_20156);
nand U27224 (N_27224,N_19099,N_20902);
xnor U27225 (N_27225,N_22933,N_21322);
nand U27226 (N_27226,N_22097,N_22144);
and U27227 (N_27227,N_20977,N_21543);
nand U27228 (N_27228,N_20506,N_18399);
and U27229 (N_27229,N_22406,N_18199);
nand U27230 (N_27230,N_22992,N_19524);
xnor U27231 (N_27231,N_22119,N_21346);
xor U27232 (N_27232,N_21080,N_19979);
nor U27233 (N_27233,N_21456,N_18269);
nand U27234 (N_27234,N_21257,N_18986);
and U27235 (N_27235,N_21613,N_22834);
and U27236 (N_27236,N_18942,N_23876);
nand U27237 (N_27237,N_21142,N_20230);
xor U27238 (N_27238,N_19998,N_23378);
xor U27239 (N_27239,N_21391,N_23428);
xnor U27240 (N_27240,N_18852,N_18923);
and U27241 (N_27241,N_22627,N_19058);
nor U27242 (N_27242,N_19554,N_19730);
nor U27243 (N_27243,N_22098,N_23815);
nand U27244 (N_27244,N_20523,N_20281);
and U27245 (N_27245,N_22127,N_23484);
nand U27246 (N_27246,N_19940,N_21183);
or U27247 (N_27247,N_18667,N_19107);
nor U27248 (N_27248,N_19701,N_19729);
xor U27249 (N_27249,N_20282,N_22716);
nor U27250 (N_27250,N_23860,N_18620);
and U27251 (N_27251,N_21917,N_21118);
nor U27252 (N_27252,N_21287,N_19223);
and U27253 (N_27253,N_18496,N_23903);
nor U27254 (N_27254,N_20322,N_23787);
or U27255 (N_27255,N_21177,N_21684);
xnor U27256 (N_27256,N_21658,N_22964);
xnor U27257 (N_27257,N_19612,N_20218);
or U27258 (N_27258,N_23670,N_20732);
nand U27259 (N_27259,N_23155,N_23799);
and U27260 (N_27260,N_19236,N_21404);
nand U27261 (N_27261,N_22870,N_21477);
nand U27262 (N_27262,N_23068,N_19949);
or U27263 (N_27263,N_22981,N_22611);
nand U27264 (N_27264,N_20978,N_21577);
or U27265 (N_27265,N_18789,N_20583);
and U27266 (N_27266,N_23187,N_18950);
and U27267 (N_27267,N_20639,N_21248);
nand U27268 (N_27268,N_22493,N_22034);
xnor U27269 (N_27269,N_20194,N_18721);
and U27270 (N_27270,N_18301,N_18165);
xor U27271 (N_27271,N_21783,N_19786);
nand U27272 (N_27272,N_19937,N_22368);
nand U27273 (N_27273,N_22334,N_21907);
nand U27274 (N_27274,N_22623,N_22950);
nand U27275 (N_27275,N_20861,N_20367);
or U27276 (N_27276,N_20774,N_20182);
xnor U27277 (N_27277,N_21925,N_18791);
nand U27278 (N_27278,N_21393,N_19035);
or U27279 (N_27279,N_21733,N_23868);
and U27280 (N_27280,N_23732,N_18994);
nand U27281 (N_27281,N_23253,N_22032);
and U27282 (N_27282,N_18488,N_20258);
nand U27283 (N_27283,N_19580,N_22428);
or U27284 (N_27284,N_21571,N_18788);
or U27285 (N_27285,N_22269,N_19895);
or U27286 (N_27286,N_19713,N_22495);
xor U27287 (N_27287,N_23188,N_22068);
xor U27288 (N_27288,N_20690,N_18933);
nor U27289 (N_27289,N_20886,N_19894);
nor U27290 (N_27290,N_22369,N_19058);
or U27291 (N_27291,N_19328,N_19079);
nor U27292 (N_27292,N_22265,N_21886);
xnor U27293 (N_27293,N_20432,N_23920);
or U27294 (N_27294,N_22677,N_19099);
xnor U27295 (N_27295,N_19190,N_19242);
and U27296 (N_27296,N_23326,N_21455);
or U27297 (N_27297,N_23057,N_18296);
and U27298 (N_27298,N_18452,N_19536);
nand U27299 (N_27299,N_19109,N_22324);
nand U27300 (N_27300,N_18364,N_20870);
or U27301 (N_27301,N_20457,N_20217);
xor U27302 (N_27302,N_18714,N_20119);
nand U27303 (N_27303,N_18425,N_21665);
or U27304 (N_27304,N_23224,N_18123);
xor U27305 (N_27305,N_18810,N_22667);
nand U27306 (N_27306,N_20448,N_23410);
and U27307 (N_27307,N_20257,N_18724);
nor U27308 (N_27308,N_22267,N_22701);
or U27309 (N_27309,N_21598,N_19855);
xor U27310 (N_27310,N_22846,N_19597);
xor U27311 (N_27311,N_19727,N_22609);
nor U27312 (N_27312,N_22910,N_18772);
or U27313 (N_27313,N_21299,N_22550);
and U27314 (N_27314,N_19081,N_23319);
nand U27315 (N_27315,N_22925,N_18587);
and U27316 (N_27316,N_22406,N_18717);
nor U27317 (N_27317,N_21967,N_23214);
nor U27318 (N_27318,N_18018,N_20260);
and U27319 (N_27319,N_22871,N_20478);
nor U27320 (N_27320,N_23919,N_21310);
nand U27321 (N_27321,N_19876,N_22379);
and U27322 (N_27322,N_19385,N_18743);
nand U27323 (N_27323,N_19133,N_18119);
or U27324 (N_27324,N_18317,N_21676);
nand U27325 (N_27325,N_18791,N_21534);
xnor U27326 (N_27326,N_20754,N_19156);
nor U27327 (N_27327,N_18366,N_20599);
nor U27328 (N_27328,N_19217,N_20804);
xor U27329 (N_27329,N_20803,N_21498);
and U27330 (N_27330,N_22844,N_19043);
and U27331 (N_27331,N_22143,N_20391);
nor U27332 (N_27332,N_21357,N_20546);
xor U27333 (N_27333,N_19849,N_22540);
nand U27334 (N_27334,N_19916,N_18948);
nand U27335 (N_27335,N_19517,N_21325);
and U27336 (N_27336,N_18692,N_18396);
and U27337 (N_27337,N_22315,N_19135);
xor U27338 (N_27338,N_19730,N_20498);
xor U27339 (N_27339,N_21353,N_23300);
nor U27340 (N_27340,N_20789,N_20796);
and U27341 (N_27341,N_21884,N_22506);
nor U27342 (N_27342,N_20997,N_22112);
nor U27343 (N_27343,N_18506,N_22361);
nand U27344 (N_27344,N_19569,N_23000);
and U27345 (N_27345,N_18126,N_21089);
or U27346 (N_27346,N_18157,N_22707);
and U27347 (N_27347,N_20814,N_19068);
xor U27348 (N_27348,N_23403,N_23595);
or U27349 (N_27349,N_18713,N_23792);
nand U27350 (N_27350,N_18543,N_19642);
xor U27351 (N_27351,N_19825,N_22837);
or U27352 (N_27352,N_18402,N_18386);
nand U27353 (N_27353,N_22612,N_21553);
or U27354 (N_27354,N_22616,N_19279);
and U27355 (N_27355,N_19126,N_21187);
xnor U27356 (N_27356,N_20142,N_19215);
nand U27357 (N_27357,N_23080,N_23397);
xnor U27358 (N_27358,N_22551,N_18001);
and U27359 (N_27359,N_19651,N_22878);
and U27360 (N_27360,N_23621,N_18628);
xor U27361 (N_27361,N_20685,N_18732);
nor U27362 (N_27362,N_19321,N_18885);
and U27363 (N_27363,N_22074,N_22587);
nand U27364 (N_27364,N_23301,N_20901);
nor U27365 (N_27365,N_20907,N_22160);
and U27366 (N_27366,N_20452,N_18512);
xnor U27367 (N_27367,N_18195,N_21438);
xor U27368 (N_27368,N_19272,N_21247);
nor U27369 (N_27369,N_21453,N_18422);
or U27370 (N_27370,N_18628,N_21583);
nand U27371 (N_27371,N_23878,N_21932);
xor U27372 (N_27372,N_21385,N_19696);
and U27373 (N_27373,N_21610,N_20963);
nand U27374 (N_27374,N_19073,N_20070);
nand U27375 (N_27375,N_19094,N_21776);
xnor U27376 (N_27376,N_20329,N_23677);
and U27377 (N_27377,N_19951,N_20232);
nor U27378 (N_27378,N_21916,N_18674);
nor U27379 (N_27379,N_22920,N_20516);
and U27380 (N_27380,N_19927,N_21822);
or U27381 (N_27381,N_21849,N_21156);
nor U27382 (N_27382,N_20029,N_20652);
nand U27383 (N_27383,N_23941,N_18474);
nor U27384 (N_27384,N_19530,N_21171);
xnor U27385 (N_27385,N_22009,N_19830);
and U27386 (N_27386,N_20369,N_19150);
or U27387 (N_27387,N_22810,N_21904);
nor U27388 (N_27388,N_20727,N_23950);
nor U27389 (N_27389,N_21323,N_18814);
xor U27390 (N_27390,N_23965,N_23611);
nor U27391 (N_27391,N_19214,N_23402);
xor U27392 (N_27392,N_22261,N_18978);
nor U27393 (N_27393,N_21026,N_19310);
or U27394 (N_27394,N_22925,N_19700);
nand U27395 (N_27395,N_18125,N_23908);
nor U27396 (N_27396,N_20871,N_22089);
xor U27397 (N_27397,N_18513,N_23883);
xnor U27398 (N_27398,N_20685,N_22764);
xor U27399 (N_27399,N_20241,N_18498);
xor U27400 (N_27400,N_19125,N_22448);
nor U27401 (N_27401,N_23581,N_23154);
xnor U27402 (N_27402,N_21147,N_21356);
or U27403 (N_27403,N_22130,N_23042);
nor U27404 (N_27404,N_19791,N_20641);
or U27405 (N_27405,N_19772,N_21679);
nand U27406 (N_27406,N_19812,N_18264);
and U27407 (N_27407,N_21387,N_19621);
or U27408 (N_27408,N_19483,N_23424);
nand U27409 (N_27409,N_23038,N_20708);
or U27410 (N_27410,N_19464,N_19997);
and U27411 (N_27411,N_20393,N_19974);
nand U27412 (N_27412,N_19368,N_19759);
xor U27413 (N_27413,N_19972,N_19931);
nand U27414 (N_27414,N_22395,N_18806);
xor U27415 (N_27415,N_21953,N_23971);
and U27416 (N_27416,N_22653,N_21153);
xnor U27417 (N_27417,N_18715,N_23111);
and U27418 (N_27418,N_18941,N_18751);
nand U27419 (N_27419,N_19643,N_19746);
nand U27420 (N_27420,N_20620,N_19196);
nand U27421 (N_27421,N_23332,N_18989);
xor U27422 (N_27422,N_22501,N_22174);
nor U27423 (N_27423,N_20824,N_18483);
nand U27424 (N_27424,N_23143,N_18537);
and U27425 (N_27425,N_21004,N_20551);
xnor U27426 (N_27426,N_20494,N_20209);
nand U27427 (N_27427,N_18402,N_19912);
nor U27428 (N_27428,N_23152,N_22630);
nor U27429 (N_27429,N_18431,N_18413);
nor U27430 (N_27430,N_20271,N_22836);
nand U27431 (N_27431,N_18121,N_19515);
xor U27432 (N_27432,N_20239,N_22222);
nor U27433 (N_27433,N_21796,N_18265);
nor U27434 (N_27434,N_21661,N_19181);
nor U27435 (N_27435,N_20933,N_22565);
xnor U27436 (N_27436,N_19396,N_20009);
xnor U27437 (N_27437,N_23131,N_19863);
or U27438 (N_27438,N_18522,N_20066);
and U27439 (N_27439,N_18679,N_18969);
and U27440 (N_27440,N_21513,N_23960);
nand U27441 (N_27441,N_20168,N_23572);
and U27442 (N_27442,N_21321,N_23691);
nand U27443 (N_27443,N_18667,N_19808);
and U27444 (N_27444,N_22338,N_23645);
nand U27445 (N_27445,N_21647,N_19601);
and U27446 (N_27446,N_23976,N_20216);
and U27447 (N_27447,N_19945,N_23597);
xor U27448 (N_27448,N_23268,N_20009);
or U27449 (N_27449,N_18933,N_19853);
and U27450 (N_27450,N_22795,N_20345);
nor U27451 (N_27451,N_23267,N_22443);
xor U27452 (N_27452,N_22289,N_18625);
nand U27453 (N_27453,N_23548,N_18179);
or U27454 (N_27454,N_23101,N_20523);
and U27455 (N_27455,N_19209,N_18614);
nor U27456 (N_27456,N_18705,N_23201);
xnor U27457 (N_27457,N_19945,N_20730);
xnor U27458 (N_27458,N_19249,N_19095);
and U27459 (N_27459,N_19689,N_22952);
or U27460 (N_27460,N_18981,N_22218);
nand U27461 (N_27461,N_21248,N_19044);
and U27462 (N_27462,N_20896,N_20836);
xor U27463 (N_27463,N_20448,N_22634);
nand U27464 (N_27464,N_18561,N_21095);
or U27465 (N_27465,N_22961,N_21289);
nor U27466 (N_27466,N_22003,N_18545);
or U27467 (N_27467,N_18826,N_18691);
nor U27468 (N_27468,N_23556,N_22987);
nor U27469 (N_27469,N_23925,N_23366);
xor U27470 (N_27470,N_19947,N_19139);
xnor U27471 (N_27471,N_19940,N_19282);
nand U27472 (N_27472,N_21636,N_20599);
nor U27473 (N_27473,N_21516,N_21167);
or U27474 (N_27474,N_19501,N_21208);
nor U27475 (N_27475,N_18040,N_19686);
xor U27476 (N_27476,N_22814,N_22594);
nand U27477 (N_27477,N_22426,N_20521);
xnor U27478 (N_27478,N_21811,N_23536);
xor U27479 (N_27479,N_20724,N_20638);
nor U27480 (N_27480,N_19262,N_21946);
xnor U27481 (N_27481,N_23936,N_20827);
and U27482 (N_27482,N_21140,N_19690);
xor U27483 (N_27483,N_19043,N_19659);
or U27484 (N_27484,N_19010,N_23286);
nand U27485 (N_27485,N_21918,N_23837);
nor U27486 (N_27486,N_20128,N_18966);
nor U27487 (N_27487,N_19213,N_22580);
and U27488 (N_27488,N_18634,N_18742);
nand U27489 (N_27489,N_21821,N_20792);
or U27490 (N_27490,N_23003,N_18111);
or U27491 (N_27491,N_18739,N_21119);
and U27492 (N_27492,N_20456,N_19000);
nand U27493 (N_27493,N_19992,N_23260);
or U27494 (N_27494,N_20351,N_20857);
and U27495 (N_27495,N_23082,N_18515);
xor U27496 (N_27496,N_19333,N_23702);
and U27497 (N_27497,N_22618,N_19679);
nor U27498 (N_27498,N_21485,N_23966);
nor U27499 (N_27499,N_22062,N_21933);
or U27500 (N_27500,N_18029,N_23682);
nand U27501 (N_27501,N_23578,N_18411);
nor U27502 (N_27502,N_22085,N_20519);
or U27503 (N_27503,N_23528,N_20880);
or U27504 (N_27504,N_18216,N_18522);
nor U27505 (N_27505,N_22062,N_18030);
xor U27506 (N_27506,N_23008,N_22334);
or U27507 (N_27507,N_21017,N_22661);
and U27508 (N_27508,N_23773,N_18320);
or U27509 (N_27509,N_22390,N_19957);
xnor U27510 (N_27510,N_23251,N_22011);
nand U27511 (N_27511,N_23864,N_21536);
and U27512 (N_27512,N_21660,N_19838);
xnor U27513 (N_27513,N_19975,N_21339);
and U27514 (N_27514,N_22919,N_22605);
or U27515 (N_27515,N_19837,N_21529);
xnor U27516 (N_27516,N_20764,N_18193);
xnor U27517 (N_27517,N_23942,N_18496);
and U27518 (N_27518,N_21226,N_19921);
nor U27519 (N_27519,N_19854,N_19731);
nand U27520 (N_27520,N_18750,N_20883);
or U27521 (N_27521,N_20478,N_20625);
xnor U27522 (N_27522,N_22154,N_18239);
nor U27523 (N_27523,N_23088,N_19107);
xnor U27524 (N_27524,N_19066,N_21159);
or U27525 (N_27525,N_19321,N_20721);
or U27526 (N_27526,N_23341,N_21325);
nor U27527 (N_27527,N_23343,N_22688);
or U27528 (N_27528,N_20622,N_23955);
nand U27529 (N_27529,N_20081,N_23404);
nor U27530 (N_27530,N_19468,N_21538);
or U27531 (N_27531,N_23053,N_19480);
nor U27532 (N_27532,N_20776,N_21367);
and U27533 (N_27533,N_23915,N_22023);
nor U27534 (N_27534,N_20145,N_23108);
xor U27535 (N_27535,N_20754,N_18978);
or U27536 (N_27536,N_19028,N_23707);
xnor U27537 (N_27537,N_19153,N_20652);
and U27538 (N_27538,N_22161,N_20459);
and U27539 (N_27539,N_22124,N_21317);
or U27540 (N_27540,N_21163,N_22502);
or U27541 (N_27541,N_23567,N_20987);
xor U27542 (N_27542,N_22726,N_19220);
nor U27543 (N_27543,N_23321,N_22674);
or U27544 (N_27544,N_22936,N_23855);
nand U27545 (N_27545,N_19396,N_18482);
and U27546 (N_27546,N_18782,N_21433);
and U27547 (N_27547,N_18460,N_19279);
nand U27548 (N_27548,N_20024,N_23531);
or U27549 (N_27549,N_19975,N_20051);
xor U27550 (N_27550,N_21241,N_21687);
or U27551 (N_27551,N_18815,N_18903);
or U27552 (N_27552,N_22454,N_18366);
xnor U27553 (N_27553,N_20741,N_19735);
xor U27554 (N_27554,N_23392,N_18791);
or U27555 (N_27555,N_21969,N_22734);
nor U27556 (N_27556,N_21289,N_19627);
xnor U27557 (N_27557,N_22213,N_19719);
nor U27558 (N_27558,N_22225,N_23752);
or U27559 (N_27559,N_23338,N_19104);
nor U27560 (N_27560,N_22529,N_18818);
xor U27561 (N_27561,N_20577,N_23647);
or U27562 (N_27562,N_21600,N_23571);
xor U27563 (N_27563,N_19498,N_18262);
nand U27564 (N_27564,N_22122,N_20923);
nand U27565 (N_27565,N_21880,N_23705);
and U27566 (N_27566,N_18431,N_18850);
or U27567 (N_27567,N_21144,N_23014);
nor U27568 (N_27568,N_18738,N_19096);
nand U27569 (N_27569,N_18531,N_22386);
and U27570 (N_27570,N_22589,N_23913);
or U27571 (N_27571,N_20148,N_18199);
and U27572 (N_27572,N_19987,N_18130);
nand U27573 (N_27573,N_18690,N_20786);
nor U27574 (N_27574,N_22637,N_22597);
xnor U27575 (N_27575,N_19119,N_20768);
or U27576 (N_27576,N_23201,N_23153);
xnor U27577 (N_27577,N_23234,N_18444);
and U27578 (N_27578,N_18138,N_21870);
nand U27579 (N_27579,N_20614,N_21551);
and U27580 (N_27580,N_18718,N_20651);
nand U27581 (N_27581,N_20753,N_19785);
or U27582 (N_27582,N_22376,N_19997);
nor U27583 (N_27583,N_21385,N_18787);
or U27584 (N_27584,N_22700,N_19189);
and U27585 (N_27585,N_20417,N_19593);
xor U27586 (N_27586,N_18361,N_22660);
or U27587 (N_27587,N_22866,N_22495);
nand U27588 (N_27588,N_18019,N_18203);
nor U27589 (N_27589,N_22137,N_19860);
and U27590 (N_27590,N_21075,N_21405);
or U27591 (N_27591,N_20627,N_19069);
or U27592 (N_27592,N_22593,N_22144);
xor U27593 (N_27593,N_18792,N_22467);
nor U27594 (N_27594,N_22155,N_21281);
and U27595 (N_27595,N_20123,N_20097);
xor U27596 (N_27596,N_19338,N_22387);
or U27597 (N_27597,N_21331,N_19806);
nand U27598 (N_27598,N_20359,N_21323);
nand U27599 (N_27599,N_19277,N_23242);
or U27600 (N_27600,N_19549,N_21943);
and U27601 (N_27601,N_22767,N_19725);
xnor U27602 (N_27602,N_20373,N_20826);
nor U27603 (N_27603,N_18665,N_23081);
nand U27604 (N_27604,N_19725,N_22882);
and U27605 (N_27605,N_22818,N_22114);
xnor U27606 (N_27606,N_20156,N_18121);
nand U27607 (N_27607,N_19417,N_22292);
nand U27608 (N_27608,N_18638,N_20643);
nor U27609 (N_27609,N_22961,N_21364);
xnor U27610 (N_27610,N_22756,N_22156);
nand U27611 (N_27611,N_21724,N_23083);
nand U27612 (N_27612,N_18055,N_18922);
nor U27613 (N_27613,N_22505,N_18336);
or U27614 (N_27614,N_22205,N_18817);
and U27615 (N_27615,N_21659,N_19452);
xnor U27616 (N_27616,N_21681,N_23367);
nand U27617 (N_27617,N_23622,N_22211);
nor U27618 (N_27618,N_23845,N_23581);
nand U27619 (N_27619,N_21055,N_23352);
xnor U27620 (N_27620,N_21050,N_23456);
nand U27621 (N_27621,N_18257,N_20020);
or U27622 (N_27622,N_22522,N_18381);
and U27623 (N_27623,N_19567,N_21116);
nor U27624 (N_27624,N_21794,N_18428);
xor U27625 (N_27625,N_22978,N_19086);
xor U27626 (N_27626,N_20136,N_18720);
and U27627 (N_27627,N_23419,N_19613);
or U27628 (N_27628,N_21884,N_18404);
or U27629 (N_27629,N_20493,N_23344);
and U27630 (N_27630,N_20339,N_20134);
nand U27631 (N_27631,N_23796,N_20885);
and U27632 (N_27632,N_23877,N_20830);
xor U27633 (N_27633,N_22421,N_20497);
xnor U27634 (N_27634,N_21851,N_23923);
nand U27635 (N_27635,N_23033,N_21634);
and U27636 (N_27636,N_19255,N_20285);
nor U27637 (N_27637,N_20239,N_23633);
xor U27638 (N_27638,N_19914,N_22988);
nand U27639 (N_27639,N_22379,N_21263);
xor U27640 (N_27640,N_21126,N_20426);
nor U27641 (N_27641,N_19026,N_21544);
xnor U27642 (N_27642,N_20308,N_20837);
nor U27643 (N_27643,N_20362,N_23647);
or U27644 (N_27644,N_23614,N_21208);
or U27645 (N_27645,N_22256,N_22837);
nor U27646 (N_27646,N_19239,N_19519);
and U27647 (N_27647,N_21867,N_19040);
xor U27648 (N_27648,N_19307,N_19023);
nor U27649 (N_27649,N_23472,N_20714);
xor U27650 (N_27650,N_20796,N_22735);
nor U27651 (N_27651,N_19067,N_21691);
xnor U27652 (N_27652,N_19448,N_20653);
nor U27653 (N_27653,N_23635,N_23661);
nand U27654 (N_27654,N_19274,N_18518);
nor U27655 (N_27655,N_18683,N_22193);
xnor U27656 (N_27656,N_18982,N_19307);
or U27657 (N_27657,N_19240,N_19421);
xor U27658 (N_27658,N_22029,N_20654);
nand U27659 (N_27659,N_20147,N_21079);
xnor U27660 (N_27660,N_20100,N_18939);
or U27661 (N_27661,N_21032,N_18962);
nand U27662 (N_27662,N_20392,N_18507);
xnor U27663 (N_27663,N_19213,N_18738);
and U27664 (N_27664,N_21175,N_23640);
xor U27665 (N_27665,N_19282,N_23518);
and U27666 (N_27666,N_20156,N_23673);
or U27667 (N_27667,N_19074,N_21211);
or U27668 (N_27668,N_18952,N_20677);
nor U27669 (N_27669,N_23751,N_20096);
or U27670 (N_27670,N_22105,N_22650);
nand U27671 (N_27671,N_22721,N_18474);
and U27672 (N_27672,N_23135,N_18776);
xor U27673 (N_27673,N_21989,N_20836);
and U27674 (N_27674,N_23783,N_21421);
nand U27675 (N_27675,N_18816,N_23816);
xor U27676 (N_27676,N_20697,N_22261);
xor U27677 (N_27677,N_18257,N_21246);
and U27678 (N_27678,N_19498,N_21613);
nand U27679 (N_27679,N_21524,N_23299);
nor U27680 (N_27680,N_22503,N_20728);
or U27681 (N_27681,N_20983,N_23980);
nand U27682 (N_27682,N_19285,N_20485);
nand U27683 (N_27683,N_21734,N_19703);
nand U27684 (N_27684,N_22863,N_21688);
nor U27685 (N_27685,N_22399,N_19081);
nor U27686 (N_27686,N_23256,N_23053);
xor U27687 (N_27687,N_23220,N_21966);
nor U27688 (N_27688,N_20281,N_23020);
nor U27689 (N_27689,N_18860,N_23483);
and U27690 (N_27690,N_22938,N_23309);
or U27691 (N_27691,N_18533,N_19222);
and U27692 (N_27692,N_20617,N_22296);
xnor U27693 (N_27693,N_23820,N_20047);
and U27694 (N_27694,N_18950,N_20415);
or U27695 (N_27695,N_23377,N_18493);
xor U27696 (N_27696,N_18558,N_19844);
or U27697 (N_27697,N_23462,N_23751);
xnor U27698 (N_27698,N_23629,N_19344);
xnor U27699 (N_27699,N_21404,N_22237);
or U27700 (N_27700,N_19379,N_19726);
nor U27701 (N_27701,N_19756,N_19332);
or U27702 (N_27702,N_23677,N_19869);
nor U27703 (N_27703,N_21929,N_23152);
nand U27704 (N_27704,N_18630,N_20176);
nand U27705 (N_27705,N_20523,N_23058);
nand U27706 (N_27706,N_21080,N_19871);
nand U27707 (N_27707,N_22593,N_18010);
xor U27708 (N_27708,N_21847,N_19317);
xnor U27709 (N_27709,N_21851,N_18063);
or U27710 (N_27710,N_18873,N_19501);
or U27711 (N_27711,N_23397,N_22471);
nand U27712 (N_27712,N_18129,N_19026);
nand U27713 (N_27713,N_18887,N_18604);
nor U27714 (N_27714,N_21308,N_23400);
xnor U27715 (N_27715,N_19618,N_20001);
nand U27716 (N_27716,N_21386,N_23641);
nand U27717 (N_27717,N_22881,N_19999);
xnor U27718 (N_27718,N_19926,N_23619);
nor U27719 (N_27719,N_22021,N_18266);
and U27720 (N_27720,N_20878,N_18021);
xor U27721 (N_27721,N_22575,N_19410);
and U27722 (N_27722,N_19921,N_18663);
xor U27723 (N_27723,N_18011,N_18877);
nand U27724 (N_27724,N_19425,N_22805);
nor U27725 (N_27725,N_18509,N_19420);
nand U27726 (N_27726,N_20789,N_19921);
or U27727 (N_27727,N_18058,N_20415);
and U27728 (N_27728,N_22135,N_21112);
nand U27729 (N_27729,N_20166,N_23652);
or U27730 (N_27730,N_20208,N_23593);
xor U27731 (N_27731,N_21735,N_22789);
or U27732 (N_27732,N_21035,N_18296);
and U27733 (N_27733,N_19426,N_23393);
or U27734 (N_27734,N_18420,N_19127);
or U27735 (N_27735,N_23517,N_22459);
or U27736 (N_27736,N_20609,N_20264);
xnor U27737 (N_27737,N_23739,N_18505);
nor U27738 (N_27738,N_20645,N_18702);
nand U27739 (N_27739,N_19140,N_23853);
and U27740 (N_27740,N_18710,N_22713);
xnor U27741 (N_27741,N_22909,N_22996);
nor U27742 (N_27742,N_19060,N_19462);
nand U27743 (N_27743,N_21722,N_19720);
nand U27744 (N_27744,N_18879,N_20057);
nor U27745 (N_27745,N_19042,N_19894);
xor U27746 (N_27746,N_22112,N_22286);
nor U27747 (N_27747,N_22721,N_20081);
or U27748 (N_27748,N_20412,N_21396);
nand U27749 (N_27749,N_23631,N_20728);
nand U27750 (N_27750,N_18461,N_19510);
xor U27751 (N_27751,N_21144,N_22845);
nor U27752 (N_27752,N_20748,N_19574);
xor U27753 (N_27753,N_21620,N_22213);
nand U27754 (N_27754,N_22488,N_21827);
nand U27755 (N_27755,N_20962,N_20783);
nand U27756 (N_27756,N_21334,N_22379);
xor U27757 (N_27757,N_21571,N_23977);
and U27758 (N_27758,N_18313,N_23269);
xnor U27759 (N_27759,N_18908,N_23508);
and U27760 (N_27760,N_21488,N_23816);
nand U27761 (N_27761,N_19570,N_22682);
or U27762 (N_27762,N_22596,N_21049);
nand U27763 (N_27763,N_18390,N_19841);
nor U27764 (N_27764,N_21960,N_19609);
xnor U27765 (N_27765,N_18947,N_20404);
nor U27766 (N_27766,N_20899,N_23664);
or U27767 (N_27767,N_18902,N_20265);
nor U27768 (N_27768,N_18369,N_19888);
nor U27769 (N_27769,N_21965,N_21013);
and U27770 (N_27770,N_20924,N_19750);
nand U27771 (N_27771,N_19858,N_22147);
xor U27772 (N_27772,N_21283,N_22073);
or U27773 (N_27773,N_19011,N_23909);
nand U27774 (N_27774,N_23508,N_22127);
nor U27775 (N_27775,N_19078,N_23782);
nor U27776 (N_27776,N_18312,N_18641);
xor U27777 (N_27777,N_22912,N_23700);
or U27778 (N_27778,N_22742,N_23486);
xor U27779 (N_27779,N_20181,N_21556);
nor U27780 (N_27780,N_21827,N_22308);
xor U27781 (N_27781,N_23265,N_19911);
nand U27782 (N_27782,N_20703,N_23807);
and U27783 (N_27783,N_23759,N_23744);
or U27784 (N_27784,N_21436,N_21578);
and U27785 (N_27785,N_21470,N_18852);
nor U27786 (N_27786,N_19602,N_18236);
and U27787 (N_27787,N_19183,N_23683);
nand U27788 (N_27788,N_22639,N_22643);
nor U27789 (N_27789,N_18083,N_19847);
or U27790 (N_27790,N_22405,N_19294);
nor U27791 (N_27791,N_19010,N_18049);
xor U27792 (N_27792,N_23194,N_21767);
and U27793 (N_27793,N_19813,N_18770);
nand U27794 (N_27794,N_23491,N_21046);
nor U27795 (N_27795,N_18500,N_18690);
xnor U27796 (N_27796,N_21414,N_18549);
and U27797 (N_27797,N_18306,N_22479);
nor U27798 (N_27798,N_22298,N_23853);
nor U27799 (N_27799,N_19680,N_23891);
nand U27800 (N_27800,N_19965,N_18655);
and U27801 (N_27801,N_20767,N_21063);
or U27802 (N_27802,N_19923,N_19534);
or U27803 (N_27803,N_19845,N_18717);
nand U27804 (N_27804,N_23848,N_23864);
nand U27805 (N_27805,N_20104,N_19829);
or U27806 (N_27806,N_23600,N_18531);
nand U27807 (N_27807,N_22983,N_22231);
and U27808 (N_27808,N_23673,N_20934);
or U27809 (N_27809,N_22457,N_23366);
or U27810 (N_27810,N_19363,N_18245);
or U27811 (N_27811,N_21866,N_22310);
or U27812 (N_27812,N_18326,N_21662);
or U27813 (N_27813,N_22896,N_23753);
nor U27814 (N_27814,N_19995,N_18037);
xnor U27815 (N_27815,N_20083,N_22318);
and U27816 (N_27816,N_23557,N_20496);
or U27817 (N_27817,N_23460,N_19410);
or U27818 (N_27818,N_22838,N_23254);
xnor U27819 (N_27819,N_20844,N_18017);
or U27820 (N_27820,N_22219,N_22896);
xnor U27821 (N_27821,N_20036,N_18418);
nor U27822 (N_27822,N_21343,N_22633);
nand U27823 (N_27823,N_19587,N_20181);
and U27824 (N_27824,N_23055,N_20882);
nor U27825 (N_27825,N_20299,N_21428);
and U27826 (N_27826,N_19860,N_23195);
and U27827 (N_27827,N_21358,N_21820);
or U27828 (N_27828,N_18861,N_21381);
nor U27829 (N_27829,N_23772,N_23545);
and U27830 (N_27830,N_22691,N_23019);
and U27831 (N_27831,N_22764,N_20555);
and U27832 (N_27832,N_19395,N_23255);
and U27833 (N_27833,N_20819,N_18194);
or U27834 (N_27834,N_20426,N_22659);
nand U27835 (N_27835,N_20701,N_23102);
xor U27836 (N_27836,N_18940,N_20042);
or U27837 (N_27837,N_18771,N_19937);
nand U27838 (N_27838,N_22776,N_18318);
nor U27839 (N_27839,N_22404,N_22883);
xnor U27840 (N_27840,N_22548,N_18938);
xor U27841 (N_27841,N_23905,N_19142);
nand U27842 (N_27842,N_19224,N_23642);
nor U27843 (N_27843,N_23219,N_19646);
nor U27844 (N_27844,N_22147,N_18580);
and U27845 (N_27845,N_20497,N_19047);
and U27846 (N_27846,N_23227,N_21835);
nor U27847 (N_27847,N_20446,N_21279);
nor U27848 (N_27848,N_19085,N_21953);
xnor U27849 (N_27849,N_20074,N_23803);
nand U27850 (N_27850,N_22586,N_22787);
and U27851 (N_27851,N_19209,N_20640);
xnor U27852 (N_27852,N_23981,N_20235);
and U27853 (N_27853,N_21196,N_23445);
nor U27854 (N_27854,N_23431,N_21690);
or U27855 (N_27855,N_23034,N_20571);
and U27856 (N_27856,N_18714,N_23537);
nand U27857 (N_27857,N_20963,N_19636);
nor U27858 (N_27858,N_19097,N_18396);
nand U27859 (N_27859,N_20462,N_23187);
nor U27860 (N_27860,N_23497,N_22085);
or U27861 (N_27861,N_20967,N_20167);
or U27862 (N_27862,N_23377,N_18925);
nand U27863 (N_27863,N_21909,N_22258);
xnor U27864 (N_27864,N_20163,N_18027);
xnor U27865 (N_27865,N_19058,N_22574);
or U27866 (N_27866,N_21739,N_21040);
or U27867 (N_27867,N_23803,N_20929);
nor U27868 (N_27868,N_18586,N_23339);
nand U27869 (N_27869,N_23947,N_18965);
and U27870 (N_27870,N_22639,N_18350);
xor U27871 (N_27871,N_18768,N_18383);
or U27872 (N_27872,N_20830,N_22663);
or U27873 (N_27873,N_21399,N_22753);
nand U27874 (N_27874,N_22317,N_21729);
xnor U27875 (N_27875,N_23790,N_22555);
nand U27876 (N_27876,N_19528,N_19182);
and U27877 (N_27877,N_20168,N_23416);
nor U27878 (N_27878,N_20853,N_23444);
and U27879 (N_27879,N_21211,N_19254);
and U27880 (N_27880,N_22135,N_23256);
and U27881 (N_27881,N_19852,N_21718);
or U27882 (N_27882,N_20210,N_19464);
nand U27883 (N_27883,N_22417,N_23206);
nor U27884 (N_27884,N_18126,N_18043);
and U27885 (N_27885,N_20618,N_18243);
or U27886 (N_27886,N_22815,N_19183);
xnor U27887 (N_27887,N_20621,N_22564);
nand U27888 (N_27888,N_20261,N_20921);
and U27889 (N_27889,N_20650,N_22286);
or U27890 (N_27890,N_19552,N_19992);
and U27891 (N_27891,N_22557,N_19775);
xnor U27892 (N_27892,N_20942,N_22601);
xnor U27893 (N_27893,N_22320,N_20218);
nand U27894 (N_27894,N_20157,N_19667);
nor U27895 (N_27895,N_22685,N_18697);
nor U27896 (N_27896,N_23298,N_20064);
and U27897 (N_27897,N_19917,N_21752);
or U27898 (N_27898,N_19304,N_22303);
nor U27899 (N_27899,N_19311,N_20871);
nor U27900 (N_27900,N_19067,N_18694);
or U27901 (N_27901,N_18467,N_20665);
nand U27902 (N_27902,N_20972,N_22371);
and U27903 (N_27903,N_23438,N_21839);
nor U27904 (N_27904,N_22662,N_23941);
xnor U27905 (N_27905,N_20948,N_22639);
and U27906 (N_27906,N_23384,N_20533);
nor U27907 (N_27907,N_22518,N_23971);
nor U27908 (N_27908,N_22200,N_23585);
nor U27909 (N_27909,N_19547,N_18400);
xnor U27910 (N_27910,N_18845,N_19424);
and U27911 (N_27911,N_21318,N_18983);
or U27912 (N_27912,N_20802,N_20668);
or U27913 (N_27913,N_19756,N_23099);
nor U27914 (N_27914,N_20743,N_19546);
xor U27915 (N_27915,N_22088,N_22011);
xnor U27916 (N_27916,N_19616,N_19249);
and U27917 (N_27917,N_22524,N_19374);
xor U27918 (N_27918,N_22402,N_19647);
xor U27919 (N_27919,N_22622,N_21750);
and U27920 (N_27920,N_20853,N_20458);
nor U27921 (N_27921,N_21201,N_20093);
xnor U27922 (N_27922,N_21414,N_18951);
or U27923 (N_27923,N_22519,N_23969);
or U27924 (N_27924,N_21604,N_23613);
or U27925 (N_27925,N_19547,N_18756);
or U27926 (N_27926,N_19444,N_23542);
and U27927 (N_27927,N_20253,N_23978);
nand U27928 (N_27928,N_21853,N_22987);
xnor U27929 (N_27929,N_19779,N_20899);
xnor U27930 (N_27930,N_18410,N_20125);
nor U27931 (N_27931,N_23594,N_20624);
nor U27932 (N_27932,N_18059,N_18394);
or U27933 (N_27933,N_22608,N_18381);
and U27934 (N_27934,N_18164,N_18532);
and U27935 (N_27935,N_19732,N_20988);
nor U27936 (N_27936,N_18289,N_23616);
or U27937 (N_27937,N_19474,N_23215);
nor U27938 (N_27938,N_18704,N_20870);
nor U27939 (N_27939,N_23208,N_20609);
or U27940 (N_27940,N_18964,N_22245);
nor U27941 (N_27941,N_18208,N_21918);
or U27942 (N_27942,N_21742,N_23496);
nand U27943 (N_27943,N_21660,N_23355);
or U27944 (N_27944,N_20597,N_22280);
nor U27945 (N_27945,N_22095,N_22131);
nor U27946 (N_27946,N_22535,N_18408);
nand U27947 (N_27947,N_20689,N_21916);
nand U27948 (N_27948,N_22426,N_18880);
nand U27949 (N_27949,N_22236,N_19581);
and U27950 (N_27950,N_23806,N_20752);
or U27951 (N_27951,N_19475,N_21421);
or U27952 (N_27952,N_20425,N_22611);
xnor U27953 (N_27953,N_22538,N_22804);
or U27954 (N_27954,N_21703,N_21038);
nor U27955 (N_27955,N_18702,N_19765);
and U27956 (N_27956,N_20874,N_20440);
and U27957 (N_27957,N_22744,N_18268);
nand U27958 (N_27958,N_18529,N_20810);
nand U27959 (N_27959,N_18863,N_18722);
xnor U27960 (N_27960,N_21891,N_18742);
xnor U27961 (N_27961,N_18815,N_20074);
and U27962 (N_27962,N_19305,N_21268);
nor U27963 (N_27963,N_22485,N_18345);
or U27964 (N_27964,N_20322,N_21340);
xnor U27965 (N_27965,N_23038,N_23434);
nand U27966 (N_27966,N_22130,N_23096);
xor U27967 (N_27967,N_19415,N_21918);
nand U27968 (N_27968,N_23868,N_23614);
or U27969 (N_27969,N_18435,N_20541);
nand U27970 (N_27970,N_22380,N_23295);
xor U27971 (N_27971,N_20233,N_22036);
nor U27972 (N_27972,N_19982,N_21434);
nand U27973 (N_27973,N_22032,N_23346);
nor U27974 (N_27974,N_19649,N_20674);
nand U27975 (N_27975,N_22030,N_21809);
or U27976 (N_27976,N_18342,N_19057);
xnor U27977 (N_27977,N_20654,N_18960);
nor U27978 (N_27978,N_22627,N_23270);
and U27979 (N_27979,N_19353,N_18572);
nand U27980 (N_27980,N_23924,N_20096);
or U27981 (N_27981,N_21360,N_21681);
or U27982 (N_27982,N_18855,N_19374);
xor U27983 (N_27983,N_23006,N_20875);
or U27984 (N_27984,N_22721,N_22291);
nor U27985 (N_27985,N_19894,N_19008);
and U27986 (N_27986,N_19441,N_19567);
or U27987 (N_27987,N_19601,N_18998);
and U27988 (N_27988,N_22052,N_18806);
xnor U27989 (N_27989,N_21319,N_22961);
nor U27990 (N_27990,N_20799,N_20954);
nor U27991 (N_27991,N_19440,N_22120);
nor U27992 (N_27992,N_22429,N_21915);
or U27993 (N_27993,N_20118,N_20979);
or U27994 (N_27994,N_18326,N_21291);
or U27995 (N_27995,N_20073,N_21323);
nor U27996 (N_27996,N_22718,N_23787);
nand U27997 (N_27997,N_19291,N_21164);
or U27998 (N_27998,N_23622,N_19566);
nor U27999 (N_27999,N_23490,N_18975);
xor U28000 (N_28000,N_22870,N_20650);
or U28001 (N_28001,N_22295,N_18764);
or U28002 (N_28002,N_18766,N_18044);
and U28003 (N_28003,N_19714,N_20751);
nand U28004 (N_28004,N_20259,N_23350);
nor U28005 (N_28005,N_20929,N_20251);
nand U28006 (N_28006,N_20331,N_19285);
xor U28007 (N_28007,N_22352,N_18817);
or U28008 (N_28008,N_19178,N_22094);
nor U28009 (N_28009,N_21603,N_23863);
nor U28010 (N_28010,N_21277,N_20857);
nand U28011 (N_28011,N_20342,N_22273);
xor U28012 (N_28012,N_22385,N_19468);
nor U28013 (N_28013,N_23312,N_19773);
nand U28014 (N_28014,N_18544,N_20621);
nand U28015 (N_28015,N_21442,N_19110);
or U28016 (N_28016,N_21864,N_22417);
or U28017 (N_28017,N_23570,N_21029);
and U28018 (N_28018,N_18695,N_22534);
nand U28019 (N_28019,N_22517,N_20936);
or U28020 (N_28020,N_20310,N_22626);
nand U28021 (N_28021,N_19392,N_21394);
or U28022 (N_28022,N_18596,N_20641);
nor U28023 (N_28023,N_23626,N_20166);
and U28024 (N_28024,N_20504,N_18647);
or U28025 (N_28025,N_18599,N_19696);
or U28026 (N_28026,N_19632,N_18169);
nor U28027 (N_28027,N_22692,N_18640);
nand U28028 (N_28028,N_21031,N_18607);
nor U28029 (N_28029,N_19610,N_23814);
xnor U28030 (N_28030,N_19365,N_19306);
or U28031 (N_28031,N_22364,N_22293);
xnor U28032 (N_28032,N_20197,N_18110);
and U28033 (N_28033,N_22894,N_21959);
nand U28034 (N_28034,N_21554,N_19007);
nand U28035 (N_28035,N_21283,N_20546);
and U28036 (N_28036,N_23583,N_18608);
or U28037 (N_28037,N_18307,N_20126);
nor U28038 (N_28038,N_21697,N_19279);
nand U28039 (N_28039,N_19286,N_20049);
or U28040 (N_28040,N_21040,N_18029);
nor U28041 (N_28041,N_20032,N_23978);
and U28042 (N_28042,N_21253,N_19307);
and U28043 (N_28043,N_22853,N_22551);
nor U28044 (N_28044,N_23174,N_20402);
nor U28045 (N_28045,N_18191,N_22903);
nand U28046 (N_28046,N_23895,N_19560);
xnor U28047 (N_28047,N_20637,N_20676);
nor U28048 (N_28048,N_22445,N_21953);
xnor U28049 (N_28049,N_18403,N_20332);
nand U28050 (N_28050,N_20490,N_18762);
or U28051 (N_28051,N_19308,N_18773);
and U28052 (N_28052,N_23894,N_22402);
and U28053 (N_28053,N_18641,N_22037);
and U28054 (N_28054,N_23002,N_18921);
or U28055 (N_28055,N_19325,N_21580);
nand U28056 (N_28056,N_19482,N_18838);
or U28057 (N_28057,N_23337,N_21716);
xor U28058 (N_28058,N_21468,N_22700);
nand U28059 (N_28059,N_23392,N_18245);
nand U28060 (N_28060,N_19847,N_21531);
xor U28061 (N_28061,N_18195,N_22539);
xor U28062 (N_28062,N_23575,N_22354);
xnor U28063 (N_28063,N_21822,N_20934);
and U28064 (N_28064,N_21029,N_18716);
nand U28065 (N_28065,N_23001,N_21821);
and U28066 (N_28066,N_21105,N_18408);
and U28067 (N_28067,N_19641,N_18131);
xor U28068 (N_28068,N_19064,N_20575);
nand U28069 (N_28069,N_21970,N_18818);
nor U28070 (N_28070,N_22700,N_22120);
or U28071 (N_28071,N_21880,N_21258);
xor U28072 (N_28072,N_23625,N_18730);
xor U28073 (N_28073,N_18152,N_22829);
nand U28074 (N_28074,N_18724,N_18272);
nor U28075 (N_28075,N_23770,N_23902);
nand U28076 (N_28076,N_22633,N_21795);
and U28077 (N_28077,N_22909,N_20946);
or U28078 (N_28078,N_21185,N_21331);
and U28079 (N_28079,N_22030,N_20431);
and U28080 (N_28080,N_20289,N_19219);
or U28081 (N_28081,N_19802,N_22542);
xnor U28082 (N_28082,N_20179,N_18257);
xnor U28083 (N_28083,N_22467,N_21467);
nand U28084 (N_28084,N_19755,N_23459);
nor U28085 (N_28085,N_21137,N_19638);
nor U28086 (N_28086,N_23131,N_18555);
xnor U28087 (N_28087,N_19568,N_23817);
nor U28088 (N_28088,N_21645,N_18135);
or U28089 (N_28089,N_22590,N_19435);
nand U28090 (N_28090,N_21889,N_21870);
and U28091 (N_28091,N_21968,N_18428);
nand U28092 (N_28092,N_18480,N_21010);
nor U28093 (N_28093,N_19939,N_22449);
or U28094 (N_28094,N_22691,N_23719);
or U28095 (N_28095,N_23716,N_18195);
xor U28096 (N_28096,N_22766,N_21724);
or U28097 (N_28097,N_20310,N_19482);
nor U28098 (N_28098,N_21431,N_23756);
and U28099 (N_28099,N_19950,N_20767);
xor U28100 (N_28100,N_20897,N_22422);
nand U28101 (N_28101,N_19848,N_21874);
nor U28102 (N_28102,N_23597,N_21208);
and U28103 (N_28103,N_20265,N_18641);
nor U28104 (N_28104,N_21192,N_23732);
and U28105 (N_28105,N_20894,N_22432);
xor U28106 (N_28106,N_18495,N_23081);
nand U28107 (N_28107,N_22383,N_21358);
and U28108 (N_28108,N_21595,N_19082);
nand U28109 (N_28109,N_18548,N_18852);
nand U28110 (N_28110,N_22042,N_19480);
and U28111 (N_28111,N_18581,N_21983);
nor U28112 (N_28112,N_19076,N_21953);
nor U28113 (N_28113,N_19616,N_20906);
xor U28114 (N_28114,N_22640,N_21668);
nor U28115 (N_28115,N_22998,N_19731);
nor U28116 (N_28116,N_18210,N_23945);
nor U28117 (N_28117,N_22704,N_18458);
and U28118 (N_28118,N_21160,N_18187);
nand U28119 (N_28119,N_23946,N_22868);
or U28120 (N_28120,N_22158,N_19918);
nor U28121 (N_28121,N_22956,N_21255);
and U28122 (N_28122,N_18163,N_18473);
or U28123 (N_28123,N_22942,N_20067);
or U28124 (N_28124,N_23606,N_19525);
or U28125 (N_28125,N_22817,N_21882);
nor U28126 (N_28126,N_18452,N_21880);
or U28127 (N_28127,N_19440,N_20890);
xor U28128 (N_28128,N_21654,N_22398);
xnor U28129 (N_28129,N_20086,N_22851);
nand U28130 (N_28130,N_20719,N_18948);
nor U28131 (N_28131,N_20345,N_19938);
xnor U28132 (N_28132,N_23872,N_23052);
or U28133 (N_28133,N_23926,N_21433);
and U28134 (N_28134,N_23019,N_21171);
xor U28135 (N_28135,N_22000,N_20499);
and U28136 (N_28136,N_20034,N_21472);
xnor U28137 (N_28137,N_20950,N_22582);
or U28138 (N_28138,N_21846,N_20496);
xor U28139 (N_28139,N_20243,N_23015);
nor U28140 (N_28140,N_19219,N_19667);
or U28141 (N_28141,N_22276,N_19351);
xor U28142 (N_28142,N_21318,N_20724);
and U28143 (N_28143,N_21061,N_23386);
and U28144 (N_28144,N_21380,N_19705);
nand U28145 (N_28145,N_18610,N_20926);
and U28146 (N_28146,N_22663,N_19670);
nor U28147 (N_28147,N_23672,N_20008);
and U28148 (N_28148,N_22945,N_19913);
xor U28149 (N_28149,N_18898,N_22113);
nand U28150 (N_28150,N_19225,N_19383);
or U28151 (N_28151,N_23857,N_23806);
xor U28152 (N_28152,N_22473,N_18196);
xor U28153 (N_28153,N_23632,N_23726);
nand U28154 (N_28154,N_21845,N_23984);
nand U28155 (N_28155,N_18711,N_18831);
xnor U28156 (N_28156,N_21178,N_23899);
and U28157 (N_28157,N_21381,N_23544);
or U28158 (N_28158,N_22544,N_21159);
xnor U28159 (N_28159,N_20914,N_22531);
xor U28160 (N_28160,N_19618,N_23917);
or U28161 (N_28161,N_18260,N_22717);
xor U28162 (N_28162,N_21792,N_23076);
nor U28163 (N_28163,N_20981,N_23604);
and U28164 (N_28164,N_21881,N_20912);
xnor U28165 (N_28165,N_22434,N_18316);
nand U28166 (N_28166,N_23330,N_18237);
and U28167 (N_28167,N_21699,N_19257);
nor U28168 (N_28168,N_22360,N_21759);
nand U28169 (N_28169,N_18845,N_21119);
or U28170 (N_28170,N_18518,N_22440);
nor U28171 (N_28171,N_19171,N_19567);
nand U28172 (N_28172,N_19084,N_23829);
or U28173 (N_28173,N_20994,N_21993);
nor U28174 (N_28174,N_19392,N_21749);
xnor U28175 (N_28175,N_23094,N_19181);
nor U28176 (N_28176,N_19312,N_19334);
or U28177 (N_28177,N_20850,N_19435);
nand U28178 (N_28178,N_23944,N_18756);
or U28179 (N_28179,N_21757,N_19290);
nor U28180 (N_28180,N_23267,N_20637);
and U28181 (N_28181,N_22531,N_21926);
or U28182 (N_28182,N_19309,N_23929);
xor U28183 (N_28183,N_18433,N_20534);
nand U28184 (N_28184,N_18997,N_22198);
nor U28185 (N_28185,N_19104,N_20901);
or U28186 (N_28186,N_23815,N_21693);
and U28187 (N_28187,N_19444,N_23034);
and U28188 (N_28188,N_20396,N_22659);
nand U28189 (N_28189,N_18919,N_21299);
and U28190 (N_28190,N_20775,N_19592);
nand U28191 (N_28191,N_21420,N_18395);
or U28192 (N_28192,N_19043,N_22836);
or U28193 (N_28193,N_19227,N_22442);
or U28194 (N_28194,N_18527,N_21438);
or U28195 (N_28195,N_23584,N_19044);
and U28196 (N_28196,N_18126,N_18108);
xnor U28197 (N_28197,N_18313,N_23777);
and U28198 (N_28198,N_18725,N_22290);
nand U28199 (N_28199,N_18511,N_23557);
and U28200 (N_28200,N_22367,N_23863);
nand U28201 (N_28201,N_19359,N_21970);
or U28202 (N_28202,N_18948,N_18578);
or U28203 (N_28203,N_23270,N_19065);
xnor U28204 (N_28204,N_19775,N_23110);
or U28205 (N_28205,N_20199,N_21240);
or U28206 (N_28206,N_18778,N_18834);
or U28207 (N_28207,N_19216,N_19930);
nor U28208 (N_28208,N_22288,N_18884);
and U28209 (N_28209,N_20502,N_23872);
xnor U28210 (N_28210,N_19803,N_20643);
or U28211 (N_28211,N_18511,N_20091);
xor U28212 (N_28212,N_20748,N_18050);
xor U28213 (N_28213,N_21961,N_18742);
and U28214 (N_28214,N_20513,N_19540);
xor U28215 (N_28215,N_18174,N_20733);
nand U28216 (N_28216,N_20206,N_23148);
and U28217 (N_28217,N_20833,N_21141);
or U28218 (N_28218,N_20852,N_20886);
and U28219 (N_28219,N_19379,N_19698);
xnor U28220 (N_28220,N_20753,N_22568);
and U28221 (N_28221,N_19928,N_19479);
nand U28222 (N_28222,N_20463,N_22491);
xnor U28223 (N_28223,N_21619,N_21266);
nand U28224 (N_28224,N_22206,N_23118);
and U28225 (N_28225,N_23193,N_23534);
xnor U28226 (N_28226,N_19022,N_19291);
nand U28227 (N_28227,N_21007,N_19267);
and U28228 (N_28228,N_21111,N_20337);
xnor U28229 (N_28229,N_18624,N_23306);
nand U28230 (N_28230,N_20605,N_23964);
and U28231 (N_28231,N_19485,N_18108);
and U28232 (N_28232,N_18912,N_23872);
and U28233 (N_28233,N_19988,N_23399);
xnor U28234 (N_28234,N_19307,N_20647);
nand U28235 (N_28235,N_19535,N_19867);
xor U28236 (N_28236,N_22739,N_19552);
and U28237 (N_28237,N_22261,N_23833);
nand U28238 (N_28238,N_21105,N_20184);
nor U28239 (N_28239,N_22059,N_23138);
nand U28240 (N_28240,N_23820,N_21404);
or U28241 (N_28241,N_18606,N_19709);
and U28242 (N_28242,N_23949,N_23168);
xor U28243 (N_28243,N_21609,N_20944);
or U28244 (N_28244,N_18127,N_18611);
nor U28245 (N_28245,N_18529,N_23066);
nor U28246 (N_28246,N_19178,N_19474);
and U28247 (N_28247,N_21076,N_23791);
nand U28248 (N_28248,N_19845,N_18319);
xor U28249 (N_28249,N_23504,N_18610);
or U28250 (N_28250,N_19078,N_21460);
or U28251 (N_28251,N_19760,N_18471);
and U28252 (N_28252,N_18818,N_20335);
and U28253 (N_28253,N_21524,N_21153);
and U28254 (N_28254,N_22918,N_22809);
nor U28255 (N_28255,N_18283,N_21700);
nand U28256 (N_28256,N_23443,N_20918);
nor U28257 (N_28257,N_20432,N_18986);
xnor U28258 (N_28258,N_21242,N_19022);
nand U28259 (N_28259,N_18901,N_21167);
and U28260 (N_28260,N_22393,N_22728);
nand U28261 (N_28261,N_19254,N_23109);
nor U28262 (N_28262,N_21075,N_18248);
nor U28263 (N_28263,N_18979,N_18586);
nor U28264 (N_28264,N_18273,N_20578);
nor U28265 (N_28265,N_22881,N_23216);
xor U28266 (N_28266,N_19683,N_19327);
nand U28267 (N_28267,N_19647,N_19488);
nor U28268 (N_28268,N_19784,N_22140);
or U28269 (N_28269,N_18110,N_20247);
and U28270 (N_28270,N_22854,N_20909);
xor U28271 (N_28271,N_23745,N_21692);
xor U28272 (N_28272,N_18603,N_19674);
nor U28273 (N_28273,N_23430,N_23107);
nand U28274 (N_28274,N_23907,N_18350);
nand U28275 (N_28275,N_23366,N_20585);
xor U28276 (N_28276,N_19931,N_23793);
nand U28277 (N_28277,N_20104,N_20551);
nor U28278 (N_28278,N_21718,N_18302);
nand U28279 (N_28279,N_22903,N_19071);
and U28280 (N_28280,N_18017,N_21614);
or U28281 (N_28281,N_19696,N_20858);
nor U28282 (N_28282,N_19921,N_21701);
xnor U28283 (N_28283,N_20359,N_22242);
nor U28284 (N_28284,N_21675,N_23763);
xor U28285 (N_28285,N_23385,N_23292);
or U28286 (N_28286,N_20758,N_19366);
and U28287 (N_28287,N_23159,N_18538);
or U28288 (N_28288,N_23266,N_21209);
nor U28289 (N_28289,N_22319,N_18663);
nor U28290 (N_28290,N_23480,N_23101);
nand U28291 (N_28291,N_18276,N_20049);
or U28292 (N_28292,N_19472,N_20264);
nand U28293 (N_28293,N_19775,N_18430);
nand U28294 (N_28294,N_23785,N_20818);
xnor U28295 (N_28295,N_21104,N_21231);
and U28296 (N_28296,N_21320,N_22809);
and U28297 (N_28297,N_22420,N_18449);
or U28298 (N_28298,N_18378,N_18211);
nor U28299 (N_28299,N_20760,N_20172);
or U28300 (N_28300,N_21337,N_23838);
or U28301 (N_28301,N_20665,N_19297);
nor U28302 (N_28302,N_18256,N_23755);
xnor U28303 (N_28303,N_22254,N_19250);
and U28304 (N_28304,N_20389,N_22654);
xnor U28305 (N_28305,N_22831,N_18244);
xnor U28306 (N_28306,N_20867,N_22238);
or U28307 (N_28307,N_23021,N_18566);
nor U28308 (N_28308,N_21588,N_23001);
and U28309 (N_28309,N_22330,N_18310);
xnor U28310 (N_28310,N_21436,N_20477);
and U28311 (N_28311,N_23782,N_22269);
xor U28312 (N_28312,N_20365,N_21042);
xnor U28313 (N_28313,N_20688,N_22669);
xnor U28314 (N_28314,N_19628,N_22239);
nand U28315 (N_28315,N_22239,N_18014);
nand U28316 (N_28316,N_19858,N_20058);
and U28317 (N_28317,N_19688,N_21720);
xor U28318 (N_28318,N_20495,N_22123);
xor U28319 (N_28319,N_20098,N_19145);
or U28320 (N_28320,N_21360,N_19166);
or U28321 (N_28321,N_18647,N_21295);
or U28322 (N_28322,N_23384,N_21983);
xor U28323 (N_28323,N_21994,N_23005);
nand U28324 (N_28324,N_18674,N_19479);
and U28325 (N_28325,N_22954,N_20091);
nor U28326 (N_28326,N_20078,N_21435);
or U28327 (N_28327,N_18118,N_22821);
nand U28328 (N_28328,N_19612,N_19646);
and U28329 (N_28329,N_18538,N_23738);
nand U28330 (N_28330,N_22908,N_22116);
nand U28331 (N_28331,N_21022,N_18264);
xnor U28332 (N_28332,N_19277,N_22339);
nor U28333 (N_28333,N_22298,N_22078);
xor U28334 (N_28334,N_22593,N_21388);
or U28335 (N_28335,N_18571,N_22657);
or U28336 (N_28336,N_23788,N_21092);
nand U28337 (N_28337,N_22682,N_18476);
xnor U28338 (N_28338,N_18518,N_23772);
xnor U28339 (N_28339,N_19263,N_20436);
nor U28340 (N_28340,N_22069,N_22224);
nand U28341 (N_28341,N_20984,N_23505);
nor U28342 (N_28342,N_22759,N_21637);
nor U28343 (N_28343,N_22058,N_22099);
nor U28344 (N_28344,N_21895,N_18881);
or U28345 (N_28345,N_21338,N_21087);
and U28346 (N_28346,N_18895,N_20418);
nand U28347 (N_28347,N_22015,N_19159);
nand U28348 (N_28348,N_23494,N_22196);
nor U28349 (N_28349,N_21993,N_22458);
nand U28350 (N_28350,N_22020,N_23208);
nor U28351 (N_28351,N_22474,N_19792);
and U28352 (N_28352,N_22568,N_20550);
and U28353 (N_28353,N_18508,N_19757);
and U28354 (N_28354,N_18211,N_23982);
xnor U28355 (N_28355,N_22911,N_22236);
nand U28356 (N_28356,N_22289,N_23942);
and U28357 (N_28357,N_23793,N_21145);
xor U28358 (N_28358,N_23823,N_19966);
xor U28359 (N_28359,N_22391,N_22663);
or U28360 (N_28360,N_21044,N_18516);
nand U28361 (N_28361,N_20855,N_23454);
nor U28362 (N_28362,N_20819,N_18247);
xnor U28363 (N_28363,N_19106,N_23018);
nand U28364 (N_28364,N_21491,N_19816);
or U28365 (N_28365,N_23937,N_21706);
xnor U28366 (N_28366,N_21380,N_20378);
and U28367 (N_28367,N_23687,N_20314);
or U28368 (N_28368,N_22348,N_21149);
and U28369 (N_28369,N_20319,N_19082);
nand U28370 (N_28370,N_19174,N_20959);
nor U28371 (N_28371,N_18091,N_22836);
nor U28372 (N_28372,N_20193,N_22839);
and U28373 (N_28373,N_19987,N_21380);
and U28374 (N_28374,N_23952,N_18781);
and U28375 (N_28375,N_21081,N_22471);
and U28376 (N_28376,N_21480,N_20238);
and U28377 (N_28377,N_23271,N_21115);
xnor U28378 (N_28378,N_21556,N_19990);
and U28379 (N_28379,N_22833,N_19207);
nor U28380 (N_28380,N_23245,N_18449);
xnor U28381 (N_28381,N_23308,N_20192);
or U28382 (N_28382,N_18506,N_23692);
xor U28383 (N_28383,N_21145,N_21405);
nand U28384 (N_28384,N_20620,N_21649);
xnor U28385 (N_28385,N_19221,N_19494);
or U28386 (N_28386,N_23558,N_22006);
nor U28387 (N_28387,N_23949,N_20291);
or U28388 (N_28388,N_22242,N_20676);
and U28389 (N_28389,N_22317,N_18379);
or U28390 (N_28390,N_18284,N_22355);
xnor U28391 (N_28391,N_23233,N_22109);
nor U28392 (N_28392,N_18365,N_19775);
or U28393 (N_28393,N_18620,N_18590);
nand U28394 (N_28394,N_22464,N_19024);
nor U28395 (N_28395,N_22201,N_22188);
xor U28396 (N_28396,N_21460,N_22585);
nand U28397 (N_28397,N_19933,N_23979);
and U28398 (N_28398,N_20286,N_21728);
nor U28399 (N_28399,N_23495,N_23508);
or U28400 (N_28400,N_19842,N_23855);
and U28401 (N_28401,N_19487,N_22650);
xnor U28402 (N_28402,N_20432,N_21710);
nand U28403 (N_28403,N_18391,N_23391);
or U28404 (N_28404,N_19615,N_19595);
and U28405 (N_28405,N_23130,N_23274);
and U28406 (N_28406,N_20256,N_19392);
and U28407 (N_28407,N_20996,N_18709);
xor U28408 (N_28408,N_22942,N_18484);
xnor U28409 (N_28409,N_20561,N_19459);
and U28410 (N_28410,N_19687,N_20190);
nand U28411 (N_28411,N_19723,N_20514);
nor U28412 (N_28412,N_22082,N_18132);
nor U28413 (N_28413,N_23106,N_20940);
xor U28414 (N_28414,N_22104,N_22350);
nor U28415 (N_28415,N_19663,N_20883);
and U28416 (N_28416,N_21060,N_20128);
nor U28417 (N_28417,N_22712,N_22595);
nand U28418 (N_28418,N_19454,N_22151);
xor U28419 (N_28419,N_18532,N_23617);
and U28420 (N_28420,N_21379,N_23296);
nand U28421 (N_28421,N_18317,N_23482);
or U28422 (N_28422,N_18688,N_22737);
xor U28423 (N_28423,N_23394,N_22138);
nand U28424 (N_28424,N_20674,N_18547);
nor U28425 (N_28425,N_21651,N_18131);
or U28426 (N_28426,N_18782,N_19604);
nor U28427 (N_28427,N_21535,N_22002);
or U28428 (N_28428,N_22290,N_22434);
or U28429 (N_28429,N_21380,N_23526);
nand U28430 (N_28430,N_18008,N_22208);
and U28431 (N_28431,N_18182,N_21769);
and U28432 (N_28432,N_20355,N_22462);
or U28433 (N_28433,N_21876,N_23864);
nand U28434 (N_28434,N_20860,N_23663);
nand U28435 (N_28435,N_22643,N_23106);
or U28436 (N_28436,N_19945,N_23030);
nand U28437 (N_28437,N_19833,N_23330);
and U28438 (N_28438,N_20670,N_22869);
nand U28439 (N_28439,N_18187,N_19563);
or U28440 (N_28440,N_20704,N_19514);
or U28441 (N_28441,N_20666,N_22646);
xor U28442 (N_28442,N_21209,N_18596);
and U28443 (N_28443,N_22130,N_19284);
or U28444 (N_28444,N_18772,N_19295);
xor U28445 (N_28445,N_21075,N_19954);
or U28446 (N_28446,N_21720,N_22223);
xor U28447 (N_28447,N_23914,N_20316);
and U28448 (N_28448,N_19991,N_20084);
xor U28449 (N_28449,N_19864,N_20890);
nand U28450 (N_28450,N_19624,N_20434);
and U28451 (N_28451,N_19741,N_22904);
and U28452 (N_28452,N_18192,N_18842);
nor U28453 (N_28453,N_21501,N_23097);
nor U28454 (N_28454,N_21155,N_22269);
nand U28455 (N_28455,N_20217,N_23141);
or U28456 (N_28456,N_19440,N_21943);
nor U28457 (N_28457,N_23524,N_19315);
and U28458 (N_28458,N_22235,N_23510);
nand U28459 (N_28459,N_21595,N_20334);
nor U28460 (N_28460,N_23066,N_19571);
xor U28461 (N_28461,N_21236,N_21318);
nand U28462 (N_28462,N_22388,N_22780);
and U28463 (N_28463,N_18970,N_19718);
nor U28464 (N_28464,N_20421,N_19728);
nand U28465 (N_28465,N_22976,N_18642);
xnor U28466 (N_28466,N_23747,N_20962);
nor U28467 (N_28467,N_22102,N_19439);
nor U28468 (N_28468,N_22185,N_18135);
nand U28469 (N_28469,N_22067,N_20804);
xor U28470 (N_28470,N_23877,N_19989);
xor U28471 (N_28471,N_19273,N_22809);
and U28472 (N_28472,N_22614,N_20445);
nor U28473 (N_28473,N_23467,N_19056);
nand U28474 (N_28474,N_18185,N_20438);
and U28475 (N_28475,N_23523,N_23991);
nand U28476 (N_28476,N_23849,N_22941);
and U28477 (N_28477,N_20501,N_18376);
or U28478 (N_28478,N_21495,N_20987);
xnor U28479 (N_28479,N_21049,N_22367);
and U28480 (N_28480,N_21495,N_20995);
nor U28481 (N_28481,N_18550,N_20461);
and U28482 (N_28482,N_20632,N_20208);
xnor U28483 (N_28483,N_21535,N_21572);
or U28484 (N_28484,N_23736,N_22801);
and U28485 (N_28485,N_23484,N_22741);
xnor U28486 (N_28486,N_23035,N_19718);
xnor U28487 (N_28487,N_18788,N_22430);
xor U28488 (N_28488,N_19438,N_20111);
or U28489 (N_28489,N_20562,N_22674);
xor U28490 (N_28490,N_22972,N_21427);
nand U28491 (N_28491,N_18495,N_20831);
and U28492 (N_28492,N_22697,N_18271);
xor U28493 (N_28493,N_20970,N_18764);
nor U28494 (N_28494,N_22130,N_18138);
or U28495 (N_28495,N_19116,N_20925);
and U28496 (N_28496,N_21962,N_20810);
nor U28497 (N_28497,N_20630,N_20678);
nor U28498 (N_28498,N_23834,N_23239);
nor U28499 (N_28499,N_18904,N_23254);
or U28500 (N_28500,N_18658,N_23339);
and U28501 (N_28501,N_22661,N_18474);
xnor U28502 (N_28502,N_19246,N_21179);
and U28503 (N_28503,N_20899,N_22889);
xor U28504 (N_28504,N_22207,N_19117);
nor U28505 (N_28505,N_18414,N_23093);
xnor U28506 (N_28506,N_20467,N_20102);
or U28507 (N_28507,N_20083,N_20220);
and U28508 (N_28508,N_18044,N_23748);
or U28509 (N_28509,N_18489,N_19263);
xor U28510 (N_28510,N_23337,N_21292);
and U28511 (N_28511,N_19084,N_23732);
xnor U28512 (N_28512,N_18630,N_19378);
xor U28513 (N_28513,N_22940,N_22636);
xnor U28514 (N_28514,N_23570,N_21937);
nor U28515 (N_28515,N_19283,N_18734);
nor U28516 (N_28516,N_20336,N_20275);
and U28517 (N_28517,N_22902,N_23347);
nand U28518 (N_28518,N_19457,N_19925);
and U28519 (N_28519,N_22175,N_18569);
and U28520 (N_28520,N_21798,N_18822);
or U28521 (N_28521,N_23710,N_20824);
or U28522 (N_28522,N_18010,N_22761);
nand U28523 (N_28523,N_18916,N_22827);
nor U28524 (N_28524,N_23439,N_20057);
and U28525 (N_28525,N_23883,N_22524);
and U28526 (N_28526,N_22379,N_19897);
and U28527 (N_28527,N_18255,N_21468);
xnor U28528 (N_28528,N_18917,N_19807);
nand U28529 (N_28529,N_20874,N_21613);
and U28530 (N_28530,N_18806,N_18680);
or U28531 (N_28531,N_21095,N_19586);
nor U28532 (N_28532,N_21266,N_21874);
nand U28533 (N_28533,N_21547,N_18754);
nor U28534 (N_28534,N_19647,N_19060);
or U28535 (N_28535,N_21648,N_23589);
nor U28536 (N_28536,N_21680,N_23657);
nor U28537 (N_28537,N_18587,N_18495);
nor U28538 (N_28538,N_19423,N_20116);
nor U28539 (N_28539,N_20969,N_22251);
nand U28540 (N_28540,N_23669,N_21470);
and U28541 (N_28541,N_22780,N_19071);
nand U28542 (N_28542,N_23985,N_23628);
xnor U28543 (N_28543,N_20825,N_23652);
and U28544 (N_28544,N_22138,N_20684);
and U28545 (N_28545,N_23243,N_22003);
xnor U28546 (N_28546,N_23787,N_20780);
nand U28547 (N_28547,N_22516,N_21794);
nor U28548 (N_28548,N_21701,N_20435);
nor U28549 (N_28549,N_20601,N_18873);
or U28550 (N_28550,N_23466,N_18101);
and U28551 (N_28551,N_22602,N_18277);
or U28552 (N_28552,N_20252,N_18424);
and U28553 (N_28553,N_22209,N_19939);
nand U28554 (N_28554,N_19070,N_21472);
xor U28555 (N_28555,N_19030,N_23505);
or U28556 (N_28556,N_22103,N_19560);
or U28557 (N_28557,N_21723,N_23814);
or U28558 (N_28558,N_20043,N_23038);
nor U28559 (N_28559,N_22830,N_21692);
or U28560 (N_28560,N_21987,N_20607);
xor U28561 (N_28561,N_20856,N_18713);
nand U28562 (N_28562,N_20908,N_18604);
or U28563 (N_28563,N_23661,N_20248);
nand U28564 (N_28564,N_20360,N_21462);
and U28565 (N_28565,N_23251,N_22907);
nor U28566 (N_28566,N_21598,N_22124);
nand U28567 (N_28567,N_19357,N_22242);
xor U28568 (N_28568,N_18031,N_20721);
and U28569 (N_28569,N_18043,N_21896);
xnor U28570 (N_28570,N_18631,N_23464);
nor U28571 (N_28571,N_23546,N_21995);
nor U28572 (N_28572,N_19489,N_23621);
and U28573 (N_28573,N_22171,N_23768);
xor U28574 (N_28574,N_20004,N_20935);
or U28575 (N_28575,N_18158,N_20086);
nor U28576 (N_28576,N_21497,N_18925);
nand U28577 (N_28577,N_20443,N_20390);
and U28578 (N_28578,N_21178,N_22662);
nor U28579 (N_28579,N_18570,N_20880);
xor U28580 (N_28580,N_19722,N_21796);
nand U28581 (N_28581,N_22587,N_18656);
nand U28582 (N_28582,N_20340,N_19608);
and U28583 (N_28583,N_23382,N_19305);
nor U28584 (N_28584,N_21704,N_19355);
nor U28585 (N_28585,N_21664,N_18395);
or U28586 (N_28586,N_20801,N_20435);
nand U28587 (N_28587,N_23051,N_19751);
nand U28588 (N_28588,N_23841,N_18563);
nand U28589 (N_28589,N_22479,N_20406);
nand U28590 (N_28590,N_21366,N_23024);
nand U28591 (N_28591,N_21790,N_21017);
nand U28592 (N_28592,N_18449,N_21936);
xnor U28593 (N_28593,N_18758,N_23288);
or U28594 (N_28594,N_23461,N_20006);
nor U28595 (N_28595,N_22689,N_23314);
and U28596 (N_28596,N_19023,N_22960);
nor U28597 (N_28597,N_23015,N_23582);
or U28598 (N_28598,N_19434,N_21459);
and U28599 (N_28599,N_23881,N_21321);
nor U28600 (N_28600,N_20571,N_18093);
xor U28601 (N_28601,N_18541,N_18846);
nor U28602 (N_28602,N_21711,N_18228);
and U28603 (N_28603,N_22333,N_22234);
and U28604 (N_28604,N_19405,N_22713);
and U28605 (N_28605,N_21493,N_18088);
and U28606 (N_28606,N_20944,N_19256);
nor U28607 (N_28607,N_19684,N_21890);
or U28608 (N_28608,N_22809,N_23529);
nor U28609 (N_28609,N_18451,N_21529);
or U28610 (N_28610,N_19727,N_23474);
and U28611 (N_28611,N_21832,N_18867);
or U28612 (N_28612,N_23189,N_21466);
xnor U28613 (N_28613,N_22368,N_23799);
nor U28614 (N_28614,N_19839,N_23320);
and U28615 (N_28615,N_22289,N_23540);
nand U28616 (N_28616,N_20402,N_21729);
nand U28617 (N_28617,N_18043,N_20097);
and U28618 (N_28618,N_20031,N_20892);
xnor U28619 (N_28619,N_21875,N_19619);
nor U28620 (N_28620,N_19186,N_22376);
and U28621 (N_28621,N_21754,N_19973);
and U28622 (N_28622,N_20671,N_21392);
or U28623 (N_28623,N_20201,N_20809);
nor U28624 (N_28624,N_22076,N_18401);
nor U28625 (N_28625,N_21046,N_23517);
nor U28626 (N_28626,N_23818,N_18468);
and U28627 (N_28627,N_19505,N_20678);
nor U28628 (N_28628,N_20665,N_22285);
or U28629 (N_28629,N_21271,N_21022);
or U28630 (N_28630,N_18725,N_21373);
nor U28631 (N_28631,N_20886,N_18301);
and U28632 (N_28632,N_19645,N_19652);
or U28633 (N_28633,N_20014,N_20026);
nor U28634 (N_28634,N_23169,N_22660);
xnor U28635 (N_28635,N_23944,N_22117);
or U28636 (N_28636,N_20152,N_20200);
xor U28637 (N_28637,N_21292,N_18017);
or U28638 (N_28638,N_18099,N_18810);
nor U28639 (N_28639,N_21153,N_19786);
nand U28640 (N_28640,N_21609,N_22014);
or U28641 (N_28641,N_18765,N_22317);
and U28642 (N_28642,N_21514,N_23581);
or U28643 (N_28643,N_23969,N_22793);
and U28644 (N_28644,N_19201,N_21809);
xor U28645 (N_28645,N_18110,N_21594);
nand U28646 (N_28646,N_18650,N_22921);
and U28647 (N_28647,N_22691,N_18799);
nor U28648 (N_28648,N_21206,N_22238);
and U28649 (N_28649,N_19248,N_20607);
nand U28650 (N_28650,N_22731,N_18730);
nand U28651 (N_28651,N_20005,N_23305);
nor U28652 (N_28652,N_23683,N_22592);
xor U28653 (N_28653,N_23015,N_21373);
nor U28654 (N_28654,N_21682,N_20415);
or U28655 (N_28655,N_18004,N_22978);
nor U28656 (N_28656,N_23254,N_19120);
and U28657 (N_28657,N_18809,N_21990);
or U28658 (N_28658,N_19324,N_22980);
nand U28659 (N_28659,N_19474,N_21092);
and U28660 (N_28660,N_23636,N_22280);
xor U28661 (N_28661,N_19102,N_23049);
xor U28662 (N_28662,N_20161,N_19462);
and U28663 (N_28663,N_20953,N_20798);
nand U28664 (N_28664,N_22053,N_21482);
xor U28665 (N_28665,N_21015,N_22581);
nor U28666 (N_28666,N_20690,N_23098);
xnor U28667 (N_28667,N_22409,N_23789);
xnor U28668 (N_28668,N_23594,N_23354);
nor U28669 (N_28669,N_21959,N_23218);
nor U28670 (N_28670,N_18379,N_22066);
xor U28671 (N_28671,N_21321,N_23956);
and U28672 (N_28672,N_20150,N_18299);
and U28673 (N_28673,N_18262,N_23763);
or U28674 (N_28674,N_21128,N_23872);
or U28675 (N_28675,N_20028,N_19573);
xor U28676 (N_28676,N_22108,N_20546);
nor U28677 (N_28677,N_22645,N_23619);
nor U28678 (N_28678,N_19018,N_22891);
nand U28679 (N_28679,N_20977,N_23432);
nor U28680 (N_28680,N_20554,N_19640);
xor U28681 (N_28681,N_19077,N_18650);
xor U28682 (N_28682,N_19425,N_18793);
or U28683 (N_28683,N_19178,N_19789);
xnor U28684 (N_28684,N_21592,N_23620);
nor U28685 (N_28685,N_23751,N_22455);
nand U28686 (N_28686,N_21039,N_18145);
or U28687 (N_28687,N_21292,N_21923);
or U28688 (N_28688,N_21429,N_23579);
nor U28689 (N_28689,N_21048,N_22397);
and U28690 (N_28690,N_19831,N_22183);
nor U28691 (N_28691,N_22111,N_23785);
xnor U28692 (N_28692,N_21550,N_20813);
xor U28693 (N_28693,N_19671,N_23881);
or U28694 (N_28694,N_20710,N_20951);
xnor U28695 (N_28695,N_21987,N_19501);
nor U28696 (N_28696,N_18897,N_18919);
or U28697 (N_28697,N_19416,N_21021);
nand U28698 (N_28698,N_23613,N_19419);
or U28699 (N_28699,N_22703,N_20590);
nand U28700 (N_28700,N_19391,N_22279);
and U28701 (N_28701,N_18890,N_20286);
xor U28702 (N_28702,N_19317,N_20509);
or U28703 (N_28703,N_18235,N_21266);
nor U28704 (N_28704,N_23793,N_22834);
nor U28705 (N_28705,N_19829,N_18559);
or U28706 (N_28706,N_20937,N_19394);
and U28707 (N_28707,N_20968,N_22577);
and U28708 (N_28708,N_20464,N_18260);
xor U28709 (N_28709,N_22165,N_19301);
xnor U28710 (N_28710,N_18484,N_20030);
and U28711 (N_28711,N_21379,N_19240);
nand U28712 (N_28712,N_23711,N_22943);
nand U28713 (N_28713,N_18359,N_18458);
and U28714 (N_28714,N_18007,N_21842);
nor U28715 (N_28715,N_23359,N_20728);
nor U28716 (N_28716,N_20884,N_22394);
nor U28717 (N_28717,N_22402,N_20744);
or U28718 (N_28718,N_23868,N_20319);
xnor U28719 (N_28719,N_18655,N_23112);
nor U28720 (N_28720,N_19669,N_23624);
xor U28721 (N_28721,N_22431,N_22533);
nor U28722 (N_28722,N_22258,N_19323);
nor U28723 (N_28723,N_19735,N_22142);
and U28724 (N_28724,N_20672,N_22132);
or U28725 (N_28725,N_18183,N_22974);
and U28726 (N_28726,N_21199,N_19838);
nand U28727 (N_28727,N_21360,N_21634);
xor U28728 (N_28728,N_19729,N_18088);
nand U28729 (N_28729,N_18248,N_23179);
xnor U28730 (N_28730,N_21970,N_18491);
xnor U28731 (N_28731,N_19251,N_20263);
or U28732 (N_28732,N_20268,N_19257);
nand U28733 (N_28733,N_20592,N_21550);
and U28734 (N_28734,N_22650,N_18583);
nor U28735 (N_28735,N_20342,N_21301);
nor U28736 (N_28736,N_23447,N_19952);
and U28737 (N_28737,N_21044,N_18938);
nor U28738 (N_28738,N_20456,N_21793);
xnor U28739 (N_28739,N_18470,N_19696);
or U28740 (N_28740,N_22744,N_18776);
xor U28741 (N_28741,N_19002,N_23863);
or U28742 (N_28742,N_20228,N_19228);
nor U28743 (N_28743,N_20600,N_21470);
and U28744 (N_28744,N_19994,N_20896);
nor U28745 (N_28745,N_20847,N_22759);
nor U28746 (N_28746,N_19439,N_20925);
and U28747 (N_28747,N_23476,N_21324);
nand U28748 (N_28748,N_23830,N_19017);
nand U28749 (N_28749,N_22145,N_19624);
or U28750 (N_28750,N_23017,N_20228);
nand U28751 (N_28751,N_20956,N_23356);
xnor U28752 (N_28752,N_21126,N_18878);
or U28753 (N_28753,N_19346,N_22162);
nand U28754 (N_28754,N_23933,N_21351);
or U28755 (N_28755,N_18731,N_20731);
and U28756 (N_28756,N_22412,N_21845);
and U28757 (N_28757,N_22087,N_22922);
nor U28758 (N_28758,N_19610,N_19882);
nand U28759 (N_28759,N_20109,N_21949);
or U28760 (N_28760,N_18380,N_18895);
xor U28761 (N_28761,N_23946,N_23182);
nor U28762 (N_28762,N_23715,N_20865);
nor U28763 (N_28763,N_23754,N_18261);
or U28764 (N_28764,N_19578,N_21771);
xnor U28765 (N_28765,N_22516,N_22903);
xor U28766 (N_28766,N_21001,N_20132);
and U28767 (N_28767,N_19248,N_22773);
and U28768 (N_28768,N_20166,N_23176);
xnor U28769 (N_28769,N_22143,N_18108);
or U28770 (N_28770,N_18982,N_23109);
and U28771 (N_28771,N_18349,N_19702);
nand U28772 (N_28772,N_22058,N_23501);
or U28773 (N_28773,N_20083,N_23106);
xnor U28774 (N_28774,N_18712,N_19633);
nand U28775 (N_28775,N_23292,N_19562);
nand U28776 (N_28776,N_23654,N_18653);
and U28777 (N_28777,N_20250,N_19165);
nand U28778 (N_28778,N_21068,N_19690);
xor U28779 (N_28779,N_19023,N_18540);
nor U28780 (N_28780,N_23741,N_23853);
or U28781 (N_28781,N_20546,N_18663);
nand U28782 (N_28782,N_19477,N_18555);
xnor U28783 (N_28783,N_23512,N_20284);
xor U28784 (N_28784,N_19143,N_21040);
xnor U28785 (N_28785,N_22832,N_20582);
nand U28786 (N_28786,N_22561,N_22018);
nand U28787 (N_28787,N_23073,N_22764);
nand U28788 (N_28788,N_19847,N_20333);
and U28789 (N_28789,N_20551,N_19732);
nand U28790 (N_28790,N_22178,N_19739);
nand U28791 (N_28791,N_22457,N_20130);
nand U28792 (N_28792,N_21666,N_23936);
xnor U28793 (N_28793,N_19124,N_20535);
and U28794 (N_28794,N_23835,N_23525);
or U28795 (N_28795,N_18585,N_22855);
nor U28796 (N_28796,N_18696,N_22720);
or U28797 (N_28797,N_21674,N_18482);
or U28798 (N_28798,N_18947,N_23835);
and U28799 (N_28799,N_19796,N_23502);
xor U28800 (N_28800,N_18644,N_20080);
xnor U28801 (N_28801,N_18231,N_21987);
or U28802 (N_28802,N_18111,N_19822);
or U28803 (N_28803,N_21678,N_19602);
xnor U28804 (N_28804,N_21736,N_22402);
nand U28805 (N_28805,N_22073,N_23683);
nand U28806 (N_28806,N_20664,N_23811);
nor U28807 (N_28807,N_18839,N_22905);
and U28808 (N_28808,N_23653,N_22811);
nor U28809 (N_28809,N_23355,N_19230);
nor U28810 (N_28810,N_23473,N_19634);
or U28811 (N_28811,N_18557,N_22043);
or U28812 (N_28812,N_22453,N_23073);
nand U28813 (N_28813,N_19237,N_21736);
nor U28814 (N_28814,N_22719,N_23549);
and U28815 (N_28815,N_18038,N_21688);
nand U28816 (N_28816,N_23614,N_19867);
nor U28817 (N_28817,N_18394,N_23755);
nand U28818 (N_28818,N_22567,N_22895);
nor U28819 (N_28819,N_23694,N_20522);
and U28820 (N_28820,N_19172,N_22310);
or U28821 (N_28821,N_23563,N_18518);
nand U28822 (N_28822,N_20627,N_23970);
or U28823 (N_28823,N_22595,N_18505);
nor U28824 (N_28824,N_23698,N_18511);
and U28825 (N_28825,N_18441,N_21760);
and U28826 (N_28826,N_20245,N_23995);
or U28827 (N_28827,N_21463,N_20460);
nor U28828 (N_28828,N_20938,N_20092);
nand U28829 (N_28829,N_20756,N_20747);
nand U28830 (N_28830,N_23165,N_20085);
xor U28831 (N_28831,N_22396,N_19176);
or U28832 (N_28832,N_22835,N_22220);
or U28833 (N_28833,N_23259,N_18938);
xor U28834 (N_28834,N_18396,N_21573);
or U28835 (N_28835,N_21221,N_18270);
and U28836 (N_28836,N_18217,N_23304);
or U28837 (N_28837,N_19175,N_22680);
xor U28838 (N_28838,N_23931,N_23187);
nor U28839 (N_28839,N_19604,N_23445);
xnor U28840 (N_28840,N_21079,N_19176);
nor U28841 (N_28841,N_22172,N_18546);
and U28842 (N_28842,N_20393,N_19097);
and U28843 (N_28843,N_23368,N_22692);
and U28844 (N_28844,N_18176,N_22435);
and U28845 (N_28845,N_20330,N_23996);
nor U28846 (N_28846,N_22539,N_20397);
nand U28847 (N_28847,N_23684,N_23372);
and U28848 (N_28848,N_18619,N_23088);
or U28849 (N_28849,N_23585,N_20567);
nand U28850 (N_28850,N_18827,N_18537);
nor U28851 (N_28851,N_20534,N_19586);
or U28852 (N_28852,N_21994,N_18650);
nor U28853 (N_28853,N_19378,N_21342);
and U28854 (N_28854,N_18371,N_23611);
xor U28855 (N_28855,N_21137,N_23451);
or U28856 (N_28856,N_19192,N_20176);
and U28857 (N_28857,N_22829,N_23856);
or U28858 (N_28858,N_19634,N_21532);
nand U28859 (N_28859,N_18694,N_20057);
nor U28860 (N_28860,N_20553,N_20175);
or U28861 (N_28861,N_18953,N_22821);
nand U28862 (N_28862,N_21781,N_20474);
or U28863 (N_28863,N_22205,N_19300);
xor U28864 (N_28864,N_20127,N_22045);
xor U28865 (N_28865,N_19889,N_21270);
and U28866 (N_28866,N_21182,N_22265);
xnor U28867 (N_28867,N_21366,N_19788);
xor U28868 (N_28868,N_20888,N_23811);
and U28869 (N_28869,N_20935,N_22563);
xnor U28870 (N_28870,N_23116,N_20243);
nand U28871 (N_28871,N_22684,N_20669);
nor U28872 (N_28872,N_22826,N_18219);
nand U28873 (N_28873,N_21250,N_18299);
or U28874 (N_28874,N_20632,N_18950);
and U28875 (N_28875,N_22248,N_19676);
nor U28876 (N_28876,N_18453,N_23667);
nor U28877 (N_28877,N_20625,N_23952);
xor U28878 (N_28878,N_19867,N_22675);
and U28879 (N_28879,N_21461,N_20893);
and U28880 (N_28880,N_22291,N_23105);
and U28881 (N_28881,N_19476,N_18204);
nor U28882 (N_28882,N_22622,N_19525);
and U28883 (N_28883,N_19351,N_18044);
nand U28884 (N_28884,N_18155,N_18415);
and U28885 (N_28885,N_21876,N_19982);
nor U28886 (N_28886,N_23852,N_20148);
nor U28887 (N_28887,N_19147,N_23259);
xnor U28888 (N_28888,N_22564,N_20740);
nand U28889 (N_28889,N_19916,N_18207);
nand U28890 (N_28890,N_20527,N_22015);
or U28891 (N_28891,N_20178,N_22187);
nor U28892 (N_28892,N_19380,N_20158);
xor U28893 (N_28893,N_22348,N_19039);
or U28894 (N_28894,N_21919,N_22312);
or U28895 (N_28895,N_18589,N_21517);
or U28896 (N_28896,N_22418,N_23239);
and U28897 (N_28897,N_18298,N_23795);
and U28898 (N_28898,N_20851,N_23837);
xnor U28899 (N_28899,N_20401,N_18972);
and U28900 (N_28900,N_19468,N_18396);
or U28901 (N_28901,N_23113,N_20863);
nand U28902 (N_28902,N_19962,N_18738);
xnor U28903 (N_28903,N_22467,N_20779);
xor U28904 (N_28904,N_19069,N_18925);
nor U28905 (N_28905,N_19522,N_20894);
xnor U28906 (N_28906,N_20193,N_23476);
and U28907 (N_28907,N_23931,N_23996);
and U28908 (N_28908,N_19682,N_22881);
or U28909 (N_28909,N_19648,N_22933);
nand U28910 (N_28910,N_19256,N_21887);
and U28911 (N_28911,N_20408,N_20502);
nor U28912 (N_28912,N_21775,N_20299);
nor U28913 (N_28913,N_18101,N_19781);
and U28914 (N_28914,N_20783,N_23829);
and U28915 (N_28915,N_20354,N_21365);
and U28916 (N_28916,N_21372,N_20366);
xnor U28917 (N_28917,N_22696,N_22874);
nand U28918 (N_28918,N_20446,N_22560);
nand U28919 (N_28919,N_21196,N_20756);
nor U28920 (N_28920,N_21528,N_20446);
and U28921 (N_28921,N_18494,N_23001);
or U28922 (N_28922,N_19172,N_21429);
nand U28923 (N_28923,N_18266,N_20414);
xnor U28924 (N_28924,N_23527,N_19558);
and U28925 (N_28925,N_22437,N_23173);
nand U28926 (N_28926,N_23564,N_21806);
nor U28927 (N_28927,N_23287,N_22878);
nor U28928 (N_28928,N_18168,N_22322);
nand U28929 (N_28929,N_21248,N_21204);
xnor U28930 (N_28930,N_19321,N_22467);
xor U28931 (N_28931,N_22367,N_18443);
xor U28932 (N_28932,N_23374,N_18469);
xnor U28933 (N_28933,N_18686,N_20475);
or U28934 (N_28934,N_18101,N_19683);
or U28935 (N_28935,N_21508,N_18662);
xor U28936 (N_28936,N_21515,N_20084);
nor U28937 (N_28937,N_18945,N_18743);
and U28938 (N_28938,N_21111,N_20731);
nor U28939 (N_28939,N_20613,N_20150);
nand U28940 (N_28940,N_18702,N_19169);
nor U28941 (N_28941,N_18348,N_23373);
nor U28942 (N_28942,N_19397,N_20066);
xnor U28943 (N_28943,N_21158,N_22959);
nand U28944 (N_28944,N_18707,N_18353);
or U28945 (N_28945,N_20840,N_20549);
xor U28946 (N_28946,N_20728,N_21504);
and U28947 (N_28947,N_20083,N_20598);
and U28948 (N_28948,N_20170,N_22920);
xor U28949 (N_28949,N_23807,N_18754);
nand U28950 (N_28950,N_20283,N_18474);
and U28951 (N_28951,N_18142,N_23700);
and U28952 (N_28952,N_21442,N_18624);
nand U28953 (N_28953,N_20147,N_21713);
or U28954 (N_28954,N_18283,N_21555);
nand U28955 (N_28955,N_22662,N_20854);
and U28956 (N_28956,N_23351,N_21710);
nor U28957 (N_28957,N_21461,N_21510);
nor U28958 (N_28958,N_23272,N_20927);
xnor U28959 (N_28959,N_23302,N_22135);
or U28960 (N_28960,N_19086,N_23297);
or U28961 (N_28961,N_19897,N_20601);
or U28962 (N_28962,N_18736,N_18381);
nor U28963 (N_28963,N_19962,N_20902);
or U28964 (N_28964,N_18364,N_21627);
and U28965 (N_28965,N_19488,N_22724);
or U28966 (N_28966,N_18116,N_22138);
and U28967 (N_28967,N_20071,N_18203);
nor U28968 (N_28968,N_23684,N_22677);
nand U28969 (N_28969,N_23099,N_18314);
nand U28970 (N_28970,N_23524,N_18652);
nor U28971 (N_28971,N_19641,N_21097);
xnor U28972 (N_28972,N_23750,N_18236);
or U28973 (N_28973,N_18535,N_19794);
or U28974 (N_28974,N_19642,N_23542);
nor U28975 (N_28975,N_20943,N_19054);
xnor U28976 (N_28976,N_19943,N_22176);
xor U28977 (N_28977,N_22861,N_18303);
nand U28978 (N_28978,N_18586,N_20375);
or U28979 (N_28979,N_23585,N_19993);
and U28980 (N_28980,N_20996,N_23794);
or U28981 (N_28981,N_20210,N_19743);
or U28982 (N_28982,N_19935,N_23471);
xor U28983 (N_28983,N_21747,N_22845);
and U28984 (N_28984,N_21975,N_22826);
nor U28985 (N_28985,N_20298,N_22834);
nor U28986 (N_28986,N_22479,N_18338);
or U28987 (N_28987,N_22836,N_20907);
or U28988 (N_28988,N_22859,N_22977);
or U28989 (N_28989,N_21651,N_23984);
xnor U28990 (N_28990,N_18379,N_20473);
nand U28991 (N_28991,N_23184,N_18032);
nor U28992 (N_28992,N_20161,N_18830);
and U28993 (N_28993,N_22598,N_21906);
xnor U28994 (N_28994,N_20898,N_23227);
or U28995 (N_28995,N_21445,N_22045);
nand U28996 (N_28996,N_18437,N_19987);
and U28997 (N_28997,N_20900,N_23308);
xnor U28998 (N_28998,N_23241,N_18067);
or U28999 (N_28999,N_20332,N_18480);
or U29000 (N_29000,N_23966,N_19903);
xnor U29001 (N_29001,N_22259,N_22331);
xor U29002 (N_29002,N_21777,N_22629);
nand U29003 (N_29003,N_22860,N_21096);
nor U29004 (N_29004,N_23939,N_20392);
and U29005 (N_29005,N_22022,N_19269);
xnor U29006 (N_29006,N_21170,N_23027);
or U29007 (N_29007,N_20732,N_19769);
xnor U29008 (N_29008,N_19211,N_18708);
xnor U29009 (N_29009,N_23826,N_19025);
nor U29010 (N_29010,N_23093,N_22279);
or U29011 (N_29011,N_23738,N_21165);
nand U29012 (N_29012,N_23394,N_23196);
nand U29013 (N_29013,N_20907,N_23909);
nand U29014 (N_29014,N_22086,N_18737);
or U29015 (N_29015,N_21678,N_22750);
nor U29016 (N_29016,N_23634,N_23266);
and U29017 (N_29017,N_21969,N_20875);
nor U29018 (N_29018,N_23797,N_18274);
xnor U29019 (N_29019,N_21901,N_19253);
xnor U29020 (N_29020,N_20539,N_21167);
or U29021 (N_29021,N_19260,N_20053);
nand U29022 (N_29022,N_23854,N_20627);
nor U29023 (N_29023,N_19415,N_23340);
and U29024 (N_29024,N_21155,N_23381);
or U29025 (N_29025,N_21749,N_21024);
nor U29026 (N_29026,N_18942,N_19977);
nor U29027 (N_29027,N_18596,N_18515);
nand U29028 (N_29028,N_22994,N_18931);
nor U29029 (N_29029,N_22986,N_18212);
nor U29030 (N_29030,N_19047,N_22224);
xor U29031 (N_29031,N_22604,N_23244);
or U29032 (N_29032,N_18822,N_19192);
xnor U29033 (N_29033,N_18390,N_20141);
xnor U29034 (N_29034,N_21725,N_21108);
and U29035 (N_29035,N_18552,N_19931);
xor U29036 (N_29036,N_21072,N_21668);
and U29037 (N_29037,N_22479,N_23045);
and U29038 (N_29038,N_21670,N_20491);
xnor U29039 (N_29039,N_20745,N_20008);
or U29040 (N_29040,N_18546,N_22865);
nor U29041 (N_29041,N_23984,N_20010);
or U29042 (N_29042,N_23310,N_18341);
xnor U29043 (N_29043,N_19616,N_21779);
or U29044 (N_29044,N_21416,N_19416);
and U29045 (N_29045,N_20657,N_20642);
and U29046 (N_29046,N_21179,N_20414);
xnor U29047 (N_29047,N_18265,N_18609);
and U29048 (N_29048,N_20045,N_23488);
xnor U29049 (N_29049,N_22391,N_22982);
or U29050 (N_29050,N_23051,N_18085);
xnor U29051 (N_29051,N_23851,N_20077);
nor U29052 (N_29052,N_20856,N_23565);
or U29053 (N_29053,N_23755,N_19572);
xnor U29054 (N_29054,N_21446,N_22564);
nand U29055 (N_29055,N_18786,N_18909);
nor U29056 (N_29056,N_22840,N_23786);
nor U29057 (N_29057,N_19623,N_23298);
or U29058 (N_29058,N_21018,N_20429);
nand U29059 (N_29059,N_21330,N_21694);
or U29060 (N_29060,N_22580,N_18559);
nand U29061 (N_29061,N_20536,N_20410);
xnor U29062 (N_29062,N_23091,N_23697);
or U29063 (N_29063,N_18030,N_21758);
xor U29064 (N_29064,N_22510,N_23668);
nor U29065 (N_29065,N_18667,N_19922);
xor U29066 (N_29066,N_23148,N_22076);
or U29067 (N_29067,N_20798,N_19415);
xnor U29068 (N_29068,N_18001,N_23399);
and U29069 (N_29069,N_18706,N_18084);
nand U29070 (N_29070,N_23840,N_20869);
xnor U29071 (N_29071,N_21979,N_18367);
xnor U29072 (N_29072,N_20190,N_19289);
nor U29073 (N_29073,N_22723,N_23480);
nor U29074 (N_29074,N_18352,N_19175);
nor U29075 (N_29075,N_22785,N_22100);
xnor U29076 (N_29076,N_18235,N_19444);
and U29077 (N_29077,N_23150,N_22700);
or U29078 (N_29078,N_21442,N_21591);
and U29079 (N_29079,N_21794,N_23171);
or U29080 (N_29080,N_19483,N_18353);
and U29081 (N_29081,N_22457,N_23951);
xnor U29082 (N_29082,N_21623,N_21245);
xnor U29083 (N_29083,N_23514,N_19592);
and U29084 (N_29084,N_21936,N_19698);
nor U29085 (N_29085,N_18726,N_19613);
nor U29086 (N_29086,N_22533,N_19731);
nor U29087 (N_29087,N_23500,N_21036);
and U29088 (N_29088,N_23460,N_21430);
nor U29089 (N_29089,N_23190,N_18774);
and U29090 (N_29090,N_19938,N_21927);
nand U29091 (N_29091,N_21548,N_22187);
xor U29092 (N_29092,N_22966,N_19277);
nor U29093 (N_29093,N_21686,N_21188);
nor U29094 (N_29094,N_20360,N_18299);
and U29095 (N_29095,N_18330,N_21626);
nand U29096 (N_29096,N_22243,N_21494);
and U29097 (N_29097,N_19305,N_22226);
and U29098 (N_29098,N_23786,N_22619);
and U29099 (N_29099,N_19206,N_21929);
nor U29100 (N_29100,N_19450,N_18834);
and U29101 (N_29101,N_22191,N_20302);
nor U29102 (N_29102,N_19212,N_23715);
nand U29103 (N_29103,N_22387,N_18386);
nor U29104 (N_29104,N_19826,N_22267);
xnor U29105 (N_29105,N_21860,N_22755);
and U29106 (N_29106,N_23478,N_21985);
xor U29107 (N_29107,N_18407,N_22063);
and U29108 (N_29108,N_20180,N_18113);
or U29109 (N_29109,N_22007,N_18095);
nor U29110 (N_29110,N_21956,N_20937);
or U29111 (N_29111,N_19513,N_23070);
xnor U29112 (N_29112,N_21939,N_18250);
and U29113 (N_29113,N_19663,N_23356);
and U29114 (N_29114,N_20415,N_20467);
and U29115 (N_29115,N_21569,N_21779);
nand U29116 (N_29116,N_23759,N_22350);
nand U29117 (N_29117,N_20427,N_18511);
xnor U29118 (N_29118,N_22034,N_23528);
xor U29119 (N_29119,N_21779,N_21999);
xnor U29120 (N_29120,N_21117,N_22346);
nor U29121 (N_29121,N_22066,N_18000);
xor U29122 (N_29122,N_22680,N_18894);
xnor U29123 (N_29123,N_20085,N_22643);
xnor U29124 (N_29124,N_23191,N_19202);
nand U29125 (N_29125,N_21968,N_20361);
or U29126 (N_29126,N_20127,N_21316);
and U29127 (N_29127,N_19741,N_19221);
xnor U29128 (N_29128,N_22346,N_22602);
xor U29129 (N_29129,N_21319,N_19862);
nor U29130 (N_29130,N_22755,N_22593);
nand U29131 (N_29131,N_22899,N_21411);
xor U29132 (N_29132,N_18781,N_18998);
or U29133 (N_29133,N_20168,N_18379);
xor U29134 (N_29134,N_19956,N_23713);
and U29135 (N_29135,N_19499,N_19596);
or U29136 (N_29136,N_18728,N_20998);
nor U29137 (N_29137,N_23483,N_23449);
xnor U29138 (N_29138,N_19485,N_23870);
xor U29139 (N_29139,N_23496,N_18642);
or U29140 (N_29140,N_23286,N_22935);
and U29141 (N_29141,N_20317,N_22678);
or U29142 (N_29142,N_19485,N_19092);
and U29143 (N_29143,N_21980,N_18476);
or U29144 (N_29144,N_19698,N_23213);
nand U29145 (N_29145,N_18174,N_22927);
or U29146 (N_29146,N_18897,N_19164);
and U29147 (N_29147,N_19643,N_19023);
or U29148 (N_29148,N_23133,N_22132);
xnor U29149 (N_29149,N_21297,N_22963);
and U29150 (N_29150,N_21281,N_18688);
nand U29151 (N_29151,N_21134,N_21082);
nor U29152 (N_29152,N_23226,N_19165);
nor U29153 (N_29153,N_22223,N_21916);
and U29154 (N_29154,N_21432,N_18222);
nor U29155 (N_29155,N_22556,N_22032);
nand U29156 (N_29156,N_22856,N_22292);
xnor U29157 (N_29157,N_18645,N_21123);
xor U29158 (N_29158,N_23141,N_21817);
nand U29159 (N_29159,N_22000,N_19781);
or U29160 (N_29160,N_20631,N_20689);
or U29161 (N_29161,N_19457,N_19389);
and U29162 (N_29162,N_22371,N_23230);
or U29163 (N_29163,N_20139,N_18837);
and U29164 (N_29164,N_23362,N_23777);
or U29165 (N_29165,N_18881,N_21149);
or U29166 (N_29166,N_20830,N_21231);
nor U29167 (N_29167,N_19175,N_23909);
nor U29168 (N_29168,N_23628,N_21067);
and U29169 (N_29169,N_23974,N_23320);
and U29170 (N_29170,N_20646,N_23370);
and U29171 (N_29171,N_19914,N_21363);
or U29172 (N_29172,N_22053,N_21674);
or U29173 (N_29173,N_21807,N_19703);
nand U29174 (N_29174,N_18449,N_22697);
xnor U29175 (N_29175,N_23646,N_23661);
xor U29176 (N_29176,N_22391,N_23663);
and U29177 (N_29177,N_18024,N_23431);
and U29178 (N_29178,N_22231,N_20082);
nand U29179 (N_29179,N_23521,N_23554);
xor U29180 (N_29180,N_21617,N_21042);
xnor U29181 (N_29181,N_22558,N_18218);
nand U29182 (N_29182,N_19545,N_21096);
and U29183 (N_29183,N_22673,N_21437);
or U29184 (N_29184,N_18115,N_21598);
and U29185 (N_29185,N_19047,N_22297);
xor U29186 (N_29186,N_19090,N_19239);
nor U29187 (N_29187,N_19620,N_21518);
xor U29188 (N_29188,N_20700,N_21287);
xnor U29189 (N_29189,N_21861,N_22628);
and U29190 (N_29190,N_18846,N_22440);
nand U29191 (N_29191,N_22149,N_20542);
or U29192 (N_29192,N_23033,N_22002);
nor U29193 (N_29193,N_19331,N_19552);
nor U29194 (N_29194,N_20368,N_22106);
nor U29195 (N_29195,N_19834,N_20931);
nor U29196 (N_29196,N_21631,N_18740);
nor U29197 (N_29197,N_18763,N_18776);
nor U29198 (N_29198,N_22745,N_20371);
and U29199 (N_29199,N_19429,N_18842);
and U29200 (N_29200,N_20664,N_21522);
xor U29201 (N_29201,N_23302,N_18819);
or U29202 (N_29202,N_23690,N_18463);
nand U29203 (N_29203,N_19354,N_19789);
xnor U29204 (N_29204,N_19874,N_23668);
xnor U29205 (N_29205,N_23184,N_20659);
xnor U29206 (N_29206,N_23870,N_20074);
nor U29207 (N_29207,N_21692,N_18844);
xor U29208 (N_29208,N_23107,N_19782);
nand U29209 (N_29209,N_23449,N_19793);
xnor U29210 (N_29210,N_18407,N_21140);
xor U29211 (N_29211,N_19523,N_21930);
xor U29212 (N_29212,N_20761,N_18539);
and U29213 (N_29213,N_20782,N_23799);
and U29214 (N_29214,N_20142,N_20689);
or U29215 (N_29215,N_19709,N_22949);
and U29216 (N_29216,N_20961,N_18144);
xnor U29217 (N_29217,N_23501,N_20993);
nor U29218 (N_29218,N_21437,N_19434);
and U29219 (N_29219,N_18567,N_19262);
or U29220 (N_29220,N_19947,N_21371);
nor U29221 (N_29221,N_19659,N_20669);
nor U29222 (N_29222,N_21927,N_20145);
xnor U29223 (N_29223,N_20167,N_21249);
nand U29224 (N_29224,N_18202,N_20392);
or U29225 (N_29225,N_20012,N_23247);
xor U29226 (N_29226,N_19953,N_22097);
xor U29227 (N_29227,N_22423,N_19333);
or U29228 (N_29228,N_23117,N_18936);
nor U29229 (N_29229,N_19792,N_20999);
or U29230 (N_29230,N_18471,N_21993);
nand U29231 (N_29231,N_20247,N_20603);
or U29232 (N_29232,N_23169,N_22318);
or U29233 (N_29233,N_20898,N_22076);
xor U29234 (N_29234,N_23246,N_22006);
nor U29235 (N_29235,N_21421,N_23172);
nand U29236 (N_29236,N_19792,N_22354);
xnor U29237 (N_29237,N_19387,N_19373);
or U29238 (N_29238,N_18869,N_18219);
nor U29239 (N_29239,N_18975,N_21311);
xor U29240 (N_29240,N_21353,N_23613);
xor U29241 (N_29241,N_21615,N_21089);
or U29242 (N_29242,N_19131,N_23776);
and U29243 (N_29243,N_22503,N_22608);
xnor U29244 (N_29244,N_19004,N_19522);
nor U29245 (N_29245,N_19046,N_18798);
nand U29246 (N_29246,N_18536,N_22247);
nor U29247 (N_29247,N_20791,N_20215);
xnor U29248 (N_29248,N_20147,N_20030);
or U29249 (N_29249,N_19987,N_22682);
nor U29250 (N_29250,N_18093,N_18432);
and U29251 (N_29251,N_22086,N_21190);
xnor U29252 (N_29252,N_22683,N_19445);
nor U29253 (N_29253,N_20361,N_19674);
nor U29254 (N_29254,N_21645,N_20632);
nor U29255 (N_29255,N_18937,N_22190);
xnor U29256 (N_29256,N_22911,N_23759);
xor U29257 (N_29257,N_22573,N_22964);
and U29258 (N_29258,N_20631,N_21380);
and U29259 (N_29259,N_20120,N_18890);
and U29260 (N_29260,N_21341,N_21608);
nand U29261 (N_29261,N_19574,N_23683);
xnor U29262 (N_29262,N_18009,N_23629);
or U29263 (N_29263,N_18252,N_22662);
and U29264 (N_29264,N_20661,N_21811);
or U29265 (N_29265,N_19379,N_22622);
nand U29266 (N_29266,N_18220,N_20756);
xnor U29267 (N_29267,N_19137,N_23344);
and U29268 (N_29268,N_18052,N_23617);
nand U29269 (N_29269,N_18388,N_19949);
xnor U29270 (N_29270,N_21707,N_22092);
nor U29271 (N_29271,N_21285,N_20291);
and U29272 (N_29272,N_18694,N_23790);
or U29273 (N_29273,N_20921,N_22349);
nand U29274 (N_29274,N_18922,N_19780);
or U29275 (N_29275,N_22963,N_20201);
nand U29276 (N_29276,N_22436,N_19460);
xnor U29277 (N_29277,N_18125,N_21746);
or U29278 (N_29278,N_20720,N_22999);
or U29279 (N_29279,N_20168,N_19158);
nand U29280 (N_29280,N_18460,N_19205);
xnor U29281 (N_29281,N_21406,N_22869);
nand U29282 (N_29282,N_23165,N_23112);
nor U29283 (N_29283,N_21358,N_23062);
xnor U29284 (N_29284,N_21682,N_20991);
xnor U29285 (N_29285,N_19111,N_23480);
nand U29286 (N_29286,N_20937,N_20474);
nor U29287 (N_29287,N_19595,N_23731);
and U29288 (N_29288,N_21228,N_23681);
and U29289 (N_29289,N_20551,N_23618);
and U29290 (N_29290,N_20918,N_22329);
and U29291 (N_29291,N_22256,N_23991);
xor U29292 (N_29292,N_21421,N_20036);
or U29293 (N_29293,N_20885,N_23039);
and U29294 (N_29294,N_18512,N_18320);
or U29295 (N_29295,N_19170,N_23866);
xor U29296 (N_29296,N_18424,N_23688);
nand U29297 (N_29297,N_23022,N_23352);
xor U29298 (N_29298,N_20360,N_23284);
xnor U29299 (N_29299,N_18725,N_22628);
or U29300 (N_29300,N_19710,N_21920);
nor U29301 (N_29301,N_18027,N_18415);
nand U29302 (N_29302,N_19246,N_19882);
nor U29303 (N_29303,N_19611,N_18607);
or U29304 (N_29304,N_22324,N_18108);
and U29305 (N_29305,N_19755,N_20819);
xnor U29306 (N_29306,N_19451,N_19468);
and U29307 (N_29307,N_20259,N_20692);
xor U29308 (N_29308,N_18091,N_23532);
nand U29309 (N_29309,N_21301,N_19367);
xnor U29310 (N_29310,N_19272,N_22499);
xnor U29311 (N_29311,N_18499,N_22255);
nand U29312 (N_29312,N_20494,N_19864);
and U29313 (N_29313,N_22688,N_20577);
nor U29314 (N_29314,N_22344,N_23447);
and U29315 (N_29315,N_18063,N_18188);
xor U29316 (N_29316,N_21828,N_19635);
xor U29317 (N_29317,N_23611,N_22266);
xnor U29318 (N_29318,N_21237,N_23426);
and U29319 (N_29319,N_19631,N_22991);
or U29320 (N_29320,N_22662,N_20332);
or U29321 (N_29321,N_18426,N_22279);
or U29322 (N_29322,N_18380,N_19743);
nand U29323 (N_29323,N_21849,N_22265);
or U29324 (N_29324,N_23876,N_22731);
xor U29325 (N_29325,N_20129,N_21480);
and U29326 (N_29326,N_18524,N_23627);
and U29327 (N_29327,N_22352,N_19220);
or U29328 (N_29328,N_22196,N_20791);
nand U29329 (N_29329,N_18727,N_18637);
or U29330 (N_29330,N_18198,N_22185);
or U29331 (N_29331,N_20287,N_20465);
or U29332 (N_29332,N_18477,N_18465);
nand U29333 (N_29333,N_22782,N_22756);
and U29334 (N_29334,N_22628,N_23907);
nand U29335 (N_29335,N_18500,N_20551);
nand U29336 (N_29336,N_18000,N_23346);
or U29337 (N_29337,N_21709,N_18111);
nor U29338 (N_29338,N_23836,N_22993);
nor U29339 (N_29339,N_19519,N_23092);
or U29340 (N_29340,N_23913,N_18770);
or U29341 (N_29341,N_19245,N_20830);
nor U29342 (N_29342,N_22341,N_20317);
xnor U29343 (N_29343,N_21471,N_22442);
nand U29344 (N_29344,N_19874,N_19022);
xor U29345 (N_29345,N_20737,N_21039);
xnor U29346 (N_29346,N_19460,N_21045);
nor U29347 (N_29347,N_21767,N_22419);
and U29348 (N_29348,N_23809,N_19612);
and U29349 (N_29349,N_23272,N_20379);
xor U29350 (N_29350,N_23132,N_19623);
and U29351 (N_29351,N_20574,N_19681);
or U29352 (N_29352,N_21066,N_23642);
and U29353 (N_29353,N_19230,N_18775);
nor U29354 (N_29354,N_20488,N_23427);
nand U29355 (N_29355,N_23213,N_21475);
and U29356 (N_29356,N_21522,N_22902);
and U29357 (N_29357,N_23207,N_20267);
and U29358 (N_29358,N_18055,N_20499);
xor U29359 (N_29359,N_19409,N_18495);
or U29360 (N_29360,N_22606,N_20829);
nor U29361 (N_29361,N_20957,N_18647);
or U29362 (N_29362,N_21290,N_18323);
nand U29363 (N_29363,N_18259,N_18010);
nand U29364 (N_29364,N_18437,N_23257);
xnor U29365 (N_29365,N_18914,N_20723);
nand U29366 (N_29366,N_21155,N_18388);
nand U29367 (N_29367,N_23370,N_18775);
and U29368 (N_29368,N_23009,N_19005);
nand U29369 (N_29369,N_19151,N_19829);
nor U29370 (N_29370,N_21502,N_23070);
or U29371 (N_29371,N_21303,N_20801);
or U29372 (N_29372,N_21867,N_22312);
nand U29373 (N_29373,N_18561,N_22963);
nand U29374 (N_29374,N_23450,N_22862);
nand U29375 (N_29375,N_18832,N_20810);
and U29376 (N_29376,N_23837,N_22244);
nand U29377 (N_29377,N_22929,N_19272);
xnor U29378 (N_29378,N_20071,N_19546);
or U29379 (N_29379,N_18265,N_21618);
and U29380 (N_29380,N_23849,N_21466);
and U29381 (N_29381,N_23856,N_20594);
and U29382 (N_29382,N_21578,N_18003);
nand U29383 (N_29383,N_21290,N_23800);
nand U29384 (N_29384,N_19238,N_23230);
and U29385 (N_29385,N_22436,N_21254);
or U29386 (N_29386,N_22485,N_18878);
or U29387 (N_29387,N_18171,N_21412);
nor U29388 (N_29388,N_23261,N_18413);
or U29389 (N_29389,N_21489,N_18420);
xnor U29390 (N_29390,N_18147,N_19899);
and U29391 (N_29391,N_20408,N_20430);
xor U29392 (N_29392,N_21969,N_19255);
nor U29393 (N_29393,N_22826,N_22444);
or U29394 (N_29394,N_19063,N_20896);
or U29395 (N_29395,N_23924,N_18407);
xor U29396 (N_29396,N_23951,N_18751);
nor U29397 (N_29397,N_22197,N_19012);
nand U29398 (N_29398,N_21680,N_20187);
and U29399 (N_29399,N_22458,N_20564);
and U29400 (N_29400,N_19766,N_23019);
nor U29401 (N_29401,N_20139,N_23154);
nand U29402 (N_29402,N_20921,N_19036);
nand U29403 (N_29403,N_18114,N_23000);
and U29404 (N_29404,N_18769,N_19270);
nand U29405 (N_29405,N_19625,N_22024);
or U29406 (N_29406,N_20923,N_19376);
nand U29407 (N_29407,N_20105,N_23147);
nor U29408 (N_29408,N_23456,N_19047);
nor U29409 (N_29409,N_20996,N_23604);
nand U29410 (N_29410,N_23242,N_21645);
xor U29411 (N_29411,N_22387,N_19667);
and U29412 (N_29412,N_23498,N_20617);
and U29413 (N_29413,N_20411,N_21982);
xnor U29414 (N_29414,N_20517,N_23339);
or U29415 (N_29415,N_20113,N_23123);
nor U29416 (N_29416,N_21577,N_19340);
and U29417 (N_29417,N_21436,N_19524);
xnor U29418 (N_29418,N_19060,N_21450);
or U29419 (N_29419,N_19163,N_19903);
or U29420 (N_29420,N_20115,N_20770);
and U29421 (N_29421,N_21935,N_20089);
nor U29422 (N_29422,N_19882,N_22041);
nor U29423 (N_29423,N_22000,N_18430);
nand U29424 (N_29424,N_18691,N_19800);
nand U29425 (N_29425,N_22221,N_22467);
xor U29426 (N_29426,N_22334,N_22516);
xnor U29427 (N_29427,N_19861,N_19070);
nor U29428 (N_29428,N_20360,N_22571);
xor U29429 (N_29429,N_19921,N_21006);
or U29430 (N_29430,N_21577,N_22794);
or U29431 (N_29431,N_19185,N_21825);
nand U29432 (N_29432,N_19401,N_23841);
or U29433 (N_29433,N_23198,N_20084);
nor U29434 (N_29434,N_20622,N_21221);
xnor U29435 (N_29435,N_23207,N_19531);
and U29436 (N_29436,N_21459,N_20320);
xnor U29437 (N_29437,N_21524,N_21138);
nor U29438 (N_29438,N_18263,N_20442);
nand U29439 (N_29439,N_18139,N_21326);
xnor U29440 (N_29440,N_19643,N_20469);
or U29441 (N_29441,N_20151,N_19034);
nand U29442 (N_29442,N_21686,N_21990);
or U29443 (N_29443,N_23930,N_20440);
nor U29444 (N_29444,N_22609,N_19911);
nand U29445 (N_29445,N_18735,N_22916);
or U29446 (N_29446,N_22143,N_19982);
xor U29447 (N_29447,N_18335,N_18181);
and U29448 (N_29448,N_22926,N_21132);
and U29449 (N_29449,N_21827,N_22882);
and U29450 (N_29450,N_21871,N_19806);
nor U29451 (N_29451,N_23190,N_18708);
nor U29452 (N_29452,N_23672,N_23220);
xor U29453 (N_29453,N_19531,N_19047);
xor U29454 (N_29454,N_19740,N_22040);
and U29455 (N_29455,N_18217,N_18655);
nor U29456 (N_29456,N_23887,N_23190);
nand U29457 (N_29457,N_19578,N_20776);
nand U29458 (N_29458,N_21300,N_18531);
nor U29459 (N_29459,N_22768,N_23243);
or U29460 (N_29460,N_20689,N_23866);
or U29461 (N_29461,N_18803,N_18601);
and U29462 (N_29462,N_22527,N_20919);
or U29463 (N_29463,N_18475,N_23435);
and U29464 (N_29464,N_22081,N_23015);
xnor U29465 (N_29465,N_23324,N_20063);
nand U29466 (N_29466,N_19403,N_22130);
nor U29467 (N_29467,N_19514,N_23263);
or U29468 (N_29468,N_23606,N_20725);
xnor U29469 (N_29469,N_22089,N_20010);
xnor U29470 (N_29470,N_20739,N_21240);
and U29471 (N_29471,N_19728,N_20360);
and U29472 (N_29472,N_22289,N_18800);
or U29473 (N_29473,N_19156,N_22933);
or U29474 (N_29474,N_19012,N_20319);
or U29475 (N_29475,N_19389,N_21489);
and U29476 (N_29476,N_19349,N_22803);
or U29477 (N_29477,N_23006,N_22939);
and U29478 (N_29478,N_18846,N_21473);
nand U29479 (N_29479,N_20515,N_18818);
or U29480 (N_29480,N_20762,N_20989);
or U29481 (N_29481,N_19151,N_21884);
xor U29482 (N_29482,N_19643,N_21174);
or U29483 (N_29483,N_21483,N_19607);
nor U29484 (N_29484,N_19870,N_23250);
nand U29485 (N_29485,N_21038,N_20473);
and U29486 (N_29486,N_19357,N_23979);
or U29487 (N_29487,N_23128,N_20253);
and U29488 (N_29488,N_19138,N_19340);
xnor U29489 (N_29489,N_21385,N_18330);
and U29490 (N_29490,N_19144,N_19562);
nand U29491 (N_29491,N_21558,N_19638);
and U29492 (N_29492,N_22264,N_18539);
and U29493 (N_29493,N_21067,N_22370);
or U29494 (N_29494,N_23179,N_21054);
and U29495 (N_29495,N_19041,N_23404);
nand U29496 (N_29496,N_19314,N_19896);
nor U29497 (N_29497,N_20920,N_18327);
xnor U29498 (N_29498,N_18733,N_18480);
or U29499 (N_29499,N_19561,N_20119);
or U29500 (N_29500,N_23304,N_22602);
and U29501 (N_29501,N_22324,N_23259);
nand U29502 (N_29502,N_18394,N_23934);
xnor U29503 (N_29503,N_23707,N_22585);
xnor U29504 (N_29504,N_21435,N_23233);
or U29505 (N_29505,N_20117,N_23356);
xor U29506 (N_29506,N_22947,N_23642);
and U29507 (N_29507,N_23691,N_20187);
and U29508 (N_29508,N_19962,N_20583);
and U29509 (N_29509,N_22291,N_21407);
nand U29510 (N_29510,N_21392,N_20285);
or U29511 (N_29511,N_21755,N_18381);
xnor U29512 (N_29512,N_23591,N_19401);
or U29513 (N_29513,N_19862,N_20790);
nand U29514 (N_29514,N_22859,N_22349);
nand U29515 (N_29515,N_22284,N_23765);
and U29516 (N_29516,N_19743,N_19300);
xnor U29517 (N_29517,N_22881,N_23064);
and U29518 (N_29518,N_22615,N_18186);
xor U29519 (N_29519,N_23293,N_22275);
nor U29520 (N_29520,N_18047,N_18599);
nor U29521 (N_29521,N_20175,N_22501);
or U29522 (N_29522,N_19183,N_22827);
nor U29523 (N_29523,N_19098,N_18864);
and U29524 (N_29524,N_22990,N_18619);
or U29525 (N_29525,N_19035,N_20105);
nor U29526 (N_29526,N_18545,N_18638);
nand U29527 (N_29527,N_19763,N_20468);
and U29528 (N_29528,N_23017,N_20289);
and U29529 (N_29529,N_21810,N_20848);
and U29530 (N_29530,N_20972,N_23322);
nand U29531 (N_29531,N_18218,N_22663);
and U29532 (N_29532,N_19468,N_21911);
xor U29533 (N_29533,N_20356,N_20149);
or U29534 (N_29534,N_20320,N_22804);
nand U29535 (N_29535,N_23427,N_23735);
or U29536 (N_29536,N_18137,N_23285);
and U29537 (N_29537,N_22920,N_19948);
nand U29538 (N_29538,N_21970,N_18352);
xnor U29539 (N_29539,N_23192,N_23460);
or U29540 (N_29540,N_21543,N_21490);
and U29541 (N_29541,N_18190,N_23729);
or U29542 (N_29542,N_18996,N_22722);
xnor U29543 (N_29543,N_18326,N_22709);
and U29544 (N_29544,N_22061,N_18492);
nor U29545 (N_29545,N_23783,N_23496);
and U29546 (N_29546,N_20032,N_21411);
nor U29547 (N_29547,N_18409,N_23425);
nor U29548 (N_29548,N_20103,N_20763);
nor U29549 (N_29549,N_21761,N_21560);
nand U29550 (N_29550,N_19406,N_19155);
xnor U29551 (N_29551,N_23887,N_22297);
nand U29552 (N_29552,N_19099,N_20825);
nor U29553 (N_29553,N_18742,N_22854);
nor U29554 (N_29554,N_20279,N_22880);
and U29555 (N_29555,N_18232,N_19948);
or U29556 (N_29556,N_20874,N_21924);
and U29557 (N_29557,N_19295,N_20019);
nor U29558 (N_29558,N_18824,N_18161);
xnor U29559 (N_29559,N_20477,N_20577);
xnor U29560 (N_29560,N_22416,N_23684);
and U29561 (N_29561,N_18601,N_19301);
nand U29562 (N_29562,N_19233,N_22757);
nand U29563 (N_29563,N_21535,N_23767);
nand U29564 (N_29564,N_20627,N_18580);
or U29565 (N_29565,N_20417,N_18504);
nand U29566 (N_29566,N_23626,N_18242);
nor U29567 (N_29567,N_19923,N_21444);
and U29568 (N_29568,N_22539,N_21180);
and U29569 (N_29569,N_22570,N_22029);
nand U29570 (N_29570,N_20374,N_18193);
xor U29571 (N_29571,N_19057,N_19428);
nor U29572 (N_29572,N_22187,N_18173);
xor U29573 (N_29573,N_23478,N_22524);
or U29574 (N_29574,N_21777,N_19876);
nor U29575 (N_29575,N_21665,N_18352);
and U29576 (N_29576,N_20810,N_19476);
and U29577 (N_29577,N_22080,N_20857);
and U29578 (N_29578,N_21777,N_21037);
xnor U29579 (N_29579,N_18437,N_21377);
xnor U29580 (N_29580,N_18126,N_23891);
nor U29581 (N_29581,N_22287,N_23394);
and U29582 (N_29582,N_21833,N_20123);
or U29583 (N_29583,N_23444,N_19390);
or U29584 (N_29584,N_20616,N_19210);
xor U29585 (N_29585,N_22922,N_22383);
nor U29586 (N_29586,N_19183,N_22668);
or U29587 (N_29587,N_22575,N_18229);
nor U29588 (N_29588,N_23326,N_18075);
and U29589 (N_29589,N_18227,N_19159);
xor U29590 (N_29590,N_21793,N_23198);
or U29591 (N_29591,N_20143,N_18163);
and U29592 (N_29592,N_19678,N_19715);
and U29593 (N_29593,N_22207,N_18290);
and U29594 (N_29594,N_21193,N_22032);
nand U29595 (N_29595,N_20792,N_20749);
xor U29596 (N_29596,N_19591,N_22950);
nor U29597 (N_29597,N_20916,N_21409);
or U29598 (N_29598,N_18861,N_23603);
nand U29599 (N_29599,N_18000,N_22380);
and U29600 (N_29600,N_19642,N_22498);
xor U29601 (N_29601,N_22962,N_23911);
nor U29602 (N_29602,N_19662,N_21625);
or U29603 (N_29603,N_18654,N_23188);
nor U29604 (N_29604,N_20660,N_23326);
xnor U29605 (N_29605,N_18700,N_22288);
nand U29606 (N_29606,N_22631,N_23353);
and U29607 (N_29607,N_18773,N_22874);
nor U29608 (N_29608,N_23776,N_19783);
nand U29609 (N_29609,N_23193,N_22590);
or U29610 (N_29610,N_23112,N_18670);
or U29611 (N_29611,N_19710,N_19824);
or U29612 (N_29612,N_18138,N_23999);
or U29613 (N_29613,N_20079,N_23715);
and U29614 (N_29614,N_23463,N_22067);
xor U29615 (N_29615,N_21884,N_23397);
and U29616 (N_29616,N_18655,N_21582);
nor U29617 (N_29617,N_19176,N_20870);
xnor U29618 (N_29618,N_23208,N_23950);
or U29619 (N_29619,N_20576,N_18219);
and U29620 (N_29620,N_20992,N_23358);
or U29621 (N_29621,N_21592,N_18200);
xnor U29622 (N_29622,N_19067,N_23915);
or U29623 (N_29623,N_21817,N_21535);
nor U29624 (N_29624,N_18362,N_23313);
xor U29625 (N_29625,N_21186,N_21113);
xor U29626 (N_29626,N_23807,N_21469);
nand U29627 (N_29627,N_21741,N_23677);
xor U29628 (N_29628,N_19314,N_21128);
or U29629 (N_29629,N_18266,N_23433);
and U29630 (N_29630,N_18992,N_23663);
xor U29631 (N_29631,N_22526,N_18436);
and U29632 (N_29632,N_19955,N_21730);
nor U29633 (N_29633,N_20109,N_20234);
nand U29634 (N_29634,N_19453,N_18257);
or U29635 (N_29635,N_19780,N_23318);
and U29636 (N_29636,N_18118,N_20269);
nand U29637 (N_29637,N_22576,N_22564);
nor U29638 (N_29638,N_20045,N_18801);
nand U29639 (N_29639,N_22312,N_21397);
nor U29640 (N_29640,N_20011,N_19218);
nor U29641 (N_29641,N_20193,N_23458);
and U29642 (N_29642,N_23218,N_23353);
nand U29643 (N_29643,N_21555,N_19333);
xnor U29644 (N_29644,N_20488,N_18613);
and U29645 (N_29645,N_20514,N_19947);
xor U29646 (N_29646,N_21552,N_23141);
nand U29647 (N_29647,N_20901,N_18104);
and U29648 (N_29648,N_23063,N_19168);
xor U29649 (N_29649,N_18293,N_22456);
nand U29650 (N_29650,N_19463,N_22725);
or U29651 (N_29651,N_21297,N_19346);
or U29652 (N_29652,N_21021,N_22233);
and U29653 (N_29653,N_19958,N_23938);
nand U29654 (N_29654,N_20589,N_18362);
nor U29655 (N_29655,N_21115,N_18017);
or U29656 (N_29656,N_21899,N_20557);
xnor U29657 (N_29657,N_22268,N_20997);
or U29658 (N_29658,N_22922,N_21486);
nor U29659 (N_29659,N_23219,N_22367);
nor U29660 (N_29660,N_21078,N_23684);
nand U29661 (N_29661,N_22881,N_19751);
nor U29662 (N_29662,N_22777,N_23141);
or U29663 (N_29663,N_23784,N_22410);
or U29664 (N_29664,N_20725,N_22636);
nor U29665 (N_29665,N_21823,N_23736);
nand U29666 (N_29666,N_19013,N_21885);
and U29667 (N_29667,N_20716,N_23775);
nor U29668 (N_29668,N_20082,N_23910);
nand U29669 (N_29669,N_18284,N_20771);
and U29670 (N_29670,N_19474,N_18679);
xnor U29671 (N_29671,N_21670,N_23545);
and U29672 (N_29672,N_23921,N_22247);
nor U29673 (N_29673,N_18545,N_22578);
or U29674 (N_29674,N_21396,N_22093);
xnor U29675 (N_29675,N_22954,N_19809);
nand U29676 (N_29676,N_23819,N_21440);
xnor U29677 (N_29677,N_22591,N_19078);
or U29678 (N_29678,N_22552,N_19479);
xnor U29679 (N_29679,N_18358,N_18002);
or U29680 (N_29680,N_23401,N_22242);
nor U29681 (N_29681,N_21883,N_20727);
or U29682 (N_29682,N_19819,N_19490);
or U29683 (N_29683,N_20024,N_18191);
xnor U29684 (N_29684,N_20999,N_19434);
or U29685 (N_29685,N_21091,N_22829);
xor U29686 (N_29686,N_20763,N_19425);
or U29687 (N_29687,N_18656,N_21212);
nor U29688 (N_29688,N_20287,N_19492);
or U29689 (N_29689,N_23268,N_22509);
xor U29690 (N_29690,N_20334,N_18841);
xor U29691 (N_29691,N_23292,N_18963);
xnor U29692 (N_29692,N_18361,N_19309);
or U29693 (N_29693,N_19576,N_23167);
or U29694 (N_29694,N_19484,N_20885);
xor U29695 (N_29695,N_20985,N_21387);
nand U29696 (N_29696,N_20216,N_20393);
and U29697 (N_29697,N_18303,N_18256);
and U29698 (N_29698,N_23619,N_22809);
nor U29699 (N_29699,N_19113,N_23661);
nand U29700 (N_29700,N_21019,N_19253);
or U29701 (N_29701,N_21637,N_20220);
nand U29702 (N_29702,N_18515,N_20009);
xnor U29703 (N_29703,N_19627,N_23731);
nand U29704 (N_29704,N_22803,N_22871);
nor U29705 (N_29705,N_21041,N_22433);
xnor U29706 (N_29706,N_18162,N_18284);
xnor U29707 (N_29707,N_19333,N_22032);
and U29708 (N_29708,N_20534,N_21766);
nor U29709 (N_29709,N_20393,N_19957);
and U29710 (N_29710,N_21479,N_22943);
xnor U29711 (N_29711,N_21379,N_21704);
nor U29712 (N_29712,N_21749,N_19924);
or U29713 (N_29713,N_23963,N_21366);
and U29714 (N_29714,N_18946,N_20165);
and U29715 (N_29715,N_22635,N_21127);
nand U29716 (N_29716,N_21157,N_18958);
and U29717 (N_29717,N_18263,N_22084);
nor U29718 (N_29718,N_21999,N_19821);
nor U29719 (N_29719,N_23706,N_22590);
or U29720 (N_29720,N_18111,N_22951);
and U29721 (N_29721,N_21987,N_19680);
nor U29722 (N_29722,N_19689,N_22019);
nand U29723 (N_29723,N_22782,N_21722);
or U29724 (N_29724,N_22652,N_23549);
nor U29725 (N_29725,N_21008,N_20558);
nand U29726 (N_29726,N_21078,N_20242);
nand U29727 (N_29727,N_23901,N_23663);
and U29728 (N_29728,N_19334,N_23025);
nand U29729 (N_29729,N_22095,N_20290);
nor U29730 (N_29730,N_23054,N_22939);
or U29731 (N_29731,N_23799,N_23158);
nand U29732 (N_29732,N_20659,N_20469);
or U29733 (N_29733,N_23134,N_21212);
xnor U29734 (N_29734,N_20276,N_18322);
or U29735 (N_29735,N_19769,N_20247);
nand U29736 (N_29736,N_19499,N_19654);
nor U29737 (N_29737,N_18613,N_20762);
nor U29738 (N_29738,N_21989,N_22691);
or U29739 (N_29739,N_23562,N_20372);
or U29740 (N_29740,N_18540,N_18542);
nand U29741 (N_29741,N_19271,N_22737);
nand U29742 (N_29742,N_23742,N_23685);
and U29743 (N_29743,N_18772,N_18945);
nor U29744 (N_29744,N_22494,N_19897);
and U29745 (N_29745,N_23345,N_22081);
or U29746 (N_29746,N_21365,N_22912);
xnor U29747 (N_29747,N_22174,N_20149);
or U29748 (N_29748,N_19298,N_20595);
nand U29749 (N_29749,N_19586,N_20622);
and U29750 (N_29750,N_23886,N_20483);
and U29751 (N_29751,N_18727,N_21981);
and U29752 (N_29752,N_23946,N_23241);
nor U29753 (N_29753,N_18105,N_21969);
nor U29754 (N_29754,N_20864,N_21424);
or U29755 (N_29755,N_23806,N_19727);
nor U29756 (N_29756,N_22306,N_18399);
or U29757 (N_29757,N_23860,N_21595);
or U29758 (N_29758,N_20049,N_18964);
xnor U29759 (N_29759,N_18325,N_20649);
and U29760 (N_29760,N_22099,N_22420);
or U29761 (N_29761,N_18424,N_18221);
and U29762 (N_29762,N_20136,N_19107);
and U29763 (N_29763,N_23529,N_19550);
or U29764 (N_29764,N_23749,N_23106);
nand U29765 (N_29765,N_18068,N_23212);
nand U29766 (N_29766,N_18052,N_21316);
nand U29767 (N_29767,N_20937,N_22080);
nand U29768 (N_29768,N_23847,N_22225);
nor U29769 (N_29769,N_18998,N_21701);
or U29770 (N_29770,N_23197,N_19802);
xnor U29771 (N_29771,N_19943,N_18985);
nor U29772 (N_29772,N_23620,N_19805);
or U29773 (N_29773,N_23308,N_19835);
nand U29774 (N_29774,N_23201,N_20100);
and U29775 (N_29775,N_22599,N_18352);
xnor U29776 (N_29776,N_21794,N_20635);
nor U29777 (N_29777,N_22006,N_20527);
nand U29778 (N_29778,N_22285,N_19672);
and U29779 (N_29779,N_23319,N_21492);
nor U29780 (N_29780,N_22103,N_21562);
and U29781 (N_29781,N_19617,N_19720);
or U29782 (N_29782,N_23454,N_21292);
and U29783 (N_29783,N_20595,N_19046);
or U29784 (N_29784,N_23621,N_18455);
xor U29785 (N_29785,N_20689,N_21412);
nand U29786 (N_29786,N_20141,N_22154);
xnor U29787 (N_29787,N_19255,N_23016);
xor U29788 (N_29788,N_21024,N_18422);
or U29789 (N_29789,N_20535,N_19578);
or U29790 (N_29790,N_18667,N_21726);
or U29791 (N_29791,N_19923,N_21455);
nor U29792 (N_29792,N_19503,N_18098);
xor U29793 (N_29793,N_22551,N_18535);
nor U29794 (N_29794,N_22141,N_22258);
nand U29795 (N_29795,N_20106,N_21245);
xnor U29796 (N_29796,N_23766,N_23232);
xnor U29797 (N_29797,N_22412,N_21596);
nand U29798 (N_29798,N_18475,N_23478);
xnor U29799 (N_29799,N_22311,N_20830);
nand U29800 (N_29800,N_22075,N_22954);
nand U29801 (N_29801,N_18290,N_23568);
xnor U29802 (N_29802,N_19963,N_23771);
xor U29803 (N_29803,N_23120,N_21255);
or U29804 (N_29804,N_20615,N_19053);
or U29805 (N_29805,N_23337,N_21060);
nor U29806 (N_29806,N_21052,N_18394);
xnor U29807 (N_29807,N_20378,N_23577);
xor U29808 (N_29808,N_18903,N_18404);
nand U29809 (N_29809,N_22614,N_20170);
nor U29810 (N_29810,N_22130,N_23984);
nand U29811 (N_29811,N_20675,N_20391);
nor U29812 (N_29812,N_20079,N_20194);
nor U29813 (N_29813,N_23527,N_18850);
nor U29814 (N_29814,N_23551,N_18104);
nor U29815 (N_29815,N_22912,N_19406);
or U29816 (N_29816,N_20816,N_20114);
nor U29817 (N_29817,N_22156,N_23069);
and U29818 (N_29818,N_23930,N_22401);
nor U29819 (N_29819,N_22865,N_20503);
xnor U29820 (N_29820,N_21745,N_18721);
and U29821 (N_29821,N_19777,N_20492);
and U29822 (N_29822,N_21336,N_22713);
and U29823 (N_29823,N_21000,N_18528);
and U29824 (N_29824,N_23226,N_20634);
xor U29825 (N_29825,N_21149,N_18158);
and U29826 (N_29826,N_22147,N_18139);
or U29827 (N_29827,N_20435,N_22473);
nand U29828 (N_29828,N_18901,N_23311);
and U29829 (N_29829,N_21521,N_21523);
nand U29830 (N_29830,N_21039,N_20938);
nor U29831 (N_29831,N_19331,N_22093);
nand U29832 (N_29832,N_20251,N_21572);
or U29833 (N_29833,N_23326,N_19016);
xor U29834 (N_29834,N_22842,N_19484);
or U29835 (N_29835,N_19778,N_23388);
xnor U29836 (N_29836,N_19073,N_23326);
nand U29837 (N_29837,N_18081,N_20785);
or U29838 (N_29838,N_22884,N_18369);
or U29839 (N_29839,N_19347,N_18830);
nand U29840 (N_29840,N_21624,N_23841);
nor U29841 (N_29841,N_18181,N_19118);
and U29842 (N_29842,N_21887,N_20566);
nor U29843 (N_29843,N_18518,N_21919);
xnor U29844 (N_29844,N_23075,N_23602);
nor U29845 (N_29845,N_22754,N_23530);
xnor U29846 (N_29846,N_18184,N_20693);
or U29847 (N_29847,N_20697,N_18380);
xnor U29848 (N_29848,N_22240,N_20597);
nor U29849 (N_29849,N_23939,N_18286);
nor U29850 (N_29850,N_22207,N_21275);
nor U29851 (N_29851,N_21958,N_19180);
nand U29852 (N_29852,N_20022,N_23638);
and U29853 (N_29853,N_23630,N_20038);
and U29854 (N_29854,N_23890,N_23120);
and U29855 (N_29855,N_18420,N_23599);
nor U29856 (N_29856,N_23986,N_20043);
nor U29857 (N_29857,N_21315,N_23765);
xnor U29858 (N_29858,N_18457,N_21331);
nand U29859 (N_29859,N_23817,N_21700);
nor U29860 (N_29860,N_20455,N_23194);
xor U29861 (N_29861,N_23730,N_18842);
xnor U29862 (N_29862,N_21767,N_19513);
nor U29863 (N_29863,N_19017,N_18709);
xor U29864 (N_29864,N_20042,N_23574);
nand U29865 (N_29865,N_21529,N_23201);
and U29866 (N_29866,N_23267,N_23006);
and U29867 (N_29867,N_20926,N_22052);
or U29868 (N_29868,N_21674,N_22936);
nor U29869 (N_29869,N_19228,N_19274);
or U29870 (N_29870,N_18234,N_21434);
or U29871 (N_29871,N_22190,N_21679);
or U29872 (N_29872,N_20208,N_18729);
nand U29873 (N_29873,N_20138,N_18565);
nand U29874 (N_29874,N_23078,N_22777);
and U29875 (N_29875,N_23799,N_23751);
and U29876 (N_29876,N_22483,N_20669);
xnor U29877 (N_29877,N_19783,N_19699);
nor U29878 (N_29878,N_23676,N_23327);
nor U29879 (N_29879,N_22869,N_23230);
or U29880 (N_29880,N_19838,N_19580);
nor U29881 (N_29881,N_19871,N_20176);
and U29882 (N_29882,N_21872,N_18581);
and U29883 (N_29883,N_21503,N_19389);
xor U29884 (N_29884,N_19976,N_20960);
or U29885 (N_29885,N_22389,N_20911);
and U29886 (N_29886,N_22009,N_20589);
nand U29887 (N_29887,N_20352,N_20984);
nand U29888 (N_29888,N_22263,N_19504);
xor U29889 (N_29889,N_23101,N_23807);
xor U29890 (N_29890,N_22421,N_18815);
xnor U29891 (N_29891,N_22832,N_22145);
nand U29892 (N_29892,N_22753,N_22100);
and U29893 (N_29893,N_23706,N_18819);
xor U29894 (N_29894,N_21723,N_20013);
nand U29895 (N_29895,N_18611,N_22928);
xor U29896 (N_29896,N_23209,N_20405);
xnor U29897 (N_29897,N_20083,N_21809);
nand U29898 (N_29898,N_18303,N_20502);
nor U29899 (N_29899,N_22344,N_22333);
nand U29900 (N_29900,N_19791,N_20504);
or U29901 (N_29901,N_18548,N_22487);
nand U29902 (N_29902,N_20320,N_22813);
nor U29903 (N_29903,N_18927,N_18857);
nor U29904 (N_29904,N_19079,N_22597);
nand U29905 (N_29905,N_19433,N_18108);
or U29906 (N_29906,N_19420,N_22809);
nand U29907 (N_29907,N_21604,N_19533);
nor U29908 (N_29908,N_19903,N_19702);
nand U29909 (N_29909,N_20930,N_23545);
or U29910 (N_29910,N_22535,N_18839);
or U29911 (N_29911,N_19223,N_20637);
or U29912 (N_29912,N_18815,N_19247);
and U29913 (N_29913,N_20156,N_19894);
nor U29914 (N_29914,N_21461,N_19635);
or U29915 (N_29915,N_21689,N_21359);
xnor U29916 (N_29916,N_19359,N_19710);
or U29917 (N_29917,N_20417,N_22564);
xor U29918 (N_29918,N_19855,N_20382);
nand U29919 (N_29919,N_23139,N_20541);
nor U29920 (N_29920,N_21338,N_20316);
and U29921 (N_29921,N_18039,N_19658);
or U29922 (N_29922,N_18000,N_18571);
or U29923 (N_29923,N_23812,N_22490);
nor U29924 (N_29924,N_23272,N_19291);
xnor U29925 (N_29925,N_18900,N_21235);
and U29926 (N_29926,N_23881,N_21658);
or U29927 (N_29927,N_23675,N_21724);
or U29928 (N_29928,N_22916,N_19116);
xor U29929 (N_29929,N_18814,N_18809);
xor U29930 (N_29930,N_19591,N_22297);
and U29931 (N_29931,N_20380,N_20709);
or U29932 (N_29932,N_19514,N_18787);
xnor U29933 (N_29933,N_21394,N_22037);
and U29934 (N_29934,N_22932,N_18925);
nand U29935 (N_29935,N_18497,N_21035);
and U29936 (N_29936,N_21811,N_19877);
nand U29937 (N_29937,N_20900,N_23358);
xor U29938 (N_29938,N_18122,N_21162);
and U29939 (N_29939,N_21850,N_21598);
xnor U29940 (N_29940,N_20907,N_20540);
and U29941 (N_29941,N_21795,N_23074);
nand U29942 (N_29942,N_20502,N_18406);
or U29943 (N_29943,N_19116,N_20282);
and U29944 (N_29944,N_19900,N_20144);
xnor U29945 (N_29945,N_18973,N_20980);
nand U29946 (N_29946,N_21744,N_19237);
nor U29947 (N_29947,N_18584,N_21708);
or U29948 (N_29948,N_20492,N_22311);
nand U29949 (N_29949,N_18111,N_20083);
xor U29950 (N_29950,N_22070,N_19159);
and U29951 (N_29951,N_21216,N_18000);
and U29952 (N_29952,N_20778,N_20793);
nor U29953 (N_29953,N_21230,N_18052);
or U29954 (N_29954,N_21384,N_20923);
or U29955 (N_29955,N_20899,N_22501);
or U29956 (N_29956,N_23322,N_21080);
nor U29957 (N_29957,N_21142,N_20021);
or U29958 (N_29958,N_21898,N_20288);
xor U29959 (N_29959,N_18784,N_22654);
or U29960 (N_29960,N_22031,N_22762);
nor U29961 (N_29961,N_20406,N_22953);
nor U29962 (N_29962,N_22711,N_18940);
nand U29963 (N_29963,N_21105,N_20566);
nand U29964 (N_29964,N_23926,N_19774);
and U29965 (N_29965,N_22865,N_23249);
xor U29966 (N_29966,N_23929,N_18957);
xnor U29967 (N_29967,N_22768,N_23392);
nor U29968 (N_29968,N_18417,N_18657);
or U29969 (N_29969,N_18406,N_21434);
nor U29970 (N_29970,N_23894,N_23568);
xnor U29971 (N_29971,N_19923,N_20838);
xnor U29972 (N_29972,N_22141,N_22742);
nand U29973 (N_29973,N_18421,N_18731);
or U29974 (N_29974,N_23062,N_21879);
xnor U29975 (N_29975,N_18128,N_20565);
xnor U29976 (N_29976,N_23370,N_22126);
nor U29977 (N_29977,N_19204,N_22253);
nor U29978 (N_29978,N_22084,N_23416);
nand U29979 (N_29979,N_22045,N_22772);
nand U29980 (N_29980,N_18286,N_23077);
nand U29981 (N_29981,N_18011,N_19427);
xor U29982 (N_29982,N_23094,N_18421);
or U29983 (N_29983,N_20212,N_19465);
and U29984 (N_29984,N_21986,N_21353);
nor U29985 (N_29985,N_23882,N_20917);
nor U29986 (N_29986,N_19891,N_23604);
nor U29987 (N_29987,N_20337,N_21376);
xor U29988 (N_29988,N_18904,N_20369);
xnor U29989 (N_29989,N_18346,N_18037);
and U29990 (N_29990,N_22281,N_22619);
xor U29991 (N_29991,N_20318,N_23226);
and U29992 (N_29992,N_21740,N_18319);
or U29993 (N_29993,N_19629,N_20817);
and U29994 (N_29994,N_20735,N_22026);
and U29995 (N_29995,N_19414,N_23296);
xnor U29996 (N_29996,N_19513,N_23955);
nand U29997 (N_29997,N_21672,N_23827);
nand U29998 (N_29998,N_18663,N_22595);
and U29999 (N_29999,N_21964,N_18410);
nor UO_0 (O_0,N_27962,N_29839);
xor UO_1 (O_1,N_24711,N_28842);
or UO_2 (O_2,N_27083,N_24193);
and UO_3 (O_3,N_27475,N_29284);
and UO_4 (O_4,N_24550,N_29663);
nor UO_5 (O_5,N_27608,N_27281);
and UO_6 (O_6,N_29218,N_27894);
or UO_7 (O_7,N_25552,N_27166);
nand UO_8 (O_8,N_29921,N_26640);
and UO_9 (O_9,N_24738,N_27792);
or UO_10 (O_10,N_28114,N_26394);
nor UO_11 (O_11,N_26905,N_24703);
nand UO_12 (O_12,N_29703,N_28780);
and UO_13 (O_13,N_27648,N_26512);
nor UO_14 (O_14,N_24413,N_26396);
nor UO_15 (O_15,N_27832,N_29176);
nor UO_16 (O_16,N_28257,N_29886);
nor UO_17 (O_17,N_25288,N_25785);
xnor UO_18 (O_18,N_26095,N_27933);
nand UO_19 (O_19,N_27161,N_24389);
xor UO_20 (O_20,N_26572,N_28392);
xnor UO_21 (O_21,N_28922,N_27163);
xnor UO_22 (O_22,N_24598,N_24937);
or UO_23 (O_23,N_28136,N_24453);
and UO_24 (O_24,N_29067,N_28358);
or UO_25 (O_25,N_25858,N_25137);
nor UO_26 (O_26,N_27004,N_26945);
and UO_27 (O_27,N_24203,N_28773);
and UO_28 (O_28,N_24974,N_25204);
nand UO_29 (O_29,N_26787,N_28928);
nor UO_30 (O_30,N_28754,N_28140);
and UO_31 (O_31,N_25131,N_24356);
nor UO_32 (O_32,N_25320,N_29336);
nor UO_33 (O_33,N_24656,N_24150);
nor UO_34 (O_34,N_25100,N_26962);
xnor UO_35 (O_35,N_24385,N_26002);
xor UO_36 (O_36,N_26858,N_25806);
and UO_37 (O_37,N_25626,N_29406);
nor UO_38 (O_38,N_24571,N_24552);
and UO_39 (O_39,N_29498,N_24543);
nand UO_40 (O_40,N_27113,N_24194);
xnor UO_41 (O_41,N_27386,N_28656);
nor UO_42 (O_42,N_26177,N_27826);
nand UO_43 (O_43,N_27794,N_25326);
xor UO_44 (O_44,N_28985,N_26405);
and UO_45 (O_45,N_28573,N_25134);
nor UO_46 (O_46,N_25817,N_27585);
or UO_47 (O_47,N_24753,N_27292);
nor UO_48 (O_48,N_24785,N_24648);
xnor UO_49 (O_49,N_27171,N_24304);
nor UO_50 (O_50,N_26598,N_24911);
nand UO_51 (O_51,N_27329,N_28121);
and UO_52 (O_52,N_25191,N_26094);
or UO_53 (O_53,N_28681,N_29053);
and UO_54 (O_54,N_26496,N_24249);
xor UO_55 (O_55,N_28889,N_29774);
xor UO_56 (O_56,N_27588,N_24374);
xnor UO_57 (O_57,N_28072,N_26412);
nand UO_58 (O_58,N_28579,N_29039);
nand UO_59 (O_59,N_25089,N_26878);
xor UO_60 (O_60,N_29057,N_25022);
and UO_61 (O_61,N_25480,N_24211);
nor UO_62 (O_62,N_27492,N_29717);
nor UO_63 (O_63,N_26350,N_24667);
nand UO_64 (O_64,N_28008,N_25487);
nand UO_65 (O_65,N_27101,N_29418);
or UO_66 (O_66,N_28520,N_27079);
xor UO_67 (O_67,N_27066,N_26319);
xnor UO_68 (O_68,N_28941,N_26497);
and UO_69 (O_69,N_24679,N_26137);
and UO_70 (O_70,N_25575,N_25498);
nand UO_71 (O_71,N_26129,N_28147);
nand UO_72 (O_72,N_29389,N_25745);
nand UO_73 (O_73,N_24814,N_29248);
nand UO_74 (O_74,N_25442,N_29182);
nand UO_75 (O_75,N_25365,N_24151);
nor UO_76 (O_76,N_27998,N_27474);
nor UO_77 (O_77,N_28923,N_25472);
nand UO_78 (O_78,N_28921,N_28296);
nand UO_79 (O_79,N_26491,N_26501);
nor UO_80 (O_80,N_25112,N_28668);
xor UO_81 (O_81,N_29226,N_25143);
or UO_82 (O_82,N_28319,N_24567);
nand UO_83 (O_83,N_29402,N_28696);
nand UO_84 (O_84,N_25666,N_24159);
or UO_85 (O_85,N_28198,N_24106);
nor UO_86 (O_86,N_24419,N_25652);
or UO_87 (O_87,N_27866,N_29925);
or UO_88 (O_88,N_28424,N_28102);
xnor UO_89 (O_89,N_25185,N_29142);
xor UO_90 (O_90,N_27736,N_29795);
xnor UO_91 (O_91,N_24474,N_24288);
nand UO_92 (O_92,N_25184,N_28789);
xnor UO_93 (O_93,N_29748,N_28628);
and UO_94 (O_94,N_25001,N_26393);
and UO_95 (O_95,N_27592,N_27486);
nor UO_96 (O_96,N_28654,N_26605);
nor UO_97 (O_97,N_26233,N_29290);
or UO_98 (O_98,N_27927,N_29278);
xor UO_99 (O_99,N_29741,N_27176);
nand UO_100 (O_100,N_25933,N_28788);
or UO_101 (O_101,N_25226,N_29954);
or UO_102 (O_102,N_27768,N_29169);
nand UO_103 (O_103,N_28717,N_27304);
xnor UO_104 (O_104,N_29983,N_27147);
nor UO_105 (O_105,N_26833,N_29249);
xor UO_106 (O_106,N_27297,N_27958);
and UO_107 (O_107,N_27373,N_24811);
or UO_108 (O_108,N_29327,N_29549);
or UO_109 (O_109,N_28253,N_28252);
nand UO_110 (O_110,N_24450,N_29118);
nand UO_111 (O_111,N_27034,N_27779);
or UO_112 (O_112,N_26173,N_25646);
and UO_113 (O_113,N_25960,N_29937);
xnor UO_114 (O_114,N_24661,N_25572);
and UO_115 (O_115,N_26447,N_25726);
nor UO_116 (O_116,N_27035,N_28208);
and UO_117 (O_117,N_28359,N_26340);
or UO_118 (O_118,N_28461,N_27765);
and UO_119 (O_119,N_24588,N_26556);
xnor UO_120 (O_120,N_24366,N_24109);
or UO_121 (O_121,N_25183,N_27547);
and UO_122 (O_122,N_25988,N_24923);
or UO_123 (O_123,N_24977,N_29240);
xnor UO_124 (O_124,N_27072,N_27482);
xnor UO_125 (O_125,N_29531,N_29130);
or UO_126 (O_126,N_26639,N_27076);
nor UO_127 (O_127,N_24171,N_28015);
xnor UO_128 (O_128,N_26433,N_26202);
nand UO_129 (O_129,N_29298,N_25418);
xnor UO_130 (O_130,N_26961,N_26462);
and UO_131 (O_131,N_25382,N_29437);
xnor UO_132 (O_132,N_29584,N_29805);
xor UO_133 (O_133,N_27200,N_29380);
nand UO_134 (O_134,N_27013,N_29850);
nand UO_135 (O_135,N_26113,N_29054);
nor UO_136 (O_136,N_24298,N_29210);
or UO_137 (O_137,N_25376,N_25065);
or UO_138 (O_138,N_27940,N_29729);
nand UO_139 (O_139,N_26187,N_29005);
nand UO_140 (O_140,N_25884,N_28423);
nor UO_141 (O_141,N_28731,N_26381);
and UO_142 (O_142,N_29334,N_28859);
nand UO_143 (O_143,N_26475,N_24485);
nand UO_144 (O_144,N_27627,N_29344);
nor UO_145 (O_145,N_28575,N_28294);
and UO_146 (O_146,N_29496,N_25297);
nand UO_147 (O_147,N_24927,N_28959);
nor UO_148 (O_148,N_27662,N_26716);
or UO_149 (O_149,N_25427,N_27495);
xor UO_150 (O_150,N_28478,N_27276);
and UO_151 (O_151,N_25470,N_25019);
xor UO_152 (O_152,N_25668,N_28713);
and UO_153 (O_153,N_26717,N_25986);
xor UO_154 (O_154,N_24457,N_26130);
nand UO_155 (O_155,N_29945,N_24227);
nor UO_156 (O_156,N_29694,N_28270);
or UO_157 (O_157,N_26244,N_27092);
nor UO_158 (O_158,N_26638,N_25166);
or UO_159 (O_159,N_26321,N_28705);
xnor UO_160 (O_160,N_27516,N_26266);
and UO_161 (O_161,N_29618,N_27974);
and UO_162 (O_162,N_26855,N_26887);
or UO_163 (O_163,N_27154,N_25816);
xor UO_164 (O_164,N_28802,N_29066);
nand UO_165 (O_165,N_29812,N_24496);
or UO_166 (O_166,N_25928,N_24783);
nand UO_167 (O_167,N_26423,N_26934);
xnor UO_168 (O_168,N_28088,N_28973);
or UO_169 (O_169,N_26697,N_28206);
nand UO_170 (O_170,N_24274,N_27942);
or UO_171 (O_171,N_27561,N_26649);
xnor UO_172 (O_172,N_28622,N_24086);
nor UO_173 (O_173,N_24842,N_24975);
or UO_174 (O_174,N_29259,N_24772);
nor UO_175 (O_175,N_26384,N_25469);
nor UO_176 (O_176,N_26546,N_29132);
nor UO_177 (O_177,N_27414,N_25605);
or UO_178 (O_178,N_26884,N_29236);
or UO_179 (O_179,N_25518,N_26227);
xnor UO_180 (O_180,N_24087,N_28778);
or UO_181 (O_181,N_27604,N_26196);
xor UO_182 (O_182,N_29956,N_26989);
xnor UO_183 (O_183,N_25386,N_29629);
and UO_184 (O_184,N_28619,N_26048);
nor UO_185 (O_185,N_25432,N_25856);
and UO_186 (O_186,N_26499,N_27714);
xnor UO_187 (O_187,N_26353,N_28398);
and UO_188 (O_188,N_27351,N_29676);
xor UO_189 (O_189,N_25950,N_26943);
or UO_190 (O_190,N_27621,N_28223);
nor UO_191 (O_191,N_29858,N_24311);
nor UO_192 (O_192,N_25701,N_24275);
or UO_193 (O_193,N_25609,N_24530);
nand UO_194 (O_194,N_28176,N_29143);
nor UO_195 (O_195,N_26775,N_29079);
nor UO_196 (O_196,N_29239,N_29711);
xnor UO_197 (O_197,N_24885,N_25830);
and UO_198 (O_198,N_25046,N_24220);
and UO_199 (O_199,N_24912,N_28758);
and UO_200 (O_200,N_25512,N_25748);
and UO_201 (O_201,N_29837,N_27746);
xor UO_202 (O_202,N_26477,N_26927);
xor UO_203 (O_203,N_24253,N_24578);
nor UO_204 (O_204,N_25892,N_25885);
and UO_205 (O_205,N_29785,N_28699);
or UO_206 (O_206,N_29173,N_29371);
nor UO_207 (O_207,N_28884,N_25828);
xnor UO_208 (O_208,N_24263,N_25583);
nand UO_209 (O_209,N_25047,N_27575);
or UO_210 (O_210,N_26300,N_25760);
and UO_211 (O_211,N_28823,N_24765);
and UO_212 (O_212,N_24320,N_26681);
xor UO_213 (O_213,N_24382,N_27945);
xnor UO_214 (O_214,N_29623,N_28847);
nand UO_215 (O_215,N_28538,N_28230);
and UO_216 (O_216,N_28032,N_27433);
nand UO_217 (O_217,N_26397,N_24947);
nor UO_218 (O_218,N_27848,N_25632);
nor UO_219 (O_219,N_27531,N_28427);
and UO_220 (O_220,N_24510,N_28352);
xor UO_221 (O_221,N_26387,N_24644);
or UO_222 (O_222,N_26761,N_24671);
nand UO_223 (O_223,N_25690,N_28625);
and UO_224 (O_224,N_26985,N_26751);
and UO_225 (O_225,N_27730,N_25150);
xnor UO_226 (O_226,N_24396,N_29340);
or UO_227 (O_227,N_27844,N_26245);
nand UO_228 (O_228,N_28969,N_29238);
or UO_229 (O_229,N_26795,N_28262);
or UO_230 (O_230,N_26867,N_28432);
nor UO_231 (O_231,N_29543,N_28081);
nand UO_232 (O_232,N_27535,N_25050);
nand UO_233 (O_233,N_29902,N_26937);
xor UO_234 (O_234,N_27272,N_25409);
nor UO_235 (O_235,N_26438,N_29510);
or UO_236 (O_236,N_26599,N_26912);
or UO_237 (O_237,N_28554,N_28500);
nor UO_238 (O_238,N_28944,N_26118);
xnor UO_239 (O_239,N_26526,N_28016);
nor UO_240 (O_240,N_26591,N_28597);
nand UO_241 (O_241,N_24969,N_24279);
and UO_242 (O_242,N_27217,N_25265);
or UO_243 (O_243,N_29760,N_24339);
or UO_244 (O_244,N_25795,N_28063);
or UO_245 (O_245,N_26217,N_26733);
nand UO_246 (O_246,N_24354,N_28836);
nand UO_247 (O_247,N_24820,N_25390);
or UO_248 (O_248,N_25940,N_27514);
xor UO_249 (O_249,N_26328,N_26410);
xnor UO_250 (O_250,N_29713,N_27082);
xor UO_251 (O_251,N_28852,N_27522);
and UO_252 (O_252,N_24500,N_27128);
or UO_253 (O_253,N_27574,N_25061);
nand UO_254 (O_254,N_25896,N_26379);
and UO_255 (O_255,N_26105,N_24930);
or UO_256 (O_256,N_25704,N_27829);
nand UO_257 (O_257,N_28553,N_26659);
xor UO_258 (O_258,N_29879,N_24407);
nand UO_259 (O_259,N_27569,N_27607);
and UO_260 (O_260,N_26239,N_28443);
and UO_261 (O_261,N_24777,N_24551);
and UO_262 (O_262,N_28824,N_24537);
nor UO_263 (O_263,N_28112,N_29749);
nor UO_264 (O_264,N_25257,N_28490);
nand UO_265 (O_265,N_28957,N_25732);
nor UO_266 (O_266,N_28099,N_29472);
xor UO_267 (O_267,N_26758,N_27371);
xor UO_268 (O_268,N_29267,N_25360);
nor UO_269 (O_269,N_28698,N_26283);
xnor UO_270 (O_270,N_29939,N_27700);
or UO_271 (O_271,N_25459,N_28195);
or UO_272 (O_272,N_26749,N_24364);
xor UO_273 (O_273,N_24846,N_27837);
nand UO_274 (O_274,N_28709,N_25304);
or UO_275 (O_275,N_25770,N_27811);
nor UO_276 (O_276,N_26949,N_29061);
nand UO_277 (O_277,N_26954,N_24649);
and UO_278 (O_278,N_29845,N_27137);
xor UO_279 (O_279,N_28547,N_27046);
nand UO_280 (O_280,N_25063,N_24998);
nand UO_281 (O_281,N_25967,N_27667);
nand UO_282 (O_282,N_29536,N_29453);
nor UO_283 (O_283,N_24318,N_26637);
xnor UO_284 (O_284,N_26752,N_26098);
nand UO_285 (O_285,N_28259,N_27151);
and UO_286 (O_286,N_24369,N_24549);
xor UO_287 (O_287,N_28239,N_29686);
nand UO_288 (O_288,N_29514,N_27177);
or UO_289 (O_289,N_24028,N_27815);
and UO_290 (O_290,N_25175,N_29517);
nand UO_291 (O_291,N_25439,N_28704);
and UO_292 (O_292,N_26581,N_26689);
and UO_293 (O_293,N_25420,N_28710);
and UO_294 (O_294,N_28061,N_29397);
nor UO_295 (O_295,N_29470,N_27632);
or UO_296 (O_296,N_26248,N_25582);
and UO_297 (O_297,N_26000,N_24860);
nor UO_298 (O_298,N_28300,N_24089);
nand UO_299 (O_299,N_25236,N_29288);
or UO_300 (O_300,N_26357,N_28994);
and UO_301 (O_301,N_29905,N_28862);
nor UO_302 (O_302,N_29491,N_29405);
and UO_303 (O_303,N_29279,N_24011);
or UO_304 (O_304,N_27047,N_27983);
or UO_305 (O_305,N_28126,N_28914);
or UO_306 (O_306,N_26722,N_27165);
xor UO_307 (O_307,N_27327,N_28761);
xor UO_308 (O_308,N_26903,N_28987);
and UO_309 (O_309,N_24733,N_29995);
or UO_310 (O_310,N_25731,N_29524);
and UO_311 (O_311,N_28456,N_29412);
or UO_312 (O_312,N_24085,N_24600);
xor UO_313 (O_313,N_28945,N_27063);
nor UO_314 (O_314,N_24380,N_26594);
or UO_315 (O_315,N_24909,N_27493);
xor UO_316 (O_316,N_28727,N_28367);
nand UO_317 (O_317,N_29677,N_26958);
or UO_318 (O_318,N_25245,N_26117);
nand UO_319 (O_319,N_27445,N_28863);
or UO_320 (O_320,N_26559,N_27709);
nor UO_321 (O_321,N_26669,N_25375);
and UO_322 (O_322,N_26871,N_27770);
or UO_323 (O_323,N_25581,N_24233);
or UO_324 (O_324,N_25914,N_28164);
or UO_325 (O_325,N_24499,N_28303);
xor UO_326 (O_326,N_26083,N_28793);
nor UO_327 (O_327,N_24949,N_29868);
and UO_328 (O_328,N_28878,N_29369);
nand UO_329 (O_329,N_27724,N_26891);
xor UO_330 (O_330,N_27847,N_25603);
xor UO_331 (O_331,N_27676,N_26342);
xor UO_332 (O_332,N_29828,N_24308);
nor UO_333 (O_333,N_27436,N_27684);
xnor UO_334 (O_334,N_25157,N_24819);
nand UO_335 (O_335,N_26760,N_26921);
nor UO_336 (O_336,N_26788,N_27630);
nor UO_337 (O_337,N_26567,N_27741);
nor UO_338 (O_338,N_27418,N_28100);
nor UO_339 (O_339,N_28501,N_26062);
nand UO_340 (O_340,N_24405,N_25311);
nand UO_341 (O_341,N_28283,N_28194);
and UO_342 (O_342,N_26316,N_26025);
xnor UO_343 (O_343,N_28122,N_26755);
or UO_344 (O_344,N_26441,N_26458);
nand UO_345 (O_345,N_24572,N_29572);
xor UO_346 (O_346,N_26773,N_25221);
xnor UO_347 (O_347,N_24816,N_28064);
nand UO_348 (O_348,N_28269,N_24726);
nand UO_349 (O_349,N_29528,N_29031);
nor UO_350 (O_350,N_26521,N_24553);
and UO_351 (O_351,N_28074,N_25984);
or UO_352 (O_352,N_28309,N_25898);
nand UO_353 (O_353,N_26508,N_29896);
nor UO_354 (O_354,N_26709,N_26885);
or UO_355 (O_355,N_24902,N_29641);
or UO_356 (O_356,N_25446,N_25557);
and UO_357 (O_357,N_24808,N_27044);
nand UO_358 (O_358,N_27571,N_29690);
nor UO_359 (O_359,N_26487,N_26005);
nand UO_360 (O_360,N_24456,N_26108);
and UO_361 (O_361,N_27477,N_27564);
and UO_362 (O_362,N_24051,N_25066);
nand UO_363 (O_363,N_27230,N_27368);
or UO_364 (O_364,N_28972,N_26116);
nor UO_365 (O_365,N_28843,N_26759);
and UO_366 (O_366,N_29798,N_24953);
and UO_367 (O_367,N_28638,N_27090);
or UO_368 (O_368,N_29165,N_25419);
nand UO_369 (O_369,N_27599,N_28976);
nor UO_370 (O_370,N_28123,N_26072);
xnor UO_371 (O_371,N_24835,N_24080);
or UO_372 (O_372,N_28240,N_26970);
or UO_373 (O_373,N_24469,N_24652);
xnor UO_374 (O_374,N_24408,N_29215);
xnor UO_375 (O_375,N_26857,N_25170);
nor UO_376 (O_376,N_29578,N_25230);
xor UO_377 (O_377,N_29923,N_28755);
xor UO_378 (O_378,N_26097,N_29184);
nand UO_379 (O_379,N_26329,N_29253);
or UO_380 (O_380,N_25758,N_26263);
nor UO_381 (O_381,N_26898,N_26152);
nor UO_382 (O_382,N_28651,N_25141);
nor UO_383 (O_383,N_29246,N_29710);
xnor UO_384 (O_384,N_26052,N_24091);
nand UO_385 (O_385,N_28026,N_27408);
or UO_386 (O_386,N_24322,N_24611);
xor UO_387 (O_387,N_26553,N_26085);
or UO_388 (O_388,N_27873,N_26159);
and UO_389 (O_389,N_29669,N_24621);
or UO_390 (O_390,N_24267,N_25925);
xor UO_391 (O_391,N_29801,N_29497);
xnor UO_392 (O_392,N_29920,N_28311);
xor UO_393 (O_393,N_27988,N_25671);
nor UO_394 (O_394,N_26136,N_24815);
and UO_395 (O_395,N_26841,N_26320);
nor UO_396 (O_396,N_27606,N_27356);
nand UO_397 (O_397,N_29871,N_25453);
and UO_398 (O_398,N_24769,N_29017);
or UO_399 (O_399,N_26420,N_24837);
xnor UO_400 (O_400,N_28066,N_27991);
nand UO_401 (O_401,N_25672,N_29223);
or UO_402 (O_402,N_27609,N_28981);
xor UO_403 (O_403,N_24447,N_27164);
or UO_404 (O_404,N_27882,N_24691);
or UO_405 (O_405,N_26818,N_29534);
nand UO_406 (O_406,N_26305,N_26902);
nor UO_407 (O_407,N_25070,N_24119);
xnor UO_408 (O_408,N_28946,N_28451);
and UO_409 (O_409,N_25207,N_28870);
nor UO_410 (O_410,N_24944,N_29291);
nor UO_411 (O_411,N_29882,N_29834);
nand UO_412 (O_412,N_26425,N_24612);
nand UO_413 (O_413,N_26194,N_27694);
or UO_414 (O_414,N_26061,N_25942);
nor UO_415 (O_415,N_26686,N_26312);
and UO_416 (O_416,N_26753,N_27924);
xnor UO_417 (O_417,N_25966,N_29894);
nand UO_418 (O_418,N_29639,N_26816);
nand UO_419 (O_419,N_28049,N_24155);
nand UO_420 (O_420,N_29044,N_28051);
or UO_421 (O_421,N_26783,N_27913);
and UO_422 (O_422,N_25804,N_24724);
xnor UO_423 (O_423,N_27687,N_28041);
xnor UO_424 (O_424,N_26003,N_26172);
or UO_425 (O_425,N_25189,N_24210);
and UO_426 (O_426,N_28357,N_28390);
nand UO_427 (O_427,N_28770,N_26247);
nor UO_428 (O_428,N_28241,N_26306);
or UO_429 (O_429,N_26925,N_27212);
and UO_430 (O_430,N_24594,N_27003);
nand UO_431 (O_431,N_24547,N_24782);
xnor UO_432 (O_432,N_28528,N_27052);
and UO_433 (O_433,N_26778,N_27935);
or UO_434 (O_434,N_24271,N_29180);
xnor UO_435 (O_435,N_24668,N_28917);
xor UO_436 (O_436,N_25330,N_29467);
or UO_437 (O_437,N_28027,N_29652);
nand UO_438 (O_438,N_24720,N_29888);
nor UO_439 (O_439,N_28650,N_24254);
nand UO_440 (O_440,N_29804,N_24146);
nor UO_441 (O_441,N_27343,N_27104);
nor UO_442 (O_442,N_28394,N_26747);
or UO_443 (O_443,N_26547,N_28700);
nand UO_444 (O_444,N_26338,N_28701);
xor UO_445 (O_445,N_24200,N_27566);
or UO_446 (O_446,N_24809,N_29052);
or UO_447 (O_447,N_29213,N_25913);
nand UO_448 (O_448,N_29416,N_28983);
or UO_449 (O_449,N_29211,N_27636);
and UO_450 (O_450,N_29294,N_27168);
nor UO_451 (O_451,N_24010,N_29823);
xnor UO_452 (O_452,N_25478,N_24859);
nor UO_453 (O_453,N_27693,N_24956);
nand UO_454 (O_454,N_27681,N_26053);
or UO_455 (O_455,N_24684,N_29880);
or UO_456 (O_456,N_24743,N_27699);
nand UO_457 (O_457,N_29311,N_24881);
nor UO_458 (O_458,N_25213,N_29171);
nand UO_459 (O_459,N_24540,N_25429);
nor UO_460 (O_460,N_27233,N_27407);
nor UO_461 (O_461,N_26740,N_24310);
or UO_462 (O_462,N_26990,N_24259);
xor UO_463 (O_463,N_26039,N_24825);
xor UO_464 (O_464,N_29985,N_24167);
nand UO_465 (O_465,N_26682,N_27633);
nand UO_466 (O_466,N_25886,N_25563);
or UO_467 (O_467,N_27325,N_27946);
and UO_468 (O_468,N_24706,N_25840);
nor UO_469 (O_469,N_27112,N_24270);
xnor UO_470 (O_470,N_26185,N_25515);
or UO_471 (O_471,N_25103,N_25058);
or UO_472 (O_472,N_29167,N_28386);
nor UO_473 (O_473,N_24730,N_26304);
nor UO_474 (O_474,N_28439,N_28465);
nor UO_475 (O_475,N_28158,N_25088);
nor UO_476 (O_476,N_24074,N_25127);
or UO_477 (O_477,N_28832,N_28982);
or UO_478 (O_478,N_28742,N_25909);
xnor UO_479 (O_479,N_26930,N_24900);
or UO_480 (O_480,N_28093,N_24431);
nor UO_481 (O_481,N_25659,N_25035);
nor UO_482 (O_482,N_28753,N_24521);
nand UO_483 (O_483,N_28658,N_28069);
and UO_484 (O_484,N_24787,N_24376);
nand UO_485 (O_485,N_24516,N_28351);
or UO_486 (O_486,N_25440,N_26707);
nand UO_487 (O_487,N_25156,N_27896);
nand UO_488 (O_488,N_25853,N_26182);
xnor UO_489 (O_489,N_26229,N_25593);
nor UO_490 (O_490,N_27133,N_25633);
and UO_491 (O_491,N_29962,N_29168);
and UO_492 (O_492,N_24643,N_26411);
xor UO_493 (O_493,N_26254,N_27043);
xor UO_494 (O_494,N_28748,N_29640);
or UO_495 (O_495,N_28070,N_28425);
xor UO_496 (O_496,N_24806,N_28502);
nor UO_497 (O_497,N_25959,N_29366);
or UO_498 (O_498,N_26474,N_24153);
or UO_499 (O_499,N_26257,N_26695);
xor UO_500 (O_500,N_29667,N_28374);
xnor UO_501 (O_501,N_27024,N_29622);
xor UO_502 (O_502,N_24163,N_24487);
nand UO_503 (O_503,N_24455,N_25708);
nand UO_504 (O_504,N_24034,N_26081);
or UO_505 (O_505,N_27185,N_24546);
xnor UO_506 (O_506,N_25433,N_28741);
nand UO_507 (O_507,N_29170,N_26799);
xnor UO_508 (O_508,N_26486,N_26401);
nor UO_509 (O_509,N_26176,N_28058);
nor UO_510 (O_510,N_29281,N_25927);
nand UO_511 (O_511,N_25105,N_25002);
or UO_512 (O_512,N_26195,N_25624);
xnor UO_513 (O_513,N_28937,N_29728);
or UO_514 (O_514,N_24370,N_24735);
and UO_515 (O_515,N_28513,N_24517);
and UO_516 (O_516,N_25550,N_29598);
and UO_517 (O_517,N_25528,N_26376);
xnor UO_518 (O_518,N_29192,N_26762);
nor UO_519 (O_519,N_25741,N_24871);
nand UO_520 (O_520,N_26088,N_27221);
xnor UO_521 (O_521,N_28422,N_26045);
xor UO_522 (O_522,N_24756,N_29110);
or UO_523 (O_523,N_27702,N_27839);
nand UO_524 (O_524,N_28286,N_24692);
nor UO_525 (O_525,N_27259,N_27258);
xor UO_526 (O_526,N_26975,N_24403);
and UO_527 (O_527,N_27409,N_25012);
nand UO_528 (O_528,N_29370,N_28315);
nand UO_529 (O_529,N_27421,N_26993);
nand UO_530 (O_530,N_26889,N_28082);
xor UO_531 (O_531,N_29904,N_29312);
nand UO_532 (O_532,N_26018,N_25024);
xor UO_533 (O_533,N_28571,N_28477);
nor UO_534 (O_534,N_27704,N_26096);
or UO_535 (O_535,N_24801,N_25696);
or UO_536 (O_536,N_27439,N_24587);
nor UO_537 (O_537,N_26210,N_28361);
xnor UO_538 (O_538,N_25756,N_28745);
xor UO_539 (O_539,N_26557,N_28737);
nor UO_540 (O_540,N_28539,N_26910);
or UO_541 (O_541,N_27091,N_29776);
and UO_542 (O_542,N_26562,N_24465);
nor UO_543 (O_543,N_28293,N_25818);
nor UO_544 (O_544,N_29262,N_24741);
or UO_545 (O_545,N_24767,N_29330);
xor UO_546 (O_546,N_24660,N_24289);
or UO_547 (O_547,N_29413,N_27838);
or UO_548 (O_548,N_27978,N_27219);
and UO_549 (O_549,N_24189,N_28810);
xor UO_550 (O_550,N_27295,N_29159);
nand UO_551 (O_551,N_26854,N_29106);
nand UO_552 (O_552,N_26922,N_24099);
nor UO_553 (O_553,N_28895,N_26798);
xor UO_554 (O_554,N_26057,N_24176);
and UO_555 (O_555,N_29917,N_24101);
xor UO_556 (O_556,N_24355,N_24458);
or UO_557 (O_557,N_24639,N_27795);
nor UO_558 (O_558,N_24983,N_28023);
and UO_559 (O_559,N_26164,N_29375);
nor UO_560 (O_560,N_28736,N_29097);
nand UO_561 (O_561,N_27858,N_25645);
nand UO_562 (O_562,N_29754,N_27193);
or UO_563 (O_563,N_25190,N_25778);
and UO_564 (O_564,N_25363,N_28885);
and UO_565 (O_565,N_26201,N_25333);
xor UO_566 (O_566,N_25314,N_28819);
nand UO_567 (O_567,N_24699,N_29131);
or UO_568 (O_568,N_26573,N_29697);
and UO_569 (O_569,N_26267,N_26706);
and UO_570 (O_570,N_27148,N_27417);
nor UO_571 (O_571,N_25312,N_28876);
and UO_572 (O_572,N_26736,N_28577);
xor UO_573 (O_573,N_29367,N_27462);
nand UO_574 (O_574,N_28178,N_25747);
and UO_575 (O_575,N_28722,N_25514);
xor UO_576 (O_576,N_24555,N_26270);
and UO_577 (O_577,N_26664,N_29377);
xor UO_578 (O_578,N_25359,N_27496);
nor UO_579 (O_579,N_26464,N_29734);
nand UO_580 (O_580,N_24577,N_24605);
and UO_581 (O_581,N_28672,N_29725);
nand UO_582 (O_582,N_29244,N_27580);
nor UO_583 (O_583,N_29579,N_29072);
and UO_584 (O_584,N_24017,N_26251);
xor UO_585 (O_585,N_24198,N_29282);
nor UO_586 (O_586,N_28242,N_24585);
or UO_587 (O_587,N_27114,N_28025);
and UO_588 (O_588,N_26679,N_24664);
and UO_589 (O_589,N_27871,N_25834);
nor UO_590 (O_590,N_25474,N_27162);
nand UO_591 (O_591,N_24887,N_29087);
or UO_592 (O_592,N_27197,N_26259);
nor UO_593 (O_593,N_27298,N_29778);
nand UO_594 (O_594,N_28867,N_29483);
nor UO_595 (O_595,N_27375,N_26745);
and UO_596 (O_596,N_29732,N_29986);
xnor UO_597 (O_597,N_27713,N_26272);
nand UO_598 (O_598,N_24103,N_25077);
nand UO_599 (O_599,N_29791,N_28010);
or UO_600 (O_600,N_26919,N_26653);
nand UO_601 (O_601,N_27348,N_28464);
or UO_602 (O_602,N_26418,N_24933);
nor UO_603 (O_603,N_25076,N_29519);
nand UO_604 (O_604,N_27404,N_28335);
nand UO_605 (O_605,N_29624,N_27352);
nor UO_606 (O_606,N_26456,N_25687);
nor UO_607 (O_607,N_26183,N_24570);
xnor UO_608 (O_608,N_24391,N_29847);
or UO_609 (O_609,N_27167,N_27199);
and UO_610 (O_610,N_26516,N_26957);
nand UO_611 (O_611,N_28882,N_27300);
and UO_612 (O_612,N_25087,N_28221);
xnor UO_613 (O_613,N_27476,N_29525);
or UO_614 (O_614,N_29657,N_27226);
nand UO_615 (O_615,N_28373,N_28919);
nand UO_616 (O_616,N_24762,N_26846);
or UO_617 (O_617,N_24070,N_28271);
nand UO_618 (O_618,N_27120,N_27428);
nand UO_619 (O_619,N_25677,N_27187);
nand UO_620 (O_620,N_28682,N_27243);
xor UO_621 (O_621,N_28666,N_25766);
nor UO_622 (O_622,N_26998,N_28362);
nor UO_623 (O_623,N_28706,N_28949);
nand UO_624 (O_624,N_24866,N_28204);
or UO_625 (O_625,N_29836,N_24793);
and UO_626 (O_626,N_24736,N_29596);
and UO_627 (O_627,N_29065,N_28336);
and UO_628 (O_628,N_25947,N_26361);
xnor UO_629 (O_629,N_28719,N_28548);
nand UO_630 (O_630,N_27358,N_27932);
and UO_631 (O_631,N_29105,N_27610);
and UO_632 (O_632,N_24357,N_27032);
nor UO_633 (O_633,N_25709,N_27989);
nand UO_634 (O_634,N_27470,N_29479);
and UO_635 (O_635,N_28779,N_28233);
or UO_636 (O_636,N_28618,N_24511);
or UO_637 (O_637,N_29951,N_26032);
nand UO_638 (O_638,N_27491,N_25541);
xnor UO_639 (O_639,N_29175,N_26200);
xnor UO_640 (O_640,N_26365,N_27579);
xnor UO_641 (O_641,N_28825,N_27626);
nand UO_642 (O_642,N_28800,N_27263);
or UO_643 (O_643,N_25669,N_25521);
nand UO_644 (O_644,N_29753,N_24162);
nand UO_645 (O_645,N_29237,N_25115);
and UO_646 (O_646,N_24876,N_27308);
and UO_647 (O_647,N_27268,N_25680);
xor UO_648 (O_648,N_27911,N_26663);
nor UO_649 (O_649,N_29123,N_26428);
xnor UO_650 (O_650,N_29093,N_26326);
nand UO_651 (O_651,N_25071,N_29862);
nor UO_652 (O_652,N_27471,N_27077);
nor UO_653 (O_653,N_24993,N_25471);
nor UO_654 (O_654,N_26124,N_28711);
and UO_655 (O_655,N_26667,N_27089);
nor UO_656 (O_656,N_26767,N_29461);
and UO_657 (O_657,N_25151,N_28615);
and UO_658 (O_658,N_25725,N_24829);
or UO_659 (O_659,N_25862,N_24423);
nor UO_660 (O_660,N_24044,N_25030);
nor UO_661 (O_661,N_27743,N_26895);
and UO_662 (O_662,N_24237,N_28726);
nand UO_663 (O_663,N_24940,N_25434);
nor UO_664 (O_664,N_25935,N_29832);
and UO_665 (O_665,N_26777,N_28613);
nor UO_666 (O_666,N_26169,N_27062);
or UO_667 (O_667,N_29559,N_26480);
nor UO_668 (O_668,N_29121,N_25727);
nor UO_669 (O_669,N_29229,N_28715);
and UO_670 (O_670,N_27503,N_28474);
nor UO_671 (O_671,N_24351,N_27129);
xnor UO_672 (O_672,N_28712,N_25428);
and UO_673 (O_673,N_24865,N_25202);
nor UO_674 (O_674,N_26206,N_25678);
xnor UO_675 (O_675,N_26240,N_26883);
nor UO_676 (O_676,N_24533,N_28521);
or UO_677 (O_677,N_26222,N_29070);
xnor UO_678 (O_678,N_28376,N_27696);
and UO_679 (O_679,N_26715,N_28892);
nand UO_680 (O_680,N_26285,N_29068);
nor UO_681 (O_681,N_24067,N_28413);
xor UO_682 (O_682,N_29621,N_25761);
and UO_683 (O_683,N_29296,N_25543);
xor UO_684 (O_684,N_28786,N_25569);
nor UO_685 (O_685,N_24794,N_28542);
xnor UO_686 (O_686,N_28034,N_27761);
or UO_687 (O_687,N_28327,N_28546);
or UO_688 (O_688,N_26971,N_25139);
nor UO_689 (O_689,N_26296,N_25140);
xor UO_690 (O_690,N_26112,N_27864);
or UO_691 (O_691,N_28683,N_27956);
xor UO_692 (O_692,N_26147,N_26158);
and UO_693 (O_693,N_25889,N_26843);
and UO_694 (O_694,N_29401,N_29944);
nand UO_695 (O_695,N_26224,N_27040);
or UO_696 (O_696,N_29318,N_24678);
nand UO_697 (O_697,N_29542,N_24315);
xnor UO_698 (O_698,N_26252,N_26021);
and UO_699 (O_699,N_25237,N_24630);
and UO_700 (O_700,N_27560,N_24161);
or UO_701 (O_701,N_26086,N_25192);
nand UO_702 (O_702,N_26119,N_28399);
or UO_703 (O_703,N_25995,N_28776);
or UO_704 (O_704,N_28809,N_24012);
nand UO_705 (O_705,N_26913,N_28028);
nand UO_706 (O_706,N_27438,N_25248);
xor UO_707 (O_707,N_24349,N_25054);
nand UO_708 (O_708,N_25225,N_26360);
and UO_709 (O_709,N_27096,N_25779);
xnor UO_710 (O_710,N_24754,N_29859);
nand UO_711 (O_711,N_26380,N_28193);
and UO_712 (O_712,N_25179,N_29515);
nor UO_713 (O_713,N_25268,N_24063);
and UO_714 (O_714,N_25777,N_24614);
or UO_715 (O_715,N_29573,N_26502);
xor UO_716 (O_716,N_27478,N_26126);
nand UO_717 (O_717,N_24886,N_29665);
nand UO_718 (O_718,N_25622,N_27314);
nand UO_719 (O_719,N_25900,N_26648);
or UO_720 (O_720,N_25064,N_27119);
nand UO_721 (O_721,N_28408,N_27405);
nor UO_722 (O_722,N_24875,N_28865);
nand UO_723 (O_723,N_28714,N_27690);
or UO_724 (O_724,N_25346,N_25017);
nand UO_725 (O_725,N_28595,N_27705);
xor UO_726 (O_726,N_26784,N_24745);
xor UO_727 (O_727,N_27947,N_26463);
and UO_728 (O_728,N_24526,N_26028);
xor UO_729 (O_729,N_27979,N_27857);
and UO_730 (O_730,N_25564,N_28047);
nand UO_731 (O_731,N_25887,N_24031);
and UO_732 (O_732,N_29004,N_29781);
xnor UO_733 (O_733,N_28075,N_25850);
or UO_734 (O_734,N_26070,N_25193);
nor UO_735 (O_735,N_24655,N_27716);
nand UO_736 (O_736,N_27149,N_28482);
nand UO_737 (O_737,N_26587,N_25369);
or UO_738 (O_738,N_28991,N_26996);
nand UO_739 (O_739,N_26630,N_27251);
nor UO_740 (O_740,N_26692,N_25338);
nor UO_741 (O_741,N_24175,N_26494);
or UO_742 (O_742,N_25352,N_25618);
and UO_743 (O_743,N_25805,N_27028);
or UO_744 (O_744,N_25837,N_25751);
nor UO_745 (O_745,N_28826,N_24117);
nand UO_746 (O_746,N_28404,N_28993);
nand UO_747 (O_747,N_25449,N_26478);
nand UO_748 (O_748,N_29512,N_28435);
xor UO_749 (O_749,N_24147,N_29893);
and UO_750 (O_750,N_27551,N_28050);
nand UO_751 (O_751,N_29129,N_27914);
or UO_752 (O_752,N_26469,N_24437);
and UO_753 (O_753,N_29362,N_26708);
and UO_754 (O_754,N_26870,N_28036);
nor UO_755 (O_755,N_24779,N_26107);
nand UO_756 (O_756,N_28631,N_25399);
nor UO_757 (O_757,N_27782,N_26043);
nor UO_758 (O_758,N_25062,N_28364);
or UO_759 (O_759,N_26860,N_29796);
nand UO_760 (O_760,N_25604,N_26786);
nor UO_761 (O_761,N_25318,N_24784);
nand UO_762 (O_762,N_24402,N_27802);
nor UO_763 (O_763,N_25211,N_26807);
and UO_764 (O_764,N_28402,N_25908);
xor UO_765 (O_765,N_26037,N_24247);
or UO_766 (O_766,N_26748,N_26955);
or UO_767 (O_767,N_25567,N_26554);
nor UO_768 (O_768,N_27403,N_27785);
nand UO_769 (O_769,N_25029,N_26207);
nand UO_770 (O_770,N_27264,N_26742);
nor UO_771 (O_771,N_26504,N_27055);
nand UO_772 (O_772,N_24569,N_24734);
and UO_773 (O_773,N_27053,N_27099);
nor UO_774 (O_774,N_28540,N_26241);
xor UO_775 (O_775,N_29285,N_27600);
or UO_776 (O_776,N_29963,N_27015);
or UO_777 (O_777,N_24810,N_24676);
xnor UO_778 (O_778,N_27182,N_28545);
and UO_779 (O_779,N_25466,N_28887);
xor UO_780 (O_780,N_27862,N_26964);
or UO_781 (O_781,N_27440,N_29113);
and UO_782 (O_782,N_25529,N_28530);
nor UO_783 (O_783,N_26994,N_26065);
nand UO_784 (O_784,N_24564,N_25901);
or UO_785 (O_785,N_25998,N_27650);
xnor UO_786 (O_786,N_24045,N_24695);
xnor UO_787 (O_787,N_29338,N_24215);
xnor UO_788 (O_788,N_26123,N_29591);
xor UO_789 (O_789,N_27755,N_25350);
nor UO_790 (O_790,N_27350,N_26135);
nor UO_791 (O_791,N_25824,N_28006);
or UO_792 (O_792,N_26577,N_26696);
and UO_793 (O_793,N_27156,N_24719);
nand UO_794 (O_794,N_25533,N_29992);
or UO_795 (O_795,N_24989,N_27992);
and UO_796 (O_796,N_29630,N_24197);
and UO_797 (O_797,N_29809,N_27139);
xor UO_798 (O_798,N_29408,N_29821);
xnor UO_799 (O_799,N_29727,N_27767);
nor UO_800 (O_800,N_24358,N_25585);
nand UO_801 (O_801,N_27831,N_27173);
nor UO_802 (O_802,N_26075,N_26063);
nand UO_803 (O_803,N_25074,N_27511);
nand UO_804 (O_804,N_24773,N_28429);
xor UO_805 (O_805,N_24716,N_29771);
and UO_806 (O_806,N_28142,N_29265);
and UO_807 (O_807,N_29872,N_26356);
nor UO_808 (O_808,N_25144,N_25187);
and UO_809 (O_809,N_29521,N_27468);
xor UO_810 (O_810,N_29916,N_26815);
xor UO_811 (O_811,N_26154,N_27645);
xnor UO_812 (O_812,N_25944,N_24891);
nor UO_813 (O_813,N_25395,N_28689);
xnor UO_814 (O_814,N_29835,N_24508);
nand UO_815 (O_815,N_27738,N_25026);
nand UO_816 (O_816,N_29661,N_27415);
nor UO_817 (O_817,N_25080,N_25767);
xor UO_818 (O_818,N_26539,N_29157);
or UO_819 (O_819,N_28459,N_28238);
xor UO_820 (O_820,N_24075,N_29452);
and UO_821 (O_821,N_29747,N_25423);
or UO_822 (O_822,N_28849,N_29372);
nor UO_823 (O_823,N_24603,N_24520);
or UO_824 (O_824,N_25681,N_28426);
xnor UO_825 (O_825,N_29190,N_25283);
nand UO_826 (O_826,N_25762,N_24061);
xnor UO_827 (O_827,N_24293,N_24132);
and UO_828 (O_828,N_27447,N_25782);
and UO_829 (O_829,N_26606,N_28920);
nor UO_830 (O_830,N_24066,N_26701);
and UO_831 (O_831,N_25473,N_25911);
or UO_832 (O_832,N_24874,N_25305);
or UO_833 (O_833,N_24645,N_29701);
xor UO_834 (O_834,N_25948,N_24127);
nor UO_835 (O_835,N_24901,N_24758);
xor UO_836 (O_836,N_26355,N_26256);
xor UO_837 (O_837,N_29731,N_27883);
and UO_838 (O_838,N_24831,N_28231);
or UO_839 (O_839,N_25639,N_26339);
nor UO_840 (O_840,N_25619,N_27917);
nand UO_841 (O_841,N_28687,N_27045);
nand UO_842 (O_842,N_26140,N_24996);
or UO_843 (O_843,N_24001,N_25068);
nor UO_844 (O_844,N_26026,N_28235);
and UO_845 (O_845,N_25576,N_28205);
nand UO_846 (O_846,N_24390,N_25821);
xor UO_847 (O_847,N_29360,N_28396);
or UO_848 (O_848,N_26331,N_25444);
nand UO_849 (O_849,N_26876,N_25553);
or UO_850 (O_850,N_24675,N_27427);
and UO_851 (O_851,N_24638,N_29691);
or UO_852 (O_852,N_29616,N_27744);
nand UO_853 (O_853,N_28492,N_29777);
nand UO_854 (O_854,N_28532,N_29547);
or UO_855 (O_855,N_24160,N_24713);
nand UO_856 (O_856,N_28130,N_27080);
or UO_857 (O_857,N_29424,N_29456);
and UO_858 (O_858,N_28214,N_24696);
or UO_859 (O_859,N_25742,N_25431);
xnor UO_860 (O_860,N_29225,N_28732);
or UO_861 (O_861,N_29434,N_28073);
nand UO_862 (O_862,N_26738,N_29436);
xor UO_863 (O_863,N_25749,N_26076);
or UO_864 (O_864,N_29802,N_26528);
or UO_865 (O_865,N_27302,N_27536);
xor UO_866 (O_866,N_28179,N_28321);
and UO_867 (O_867,N_25848,N_28781);
and UO_868 (O_868,N_28762,N_29286);
or UO_869 (O_869,N_24617,N_27625);
nand UO_870 (O_870,N_29928,N_25172);
xnor UO_871 (O_871,N_28052,N_24910);
or UO_872 (O_872,N_25579,N_25475);
nand UO_873 (O_873,N_29420,N_24663);
and UO_874 (O_874,N_24000,N_28391);
and UO_875 (O_875,N_24967,N_27643);
or UO_876 (O_876,N_26864,N_28044);
and UO_877 (O_877,N_25822,N_28926);
xor UO_878 (O_878,N_24799,N_25912);
nand UO_879 (O_879,N_26235,N_27961);
or UO_880 (O_880,N_29503,N_28278);
and UO_881 (O_881,N_25344,N_27619);
nand UO_882 (O_882,N_27396,N_26317);
nor UO_883 (O_883,N_25744,N_26666);
nor UO_884 (O_884,N_25490,N_28014);
and UO_885 (O_885,N_24602,N_26875);
xor UO_886 (O_886,N_24867,N_25711);
nor UO_887 (O_887,N_29866,N_25339);
nand UO_888 (O_888,N_26897,N_28078);
xor UO_889 (O_889,N_29335,N_25496);
and UO_890 (O_890,N_27441,N_25094);
and UO_891 (O_891,N_26909,N_24367);
or UO_892 (O_892,N_25654,N_27903);
xnor UO_893 (O_893,N_28551,N_24920);
or UO_894 (O_894,N_25208,N_27678);
and UO_895 (O_895,N_27584,N_24725);
nor UO_896 (O_896,N_28671,N_24169);
nand UO_897 (O_897,N_28763,N_29910);
and UO_898 (O_898,N_29425,N_29144);
or UO_899 (O_899,N_29325,N_24344);
and UO_900 (O_900,N_24841,N_24330);
and UO_901 (O_901,N_28868,N_28989);
xnor UO_902 (O_902,N_27073,N_26803);
nor UO_903 (O_903,N_28079,N_26228);
nor UO_904 (O_904,N_29009,N_29977);
and UO_905 (O_905,N_28648,N_27027);
and UO_906 (O_906,N_26277,N_25345);
nor UO_907 (O_907,N_24890,N_28695);
nor UO_908 (O_908,N_29989,N_24348);
nor UO_909 (O_909,N_28844,N_25547);
nand UO_910 (O_910,N_27562,N_27267);
nor UO_911 (O_911,N_24513,N_28602);
and UO_912 (O_912,N_25982,N_27454);
xor UO_913 (O_913,N_28643,N_25964);
xnor UO_914 (O_914,N_27615,N_25010);
and UO_915 (O_915,N_29141,N_27106);
nand UO_916 (O_916,N_28317,N_24328);
nor UO_917 (O_917,N_29876,N_25794);
nand UO_918 (O_918,N_26344,N_27442);
and UO_919 (O_919,N_26424,N_26541);
xor UO_920 (O_920,N_28106,N_24096);
and UO_921 (O_921,N_26264,N_26560);
or UO_922 (O_922,N_26907,N_26178);
nor UO_923 (O_923,N_29179,N_27706);
xor UO_924 (O_924,N_28022,N_24042);
and UO_925 (O_925,N_27557,N_28249);
or UO_926 (O_926,N_24049,N_24375);
and UO_927 (O_927,N_25148,N_29202);
or UO_928 (O_928,N_28043,N_24545);
and UO_929 (O_929,N_28953,N_27150);
and UO_930 (O_930,N_25476,N_25142);
or UO_931 (O_931,N_26268,N_28662);
nor UO_932 (O_932,N_27817,N_28686);
and UO_933 (O_933,N_29100,N_28854);
or UO_934 (O_934,N_27601,N_27257);
or UO_935 (O_935,N_24319,N_29447);
nor UO_936 (O_936,N_25823,N_28450);
or UO_937 (O_937,N_25307,N_27907);
nor UO_938 (O_938,N_27937,N_29076);
or UO_939 (O_939,N_24238,N_26916);
and UO_940 (O_940,N_25397,N_28557);
nor UO_941 (O_941,N_28104,N_26148);
nand UO_942 (O_942,N_27419,N_29484);
and UO_943 (O_943,N_25730,N_26362);
nor UO_944 (O_944,N_26789,N_27955);
and UO_945 (O_945,N_29935,N_28570);
nand UO_946 (O_946,N_24343,N_26352);
nand UO_947 (O_947,N_29763,N_29541);
xnor UO_948 (O_948,N_25717,N_28735);
and UO_949 (O_949,N_28108,N_29181);
and UO_950 (O_950,N_27980,N_26050);
or UO_951 (O_951,N_25154,N_27533);
and UO_952 (O_952,N_24016,N_29645);
and UO_953 (O_953,N_28254,N_29458);
and UO_954 (O_954,N_24942,N_29537);
xor UO_955 (O_955,N_25284,N_25875);
and UO_956 (O_956,N_26721,N_26963);
nand UO_957 (O_957,N_24068,N_27041);
xor UO_958 (O_958,N_26586,N_27435);
nand UO_959 (O_959,N_27220,N_29833);
nor UO_960 (O_960,N_27234,N_28216);
or UO_961 (O_961,N_26644,N_28485);
or UO_962 (O_962,N_25355,N_29689);
or UO_963 (O_963,N_24971,N_25282);
or UO_964 (O_964,N_29462,N_29926);
or UO_965 (O_965,N_24291,N_24043);
or UO_966 (O_966,N_26657,N_25736);
nor UO_967 (O_967,N_28600,N_24243);
nor UO_968 (O_968,N_29140,N_25111);
and UO_969 (O_969,N_28113,N_25849);
and UO_970 (O_970,N_26534,N_26704);
nor UO_971 (O_971,N_26121,N_28637);
xor UO_972 (O_972,N_26280,N_24763);
or UO_973 (O_973,N_24480,N_28558);
nand UO_974 (O_974,N_27050,N_26181);
and UO_975 (O_975,N_24579,N_26568);
or UO_976 (O_976,N_25735,N_25768);
nor UO_977 (O_977,N_27132,N_24751);
xor UO_978 (O_978,N_27532,N_28730);
nor UO_979 (O_979,N_27668,N_29432);
nor UO_980 (O_980,N_25099,N_25962);
nor UO_981 (O_981,N_26634,N_29590);
xnor UO_982 (O_982,N_28224,N_27347);
nand UO_983 (O_983,N_27381,N_24143);
nand UO_984 (O_984,N_26678,N_24821);
nand UO_985 (O_985,N_28861,N_24324);
and UO_986 (O_986,N_29151,N_28999);
nand UO_987 (O_987,N_27413,N_29049);
and UO_988 (O_988,N_24399,N_29321);
nand UO_989 (O_989,N_27054,N_29200);
nand UO_990 (O_990,N_28883,N_28567);
nand UO_991 (O_991,N_29251,N_24273);
and UO_992 (O_992,N_25536,N_29878);
or UO_993 (O_993,N_24582,N_25562);
nand UO_994 (O_994,N_27393,N_28533);
and UO_995 (O_995,N_27189,N_25943);
xor UO_996 (O_996,N_26170,N_25153);
nor UO_997 (O_997,N_27874,N_25755);
and UO_998 (O_998,N_27499,N_24260);
and UO_999 (O_999,N_25750,N_27153);
xor UO_1000 (O_1000,N_28288,N_29838);
or UO_1001 (O_1001,N_27799,N_24807);
nor UO_1002 (O_1002,N_24904,N_25532);
nor UO_1003 (O_1003,N_29704,N_24670);
xor UO_1004 (O_1004,N_29492,N_29599);
nand UO_1005 (O_1005,N_26218,N_27181);
or UO_1006 (O_1006,N_28936,N_26503);
nor UO_1007 (O_1007,N_28347,N_26768);
and UO_1008 (O_1008,N_27814,N_25306);
nor UO_1009 (O_1009,N_27611,N_24759);
and UO_1010 (O_1010,N_27222,N_28132);
nand UO_1011 (O_1011,N_26226,N_28636);
nor UO_1012 (O_1012,N_27056,N_27556);
or UO_1013 (O_1013,N_24915,N_29365);
xor UO_1014 (O_1014,N_29915,N_29230);
nor UO_1015 (O_1015,N_28133,N_27293);
nand UO_1016 (O_1016,N_28646,N_25916);
xnor UO_1017 (O_1017,N_26558,N_27289);
xor UO_1018 (O_1018,N_26952,N_29526);
and UO_1019 (O_1019,N_27122,N_25168);
or UO_1020 (O_1020,N_29016,N_24418);
or UO_1021 (O_1021,N_28417,N_27074);
or UO_1022 (O_1022,N_28494,N_29011);
nor UO_1023 (O_1023,N_26373,N_28840);
or UO_1024 (O_1024,N_28274,N_24173);
or UO_1025 (O_1025,N_28939,N_24978);
nand UO_1026 (O_1026,N_29489,N_26019);
or UO_1027 (O_1027,N_28992,N_27587);
or UO_1028 (O_1028,N_24905,N_29247);
and UO_1029 (O_1029,N_25923,N_25601);
nor UO_1030 (O_1030,N_25041,N_27449);
xnor UO_1031 (O_1031,N_24409,N_28799);
and UO_1032 (O_1032,N_24331,N_24620);
nor UO_1033 (O_1033,N_27904,N_29605);
nor UO_1034 (O_1034,N_26950,N_25506);
nand UO_1035 (O_1035,N_28096,N_24337);
xor UO_1036 (O_1036,N_27975,N_27344);
xor UO_1037 (O_1037,N_24095,N_26674);
and UO_1038 (O_1038,N_28766,N_28412);
nor UO_1039 (O_1039,N_26324,N_25763);
or UO_1040 (O_1040,N_26077,N_26238);
or UO_1041 (O_1041,N_24817,N_24593);
nand UO_1042 (O_1042,N_28030,N_29233);
and UO_1043 (O_1043,N_27519,N_29997);
nand UO_1044 (O_1044,N_24938,N_26811);
or UO_1045 (O_1045,N_27145,N_25937);
xor UO_1046 (O_1046,N_28146,N_25993);
xor UO_1047 (O_1047,N_27948,N_24223);
nand UO_1048 (O_1048,N_28750,N_28103);
xnor UO_1049 (O_1049,N_27590,N_28420);
or UO_1050 (O_1050,N_25548,N_24239);
nor UO_1051 (O_1051,N_24461,N_24277);
xnor UO_1052 (O_1052,N_27622,N_26873);
or UO_1053 (O_1053,N_24255,N_29448);
and UO_1054 (O_1054,N_25085,N_25705);
and UO_1055 (O_1055,N_24637,N_26089);
nor UO_1056 (O_1056,N_25780,N_27107);
and UO_1057 (O_1057,N_26237,N_26519);
nand UO_1058 (O_1058,N_27064,N_24872);
and UO_1059 (O_1059,N_29274,N_26585);
and UO_1060 (O_1060,N_24723,N_24436);
nor UO_1061 (O_1061,N_27644,N_25027);
xnor UO_1062 (O_1062,N_25803,N_27919);
xnor UO_1063 (O_1063,N_26345,N_28634);
or UO_1064 (O_1064,N_25728,N_28246);
or UO_1065 (O_1065,N_24098,N_29784);
xnor UO_1066 (O_1066,N_25276,N_29047);
nand UO_1067 (O_1067,N_26804,N_25130);
xor UO_1068 (O_1068,N_26467,N_24201);
or UO_1069 (O_1069,N_28931,N_27109);
and UO_1070 (O_1070,N_27432,N_24426);
and UO_1071 (O_1071,N_24406,N_26651);
or UO_1072 (O_1072,N_28284,N_27775);
and UO_1073 (O_1073,N_29714,N_27203);
and UO_1074 (O_1074,N_29780,N_27284);
xor UO_1075 (O_1075,N_24222,N_26999);
and UO_1076 (O_1076,N_26090,N_27270);
or UO_1077 (O_1077,N_26156,N_24199);
or UO_1078 (O_1078,N_26714,N_27218);
xor UO_1079 (O_1079,N_25739,N_25031);
xor UO_1080 (O_1080,N_25724,N_28971);
nor UO_1081 (O_1081,N_29114,N_27602);
xor UO_1082 (O_1082,N_24269,N_29363);
and UO_1083 (O_1083,N_24776,N_28940);
or UO_1084 (O_1084,N_24149,N_27786);
nand UO_1085 (O_1085,N_24165,N_28149);
nand UO_1086 (O_1086,N_28410,N_25827);
xnor UO_1087 (O_1087,N_26956,N_26621);
nor UO_1088 (O_1088,N_26834,N_28222);
xor UO_1089 (O_1089,N_24299,N_29908);
or UO_1090 (O_1090,N_26705,N_27926);
nor UO_1091 (O_1091,N_25819,N_29313);
or UO_1092 (O_1092,N_25607,N_27843);
nor UO_1093 (O_1093,N_26987,N_28228);
and UO_1094 (O_1094,N_24116,N_27169);
nor UO_1095 (O_1095,N_28675,N_29368);
nand UO_1096 (O_1096,N_26429,N_27017);
xnor UO_1097 (O_1097,N_25555,N_29032);
xnor UO_1098 (O_1098,N_27241,N_28446);
xor UO_1099 (O_1099,N_29889,N_25903);
nand UO_1100 (O_1100,N_27126,N_24925);
or UO_1101 (O_1101,N_25847,N_26231);
or UO_1102 (O_1102,N_26859,N_27897);
or UO_1103 (O_1103,N_28251,N_26036);
nor UO_1104 (O_1104,N_27127,N_24929);
nand UO_1105 (O_1105,N_28970,N_28838);
xnor UO_1106 (O_1106,N_28101,N_24301);
xor UO_1107 (O_1107,N_25164,N_25238);
nor UO_1108 (O_1108,N_26253,N_25009);
nor UO_1109 (O_1109,N_26935,N_26680);
or UO_1110 (O_1110,N_25285,N_24145);
nand UO_1111 (O_1111,N_29352,N_25924);
or UO_1112 (O_1112,N_28304,N_26354);
or UO_1113 (O_1113,N_28166,N_26792);
xor UO_1114 (O_1114,N_26590,N_25854);
nor UO_1115 (O_1115,N_28664,N_25273);
xnor UO_1116 (O_1116,N_29258,N_26455);
or UO_1117 (O_1117,N_26102,N_29115);
nor UO_1118 (O_1118,N_26540,N_25145);
or UO_1119 (O_1119,N_28795,N_24334);
nor UO_1120 (O_1120,N_27262,N_24705);
nand UO_1121 (O_1121,N_29724,N_24126);
or UO_1122 (O_1122,N_27364,N_25519);
nand UO_1123 (O_1123,N_24093,N_28340);
xor UO_1124 (O_1124,N_27671,N_29651);
nand UO_1125 (O_1125,N_26655,N_28171);
and UO_1126 (O_1126,N_26415,N_29744);
nor UO_1127 (O_1127,N_28503,N_24541);
nor UO_1128 (O_1128,N_26297,N_27583);
xor UO_1129 (O_1129,N_29188,N_26658);
nand UO_1130 (O_1130,N_29968,N_27663);
xor UO_1131 (O_1131,N_27578,N_27466);
or UO_1132 (O_1132,N_27071,N_26236);
or UO_1133 (O_1133,N_28641,N_25723);
xor UO_1134 (O_1134,N_29856,N_29495);
nand UO_1135 (O_1135,N_25393,N_27174);
nand UO_1136 (O_1136,N_27131,N_29395);
xor UO_1137 (O_1137,N_28219,N_28324);
or UO_1138 (O_1138,N_24347,N_28633);
nand UO_1139 (O_1139,N_29329,N_25461);
xnor UO_1140 (O_1140,N_25863,N_24964);
or UO_1141 (O_1141,N_29586,N_28801);
xor UO_1142 (O_1142,N_25465,N_25201);
nor UO_1143 (O_1143,N_28265,N_24383);
nor UO_1144 (O_1144,N_29852,N_24467);
nor UO_1145 (O_1145,N_27910,N_28174);
or UO_1146 (O_1146,N_27378,N_24092);
nor UO_1147 (O_1147,N_26084,N_29650);
and UO_1148 (O_1148,N_29419,N_27481);
and UO_1149 (O_1149,N_28203,N_28445);
nor UO_1150 (O_1150,N_26612,N_28544);
nand UO_1151 (O_1151,N_28837,N_26056);
nand UO_1152 (O_1152,N_27969,N_28729);
and UO_1153 (O_1153,N_26215,N_29881);
nand UO_1154 (O_1154,N_24039,N_24800);
nor UO_1155 (O_1155,N_27196,N_28804);
and UO_1156 (O_1156,N_29611,N_25504);
or UO_1157 (O_1157,N_29091,N_25643);
nand UO_1158 (O_1158,N_27823,N_25385);
or UO_1159 (O_1159,N_27306,N_27976);
nand UO_1160 (O_1160,N_25023,N_29972);
nand UO_1161 (O_1161,N_26030,N_26588);
xnor UO_1162 (O_1162,N_24628,N_28247);
xor UO_1163 (O_1163,N_27594,N_26041);
and UO_1164 (O_1164,N_29826,N_25846);
xor UO_1165 (O_1165,N_25025,N_27188);
or UO_1166 (O_1166,N_27389,N_25075);
xnor UO_1167 (O_1167,N_25649,N_26191);
and UO_1168 (O_1168,N_28244,N_29156);
xor UO_1169 (O_1169,N_29750,N_28690);
and UO_1170 (O_1170,N_24004,N_24481);
nand UO_1171 (O_1171,N_29478,N_28348);
or UO_1172 (O_1172,N_27646,N_28366);
nor UO_1173 (O_1173,N_25949,N_29884);
nor UO_1174 (O_1174,N_29073,N_24462);
and UO_1175 (O_1175,N_27783,N_25057);
or UO_1176 (O_1176,N_29602,N_27542);
or UO_1177 (O_1177,N_24632,N_27022);
xnor UO_1178 (O_1178,N_25244,N_24110);
nand UO_1179 (O_1179,N_26101,N_29505);
nor UO_1180 (O_1180,N_29374,N_26216);
xor UO_1181 (O_1181,N_26444,N_29064);
nand UO_1182 (O_1182,N_29646,N_26466);
xnor UO_1183 (O_1183,N_26413,N_25978);
nor UO_1184 (O_1184,N_26734,N_24640);
or UO_1185 (O_1185,N_29431,N_25997);
or UO_1186 (O_1186,N_24659,N_27485);
xnor UO_1187 (O_1187,N_26290,N_25126);
nand UO_1188 (O_1188,N_24917,N_29050);
or UO_1189 (O_1189,N_27400,N_25368);
xnor UO_1190 (O_1190,N_27049,N_28517);
nand UO_1191 (O_1191,N_26445,N_24498);
and UO_1192 (O_1192,N_28893,N_26485);
or UO_1193 (O_1193,N_28585,N_25946);
nand UO_1194 (O_1194,N_26570,N_24371);
nand UO_1195 (O_1195,N_24932,N_25408);
or UO_1196 (O_1196,N_28018,N_28565);
or UO_1197 (O_1197,N_24698,N_24803);
or UO_1198 (O_1198,N_24284,N_24439);
nand UO_1199 (O_1199,N_25203,N_27277);
nor UO_1200 (O_1200,N_29104,N_26435);
nand UO_1201 (O_1201,N_24928,N_24417);
and UO_1202 (O_1202,N_24084,N_27841);
or UO_1203 (O_1203,N_26622,N_25215);
and UO_1204 (O_1204,N_24580,N_25256);
and UO_1205 (O_1205,N_29563,N_29075);
nand UO_1206 (O_1206,N_28509,N_24654);
nand UO_1207 (O_1207,N_25327,N_28145);
and UO_1208 (O_1208,N_25969,N_28314);
nor UO_1209 (O_1209,N_24342,N_28060);
xnor UO_1210 (O_1210,N_25000,N_27038);
xor UO_1211 (O_1211,N_26106,N_28380);
nand UO_1212 (O_1212,N_25613,N_25799);
and UO_1213 (O_1213,N_25807,N_25438);
and UO_1214 (O_1214,N_25138,N_27929);
xor UO_1215 (O_1215,N_27689,N_24083);
xor UO_1216 (O_1216,N_25963,N_24610);
nor UO_1217 (O_1217,N_26641,N_28617);
nor UO_1218 (O_1218,N_29742,N_28984);
and UO_1219 (O_1219,N_28720,N_27920);
xnor UO_1220 (O_1220,N_29870,N_25329);
xor UO_1221 (O_1221,N_24855,N_27939);
xor UO_1222 (O_1222,N_24401,N_29255);
nand UO_1223 (O_1223,N_28594,N_29302);
xnor UO_1224 (O_1224,N_26465,N_25396);
and UO_1225 (O_1225,N_27887,N_28872);
nand UO_1226 (O_1226,N_27321,N_28856);
and UO_1227 (O_1227,N_29466,N_24120);
nor UO_1228 (O_1228,N_24623,N_27888);
nor UO_1229 (O_1229,N_28968,N_28744);
xnor UO_1230 (O_1230,N_29726,N_25162);
xor UO_1231 (O_1231,N_25098,N_25082);
xor UO_1232 (O_1232,N_24258,N_26261);
or UO_1233 (O_1233,N_28508,N_29078);
or UO_1234 (O_1234,N_27635,N_24475);
xnor UO_1235 (O_1235,N_27138,N_29193);
and UO_1236 (O_1236,N_24226,N_25452);
xor UO_1237 (O_1237,N_26013,N_25454);
nand UO_1238 (O_1238,N_24775,N_26143);
nand UO_1239 (O_1239,N_28962,N_28821);
nor UO_1240 (O_1240,N_25021,N_28379);
and UO_1241 (O_1241,N_25973,N_25260);
or UO_1242 (O_1242,N_27568,N_24241);
xnor UO_1243 (O_1243,N_25676,N_29081);
nand UO_1244 (O_1244,N_24868,N_25093);
xor UO_1245 (O_1245,N_29349,N_29385);
nor UO_1246 (O_1246,N_29993,N_26685);
or UO_1247 (O_1247,N_25242,N_24709);
nor UO_1248 (O_1248,N_26538,N_27729);
nand UO_1249 (O_1249,N_25599,N_26974);
xor UO_1250 (O_1250,N_26479,N_26403);
and UO_1251 (O_1251,N_29817,N_29913);
or UO_1252 (O_1252,N_24818,N_24490);
xor UO_1253 (O_1253,N_27207,N_27836);
xor UO_1254 (O_1254,N_29499,N_27544);
or UO_1255 (O_1255,N_27780,N_24429);
nand UO_1256 (O_1256,N_29197,N_25133);
nor UO_1257 (O_1257,N_24410,N_26615);
or UO_1258 (O_1258,N_26725,N_25630);
and UO_1259 (O_1259,N_25955,N_27102);
nand UO_1260 (O_1260,N_24228,N_24144);
nor UO_1261 (O_1261,N_24040,N_28467);
nor UO_1262 (O_1262,N_24943,N_26566);
nor UO_1263 (O_1263,N_25371,N_29535);
xor UO_1264 (O_1264,N_29772,N_28080);
nor UO_1265 (O_1265,N_29149,N_28167);
and UO_1266 (O_1266,N_29634,N_28415);
and UO_1267 (O_1267,N_26139,N_25623);
and UO_1268 (O_1268,N_24335,N_29345);
or UO_1269 (O_1269,N_28559,N_27342);
xor UO_1270 (O_1270,N_27206,N_27152);
nand UO_1271 (O_1271,N_25007,N_27385);
or UO_1272 (O_1272,N_25573,N_25361);
xnor UO_1273 (O_1273,N_27548,N_26163);
or UO_1274 (O_1274,N_26853,N_26911);
nand UO_1275 (O_1275,N_25481,N_29101);
and UO_1276 (O_1276,N_29975,N_25500);
nor UO_1277 (O_1277,N_26142,N_28094);
and UO_1278 (O_1278,N_29486,N_27921);
or UO_1279 (O_1279,N_24506,N_24869);
xnor UO_1280 (O_1280,N_29473,N_28276);
nor UO_1281 (O_1281,N_29150,N_26392);
xnor UO_1282 (O_1282,N_27225,N_28211);
nand UO_1283 (O_1283,N_26378,N_29404);
nor UO_1284 (O_1284,N_27058,N_25864);
nor UO_1285 (O_1285,N_28411,N_26437);
nor UO_1286 (O_1286,N_26620,N_24294);
xor UO_1287 (O_1287,N_24575,N_28812);
or UO_1288 (O_1288,N_24830,N_26782);
or UO_1289 (O_1289,N_28038,N_25951);
or UO_1290 (O_1290,N_26225,N_27641);
and UO_1291 (O_1291,N_25865,N_28679);
xor UO_1292 (O_1292,N_24750,N_26203);
xor UO_1293 (O_1293,N_27186,N_25956);
xnor UO_1294 (O_1294,N_25653,N_24804);
nor UO_1295 (O_1295,N_27191,N_27776);
or UO_1296 (O_1296,N_25090,N_27146);
or UO_1297 (O_1297,N_28568,N_26209);
and UO_1298 (O_1298,N_28655,N_26942);
nand UO_1299 (O_1299,N_25275,N_27213);
nor UO_1300 (O_1300,N_26276,N_26941);
xor UO_1301 (O_1301,N_26448,N_26167);
or UO_1302 (O_1302,N_29194,N_24936);
and UO_1303 (O_1303,N_24888,N_26847);
xnor UO_1304 (O_1304,N_24535,N_29971);
and UO_1305 (O_1305,N_26618,N_29508);
and UO_1306 (O_1306,N_29108,N_29565);
or UO_1307 (O_1307,N_26265,N_29819);
nand UO_1308 (O_1308,N_24501,N_27208);
or UO_1309 (O_1309,N_28504,N_24681);
xor UO_1310 (O_1310,N_25938,N_27620);
and UO_1311 (O_1311,N_26212,N_24822);
xor UO_1312 (O_1312,N_27305,N_29664);
or UO_1313 (O_1313,N_25608,N_25648);
xnor UO_1314 (O_1314,N_24114,N_29987);
nand UO_1315 (O_1315,N_25235,N_27581);
xnor UO_1316 (O_1316,N_25907,N_26670);
nor UO_1317 (O_1317,N_24519,N_26278);
nor UO_1318 (O_1318,N_25707,N_28307);
xnor UO_1319 (O_1319,N_29007,N_27136);
xnor UO_1320 (O_1320,N_24616,N_24240);
and UO_1321 (O_1321,N_28693,N_24747);
or UO_1322 (O_1322,N_24926,N_25167);
or UO_1323 (O_1323,N_24771,N_25781);
and UO_1324 (O_1324,N_27025,N_25740);
and UO_1325 (O_1325,N_27184,N_27242);
xor UO_1326 (O_1326,N_26796,N_26984);
or UO_1327 (O_1327,N_26500,N_25436);
or UO_1328 (O_1328,N_29013,N_29787);
nor UO_1329 (O_1329,N_27322,N_24544);
and UO_1330 (O_1330,N_28684,N_29277);
and UO_1331 (O_1331,N_26336,N_24362);
or UO_1332 (O_1332,N_25006,N_29900);
nand UO_1333 (O_1333,N_28177,N_25658);
nor UO_1334 (O_1334,N_28331,N_26966);
xnor UO_1335 (O_1335,N_27157,N_29355);
and UO_1336 (O_1336,N_27521,N_24014);
nand UO_1337 (O_1337,N_27915,N_27754);
or UO_1338 (O_1338,N_24636,N_28911);
nor UO_1339 (O_1339,N_28965,N_25673);
and UO_1340 (O_1340,N_26104,N_28213);
nand UO_1341 (O_1341,N_27720,N_26289);
and UO_1342 (O_1342,N_24690,N_29056);
nor UO_1343 (O_1343,N_27510,N_27682);
and UO_1344 (O_1344,N_27100,N_28586);
and UO_1345 (O_1345,N_27201,N_25011);
xnor UO_1346 (O_1346,N_25531,N_27085);
nor UO_1347 (O_1347,N_29831,N_25899);
xor UO_1348 (O_1348,N_26452,N_24183);
and UO_1349 (O_1349,N_25965,N_25296);
and UO_1350 (O_1350,N_25477,N_29010);
or UO_1351 (O_1351,N_26409,N_26291);
or UO_1352 (O_1352,N_26308,N_29873);
or UO_1353 (O_1353,N_27211,N_24156);
nor UO_1354 (O_1354,N_27796,N_26839);
nand UO_1355 (O_1355,N_26067,N_26603);
nor UO_1356 (O_1356,N_29768,N_25754);
and UO_1357 (O_1357,N_28621,N_25389);
or UO_1358 (O_1358,N_29487,N_25616);
nand UO_1359 (O_1359,N_28156,N_25210);
nor UO_1360 (O_1360,N_27324,N_28029);
xor UO_1361 (O_1361,N_25176,N_26166);
and UO_1362 (O_1362,N_24325,N_27088);
and UO_1363 (O_1363,N_29241,N_28039);
and UO_1364 (O_1364,N_25411,N_25841);
or UO_1365 (O_1365,N_24135,N_24527);
nor UO_1366 (O_1366,N_26472,N_29555);
and UO_1367 (O_1367,N_24752,N_29800);
or UO_1368 (O_1368,N_28255,N_25197);
or UO_1369 (O_1369,N_24048,N_29220);
or UO_1370 (O_1370,N_25114,N_27453);
nor UO_1371 (O_1371,N_28312,N_28301);
nor UO_1372 (O_1372,N_27291,N_28948);
and UO_1373 (O_1373,N_29292,N_25059);
and UO_1374 (O_1374,N_29843,N_26576);
and UO_1375 (O_1375,N_26703,N_29609);
nor UO_1376 (O_1376,N_25259,N_27598);
and UO_1377 (O_1377,N_27877,N_25300);
xnor UO_1378 (O_1378,N_26133,N_26171);
xnor UO_1379 (O_1379,N_27287,N_26848);
nor UO_1380 (O_1380,N_29088,N_25413);
nand UO_1381 (O_1381,N_25467,N_28519);
nand UO_1382 (O_1382,N_24985,N_28829);
xor UO_1383 (O_1383,N_27819,N_26607);
or UO_1384 (O_1384,N_27204,N_24245);
nor UO_1385 (O_1385,N_25401,N_27501);
xor UO_1386 (O_1386,N_28263,N_24812);
or UO_1387 (O_1387,N_24647,N_27773);
or UO_1388 (O_1388,N_24460,N_28784);
nand UO_1389 (O_1389,N_25571,N_25825);
and UO_1390 (O_1390,N_29501,N_24090);
and UO_1391 (O_1391,N_29827,N_29471);
nor UO_1392 (O_1392,N_29527,N_28563);
nor UO_1393 (O_1393,N_29227,N_27235);
nor UO_1394 (O_1394,N_26313,N_29046);
or UO_1395 (O_1395,N_26614,N_26874);
nand UO_1396 (O_1396,N_26029,N_25412);
nand UO_1397 (O_1397,N_24148,N_24914);
and UO_1398 (O_1398,N_27995,N_24682);
and UO_1399 (O_1399,N_24994,N_27860);
xor UO_1400 (O_1400,N_28871,N_24710);
xor UO_1401 (O_1401,N_26439,N_27500);
and UO_1402 (O_1402,N_26080,N_29779);
nand UO_1403 (O_1403,N_24209,N_28550);
or UO_1404 (O_1404,N_24073,N_26719);
xor UO_1405 (O_1405,N_24542,N_26165);
nand UO_1406 (O_1406,N_29480,N_24574);
nand UO_1407 (O_1407,N_27810,N_26593);
nand UO_1408 (O_1408,N_26087,N_27647);
nand UO_1409 (O_1409,N_25617,N_28452);
nand UO_1410 (O_1410,N_26780,N_28371);
and UO_1411 (O_1411,N_24746,N_27256);
nand UO_1412 (O_1412,N_25719,N_27031);
nor UO_1413 (O_1413,N_28659,N_27789);
xnor UO_1414 (O_1414,N_28031,N_24565);
nand UO_1415 (O_1415,N_25104,N_26162);
nor UO_1416 (O_1416,N_26457,N_24007);
nor UO_1417 (O_1417,N_29507,N_29195);
or UO_1418 (O_1418,N_25123,N_27900);
xnor UO_1419 (O_1419,N_26031,N_29658);
xnor UO_1420 (O_1420,N_28596,N_24861);
nor UO_1421 (O_1421,N_29875,N_26334);
or UO_1422 (O_1422,N_28363,N_29059);
nand UO_1423 (O_1423,N_28583,N_25631);
nor UO_1424 (O_1424,N_26776,N_24139);
nand UO_1425 (O_1425,N_29681,N_27261);
xor UO_1426 (O_1426,N_29219,N_26358);
nor UO_1427 (O_1427,N_27144,N_25325);
nor UO_1428 (O_1428,N_29619,N_25981);
or UO_1429 (O_1429,N_29699,N_27332);
and UO_1430 (O_1430,N_29392,N_29998);
xnor UO_1431 (O_1431,N_24323,N_29636);
or UO_1432 (O_1432,N_24615,N_25872);
nand UO_1433 (O_1433,N_28783,N_28433);
or UO_1434 (O_1434,N_28888,N_25110);
or UO_1435 (O_1435,N_29764,N_29445);
or UO_1436 (O_1436,N_29688,N_29015);
nor UO_1437 (O_1437,N_25056,N_25146);
xnor UO_1438 (O_1438,N_26524,N_29822);
and UO_1439 (O_1439,N_28199,N_27430);
and UO_1440 (O_1440,N_28170,N_29122);
or UO_1441 (O_1441,N_24187,N_26199);
nor UO_1442 (O_1442,N_24608,N_24958);
or UO_1443 (O_1443,N_27642,N_24715);
or UO_1444 (O_1444,N_24505,N_24976);
nand UO_1445 (O_1445,N_26008,N_29199);
and UO_1446 (O_1446,N_28816,N_26011);
nand UO_1447 (O_1447,N_27708,N_27280);
nand UO_1448 (O_1448,N_29337,N_27930);
nor UO_1449 (O_1449,N_24278,N_26493);
or UO_1450 (O_1450,N_28381,N_24984);
or UO_1451 (O_1451,N_24055,N_24972);
and UO_1452 (O_1452,N_27086,N_28796);
or UO_1453 (O_1453,N_28470,N_26779);
nand UO_1454 (O_1454,N_27472,N_25545);
or UO_1455 (O_1455,N_29592,N_25871);
or UO_1456 (O_1456,N_27360,N_25231);
nand UO_1457 (O_1457,N_25656,N_29391);
nor UO_1458 (O_1458,N_24478,N_29250);
xnor UO_1459 (O_1459,N_25644,N_27029);
or UO_1460 (O_1460,N_27971,N_28090);
and UO_1461 (O_1461,N_26442,N_27891);
nor UO_1462 (O_1462,N_25264,N_26694);
xnor UO_1463 (O_1463,N_27255,N_24262);
and UO_1464 (O_1464,N_27340,N_25258);
nor UO_1465 (O_1465,N_29124,N_28835);
and UO_1466 (O_1466,N_29062,N_25600);
or UO_1467 (O_1467,N_28505,N_26813);
nor UO_1468 (O_1468,N_27790,N_27842);
or UO_1469 (O_1469,N_29953,N_25482);
or UO_1470 (O_1470,N_26468,N_27311);
and UO_1471 (O_1471,N_29423,N_27429);
or UO_1472 (O_1472,N_25771,N_27546);
or UO_1473 (O_1473,N_29378,N_24438);
and UO_1474 (O_1474,N_27384,N_25421);
and UO_1475 (O_1475,N_25990,N_26427);
nor UO_1476 (O_1476,N_28874,N_29849);
xor UO_1477 (O_1477,N_25611,N_28483);
or UO_1478 (O_1478,N_26382,N_26066);
or UO_1479 (O_1479,N_26451,N_29815);
and UO_1480 (O_1480,N_24884,N_28454);
and UO_1481 (O_1481,N_28975,N_27008);
xor UO_1482 (O_1482,N_24677,N_24333);
and UO_1483 (O_1483,N_27498,N_28349);
nand UO_1484 (O_1484,N_26481,N_29504);
nor UO_1485 (O_1485,N_27617,N_26625);
and UO_1486 (O_1486,N_25488,N_25926);
and UO_1487 (O_1487,N_25272,N_24642);
or UO_1488 (O_1488,N_25299,N_27964);
nor UO_1489 (O_1489,N_24563,N_29006);
nor UO_1490 (O_1490,N_29532,N_29216);
nand UO_1491 (O_1491,N_25317,N_27117);
or UO_1492 (O_1492,N_26131,N_27732);
and UO_1493 (O_1493,N_24283,N_26369);
xor UO_1494 (O_1494,N_29960,N_29758);
and UO_1495 (O_1495,N_29970,N_29617);
or UO_1496 (O_1496,N_29973,N_28723);
or UO_1497 (O_1497,N_29705,N_26179);
nand UO_1498 (O_1498,N_29094,N_29411);
or UO_1499 (O_1499,N_29550,N_26713);
xor UO_1500 (O_1500,N_28587,N_25323);
xnor UO_1501 (O_1501,N_29846,N_24026);
xnor UO_1502 (O_1502,N_26303,N_24494);
and UO_1503 (O_1503,N_25107,N_28448);
xnor UO_1504 (O_1504,N_28200,N_24107);
and UO_1505 (O_1505,N_29919,N_29382);
xnor UO_1506 (O_1506,N_24685,N_29583);
or UO_1507 (O_1507,N_29675,N_24261);
nand UO_1508 (O_1508,N_27391,N_26537);
nor UO_1509 (O_1509,N_24633,N_29400);
nor UO_1510 (O_1510,N_25051,N_27820);
and UO_1511 (O_1511,N_28649,N_29544);
nor UO_1512 (O_1512,N_26422,N_29943);
and UO_1513 (O_1513,N_24130,N_27715);
or UO_1514 (O_1514,N_25279,N_26561);
nor UO_1515 (O_1515,N_24321,N_29715);
nor UO_1516 (O_1516,N_29511,N_26273);
or UO_1517 (O_1517,N_28905,N_27214);
xor UO_1518 (O_1518,N_27909,N_27655);
nor UO_1519 (O_1519,N_26924,N_27246);
nand UO_1520 (O_1520,N_29718,N_24378);
nand UO_1521 (O_1521,N_29500,N_28511);
xor UO_1522 (O_1522,N_29069,N_25136);
nand UO_1523 (O_1523,N_28774,N_29222);
and UO_1524 (O_1524,N_26017,N_24562);
nand UO_1525 (O_1525,N_27778,N_29469);
nand UO_1526 (O_1526,N_29948,N_24778);
or UO_1527 (O_1527,N_25790,N_24124);
nor UO_1528 (O_1528,N_27020,N_29568);
xor UO_1529 (O_1529,N_29647,N_29117);
nand UO_1530 (O_1530,N_25893,N_29112);
or UO_1531 (O_1531,N_29136,N_27357);
nand UO_1532 (O_1532,N_26404,N_25561);
nor UO_1533 (O_1533,N_26812,N_25435);
nor UO_1534 (O_1534,N_28486,N_24186);
xnor UO_1535 (O_1535,N_25147,N_29957);
or UO_1536 (O_1536,N_26284,N_25291);
nor UO_1537 (O_1537,N_27275,N_28440);
and UO_1538 (O_1538,N_24599,N_26829);
xnor UO_1539 (O_1539,N_25120,N_29051);
and UO_1540 (O_1540,N_25253,N_24986);
or UO_1541 (O_1541,N_28626,N_28721);
nor UO_1542 (O_1542,N_27570,N_26991);
xor UO_1543 (O_1543,N_27036,N_29224);
nor UO_1544 (O_1544,N_24264,N_24805);
nor UO_1545 (O_1545,N_24538,N_26877);
nand UO_1546 (O_1546,N_26596,N_28157);
nand UO_1547 (O_1547,N_29818,N_27901);
or UO_1548 (O_1548,N_25706,N_27923);
or UO_1549 (O_1549,N_28161,N_25495);
or UO_1550 (O_1550,N_26060,N_29198);
nand UO_1551 (O_1551,N_27670,N_25920);
nor UO_1552 (O_1552,N_26507,N_28065);
nor UO_1553 (O_1553,N_25016,N_29446);
or UO_1554 (O_1554,N_29270,N_27135);
or UO_1555 (O_1555,N_27108,N_27763);
or UO_1556 (O_1556,N_29587,N_27140);
and UO_1557 (O_1557,N_27081,N_28298);
and UO_1558 (O_1558,N_26532,N_25483);
or UO_1559 (O_1559,N_29454,N_24728);
nand UO_1560 (O_1560,N_24111,N_28444);
or UO_1561 (O_1561,N_25079,N_27443);
nor UO_1562 (O_1562,N_28215,N_24332);
nand UO_1563 (O_1563,N_25738,N_25018);
xor UO_1564 (O_1564,N_29485,N_27905);
nand UO_1565 (O_1565,N_24507,N_29952);
nor UO_1566 (O_1566,N_27367,N_26388);
and UO_1567 (O_1567,N_28771,N_25764);
xor UO_1568 (O_1568,N_27098,N_25831);
and UO_1569 (O_1569,N_28181,N_25455);
nor UO_1570 (O_1570,N_26190,N_26269);
xor UO_1571 (O_1571,N_27070,N_26918);
nand UO_1572 (O_1572,N_29912,N_27192);
or UO_1573 (O_1573,N_28751,N_25851);
xor UO_1574 (O_1574,N_26490,N_28929);
and UO_1575 (O_1575,N_27534,N_25941);
nand UO_1576 (O_1576,N_29678,N_27737);
xnor UO_1577 (O_1577,N_26724,N_26406);
nor UO_1578 (O_1578,N_26574,N_25044);
nor UO_1579 (O_1579,N_26866,N_28339);
xnor UO_1580 (O_1580,N_25682,N_24216);
xor UO_1581 (O_1581,N_25974,N_29264);
nor UO_1582 (O_1582,N_24606,N_28436);
xor UO_1583 (O_1583,N_28531,N_24327);
xnor UO_1584 (O_1584,N_26826,N_28574);
or UO_1585 (O_1585,N_29558,N_25720);
xor UO_1586 (O_1586,N_25460,N_26851);
nor UO_1587 (O_1587,N_28966,N_28037);
and UO_1588 (O_1588,N_24421,N_26125);
xnor UO_1589 (O_1589,N_27908,N_24191);
and UO_1590 (O_1590,N_24428,N_27248);
xor UO_1591 (O_1591,N_24064,N_27504);
xor UO_1592 (O_1592,N_26688,N_29383);
and UO_1593 (O_1593,N_24047,N_25558);
nand UO_1594 (O_1594,N_26132,N_28588);
xor UO_1595 (O_1595,N_24297,N_29263);
or UO_1596 (O_1596,N_28676,N_28990);
nor UO_1597 (O_1597,N_27359,N_24658);
or UO_1598 (O_1598,N_26069,N_24838);
or UO_1599 (O_1599,N_29333,N_28279);
xor UO_1600 (O_1600,N_24483,N_24788);
xnor UO_1601 (O_1601,N_26536,N_25028);
and UO_1602 (O_1602,N_27093,N_26221);
or UO_1603 (O_1603,N_25539,N_29147);
or UO_1604 (O_1604,N_29863,N_24489);
nand UO_1605 (O_1605,N_27007,N_26509);
or UO_1606 (O_1606,N_26155,N_24218);
nand UO_1607 (O_1607,N_29315,N_28318);
nor UO_1608 (O_1608,N_24813,N_24607);
xor UO_1609 (O_1609,N_24523,N_27685);
xor UO_1610 (O_1610,N_29232,N_28692);
xnor UO_1611 (O_1611,N_29608,N_24464);
and UO_1612 (O_1612,N_26180,N_28757);
nand UO_1613 (O_1613,N_25877,N_24112);
or UO_1614 (O_1614,N_26064,N_29373);
xor UO_1615 (O_1615,N_29803,N_28912);
nor UO_1616 (O_1616,N_28526,N_28305);
or UO_1617 (O_1617,N_26929,N_28739);
xnor UO_1618 (O_1618,N_28086,N_29540);
nand UO_1619 (O_1619,N_29967,N_28627);
xnor UO_1620 (O_1620,N_28902,N_27448);
nor UO_1621 (O_1621,N_26730,N_25020);
nand UO_1622 (O_1622,N_24897,N_27508);
xnor UO_1623 (O_1623,N_24786,N_25331);
nand UO_1624 (O_1624,N_29533,N_28141);
xnor UO_1625 (O_1625,N_29212,N_28005);
or UO_1626 (O_1626,N_28344,N_24313);
nand UO_1627 (O_1627,N_24444,N_26969);
or UO_1628 (O_1628,N_28488,N_24192);
nor UO_1629 (O_1629,N_28220,N_26529);
xnor UO_1630 (O_1630,N_27769,N_26861);
and UO_1631 (O_1631,N_28189,N_29706);
nand UO_1632 (O_1632,N_29414,N_24729);
xor UO_1633 (O_1633,N_28124,N_29797);
or UO_1634 (O_1634,N_28000,N_24281);
and UO_1635 (O_1635,N_28673,N_26014);
xnor UO_1636 (O_1636,N_24424,N_24341);
nor UO_1637 (O_1637,N_28306,N_29347);
or UO_1638 (O_1638,N_26896,N_25702);
nand UO_1639 (O_1639,N_28645,N_28660);
nor UO_1640 (O_1640,N_26808,N_28153);
nand UO_1641 (O_1641,N_25888,N_24836);
or UO_1642 (O_1642,N_27797,N_28667);
nor UO_1643 (O_1643,N_25186,N_26764);
or UO_1644 (O_1644,N_28537,N_29086);
xnor UO_1645 (O_1645,N_25358,N_27634);
and UO_1646 (O_1646,N_25388,N_26840);
nand UO_1647 (O_1647,N_27527,N_29036);
and UO_1648 (O_1648,N_28003,N_26677);
or UO_1649 (O_1649,N_26407,N_27898);
xnor UO_1650 (O_1650,N_26613,N_24988);
or UO_1651 (O_1651,N_26330,N_24442);
nor UO_1652 (O_1652,N_25881,N_29755);
xor UO_1653 (O_1653,N_26842,N_24317);
nor UO_1654 (O_1654,N_28707,N_29305);
or UO_1655 (O_1655,N_27824,N_27875);
nor UO_1656 (O_1656,N_27966,N_25499);
xor UO_1657 (O_1657,N_25492,N_25637);
and UO_1658 (O_1658,N_26988,N_29026);
or UO_1659 (O_1659,N_25693,N_29723);
nand UO_1660 (O_1660,N_28383,N_26530);
xnor UO_1661 (O_1661,N_25042,N_28814);
and UO_1662 (O_1662,N_28747,N_24951);
xor UO_1663 (O_1663,N_28055,N_26608);
or UO_1664 (O_1664,N_25277,N_28576);
xnor UO_1665 (O_1665,N_26314,N_29307);
or UO_1666 (O_1666,N_26785,N_25526);
nand UO_1667 (O_1667,N_29670,N_24207);
nor UO_1668 (O_1668,N_24038,N_28584);
and UO_1669 (O_1669,N_25556,N_29482);
and UO_1670 (O_1670,N_26690,N_27853);
and UO_1671 (O_1671,N_28963,N_24025);
and UO_1672 (O_1672,N_29840,N_25796);
and UO_1673 (O_1673,N_24079,N_25635);
nand UO_1674 (O_1674,N_27155,N_24359);
or UO_1675 (O_1675,N_27296,N_26569);
nand UO_1676 (O_1676,N_29394,N_24303);
nor UO_1677 (O_1677,N_24123,N_24195);
nand UO_1678 (O_1678,N_25121,N_29516);
nor UO_1679 (O_1679,N_25629,N_28612);
and UO_1680 (O_1680,N_27993,N_28409);
or UO_1681 (O_1681,N_24798,N_25615);
nand UO_1682 (O_1682,N_29271,N_26363);
nand UO_1683 (O_1683,N_28185,N_25052);
or UO_1684 (O_1684,N_27748,N_26459);
nor UO_1685 (O_1685,N_25718,N_29092);
xor UO_1686 (O_1686,N_27549,N_24115);
nor UO_1687 (O_1687,N_28388,N_29158);
and UO_1688 (O_1688,N_29567,N_26584);
and UO_1689 (O_1689,N_25377,N_26879);
and UO_1690 (O_1690,N_25328,N_24707);
nor UO_1691 (O_1691,N_27288,N_25859);
nor UO_1692 (O_1692,N_29895,N_28908);
and UO_1693 (O_1693,N_29041,N_24624);
nand UO_1694 (O_1694,N_28522,N_27806);
or UO_1695 (O_1695,N_29107,N_24631);
nand UO_1696 (O_1696,N_29739,N_29773);
or UO_1697 (O_1697,N_26109,N_25897);
or UO_1698 (O_1698,N_29580,N_26120);
nand UO_1699 (O_1699,N_24981,N_28562);
nor UO_1700 (O_1700,N_25218,N_24296);
nand UO_1701 (O_1701,N_29927,N_26899);
nor UO_1702 (O_1702,N_27488,N_28900);
and UO_1703 (O_1703,N_28592,N_29357);
and UO_1704 (O_1704,N_28355,N_29012);
nand UO_1705 (O_1705,N_24466,N_25628);
xnor UO_1706 (O_1706,N_28493,N_29396);
or UO_1707 (O_1707,N_26542,N_28162);
nand UO_1708 (O_1708,N_26022,N_27518);
xnor UO_1709 (O_1709,N_28111,N_28848);
nor UO_1710 (O_1710,N_26416,N_26242);
and UO_1711 (O_1711,N_25416,N_28419);
xnor UO_1712 (O_1712,N_25769,N_25391);
nand UO_1713 (O_1713,N_25664,N_24302);
or UO_1714 (O_1714,N_26675,N_26635);
nand UO_1715 (O_1715,N_28873,N_28708);
nand UO_1716 (O_1716,N_25417,N_29539);
xor UO_1717 (O_1717,N_29421,N_26298);
nor UO_1718 (O_1718,N_28290,N_24468);
nand UO_1719 (O_1719,N_29280,N_26619);
nor UO_1720 (O_1720,N_24336,N_29125);
nor UO_1721 (O_1721,N_24877,N_28808);
or UO_1722 (O_1722,N_28476,N_28986);
and UO_1723 (O_1723,N_25688,N_27695);
xor UO_1724 (O_1724,N_24739,N_29656);
or UO_1725 (O_1725,N_29782,N_24629);
xnor UO_1726 (O_1726,N_28091,N_27067);
nand UO_1727 (O_1727,N_29588,N_27123);
xnor UO_1728 (O_1728,N_25262,N_28406);
or UO_1729 (O_1729,N_29901,N_24381);
and UO_1730 (O_1730,N_28042,N_27984);
or UO_1731 (O_1731,N_24027,N_28881);
and UO_1732 (O_1732,N_29440,N_25182);
nand UO_1733 (O_1733,N_29415,N_28119);
nor UO_1734 (O_1734,N_27111,N_29737);
or UO_1735 (O_1735,N_26010,N_25902);
nor UO_1736 (O_1736,N_29883,N_28407);
nand UO_1737 (O_1737,N_27142,N_25710);
or UO_1738 (O_1738,N_29021,N_25538);
nand UO_1739 (O_1739,N_28797,N_25289);
nor UO_1740 (O_1740,N_29252,N_28110);
or UO_1741 (O_1741,N_29844,N_29037);
nor UO_1742 (O_1742,N_24152,N_29682);
xor UO_1743 (O_1743,N_25060,N_28768);
nand UO_1744 (O_1744,N_25223,N_26968);
or UO_1745 (O_1745,N_25544,N_27237);
xnor UO_1746 (O_1746,N_29929,N_24225);
or UO_1747 (O_1747,N_28326,N_24892);
and UO_1748 (O_1748,N_26980,N_24625);
or UO_1749 (O_1749,N_27952,N_24894);
and UO_1750 (O_1750,N_25952,N_24213);
and UO_1751 (O_1751,N_29299,N_28202);
nand UO_1752 (O_1752,N_24827,N_25106);
nor UO_1753 (O_1753,N_24823,N_29906);
or UO_1754 (O_1754,N_24826,N_26995);
and UO_1755 (O_1755,N_25373,N_29684);
and UO_1756 (O_1756,N_24184,N_29890);
and UO_1757 (O_1757,N_29824,N_28159);
or UO_1758 (O_1758,N_28416,N_28879);
xor UO_1759 (O_1759,N_27916,N_26093);
xnor UO_1760 (O_1760,N_27018,N_29740);
nand UO_1761 (O_1761,N_25116,N_28535);
or UO_1762 (O_1762,N_28057,N_27639);
nor UO_1763 (O_1763,N_27781,N_28232);
and UO_1764 (O_1764,N_28589,N_27688);
and UO_1765 (O_1765,N_29272,N_27180);
xnor UO_1766 (O_1766,N_29865,N_29403);
xor UO_1767 (O_1767,N_24862,N_29342);
and UO_1768 (O_1768,N_28834,N_26307);
nor UO_1769 (O_1769,N_24368,N_24992);
nand UO_1770 (O_1770,N_24196,N_29386);
and UO_1771 (O_1771,N_24121,N_26739);
or UO_1772 (O_1772,N_28785,N_28853);
xor UO_1773 (O_1773,N_24634,N_27458);
nor UO_1774 (O_1774,N_26220,N_24306);
nand UO_1775 (O_1775,N_26015,N_29189);
and UO_1776 (O_1776,N_25250,N_25559);
nor UO_1777 (O_1777,N_29722,N_27103);
nand UO_1778 (O_1778,N_25463,N_27777);
or UO_1779 (O_1779,N_28716,N_25985);
xnor UO_1780 (O_1780,N_25069,N_29358);
xnor UO_1781 (O_1781,N_28040,N_28173);
xnor UO_1782 (O_1782,N_29161,N_28021);
xor UO_1783 (O_1783,N_27943,N_27240);
nand UO_1784 (O_1784,N_24590,N_24924);
nor UO_1785 (O_1785,N_27353,N_26295);
and UO_1786 (O_1786,N_27370,N_26184);
xnor UO_1787 (O_1787,N_25522,N_26079);
xor UO_1788 (O_1788,N_26838,N_24834);
nand UO_1789 (O_1789,N_25868,N_27473);
nor UO_1790 (O_1790,N_28172,N_29477);
or UO_1791 (O_1791,N_24057,N_25055);
xnor UO_1792 (O_1792,N_28541,N_24721);
nand UO_1793 (O_1793,N_29063,N_27228);
nand UO_1794 (O_1794,N_29829,N_27963);
and UO_1795 (O_1795,N_26286,N_28598);
xnor UO_1796 (O_1796,N_28610,N_26288);
nor UO_1797 (O_1797,N_24791,N_24946);
nand UO_1798 (O_1798,N_26073,N_24166);
nor UO_1799 (O_1799,N_25996,N_25975);
xnor UO_1800 (O_1800,N_28967,N_25679);
nor UO_1801 (O_1801,N_26600,N_25101);
and UO_1802 (O_1802,N_24509,N_25765);
xnor UO_1803 (O_1803,N_26662,N_27801);
nand UO_1804 (O_1804,N_26650,N_26197);
nor UO_1805 (O_1805,N_27115,N_28869);
nand UO_1806 (O_1806,N_27323,N_26699);
or UO_1807 (O_1807,N_25254,N_24392);
nor UO_1808 (O_1808,N_25270,N_25462);
or UO_1809 (O_1809,N_26506,N_25882);
or UO_1810 (O_1810,N_28393,N_25366);
nor UO_1811 (O_1811,N_29160,N_28897);
nand UO_1812 (O_1812,N_24248,N_27392);
nor UO_1813 (O_1813,N_25606,N_27949);
nand UO_1814 (O_1814,N_25132,N_29643);
and UO_1815 (O_1815,N_27354,N_28815);
or UO_1816 (O_1816,N_25577,N_28694);
or UO_1817 (O_1817,N_25310,N_26399);
or UO_1818 (O_1818,N_25406,N_25108);
or UO_1819 (O_1819,N_29752,N_28337);
nand UO_1820 (O_1820,N_27084,N_25309);
or UO_1821 (O_1821,N_24076,N_24857);
and UO_1822 (O_1822,N_25542,N_25241);
and UO_1823 (O_1823,N_25774,N_27550);
nor UO_1824 (O_1824,N_27009,N_25523);
nand UO_1825 (O_1825,N_28431,N_25422);
or UO_1826 (O_1826,N_26110,N_26246);
nor UO_1827 (O_1827,N_26161,N_25712);
nor UO_1828 (O_1828,N_27664,N_28489);
nor UO_1829 (O_1829,N_27784,N_28764);
or UO_1830 (O_1830,N_26511,N_28725);
and UO_1831 (O_1831,N_28481,N_28127);
xor UO_1832 (O_1832,N_26046,N_26901);
xor UO_1833 (O_1833,N_24230,N_28514);
and UO_1834 (O_1834,N_26654,N_26027);
or UO_1835 (O_1835,N_27673,N_29899);
xnor UO_1836 (O_1836,N_27355,N_25590);
or UO_1837 (O_1837,N_24497,N_27105);
nand UO_1838 (O_1838,N_26623,N_25224);
nor UO_1839 (O_1839,N_28462,N_27023);
and UO_1840 (O_1840,N_24400,N_28979);
and UO_1841 (O_1841,N_27572,N_24870);
and UO_1842 (O_1842,N_29702,N_29965);
or UO_1843 (O_1843,N_24960,N_27760);
or UO_1844 (O_1844,N_25228,N_27807);
nor UO_1845 (O_1845,N_26035,N_29708);
nand UO_1846 (O_1846,N_24276,N_29451);
or UO_1847 (O_1847,N_28118,N_26948);
nor UO_1848 (O_1848,N_27931,N_29326);
nor UO_1849 (O_1849,N_27674,N_29806);
nand UO_1850 (O_1850,N_28475,N_25267);
nand UO_1851 (O_1851,N_24024,N_26260);
and UO_1852 (O_1852,N_29693,N_26938);
nand UO_1853 (O_1853,N_29324,N_26888);
and UO_1854 (O_1854,N_26794,N_29254);
nor UO_1855 (O_1855,N_27238,N_25336);
or UO_1856 (O_1856,N_26823,N_28524);
and UO_1857 (O_1857,N_29490,N_24256);
nand UO_1858 (O_1858,N_29712,N_24635);
or UO_1859 (O_1859,N_27603,N_28236);
and UO_1860 (O_1860,N_27703,N_27613);
xor UO_1861 (O_1861,N_24020,N_26624);
nor UO_1862 (O_1862,N_24950,N_29766);
nor UO_1863 (O_1863,N_26806,N_27528);
or UO_1864 (O_1864,N_27236,N_25486);
nand UO_1865 (O_1865,N_28210,N_29502);
xnor UO_1866 (O_1866,N_26430,N_28053);
or UO_1867 (O_1867,N_26673,N_28955);
xor UO_1868 (O_1868,N_28860,N_25128);
nor UO_1869 (O_1869,N_27266,N_26698);
xor UO_1870 (O_1870,N_27336,N_29417);
nor UO_1871 (O_1871,N_25832,N_25524);
and UO_1872 (O_1872,N_24613,N_29018);
and UO_1873 (O_1873,N_29589,N_24340);
or UO_1874 (O_1874,N_27808,N_26193);
and UO_1875 (O_1875,N_27959,N_27525);
xor UO_1876 (O_1876,N_29348,N_25689);
nor UO_1877 (O_1877,N_25759,N_25073);
or UO_1878 (O_1878,N_26115,N_25479);
or UO_1879 (O_1879,N_26016,N_28516);
nor UO_1880 (O_1880,N_27800,N_27512);
or UO_1881 (O_1881,N_24893,N_27545);
and UO_1882 (O_1882,N_28933,N_24202);
or UO_1883 (O_1883,N_29633,N_28916);
nand UO_1884 (O_1884,N_28880,N_24448);
xnor UO_1885 (O_1885,N_24957,N_24504);
nor UO_1886 (O_1886,N_26332,N_26723);
and UO_1887 (O_1887,N_26055,N_28767);
and UO_1888 (O_1888,N_25597,N_28927);
nand UO_1889 (O_1889,N_26720,N_27209);
xor UO_1890 (O_1890,N_28148,N_25067);
and UO_1891 (O_1891,N_29556,N_25374);
or UO_1892 (O_1892,N_24973,N_29743);
nor UO_1893 (O_1893,N_24755,N_26144);
xnor UO_1894 (O_1894,N_28184,N_27065);
nor UO_1895 (O_1895,N_25234,N_24053);
xor UO_1896 (O_1896,N_27380,N_26299);
or UO_1897 (O_1897,N_24895,N_24673);
or UO_1898 (O_1898,N_24206,N_28085);
and UO_1899 (O_1899,N_26470,N_29116);
xnor UO_1900 (O_1900,N_26800,N_26827);
or UO_1901 (O_1901,N_29163,N_29481);
nand UO_1902 (O_1902,N_29594,N_28851);
nor UO_1903 (O_1903,N_25161,N_25217);
nor UO_1904 (O_1904,N_26450,N_24062);
xor UO_1905 (O_1905,N_25866,N_27941);
nand UO_1906 (O_1906,N_29631,N_27559);
xor UO_1907 (O_1907,N_25776,N_29174);
xnor UO_1908 (O_1908,N_26890,N_29958);
or UO_1909 (O_1909,N_27460,N_24518);
and UO_1910 (O_1910,N_25160,N_29103);
xnor UO_1911 (O_1911,N_26417,N_27318);
nor UO_1912 (O_1912,N_29309,N_28934);
nand UO_1913 (O_1913,N_28197,N_24561);
and UO_1914 (O_1914,N_26471,N_29783);
and UO_1915 (O_1915,N_27985,N_29465);
and UO_1916 (O_1916,N_28738,N_24486);
or UO_1917 (O_1917,N_27513,N_29961);
nor UO_1918 (O_1918,N_24484,N_27889);
or UO_1919 (O_1919,N_26982,N_25149);
nor UO_1920 (O_1920,N_25977,N_24412);
and UO_1921 (O_1921,N_25081,N_29626);
nor UO_1922 (O_1922,N_28903,N_25815);
and UO_1923 (O_1923,N_27434,N_29409);
nor UO_1924 (O_1924,N_29410,N_27042);
nand UO_1925 (O_1925,N_25220,N_24697);
and UO_1926 (O_1926,N_28007,N_26543);
and UO_1927 (O_1927,N_28001,N_27679);
or UO_1928 (O_1928,N_24727,N_29582);
nor UO_1929 (O_1929,N_26128,N_29289);
and UO_1930 (O_1930,N_25072,N_25922);
nand UO_1931 (O_1931,N_26302,N_28642);
nand UO_1932 (O_1932,N_24234,N_24190);
or UO_1933 (O_1933,N_28998,N_24134);
nor UO_1934 (O_1934,N_26517,N_29435);
and UO_1935 (O_1935,N_26153,N_28616);
xnor UO_1936 (O_1936,N_24718,N_28950);
or UO_1937 (O_1937,N_25243,N_29356);
xor UO_1938 (O_1938,N_27759,N_26292);
or UO_1939 (O_1939,N_27972,N_24843);
and UO_1940 (O_1940,N_29134,N_24188);
xnor UO_1941 (O_1941,N_24934,N_29969);
nor UO_1942 (O_1942,N_26301,N_27563);
or UO_1943 (O_1943,N_27494,N_27723);
or UO_1944 (O_1944,N_28639,N_26492);
xor UO_1945 (O_1945,N_24896,N_28128);
nor UO_1946 (O_1946,N_25757,N_28980);
or UO_1947 (O_1947,N_24440,N_24125);
xor UO_1948 (O_1948,N_28201,N_29897);
or UO_1949 (O_1949,N_24712,N_25566);
xor UO_1950 (O_1950,N_25194,N_24609);
nor UO_1951 (O_1951,N_24627,N_26550);
xnor UO_1952 (O_1952,N_26881,N_29931);
and UO_1953 (O_1953,N_27697,N_28552);
nor UO_1954 (O_1954,N_27629,N_29668);
nand UO_1955 (O_1955,N_25905,N_25588);
nand UO_1956 (O_1956,N_29029,N_25489);
nor UO_1957 (O_1957,N_26579,N_28437);
nand UO_1958 (O_1958,N_28155,N_28918);
xor UO_1959 (O_1959,N_28256,N_26781);
and UO_1960 (O_1960,N_28077,N_26370);
nor UO_1961 (O_1961,N_28117,N_27509);
and UO_1962 (O_1962,N_28217,N_27651);
nor UO_1963 (O_1963,N_24832,N_26731);
and UO_1964 (O_1964,N_27245,N_24446);
nand UO_1965 (O_1965,N_28237,N_27490);
xnor UO_1966 (O_1966,N_24251,N_28421);
or UO_1967 (O_1967,N_26926,N_26287);
nand UO_1968 (O_1968,N_28385,N_24434);
nor UO_1969 (O_1969,N_25155,N_26168);
xnor UO_1970 (O_1970,N_24280,N_27658);
or UO_1971 (O_1971,N_24142,N_25038);
or UO_1972 (O_1972,N_24433,N_28430);
nor UO_1973 (O_1973,N_25989,N_24952);
nand UO_1974 (O_1974,N_26992,N_27456);
nor UO_1975 (O_1975,N_24266,N_29008);
nand UO_1976 (O_1976,N_27422,N_25083);
and UO_1977 (O_1977,N_27728,N_28827);
or UO_1978 (O_1978,N_25177,N_28087);
and UO_1979 (O_1979,N_29603,N_28915);
xnor UO_1980 (O_1980,N_28234,N_27294);
nor UO_1981 (O_1981,N_24008,N_27726);
nor UO_1982 (O_1982,N_26395,N_28137);
xnor UO_1983 (O_1983,N_27623,N_25040);
or UO_1984 (O_1984,N_24404,N_27870);
nand UO_1985 (O_1985,N_27879,N_27397);
nand UO_1986 (O_1986,N_29981,N_29217);
or UO_1987 (O_1987,N_29381,N_25792);
xnor UO_1988 (O_1988,N_27787,N_27657);
and UO_1989 (O_1989,N_25113,N_26198);
xnor UO_1990 (O_1990,N_29155,N_27950);
xor UO_1991 (O_1991,N_29907,N_24899);
or UO_1992 (O_1992,N_26671,N_28338);
nor UO_1993 (O_1993,N_29625,N_24463);
nor UO_1994 (O_1994,N_29793,N_29019);
or UO_1995 (O_1995,N_24235,N_28543);
nor UO_1996 (O_1996,N_28818,N_26520);
or UO_1997 (O_1997,N_27369,N_28024);
nor UO_1998 (O_1998,N_28105,N_25457);
nand UO_1999 (O_1999,N_28395,N_28168);
and UO_2000 (O_2000,N_27125,N_25426);
nor UO_2001 (O_2001,N_27130,N_25205);
and UO_2002 (O_2002,N_26647,N_28839);
nor UO_2003 (O_2003,N_24372,N_25404);
nor UO_2004 (O_2004,N_26219,N_27968);
xor UO_2005 (O_2005,N_27856,N_26482);
nand UO_2006 (O_2006,N_28760,N_27692);
or UO_2007 (O_2007,N_27010,N_26175);
or UO_2008 (O_2008,N_29014,N_28756);
and UO_2009 (O_2009,N_28877,N_28898);
xnor UO_2010 (O_2010,N_25443,N_26746);
nand UO_2011 (O_2011,N_29860,N_24849);
or UO_2012 (O_2012,N_26449,N_24122);
nor UO_2013 (O_2013,N_25784,N_25880);
and UO_2014 (O_2014,N_24852,N_27399);
or UO_2015 (O_2015,N_25589,N_29930);
or UO_2016 (O_2016,N_27751,N_25714);
xnor UO_2017 (O_2017,N_27710,N_28746);
or UO_2018 (O_2018,N_27048,N_25274);
xor UO_2019 (O_2019,N_25980,N_29593);
nand UO_2020 (O_2020,N_29276,N_27484);
or UO_2021 (O_2021,N_24962,N_29438);
xor UO_2022 (O_2022,N_24789,N_27852);
or UO_2023 (O_2023,N_26483,N_27878);
or UO_2024 (O_2024,N_25535,N_25598);
nor UO_2025 (O_2025,N_26527,N_27936);
nor UO_2026 (O_2026,N_27116,N_29152);
nand UO_2027 (O_2027,N_25587,N_24515);
and UO_2028 (O_2028,N_25527,N_26790);
or UO_2029 (O_2029,N_28377,N_28647);
and UO_2030 (O_2030,N_26886,N_28479);
nand UO_2031 (O_2031,N_25509,N_29825);
nor UO_2032 (O_2032,N_29172,N_24780);
and UO_2033 (O_2033,N_27202,N_29393);
and UO_2034 (O_2034,N_28192,N_27198);
nor UO_2035 (O_2035,N_29794,N_25869);
nor UO_2036 (O_2036,N_27529,N_27377);
nand UO_2037 (O_2037,N_29127,N_27019);
nor UO_2038 (O_2038,N_28332,N_27999);
nand UO_2039 (O_2039,N_25787,N_27012);
and UO_2040 (O_2040,N_29982,N_27283);
nand UO_2041 (O_2041,N_28961,N_29201);
xnor UO_2042 (O_2042,N_29648,N_28997);
nor UO_2043 (O_2043,N_24232,N_29040);
and UO_2044 (O_2044,N_25292,N_26687);
xor UO_2045 (O_2045,N_24584,N_28724);
xor UO_2046 (O_2046,N_26983,N_25117);
nand UO_2047 (O_2047,N_27057,N_26973);
nand UO_2048 (O_2048,N_26402,N_29759);
nand UO_2049 (O_2049,N_27339,N_25322);
nand UO_2050 (O_2050,N_29137,N_24848);
or UO_2051 (O_2051,N_28525,N_28441);
and UO_2052 (O_2052,N_28227,N_24781);
nand UO_2053 (O_2053,N_29208,N_26727);
nand UO_2054 (O_2054,N_24532,N_28260);
nor UO_2055 (O_2055,N_24854,N_28864);
nand UO_2056 (O_2056,N_28212,N_28183);
xnor UO_2057 (O_2057,N_28775,N_27987);
or UO_2058 (O_2058,N_26293,N_26059);
nand UO_2059 (O_2059,N_24105,N_25349);
xor UO_2060 (O_2060,N_28886,N_25665);
nor UO_2061 (O_2061,N_24604,N_26213);
and UO_2062 (O_2062,N_28369,N_28447);
and UO_2063 (O_2063,N_25534,N_27320);
and UO_2064 (O_2064,N_24666,N_27938);
and UO_2065 (O_2065,N_27526,N_27134);
and UO_2066 (O_2066,N_24041,N_29655);
nor UO_2067 (O_2067,N_25392,N_29685);
or UO_2068 (O_2068,N_29709,N_24653);
nor UO_2069 (O_2069,N_26390,N_26552);
xnor UO_2070 (O_2070,N_29562,N_29153);
and UO_2071 (O_2071,N_27925,N_28084);
or UO_2072 (O_2072,N_28857,N_26819);
nand UO_2073 (O_2073,N_26668,N_29085);
nor UO_2074 (O_2074,N_25251,N_24503);
and UO_2075 (O_2075,N_24589,N_26145);
nor UO_2076 (O_2076,N_29942,N_28004);
nor UO_2077 (O_2077,N_29529,N_25095);
and UO_2078 (O_2078,N_24913,N_26255);
nand UO_2079 (O_2079,N_27285,N_29530);
xor UO_2080 (O_2080,N_27895,N_29300);
nand UO_2081 (O_2081,N_27827,N_24268);
and UO_2082 (O_2082,N_26174,N_25713);
nand UO_2083 (O_2083,N_28740,N_29991);
nand UO_2084 (O_2084,N_24212,N_29045);
or UO_2085 (O_2085,N_25525,N_25932);
or UO_2086 (O_2086,N_29186,N_25640);
nand UO_2087 (O_2087,N_27859,N_25271);
and UO_2088 (O_2088,N_25861,N_25670);
nand UO_2089 (O_2089,N_25560,N_25578);
nor UO_2090 (O_2090,N_26074,N_26341);
or UO_2091 (O_2091,N_27593,N_27996);
xor UO_2092 (O_2092,N_29994,N_29653);
or UO_2093 (O_2093,N_28960,N_24921);
nor UO_2094 (O_2094,N_25491,N_27735);
or UO_2095 (O_2095,N_28803,N_29350);
and UO_2096 (O_2096,N_25458,N_28089);
nor UO_2097 (O_2097,N_27061,N_29343);
nor UO_2098 (O_2098,N_28083,N_28457);
xnor UO_2099 (O_2099,N_28904,N_26315);
xnor UO_2100 (O_2100,N_28791,N_27753);
xor UO_2101 (O_2101,N_25456,N_25129);
and UO_2102 (O_2102,N_26965,N_29946);
or UO_2103 (O_2103,N_27006,N_24864);
and UO_2104 (O_2104,N_26904,N_29807);
nor UO_2105 (O_2105,N_28310,N_29887);
nor UO_2106 (O_2106,N_26157,N_25233);
nor UO_2107 (O_2107,N_27803,N_25812);
and UO_2108 (O_2108,N_27420,N_28180);
or UO_2109 (O_2109,N_28151,N_26791);
or UO_2110 (O_2110,N_25097,N_26189);
or UO_2111 (O_2111,N_28323,N_27967);
nand UO_2112 (O_2112,N_24669,N_28343);
or UO_2113 (O_2113,N_26908,N_24292);
xnor UO_2114 (O_2114,N_27026,N_28828);
or UO_2115 (O_2115,N_28011,N_24006);
nor UO_2116 (O_2116,N_24916,N_28556);
nor UO_2117 (O_2117,N_24015,N_24472);
or UO_2118 (O_2118,N_25370,N_24244);
nand UO_2119 (O_2119,N_28138,N_24352);
nand UO_2120 (O_2120,N_27742,N_28807);
nand UO_2121 (O_2121,N_29139,N_25286);
nand UO_2122 (O_2122,N_25511,N_29613);
nand UO_2123 (O_2123,N_27252,N_24272);
or UO_2124 (O_2124,N_24674,N_26262);
or UO_2125 (O_2125,N_29869,N_29177);
or UO_2126 (O_2126,N_25844,N_28951);
and UO_2127 (O_2127,N_29695,N_26071);
nand UO_2128 (O_2128,N_26333,N_27554);
xor UO_2129 (O_2129,N_26434,N_28468);
xor UO_2130 (O_2130,N_26141,N_29390);
nor UO_2131 (O_2131,N_26555,N_27372);
nand UO_2132 (O_2132,N_28906,N_27087);
nor UO_2133 (O_2133,N_25378,N_26391);
and UO_2134 (O_2134,N_28048,N_29111);
or UO_2135 (O_2135,N_27143,N_28020);
or UO_2136 (O_2136,N_25991,N_27179);
nor UO_2137 (O_2137,N_24242,N_24476);
xor UO_2138 (O_2138,N_25503,N_25800);
xor UO_2139 (O_2139,N_27552,N_27183);
nor UO_2140 (O_2140,N_27279,N_25303);
nand UO_2141 (O_2141,N_29119,N_28056);
or UO_2142 (O_2142,N_29000,N_28428);
or UO_2143 (O_2143,N_28947,N_26917);
nor UO_2144 (O_2144,N_29561,N_24907);
and UO_2145 (O_2145,N_27793,N_25953);
xnor UO_2146 (O_2146,N_25163,N_29038);
xor UO_2147 (O_2147,N_26421,N_28591);
or UO_2148 (O_2148,N_28292,N_25833);
xnor UO_2149 (O_2149,N_25180,N_24454);
xnor UO_2150 (O_2150,N_25353,N_24360);
xor UO_2151 (O_2151,N_25835,N_26933);
xnor UO_2152 (O_2152,N_25703,N_29885);
and UO_2153 (O_2153,N_29022,N_28471);
xnor UO_2154 (O_2154,N_26004,N_26294);
nor UO_2155 (O_2155,N_25910,N_25546);
xor UO_2156 (O_2156,N_24665,N_24492);
nor UO_2157 (O_2157,N_26234,N_26281);
nor UO_2158 (O_2158,N_29786,N_29166);
and UO_2159 (O_2159,N_26947,N_24397);
or UO_2160 (O_2160,N_27376,N_24757);
nand UO_2161 (O_2161,N_26809,N_25634);
and UO_2162 (O_2162,N_26769,N_27455);
or UO_2163 (O_2163,N_29443,N_26211);
or UO_2164 (O_2164,N_25014,N_27672);
or UO_2165 (O_2165,N_24991,N_24708);
xor UO_2166 (O_2166,N_27833,N_28226);
and UO_2167 (O_2167,N_25301,N_26580);
and UO_2168 (O_2168,N_27229,N_29564);
nand UO_2169 (O_2169,N_26729,N_27791);
and UO_2170 (O_2170,N_25122,N_28046);
or UO_2171 (O_2171,N_24104,N_27541);
and UO_2172 (O_2172,N_28308,N_24036);
nor UO_2173 (O_2173,N_25497,N_28497);
xnor UO_2174 (O_2174,N_28280,N_24069);
and UO_2175 (O_2175,N_24732,N_29808);
xor UO_2176 (O_2176,N_27502,N_28152);
nand UO_2177 (O_2177,N_26944,N_28160);
and UO_2178 (O_2178,N_24573,N_26831);
nand UO_2179 (O_2179,N_25809,N_26518);
or UO_2180 (O_2180,N_27973,N_27721);
xnor UO_2181 (O_2181,N_25614,N_25169);
and UO_2182 (O_2182,N_29911,N_28342);
or UO_2183 (O_2183,N_24246,N_28845);
and UO_2184 (O_2184,N_28527,N_27464);
and UO_2185 (O_2185,N_27479,N_25873);
nor UO_2186 (O_2186,N_29074,N_28328);
nand UO_2187 (O_2187,N_28275,N_25403);
nand UO_2188 (O_2188,N_24796,N_28302);
xor UO_2189 (O_2189,N_24411,N_28512);
xor UO_2190 (O_2190,N_25874,N_25295);
and UO_2191 (O_2191,N_28607,N_28282);
and UO_2192 (O_2192,N_26488,N_28769);
xor UO_2193 (O_2193,N_29099,N_24556);
nor UO_2194 (O_2194,N_29933,N_27821);
nor UO_2195 (O_2195,N_29792,N_28777);
or UO_2196 (O_2196,N_26049,N_27669);
and UO_2197 (O_2197,N_24999,N_24557);
nor UO_2198 (O_2198,N_27739,N_24300);
xor UO_2199 (O_2199,N_29077,N_26040);
and UO_2200 (O_2200,N_24338,N_29234);
nor UO_2201 (O_2201,N_29242,N_28329);
and UO_2202 (O_2202,N_24595,N_26258);
nor UO_2203 (O_2203,N_28792,N_27480);
xor UO_2204 (O_2204,N_27928,N_26631);
or UO_2205 (O_2205,N_26868,N_29433);
nand UO_2206 (O_2206,N_29055,N_25092);
xnor UO_2207 (O_2207,N_29964,N_24764);
nand UO_2208 (O_2208,N_27818,N_29048);
nand UO_2209 (O_2209,N_27638,N_24129);
and UO_2210 (O_2210,N_29635,N_24491);
or UO_2211 (O_2211,N_26801,N_27752);
or UO_2212 (O_2212,N_28833,N_28609);
nand UO_2213 (O_2213,N_29788,N_26371);
and UO_2214 (O_2214,N_24178,N_24021);
or UO_2215 (O_2215,N_25976,N_25580);
nor UO_2216 (O_2216,N_27558,N_27423);
or UO_2217 (O_2217,N_29027,N_25921);
nand UO_2218 (O_2218,N_26750,N_29196);
nand UO_2219 (O_2219,N_25178,N_26204);
xor UO_2220 (O_2220,N_27997,N_24345);
nor UO_2221 (O_2221,N_29133,N_27717);
nand UO_2222 (O_2222,N_28924,N_26865);
nor UO_2223 (O_2223,N_27260,N_26188);
nand UO_2224 (O_2224,N_29607,N_29260);
xor UO_2225 (O_2225,N_29934,N_27346);
nor UO_2226 (O_2226,N_27005,N_29716);
nor UO_2227 (O_2227,N_28685,N_26068);
nand UO_2228 (O_2228,N_24286,N_27124);
xor UO_2229 (O_2229,N_25402,N_26979);
nor UO_2230 (O_2230,N_25695,N_26845);
nand UO_2231 (O_2231,N_27750,N_27412);
and UO_2232 (O_2232,N_24136,N_25811);
nor UO_2233 (O_2233,N_28472,N_25091);
nand UO_2234 (O_2234,N_26691,N_28196);
nor UO_2235 (O_2235,N_29235,N_27239);
or UO_2236 (O_2236,N_24722,N_29976);
and UO_2237 (O_2237,N_26385,N_28316);
nor UO_2238 (O_2238,N_26311,N_24744);
or UO_2239 (O_2239,N_24879,N_29506);
or UO_2240 (O_2240,N_25979,N_27011);
or UO_2241 (O_2241,N_24672,N_26892);
or UO_2242 (O_2242,N_26551,N_25501);
and UO_2243 (O_2243,N_24221,N_29308);
xor UO_2244 (O_2244,N_24583,N_28703);
nand UO_2245 (O_2245,N_25337,N_28910);
xor UO_2246 (O_2246,N_28644,N_28229);
xor UO_2247 (O_2247,N_26377,N_25642);
nor UO_2248 (O_2248,N_28378,N_28956);
nand UO_2249 (O_2249,N_25425,N_24427);
nand UO_2250 (O_2250,N_24154,N_24651);
or UO_2251 (O_2251,N_24257,N_29765);
nand UO_2252 (O_2252,N_29932,N_29398);
xnor UO_2253 (O_2253,N_24657,N_24353);
xor UO_2254 (O_2254,N_25298,N_26774);
and UO_2255 (O_2255,N_27398,N_24164);
or UO_2256 (O_2256,N_25667,N_28572);
or UO_2257 (O_2257,N_29761,N_28353);
or UO_2258 (O_2258,N_27850,N_26510);
and UO_2259 (O_2259,N_26514,N_25994);
or UO_2260 (O_2260,N_24693,N_25280);
xor UO_2261 (O_2261,N_29941,N_29614);
nor UO_2262 (O_2262,N_24471,N_28866);
nor UO_2263 (O_2263,N_25838,N_29721);
nor UO_2264 (O_2264,N_26020,N_29388);
nand UO_2265 (O_2265,N_27774,N_24704);
or UO_2266 (O_2266,N_27390,N_24873);
or UO_2267 (O_2267,N_24539,N_25485);
nand UO_2268 (O_2268,N_26793,N_28109);
and UO_2269 (O_2269,N_25037,N_24833);
xor UO_2270 (O_2270,N_26374,N_26495);
or UO_2271 (O_2271,N_28186,N_24889);
and UO_2272 (O_2272,N_29538,N_24847);
and UO_2273 (O_2273,N_26454,N_28670);
nor UO_2274 (O_2274,N_28330,N_28484);
nand UO_2275 (O_2275,N_26505,N_28134);
xnor UO_2276 (O_2276,N_24863,N_24398);
and UO_2277 (O_2277,N_24009,N_27649);
xor UO_2278 (O_2278,N_24714,N_28384);
nand UO_2279 (O_2279,N_25845,N_27589);
and UO_2280 (O_2280,N_27520,N_28978);
nor UO_2281 (O_2281,N_24701,N_27457);
or UO_2282 (O_2282,N_26230,N_28285);
nand UO_2283 (O_2283,N_24536,N_29918);
xnor UO_2284 (O_2284,N_24373,N_27660);
nor UO_2285 (O_2285,N_27880,N_29306);
nand UO_2286 (O_2286,N_27328,N_28813);
and UO_2287 (O_2287,N_25857,N_26814);
and UO_2288 (O_2288,N_24554,N_24394);
and UO_2289 (O_2289,N_24618,N_27247);
or UO_2290 (O_2290,N_27665,N_27001);
or UO_2291 (O_2291,N_29615,N_24451);
xnor UO_2292 (O_2292,N_29426,N_25510);
nor UO_2293 (O_2293,N_24082,N_26232);
nor UO_2294 (O_2294,N_29909,N_29736);
xor UO_2295 (O_2295,N_28209,N_28691);
xnor UO_2296 (O_2296,N_25039,N_25697);
nor UO_2297 (O_2297,N_25894,N_26058);
or UO_2298 (O_2298,N_26134,N_25692);
nand UO_2299 (O_2299,N_27652,N_26797);
or UO_2300 (O_2300,N_29475,N_27922);
and UO_2301 (O_2301,N_25638,N_28135);
nand UO_2302 (O_2302,N_26460,N_27095);
and UO_2303 (O_2303,N_24880,N_27431);
xor UO_2304 (O_2304,N_29841,N_29084);
or UO_2305 (O_2305,N_26426,N_27121);
nand UO_2306 (O_2306,N_27960,N_24766);
nand UO_2307 (O_2307,N_29468,N_29638);
nor UO_2308 (O_2308,N_25733,N_29820);
xnor UO_2309 (O_2309,N_26849,N_25775);
nand UO_2310 (O_2310,N_27215,N_24731);
nor UO_2311 (O_2311,N_25053,N_24416);
nor UO_2312 (O_2312,N_25335,N_29319);
nand UO_2313 (O_2313,N_24576,N_27039);
or UO_2314 (O_2314,N_28261,N_25663);
nand UO_2315 (O_2315,N_27902,N_29601);
and UO_2316 (O_2316,N_28460,N_29980);
or UO_2317 (O_2317,N_24420,N_26765);
xor UO_2318 (O_2318,N_29035,N_26617);
xor UO_2319 (O_2319,N_29316,N_29399);
nand UO_2320 (O_2320,N_24282,N_25650);
xnor UO_2321 (O_2321,N_28182,N_28518);
nand UO_2322 (O_2322,N_29261,N_25430);
nor UO_2323 (O_2323,N_27944,N_27537);
and UO_2324 (O_2324,N_24586,N_25332);
nand UO_2325 (O_2325,N_25839,N_25003);
xor UO_2326 (O_2326,N_25033,N_26589);
nor UO_2327 (O_2327,N_28190,N_27631);
nor UO_2328 (O_2328,N_24236,N_29548);
nand UO_2329 (O_2329,N_26602,N_26149);
nor UO_2330 (O_2330,N_28495,N_26372);
xor UO_2331 (O_2331,N_25045,N_25125);
nor UO_2332 (O_2332,N_28165,N_25032);
xnor UO_2333 (O_2333,N_28397,N_26656);
and UO_2334 (O_2334,N_27954,N_26923);
or UO_2335 (O_2335,N_28017,N_25261);
xnor UO_2336 (O_2336,N_29874,N_24662);
nor UO_2337 (O_2337,N_26533,N_28765);
nand UO_2338 (O_2338,N_27483,N_25229);
nand UO_2339 (O_2339,N_28830,N_27411);
or UO_2340 (O_2340,N_26597,N_24170);
nand UO_2341 (O_2341,N_25786,N_25351);
nand UO_2342 (O_2342,N_26821,N_27402);
nor UO_2343 (O_2343,N_26702,N_29450);
nand UO_2344 (O_2344,N_27712,N_25247);
and UO_2345 (O_2345,N_28299,N_26844);
nand UO_2346 (O_2346,N_27881,N_26960);
or UO_2347 (O_2347,N_27014,N_28438);
nor UO_2348 (O_2348,N_26928,N_28611);
nor UO_2349 (O_2349,N_28787,N_26009);
and UO_2350 (O_2350,N_27210,N_26111);
and UO_2351 (O_2351,N_29959,N_27341);
nand UO_2352 (O_2352,N_25753,N_25199);
nand UO_2353 (O_2353,N_27379,N_24443);
xor UO_2354 (O_2354,N_27394,N_29974);
and UO_2355 (O_2355,N_28988,N_24316);
nand UO_2356 (O_2356,N_27362,N_28855);
nor UO_2357 (O_2357,N_25447,N_29314);
and UO_2358 (O_2358,N_26652,N_26366);
nor UO_2359 (O_2359,N_28131,N_24388);
xor UO_2360 (O_2360,N_25517,N_29145);
nand UO_2361 (O_2361,N_24100,N_28995);
or UO_2362 (O_2362,N_29746,N_27876);
xnor UO_2363 (O_2363,N_25450,N_27540);
nor UO_2364 (O_2364,N_24740,N_28453);
xor UO_2365 (O_2365,N_25451,N_29428);
or UO_2366 (O_2366,N_25612,N_29571);
nor UO_2367 (O_2367,N_26824,N_24140);
and UO_2368 (O_2368,N_29692,N_27159);
or UO_2369 (O_2369,N_24482,N_24445);
or UO_2370 (O_2370,N_25929,N_26318);
nand UO_2371 (O_2371,N_29790,N_24689);
nor UO_2372 (O_2372,N_29341,N_29576);
or UO_2373 (O_2373,N_29376,N_25551);
xor UO_2374 (O_2374,N_27953,N_24138);
nand UO_2375 (O_2375,N_29947,N_26817);
nor UO_2376 (O_2376,N_29023,N_29460);
and UO_2377 (O_2377,N_28277,N_27764);
xor UO_2378 (O_2378,N_27160,N_26894);
nand UO_2379 (O_2379,N_28674,N_27640);
and UO_2380 (O_2380,N_29301,N_25173);
xnor UO_2381 (O_2381,N_26054,N_25970);
nand UO_2382 (O_2382,N_24023,N_26642);
nor UO_2383 (O_2383,N_28250,N_25372);
and UO_2384 (O_2384,N_27337,N_26997);
nand UO_2385 (O_2385,N_27097,N_25983);
and UO_2386 (O_2386,N_29339,N_28523);
xor UO_2387 (O_2387,N_29733,N_29566);
nor UO_2388 (O_2388,N_28372,N_24056);
nand UO_2389 (O_2389,N_25591,N_27410);
nand UO_2390 (O_2390,N_29203,N_28653);
nor UO_2391 (O_2391,N_28243,N_29769);
xor UO_2392 (O_2392,N_25698,N_27986);
xnor UO_2393 (O_2393,N_28334,N_29231);
nor UO_2394 (O_2394,N_26548,N_24760);
nor UO_2395 (O_2395,N_25308,N_27691);
nand UO_2396 (O_2396,N_26346,N_24512);
and UO_2397 (O_2397,N_24922,N_24449);
nand UO_2398 (O_2398,N_27282,N_29984);
xor UO_2399 (O_2399,N_28322,N_24035);
nor UO_2400 (O_2400,N_24954,N_25394);
or UO_2401 (O_2401,N_26718,N_26249);
nand UO_2402 (O_2402,N_24177,N_25484);
xor UO_2403 (O_2403,N_24919,N_24470);
or UO_2404 (O_2404,N_27317,N_28002);
nand UO_2405 (O_2405,N_28938,N_29268);
nand UO_2406 (O_2406,N_26436,N_25662);
nand UO_2407 (O_2407,N_25008,N_24495);
nand UO_2408 (O_2408,N_28590,N_24683);
nor UO_2409 (O_2409,N_24013,N_25015);
and UO_2410 (O_2410,N_24133,N_25342);
and UO_2411 (O_2411,N_25357,N_26632);
nand UO_2412 (O_2412,N_26347,N_27965);
xor UO_2413 (O_2413,N_29707,N_27994);
xnor UO_2414 (O_2414,N_27893,N_25048);
xnor UO_2415 (O_2415,N_26351,N_25343);
nand UO_2416 (O_2416,N_28418,N_27021);
nand UO_2417 (O_2417,N_29331,N_25159);
xor UO_2418 (O_2418,N_28930,N_29627);
nor UO_2419 (O_2419,N_26660,N_25013);
or UO_2420 (O_2420,N_24452,N_26978);
and UO_2421 (O_2421,N_24393,N_24883);
nor UO_2422 (O_2422,N_29978,N_29135);
nor UO_2423 (O_2423,N_25118,N_29854);
nand UO_2424 (O_2424,N_24858,N_27890);
nand UO_2425 (O_2425,N_25102,N_27912);
or UO_2426 (O_2426,N_25602,N_29673);
nor UO_2427 (O_2427,N_29204,N_24850);
xnor UO_2428 (O_2428,N_28811,N_24770);
nor UO_2429 (O_2429,N_26683,N_29082);
nor UO_2430 (O_2430,N_27489,N_25086);
nand UO_2431 (O_2431,N_25278,N_28640);
xor UO_2432 (O_2432,N_26665,N_24307);
or UO_2433 (O_2433,N_24473,N_26735);
nand UO_2434 (O_2434,N_27596,N_26880);
nor UO_2435 (O_2435,N_26343,N_26578);
and UO_2436 (O_2436,N_26766,N_27825);
and UO_2437 (O_2437,N_24968,N_28891);
nand UO_2438 (O_2438,N_26741,N_24488);
nor UO_2439 (O_2439,N_28688,N_25354);
nor UO_2440 (O_2440,N_29898,N_28013);
and UO_2441 (O_2441,N_27309,N_27772);
and UO_2442 (O_2442,N_24566,N_24384);
nand UO_2443 (O_2443,N_26349,N_29463);
or UO_2444 (O_2444,N_28169,N_25783);
or UO_2445 (O_2445,N_29359,N_26375);
or UO_2446 (O_2446,N_25171,N_29671);
and UO_2447 (O_2447,N_24314,N_26906);
and UO_2448 (O_2448,N_25302,N_29924);
and UO_2449 (O_2449,N_26038,N_28387);
or UO_2450 (O_2450,N_26626,N_28529);
nor UO_2451 (O_2451,N_29560,N_26981);
xnor UO_2452 (O_2452,N_28506,N_28896);
or UO_2453 (O_2453,N_29205,N_24524);
or UO_2454 (O_2454,N_25222,N_24522);
xnor UO_2455 (O_2455,N_24365,N_29940);
or UO_2456 (O_2456,N_26986,N_28150);
or UO_2457 (O_2457,N_26327,N_29649);
nand UO_2458 (O_2458,N_29206,N_25586);
or UO_2459 (O_2459,N_27110,N_25647);
or UO_2460 (O_2460,N_28515,N_24157);
or UO_2461 (O_2461,N_27766,N_25867);
nor UO_2462 (O_2462,N_26862,N_24387);
nand UO_2463 (O_2463,N_26744,N_27861);
nor UO_2464 (O_2464,N_26271,N_25407);
or UO_2465 (O_2465,N_28144,N_28697);
and UO_2466 (O_2466,N_27452,N_25657);
or UO_2467 (O_2467,N_27330,N_29273);
nand UO_2468 (O_2468,N_24432,N_28932);
and UO_2469 (O_2469,N_24141,N_24802);
nor UO_2470 (O_2470,N_28677,N_27614);
and UO_2471 (O_2471,N_27758,N_26684);
nand UO_2472 (O_2472,N_28623,N_29644);
and UO_2473 (O_2473,N_24797,N_25621);
or UO_2474 (O_2474,N_27426,N_24214);
xnor UO_2475 (O_2475,N_28794,N_28370);
and UO_2476 (O_2476,N_29595,N_29666);
nor UO_2477 (O_2477,N_24965,N_26208);
xnor UO_2478 (O_2478,N_25954,N_24558);
nor UO_2479 (O_2479,N_29191,N_29745);
and UO_2480 (O_2480,N_27016,N_25513);
or UO_2481 (O_2481,N_26646,N_29287);
xnor UO_2482 (O_2482,N_26946,N_26205);
xor UO_2483 (O_2483,N_29060,N_24217);
or UO_2484 (O_2484,N_25891,N_26335);
and UO_2485 (O_2485,N_24005,N_27605);
or UO_2486 (O_2486,N_25917,N_26571);
or UO_2487 (O_2487,N_29513,N_27446);
nand UO_2488 (O_2488,N_28062,N_25387);
nand UO_2489 (O_2489,N_29600,N_26830);
and UO_2490 (O_2490,N_28401,N_27190);
or UO_2491 (O_2491,N_24479,N_25570);
or UO_2492 (O_2492,N_29552,N_29632);
or UO_2493 (O_2493,N_25195,N_25109);
xor UO_2494 (O_2494,N_28033,N_29522);
or UO_2495 (O_2495,N_25293,N_29293);
and UO_2496 (O_2496,N_29679,N_27395);
or UO_2497 (O_2497,N_29449,N_28743);
nand UO_2498 (O_2498,N_29269,N_29620);
and UO_2499 (O_2499,N_26389,N_29384);
nand UO_2500 (O_2500,N_25660,N_27517);
nor UO_2501 (O_2501,N_25683,N_26852);
nand UO_2502 (O_2502,N_26364,N_24945);
xor UO_2503 (O_2503,N_28817,N_28964);
and UO_2504 (O_2504,N_29557,N_24081);
and UO_2505 (O_2505,N_28045,N_28805);
nor UO_2506 (O_2506,N_27835,N_29775);
and UO_2507 (O_2507,N_27345,N_24840);
nand UO_2508 (O_2508,N_24435,N_24717);
and UO_2509 (O_2509,N_25685,N_26398);
xor UO_2510 (O_2510,N_28728,N_24019);
and UO_2511 (O_2511,N_26836,N_24231);
and UO_2512 (O_2512,N_26523,N_24882);
or UO_2513 (O_2513,N_27675,N_27899);
or UO_2514 (O_2514,N_24687,N_25814);
nand UO_2515 (O_2515,N_28116,N_27444);
nand UO_2516 (O_2516,N_24204,N_26825);
and UO_2517 (O_2517,N_27273,N_25437);
nand UO_2518 (O_2518,N_26939,N_29687);
nand UO_2519 (O_2519,N_24529,N_26386);
xor UO_2520 (O_2520,N_25240,N_29043);
and UO_2521 (O_2521,N_28566,N_26033);
nand UO_2522 (O_2522,N_26837,N_25842);
or UO_2523 (O_2523,N_25381,N_26275);
nand UO_2524 (O_2524,N_25400,N_24071);
xnor UO_2525 (O_2525,N_27425,N_29979);
and UO_2526 (O_2526,N_27271,N_25124);
xnor UO_2527 (O_2527,N_25043,N_29738);
nor UO_2528 (O_2528,N_25855,N_26914);
nand UO_2529 (O_2529,N_25200,N_24287);
or UO_2530 (O_2530,N_29297,N_26893);
xor UO_2531 (O_2531,N_27863,N_26309);
nor UO_2532 (O_2532,N_27686,N_28360);
nor UO_2533 (O_2533,N_26661,N_26223);
or UO_2534 (O_2534,N_26931,N_27141);
or UO_2535 (O_2535,N_26431,N_27437);
nand UO_2536 (O_2536,N_25356,N_27487);
nand UO_2537 (O_2537,N_25852,N_25915);
nand UO_2538 (O_2538,N_27567,N_24761);
nor UO_2539 (O_2539,N_26672,N_26712);
xnor UO_2540 (O_2540,N_27366,N_27740);
nand UO_2541 (O_2541,N_27333,N_27867);
xnor UO_2542 (O_2542,N_24305,N_24548);
or UO_2543 (O_2543,N_24851,N_25410);
nor UO_2544 (O_2544,N_24290,N_28067);
and UO_2545 (O_2545,N_24641,N_24250);
nand UO_2546 (O_2546,N_27523,N_24128);
or UO_2547 (O_2547,N_29146,N_24596);
nand UO_2548 (O_2548,N_25627,N_27313);
nand UO_2549 (O_2549,N_26595,N_28120);
and UO_2550 (O_2550,N_25078,N_25595);
nor UO_2551 (O_2551,N_25266,N_29756);
and UO_2552 (O_2552,N_24059,N_29936);
nor UO_2553 (O_2553,N_29001,N_29071);
nand UO_2554 (O_2554,N_28368,N_24737);
or UO_2555 (O_2555,N_29662,N_27290);
nand UO_2556 (O_2556,N_25810,N_24363);
nand UO_2557 (O_2557,N_28858,N_24966);
xor UO_2558 (O_2558,N_24179,N_26850);
and UO_2559 (O_2559,N_25379,N_25592);
or UO_2560 (O_2560,N_29183,N_24795);
or UO_2561 (O_2561,N_25737,N_29185);
nand UO_2562 (O_2562,N_25987,N_29813);
or UO_2563 (O_2563,N_29520,N_26604);
or UO_2564 (O_2564,N_26728,N_24828);
nor UO_2565 (O_2565,N_28297,N_28875);
or UO_2566 (O_2566,N_28076,N_24774);
nor UO_2567 (O_2567,N_29891,N_29672);
or UO_2568 (O_2568,N_24853,N_27830);
nand UO_2569 (O_2569,N_25565,N_27416);
or UO_2570 (O_2570,N_24113,N_26044);
or UO_2571 (O_2571,N_26953,N_29003);
or UO_2572 (O_2572,N_27078,N_24906);
nand UO_2573 (O_2573,N_25936,N_27884);
xnor UO_2574 (O_2574,N_24941,N_26920);
or UO_2575 (O_2575,N_28996,N_29207);
xor UO_2576 (O_2576,N_25829,N_29999);
xor UO_2577 (O_2577,N_28115,N_25957);
or UO_2578 (O_2578,N_25239,N_26192);
xor UO_2579 (O_2579,N_24982,N_26976);
nor UO_2580 (O_2580,N_27312,N_27659);
xnor UO_2581 (O_2581,N_26951,N_29938);
nand UO_2582 (O_2582,N_28958,N_28942);
or UO_2583 (O_2583,N_29903,N_28059);
or UO_2584 (O_2584,N_28487,N_27733);
xor UO_2585 (O_2585,N_27319,N_29444);
nand UO_2586 (O_2586,N_25594,N_29407);
nor UO_2587 (O_2587,N_27849,N_24995);
nand UO_2588 (O_2588,N_27812,N_29178);
xor UO_2589 (O_2589,N_24531,N_25895);
nand UO_2590 (O_2590,N_24702,N_24824);
nor UO_2591 (O_2591,N_26440,N_26082);
xnor UO_2592 (O_2592,N_27573,N_26400);
nor UO_2593 (O_2593,N_25181,N_26977);
nand UO_2594 (O_2594,N_24377,N_26710);
or UO_2595 (O_2595,N_28218,N_28913);
and UO_2596 (O_2596,N_28663,N_24918);
or UO_2597 (O_2597,N_24172,N_24459);
xor UO_2598 (O_2598,N_26325,N_24839);
nand UO_2599 (O_2599,N_27326,N_29332);
or UO_2600 (O_2600,N_25972,N_28272);
xor UO_2601 (O_2601,N_28734,N_28107);
or UO_2602 (O_2602,N_25931,N_28267);
xnor UO_2603 (O_2603,N_28678,N_29735);
nand UO_2604 (O_2604,N_29816,N_29575);
or UO_2605 (O_2605,N_28733,N_28669);
nand UO_2606 (O_2606,N_28555,N_26151);
xor UO_2607 (O_2607,N_26544,N_26012);
or UO_2608 (O_2608,N_25554,N_28469);
nor UO_2609 (O_2609,N_25930,N_24108);
or UO_2610 (O_2610,N_27725,N_27060);
xnor UO_2611 (O_2611,N_28356,N_27382);
nor UO_2612 (O_2612,N_26323,N_27254);
or UO_2613 (O_2613,N_29042,N_27591);
and UO_2614 (O_2614,N_28291,N_24030);
xor UO_2615 (O_2615,N_29221,N_28661);
nor UO_2616 (O_2616,N_28382,N_27158);
nand UO_2617 (O_2617,N_27530,N_26484);
xnor UO_2618 (O_2618,N_27618,N_25380);
nor UO_2619 (O_2619,N_27363,N_27539);
nor UO_2620 (O_2620,N_24845,N_27951);
nor UO_2621 (O_2621,N_28593,N_26610);
nor UO_2622 (O_2622,N_25722,N_27555);
nor UO_2623 (O_2623,N_27118,N_26443);
or UO_2624 (O_2624,N_27497,N_28925);
nor UO_2625 (O_2625,N_27680,N_27595);
xor UO_2626 (O_2626,N_26383,N_29353);
and UO_2627 (O_2627,N_29848,N_25843);
nor UO_2628 (O_2628,N_28624,N_27865);
xor UO_2629 (O_2629,N_27244,N_24054);
nor UO_2630 (O_2630,N_28790,N_29102);
nand UO_2631 (O_2631,N_29719,N_26243);
xor UO_2632 (O_2632,N_27000,N_27059);
nand UO_2633 (O_2633,N_24182,N_29257);
and UO_2634 (O_2634,N_29892,N_29317);
xor UO_2635 (O_2635,N_29024,N_28071);
nor UO_2636 (O_2636,N_27224,N_24686);
nor UO_2637 (O_2637,N_24265,N_28414);
nor UO_2638 (O_2638,N_29098,N_29361);
or UO_2639 (O_2639,N_25152,N_24619);
nand UO_2640 (O_2640,N_27804,N_27707);
and UO_2641 (O_2641,N_24700,N_29148);
and UO_2642 (O_2642,N_24856,N_28325);
nand UO_2643 (O_2643,N_26274,N_28466);
xor UO_2644 (O_2644,N_24329,N_29551);
xor UO_2645 (O_2645,N_29441,N_29429);
nor UO_2646 (O_2646,N_27597,N_27278);
or UO_2647 (O_2647,N_29080,N_26489);
xor UO_2648 (O_2648,N_25674,N_27834);
and UO_2649 (O_2649,N_29138,N_28635);
or UO_2650 (O_2650,N_27582,N_28350);
and UO_2651 (O_2651,N_25493,N_26700);
nand UO_2652 (O_2652,N_28605,N_25961);
nand UO_2653 (O_2653,N_25096,N_29628);
or UO_2654 (O_2654,N_26592,N_24559);
nand UO_2655 (O_2655,N_27788,N_25158);
nand UO_2656 (O_2656,N_25313,N_26583);
xor UO_2657 (O_2657,N_28175,N_27885);
nor UO_2658 (O_2658,N_29455,N_25508);
nor UO_2659 (O_2659,N_27232,N_28564);
nand UO_2660 (O_2660,N_26805,N_25999);
xor UO_2661 (O_2661,N_26882,N_28954);
xnor UO_2662 (O_2662,N_29020,N_28191);
and UO_2663 (O_2663,N_25715,N_27805);
or UO_2664 (O_2664,N_26856,N_28068);
nand UO_2665 (O_2665,N_26869,N_24131);
nor UO_2666 (O_2666,N_27383,N_29328);
and UO_2667 (O_2667,N_24430,N_25502);
or UO_2668 (O_2668,N_24395,N_26337);
nor UO_2669 (O_2669,N_25294,N_26601);
and UO_2670 (O_2670,N_25610,N_26476);
and UO_2671 (O_2671,N_28139,N_26832);
and UO_2672 (O_2672,N_24285,N_24768);
or UO_2673 (O_2673,N_24935,N_27828);
xor UO_2674 (O_2674,N_25424,N_24560);
xor UO_2675 (O_2675,N_29700,N_24022);
or UO_2676 (O_2676,N_28163,N_29379);
and UO_2677 (O_2677,N_28549,N_27223);
or UO_2678 (O_2678,N_27249,N_27661);
nor UO_2679 (O_2679,N_24790,N_24046);
nor UO_2680 (O_2680,N_27892,N_28403);
or UO_2681 (O_2681,N_25324,N_28772);
and UO_2682 (O_2682,N_24350,N_24844);
and UO_2683 (O_2683,N_24361,N_28806);
and UO_2684 (O_2684,N_25801,N_25878);
xor UO_2685 (O_2685,N_25232,N_26726);
nand UO_2686 (O_2686,N_24018,N_25879);
and UO_2687 (O_2687,N_29720,N_27250);
xor UO_2688 (O_2688,N_28943,N_27331);
nor UO_2689 (O_2689,N_27872,N_29810);
xor UO_2690 (O_2690,N_25219,N_25537);
xor UO_2691 (O_2691,N_27194,N_29266);
nor UO_2692 (O_2692,N_27538,N_28498);
xor UO_2693 (O_2693,N_26629,N_28680);
and UO_2694 (O_2694,N_29762,N_29154);
nand UO_2695 (O_2695,N_29654,N_25661);
xor UO_2696 (O_2696,N_26616,N_27507);
nand UO_2697 (O_2697,N_24688,N_29955);
or UO_2698 (O_2698,N_28759,N_25246);
or UO_2699 (O_2699,N_26359,N_28389);
or UO_2700 (O_2700,N_29283,N_28822);
nand UO_2701 (O_2701,N_24650,N_28614);
nand UO_2702 (O_2702,N_25321,N_24050);
and UO_2703 (O_2703,N_29659,N_26633);
nor UO_2704 (O_2704,N_24601,N_26772);
xnor UO_2705 (O_2705,N_26959,N_25334);
or UO_2706 (O_2706,N_24229,N_24174);
xnor UO_2707 (O_2707,N_29025,N_26446);
nor UO_2708 (O_2708,N_28560,N_27565);
nand UO_2709 (O_2709,N_29574,N_27388);
or UO_2710 (O_2710,N_29457,N_29430);
nor UO_2711 (O_2711,N_28092,N_28841);
or UO_2712 (O_2712,N_26582,N_25494);
or UO_2713 (O_2713,N_29109,N_28507);
and UO_2714 (O_2714,N_25281,N_29877);
nand UO_2715 (O_2715,N_25574,N_27749);
nor UO_2716 (O_2716,N_28346,N_25890);
nor UO_2717 (O_2717,N_27451,N_28458);
nand UO_2718 (O_2718,N_25789,N_28561);
xor UO_2719 (O_2719,N_26047,N_27469);
xor UO_2720 (O_2720,N_24568,N_27727);
xnor UO_2721 (O_2721,N_28375,N_28442);
or UO_2722 (O_2722,N_27216,N_26531);
and UO_2723 (O_2723,N_25206,N_27506);
nor UO_2724 (O_2724,N_25209,N_28345);
nor UO_2725 (O_2725,N_26186,N_28581);
nand UO_2726 (O_2726,N_27840,N_29459);
xor UO_2727 (O_2727,N_27315,N_24592);
and UO_2728 (O_2728,N_24502,N_29751);
nand UO_2729 (O_2729,N_25034,N_25945);
and UO_2730 (O_2730,N_27172,N_27734);
nor UO_2731 (O_2731,N_24414,N_25212);
or UO_2732 (O_2732,N_28850,N_29914);
nand UO_2733 (O_2733,N_26972,N_25700);
nor UO_2734 (O_2734,N_26279,N_27231);
nor UO_2735 (O_2735,N_25049,N_25934);
or UO_2736 (O_2736,N_29187,N_27798);
and UO_2737 (O_2737,N_25968,N_26828);
and UO_2738 (O_2738,N_26150,N_28129);
xor UO_2739 (O_2739,N_28400,N_26138);
nor UO_2740 (O_2740,N_27374,N_25214);
nand UO_2741 (O_2741,N_26810,N_24029);
or UO_2742 (O_2742,N_25820,N_29323);
xnor UO_2743 (O_2743,N_24961,N_26737);
xor UO_2744 (O_2744,N_28098,N_29554);
nand UO_2745 (O_2745,N_27068,N_25004);
nand UO_2746 (O_2746,N_27813,N_26322);
xnor UO_2747 (O_2747,N_28248,N_24597);
or UO_2748 (O_2748,N_28019,N_28578);
or UO_2749 (O_2749,N_24032,N_26565);
nor UO_2750 (O_2750,N_27465,N_25788);
nor UO_2751 (O_2751,N_27274,N_26515);
nor UO_2752 (O_2752,N_29990,N_26513);
xnor UO_2753 (O_2753,N_29789,N_28207);
or UO_2754 (O_2754,N_29966,N_24878);
xor UO_2755 (O_2755,N_29245,N_26214);
nor UO_2756 (O_2756,N_24626,N_28225);
nand UO_2757 (O_2757,N_25904,N_28632);
and UO_2758 (O_2758,N_27459,N_29767);
nor UO_2759 (O_2759,N_28894,N_27851);
and UO_2760 (O_2760,N_25836,N_25958);
nor UO_2761 (O_2761,N_26757,N_26754);
nand UO_2762 (O_2762,N_28268,N_28909);
xnor UO_2763 (O_2763,N_29569,N_29209);
nand UO_2764 (O_2764,N_25675,N_25347);
nand UO_2765 (O_2765,N_28143,N_25620);
and UO_2766 (O_2766,N_28604,N_25341);
or UO_2767 (O_2767,N_25255,N_25119);
xnor UO_2768 (O_2768,N_25568,N_28798);
and UO_2769 (O_2769,N_24077,N_29256);
or UO_2770 (O_2770,N_28536,N_25813);
and UO_2771 (O_2771,N_26628,N_27698);
or UO_2772 (O_2772,N_27718,N_25826);
nand UO_2773 (O_2773,N_24997,N_26915);
and UO_2774 (O_2774,N_25445,N_25729);
nor UO_2775 (O_2775,N_29597,N_28266);
nor UO_2776 (O_2776,N_28463,N_28333);
xor UO_2777 (O_2777,N_26609,N_24422);
or UO_2778 (O_2778,N_29090,N_28012);
and UO_2779 (O_2779,N_25797,N_25348);
nand UO_2780 (O_2780,N_24033,N_28449);
and UO_2781 (O_2781,N_27424,N_25340);
xnor UO_2782 (O_2782,N_27616,N_26100);
nand UO_2783 (O_2783,N_26743,N_27515);
or UO_2784 (O_2784,N_27170,N_29570);
and UO_2785 (O_2785,N_26001,N_25919);
and UO_2786 (O_2786,N_28258,N_26250);
nand UO_2787 (O_2787,N_29304,N_27463);
and UO_2788 (O_2788,N_24591,N_26802);
or UO_2789 (O_2789,N_28313,N_24185);
nand UO_2790 (O_2790,N_27461,N_24102);
and UO_2791 (O_2791,N_26006,N_29546);
xor UO_2792 (O_2792,N_27033,N_25876);
xor UO_2793 (O_2793,N_28974,N_28245);
and UO_2794 (O_2794,N_25549,N_27722);
and UO_2795 (O_2795,N_27747,N_29387);
or UO_2796 (O_2796,N_25520,N_26498);
and UO_2797 (O_2797,N_26024,N_24987);
or UO_2798 (O_2798,N_26282,N_28580);
xor UO_2799 (O_2799,N_25939,N_29295);
and UO_2800 (O_2800,N_28652,N_28718);
xnor UO_2801 (O_2801,N_25319,N_28341);
xor UO_2802 (O_2802,N_29364,N_27301);
and UO_2803 (O_2803,N_27757,N_24646);
xor UO_2804 (O_2804,N_24309,N_27175);
and UO_2805 (O_2805,N_25415,N_28125);
and UO_2806 (O_2806,N_28890,N_28782);
nor UO_2807 (O_2807,N_24477,N_27868);
nor UO_2808 (O_2808,N_25596,N_27970);
xor UO_2809 (O_2809,N_27467,N_29757);
or UO_2810 (O_2810,N_25227,N_29996);
xnor UO_2811 (O_2811,N_26611,N_25398);
and UO_2812 (O_2812,N_26711,N_27981);
nor UO_2813 (O_2813,N_28009,N_28320);
nand UO_2814 (O_2814,N_29864,N_25641);
or UO_2815 (O_2815,N_29427,N_27387);
nor UO_2816 (O_2816,N_29028,N_29120);
nand UO_2817 (O_2817,N_28606,N_25694);
and UO_2818 (O_2818,N_24002,N_26473);
and UO_2819 (O_2819,N_25691,N_28281);
nand UO_2820 (O_2820,N_29642,N_24037);
and UO_2821 (O_2821,N_29855,N_28295);
and UO_2822 (O_2822,N_27450,N_27762);
nand UO_2823 (O_2823,N_29830,N_25290);
xor UO_2824 (O_2824,N_24052,N_26822);
or UO_2825 (O_2825,N_26099,N_28569);
or UO_2826 (O_2826,N_29030,N_28154);
nor UO_2827 (O_2827,N_29637,N_29545);
nor UO_2828 (O_2828,N_29683,N_25992);
nand UO_2829 (O_2829,N_26936,N_29610);
or UO_2830 (O_2830,N_29585,N_25870);
nand UO_2831 (O_2831,N_26676,N_25252);
or UO_2832 (O_2832,N_25883,N_26732);
nor UO_2833 (O_2833,N_24939,N_25793);
or UO_2834 (O_2834,N_25505,N_29660);
or UO_2835 (O_2835,N_26160,N_28473);
nand UO_2836 (O_2836,N_26693,N_28831);
nor UO_2837 (O_2837,N_26461,N_29696);
xor UO_2838 (O_2838,N_28491,N_25448);
nor UO_2839 (O_2839,N_25860,N_28354);
xor UO_2840 (O_2840,N_29680,N_24514);
nor UO_2841 (O_2841,N_25752,N_27816);
nor UO_2842 (O_2842,N_26525,N_25772);
and UO_2843 (O_2843,N_27731,N_28534);
xnor UO_2844 (O_2844,N_28510,N_27030);
nor UO_2845 (O_2845,N_29351,N_29814);
xor UO_2846 (O_2846,N_27612,N_29606);
and UO_2847 (O_2847,N_24622,N_29509);
and UO_2848 (O_2848,N_28601,N_29476);
or UO_2849 (O_2849,N_27654,N_24581);
and UO_2850 (O_2850,N_29442,N_25135);
nand UO_2851 (O_2851,N_27543,N_24903);
xnor UO_2852 (O_2852,N_25165,N_25716);
xor UO_2853 (O_2853,N_26932,N_24948);
or UO_2854 (O_2854,N_27586,N_26007);
or UO_2855 (O_2855,N_26967,N_29857);
nand UO_2856 (O_2856,N_26367,N_27719);
nor UO_2857 (O_2857,N_25791,N_29553);
xor UO_2858 (O_2858,N_29275,N_25384);
or UO_2859 (O_2859,N_27406,N_25405);
or UO_2860 (O_2860,N_28287,N_27869);
or UO_2861 (O_2861,N_27957,N_27303);
xnor UO_2862 (O_2862,N_28603,N_28620);
xnor UO_2863 (O_2863,N_27677,N_29228);
nor UO_2864 (O_2864,N_28977,N_29128);
and UO_2865 (O_2865,N_24065,N_29604);
and UO_2866 (O_2866,N_29083,N_29853);
xnor UO_2867 (O_2867,N_27401,N_27286);
xnor UO_2868 (O_2868,N_27265,N_27653);
xnor UO_2869 (O_2869,N_25808,N_28630);
xor UO_2870 (O_2870,N_29354,N_27745);
and UO_2871 (O_2871,N_28952,N_28657);
and UO_2872 (O_2872,N_25971,N_28899);
or UO_2873 (O_2873,N_24415,N_26771);
nand UO_2874 (O_2874,N_25798,N_24792);
or UO_2875 (O_2875,N_24742,N_27338);
nor UO_2876 (O_2876,N_25036,N_27002);
xor UO_2877 (O_2877,N_25468,N_26636);
xor UO_2878 (O_2878,N_27253,N_28629);
or UO_2879 (O_2879,N_29346,N_25651);
nor UO_2880 (O_2880,N_27934,N_26078);
nor UO_2881 (O_2881,N_27094,N_24680);
or UO_2882 (O_2882,N_27310,N_25530);
xnor UO_2883 (O_2883,N_26940,N_27075);
nand UO_2884 (O_2884,N_26763,N_26414);
nand UO_2885 (O_2885,N_28264,N_29439);
xnor UO_2886 (O_2886,N_27846,N_27361);
and UO_2887 (O_2887,N_25188,N_25625);
nand UO_2888 (O_2888,N_29095,N_27269);
or UO_2889 (O_2889,N_28935,N_29988);
and UO_2890 (O_2890,N_26432,N_25196);
and UO_2891 (O_2891,N_27524,N_25918);
nand UO_2892 (O_2892,N_26563,N_29464);
nor UO_2893 (O_2893,N_29089,N_26545);
and UO_2894 (O_2894,N_26535,N_29698);
or UO_2895 (O_2895,N_27854,N_27701);
or UO_2896 (O_2896,N_26419,N_28035);
nand UO_2897 (O_2897,N_24078,N_24528);
nand UO_2898 (O_2898,N_24252,N_28582);
xnor UO_2899 (O_2899,N_25507,N_27990);
and UO_2900 (O_2900,N_28496,N_25655);
nand UO_2901 (O_2901,N_24060,N_28907);
xnor UO_2902 (O_2902,N_26114,N_25174);
xor UO_2903 (O_2903,N_24748,N_27683);
and UO_2904 (O_2904,N_29320,N_26368);
and UO_2905 (O_2905,N_29811,N_28749);
and UO_2906 (O_2906,N_26092,N_26549);
and UO_2907 (O_2907,N_27307,N_27982);
nand UO_2908 (O_2908,N_29243,N_27886);
nand UO_2909 (O_2909,N_29058,N_28188);
nor UO_2910 (O_2910,N_25699,N_25441);
xnor UO_2911 (O_2911,N_25367,N_27918);
nand UO_2912 (O_2912,N_24088,N_25362);
nand UO_2913 (O_2913,N_28365,N_24295);
xor UO_2914 (O_2914,N_29799,N_29164);
or UO_2915 (O_2915,N_24224,N_27576);
and UO_2916 (O_2916,N_28480,N_29867);
and UO_2917 (O_2917,N_25414,N_26103);
nand UO_2918 (O_2918,N_24979,N_27822);
xor UO_2919 (O_2919,N_25584,N_24158);
or UO_2920 (O_2920,N_25906,N_27628);
nand UO_2921 (O_2921,N_29002,N_25084);
nand UO_2922 (O_2922,N_24898,N_28665);
or UO_2923 (O_2923,N_27334,N_28187);
and UO_2924 (O_2924,N_29493,N_28608);
or UO_2925 (O_2925,N_24908,N_24980);
nand UO_2926 (O_2926,N_27656,N_29518);
xnor UO_2927 (O_2927,N_25721,N_25005);
nor UO_2928 (O_2928,N_27809,N_24931);
xor UO_2929 (O_2929,N_27051,N_24205);
or UO_2930 (O_2930,N_24072,N_28273);
nand UO_2931 (O_2931,N_27178,N_29322);
nor UO_2932 (O_2932,N_28820,N_25540);
nor UO_2933 (O_2933,N_24955,N_25773);
xor UO_2934 (O_2934,N_28289,N_29770);
or UO_2935 (O_2935,N_29474,N_26627);
xnor UO_2936 (O_2936,N_24386,N_28434);
or UO_2937 (O_2937,N_27316,N_25287);
xnor UO_2938 (O_2938,N_26575,N_26042);
nand UO_2939 (O_2939,N_27771,N_24180);
xnor UO_2940 (O_2940,N_25249,N_26408);
or UO_2941 (O_2941,N_24694,N_24346);
and UO_2942 (O_2942,N_26034,N_27365);
or UO_2943 (O_2943,N_26127,N_29950);
nand UO_2944 (O_2944,N_27205,N_24137);
and UO_2945 (O_2945,N_27505,N_24493);
or UO_2946 (O_2946,N_25263,N_29096);
and UO_2947 (O_2947,N_27855,N_26023);
nand UO_2948 (O_2948,N_29033,N_26453);
xor UO_2949 (O_2949,N_26770,N_28405);
and UO_2950 (O_2950,N_28095,N_24003);
nor UO_2951 (O_2951,N_26522,N_24749);
nor UO_2952 (O_2952,N_29577,N_29730);
nand UO_2953 (O_2953,N_25802,N_29612);
nand UO_2954 (O_2954,N_27577,N_26645);
xor UO_2955 (O_2955,N_24425,N_29494);
nand UO_2956 (O_2956,N_25216,N_24058);
nand UO_2957 (O_2957,N_27349,N_27069);
nand UO_2958 (O_2958,N_27906,N_27195);
xnor UO_2959 (O_2959,N_24168,N_27666);
and UO_2960 (O_2960,N_29949,N_24379);
and UO_2961 (O_2961,N_29422,N_27553);
nor UO_2962 (O_2962,N_24534,N_28702);
and UO_2963 (O_2963,N_24959,N_24094);
or UO_2964 (O_2964,N_26872,N_27756);
nand UO_2965 (O_2965,N_26900,N_25734);
xnor UO_2966 (O_2966,N_27845,N_26122);
nor UO_2967 (O_2967,N_25464,N_27227);
xor UO_2968 (O_2968,N_26051,N_25636);
and UO_2969 (O_2969,N_27037,N_28054);
nor UO_2970 (O_2970,N_27637,N_24970);
or UO_2971 (O_2971,N_24181,N_29488);
nor UO_2972 (O_2972,N_25746,N_29581);
and UO_2973 (O_2973,N_26310,N_25383);
and UO_2974 (O_2974,N_24118,N_29922);
xnor UO_2975 (O_2975,N_24441,N_28599);
and UO_2976 (O_2976,N_29523,N_29126);
nor UO_2977 (O_2977,N_27335,N_28752);
or UO_2978 (O_2978,N_27711,N_29303);
and UO_2979 (O_2979,N_25315,N_28455);
xnor UO_2980 (O_2980,N_27299,N_25516);
nor UO_2981 (O_2981,N_24990,N_26756);
xnor UO_2982 (O_2982,N_27977,N_28097);
or UO_2983 (O_2983,N_24219,N_25743);
xnor UO_2984 (O_2984,N_25684,N_26146);
nor UO_2985 (O_2985,N_28846,N_29674);
nand UO_2986 (O_2986,N_26091,N_26348);
xnor UO_2987 (O_2987,N_24097,N_29162);
nand UO_2988 (O_2988,N_29034,N_25364);
nand UO_2989 (O_2989,N_26863,N_24208);
nor UO_2990 (O_2990,N_24326,N_29214);
nand UO_2991 (O_2991,N_29861,N_28499);
and UO_2992 (O_2992,N_26564,N_25686);
or UO_2993 (O_2993,N_25316,N_25269);
nand UO_2994 (O_2994,N_26820,N_26835);
or UO_2995 (O_2995,N_25198,N_24963);
or UO_2996 (O_2996,N_27624,N_29842);
xor UO_2997 (O_2997,N_26643,N_29851);
nor UO_2998 (O_2998,N_24312,N_28901);
and UO_2999 (O_2999,N_24525,N_29310);
and UO_3000 (O_3000,N_27092,N_25278);
nor UO_3001 (O_3001,N_29178,N_28739);
and UO_3002 (O_3002,N_29500,N_24886);
and UO_3003 (O_3003,N_24588,N_28118);
xnor UO_3004 (O_3004,N_24278,N_29459);
and UO_3005 (O_3005,N_27122,N_25697);
and UO_3006 (O_3006,N_25080,N_25626);
and UO_3007 (O_3007,N_25338,N_27302);
xor UO_3008 (O_3008,N_29668,N_29272);
nor UO_3009 (O_3009,N_24225,N_25051);
and UO_3010 (O_3010,N_28835,N_24548);
nand UO_3011 (O_3011,N_28679,N_29756);
xor UO_3012 (O_3012,N_27959,N_26380);
and UO_3013 (O_3013,N_24371,N_27496);
and UO_3014 (O_3014,N_26939,N_25583);
nand UO_3015 (O_3015,N_27490,N_24607);
xor UO_3016 (O_3016,N_27075,N_27635);
nor UO_3017 (O_3017,N_28241,N_25114);
xor UO_3018 (O_3018,N_27467,N_25909);
nor UO_3019 (O_3019,N_29379,N_25287);
or UO_3020 (O_3020,N_29370,N_24696);
and UO_3021 (O_3021,N_24922,N_27588);
xnor UO_3022 (O_3022,N_29362,N_25048);
and UO_3023 (O_3023,N_27140,N_24706);
or UO_3024 (O_3024,N_24091,N_24105);
nand UO_3025 (O_3025,N_29057,N_24797);
xor UO_3026 (O_3026,N_25993,N_29313);
xnor UO_3027 (O_3027,N_26248,N_28076);
nor UO_3028 (O_3028,N_28173,N_26356);
xnor UO_3029 (O_3029,N_29202,N_27257);
xnor UO_3030 (O_3030,N_26866,N_28229);
xor UO_3031 (O_3031,N_28963,N_26577);
nand UO_3032 (O_3032,N_25205,N_26520);
nor UO_3033 (O_3033,N_28893,N_26465);
nand UO_3034 (O_3034,N_26771,N_29184);
and UO_3035 (O_3035,N_25494,N_28739);
or UO_3036 (O_3036,N_26632,N_27973);
xnor UO_3037 (O_3037,N_26622,N_28430);
xor UO_3038 (O_3038,N_27734,N_26134);
xor UO_3039 (O_3039,N_25060,N_25857);
nor UO_3040 (O_3040,N_29213,N_26372);
nor UO_3041 (O_3041,N_25899,N_25136);
xor UO_3042 (O_3042,N_27465,N_25085);
nor UO_3043 (O_3043,N_26084,N_24119);
or UO_3044 (O_3044,N_24048,N_25008);
and UO_3045 (O_3045,N_27472,N_29741);
or UO_3046 (O_3046,N_26653,N_24202);
or UO_3047 (O_3047,N_24214,N_29141);
nor UO_3048 (O_3048,N_24102,N_24927);
xor UO_3049 (O_3049,N_24336,N_29179);
nand UO_3050 (O_3050,N_28869,N_24916);
and UO_3051 (O_3051,N_29382,N_25326);
nand UO_3052 (O_3052,N_24033,N_29933);
or UO_3053 (O_3053,N_24993,N_24805);
or UO_3054 (O_3054,N_28284,N_25121);
or UO_3055 (O_3055,N_25193,N_28030);
xor UO_3056 (O_3056,N_29095,N_27767);
xnor UO_3057 (O_3057,N_27168,N_28003);
xnor UO_3058 (O_3058,N_24267,N_24375);
and UO_3059 (O_3059,N_29865,N_28753);
nor UO_3060 (O_3060,N_28472,N_27094);
nor UO_3061 (O_3061,N_29545,N_24926);
xor UO_3062 (O_3062,N_29954,N_26923);
or UO_3063 (O_3063,N_28132,N_29974);
and UO_3064 (O_3064,N_28819,N_26892);
xor UO_3065 (O_3065,N_24889,N_26891);
nand UO_3066 (O_3066,N_27954,N_24871);
and UO_3067 (O_3067,N_26055,N_25588);
xnor UO_3068 (O_3068,N_24373,N_25517);
xor UO_3069 (O_3069,N_26791,N_26907);
and UO_3070 (O_3070,N_25115,N_27921);
and UO_3071 (O_3071,N_24372,N_26782);
or UO_3072 (O_3072,N_26899,N_24251);
xnor UO_3073 (O_3073,N_24978,N_28055);
or UO_3074 (O_3074,N_25577,N_29159);
nor UO_3075 (O_3075,N_28535,N_26113);
xor UO_3076 (O_3076,N_25411,N_27379);
nor UO_3077 (O_3077,N_28619,N_29266);
nand UO_3078 (O_3078,N_26239,N_24986);
xor UO_3079 (O_3079,N_27040,N_27977);
xor UO_3080 (O_3080,N_25877,N_24285);
and UO_3081 (O_3081,N_24127,N_29054);
nor UO_3082 (O_3082,N_27293,N_29231);
nor UO_3083 (O_3083,N_29604,N_26694);
nand UO_3084 (O_3084,N_24154,N_25192);
or UO_3085 (O_3085,N_25035,N_24062);
or UO_3086 (O_3086,N_29475,N_28973);
or UO_3087 (O_3087,N_29254,N_27917);
xnor UO_3088 (O_3088,N_24199,N_28490);
xor UO_3089 (O_3089,N_29117,N_25595);
nand UO_3090 (O_3090,N_26564,N_27401);
nor UO_3091 (O_3091,N_27860,N_29693);
nand UO_3092 (O_3092,N_24774,N_25329);
nand UO_3093 (O_3093,N_26679,N_28111);
xnor UO_3094 (O_3094,N_25304,N_28507);
xnor UO_3095 (O_3095,N_24837,N_27903);
and UO_3096 (O_3096,N_28356,N_25666);
nor UO_3097 (O_3097,N_28540,N_26897);
or UO_3098 (O_3098,N_25110,N_27779);
xor UO_3099 (O_3099,N_24727,N_25021);
nor UO_3100 (O_3100,N_27964,N_25849);
and UO_3101 (O_3101,N_27514,N_24994);
xor UO_3102 (O_3102,N_28600,N_24643);
nor UO_3103 (O_3103,N_26229,N_25489);
nor UO_3104 (O_3104,N_26934,N_29531);
nor UO_3105 (O_3105,N_29320,N_26780);
and UO_3106 (O_3106,N_26832,N_25056);
nand UO_3107 (O_3107,N_29837,N_27523);
and UO_3108 (O_3108,N_24817,N_24274);
nor UO_3109 (O_3109,N_26977,N_25308);
and UO_3110 (O_3110,N_27270,N_28068);
nand UO_3111 (O_3111,N_29548,N_26064);
xor UO_3112 (O_3112,N_24155,N_26804);
or UO_3113 (O_3113,N_26070,N_28988);
or UO_3114 (O_3114,N_29612,N_24351);
or UO_3115 (O_3115,N_25820,N_26854);
and UO_3116 (O_3116,N_28595,N_29419);
xnor UO_3117 (O_3117,N_29739,N_26953);
and UO_3118 (O_3118,N_24692,N_29782);
or UO_3119 (O_3119,N_28373,N_25593);
nand UO_3120 (O_3120,N_27019,N_29637);
nand UO_3121 (O_3121,N_25479,N_27263);
nand UO_3122 (O_3122,N_25412,N_27719);
and UO_3123 (O_3123,N_24110,N_24800);
and UO_3124 (O_3124,N_24058,N_27802);
nor UO_3125 (O_3125,N_28391,N_26437);
nor UO_3126 (O_3126,N_27263,N_25369);
xor UO_3127 (O_3127,N_27306,N_29383);
xnor UO_3128 (O_3128,N_27987,N_29094);
nor UO_3129 (O_3129,N_27882,N_24512);
nor UO_3130 (O_3130,N_27792,N_25052);
nor UO_3131 (O_3131,N_28005,N_25504);
xnor UO_3132 (O_3132,N_26895,N_24752);
or UO_3133 (O_3133,N_24019,N_29310);
and UO_3134 (O_3134,N_29127,N_24084);
nand UO_3135 (O_3135,N_28677,N_25645);
or UO_3136 (O_3136,N_24066,N_28581);
xnor UO_3137 (O_3137,N_24374,N_25663);
nor UO_3138 (O_3138,N_29888,N_27812);
nand UO_3139 (O_3139,N_26175,N_29682);
or UO_3140 (O_3140,N_25318,N_24409);
and UO_3141 (O_3141,N_29202,N_26118);
nor UO_3142 (O_3142,N_24999,N_27233);
nand UO_3143 (O_3143,N_27784,N_24563);
or UO_3144 (O_3144,N_24947,N_28165);
and UO_3145 (O_3145,N_28550,N_28128);
xor UO_3146 (O_3146,N_25125,N_29048);
nand UO_3147 (O_3147,N_27799,N_27559);
or UO_3148 (O_3148,N_29958,N_28474);
xnor UO_3149 (O_3149,N_29131,N_24590);
nor UO_3150 (O_3150,N_25438,N_27651);
or UO_3151 (O_3151,N_28261,N_25856);
or UO_3152 (O_3152,N_26436,N_27948);
and UO_3153 (O_3153,N_26431,N_29106);
or UO_3154 (O_3154,N_25783,N_29307);
nor UO_3155 (O_3155,N_24984,N_27622);
xnor UO_3156 (O_3156,N_24394,N_27394);
xor UO_3157 (O_3157,N_25154,N_27711);
and UO_3158 (O_3158,N_26650,N_28086);
or UO_3159 (O_3159,N_26420,N_26894);
or UO_3160 (O_3160,N_24389,N_24281);
and UO_3161 (O_3161,N_29956,N_29490);
nand UO_3162 (O_3162,N_29348,N_26587);
and UO_3163 (O_3163,N_24830,N_27961);
nor UO_3164 (O_3164,N_24522,N_29226);
nand UO_3165 (O_3165,N_25760,N_28857);
and UO_3166 (O_3166,N_28918,N_24456);
or UO_3167 (O_3167,N_28344,N_25765);
or UO_3168 (O_3168,N_26900,N_29349);
or UO_3169 (O_3169,N_25756,N_24753);
or UO_3170 (O_3170,N_28436,N_25283);
nand UO_3171 (O_3171,N_26159,N_28054);
nand UO_3172 (O_3172,N_24304,N_27221);
and UO_3173 (O_3173,N_25755,N_26904);
xor UO_3174 (O_3174,N_24545,N_24473);
nor UO_3175 (O_3175,N_28845,N_26881);
xnor UO_3176 (O_3176,N_26467,N_24335);
xnor UO_3177 (O_3177,N_27162,N_24340);
nor UO_3178 (O_3178,N_24116,N_29047);
or UO_3179 (O_3179,N_26148,N_25578);
xnor UO_3180 (O_3180,N_28558,N_28683);
nor UO_3181 (O_3181,N_27819,N_24013);
and UO_3182 (O_3182,N_26370,N_26568);
or UO_3183 (O_3183,N_24953,N_29933);
or UO_3184 (O_3184,N_29097,N_28643);
nand UO_3185 (O_3185,N_24063,N_24486);
xnor UO_3186 (O_3186,N_25657,N_24284);
nand UO_3187 (O_3187,N_27675,N_25758);
nor UO_3188 (O_3188,N_26429,N_25225);
nor UO_3189 (O_3189,N_27221,N_26262);
xnor UO_3190 (O_3190,N_25696,N_24890);
and UO_3191 (O_3191,N_28552,N_25153);
xnor UO_3192 (O_3192,N_29873,N_29392);
nor UO_3193 (O_3193,N_27452,N_25518);
xnor UO_3194 (O_3194,N_28461,N_25980);
nor UO_3195 (O_3195,N_27612,N_27311);
nand UO_3196 (O_3196,N_25193,N_24258);
nor UO_3197 (O_3197,N_28183,N_26149);
nand UO_3198 (O_3198,N_26292,N_29059);
nand UO_3199 (O_3199,N_24893,N_24753);
or UO_3200 (O_3200,N_28200,N_28231);
xnor UO_3201 (O_3201,N_29456,N_25030);
and UO_3202 (O_3202,N_24394,N_25473);
and UO_3203 (O_3203,N_26569,N_25736);
and UO_3204 (O_3204,N_29924,N_27932);
or UO_3205 (O_3205,N_24641,N_29836);
or UO_3206 (O_3206,N_28516,N_24681);
and UO_3207 (O_3207,N_28637,N_24730);
xnor UO_3208 (O_3208,N_25529,N_29357);
nor UO_3209 (O_3209,N_28148,N_28933);
or UO_3210 (O_3210,N_29186,N_24102);
nand UO_3211 (O_3211,N_26472,N_27766);
and UO_3212 (O_3212,N_28055,N_28953);
nand UO_3213 (O_3213,N_28974,N_29260);
or UO_3214 (O_3214,N_28046,N_25348);
xor UO_3215 (O_3215,N_28609,N_29306);
and UO_3216 (O_3216,N_24001,N_27190);
or UO_3217 (O_3217,N_27837,N_29321);
xor UO_3218 (O_3218,N_26316,N_26589);
and UO_3219 (O_3219,N_29752,N_29116);
xnor UO_3220 (O_3220,N_25899,N_26772);
or UO_3221 (O_3221,N_26386,N_26518);
nor UO_3222 (O_3222,N_28882,N_29800);
and UO_3223 (O_3223,N_24267,N_26404);
and UO_3224 (O_3224,N_25659,N_24754);
nand UO_3225 (O_3225,N_24279,N_24481);
and UO_3226 (O_3226,N_26443,N_29660);
nor UO_3227 (O_3227,N_25749,N_27555);
xnor UO_3228 (O_3228,N_27279,N_29164);
and UO_3229 (O_3229,N_27092,N_28197);
and UO_3230 (O_3230,N_27387,N_28380);
nor UO_3231 (O_3231,N_28635,N_27102);
nor UO_3232 (O_3232,N_27240,N_28111);
nor UO_3233 (O_3233,N_25074,N_29220);
xnor UO_3234 (O_3234,N_26390,N_25239);
nor UO_3235 (O_3235,N_25626,N_29935);
and UO_3236 (O_3236,N_28135,N_25086);
or UO_3237 (O_3237,N_27473,N_27758);
xnor UO_3238 (O_3238,N_27021,N_28605);
xor UO_3239 (O_3239,N_24913,N_25839);
xnor UO_3240 (O_3240,N_25096,N_24741);
nand UO_3241 (O_3241,N_25609,N_29426);
nand UO_3242 (O_3242,N_27986,N_26275);
or UO_3243 (O_3243,N_24615,N_26265);
and UO_3244 (O_3244,N_29666,N_29071);
xnor UO_3245 (O_3245,N_27858,N_28018);
nand UO_3246 (O_3246,N_24650,N_27556);
and UO_3247 (O_3247,N_26393,N_25430);
or UO_3248 (O_3248,N_28019,N_24565);
xor UO_3249 (O_3249,N_24230,N_24814);
nor UO_3250 (O_3250,N_27727,N_29101);
xnor UO_3251 (O_3251,N_28223,N_24882);
nand UO_3252 (O_3252,N_25810,N_27940);
nor UO_3253 (O_3253,N_29348,N_26220);
xor UO_3254 (O_3254,N_26274,N_29252);
or UO_3255 (O_3255,N_26283,N_24572);
nor UO_3256 (O_3256,N_28194,N_27301);
xnor UO_3257 (O_3257,N_24138,N_26227);
xor UO_3258 (O_3258,N_29188,N_29318);
or UO_3259 (O_3259,N_25140,N_24831);
and UO_3260 (O_3260,N_26450,N_25092);
xor UO_3261 (O_3261,N_26043,N_29419);
or UO_3262 (O_3262,N_24684,N_27313);
nand UO_3263 (O_3263,N_26390,N_27589);
or UO_3264 (O_3264,N_28505,N_24223);
nor UO_3265 (O_3265,N_26875,N_26858);
nor UO_3266 (O_3266,N_24086,N_29032);
or UO_3267 (O_3267,N_26332,N_25992);
and UO_3268 (O_3268,N_27930,N_27048);
or UO_3269 (O_3269,N_24380,N_25307);
nor UO_3270 (O_3270,N_24959,N_27957);
and UO_3271 (O_3271,N_28459,N_25900);
or UO_3272 (O_3272,N_24231,N_24276);
or UO_3273 (O_3273,N_29566,N_27320);
or UO_3274 (O_3274,N_24435,N_29805);
nand UO_3275 (O_3275,N_29197,N_25923);
nand UO_3276 (O_3276,N_27342,N_28209);
nand UO_3277 (O_3277,N_24797,N_24214);
xor UO_3278 (O_3278,N_28159,N_28840);
nand UO_3279 (O_3279,N_27780,N_29777);
nand UO_3280 (O_3280,N_24476,N_28668);
and UO_3281 (O_3281,N_26014,N_27440);
and UO_3282 (O_3282,N_28154,N_24777);
and UO_3283 (O_3283,N_27408,N_26641);
xor UO_3284 (O_3284,N_26246,N_29319);
or UO_3285 (O_3285,N_28536,N_26605);
nor UO_3286 (O_3286,N_24284,N_29746);
or UO_3287 (O_3287,N_28548,N_27642);
xnor UO_3288 (O_3288,N_25257,N_25044);
and UO_3289 (O_3289,N_25401,N_28125);
or UO_3290 (O_3290,N_25695,N_24815);
xor UO_3291 (O_3291,N_27707,N_25046);
xor UO_3292 (O_3292,N_28143,N_27861);
xor UO_3293 (O_3293,N_29029,N_25211);
or UO_3294 (O_3294,N_26811,N_24958);
nand UO_3295 (O_3295,N_28449,N_24730);
xor UO_3296 (O_3296,N_25088,N_28088);
xor UO_3297 (O_3297,N_25406,N_28952);
nand UO_3298 (O_3298,N_27927,N_25933);
xor UO_3299 (O_3299,N_24340,N_27291);
nor UO_3300 (O_3300,N_28377,N_28011);
and UO_3301 (O_3301,N_26052,N_29647);
nand UO_3302 (O_3302,N_27962,N_25655);
nand UO_3303 (O_3303,N_25931,N_26392);
or UO_3304 (O_3304,N_27842,N_24913);
nand UO_3305 (O_3305,N_25759,N_27896);
nor UO_3306 (O_3306,N_26895,N_28963);
nand UO_3307 (O_3307,N_25021,N_25433);
or UO_3308 (O_3308,N_25092,N_29267);
and UO_3309 (O_3309,N_25348,N_24215);
nor UO_3310 (O_3310,N_26510,N_27317);
nand UO_3311 (O_3311,N_25741,N_25839);
and UO_3312 (O_3312,N_27721,N_25874);
and UO_3313 (O_3313,N_28939,N_26030);
and UO_3314 (O_3314,N_24231,N_25930);
nand UO_3315 (O_3315,N_27817,N_25203);
and UO_3316 (O_3316,N_26581,N_25126);
xnor UO_3317 (O_3317,N_27041,N_28257);
xor UO_3318 (O_3318,N_25472,N_25143);
nand UO_3319 (O_3319,N_25150,N_24332);
or UO_3320 (O_3320,N_29351,N_26222);
xor UO_3321 (O_3321,N_24594,N_25149);
nor UO_3322 (O_3322,N_26232,N_27826);
nor UO_3323 (O_3323,N_26652,N_26765);
or UO_3324 (O_3324,N_28300,N_27596);
nor UO_3325 (O_3325,N_26119,N_29362);
xor UO_3326 (O_3326,N_25688,N_24174);
xnor UO_3327 (O_3327,N_26614,N_26357);
or UO_3328 (O_3328,N_27796,N_28383);
and UO_3329 (O_3329,N_25171,N_28230);
nand UO_3330 (O_3330,N_27463,N_28739);
nor UO_3331 (O_3331,N_25951,N_29583);
xor UO_3332 (O_3332,N_28706,N_26792);
nand UO_3333 (O_3333,N_26124,N_28561);
xnor UO_3334 (O_3334,N_28116,N_27543);
and UO_3335 (O_3335,N_26381,N_28861);
nor UO_3336 (O_3336,N_27618,N_27037);
or UO_3337 (O_3337,N_28646,N_25874);
or UO_3338 (O_3338,N_27594,N_27529);
and UO_3339 (O_3339,N_25197,N_28006);
nor UO_3340 (O_3340,N_27145,N_28441);
and UO_3341 (O_3341,N_25468,N_28902);
nor UO_3342 (O_3342,N_29529,N_26026);
xnor UO_3343 (O_3343,N_24917,N_25312);
nand UO_3344 (O_3344,N_27731,N_25498);
nor UO_3345 (O_3345,N_27217,N_24321);
xnor UO_3346 (O_3346,N_26601,N_29986);
or UO_3347 (O_3347,N_29767,N_29603);
nor UO_3348 (O_3348,N_29895,N_29012);
nor UO_3349 (O_3349,N_24901,N_28255);
and UO_3350 (O_3350,N_29712,N_29661);
nor UO_3351 (O_3351,N_27360,N_27988);
or UO_3352 (O_3352,N_25805,N_24269);
nand UO_3353 (O_3353,N_28164,N_28915);
or UO_3354 (O_3354,N_27000,N_25289);
or UO_3355 (O_3355,N_27756,N_25181);
nand UO_3356 (O_3356,N_28498,N_28207);
or UO_3357 (O_3357,N_29765,N_25696);
or UO_3358 (O_3358,N_28281,N_26574);
xor UO_3359 (O_3359,N_28500,N_27062);
nor UO_3360 (O_3360,N_28171,N_27606);
nand UO_3361 (O_3361,N_24961,N_28508);
nor UO_3362 (O_3362,N_28362,N_25773);
xor UO_3363 (O_3363,N_24120,N_29587);
or UO_3364 (O_3364,N_24641,N_25976);
nor UO_3365 (O_3365,N_27666,N_25673);
or UO_3366 (O_3366,N_27812,N_29451);
and UO_3367 (O_3367,N_28305,N_27579);
nand UO_3368 (O_3368,N_29652,N_24415);
nor UO_3369 (O_3369,N_27885,N_26519);
nand UO_3370 (O_3370,N_28058,N_26921);
or UO_3371 (O_3371,N_27020,N_26909);
nor UO_3372 (O_3372,N_25410,N_26968);
nor UO_3373 (O_3373,N_29618,N_24517);
xor UO_3374 (O_3374,N_29412,N_27262);
and UO_3375 (O_3375,N_24189,N_26261);
and UO_3376 (O_3376,N_24160,N_26574);
nand UO_3377 (O_3377,N_28782,N_29832);
nor UO_3378 (O_3378,N_25047,N_27176);
or UO_3379 (O_3379,N_29780,N_27554);
nand UO_3380 (O_3380,N_29790,N_29473);
xor UO_3381 (O_3381,N_27148,N_25640);
nor UO_3382 (O_3382,N_25333,N_24118);
xnor UO_3383 (O_3383,N_24714,N_27915);
nor UO_3384 (O_3384,N_24700,N_24540);
and UO_3385 (O_3385,N_25955,N_24869);
nor UO_3386 (O_3386,N_26794,N_26858);
xnor UO_3387 (O_3387,N_27214,N_26728);
xnor UO_3388 (O_3388,N_28871,N_24565);
nor UO_3389 (O_3389,N_25482,N_26838);
or UO_3390 (O_3390,N_26175,N_26274);
and UO_3391 (O_3391,N_26469,N_29198);
or UO_3392 (O_3392,N_29787,N_25791);
xor UO_3393 (O_3393,N_24273,N_28189);
and UO_3394 (O_3394,N_26407,N_25256);
and UO_3395 (O_3395,N_26830,N_27640);
nand UO_3396 (O_3396,N_29011,N_29286);
and UO_3397 (O_3397,N_27698,N_28994);
nand UO_3398 (O_3398,N_27553,N_27248);
nand UO_3399 (O_3399,N_26798,N_24070);
or UO_3400 (O_3400,N_27222,N_27952);
and UO_3401 (O_3401,N_24311,N_27665);
xor UO_3402 (O_3402,N_24018,N_24600);
xnor UO_3403 (O_3403,N_24104,N_28828);
or UO_3404 (O_3404,N_24390,N_29565);
or UO_3405 (O_3405,N_27174,N_26333);
and UO_3406 (O_3406,N_27698,N_29330);
nor UO_3407 (O_3407,N_28916,N_29625);
and UO_3408 (O_3408,N_29078,N_25871);
and UO_3409 (O_3409,N_25757,N_29947);
nor UO_3410 (O_3410,N_27922,N_29041);
or UO_3411 (O_3411,N_24587,N_29376);
nor UO_3412 (O_3412,N_28490,N_29080);
or UO_3413 (O_3413,N_28383,N_27168);
nand UO_3414 (O_3414,N_28734,N_26959);
and UO_3415 (O_3415,N_27606,N_27840);
xnor UO_3416 (O_3416,N_24107,N_25979);
xor UO_3417 (O_3417,N_27323,N_27824);
or UO_3418 (O_3418,N_27929,N_24352);
or UO_3419 (O_3419,N_26753,N_26501);
and UO_3420 (O_3420,N_25475,N_26808);
or UO_3421 (O_3421,N_24036,N_25911);
xor UO_3422 (O_3422,N_25221,N_29727);
or UO_3423 (O_3423,N_26291,N_24324);
xor UO_3424 (O_3424,N_26592,N_29462);
nand UO_3425 (O_3425,N_24976,N_26885);
nor UO_3426 (O_3426,N_27820,N_29560);
and UO_3427 (O_3427,N_28551,N_28185);
or UO_3428 (O_3428,N_26658,N_24180);
or UO_3429 (O_3429,N_25830,N_29375);
and UO_3430 (O_3430,N_24192,N_25185);
nor UO_3431 (O_3431,N_29154,N_29350);
or UO_3432 (O_3432,N_25516,N_25957);
or UO_3433 (O_3433,N_25239,N_29672);
or UO_3434 (O_3434,N_24877,N_26985);
and UO_3435 (O_3435,N_27818,N_25857);
xor UO_3436 (O_3436,N_25324,N_24692);
or UO_3437 (O_3437,N_28017,N_25829);
xnor UO_3438 (O_3438,N_25055,N_26971);
xor UO_3439 (O_3439,N_24968,N_28585);
or UO_3440 (O_3440,N_27084,N_25129);
nor UO_3441 (O_3441,N_28206,N_29677);
and UO_3442 (O_3442,N_28242,N_28526);
nor UO_3443 (O_3443,N_27551,N_25645);
nand UO_3444 (O_3444,N_26874,N_29804);
or UO_3445 (O_3445,N_25652,N_29525);
xnor UO_3446 (O_3446,N_28417,N_27892);
nor UO_3447 (O_3447,N_24349,N_29886);
and UO_3448 (O_3448,N_29556,N_28019);
or UO_3449 (O_3449,N_29083,N_28026);
nor UO_3450 (O_3450,N_29855,N_24690);
nor UO_3451 (O_3451,N_27048,N_28872);
nand UO_3452 (O_3452,N_26258,N_25291);
xor UO_3453 (O_3453,N_26153,N_29672);
and UO_3454 (O_3454,N_29180,N_29781);
nor UO_3455 (O_3455,N_24513,N_25868);
xor UO_3456 (O_3456,N_26198,N_27156);
and UO_3457 (O_3457,N_24510,N_25915);
nor UO_3458 (O_3458,N_25349,N_25940);
nand UO_3459 (O_3459,N_27801,N_26628);
and UO_3460 (O_3460,N_26414,N_28929);
xor UO_3461 (O_3461,N_27200,N_27315);
nor UO_3462 (O_3462,N_25043,N_29524);
or UO_3463 (O_3463,N_28262,N_29874);
nand UO_3464 (O_3464,N_29517,N_25125);
nand UO_3465 (O_3465,N_26488,N_29802);
and UO_3466 (O_3466,N_25038,N_28870);
or UO_3467 (O_3467,N_29289,N_25875);
nor UO_3468 (O_3468,N_29426,N_25058);
xor UO_3469 (O_3469,N_29303,N_24976);
xnor UO_3470 (O_3470,N_28377,N_24614);
nand UO_3471 (O_3471,N_25083,N_24661);
xnor UO_3472 (O_3472,N_29448,N_26017);
nand UO_3473 (O_3473,N_28043,N_27430);
nor UO_3474 (O_3474,N_28901,N_24911);
or UO_3475 (O_3475,N_26484,N_26971);
nand UO_3476 (O_3476,N_29242,N_27277);
and UO_3477 (O_3477,N_25677,N_24326);
and UO_3478 (O_3478,N_25041,N_27082);
xor UO_3479 (O_3479,N_24740,N_26455);
nor UO_3480 (O_3480,N_28840,N_24119);
xor UO_3481 (O_3481,N_27049,N_27034);
and UO_3482 (O_3482,N_27189,N_28082);
and UO_3483 (O_3483,N_27433,N_27444);
xor UO_3484 (O_3484,N_27718,N_24477);
nand UO_3485 (O_3485,N_24054,N_25045);
and UO_3486 (O_3486,N_29244,N_26916);
nor UO_3487 (O_3487,N_29081,N_26273);
and UO_3488 (O_3488,N_29642,N_28344);
nor UO_3489 (O_3489,N_25326,N_25504);
xnor UO_3490 (O_3490,N_24354,N_29637);
nand UO_3491 (O_3491,N_28152,N_26961);
nand UO_3492 (O_3492,N_28832,N_26682);
or UO_3493 (O_3493,N_24227,N_28769);
xor UO_3494 (O_3494,N_29833,N_25721);
nor UO_3495 (O_3495,N_28775,N_24261);
nor UO_3496 (O_3496,N_29206,N_25383);
or UO_3497 (O_3497,N_24168,N_25118);
nor UO_3498 (O_3498,N_28410,N_28547);
and UO_3499 (O_3499,N_24323,N_27307);
endmodule