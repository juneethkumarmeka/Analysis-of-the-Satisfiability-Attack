module basic_750_5000_1000_5_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_175,In_608);
xor U1 (N_1,In_579,In_462);
xor U2 (N_2,In_716,In_406);
or U3 (N_3,In_52,In_21);
nor U4 (N_4,In_152,In_90);
or U5 (N_5,In_454,In_495);
nand U6 (N_6,In_425,In_366);
nand U7 (N_7,In_459,In_563);
nand U8 (N_8,In_507,In_746);
or U9 (N_9,In_650,In_356);
nand U10 (N_10,In_196,In_566);
xnor U11 (N_11,In_157,In_497);
xnor U12 (N_12,In_538,In_150);
and U13 (N_13,In_231,In_270);
nor U14 (N_14,In_197,In_153);
and U15 (N_15,In_685,In_77);
or U16 (N_16,In_728,In_391);
and U17 (N_17,In_480,In_34);
or U18 (N_18,In_656,In_645);
and U19 (N_19,In_431,In_239);
nor U20 (N_20,In_542,In_596);
nand U21 (N_21,In_474,In_46);
and U22 (N_22,In_369,In_230);
nor U23 (N_23,In_419,In_570);
nor U24 (N_24,In_509,In_345);
and U25 (N_25,In_501,In_553);
nand U26 (N_26,In_211,In_300);
nor U27 (N_27,In_529,In_268);
or U28 (N_28,In_521,In_254);
nor U29 (N_29,In_56,In_400);
or U30 (N_30,In_636,In_149);
or U31 (N_31,In_25,In_232);
nand U32 (N_32,In_452,In_671);
nand U33 (N_33,In_591,In_110);
or U34 (N_34,In_496,In_238);
and U35 (N_35,In_629,In_445);
and U36 (N_36,In_7,In_535);
or U37 (N_37,In_304,In_5);
nand U38 (N_38,In_471,In_590);
nor U39 (N_39,In_35,In_381);
nor U40 (N_40,In_531,In_422);
or U41 (N_41,In_520,In_33);
nor U42 (N_42,In_528,In_460);
and U43 (N_43,In_14,In_205);
nand U44 (N_44,In_301,In_67);
nand U45 (N_45,In_715,In_255);
or U46 (N_46,In_470,In_24);
or U47 (N_47,In_588,In_720);
or U48 (N_48,In_198,In_360);
or U49 (N_49,In_731,In_286);
nand U50 (N_50,In_659,In_705);
or U51 (N_51,In_107,In_66);
nor U52 (N_52,In_556,In_517);
nand U53 (N_53,In_453,In_672);
nor U54 (N_54,In_287,In_281);
nor U55 (N_55,In_245,In_83);
xnor U56 (N_56,In_547,In_280);
and U57 (N_57,In_614,In_225);
or U58 (N_58,In_514,In_203);
or U59 (N_59,In_584,In_267);
nor U60 (N_60,In_616,In_694);
nor U61 (N_61,In_623,In_260);
xor U62 (N_62,In_54,In_108);
nand U63 (N_63,In_394,In_367);
or U64 (N_64,In_427,In_617);
or U65 (N_65,In_26,In_475);
and U66 (N_66,In_371,In_111);
or U67 (N_67,In_456,In_9);
or U68 (N_68,In_562,In_69);
nor U69 (N_69,In_45,In_607);
nor U70 (N_70,In_654,In_236);
nand U71 (N_71,In_76,In_147);
or U72 (N_72,In_8,In_493);
nand U73 (N_73,In_557,In_692);
or U74 (N_74,In_649,In_161);
nor U75 (N_75,In_707,In_122);
and U76 (N_76,In_540,In_183);
nor U77 (N_77,In_741,In_179);
and U78 (N_78,In_549,In_372);
or U79 (N_79,In_327,In_580);
and U80 (N_80,In_613,In_303);
and U81 (N_81,In_17,In_305);
and U82 (N_82,In_13,In_701);
or U83 (N_83,In_389,In_95);
nor U84 (N_84,In_710,In_133);
nor U85 (N_85,In_146,In_444);
nor U86 (N_86,In_703,In_120);
nor U87 (N_87,In_63,In_128);
or U88 (N_88,In_651,In_719);
or U89 (N_89,In_567,In_240);
nand U90 (N_90,In_58,In_555);
nand U91 (N_91,In_169,In_730);
and U92 (N_92,In_530,In_598);
nor U93 (N_93,In_484,In_693);
nor U94 (N_94,In_100,In_515);
and U95 (N_95,In_334,In_634);
nand U96 (N_96,In_278,In_355);
or U97 (N_97,In_505,In_660);
nand U98 (N_98,In_718,In_154);
nor U99 (N_99,In_177,In_439);
or U100 (N_100,In_626,In_575);
and U101 (N_101,In_510,In_408);
xor U102 (N_102,In_243,In_506);
or U103 (N_103,In_450,In_51);
nand U104 (N_104,In_134,In_62);
nand U105 (N_105,In_87,In_277);
xnor U106 (N_106,In_48,In_269);
and U107 (N_107,In_604,In_441);
nor U108 (N_108,In_461,In_415);
nor U109 (N_109,In_679,In_383);
nor U110 (N_110,In_47,In_544);
nand U111 (N_111,In_131,In_306);
or U112 (N_112,In_477,In_112);
nand U113 (N_113,In_215,In_190);
xor U114 (N_114,In_30,In_424);
and U115 (N_115,In_399,In_709);
nand U116 (N_116,In_683,In_57);
or U117 (N_117,In_195,In_740);
nor U118 (N_118,In_413,In_465);
xnor U119 (N_119,In_343,In_224);
nor U120 (N_120,In_294,In_658);
nor U121 (N_121,In_368,In_302);
xnor U122 (N_122,In_96,In_323);
and U123 (N_123,In_361,In_696);
and U124 (N_124,In_137,In_621);
or U125 (N_125,In_89,In_65);
nor U126 (N_126,In_226,In_677);
or U127 (N_127,In_583,In_353);
nand U128 (N_128,In_485,In_572);
xor U129 (N_129,In_235,In_148);
or U130 (N_130,In_274,In_324);
or U131 (N_131,In_565,In_129);
nand U132 (N_132,In_188,In_299);
and U133 (N_133,In_186,In_401);
nor U134 (N_134,In_712,In_700);
nand U135 (N_135,In_307,In_143);
and U136 (N_136,In_734,In_749);
or U137 (N_137,In_545,In_657);
or U138 (N_138,In_74,In_603);
nand U139 (N_139,In_136,In_392);
nor U140 (N_140,In_536,In_142);
nor U141 (N_141,In_443,In_352);
or U142 (N_142,In_378,In_99);
nor U143 (N_143,In_28,In_486);
and U144 (N_144,In_446,In_216);
or U145 (N_145,In_248,In_118);
nand U146 (N_146,In_331,In_407);
nor U147 (N_147,In_275,In_249);
nor U148 (N_148,In_676,In_180);
nor U149 (N_149,In_222,In_476);
or U150 (N_150,In_468,In_365);
and U151 (N_151,In_288,In_639);
or U152 (N_152,In_398,In_15);
nor U153 (N_153,In_346,In_606);
nor U154 (N_154,In_397,In_79);
nand U155 (N_155,In_500,In_519);
and U156 (N_156,In_194,In_404);
nand U157 (N_157,In_193,In_263);
and U158 (N_158,In_541,In_257);
nand U159 (N_159,In_729,In_674);
and U160 (N_160,In_589,In_289);
nor U161 (N_161,In_258,In_262);
nor U162 (N_162,In_627,In_440);
nor U163 (N_163,In_127,In_647);
xor U164 (N_164,In_185,In_247);
and U165 (N_165,In_502,In_246);
and U166 (N_166,In_576,In_335);
nand U167 (N_167,In_166,In_348);
or U168 (N_168,In_70,In_388);
nor U169 (N_169,In_457,In_312);
or U170 (N_170,In_373,In_410);
nor U171 (N_171,In_420,In_726);
and U172 (N_172,In_393,In_174);
and U173 (N_173,In_577,In_91);
nand U174 (N_174,In_336,In_681);
nand U175 (N_175,In_283,In_158);
nor U176 (N_176,In_81,In_537);
or U177 (N_177,In_375,In_554);
nand U178 (N_178,In_724,In_64);
nand U179 (N_179,In_582,In_578);
nand U180 (N_180,In_237,In_571);
xnor U181 (N_181,In_494,In_665);
nand U182 (N_182,In_295,In_98);
or U183 (N_183,In_581,In_736);
or U184 (N_184,In_738,In_702);
or U185 (N_185,In_344,In_272);
and U186 (N_186,In_244,In_0);
xor U187 (N_187,In_472,In_80);
and U188 (N_188,In_314,In_684);
nand U189 (N_189,In_744,In_722);
xnor U190 (N_190,In_503,In_455);
and U191 (N_191,In_653,In_691);
xnor U192 (N_192,In_159,In_414);
nor U193 (N_193,In_221,In_43);
and U194 (N_194,In_207,In_699);
nand U195 (N_195,In_178,In_527);
or U196 (N_196,In_273,In_139);
xor U197 (N_197,In_206,In_121);
nor U198 (N_198,In_347,In_560);
and U199 (N_199,In_745,In_594);
or U200 (N_200,In_214,In_362);
or U201 (N_201,In_191,In_643);
nand U202 (N_202,In_85,In_669);
and U203 (N_203,In_102,In_698);
and U204 (N_204,In_522,In_322);
nand U205 (N_205,In_310,In_619);
xor U206 (N_206,In_411,In_36);
nor U207 (N_207,In_330,In_370);
and U208 (N_208,In_640,In_39);
nand U209 (N_209,In_22,In_298);
and U210 (N_210,In_680,In_377);
and U211 (N_211,In_204,In_27);
nor U212 (N_212,In_668,In_417);
and U213 (N_213,In_104,In_747);
nand U214 (N_214,In_340,In_71);
xnor U215 (N_215,In_141,In_435);
nand U216 (N_216,In_721,In_635);
nor U217 (N_217,In_358,In_678);
nor U218 (N_218,In_597,In_548);
and U219 (N_219,In_297,In_11);
and U220 (N_220,In_708,In_176);
and U221 (N_221,In_126,In_227);
or U222 (N_222,In_124,In_717);
xnor U223 (N_223,In_184,In_428);
or U224 (N_224,In_610,In_88);
nand U225 (N_225,In_573,In_469);
nor U226 (N_226,In_130,In_292);
nand U227 (N_227,In_326,In_374);
nand U228 (N_228,In_516,In_97);
or U229 (N_229,In_84,In_385);
or U230 (N_230,In_316,In_50);
nor U231 (N_231,In_132,In_200);
xnor U232 (N_232,In_181,In_103);
or U233 (N_233,In_293,In_172);
nand U234 (N_234,In_585,In_402);
nand U235 (N_235,In_412,In_586);
xor U236 (N_236,In_479,In_686);
and U237 (N_237,In_119,In_713);
xnor U238 (N_238,In_363,In_201);
or U239 (N_239,In_72,In_689);
xor U240 (N_240,In_308,In_6);
nor U241 (N_241,In_382,In_376);
and U242 (N_242,In_223,In_504);
and U243 (N_243,In_395,In_449);
nand U244 (N_244,In_364,In_266);
nor U245 (N_245,In_115,In_209);
or U246 (N_246,In_637,In_41);
nor U247 (N_247,In_725,In_165);
nor U248 (N_248,In_727,In_135);
xor U249 (N_249,In_212,In_49);
or U250 (N_250,In_624,In_271);
and U251 (N_251,In_546,In_40);
xor U252 (N_252,In_279,In_426);
nand U253 (N_253,In_329,In_42);
and U254 (N_254,In_18,In_284);
nand U255 (N_255,In_220,In_673);
nor U256 (N_256,In_655,In_187);
and U257 (N_257,In_93,In_646);
nand U258 (N_258,In_4,In_574);
and U259 (N_259,In_379,In_265);
or U260 (N_260,In_202,In_276);
and U261 (N_261,In_290,In_78);
or U262 (N_262,In_662,In_61);
nor U263 (N_263,In_10,In_349);
and U264 (N_264,In_447,In_233);
xor U265 (N_265,In_38,In_44);
or U266 (N_266,In_113,In_687);
xor U267 (N_267,In_595,In_387);
and U268 (N_268,In_630,In_518);
nor U269 (N_269,In_442,In_632);
nand U270 (N_270,In_587,In_341);
or U271 (N_271,In_733,In_155);
or U272 (N_272,In_438,In_593);
nor U273 (N_273,In_667,In_320);
or U274 (N_274,In_511,In_605);
and U275 (N_275,In_86,In_32);
or U276 (N_276,In_430,In_105);
nand U277 (N_277,In_94,In_92);
or U278 (N_278,In_251,In_338);
and U279 (N_279,In_55,In_448);
or U280 (N_280,In_332,In_210);
nor U281 (N_281,In_140,In_473);
nor U282 (N_282,In_217,In_1);
nor U283 (N_283,In_380,In_524);
or U284 (N_284,In_481,In_483);
nand U285 (N_285,In_612,In_551);
nand U286 (N_286,In_688,In_592);
nand U287 (N_287,In_458,In_351);
and U288 (N_288,In_532,In_23);
or U289 (N_289,In_600,In_234);
and U290 (N_290,In_315,In_642);
and U291 (N_291,In_250,In_433);
or U292 (N_292,In_321,In_123);
or U293 (N_293,In_2,In_568);
xor U294 (N_294,In_464,In_218);
nand U295 (N_295,In_615,In_609);
xor U296 (N_296,In_421,In_666);
or U297 (N_297,In_489,In_282);
or U298 (N_298,In_523,In_116);
nor U299 (N_299,In_59,In_317);
and U300 (N_300,In_164,In_163);
and U301 (N_301,In_423,In_418);
nand U302 (N_302,In_313,In_436);
xnor U303 (N_303,In_539,In_342);
nand U304 (N_304,In_309,In_704);
or U305 (N_305,In_543,In_167);
nor U306 (N_306,In_697,In_339);
nor U307 (N_307,In_625,In_737);
nand U308 (N_308,In_396,In_559);
or U309 (N_309,In_525,In_467);
or U310 (N_310,In_242,In_618);
and U311 (N_311,In_735,In_558);
or U312 (N_312,In_602,In_82);
nand U313 (N_313,In_601,In_534);
or U314 (N_314,In_291,In_644);
nor U315 (N_315,In_695,In_409);
and U316 (N_316,In_73,In_611);
or U317 (N_317,In_264,In_106);
nor U318 (N_318,In_550,In_285);
and U319 (N_319,In_173,In_466);
or U320 (N_320,In_319,In_318);
or U321 (N_321,In_633,In_690);
nand U322 (N_322,In_569,In_125);
nor U323 (N_323,In_664,In_513);
or U324 (N_324,In_463,In_359);
and U325 (N_325,In_482,In_259);
nor U326 (N_326,In_739,In_512);
nand U327 (N_327,In_37,In_492);
nand U328 (N_328,In_3,In_138);
nand U329 (N_329,In_333,In_638);
or U330 (N_330,In_337,In_732);
and U331 (N_331,In_552,In_487);
and U332 (N_332,In_60,In_416);
nor U333 (N_333,In_357,In_682);
nor U334 (N_334,In_19,In_561);
and U335 (N_335,In_53,In_488);
or U336 (N_336,In_160,In_533);
nand U337 (N_337,In_328,In_661);
nand U338 (N_338,In_162,In_491);
and U339 (N_339,In_620,In_490);
xnor U340 (N_340,In_171,In_168);
or U341 (N_341,In_498,In_648);
or U342 (N_342,In_748,In_711);
or U343 (N_343,In_706,In_252);
and U344 (N_344,In_114,In_675);
xnor U345 (N_345,In_354,In_564);
nor U346 (N_346,In_499,In_403);
and U347 (N_347,In_743,In_156);
nor U348 (N_348,In_723,In_631);
xor U349 (N_349,In_101,In_16);
nor U350 (N_350,In_670,In_350);
nor U351 (N_351,In_151,In_229);
nand U352 (N_352,In_68,In_109);
xnor U353 (N_353,In_429,In_192);
and U354 (N_354,In_228,In_12);
and U355 (N_355,In_405,In_325);
nand U356 (N_356,In_628,In_208);
and U357 (N_357,In_478,In_145);
or U358 (N_358,In_182,In_256);
nand U359 (N_359,In_213,In_508);
or U360 (N_360,In_31,In_451);
nand U361 (N_361,In_241,In_29);
and U362 (N_362,In_219,In_386);
or U363 (N_363,In_170,In_296);
or U364 (N_364,In_390,In_117);
or U365 (N_365,In_599,In_434);
nand U366 (N_366,In_384,In_622);
and U367 (N_367,In_526,In_189);
nand U368 (N_368,In_75,In_652);
xor U369 (N_369,In_199,In_742);
nor U370 (N_370,In_714,In_261);
and U371 (N_371,In_663,In_311);
xnor U372 (N_372,In_437,In_253);
and U373 (N_373,In_641,In_20);
and U374 (N_374,In_144,In_432);
and U375 (N_375,In_345,In_716);
and U376 (N_376,In_674,In_646);
or U377 (N_377,In_636,In_683);
nor U378 (N_378,In_691,In_561);
or U379 (N_379,In_687,In_633);
nor U380 (N_380,In_23,In_531);
or U381 (N_381,In_134,In_653);
and U382 (N_382,In_135,In_73);
nor U383 (N_383,In_551,In_572);
or U384 (N_384,In_383,In_196);
nand U385 (N_385,In_255,In_514);
nor U386 (N_386,In_433,In_692);
or U387 (N_387,In_163,In_75);
nand U388 (N_388,In_424,In_172);
nand U389 (N_389,In_202,In_414);
nand U390 (N_390,In_357,In_439);
xor U391 (N_391,In_56,In_170);
nand U392 (N_392,In_167,In_82);
and U393 (N_393,In_397,In_578);
or U394 (N_394,In_515,In_485);
nor U395 (N_395,In_385,In_672);
nand U396 (N_396,In_92,In_51);
and U397 (N_397,In_0,In_549);
nand U398 (N_398,In_405,In_318);
nand U399 (N_399,In_457,In_121);
nand U400 (N_400,In_389,In_497);
or U401 (N_401,In_530,In_442);
nor U402 (N_402,In_368,In_540);
or U403 (N_403,In_303,In_209);
or U404 (N_404,In_50,In_119);
or U405 (N_405,In_692,In_681);
nand U406 (N_406,In_723,In_457);
and U407 (N_407,In_57,In_711);
nor U408 (N_408,In_480,In_434);
xor U409 (N_409,In_47,In_718);
and U410 (N_410,In_708,In_569);
and U411 (N_411,In_618,In_113);
nor U412 (N_412,In_175,In_115);
or U413 (N_413,In_53,In_390);
nor U414 (N_414,In_337,In_210);
xor U415 (N_415,In_175,In_422);
nor U416 (N_416,In_729,In_496);
nor U417 (N_417,In_90,In_617);
or U418 (N_418,In_237,In_387);
xnor U419 (N_419,In_539,In_565);
and U420 (N_420,In_500,In_0);
nor U421 (N_421,In_495,In_197);
and U422 (N_422,In_543,In_222);
xor U423 (N_423,In_203,In_547);
and U424 (N_424,In_338,In_413);
and U425 (N_425,In_464,In_568);
or U426 (N_426,In_535,In_624);
xor U427 (N_427,In_597,In_473);
xor U428 (N_428,In_109,In_99);
nand U429 (N_429,In_433,In_640);
and U430 (N_430,In_341,In_556);
or U431 (N_431,In_464,In_498);
nand U432 (N_432,In_385,In_387);
nand U433 (N_433,In_709,In_169);
and U434 (N_434,In_45,In_632);
or U435 (N_435,In_366,In_235);
nor U436 (N_436,In_680,In_59);
and U437 (N_437,In_446,In_509);
nor U438 (N_438,In_201,In_678);
xnor U439 (N_439,In_166,In_235);
or U440 (N_440,In_51,In_543);
and U441 (N_441,In_529,In_577);
nand U442 (N_442,In_202,In_525);
nor U443 (N_443,In_606,In_650);
or U444 (N_444,In_159,In_283);
nand U445 (N_445,In_592,In_62);
or U446 (N_446,In_443,In_318);
xnor U447 (N_447,In_134,In_388);
and U448 (N_448,In_80,In_171);
nor U449 (N_449,In_377,In_719);
or U450 (N_450,In_520,In_389);
or U451 (N_451,In_309,In_717);
and U452 (N_452,In_392,In_648);
and U453 (N_453,In_627,In_395);
nand U454 (N_454,In_345,In_393);
nor U455 (N_455,In_71,In_706);
nand U456 (N_456,In_188,In_671);
nor U457 (N_457,In_437,In_670);
and U458 (N_458,In_21,In_0);
or U459 (N_459,In_207,In_108);
or U460 (N_460,In_726,In_473);
xnor U461 (N_461,In_303,In_323);
nand U462 (N_462,In_487,In_18);
nand U463 (N_463,In_504,In_300);
nor U464 (N_464,In_27,In_202);
or U465 (N_465,In_28,In_512);
xor U466 (N_466,In_370,In_85);
nand U467 (N_467,In_446,In_170);
nand U468 (N_468,In_645,In_618);
and U469 (N_469,In_438,In_275);
and U470 (N_470,In_340,In_220);
xor U471 (N_471,In_84,In_359);
nor U472 (N_472,In_481,In_106);
or U473 (N_473,In_1,In_225);
nand U474 (N_474,In_376,In_172);
nand U475 (N_475,In_512,In_70);
nand U476 (N_476,In_82,In_324);
and U477 (N_477,In_194,In_644);
nand U478 (N_478,In_406,In_520);
nor U479 (N_479,In_646,In_208);
nand U480 (N_480,In_605,In_414);
or U481 (N_481,In_191,In_506);
nor U482 (N_482,In_367,In_438);
nor U483 (N_483,In_560,In_182);
nand U484 (N_484,In_168,In_438);
nand U485 (N_485,In_344,In_480);
xnor U486 (N_486,In_466,In_230);
nor U487 (N_487,In_529,In_198);
or U488 (N_488,In_591,In_50);
or U489 (N_489,In_325,In_482);
and U490 (N_490,In_307,In_560);
nor U491 (N_491,In_495,In_682);
and U492 (N_492,In_358,In_747);
nand U493 (N_493,In_166,In_423);
and U494 (N_494,In_52,In_554);
nor U495 (N_495,In_520,In_557);
or U496 (N_496,In_692,In_54);
nand U497 (N_497,In_611,In_308);
or U498 (N_498,In_743,In_275);
or U499 (N_499,In_629,In_330);
nor U500 (N_500,In_662,In_201);
and U501 (N_501,In_640,In_362);
or U502 (N_502,In_224,In_498);
nand U503 (N_503,In_693,In_54);
or U504 (N_504,In_56,In_77);
or U505 (N_505,In_390,In_45);
nor U506 (N_506,In_320,In_608);
or U507 (N_507,In_504,In_488);
nor U508 (N_508,In_356,In_549);
and U509 (N_509,In_569,In_431);
nor U510 (N_510,In_44,In_505);
nor U511 (N_511,In_293,In_269);
and U512 (N_512,In_529,In_394);
xnor U513 (N_513,In_251,In_666);
nand U514 (N_514,In_110,In_595);
or U515 (N_515,In_365,In_163);
nand U516 (N_516,In_297,In_107);
or U517 (N_517,In_62,In_612);
or U518 (N_518,In_617,In_485);
and U519 (N_519,In_129,In_298);
nor U520 (N_520,In_259,In_718);
or U521 (N_521,In_613,In_436);
and U522 (N_522,In_291,In_695);
and U523 (N_523,In_591,In_505);
nand U524 (N_524,In_299,In_75);
or U525 (N_525,In_445,In_42);
nor U526 (N_526,In_747,In_138);
nand U527 (N_527,In_354,In_395);
nor U528 (N_528,In_417,In_504);
and U529 (N_529,In_361,In_742);
and U530 (N_530,In_26,In_338);
nor U531 (N_531,In_177,In_283);
or U532 (N_532,In_550,In_466);
nand U533 (N_533,In_29,In_561);
nor U534 (N_534,In_742,In_450);
nand U535 (N_535,In_699,In_350);
and U536 (N_536,In_360,In_180);
nand U537 (N_537,In_205,In_438);
or U538 (N_538,In_112,In_255);
nor U539 (N_539,In_306,In_136);
or U540 (N_540,In_742,In_594);
and U541 (N_541,In_260,In_311);
and U542 (N_542,In_739,In_344);
nor U543 (N_543,In_10,In_410);
or U544 (N_544,In_429,In_609);
nor U545 (N_545,In_343,In_350);
or U546 (N_546,In_342,In_12);
nand U547 (N_547,In_534,In_322);
and U548 (N_548,In_112,In_622);
and U549 (N_549,In_250,In_690);
and U550 (N_550,In_478,In_530);
nor U551 (N_551,In_736,In_407);
and U552 (N_552,In_670,In_111);
or U553 (N_553,In_609,In_563);
nor U554 (N_554,In_636,In_439);
nand U555 (N_555,In_420,In_670);
xor U556 (N_556,In_485,In_283);
nor U557 (N_557,In_484,In_567);
nor U558 (N_558,In_236,In_622);
or U559 (N_559,In_661,In_420);
and U560 (N_560,In_428,In_324);
nor U561 (N_561,In_739,In_79);
or U562 (N_562,In_374,In_420);
nor U563 (N_563,In_521,In_600);
and U564 (N_564,In_137,In_468);
nor U565 (N_565,In_219,In_508);
and U566 (N_566,In_28,In_344);
nor U567 (N_567,In_575,In_468);
nor U568 (N_568,In_239,In_321);
xnor U569 (N_569,In_255,In_511);
xor U570 (N_570,In_445,In_447);
nor U571 (N_571,In_277,In_572);
nand U572 (N_572,In_115,In_256);
nor U573 (N_573,In_742,In_596);
nand U574 (N_574,In_284,In_612);
or U575 (N_575,In_263,In_514);
xnor U576 (N_576,In_314,In_526);
nand U577 (N_577,In_583,In_170);
nor U578 (N_578,In_619,In_448);
and U579 (N_579,In_615,In_332);
nand U580 (N_580,In_105,In_476);
xnor U581 (N_581,In_281,In_421);
or U582 (N_582,In_477,In_303);
nor U583 (N_583,In_267,In_348);
or U584 (N_584,In_111,In_297);
nor U585 (N_585,In_590,In_182);
or U586 (N_586,In_678,In_722);
nand U587 (N_587,In_205,In_1);
nand U588 (N_588,In_687,In_512);
and U589 (N_589,In_297,In_474);
nor U590 (N_590,In_381,In_496);
nand U591 (N_591,In_677,In_104);
xnor U592 (N_592,In_561,In_248);
nor U593 (N_593,In_554,In_34);
or U594 (N_594,In_741,In_206);
nand U595 (N_595,In_720,In_668);
or U596 (N_596,In_586,In_321);
nand U597 (N_597,In_381,In_437);
and U598 (N_598,In_401,In_485);
nor U599 (N_599,In_586,In_513);
nand U600 (N_600,In_517,In_427);
and U601 (N_601,In_125,In_289);
nand U602 (N_602,In_397,In_549);
nand U603 (N_603,In_368,In_525);
xnor U604 (N_604,In_138,In_202);
nand U605 (N_605,In_506,In_75);
nand U606 (N_606,In_323,In_576);
nand U607 (N_607,In_46,In_20);
or U608 (N_608,In_115,In_553);
and U609 (N_609,In_87,In_283);
or U610 (N_610,In_721,In_358);
and U611 (N_611,In_421,In_594);
or U612 (N_612,In_624,In_747);
and U613 (N_613,In_628,In_188);
and U614 (N_614,In_39,In_453);
nor U615 (N_615,In_664,In_45);
nand U616 (N_616,In_384,In_683);
xor U617 (N_617,In_736,In_66);
nor U618 (N_618,In_87,In_65);
nand U619 (N_619,In_710,In_192);
and U620 (N_620,In_525,In_495);
nand U621 (N_621,In_490,In_501);
nor U622 (N_622,In_159,In_540);
and U623 (N_623,In_506,In_370);
nand U624 (N_624,In_171,In_353);
and U625 (N_625,In_42,In_45);
nor U626 (N_626,In_40,In_107);
nand U627 (N_627,In_444,In_273);
and U628 (N_628,In_62,In_376);
or U629 (N_629,In_280,In_565);
nor U630 (N_630,In_328,In_270);
nand U631 (N_631,In_358,In_156);
or U632 (N_632,In_452,In_164);
or U633 (N_633,In_145,In_136);
or U634 (N_634,In_492,In_7);
nor U635 (N_635,In_566,In_230);
nand U636 (N_636,In_741,In_135);
or U637 (N_637,In_642,In_660);
nand U638 (N_638,In_623,In_651);
or U639 (N_639,In_358,In_198);
nor U640 (N_640,In_209,In_98);
or U641 (N_641,In_583,In_65);
nor U642 (N_642,In_358,In_144);
and U643 (N_643,In_330,In_671);
or U644 (N_644,In_324,In_465);
nor U645 (N_645,In_160,In_112);
or U646 (N_646,In_148,In_592);
xor U647 (N_647,In_532,In_133);
or U648 (N_648,In_747,In_43);
nand U649 (N_649,In_92,In_560);
and U650 (N_650,In_204,In_152);
xnor U651 (N_651,In_673,In_238);
nand U652 (N_652,In_69,In_284);
or U653 (N_653,In_472,In_741);
nor U654 (N_654,In_462,In_464);
xnor U655 (N_655,In_64,In_147);
nand U656 (N_656,In_537,In_443);
nand U657 (N_657,In_359,In_694);
or U658 (N_658,In_67,In_496);
and U659 (N_659,In_121,In_624);
or U660 (N_660,In_236,In_531);
or U661 (N_661,In_250,In_194);
nand U662 (N_662,In_36,In_340);
or U663 (N_663,In_26,In_302);
and U664 (N_664,In_101,In_421);
or U665 (N_665,In_192,In_250);
nor U666 (N_666,In_493,In_371);
or U667 (N_667,In_491,In_694);
and U668 (N_668,In_742,In_293);
or U669 (N_669,In_540,In_197);
and U670 (N_670,In_14,In_517);
nand U671 (N_671,In_383,In_370);
and U672 (N_672,In_513,In_556);
and U673 (N_673,In_89,In_498);
and U674 (N_674,In_237,In_677);
nand U675 (N_675,In_677,In_577);
nand U676 (N_676,In_367,In_460);
nand U677 (N_677,In_632,In_118);
nor U678 (N_678,In_5,In_138);
or U679 (N_679,In_689,In_591);
nand U680 (N_680,In_462,In_732);
or U681 (N_681,In_708,In_456);
and U682 (N_682,In_323,In_305);
nand U683 (N_683,In_606,In_78);
and U684 (N_684,In_82,In_462);
nor U685 (N_685,In_373,In_392);
nand U686 (N_686,In_93,In_187);
xnor U687 (N_687,In_233,In_374);
and U688 (N_688,In_60,In_241);
and U689 (N_689,In_554,In_104);
nand U690 (N_690,In_403,In_622);
nand U691 (N_691,In_632,In_385);
nand U692 (N_692,In_605,In_608);
nand U693 (N_693,In_447,In_81);
nand U694 (N_694,In_444,In_246);
nand U695 (N_695,In_569,In_370);
and U696 (N_696,In_662,In_529);
or U697 (N_697,In_678,In_707);
and U698 (N_698,In_693,In_490);
xor U699 (N_699,In_665,In_280);
xnor U700 (N_700,In_367,In_356);
or U701 (N_701,In_675,In_575);
xnor U702 (N_702,In_469,In_682);
or U703 (N_703,In_372,In_579);
or U704 (N_704,In_530,In_617);
nor U705 (N_705,In_245,In_333);
nor U706 (N_706,In_321,In_503);
nor U707 (N_707,In_411,In_164);
nand U708 (N_708,In_356,In_118);
nor U709 (N_709,In_535,In_405);
or U710 (N_710,In_524,In_421);
and U711 (N_711,In_374,In_334);
xor U712 (N_712,In_566,In_290);
and U713 (N_713,In_502,In_563);
nor U714 (N_714,In_695,In_81);
and U715 (N_715,In_700,In_402);
nor U716 (N_716,In_594,In_702);
nor U717 (N_717,In_552,In_352);
or U718 (N_718,In_505,In_203);
or U719 (N_719,In_528,In_135);
xor U720 (N_720,In_670,In_121);
nor U721 (N_721,In_229,In_230);
xor U722 (N_722,In_290,In_709);
nand U723 (N_723,In_678,In_534);
and U724 (N_724,In_392,In_88);
and U725 (N_725,In_673,In_303);
nand U726 (N_726,In_494,In_655);
nor U727 (N_727,In_555,In_513);
nor U728 (N_728,In_30,In_707);
nor U729 (N_729,In_636,In_698);
nand U730 (N_730,In_618,In_342);
xor U731 (N_731,In_116,In_126);
and U732 (N_732,In_691,In_602);
or U733 (N_733,In_730,In_157);
xnor U734 (N_734,In_174,In_432);
nand U735 (N_735,In_253,In_29);
and U736 (N_736,In_393,In_7);
nand U737 (N_737,In_236,In_687);
nor U738 (N_738,In_140,In_42);
and U739 (N_739,In_727,In_312);
and U740 (N_740,In_43,In_200);
nand U741 (N_741,In_696,In_426);
nand U742 (N_742,In_261,In_540);
and U743 (N_743,In_3,In_62);
nand U744 (N_744,In_511,In_219);
and U745 (N_745,In_40,In_153);
nor U746 (N_746,In_55,In_529);
and U747 (N_747,In_110,In_708);
or U748 (N_748,In_681,In_51);
or U749 (N_749,In_39,In_358);
nand U750 (N_750,In_230,In_270);
and U751 (N_751,In_484,In_11);
or U752 (N_752,In_64,In_131);
nand U753 (N_753,In_684,In_673);
and U754 (N_754,In_297,In_469);
nand U755 (N_755,In_0,In_453);
or U756 (N_756,In_438,In_729);
or U757 (N_757,In_54,In_740);
nand U758 (N_758,In_308,In_99);
or U759 (N_759,In_381,In_126);
and U760 (N_760,In_55,In_245);
or U761 (N_761,In_271,In_98);
nor U762 (N_762,In_317,In_94);
nor U763 (N_763,In_691,In_730);
nand U764 (N_764,In_382,In_691);
nor U765 (N_765,In_305,In_60);
and U766 (N_766,In_664,In_221);
nor U767 (N_767,In_564,In_29);
nand U768 (N_768,In_306,In_557);
and U769 (N_769,In_580,In_704);
nor U770 (N_770,In_651,In_499);
and U771 (N_771,In_686,In_115);
nor U772 (N_772,In_671,In_402);
nand U773 (N_773,In_230,In_536);
and U774 (N_774,In_443,In_39);
nand U775 (N_775,In_74,In_16);
and U776 (N_776,In_557,In_518);
nor U777 (N_777,In_369,In_106);
and U778 (N_778,In_244,In_701);
xnor U779 (N_779,In_419,In_537);
nand U780 (N_780,In_654,In_54);
nor U781 (N_781,In_78,In_417);
and U782 (N_782,In_195,In_56);
or U783 (N_783,In_397,In_34);
or U784 (N_784,In_260,In_127);
and U785 (N_785,In_440,In_694);
and U786 (N_786,In_183,In_720);
and U787 (N_787,In_329,In_540);
nand U788 (N_788,In_110,In_671);
or U789 (N_789,In_599,In_695);
nor U790 (N_790,In_738,In_202);
nand U791 (N_791,In_189,In_144);
nand U792 (N_792,In_705,In_632);
nor U793 (N_793,In_53,In_224);
or U794 (N_794,In_60,In_231);
nand U795 (N_795,In_626,In_666);
or U796 (N_796,In_192,In_513);
or U797 (N_797,In_244,In_553);
nor U798 (N_798,In_716,In_311);
or U799 (N_799,In_10,In_118);
xor U800 (N_800,In_123,In_254);
nor U801 (N_801,In_637,In_621);
or U802 (N_802,In_507,In_479);
and U803 (N_803,In_182,In_310);
and U804 (N_804,In_134,In_694);
xor U805 (N_805,In_159,In_362);
and U806 (N_806,In_274,In_293);
and U807 (N_807,In_173,In_568);
nand U808 (N_808,In_372,In_147);
or U809 (N_809,In_303,In_528);
or U810 (N_810,In_694,In_650);
nand U811 (N_811,In_470,In_723);
nand U812 (N_812,In_314,In_318);
nand U813 (N_813,In_586,In_409);
or U814 (N_814,In_416,In_424);
and U815 (N_815,In_63,In_328);
and U816 (N_816,In_360,In_176);
nor U817 (N_817,In_574,In_246);
nor U818 (N_818,In_446,In_724);
or U819 (N_819,In_397,In_369);
nor U820 (N_820,In_399,In_397);
nand U821 (N_821,In_730,In_357);
and U822 (N_822,In_674,In_135);
or U823 (N_823,In_717,In_715);
or U824 (N_824,In_626,In_371);
and U825 (N_825,In_703,In_495);
xor U826 (N_826,In_420,In_246);
nand U827 (N_827,In_81,In_173);
nor U828 (N_828,In_281,In_107);
or U829 (N_829,In_196,In_261);
and U830 (N_830,In_106,In_72);
nor U831 (N_831,In_188,In_167);
nand U832 (N_832,In_606,In_704);
nor U833 (N_833,In_43,In_595);
nand U834 (N_834,In_334,In_575);
nor U835 (N_835,In_164,In_465);
nor U836 (N_836,In_473,In_437);
nor U837 (N_837,In_200,In_621);
or U838 (N_838,In_157,In_245);
nor U839 (N_839,In_748,In_309);
nor U840 (N_840,In_479,In_302);
nor U841 (N_841,In_261,In_228);
and U842 (N_842,In_612,In_420);
xnor U843 (N_843,In_358,In_510);
and U844 (N_844,In_359,In_88);
nor U845 (N_845,In_446,In_82);
or U846 (N_846,In_320,In_377);
xnor U847 (N_847,In_93,In_680);
or U848 (N_848,In_697,In_592);
xnor U849 (N_849,In_735,In_749);
nand U850 (N_850,In_39,In_35);
nor U851 (N_851,In_656,In_88);
nor U852 (N_852,In_736,In_272);
nor U853 (N_853,In_702,In_627);
or U854 (N_854,In_56,In_51);
nand U855 (N_855,In_157,In_516);
and U856 (N_856,In_178,In_618);
or U857 (N_857,In_45,In_195);
nor U858 (N_858,In_379,In_158);
nor U859 (N_859,In_260,In_444);
or U860 (N_860,In_97,In_170);
or U861 (N_861,In_355,In_646);
nor U862 (N_862,In_705,In_306);
and U863 (N_863,In_240,In_297);
and U864 (N_864,In_645,In_544);
xor U865 (N_865,In_646,In_588);
nand U866 (N_866,In_483,In_182);
nor U867 (N_867,In_547,In_170);
and U868 (N_868,In_684,In_19);
and U869 (N_869,In_661,In_557);
and U870 (N_870,In_690,In_336);
and U871 (N_871,In_432,In_342);
nand U872 (N_872,In_42,In_262);
or U873 (N_873,In_487,In_235);
nor U874 (N_874,In_412,In_634);
or U875 (N_875,In_0,In_541);
nand U876 (N_876,In_675,In_552);
nor U877 (N_877,In_106,In_252);
and U878 (N_878,In_558,In_168);
or U879 (N_879,In_644,In_344);
and U880 (N_880,In_716,In_727);
or U881 (N_881,In_366,In_373);
nand U882 (N_882,In_235,In_382);
or U883 (N_883,In_81,In_550);
nor U884 (N_884,In_743,In_492);
nor U885 (N_885,In_25,In_617);
and U886 (N_886,In_579,In_115);
and U887 (N_887,In_92,In_290);
or U888 (N_888,In_101,In_562);
nor U889 (N_889,In_100,In_383);
and U890 (N_890,In_249,In_188);
or U891 (N_891,In_459,In_267);
and U892 (N_892,In_90,In_404);
nor U893 (N_893,In_352,In_215);
nor U894 (N_894,In_4,In_168);
and U895 (N_895,In_492,In_719);
nor U896 (N_896,In_637,In_405);
and U897 (N_897,In_564,In_365);
or U898 (N_898,In_592,In_644);
xnor U899 (N_899,In_145,In_530);
xor U900 (N_900,In_726,In_107);
nor U901 (N_901,In_673,In_585);
and U902 (N_902,In_635,In_409);
and U903 (N_903,In_461,In_288);
or U904 (N_904,In_387,In_608);
and U905 (N_905,In_622,In_368);
or U906 (N_906,In_28,In_541);
nor U907 (N_907,In_146,In_66);
and U908 (N_908,In_353,In_262);
nor U909 (N_909,In_630,In_99);
nor U910 (N_910,In_18,In_104);
nor U911 (N_911,In_656,In_708);
nand U912 (N_912,In_327,In_160);
or U913 (N_913,In_317,In_101);
nor U914 (N_914,In_731,In_423);
nand U915 (N_915,In_462,In_333);
xnor U916 (N_916,In_565,In_514);
nor U917 (N_917,In_705,In_432);
nand U918 (N_918,In_640,In_448);
nand U919 (N_919,In_741,In_624);
nor U920 (N_920,In_341,In_676);
and U921 (N_921,In_471,In_186);
nand U922 (N_922,In_250,In_697);
xnor U923 (N_923,In_721,In_380);
nand U924 (N_924,In_97,In_30);
nand U925 (N_925,In_458,In_678);
xor U926 (N_926,In_674,In_414);
xnor U927 (N_927,In_31,In_188);
or U928 (N_928,In_60,In_646);
or U929 (N_929,In_309,In_610);
and U930 (N_930,In_560,In_669);
nand U931 (N_931,In_287,In_208);
xnor U932 (N_932,In_643,In_507);
nor U933 (N_933,In_386,In_633);
nand U934 (N_934,In_151,In_313);
xnor U935 (N_935,In_419,In_611);
nor U936 (N_936,In_186,In_544);
nor U937 (N_937,In_285,In_545);
and U938 (N_938,In_259,In_588);
nor U939 (N_939,In_443,In_247);
and U940 (N_940,In_81,In_1);
or U941 (N_941,In_733,In_461);
nor U942 (N_942,In_277,In_745);
xor U943 (N_943,In_137,In_605);
nand U944 (N_944,In_102,In_501);
and U945 (N_945,In_272,In_570);
and U946 (N_946,In_3,In_544);
or U947 (N_947,In_518,In_331);
or U948 (N_948,In_520,In_594);
and U949 (N_949,In_149,In_334);
nand U950 (N_950,In_328,In_45);
and U951 (N_951,In_516,In_541);
nand U952 (N_952,In_85,In_735);
and U953 (N_953,In_379,In_319);
and U954 (N_954,In_684,In_539);
nand U955 (N_955,In_721,In_354);
and U956 (N_956,In_223,In_455);
and U957 (N_957,In_52,In_722);
xnor U958 (N_958,In_37,In_79);
and U959 (N_959,In_330,In_72);
and U960 (N_960,In_243,In_695);
or U961 (N_961,In_570,In_525);
and U962 (N_962,In_729,In_645);
nand U963 (N_963,In_163,In_604);
nor U964 (N_964,In_188,In_79);
or U965 (N_965,In_117,In_147);
and U966 (N_966,In_726,In_733);
nor U967 (N_967,In_650,In_680);
nor U968 (N_968,In_637,In_623);
nor U969 (N_969,In_584,In_512);
or U970 (N_970,In_420,In_430);
nand U971 (N_971,In_282,In_567);
or U972 (N_972,In_533,In_682);
nor U973 (N_973,In_363,In_86);
and U974 (N_974,In_630,In_510);
nand U975 (N_975,In_564,In_687);
nand U976 (N_976,In_740,In_668);
nand U977 (N_977,In_496,In_679);
nor U978 (N_978,In_34,In_393);
and U979 (N_979,In_19,In_114);
nor U980 (N_980,In_651,In_52);
nand U981 (N_981,In_704,In_556);
or U982 (N_982,In_158,In_483);
nand U983 (N_983,In_289,In_680);
nor U984 (N_984,In_229,In_685);
nand U985 (N_985,In_229,In_219);
nand U986 (N_986,In_569,In_64);
or U987 (N_987,In_331,In_120);
and U988 (N_988,In_738,In_330);
nor U989 (N_989,In_349,In_604);
or U990 (N_990,In_18,In_163);
and U991 (N_991,In_214,In_176);
and U992 (N_992,In_309,In_333);
xor U993 (N_993,In_147,In_9);
xnor U994 (N_994,In_729,In_300);
and U995 (N_995,In_72,In_646);
or U996 (N_996,In_247,In_510);
nor U997 (N_997,In_29,In_395);
nand U998 (N_998,In_130,In_684);
or U999 (N_999,In_680,In_599);
nor U1000 (N_1000,N_2,N_632);
nand U1001 (N_1001,N_569,N_488);
nor U1002 (N_1002,N_521,N_34);
and U1003 (N_1003,N_360,N_161);
and U1004 (N_1004,N_480,N_247);
and U1005 (N_1005,N_182,N_795);
and U1006 (N_1006,N_841,N_450);
and U1007 (N_1007,N_53,N_503);
xor U1008 (N_1008,N_747,N_297);
and U1009 (N_1009,N_60,N_740);
nor U1010 (N_1010,N_773,N_870);
nor U1011 (N_1011,N_261,N_669);
and U1012 (N_1012,N_670,N_411);
nand U1013 (N_1013,N_915,N_932);
nor U1014 (N_1014,N_304,N_666);
nand U1015 (N_1015,N_933,N_968);
and U1016 (N_1016,N_995,N_487);
nor U1017 (N_1017,N_862,N_241);
or U1018 (N_1018,N_484,N_931);
or U1019 (N_1019,N_680,N_955);
nand U1020 (N_1020,N_463,N_86);
and U1021 (N_1021,N_930,N_564);
and U1022 (N_1022,N_17,N_949);
nor U1023 (N_1023,N_965,N_597);
nor U1024 (N_1024,N_8,N_687);
or U1025 (N_1025,N_836,N_539);
and U1026 (N_1026,N_631,N_111);
or U1027 (N_1027,N_115,N_353);
or U1028 (N_1028,N_603,N_784);
or U1029 (N_1029,N_529,N_978);
and U1030 (N_1030,N_590,N_122);
nand U1031 (N_1031,N_81,N_894);
and U1032 (N_1032,N_377,N_82);
nor U1033 (N_1033,N_490,N_306);
or U1034 (N_1034,N_725,N_544);
and U1035 (N_1035,N_628,N_924);
and U1036 (N_1036,N_741,N_589);
nor U1037 (N_1037,N_758,N_262);
nand U1038 (N_1038,N_872,N_658);
or U1039 (N_1039,N_882,N_588);
nor U1040 (N_1040,N_259,N_593);
nor U1041 (N_1041,N_971,N_433);
nor U1042 (N_1042,N_298,N_394);
and U1043 (N_1043,N_289,N_76);
nor U1044 (N_1044,N_581,N_614);
nor U1045 (N_1045,N_726,N_23);
nand U1046 (N_1046,N_660,N_234);
xnor U1047 (N_1047,N_209,N_442);
nand U1048 (N_1048,N_876,N_422);
nand U1049 (N_1049,N_63,N_87);
nor U1050 (N_1050,N_158,N_623);
and U1051 (N_1051,N_154,N_483);
nor U1052 (N_1052,N_399,N_721);
nor U1053 (N_1053,N_429,N_390);
and U1054 (N_1054,N_333,N_130);
and U1055 (N_1055,N_796,N_938);
and U1056 (N_1056,N_587,N_4);
or U1057 (N_1057,N_155,N_681);
or U1058 (N_1058,N_863,N_541);
and U1059 (N_1059,N_54,N_743);
or U1060 (N_1060,N_120,N_799);
and U1061 (N_1061,N_129,N_214);
nand U1062 (N_1062,N_531,N_465);
or U1063 (N_1063,N_400,N_185);
and U1064 (N_1064,N_170,N_676);
and U1065 (N_1065,N_361,N_335);
nor U1066 (N_1066,N_272,N_626);
nor U1067 (N_1067,N_838,N_921);
nand U1068 (N_1068,N_640,N_139);
and U1069 (N_1069,N_816,N_576);
nor U1070 (N_1070,N_926,N_582);
and U1071 (N_1071,N_156,N_16);
nor U1072 (N_1072,N_98,N_338);
nor U1073 (N_1073,N_489,N_874);
nand U1074 (N_1074,N_309,N_387);
or U1075 (N_1075,N_523,N_157);
nor U1076 (N_1076,N_977,N_513);
or U1077 (N_1077,N_116,N_555);
nor U1078 (N_1078,N_35,N_705);
nand U1079 (N_1079,N_595,N_347);
or U1080 (N_1080,N_211,N_601);
nand U1081 (N_1081,N_898,N_786);
nor U1082 (N_1082,N_510,N_383);
nand U1083 (N_1083,N_195,N_800);
or U1084 (N_1084,N_787,N_303);
nor U1085 (N_1085,N_911,N_388);
nor U1086 (N_1086,N_431,N_11);
nand U1087 (N_1087,N_830,N_228);
and U1088 (N_1088,N_985,N_964);
nor U1089 (N_1089,N_177,N_811);
xnor U1090 (N_1090,N_495,N_914);
or U1091 (N_1091,N_236,N_724);
nor U1092 (N_1092,N_918,N_763);
nand U1093 (N_1093,N_974,N_29);
xor U1094 (N_1094,N_118,N_927);
nor U1095 (N_1095,N_697,N_814);
and U1096 (N_1096,N_641,N_448);
and U1097 (N_1097,N_615,N_672);
nand U1098 (N_1098,N_67,N_493);
xor U1099 (N_1099,N_50,N_172);
nand U1100 (N_1100,N_80,N_37);
or U1101 (N_1101,N_485,N_551);
and U1102 (N_1102,N_913,N_861);
nand U1103 (N_1103,N_679,N_412);
or U1104 (N_1104,N_423,N_25);
or U1105 (N_1105,N_886,N_406);
nor U1106 (N_1106,N_871,N_478);
and U1107 (N_1107,N_382,N_56);
nand U1108 (N_1108,N_415,N_884);
nor U1109 (N_1109,N_829,N_418);
and U1110 (N_1110,N_230,N_526);
or U1111 (N_1111,N_878,N_109);
nor U1112 (N_1112,N_849,N_84);
nor U1113 (N_1113,N_151,N_408);
nor U1114 (N_1114,N_584,N_255);
nand U1115 (N_1115,N_941,N_976);
or U1116 (N_1116,N_100,N_742);
and U1117 (N_1117,N_516,N_966);
nor U1118 (N_1118,N_421,N_290);
nor U1119 (N_1119,N_715,N_344);
nand U1120 (N_1120,N_504,N_745);
nand U1121 (N_1121,N_835,N_245);
or U1122 (N_1122,N_103,N_983);
and U1123 (N_1123,N_123,N_470);
nor U1124 (N_1124,N_690,N_179);
or U1125 (N_1125,N_622,N_780);
xnor U1126 (N_1126,N_43,N_206);
nand U1127 (N_1127,N_253,N_356);
and U1128 (N_1128,N_507,N_282);
and U1129 (N_1129,N_216,N_193);
and U1130 (N_1130,N_580,N_712);
and U1131 (N_1131,N_358,N_897);
and U1132 (N_1132,N_919,N_770);
nor U1133 (N_1133,N_646,N_973);
or U1134 (N_1134,N_847,N_311);
nand U1135 (N_1135,N_858,N_577);
xnor U1136 (N_1136,N_368,N_227);
nor U1137 (N_1137,N_165,N_611);
nor U1138 (N_1138,N_686,N_126);
and U1139 (N_1139,N_990,N_895);
nand U1140 (N_1140,N_354,N_890);
or U1141 (N_1141,N_912,N_530);
or U1142 (N_1142,N_349,N_393);
and U1143 (N_1143,N_567,N_496);
nor U1144 (N_1144,N_506,N_980);
and U1145 (N_1145,N_152,N_416);
and U1146 (N_1146,N_452,N_425);
and U1147 (N_1147,N_27,N_583);
xor U1148 (N_1148,N_99,N_307);
or U1149 (N_1149,N_762,N_559);
or U1150 (N_1150,N_554,N_606);
and U1151 (N_1151,N_637,N_944);
nand U1152 (N_1152,N_337,N_128);
nand U1153 (N_1153,N_322,N_198);
nand U1154 (N_1154,N_843,N_839);
or U1155 (N_1155,N_119,N_385);
nor U1156 (N_1156,N_899,N_239);
and U1157 (N_1157,N_929,N_834);
xnor U1158 (N_1158,N_557,N_420);
and U1159 (N_1159,N_533,N_808);
nand U1160 (N_1160,N_859,N_407);
xnor U1161 (N_1161,N_276,N_534);
nand U1162 (N_1162,N_437,N_466);
or U1163 (N_1163,N_376,N_246);
or U1164 (N_1164,N_620,N_95);
and U1165 (N_1165,N_879,N_864);
and U1166 (N_1166,N_928,N_956);
and U1167 (N_1167,N_194,N_815);
and U1168 (N_1168,N_362,N_730);
xnor U1169 (N_1169,N_210,N_468);
nor U1170 (N_1170,N_942,N_826);
nor U1171 (N_1171,N_969,N_136);
nand U1172 (N_1172,N_867,N_267);
nand U1173 (N_1173,N_30,N_243);
nor U1174 (N_1174,N_249,N_852);
and U1175 (N_1175,N_453,N_375);
nand U1176 (N_1176,N_21,N_695);
and U1177 (N_1177,N_204,N_438);
nand U1178 (N_1178,N_748,N_674);
or U1179 (N_1179,N_779,N_134);
nor U1180 (N_1180,N_117,N_947);
nor U1181 (N_1181,N_51,N_305);
nand U1182 (N_1182,N_760,N_265);
or U1183 (N_1183,N_939,N_909);
and U1184 (N_1184,N_698,N_288);
xnor U1185 (N_1185,N_612,N_877);
or U1186 (N_1186,N_967,N_473);
and U1187 (N_1187,N_316,N_600);
or U1188 (N_1188,N_471,N_240);
nor U1189 (N_1189,N_367,N_945);
or U1190 (N_1190,N_527,N_553);
and U1191 (N_1191,N_732,N_220);
nor U1192 (N_1192,N_853,N_958);
or U1193 (N_1193,N_295,N_64);
nand U1194 (N_1194,N_410,N_824);
nor U1195 (N_1195,N_112,N_657);
or U1196 (N_1196,N_97,N_456);
xor U1197 (N_1197,N_723,N_47);
or U1198 (N_1198,N_906,N_998);
nand U1199 (N_1199,N_270,N_371);
nor U1200 (N_1200,N_359,N_801);
xnor U1201 (N_1201,N_684,N_910);
nor U1202 (N_1202,N_443,N_166);
xor U1203 (N_1203,N_634,N_257);
or U1204 (N_1204,N_761,N_6);
nand U1205 (N_1205,N_644,N_201);
xor U1206 (N_1206,N_819,N_296);
nand U1207 (N_1207,N_92,N_737);
or U1208 (N_1208,N_266,N_391);
nand U1209 (N_1209,N_192,N_806);
xnor U1210 (N_1210,N_324,N_24);
or U1211 (N_1211,N_750,N_778);
nor U1212 (N_1212,N_792,N_444);
and U1213 (N_1213,N_202,N_685);
nor U1214 (N_1214,N_341,N_759);
nor U1215 (N_1215,N_619,N_844);
nand U1216 (N_1216,N_804,N_823);
and U1217 (N_1217,N_273,N_302);
nor U1218 (N_1218,N_275,N_738);
or U1219 (N_1219,N_617,N_153);
or U1220 (N_1220,N_217,N_548);
nand U1221 (N_1221,N_701,N_511);
xor U1222 (N_1222,N_960,N_163);
nand U1223 (N_1223,N_774,N_52);
or U1224 (N_1224,N_594,N_552);
nand U1225 (N_1225,N_613,N_293);
or U1226 (N_1226,N_714,N_868);
and U1227 (N_1227,N_866,N_661);
nand U1228 (N_1228,N_363,N_260);
and U1229 (N_1229,N_954,N_89);
nor U1230 (N_1230,N_491,N_809);
nor U1231 (N_1231,N_268,N_310);
and U1232 (N_1232,N_769,N_467);
nand U1233 (N_1233,N_219,N_566);
xor U1234 (N_1234,N_199,N_332);
and U1235 (N_1235,N_596,N_540);
or U1236 (N_1236,N_9,N_428);
and U1237 (N_1237,N_475,N_215);
xnor U1238 (N_1238,N_846,N_916);
nand U1239 (N_1239,N_55,N_319);
and U1240 (N_1240,N_820,N_384);
nor U1241 (N_1241,N_851,N_765);
and U1242 (N_1242,N_148,N_213);
nand U1243 (N_1243,N_900,N_401);
or U1244 (N_1244,N_574,N_678);
and U1245 (N_1245,N_604,N_258);
nor U1246 (N_1246,N_934,N_183);
nor U1247 (N_1247,N_91,N_190);
xnor U1248 (N_1248,N_984,N_951);
xnor U1249 (N_1249,N_147,N_515);
nand U1250 (N_1250,N_405,N_875);
nand U1251 (N_1251,N_789,N_563);
nor U1252 (N_1252,N_937,N_850);
nor U1253 (N_1253,N_682,N_396);
and U1254 (N_1254,N_430,N_517);
nor U1255 (N_1255,N_378,N_469);
xor U1256 (N_1256,N_39,N_284);
and U1257 (N_1257,N_345,N_226);
or U1258 (N_1258,N_776,N_83);
or U1259 (N_1259,N_535,N_212);
nand U1260 (N_1260,N_197,N_72);
or U1261 (N_1261,N_790,N_221);
nor U1262 (N_1262,N_766,N_164);
and U1263 (N_1263,N_102,N_48);
and U1264 (N_1264,N_710,N_188);
nor U1265 (N_1265,N_69,N_627);
or U1266 (N_1266,N_281,N_231);
and U1267 (N_1267,N_610,N_373);
nand U1268 (N_1268,N_381,N_696);
nor U1269 (N_1269,N_328,N_413);
nand U1270 (N_1270,N_549,N_963);
xnor U1271 (N_1271,N_315,N_218);
and U1272 (N_1272,N_739,N_271);
nor U1273 (N_1273,N_318,N_832);
xnor U1274 (N_1274,N_15,N_274);
or U1275 (N_1275,N_108,N_114);
nor U1276 (N_1276,N_720,N_896);
or U1277 (N_1277,N_520,N_543);
nand U1278 (N_1278,N_427,N_837);
and U1279 (N_1279,N_810,N_744);
xor U1280 (N_1280,N_477,N_751);
or U1281 (N_1281,N_570,N_472);
nand U1282 (N_1282,N_462,N_975);
nor U1283 (N_1283,N_825,N_326);
nor U1284 (N_1284,N_336,N_334);
nand U1285 (N_1285,N_145,N_793);
nand U1286 (N_1286,N_424,N_280);
or U1287 (N_1287,N_350,N_77);
or U1288 (N_1288,N_981,N_142);
nand U1289 (N_1289,N_831,N_550);
xor U1290 (N_1290,N_512,N_772);
nand U1291 (N_1291,N_633,N_364);
or U1292 (N_1292,N_970,N_572);
nand U1293 (N_1293,N_591,N_460);
and U1294 (N_1294,N_12,N_66);
and U1295 (N_1295,N_88,N_771);
nor U1296 (N_1296,N_5,N_323);
nor U1297 (N_1297,N_486,N_536);
nand U1298 (N_1298,N_609,N_673);
and U1299 (N_1299,N_372,N_149);
and U1300 (N_1300,N_713,N_414);
nor U1301 (N_1301,N_854,N_439);
nand U1302 (N_1302,N_251,N_175);
nor U1303 (N_1303,N_936,N_464);
nand U1304 (N_1304,N_294,N_41);
nor U1305 (N_1305,N_224,N_665);
nor U1306 (N_1306,N_287,N_822);
or U1307 (N_1307,N_561,N_65);
xnor U1308 (N_1308,N_888,N_893);
nor U1309 (N_1309,N_313,N_250);
and U1310 (N_1310,N_651,N_370);
nor U1311 (N_1311,N_707,N_575);
nand U1312 (N_1312,N_683,N_321);
nor U1313 (N_1313,N_45,N_263);
nand U1314 (N_1314,N_671,N_101);
nor U1315 (N_1315,N_432,N_991);
nor U1316 (N_1316,N_106,N_812);
and U1317 (N_1317,N_920,N_445);
or U1318 (N_1318,N_200,N_621);
nand U1319 (N_1319,N_827,N_805);
nor U1320 (N_1320,N_127,N_178);
or U1321 (N_1321,N_592,N_833);
nand U1322 (N_1322,N_719,N_18);
xnor U1323 (N_1323,N_988,N_571);
or U1324 (N_1324,N_755,N_994);
nand U1325 (N_1325,N_568,N_62);
or U1326 (N_1326,N_892,N_386);
xor U1327 (N_1327,N_642,N_923);
and U1328 (N_1328,N_279,N_379);
nand U1329 (N_1329,N_499,N_777);
xor U1330 (N_1330,N_693,N_317);
and U1331 (N_1331,N_500,N_855);
and U1332 (N_1332,N_208,N_889);
and U1333 (N_1333,N_643,N_180);
and U1334 (N_1334,N_61,N_143);
and U1335 (N_1335,N_653,N_494);
and U1336 (N_1336,N_135,N_229);
nand U1337 (N_1337,N_299,N_881);
xor U1338 (N_1338,N_817,N_74);
or U1339 (N_1339,N_922,N_668);
nor U1340 (N_1340,N_320,N_982);
and U1341 (N_1341,N_972,N_946);
or U1342 (N_1342,N_343,N_402);
or U1343 (N_1343,N_70,N_33);
nand U1344 (N_1344,N_753,N_395);
nor U1345 (N_1345,N_121,N_357);
or U1346 (N_1346,N_264,N_254);
nand U1347 (N_1347,N_524,N_222);
and U1348 (N_1348,N_542,N_798);
and U1349 (N_1349,N_807,N_556);
nand U1350 (N_1350,N_578,N_840);
nand U1351 (N_1351,N_191,N_441);
and U1352 (N_1352,N_174,N_40);
or U1353 (N_1353,N_959,N_140);
nor U1354 (N_1354,N_461,N_797);
nor U1355 (N_1355,N_447,N_256);
nor U1356 (N_1356,N_625,N_857);
and U1357 (N_1357,N_398,N_419);
or U1358 (N_1358,N_308,N_706);
or U1359 (N_1359,N_986,N_953);
and U1360 (N_1360,N_546,N_505);
nand U1361 (N_1361,N_436,N_821);
nand U1362 (N_1362,N_689,N_525);
nor U1363 (N_1363,N_342,N_252);
and U1364 (N_1364,N_891,N_278);
or U1365 (N_1365,N_699,N_781);
nand U1366 (N_1366,N_989,N_996);
or U1367 (N_1367,N_736,N_374);
and U1368 (N_1368,N_292,N_187);
or U1369 (N_1369,N_537,N_629);
or U1370 (N_1370,N_46,N_788);
or U1371 (N_1371,N_365,N_655);
or U1372 (N_1372,N_901,N_708);
nor U1373 (N_1373,N_688,N_286);
and U1374 (N_1374,N_325,N_173);
xnor U1375 (N_1375,N_746,N_189);
nand U1376 (N_1376,N_474,N_141);
nand U1377 (N_1377,N_79,N_44);
xor U1378 (N_1378,N_560,N_403);
or U1379 (N_1379,N_664,N_94);
nand U1380 (N_1380,N_987,N_691);
nand U1381 (N_1381,N_454,N_476);
and U1382 (N_1382,N_828,N_20);
nand U1383 (N_1383,N_301,N_205);
nor U1384 (N_1384,N_32,N_481);
and U1385 (N_1385,N_501,N_355);
nand U1386 (N_1386,N_925,N_950);
nor U1387 (N_1387,N_242,N_75);
nor U1388 (N_1388,N_283,N_171);
nand U1389 (N_1389,N_733,N_366);
and U1390 (N_1390,N_782,N_1);
or U1391 (N_1391,N_734,N_107);
or U1392 (N_1392,N_314,N_348);
xor U1393 (N_1393,N_562,N_482);
or U1394 (N_1394,N_785,N_993);
and U1395 (N_1395,N_729,N_608);
or U1396 (N_1396,N_42,N_794);
or U1397 (N_1397,N_168,N_113);
and U1398 (N_1398,N_508,N_137);
or U1399 (N_1399,N_3,N_639);
nand U1400 (N_1400,N_13,N_0);
or U1401 (N_1401,N_14,N_331);
xor U1402 (N_1402,N_943,N_150);
nor U1403 (N_1403,N_38,N_196);
and U1404 (N_1404,N_455,N_749);
xnor U1405 (N_1405,N_409,N_392);
or U1406 (N_1406,N_885,N_248);
nor U1407 (N_1407,N_186,N_397);
nand U1408 (N_1408,N_767,N_19);
and U1409 (N_1409,N_96,N_160);
nor U1410 (N_1410,N_652,N_791);
nor U1411 (N_1411,N_694,N_638);
or U1412 (N_1412,N_110,N_514);
and U1413 (N_1413,N_607,N_908);
nor U1414 (N_1414,N_59,N_404);
nor U1415 (N_1415,N_545,N_579);
nand U1416 (N_1416,N_232,N_235);
or U1417 (N_1417,N_667,N_848);
or U1418 (N_1418,N_647,N_756);
and U1419 (N_1419,N_167,N_434);
nand U1420 (N_1420,N_71,N_340);
nand U1421 (N_1421,N_327,N_702);
nor U1422 (N_1422,N_602,N_869);
and U1423 (N_1423,N_764,N_865);
nor U1424 (N_1424,N_184,N_711);
xor U1425 (N_1425,N_532,N_451);
and U1426 (N_1426,N_7,N_479);
nor U1427 (N_1427,N_624,N_440);
nor U1428 (N_1428,N_775,N_692);
and U1429 (N_1429,N_104,N_459);
and U1430 (N_1430,N_28,N_300);
nand U1431 (N_1431,N_917,N_961);
or U1432 (N_1432,N_144,N_49);
nor U1433 (N_1433,N_146,N_518);
or U1434 (N_1434,N_645,N_58);
or U1435 (N_1435,N_757,N_352);
and U1436 (N_1436,N_31,N_329);
or U1437 (N_1437,N_880,N_457);
nor U1438 (N_1438,N_803,N_57);
and U1439 (N_1439,N_717,N_346);
or U1440 (N_1440,N_519,N_999);
nor U1441 (N_1441,N_635,N_538);
or U1442 (N_1442,N_905,N_818);
or U1443 (N_1443,N_903,N_573);
or U1444 (N_1444,N_36,N_649);
nand U1445 (N_1445,N_138,N_169);
or U1446 (N_1446,N_93,N_585);
and U1447 (N_1447,N_731,N_856);
nor U1448 (N_1448,N_845,N_547);
nand U1449 (N_1449,N_22,N_716);
and U1450 (N_1450,N_449,N_599);
xnor U1451 (N_1451,N_887,N_813);
and U1452 (N_1452,N_718,N_426);
nor U1453 (N_1453,N_389,N_904);
nor U1454 (N_1454,N_330,N_997);
nand U1455 (N_1455,N_417,N_233);
and U1456 (N_1456,N_105,N_957);
or U1457 (N_1457,N_558,N_312);
nor U1458 (N_1458,N_238,N_446);
or U1459 (N_1459,N_78,N_277);
and U1460 (N_1460,N_802,N_90);
and U1461 (N_1461,N_269,N_616);
nand U1462 (N_1462,N_73,N_992);
or U1463 (N_1463,N_703,N_709);
and U1464 (N_1464,N_948,N_598);
nand U1465 (N_1465,N_124,N_509);
nor U1466 (N_1466,N_618,N_162);
nor U1467 (N_1467,N_940,N_502);
or U1468 (N_1468,N_704,N_605);
xnor U1469 (N_1469,N_979,N_962);
nand U1470 (N_1470,N_244,N_369);
nor U1471 (N_1471,N_339,N_636);
xor U1472 (N_1472,N_902,N_656);
and U1473 (N_1473,N_663,N_132);
nand U1474 (N_1474,N_727,N_181);
and U1475 (N_1475,N_68,N_700);
or U1476 (N_1476,N_203,N_26);
or U1477 (N_1477,N_176,N_883);
nor U1478 (N_1478,N_492,N_728);
nor U1479 (N_1479,N_752,N_85);
nand U1480 (N_1480,N_522,N_10);
nor U1481 (N_1481,N_662,N_435);
nand U1482 (N_1482,N_285,N_225);
nor U1483 (N_1483,N_735,N_159);
nor U1484 (N_1484,N_654,N_754);
nor U1485 (N_1485,N_458,N_291);
nand U1486 (N_1486,N_565,N_659);
nor U1487 (N_1487,N_133,N_952);
or U1488 (N_1488,N_648,N_783);
nand U1489 (N_1489,N_860,N_223);
nand U1490 (N_1490,N_907,N_935);
nor U1491 (N_1491,N_237,N_675);
or U1492 (N_1492,N_125,N_650);
nand U1493 (N_1493,N_768,N_207);
nor U1494 (N_1494,N_528,N_351);
or U1495 (N_1495,N_586,N_722);
nor U1496 (N_1496,N_842,N_131);
nor U1497 (N_1497,N_497,N_677);
or U1498 (N_1498,N_873,N_630);
nor U1499 (N_1499,N_380,N_498);
and U1500 (N_1500,N_798,N_474);
and U1501 (N_1501,N_898,N_224);
and U1502 (N_1502,N_187,N_579);
nand U1503 (N_1503,N_519,N_99);
or U1504 (N_1504,N_538,N_528);
and U1505 (N_1505,N_308,N_700);
and U1506 (N_1506,N_382,N_25);
nor U1507 (N_1507,N_277,N_802);
or U1508 (N_1508,N_751,N_855);
xnor U1509 (N_1509,N_549,N_67);
nor U1510 (N_1510,N_89,N_580);
or U1511 (N_1511,N_641,N_309);
and U1512 (N_1512,N_662,N_25);
and U1513 (N_1513,N_166,N_760);
or U1514 (N_1514,N_615,N_287);
or U1515 (N_1515,N_651,N_539);
and U1516 (N_1516,N_422,N_947);
and U1517 (N_1517,N_57,N_287);
and U1518 (N_1518,N_690,N_265);
and U1519 (N_1519,N_535,N_632);
nor U1520 (N_1520,N_670,N_725);
and U1521 (N_1521,N_601,N_110);
and U1522 (N_1522,N_611,N_850);
or U1523 (N_1523,N_549,N_510);
and U1524 (N_1524,N_215,N_933);
xor U1525 (N_1525,N_63,N_305);
and U1526 (N_1526,N_148,N_314);
nor U1527 (N_1527,N_763,N_22);
or U1528 (N_1528,N_236,N_448);
and U1529 (N_1529,N_796,N_566);
or U1530 (N_1530,N_580,N_686);
and U1531 (N_1531,N_496,N_587);
nand U1532 (N_1532,N_752,N_964);
nand U1533 (N_1533,N_149,N_124);
nand U1534 (N_1534,N_451,N_4);
nor U1535 (N_1535,N_149,N_844);
or U1536 (N_1536,N_793,N_938);
and U1537 (N_1537,N_50,N_76);
xnor U1538 (N_1538,N_17,N_644);
nor U1539 (N_1539,N_563,N_284);
xnor U1540 (N_1540,N_979,N_858);
nor U1541 (N_1541,N_802,N_729);
nand U1542 (N_1542,N_114,N_901);
nand U1543 (N_1543,N_839,N_181);
nand U1544 (N_1544,N_427,N_228);
or U1545 (N_1545,N_300,N_15);
and U1546 (N_1546,N_685,N_364);
nand U1547 (N_1547,N_212,N_275);
or U1548 (N_1548,N_417,N_484);
and U1549 (N_1549,N_532,N_517);
nand U1550 (N_1550,N_204,N_663);
or U1551 (N_1551,N_34,N_993);
and U1552 (N_1552,N_880,N_378);
and U1553 (N_1553,N_835,N_33);
nor U1554 (N_1554,N_21,N_608);
nand U1555 (N_1555,N_506,N_831);
or U1556 (N_1556,N_435,N_668);
xnor U1557 (N_1557,N_148,N_474);
nand U1558 (N_1558,N_503,N_971);
nor U1559 (N_1559,N_395,N_986);
and U1560 (N_1560,N_291,N_511);
and U1561 (N_1561,N_624,N_854);
or U1562 (N_1562,N_251,N_838);
nor U1563 (N_1563,N_492,N_242);
nor U1564 (N_1564,N_956,N_45);
and U1565 (N_1565,N_939,N_207);
and U1566 (N_1566,N_381,N_495);
nand U1567 (N_1567,N_529,N_676);
xnor U1568 (N_1568,N_529,N_92);
or U1569 (N_1569,N_240,N_863);
and U1570 (N_1570,N_52,N_640);
nand U1571 (N_1571,N_690,N_803);
nor U1572 (N_1572,N_522,N_488);
or U1573 (N_1573,N_838,N_226);
and U1574 (N_1574,N_336,N_406);
nor U1575 (N_1575,N_685,N_865);
xnor U1576 (N_1576,N_310,N_382);
and U1577 (N_1577,N_518,N_780);
nand U1578 (N_1578,N_389,N_831);
and U1579 (N_1579,N_373,N_377);
and U1580 (N_1580,N_778,N_747);
and U1581 (N_1581,N_411,N_675);
xnor U1582 (N_1582,N_6,N_445);
and U1583 (N_1583,N_71,N_816);
nand U1584 (N_1584,N_915,N_787);
xor U1585 (N_1585,N_854,N_735);
and U1586 (N_1586,N_640,N_937);
or U1587 (N_1587,N_665,N_558);
nor U1588 (N_1588,N_42,N_488);
and U1589 (N_1589,N_152,N_114);
and U1590 (N_1590,N_317,N_182);
nor U1591 (N_1591,N_143,N_697);
nand U1592 (N_1592,N_310,N_255);
nor U1593 (N_1593,N_748,N_685);
or U1594 (N_1594,N_151,N_615);
nand U1595 (N_1595,N_855,N_622);
and U1596 (N_1596,N_472,N_669);
or U1597 (N_1597,N_118,N_362);
nor U1598 (N_1598,N_770,N_675);
nor U1599 (N_1599,N_316,N_368);
nand U1600 (N_1600,N_339,N_268);
and U1601 (N_1601,N_288,N_633);
or U1602 (N_1602,N_788,N_359);
nand U1603 (N_1603,N_318,N_723);
nand U1604 (N_1604,N_412,N_65);
or U1605 (N_1605,N_152,N_360);
nor U1606 (N_1606,N_192,N_656);
or U1607 (N_1607,N_291,N_643);
nor U1608 (N_1608,N_186,N_553);
nor U1609 (N_1609,N_326,N_503);
nand U1610 (N_1610,N_208,N_571);
and U1611 (N_1611,N_935,N_556);
and U1612 (N_1612,N_626,N_3);
nand U1613 (N_1613,N_36,N_736);
nand U1614 (N_1614,N_558,N_796);
xor U1615 (N_1615,N_7,N_556);
xor U1616 (N_1616,N_293,N_806);
nor U1617 (N_1617,N_93,N_766);
xnor U1618 (N_1618,N_710,N_664);
or U1619 (N_1619,N_12,N_49);
or U1620 (N_1620,N_431,N_920);
nand U1621 (N_1621,N_227,N_278);
nor U1622 (N_1622,N_547,N_387);
nand U1623 (N_1623,N_615,N_431);
and U1624 (N_1624,N_35,N_577);
and U1625 (N_1625,N_496,N_730);
nand U1626 (N_1626,N_759,N_63);
or U1627 (N_1627,N_978,N_16);
or U1628 (N_1628,N_180,N_247);
nand U1629 (N_1629,N_936,N_148);
and U1630 (N_1630,N_588,N_810);
nand U1631 (N_1631,N_554,N_119);
and U1632 (N_1632,N_586,N_977);
and U1633 (N_1633,N_593,N_37);
or U1634 (N_1634,N_453,N_264);
or U1635 (N_1635,N_976,N_870);
nand U1636 (N_1636,N_115,N_278);
and U1637 (N_1637,N_367,N_144);
or U1638 (N_1638,N_588,N_874);
and U1639 (N_1639,N_59,N_279);
and U1640 (N_1640,N_135,N_172);
xnor U1641 (N_1641,N_404,N_460);
or U1642 (N_1642,N_208,N_110);
xnor U1643 (N_1643,N_240,N_247);
nand U1644 (N_1644,N_773,N_227);
and U1645 (N_1645,N_930,N_979);
nand U1646 (N_1646,N_575,N_280);
nor U1647 (N_1647,N_551,N_809);
nor U1648 (N_1648,N_47,N_17);
nor U1649 (N_1649,N_179,N_111);
nor U1650 (N_1650,N_618,N_583);
or U1651 (N_1651,N_950,N_144);
xnor U1652 (N_1652,N_899,N_695);
nor U1653 (N_1653,N_789,N_265);
nor U1654 (N_1654,N_569,N_677);
or U1655 (N_1655,N_256,N_10);
nor U1656 (N_1656,N_382,N_488);
or U1657 (N_1657,N_263,N_840);
nor U1658 (N_1658,N_271,N_620);
nor U1659 (N_1659,N_421,N_15);
or U1660 (N_1660,N_925,N_203);
or U1661 (N_1661,N_320,N_590);
xnor U1662 (N_1662,N_30,N_128);
or U1663 (N_1663,N_717,N_969);
and U1664 (N_1664,N_135,N_599);
nor U1665 (N_1665,N_514,N_844);
and U1666 (N_1666,N_243,N_523);
xor U1667 (N_1667,N_717,N_646);
or U1668 (N_1668,N_289,N_836);
nor U1669 (N_1669,N_394,N_749);
and U1670 (N_1670,N_148,N_778);
xor U1671 (N_1671,N_794,N_818);
and U1672 (N_1672,N_647,N_83);
and U1673 (N_1673,N_330,N_165);
and U1674 (N_1674,N_151,N_160);
nor U1675 (N_1675,N_543,N_160);
or U1676 (N_1676,N_369,N_139);
nor U1677 (N_1677,N_597,N_638);
nor U1678 (N_1678,N_534,N_241);
and U1679 (N_1679,N_995,N_17);
nand U1680 (N_1680,N_306,N_378);
and U1681 (N_1681,N_716,N_636);
or U1682 (N_1682,N_67,N_160);
nand U1683 (N_1683,N_808,N_770);
nand U1684 (N_1684,N_400,N_513);
or U1685 (N_1685,N_419,N_191);
and U1686 (N_1686,N_224,N_647);
nand U1687 (N_1687,N_961,N_399);
and U1688 (N_1688,N_626,N_652);
nand U1689 (N_1689,N_126,N_900);
or U1690 (N_1690,N_480,N_569);
and U1691 (N_1691,N_558,N_808);
nand U1692 (N_1692,N_304,N_137);
nor U1693 (N_1693,N_369,N_306);
nand U1694 (N_1694,N_738,N_784);
or U1695 (N_1695,N_148,N_975);
nor U1696 (N_1696,N_395,N_426);
nand U1697 (N_1697,N_214,N_169);
xor U1698 (N_1698,N_374,N_117);
and U1699 (N_1699,N_806,N_372);
xor U1700 (N_1700,N_333,N_314);
nand U1701 (N_1701,N_969,N_829);
nor U1702 (N_1702,N_714,N_451);
and U1703 (N_1703,N_408,N_522);
and U1704 (N_1704,N_919,N_31);
and U1705 (N_1705,N_518,N_712);
nor U1706 (N_1706,N_65,N_431);
nor U1707 (N_1707,N_62,N_896);
nor U1708 (N_1708,N_679,N_521);
xnor U1709 (N_1709,N_580,N_739);
nand U1710 (N_1710,N_295,N_300);
and U1711 (N_1711,N_794,N_810);
or U1712 (N_1712,N_259,N_696);
nand U1713 (N_1713,N_86,N_979);
nor U1714 (N_1714,N_596,N_514);
nor U1715 (N_1715,N_342,N_607);
xor U1716 (N_1716,N_348,N_930);
nor U1717 (N_1717,N_300,N_768);
nand U1718 (N_1718,N_632,N_393);
xor U1719 (N_1719,N_847,N_894);
nand U1720 (N_1720,N_773,N_976);
and U1721 (N_1721,N_76,N_966);
xnor U1722 (N_1722,N_492,N_135);
and U1723 (N_1723,N_673,N_780);
and U1724 (N_1724,N_253,N_193);
nor U1725 (N_1725,N_887,N_819);
xnor U1726 (N_1726,N_897,N_505);
and U1727 (N_1727,N_435,N_105);
or U1728 (N_1728,N_50,N_128);
nand U1729 (N_1729,N_850,N_16);
or U1730 (N_1730,N_359,N_138);
nor U1731 (N_1731,N_587,N_852);
and U1732 (N_1732,N_144,N_564);
nand U1733 (N_1733,N_39,N_717);
xnor U1734 (N_1734,N_299,N_528);
or U1735 (N_1735,N_769,N_406);
and U1736 (N_1736,N_220,N_411);
and U1737 (N_1737,N_326,N_0);
nand U1738 (N_1738,N_378,N_835);
nand U1739 (N_1739,N_948,N_206);
and U1740 (N_1740,N_54,N_800);
or U1741 (N_1741,N_558,N_896);
nand U1742 (N_1742,N_236,N_523);
and U1743 (N_1743,N_798,N_294);
nand U1744 (N_1744,N_826,N_934);
and U1745 (N_1745,N_223,N_298);
nor U1746 (N_1746,N_932,N_141);
nor U1747 (N_1747,N_114,N_460);
and U1748 (N_1748,N_991,N_738);
nor U1749 (N_1749,N_469,N_0);
or U1750 (N_1750,N_886,N_728);
nor U1751 (N_1751,N_617,N_334);
xnor U1752 (N_1752,N_428,N_921);
and U1753 (N_1753,N_191,N_399);
or U1754 (N_1754,N_798,N_270);
and U1755 (N_1755,N_872,N_472);
nand U1756 (N_1756,N_273,N_279);
nand U1757 (N_1757,N_647,N_154);
or U1758 (N_1758,N_125,N_312);
nor U1759 (N_1759,N_809,N_1);
nor U1760 (N_1760,N_582,N_472);
nand U1761 (N_1761,N_370,N_41);
nor U1762 (N_1762,N_965,N_399);
nand U1763 (N_1763,N_696,N_557);
nand U1764 (N_1764,N_599,N_140);
nor U1765 (N_1765,N_123,N_149);
and U1766 (N_1766,N_20,N_292);
and U1767 (N_1767,N_100,N_823);
and U1768 (N_1768,N_288,N_363);
nor U1769 (N_1769,N_266,N_876);
nor U1770 (N_1770,N_795,N_809);
and U1771 (N_1771,N_56,N_810);
or U1772 (N_1772,N_566,N_295);
and U1773 (N_1773,N_476,N_121);
nor U1774 (N_1774,N_420,N_760);
and U1775 (N_1775,N_291,N_393);
or U1776 (N_1776,N_980,N_244);
xor U1777 (N_1777,N_887,N_194);
nand U1778 (N_1778,N_820,N_105);
nand U1779 (N_1779,N_30,N_298);
xor U1780 (N_1780,N_393,N_398);
xnor U1781 (N_1781,N_345,N_612);
nand U1782 (N_1782,N_424,N_802);
and U1783 (N_1783,N_73,N_317);
nand U1784 (N_1784,N_888,N_964);
nor U1785 (N_1785,N_282,N_448);
or U1786 (N_1786,N_210,N_273);
or U1787 (N_1787,N_667,N_868);
or U1788 (N_1788,N_816,N_814);
xor U1789 (N_1789,N_662,N_306);
and U1790 (N_1790,N_121,N_555);
nor U1791 (N_1791,N_906,N_788);
xor U1792 (N_1792,N_831,N_724);
nor U1793 (N_1793,N_274,N_473);
and U1794 (N_1794,N_57,N_344);
or U1795 (N_1795,N_162,N_95);
and U1796 (N_1796,N_405,N_725);
and U1797 (N_1797,N_612,N_896);
nor U1798 (N_1798,N_763,N_35);
nand U1799 (N_1799,N_658,N_937);
nor U1800 (N_1800,N_614,N_448);
nor U1801 (N_1801,N_903,N_213);
nor U1802 (N_1802,N_604,N_342);
and U1803 (N_1803,N_684,N_957);
nand U1804 (N_1804,N_128,N_820);
xor U1805 (N_1805,N_807,N_648);
nor U1806 (N_1806,N_885,N_508);
and U1807 (N_1807,N_988,N_631);
nor U1808 (N_1808,N_534,N_621);
nand U1809 (N_1809,N_121,N_280);
or U1810 (N_1810,N_858,N_275);
or U1811 (N_1811,N_698,N_375);
or U1812 (N_1812,N_540,N_88);
and U1813 (N_1813,N_456,N_840);
nand U1814 (N_1814,N_450,N_558);
and U1815 (N_1815,N_164,N_319);
nand U1816 (N_1816,N_48,N_914);
nor U1817 (N_1817,N_289,N_378);
or U1818 (N_1818,N_608,N_451);
nor U1819 (N_1819,N_977,N_621);
nand U1820 (N_1820,N_871,N_413);
xnor U1821 (N_1821,N_789,N_780);
and U1822 (N_1822,N_702,N_37);
nor U1823 (N_1823,N_475,N_694);
xor U1824 (N_1824,N_97,N_663);
nor U1825 (N_1825,N_597,N_466);
or U1826 (N_1826,N_203,N_400);
nand U1827 (N_1827,N_162,N_556);
or U1828 (N_1828,N_54,N_67);
nor U1829 (N_1829,N_393,N_438);
nand U1830 (N_1830,N_109,N_755);
and U1831 (N_1831,N_369,N_919);
or U1832 (N_1832,N_821,N_285);
nand U1833 (N_1833,N_559,N_697);
nand U1834 (N_1834,N_699,N_240);
nor U1835 (N_1835,N_83,N_82);
nand U1836 (N_1836,N_955,N_257);
xnor U1837 (N_1837,N_397,N_644);
nor U1838 (N_1838,N_276,N_968);
nand U1839 (N_1839,N_715,N_618);
and U1840 (N_1840,N_129,N_963);
nand U1841 (N_1841,N_460,N_564);
and U1842 (N_1842,N_453,N_268);
nor U1843 (N_1843,N_599,N_270);
nor U1844 (N_1844,N_571,N_709);
nor U1845 (N_1845,N_191,N_424);
nand U1846 (N_1846,N_50,N_990);
and U1847 (N_1847,N_106,N_495);
nand U1848 (N_1848,N_125,N_568);
nor U1849 (N_1849,N_282,N_214);
or U1850 (N_1850,N_86,N_531);
nand U1851 (N_1851,N_208,N_194);
and U1852 (N_1852,N_745,N_310);
nor U1853 (N_1853,N_117,N_241);
nor U1854 (N_1854,N_108,N_486);
and U1855 (N_1855,N_292,N_867);
or U1856 (N_1856,N_767,N_148);
and U1857 (N_1857,N_687,N_267);
or U1858 (N_1858,N_282,N_644);
or U1859 (N_1859,N_50,N_279);
xor U1860 (N_1860,N_111,N_414);
nand U1861 (N_1861,N_168,N_358);
nor U1862 (N_1862,N_644,N_234);
and U1863 (N_1863,N_268,N_679);
and U1864 (N_1864,N_92,N_872);
or U1865 (N_1865,N_890,N_249);
nor U1866 (N_1866,N_952,N_774);
or U1867 (N_1867,N_88,N_527);
nand U1868 (N_1868,N_794,N_859);
or U1869 (N_1869,N_825,N_807);
or U1870 (N_1870,N_940,N_70);
nand U1871 (N_1871,N_567,N_861);
nor U1872 (N_1872,N_148,N_345);
or U1873 (N_1873,N_431,N_131);
nor U1874 (N_1874,N_936,N_932);
nand U1875 (N_1875,N_776,N_610);
nand U1876 (N_1876,N_734,N_680);
xnor U1877 (N_1877,N_747,N_989);
and U1878 (N_1878,N_303,N_877);
nor U1879 (N_1879,N_978,N_835);
nand U1880 (N_1880,N_421,N_191);
or U1881 (N_1881,N_241,N_920);
and U1882 (N_1882,N_195,N_662);
nor U1883 (N_1883,N_958,N_932);
and U1884 (N_1884,N_738,N_728);
nand U1885 (N_1885,N_557,N_350);
and U1886 (N_1886,N_871,N_676);
or U1887 (N_1887,N_357,N_321);
nor U1888 (N_1888,N_72,N_429);
and U1889 (N_1889,N_356,N_797);
or U1890 (N_1890,N_33,N_619);
nand U1891 (N_1891,N_499,N_368);
or U1892 (N_1892,N_148,N_295);
or U1893 (N_1893,N_124,N_159);
and U1894 (N_1894,N_466,N_281);
or U1895 (N_1895,N_77,N_542);
nor U1896 (N_1896,N_74,N_499);
nand U1897 (N_1897,N_573,N_535);
and U1898 (N_1898,N_114,N_43);
and U1899 (N_1899,N_695,N_501);
and U1900 (N_1900,N_373,N_296);
nand U1901 (N_1901,N_779,N_857);
xnor U1902 (N_1902,N_396,N_967);
nor U1903 (N_1903,N_321,N_894);
and U1904 (N_1904,N_190,N_56);
nor U1905 (N_1905,N_666,N_653);
xnor U1906 (N_1906,N_464,N_827);
or U1907 (N_1907,N_743,N_207);
nor U1908 (N_1908,N_60,N_923);
or U1909 (N_1909,N_608,N_480);
nor U1910 (N_1910,N_515,N_142);
nand U1911 (N_1911,N_764,N_568);
nor U1912 (N_1912,N_795,N_224);
nor U1913 (N_1913,N_705,N_641);
or U1914 (N_1914,N_686,N_903);
xnor U1915 (N_1915,N_991,N_230);
nand U1916 (N_1916,N_695,N_503);
or U1917 (N_1917,N_960,N_4);
nor U1918 (N_1918,N_706,N_136);
or U1919 (N_1919,N_34,N_122);
and U1920 (N_1920,N_762,N_293);
nand U1921 (N_1921,N_773,N_609);
or U1922 (N_1922,N_747,N_562);
nor U1923 (N_1923,N_878,N_320);
nand U1924 (N_1924,N_565,N_802);
xnor U1925 (N_1925,N_702,N_79);
and U1926 (N_1926,N_188,N_51);
nor U1927 (N_1927,N_29,N_529);
and U1928 (N_1928,N_149,N_550);
xor U1929 (N_1929,N_35,N_769);
and U1930 (N_1930,N_442,N_436);
or U1931 (N_1931,N_614,N_496);
or U1932 (N_1932,N_819,N_36);
xnor U1933 (N_1933,N_896,N_521);
and U1934 (N_1934,N_342,N_84);
nand U1935 (N_1935,N_705,N_426);
nor U1936 (N_1936,N_793,N_260);
or U1937 (N_1937,N_224,N_411);
and U1938 (N_1938,N_10,N_881);
or U1939 (N_1939,N_862,N_118);
nor U1940 (N_1940,N_887,N_570);
nand U1941 (N_1941,N_311,N_263);
nand U1942 (N_1942,N_42,N_120);
nor U1943 (N_1943,N_500,N_934);
or U1944 (N_1944,N_872,N_742);
xor U1945 (N_1945,N_255,N_94);
and U1946 (N_1946,N_740,N_334);
xor U1947 (N_1947,N_340,N_492);
nor U1948 (N_1948,N_691,N_175);
nand U1949 (N_1949,N_209,N_246);
or U1950 (N_1950,N_888,N_728);
nor U1951 (N_1951,N_458,N_647);
and U1952 (N_1952,N_440,N_630);
xor U1953 (N_1953,N_29,N_237);
nand U1954 (N_1954,N_549,N_33);
or U1955 (N_1955,N_703,N_362);
and U1956 (N_1956,N_936,N_376);
and U1957 (N_1957,N_551,N_886);
xor U1958 (N_1958,N_661,N_986);
or U1959 (N_1959,N_566,N_715);
nand U1960 (N_1960,N_404,N_953);
and U1961 (N_1961,N_469,N_70);
and U1962 (N_1962,N_506,N_604);
or U1963 (N_1963,N_140,N_14);
nand U1964 (N_1964,N_171,N_376);
nand U1965 (N_1965,N_2,N_555);
nand U1966 (N_1966,N_644,N_480);
and U1967 (N_1967,N_120,N_188);
or U1968 (N_1968,N_772,N_625);
nor U1969 (N_1969,N_794,N_763);
nand U1970 (N_1970,N_454,N_960);
and U1971 (N_1971,N_323,N_724);
nand U1972 (N_1972,N_672,N_572);
nand U1973 (N_1973,N_450,N_89);
nand U1974 (N_1974,N_952,N_858);
and U1975 (N_1975,N_403,N_91);
or U1976 (N_1976,N_313,N_445);
nor U1977 (N_1977,N_524,N_91);
or U1978 (N_1978,N_64,N_426);
and U1979 (N_1979,N_829,N_920);
nand U1980 (N_1980,N_654,N_911);
nor U1981 (N_1981,N_228,N_873);
nand U1982 (N_1982,N_912,N_430);
nand U1983 (N_1983,N_628,N_914);
or U1984 (N_1984,N_481,N_105);
xor U1985 (N_1985,N_700,N_919);
nor U1986 (N_1986,N_292,N_962);
nand U1987 (N_1987,N_482,N_208);
nand U1988 (N_1988,N_421,N_253);
nand U1989 (N_1989,N_729,N_138);
nand U1990 (N_1990,N_596,N_17);
and U1991 (N_1991,N_439,N_495);
and U1992 (N_1992,N_349,N_267);
nor U1993 (N_1993,N_217,N_204);
nor U1994 (N_1994,N_492,N_303);
xor U1995 (N_1995,N_295,N_764);
xor U1996 (N_1996,N_247,N_61);
or U1997 (N_1997,N_719,N_219);
nor U1998 (N_1998,N_211,N_662);
nor U1999 (N_1999,N_479,N_506);
nor U2000 (N_2000,N_1821,N_1755);
nor U2001 (N_2001,N_1568,N_1324);
or U2002 (N_2002,N_1677,N_1564);
nor U2003 (N_2003,N_1203,N_1199);
nor U2004 (N_2004,N_1849,N_1365);
nand U2005 (N_2005,N_1599,N_1942);
nor U2006 (N_2006,N_1055,N_1245);
nand U2007 (N_2007,N_1156,N_1391);
xor U2008 (N_2008,N_1373,N_1032);
nor U2009 (N_2009,N_1516,N_1817);
nor U2010 (N_2010,N_1155,N_1865);
xor U2011 (N_2011,N_1027,N_1533);
nand U2012 (N_2012,N_1911,N_1746);
or U2013 (N_2013,N_1527,N_1308);
and U2014 (N_2014,N_1971,N_1885);
or U2015 (N_2015,N_1358,N_1503);
and U2016 (N_2016,N_1253,N_1833);
xnor U2017 (N_2017,N_1091,N_1784);
nor U2018 (N_2018,N_1222,N_1067);
nor U2019 (N_2019,N_1743,N_1194);
nor U2020 (N_2020,N_1707,N_1600);
or U2021 (N_2021,N_1827,N_1400);
nand U2022 (N_2022,N_1948,N_1133);
nand U2023 (N_2023,N_1963,N_1584);
nor U2024 (N_2024,N_1349,N_1529);
nor U2025 (N_2025,N_1770,N_1140);
or U2026 (N_2026,N_1699,N_1454);
and U2027 (N_2027,N_1730,N_1748);
or U2028 (N_2028,N_1830,N_1030);
and U2029 (N_2029,N_1659,N_1983);
nor U2030 (N_2030,N_1357,N_1112);
or U2031 (N_2031,N_1145,N_1386);
nor U2032 (N_2032,N_1103,N_1306);
nand U2033 (N_2033,N_1094,N_1903);
nor U2034 (N_2034,N_1513,N_1955);
nor U2035 (N_2035,N_1325,N_1902);
or U2036 (N_2036,N_1774,N_1406);
or U2037 (N_2037,N_1348,N_1184);
and U2038 (N_2038,N_1065,N_1340);
or U2039 (N_2039,N_1173,N_1123);
and U2040 (N_2040,N_1058,N_1138);
nand U2041 (N_2041,N_1613,N_1546);
or U2042 (N_2042,N_1897,N_1064);
nand U2043 (N_2043,N_1536,N_1585);
and U2044 (N_2044,N_1303,N_1795);
or U2045 (N_2045,N_1976,N_1650);
or U2046 (N_2046,N_1152,N_1174);
and U2047 (N_2047,N_1680,N_1692);
nand U2048 (N_2048,N_1139,N_1968);
nor U2049 (N_2049,N_1854,N_1118);
or U2050 (N_2050,N_1204,N_1090);
nand U2051 (N_2051,N_1061,N_1025);
nand U2052 (N_2052,N_1809,N_1832);
nand U2053 (N_2053,N_1352,N_1858);
nor U2054 (N_2054,N_1190,N_1507);
and U2055 (N_2055,N_1719,N_1760);
nand U2056 (N_2056,N_1597,N_1432);
nor U2057 (N_2057,N_1390,N_1732);
and U2058 (N_2058,N_1250,N_1901);
nand U2059 (N_2059,N_1430,N_1193);
nand U2060 (N_2060,N_1860,N_1724);
nand U2061 (N_2061,N_1814,N_1292);
and U2062 (N_2062,N_1894,N_1281);
nor U2063 (N_2063,N_1812,N_1326);
nand U2064 (N_2064,N_1410,N_1371);
or U2065 (N_2065,N_1399,N_1289);
and U2066 (N_2066,N_1653,N_1550);
xnor U2067 (N_2067,N_1455,N_1823);
xor U2068 (N_2068,N_1962,N_1904);
or U2069 (N_2069,N_1187,N_1670);
nor U2070 (N_2070,N_1016,N_1512);
nor U2071 (N_2071,N_1481,N_1877);
xnor U2072 (N_2072,N_1021,N_1488);
or U2073 (N_2073,N_1201,N_1886);
and U2074 (N_2074,N_1736,N_1310);
or U2075 (N_2075,N_1034,N_1551);
xor U2076 (N_2076,N_1500,N_1701);
xnor U2077 (N_2077,N_1739,N_1323);
and U2078 (N_2078,N_1618,N_1175);
xor U2079 (N_2079,N_1850,N_1007);
nand U2080 (N_2080,N_1367,N_1179);
and U2081 (N_2081,N_1335,N_1652);
and U2082 (N_2082,N_1545,N_1624);
nand U2083 (N_2083,N_1511,N_1638);
and U2084 (N_2084,N_1940,N_1045);
and U2085 (N_2085,N_1200,N_1334);
and U2086 (N_2086,N_1900,N_1177);
nor U2087 (N_2087,N_1210,N_1189);
nor U2088 (N_2088,N_1986,N_1341);
and U2089 (N_2089,N_1101,N_1110);
nand U2090 (N_2090,N_1398,N_1567);
nand U2091 (N_2091,N_1429,N_1437);
nor U2092 (N_2092,N_1845,N_1696);
or U2093 (N_2093,N_1231,N_1839);
and U2094 (N_2094,N_1104,N_1427);
or U2095 (N_2095,N_1689,N_1959);
xnor U2096 (N_2096,N_1001,N_1219);
nor U2097 (N_2097,N_1887,N_1148);
nand U2098 (N_2098,N_1977,N_1772);
nor U2099 (N_2099,N_1428,N_1908);
and U2100 (N_2100,N_1077,N_1588);
nor U2101 (N_2101,N_1128,N_1444);
nand U2102 (N_2102,N_1998,N_1220);
nand U2103 (N_2103,N_1987,N_1873);
or U2104 (N_2104,N_1799,N_1441);
or U2105 (N_2105,N_1169,N_1327);
nor U2106 (N_2106,N_1017,N_1785);
and U2107 (N_2107,N_1688,N_1251);
or U2108 (N_2108,N_1861,N_1452);
and U2109 (N_2109,N_1708,N_1639);
nor U2110 (N_2110,N_1403,N_1848);
and U2111 (N_2111,N_1037,N_1338);
nand U2112 (N_2112,N_1046,N_1615);
nand U2113 (N_2113,N_1402,N_1616);
or U2114 (N_2114,N_1182,N_1658);
nand U2115 (N_2115,N_1686,N_1288);
xor U2116 (N_2116,N_1703,N_1996);
nor U2117 (N_2117,N_1763,N_1394);
xnor U2118 (N_2118,N_1361,N_1066);
nand U2119 (N_2119,N_1872,N_1217);
or U2120 (N_2120,N_1125,N_1715);
xnor U2121 (N_2121,N_1496,N_1958);
or U2122 (N_2122,N_1824,N_1723);
nand U2123 (N_2123,N_1997,N_1646);
and U2124 (N_2124,N_1153,N_1293);
xor U2125 (N_2125,N_1137,N_1075);
nor U2126 (N_2126,N_1891,N_1031);
nor U2127 (N_2127,N_1793,N_1810);
nor U2128 (N_2128,N_1295,N_1018);
and U2129 (N_2129,N_1636,N_1521);
nand U2130 (N_2130,N_1411,N_1022);
nand U2131 (N_2131,N_1279,N_1236);
nor U2132 (N_2132,N_1843,N_1314);
or U2133 (N_2133,N_1859,N_1211);
and U2134 (N_2134,N_1144,N_1028);
nand U2135 (N_2135,N_1705,N_1426);
or U2136 (N_2136,N_1353,N_1079);
and U2137 (N_2137,N_1518,N_1741);
nor U2138 (N_2138,N_1434,N_1157);
and U2139 (N_2139,N_1811,N_1769);
xnor U2140 (N_2140,N_1890,N_1667);
nor U2141 (N_2141,N_1524,N_1019);
or U2142 (N_2142,N_1423,N_1299);
nor U2143 (N_2143,N_1060,N_1643);
and U2144 (N_2144,N_1913,N_1246);
nor U2145 (N_2145,N_1242,N_1970);
and U2146 (N_2146,N_1068,N_1951);
or U2147 (N_2147,N_1498,N_1825);
or U2148 (N_2148,N_1501,N_1796);
nor U2149 (N_2149,N_1284,N_1583);
nor U2150 (N_2150,N_1465,N_1176);
and U2151 (N_2151,N_1267,N_1107);
nand U2152 (N_2152,N_1582,N_1440);
nor U2153 (N_2153,N_1526,N_1505);
and U2154 (N_2154,N_1758,N_1035);
nand U2155 (N_2155,N_1062,N_1744);
or U2156 (N_2156,N_1893,N_1491);
or U2157 (N_2157,N_1054,N_1617);
nand U2158 (N_2158,N_1072,N_1591);
and U2159 (N_2159,N_1554,N_1366);
xor U2160 (N_2160,N_1806,N_1544);
or U2161 (N_2161,N_1604,N_1606);
or U2162 (N_2162,N_1563,N_1180);
nor U2163 (N_2163,N_1842,N_1074);
and U2164 (N_2164,N_1671,N_1385);
nor U2165 (N_2165,N_1662,N_1960);
xnor U2166 (N_2166,N_1837,N_1502);
or U2167 (N_2167,N_1108,N_1188);
and U2168 (N_2168,N_1649,N_1642);
nand U2169 (N_2169,N_1761,N_1487);
nor U2170 (N_2170,N_1376,N_1298);
or U2171 (N_2171,N_1871,N_1504);
nor U2172 (N_2172,N_1548,N_1451);
nor U2173 (N_2173,N_1731,N_1834);
nand U2174 (N_2174,N_1905,N_1863);
or U2175 (N_2175,N_1151,N_1207);
xnor U2176 (N_2176,N_1921,N_1640);
nor U2177 (N_2177,N_1360,N_1126);
nor U2178 (N_2178,N_1425,N_1186);
and U2179 (N_2179,N_1950,N_1209);
nand U2180 (N_2180,N_1438,N_1939);
nand U2181 (N_2181,N_1866,N_1764);
nor U2182 (N_2182,N_1473,N_1978);
xnor U2183 (N_2183,N_1135,N_1721);
xor U2184 (N_2184,N_1408,N_1880);
nor U2185 (N_2185,N_1573,N_1931);
and U2186 (N_2186,N_1934,N_1695);
nor U2187 (N_2187,N_1131,N_1124);
and U2188 (N_2188,N_1556,N_1879);
nand U2189 (N_2189,N_1274,N_1710);
xnor U2190 (N_2190,N_1059,N_1552);
xor U2191 (N_2191,N_1611,N_1170);
and U2192 (N_2192,N_1844,N_1047);
nand U2193 (N_2193,N_1085,N_1006);
nor U2194 (N_2194,N_1127,N_1183);
nand U2195 (N_2195,N_1776,N_1712);
and U2196 (N_2196,N_1633,N_1766);
xnor U2197 (N_2197,N_1413,N_1419);
and U2198 (N_2198,N_1494,N_1792);
xor U2199 (N_2199,N_1244,N_1158);
nor U2200 (N_2200,N_1078,N_1212);
and U2201 (N_2201,N_1927,N_1716);
xor U2202 (N_2202,N_1531,N_1223);
or U2203 (N_2203,N_1694,N_1422);
or U2204 (N_2204,N_1480,N_1215);
nand U2205 (N_2205,N_1742,N_1956);
and U2206 (N_2206,N_1704,N_1973);
nand U2207 (N_2207,N_1459,N_1275);
nand U2208 (N_2208,N_1778,N_1549);
or U2209 (N_2209,N_1383,N_1964);
and U2210 (N_2210,N_1530,N_1162);
or U2211 (N_2211,N_1555,N_1424);
and U2212 (N_2212,N_1664,N_1302);
nand U2213 (N_2213,N_1097,N_1575);
nand U2214 (N_2214,N_1994,N_1256);
nor U2215 (N_2215,N_1629,N_1924);
and U2216 (N_2216,N_1661,N_1294);
nor U2217 (N_2217,N_1490,N_1953);
or U2218 (N_2218,N_1278,N_1166);
nor U2219 (N_2219,N_1840,N_1593);
nand U2220 (N_2220,N_1336,N_1630);
nand U2221 (N_2221,N_1375,N_1925);
nor U2222 (N_2222,N_1813,N_1782);
or U2223 (N_2223,N_1102,N_1938);
nand U2224 (N_2224,N_1343,N_1095);
nand U2225 (N_2225,N_1816,N_1651);
nor U2226 (N_2226,N_1315,N_1759);
nor U2227 (N_2227,N_1836,N_1405);
nand U2228 (N_2228,N_1240,N_1436);
or U2229 (N_2229,N_1468,N_1557);
xor U2230 (N_2230,N_1098,N_1087);
nand U2231 (N_2231,N_1851,N_1198);
and U2232 (N_2232,N_1989,N_1482);
nand U2233 (N_2233,N_1446,N_1589);
nor U2234 (N_2234,N_1797,N_1846);
nor U2235 (N_2235,N_1355,N_1111);
or U2236 (N_2236,N_1635,N_1421);
nand U2237 (N_2237,N_1416,N_1679);
and U2238 (N_2238,N_1063,N_1196);
or U2239 (N_2239,N_1726,N_1002);
nand U2240 (N_2240,N_1547,N_1882);
or U2241 (N_2241,N_1450,N_1614);
or U2242 (N_2242,N_1579,N_1261);
xor U2243 (N_2243,N_1449,N_1191);
or U2244 (N_2244,N_1999,N_1388);
or U2245 (N_2245,N_1313,N_1907);
nor U2246 (N_2246,N_1870,N_1684);
nor U2247 (N_2247,N_1808,N_1457);
or U2248 (N_2248,N_1309,N_1172);
or U2249 (N_2249,N_1566,N_1243);
or U2250 (N_2250,N_1841,N_1147);
nand U2251 (N_2251,N_1706,N_1625);
or U2252 (N_2252,N_1478,N_1775);
xor U2253 (N_2253,N_1750,N_1409);
nor U2254 (N_2254,N_1470,N_1733);
and U2255 (N_2255,N_1937,N_1881);
nor U2256 (N_2256,N_1690,N_1892);
nor U2257 (N_2257,N_1722,N_1165);
and U2258 (N_2258,N_1985,N_1666);
nand U2259 (N_2259,N_1300,N_1668);
nor U2260 (N_2260,N_1864,N_1751);
and U2261 (N_2261,N_1113,N_1943);
xor U2262 (N_2262,N_1915,N_1917);
nand U2263 (N_2263,N_1254,N_1202);
nand U2264 (N_2264,N_1637,N_1559);
or U2265 (N_2265,N_1051,N_1561);
nand U2266 (N_2266,N_1757,N_1869);
and U2267 (N_2267,N_1601,N_1673);
or U2268 (N_2268,N_1713,N_1944);
nor U2269 (N_2269,N_1607,N_1081);
nor U2270 (N_2270,N_1076,N_1266);
xor U2271 (N_2271,N_1477,N_1280);
nand U2272 (N_2272,N_1804,N_1070);
and U2273 (N_2273,N_1936,N_1312);
nor U2274 (N_2274,N_1012,N_1855);
nor U2275 (N_2275,N_1458,N_1935);
xor U2276 (N_2276,N_1484,N_1558);
nand U2277 (N_2277,N_1628,N_1933);
or U2278 (N_2278,N_1553,N_1020);
and U2279 (N_2279,N_1768,N_1291);
and U2280 (N_2280,N_1486,N_1163);
nor U2281 (N_2281,N_1109,N_1359);
and U2282 (N_2282,N_1004,N_1515);
nor U2283 (N_2283,N_1205,N_1213);
and U2284 (N_2284,N_1053,N_1578);
or U2285 (N_2285,N_1456,N_1984);
and U2286 (N_2286,N_1218,N_1050);
and U2287 (N_2287,N_1702,N_1073);
nand U2288 (N_2288,N_1290,N_1522);
nand U2289 (N_2289,N_1332,N_1619);
nor U2290 (N_2290,N_1401,N_1479);
and U2291 (N_2291,N_1467,N_1594);
nor U2292 (N_2292,N_1899,N_1117);
and U2293 (N_2293,N_1418,N_1232);
nand U2294 (N_2294,N_1700,N_1822);
nand U2295 (N_2295,N_1954,N_1499);
or U2296 (N_2296,N_1675,N_1756);
or U2297 (N_2297,N_1453,N_1096);
or U2298 (N_2298,N_1698,N_1374);
and U2299 (N_2299,N_1678,N_1273);
nor U2300 (N_2300,N_1168,N_1415);
or U2301 (N_2301,N_1146,N_1981);
or U2302 (N_2302,N_1687,N_1788);
nand U2303 (N_2303,N_1929,N_1142);
or U2304 (N_2304,N_1762,N_1008);
or U2305 (N_2305,N_1041,N_1161);
xnor U2306 (N_2306,N_1884,N_1495);
xnor U2307 (N_2307,N_1779,N_1829);
and U2308 (N_2308,N_1995,N_1377);
nor U2309 (N_2309,N_1777,N_1270);
nand U2310 (N_2310,N_1230,N_1791);
and U2311 (N_2311,N_1447,N_1979);
and U2312 (N_2312,N_1141,N_1697);
or U2313 (N_2313,N_1036,N_1043);
and U2314 (N_2314,N_1026,N_1525);
nand U2315 (N_2315,N_1681,N_1178);
nor U2316 (N_2316,N_1268,N_1462);
and U2317 (N_2317,N_1412,N_1317);
nand U2318 (N_2318,N_1598,N_1541);
nor U2319 (N_2319,N_1815,N_1534);
nand U2320 (N_2320,N_1714,N_1003);
nor U2321 (N_2321,N_1347,N_1439);
and U2322 (N_2322,N_1862,N_1835);
or U2323 (N_2323,N_1789,N_1656);
nand U2324 (N_2324,N_1234,N_1519);
nor U2325 (N_2325,N_1605,N_1923);
or U2326 (N_2326,N_1263,N_1537);
xor U2327 (N_2327,N_1116,N_1057);
nor U2328 (N_2328,N_1602,N_1532);
and U2329 (N_2329,N_1920,N_1644);
nor U2330 (N_2330,N_1328,N_1171);
xor U2331 (N_2331,N_1595,N_1647);
and U2332 (N_2332,N_1596,N_1330);
and U2333 (N_2333,N_1233,N_1181);
and U2334 (N_2334,N_1195,N_1569);
nand U2335 (N_2335,N_1826,N_1350);
and U2336 (N_2336,N_1622,N_1961);
nor U2337 (N_2337,N_1928,N_1331);
and U2338 (N_2338,N_1105,N_1329);
nand U2339 (N_2339,N_1780,N_1235);
and U2340 (N_2340,N_1922,N_1720);
and U2341 (N_2341,N_1346,N_1926);
or U2342 (N_2342,N_1800,N_1773);
nand U2343 (N_2343,N_1991,N_1319);
nand U2344 (N_2344,N_1645,N_1287);
nor U2345 (N_2345,N_1572,N_1868);
nand U2346 (N_2346,N_1807,N_1492);
and U2347 (N_2347,N_1787,N_1039);
nand U2348 (N_2348,N_1693,N_1307);
and U2349 (N_2349,N_1794,N_1208);
or U2350 (N_2350,N_1129,N_1009);
nand U2351 (N_2351,N_1587,N_1949);
or U2352 (N_2352,N_1754,N_1150);
nand U2353 (N_2353,N_1276,N_1100);
nand U2354 (N_2354,N_1819,N_1257);
and U2355 (N_2355,N_1586,N_1167);
nand U2356 (N_2356,N_1185,N_1623);
or U2357 (N_2357,N_1119,N_1655);
and U2358 (N_2358,N_1729,N_1691);
and U2359 (N_2359,N_1069,N_1044);
nand U2360 (N_2360,N_1369,N_1672);
nor U2361 (N_2361,N_1363,N_1471);
and U2362 (N_2362,N_1115,N_1433);
and U2363 (N_2363,N_1539,N_1771);
or U2364 (N_2364,N_1005,N_1466);
xor U2365 (N_2365,N_1576,N_1874);
nand U2366 (N_2366,N_1483,N_1620);
nand U2367 (N_2367,N_1737,N_1380);
nor U2368 (N_2368,N_1896,N_1241);
nor U2369 (N_2369,N_1420,N_1475);
and U2370 (N_2370,N_1038,N_1608);
xor U2371 (N_2371,N_1321,N_1990);
and U2372 (N_2372,N_1626,N_1838);
nor U2373 (N_2373,N_1918,N_1969);
nor U2374 (N_2374,N_1445,N_1083);
nor U2375 (N_2375,N_1497,N_1192);
or U2376 (N_2376,N_1510,N_1734);
nor U2377 (N_2377,N_1485,N_1122);
and U2378 (N_2378,N_1206,N_1802);
nand U2379 (N_2379,N_1876,N_1946);
or U2380 (N_2380,N_1000,N_1229);
and U2381 (N_2381,N_1238,N_1283);
or U2382 (N_2382,N_1344,N_1381);
or U2383 (N_2383,N_1082,N_1049);
and U2384 (N_2384,N_1581,N_1752);
xnor U2385 (N_2385,N_1297,N_1803);
nor U2386 (N_2386,N_1029,N_1945);
nand U2387 (N_2387,N_1387,N_1224);
xor U2388 (N_2388,N_1023,N_1010);
nand U2389 (N_2389,N_1783,N_1506);
or U2390 (N_2390,N_1271,N_1443);
nor U2391 (N_2391,N_1852,N_1080);
and U2392 (N_2392,N_1669,N_1609);
nor U2393 (N_2393,N_1011,N_1132);
nand U2394 (N_2394,N_1489,N_1033);
xor U2395 (N_2395,N_1590,N_1048);
nand U2396 (N_2396,N_1382,N_1464);
nor U2397 (N_2397,N_1379,N_1024);
nor U2398 (N_2398,N_1318,N_1895);
and U2399 (N_2399,N_1831,N_1260);
nor U2400 (N_2400,N_1368,N_1747);
nor U2401 (N_2401,N_1898,N_1265);
nor U2402 (N_2402,N_1397,N_1711);
nand U2403 (N_2403,N_1974,N_1717);
or U2404 (N_2404,N_1745,N_1889);
or U2405 (N_2405,N_1565,N_1941);
or U2406 (N_2406,N_1930,N_1610);
nor U2407 (N_2407,N_1296,N_1740);
nor U2408 (N_2408,N_1627,N_1992);
or U2409 (N_2409,N_1857,N_1654);
or U2410 (N_2410,N_1523,N_1682);
and U2411 (N_2411,N_1916,N_1237);
nor U2412 (N_2412,N_1648,N_1538);
and U2413 (N_2413,N_1683,N_1993);
nor U2414 (N_2414,N_1988,N_1632);
nand U2415 (N_2415,N_1226,N_1906);
and U2416 (N_2416,N_1476,N_1560);
nand U2417 (N_2417,N_1781,N_1417);
and U2418 (N_2418,N_1339,N_1372);
and U2419 (N_2419,N_1227,N_1965);
and U2420 (N_2420,N_1134,N_1042);
nand U2421 (N_2421,N_1216,N_1092);
nand U2422 (N_2422,N_1252,N_1255);
nand U2423 (N_2423,N_1738,N_1362);
and U2424 (N_2424,N_1249,N_1801);
and U2425 (N_2425,N_1910,N_1258);
or U2426 (N_2426,N_1542,N_1316);
nor U2427 (N_2427,N_1725,N_1214);
nor U2428 (N_2428,N_1665,N_1393);
or U2429 (N_2429,N_1463,N_1728);
or U2430 (N_2430,N_1735,N_1269);
and U2431 (N_2431,N_1089,N_1520);
and U2432 (N_2432,N_1320,N_1407);
or U2433 (N_2433,N_1972,N_1197);
and U2434 (N_2434,N_1957,N_1143);
or U2435 (N_2435,N_1088,N_1878);
nand U2436 (N_2436,N_1574,N_1389);
nor U2437 (N_2437,N_1460,N_1370);
or U2438 (N_2438,N_1947,N_1718);
or U2439 (N_2439,N_1818,N_1277);
and U2440 (N_2440,N_1571,N_1514);
nand U2441 (N_2441,N_1099,N_1975);
xnor U2442 (N_2442,N_1786,N_1404);
nor U2443 (N_2443,N_1631,N_1322);
or U2444 (N_2444,N_1262,N_1493);
nor U2445 (N_2445,N_1674,N_1474);
nand U2446 (N_2446,N_1392,N_1264);
and U2447 (N_2447,N_1888,N_1071);
and U2448 (N_2448,N_1120,N_1982);
nor U2449 (N_2449,N_1286,N_1753);
nand U2450 (N_2450,N_1106,N_1966);
and U2451 (N_2451,N_1384,N_1912);
nor U2452 (N_2452,N_1364,N_1657);
or U2453 (N_2453,N_1304,N_1228);
and U2454 (N_2454,N_1621,N_1749);
nor U2455 (N_2455,N_1121,N_1847);
nor U2456 (N_2456,N_1448,N_1867);
or U2457 (N_2457,N_1272,N_1580);
nand U2458 (N_2458,N_1875,N_1056);
and U2459 (N_2459,N_1154,N_1562);
or U2460 (N_2460,N_1040,N_1239);
and U2461 (N_2461,N_1472,N_1798);
and U2462 (N_2462,N_1767,N_1932);
or U2463 (N_2463,N_1820,N_1805);
or U2464 (N_2464,N_1337,N_1414);
or U2465 (N_2465,N_1221,N_1356);
nand U2466 (N_2466,N_1952,N_1709);
and U2467 (N_2467,N_1285,N_1114);
nor U2468 (N_2468,N_1282,N_1435);
and U2469 (N_2469,N_1311,N_1431);
and U2470 (N_2470,N_1225,N_1663);
or U2471 (N_2471,N_1164,N_1790);
and U2472 (N_2472,N_1685,N_1084);
nor U2473 (N_2473,N_1828,N_1914);
xnor U2474 (N_2474,N_1469,N_1015);
or U2475 (N_2475,N_1013,N_1136);
xor U2476 (N_2476,N_1508,N_1676);
nand U2477 (N_2477,N_1612,N_1093);
and U2478 (N_2478,N_1641,N_1461);
nand U2479 (N_2479,N_1919,N_1351);
or U2480 (N_2480,N_1345,N_1577);
and U2481 (N_2481,N_1378,N_1509);
nor U2482 (N_2482,N_1592,N_1765);
nand U2483 (N_2483,N_1333,N_1354);
nor U2484 (N_2484,N_1248,N_1086);
xnor U2485 (N_2485,N_1159,N_1259);
nor U2486 (N_2486,N_1342,N_1014);
and U2487 (N_2487,N_1660,N_1543);
and U2488 (N_2488,N_1301,N_1130);
xnor U2489 (N_2489,N_1856,N_1535);
and U2490 (N_2490,N_1980,N_1883);
and U2491 (N_2491,N_1395,N_1528);
nor U2492 (N_2492,N_1570,N_1540);
and U2493 (N_2493,N_1160,N_1634);
or U2494 (N_2494,N_1052,N_1603);
nand U2495 (N_2495,N_1517,N_1442);
or U2496 (N_2496,N_1967,N_1909);
nor U2497 (N_2497,N_1853,N_1305);
or U2498 (N_2498,N_1396,N_1727);
and U2499 (N_2499,N_1247,N_1149);
or U2500 (N_2500,N_1990,N_1388);
nand U2501 (N_2501,N_1502,N_1602);
and U2502 (N_2502,N_1912,N_1009);
or U2503 (N_2503,N_1718,N_1720);
or U2504 (N_2504,N_1232,N_1017);
nand U2505 (N_2505,N_1750,N_1857);
nor U2506 (N_2506,N_1963,N_1692);
nor U2507 (N_2507,N_1988,N_1206);
or U2508 (N_2508,N_1438,N_1606);
and U2509 (N_2509,N_1957,N_1884);
nor U2510 (N_2510,N_1225,N_1750);
xnor U2511 (N_2511,N_1766,N_1683);
nand U2512 (N_2512,N_1004,N_1894);
nor U2513 (N_2513,N_1882,N_1939);
nand U2514 (N_2514,N_1796,N_1865);
nor U2515 (N_2515,N_1021,N_1663);
nor U2516 (N_2516,N_1201,N_1457);
or U2517 (N_2517,N_1207,N_1579);
and U2518 (N_2518,N_1839,N_1068);
nor U2519 (N_2519,N_1439,N_1867);
and U2520 (N_2520,N_1907,N_1366);
and U2521 (N_2521,N_1619,N_1649);
nand U2522 (N_2522,N_1076,N_1628);
nand U2523 (N_2523,N_1460,N_1329);
and U2524 (N_2524,N_1870,N_1025);
nand U2525 (N_2525,N_1195,N_1951);
nor U2526 (N_2526,N_1831,N_1667);
nor U2527 (N_2527,N_1169,N_1038);
and U2528 (N_2528,N_1160,N_1678);
nand U2529 (N_2529,N_1467,N_1054);
nand U2530 (N_2530,N_1709,N_1439);
nand U2531 (N_2531,N_1804,N_1972);
and U2532 (N_2532,N_1934,N_1976);
xor U2533 (N_2533,N_1880,N_1753);
nor U2534 (N_2534,N_1021,N_1685);
and U2535 (N_2535,N_1194,N_1090);
and U2536 (N_2536,N_1328,N_1128);
nor U2537 (N_2537,N_1028,N_1796);
nor U2538 (N_2538,N_1553,N_1936);
and U2539 (N_2539,N_1250,N_1209);
nand U2540 (N_2540,N_1015,N_1172);
nor U2541 (N_2541,N_1631,N_1973);
and U2542 (N_2542,N_1034,N_1161);
and U2543 (N_2543,N_1735,N_1975);
nand U2544 (N_2544,N_1977,N_1244);
nor U2545 (N_2545,N_1639,N_1053);
or U2546 (N_2546,N_1329,N_1935);
nand U2547 (N_2547,N_1366,N_1901);
nor U2548 (N_2548,N_1313,N_1995);
nand U2549 (N_2549,N_1344,N_1862);
or U2550 (N_2550,N_1143,N_1783);
and U2551 (N_2551,N_1041,N_1272);
nor U2552 (N_2552,N_1832,N_1604);
and U2553 (N_2553,N_1247,N_1883);
nand U2554 (N_2554,N_1595,N_1619);
nand U2555 (N_2555,N_1662,N_1485);
nor U2556 (N_2556,N_1239,N_1506);
xor U2557 (N_2557,N_1494,N_1892);
and U2558 (N_2558,N_1751,N_1080);
or U2559 (N_2559,N_1820,N_1040);
or U2560 (N_2560,N_1634,N_1343);
or U2561 (N_2561,N_1834,N_1909);
nand U2562 (N_2562,N_1036,N_1555);
or U2563 (N_2563,N_1915,N_1952);
xor U2564 (N_2564,N_1175,N_1958);
and U2565 (N_2565,N_1920,N_1221);
and U2566 (N_2566,N_1466,N_1456);
or U2567 (N_2567,N_1599,N_1541);
nor U2568 (N_2568,N_1964,N_1269);
and U2569 (N_2569,N_1555,N_1919);
or U2570 (N_2570,N_1624,N_1617);
and U2571 (N_2571,N_1036,N_1965);
nor U2572 (N_2572,N_1018,N_1822);
xor U2573 (N_2573,N_1437,N_1726);
and U2574 (N_2574,N_1856,N_1985);
and U2575 (N_2575,N_1262,N_1260);
and U2576 (N_2576,N_1593,N_1579);
nor U2577 (N_2577,N_1409,N_1570);
nor U2578 (N_2578,N_1316,N_1161);
nor U2579 (N_2579,N_1137,N_1500);
and U2580 (N_2580,N_1898,N_1996);
and U2581 (N_2581,N_1798,N_1096);
nor U2582 (N_2582,N_1802,N_1431);
and U2583 (N_2583,N_1765,N_1898);
nand U2584 (N_2584,N_1499,N_1360);
nand U2585 (N_2585,N_1271,N_1821);
nand U2586 (N_2586,N_1219,N_1814);
or U2587 (N_2587,N_1393,N_1146);
nor U2588 (N_2588,N_1133,N_1211);
and U2589 (N_2589,N_1192,N_1147);
or U2590 (N_2590,N_1097,N_1959);
nor U2591 (N_2591,N_1095,N_1197);
or U2592 (N_2592,N_1304,N_1591);
xor U2593 (N_2593,N_1301,N_1786);
nor U2594 (N_2594,N_1327,N_1205);
and U2595 (N_2595,N_1773,N_1294);
nand U2596 (N_2596,N_1234,N_1749);
nor U2597 (N_2597,N_1690,N_1139);
xnor U2598 (N_2598,N_1762,N_1162);
and U2599 (N_2599,N_1921,N_1367);
nand U2600 (N_2600,N_1502,N_1534);
nor U2601 (N_2601,N_1398,N_1542);
nand U2602 (N_2602,N_1576,N_1288);
nor U2603 (N_2603,N_1303,N_1350);
and U2604 (N_2604,N_1230,N_1449);
xnor U2605 (N_2605,N_1740,N_1313);
and U2606 (N_2606,N_1020,N_1000);
and U2607 (N_2607,N_1838,N_1786);
or U2608 (N_2608,N_1207,N_1717);
and U2609 (N_2609,N_1112,N_1513);
or U2610 (N_2610,N_1143,N_1268);
xor U2611 (N_2611,N_1142,N_1761);
nor U2612 (N_2612,N_1744,N_1173);
nand U2613 (N_2613,N_1785,N_1497);
nand U2614 (N_2614,N_1287,N_1736);
and U2615 (N_2615,N_1001,N_1330);
nand U2616 (N_2616,N_1414,N_1140);
or U2617 (N_2617,N_1014,N_1711);
and U2618 (N_2618,N_1281,N_1184);
or U2619 (N_2619,N_1673,N_1575);
and U2620 (N_2620,N_1314,N_1371);
xor U2621 (N_2621,N_1979,N_1629);
nand U2622 (N_2622,N_1581,N_1995);
or U2623 (N_2623,N_1359,N_1775);
xnor U2624 (N_2624,N_1894,N_1640);
or U2625 (N_2625,N_1197,N_1855);
nand U2626 (N_2626,N_1096,N_1655);
and U2627 (N_2627,N_1479,N_1732);
and U2628 (N_2628,N_1309,N_1244);
xor U2629 (N_2629,N_1676,N_1262);
and U2630 (N_2630,N_1443,N_1696);
or U2631 (N_2631,N_1590,N_1232);
nand U2632 (N_2632,N_1519,N_1459);
or U2633 (N_2633,N_1418,N_1779);
nand U2634 (N_2634,N_1508,N_1390);
and U2635 (N_2635,N_1289,N_1336);
or U2636 (N_2636,N_1610,N_1536);
nand U2637 (N_2637,N_1432,N_1338);
nand U2638 (N_2638,N_1641,N_1435);
and U2639 (N_2639,N_1530,N_1653);
and U2640 (N_2640,N_1412,N_1594);
nand U2641 (N_2641,N_1926,N_1431);
nor U2642 (N_2642,N_1337,N_1440);
or U2643 (N_2643,N_1028,N_1294);
nand U2644 (N_2644,N_1518,N_1958);
nand U2645 (N_2645,N_1985,N_1464);
nor U2646 (N_2646,N_1129,N_1287);
nand U2647 (N_2647,N_1603,N_1382);
nand U2648 (N_2648,N_1109,N_1364);
nor U2649 (N_2649,N_1393,N_1448);
nand U2650 (N_2650,N_1149,N_1117);
xor U2651 (N_2651,N_1408,N_1055);
and U2652 (N_2652,N_1279,N_1668);
nor U2653 (N_2653,N_1322,N_1915);
and U2654 (N_2654,N_1576,N_1575);
nor U2655 (N_2655,N_1831,N_1077);
nor U2656 (N_2656,N_1061,N_1087);
nor U2657 (N_2657,N_1852,N_1149);
or U2658 (N_2658,N_1932,N_1592);
nor U2659 (N_2659,N_1205,N_1961);
and U2660 (N_2660,N_1513,N_1046);
and U2661 (N_2661,N_1866,N_1760);
nand U2662 (N_2662,N_1206,N_1179);
or U2663 (N_2663,N_1319,N_1059);
nand U2664 (N_2664,N_1709,N_1412);
or U2665 (N_2665,N_1792,N_1277);
nor U2666 (N_2666,N_1158,N_1022);
nand U2667 (N_2667,N_1687,N_1550);
nand U2668 (N_2668,N_1659,N_1259);
and U2669 (N_2669,N_1328,N_1557);
and U2670 (N_2670,N_1795,N_1460);
nor U2671 (N_2671,N_1720,N_1978);
nor U2672 (N_2672,N_1673,N_1660);
xor U2673 (N_2673,N_1069,N_1100);
and U2674 (N_2674,N_1369,N_1042);
nand U2675 (N_2675,N_1995,N_1460);
xnor U2676 (N_2676,N_1651,N_1206);
and U2677 (N_2677,N_1812,N_1250);
or U2678 (N_2678,N_1843,N_1155);
nand U2679 (N_2679,N_1484,N_1103);
or U2680 (N_2680,N_1537,N_1148);
nor U2681 (N_2681,N_1107,N_1835);
and U2682 (N_2682,N_1282,N_1630);
nand U2683 (N_2683,N_1107,N_1996);
and U2684 (N_2684,N_1361,N_1046);
nor U2685 (N_2685,N_1897,N_1930);
nor U2686 (N_2686,N_1298,N_1386);
nor U2687 (N_2687,N_1057,N_1049);
nand U2688 (N_2688,N_1129,N_1744);
and U2689 (N_2689,N_1794,N_1173);
nand U2690 (N_2690,N_1988,N_1976);
or U2691 (N_2691,N_1976,N_1420);
or U2692 (N_2692,N_1686,N_1930);
and U2693 (N_2693,N_1824,N_1724);
nor U2694 (N_2694,N_1553,N_1543);
and U2695 (N_2695,N_1904,N_1718);
xor U2696 (N_2696,N_1622,N_1037);
or U2697 (N_2697,N_1805,N_1894);
xnor U2698 (N_2698,N_1687,N_1079);
or U2699 (N_2699,N_1156,N_1781);
and U2700 (N_2700,N_1507,N_1724);
or U2701 (N_2701,N_1181,N_1483);
nor U2702 (N_2702,N_1352,N_1532);
or U2703 (N_2703,N_1496,N_1130);
nand U2704 (N_2704,N_1575,N_1475);
nand U2705 (N_2705,N_1227,N_1608);
nor U2706 (N_2706,N_1629,N_1639);
or U2707 (N_2707,N_1931,N_1064);
and U2708 (N_2708,N_1596,N_1927);
and U2709 (N_2709,N_1293,N_1481);
and U2710 (N_2710,N_1495,N_1059);
and U2711 (N_2711,N_1323,N_1793);
nor U2712 (N_2712,N_1867,N_1544);
and U2713 (N_2713,N_1380,N_1141);
or U2714 (N_2714,N_1802,N_1094);
nor U2715 (N_2715,N_1730,N_1516);
nor U2716 (N_2716,N_1769,N_1800);
xnor U2717 (N_2717,N_1380,N_1144);
or U2718 (N_2718,N_1278,N_1124);
xnor U2719 (N_2719,N_1080,N_1621);
or U2720 (N_2720,N_1021,N_1559);
nand U2721 (N_2721,N_1576,N_1537);
or U2722 (N_2722,N_1726,N_1975);
nor U2723 (N_2723,N_1149,N_1658);
nand U2724 (N_2724,N_1356,N_1666);
nor U2725 (N_2725,N_1003,N_1927);
nor U2726 (N_2726,N_1512,N_1920);
or U2727 (N_2727,N_1027,N_1564);
and U2728 (N_2728,N_1227,N_1188);
nand U2729 (N_2729,N_1862,N_1940);
or U2730 (N_2730,N_1000,N_1003);
or U2731 (N_2731,N_1947,N_1365);
and U2732 (N_2732,N_1921,N_1157);
or U2733 (N_2733,N_1589,N_1342);
and U2734 (N_2734,N_1419,N_1500);
nor U2735 (N_2735,N_1091,N_1762);
or U2736 (N_2736,N_1199,N_1262);
nand U2737 (N_2737,N_1398,N_1496);
nor U2738 (N_2738,N_1090,N_1333);
or U2739 (N_2739,N_1170,N_1179);
and U2740 (N_2740,N_1553,N_1962);
nor U2741 (N_2741,N_1001,N_1329);
xor U2742 (N_2742,N_1672,N_1506);
or U2743 (N_2743,N_1897,N_1146);
nand U2744 (N_2744,N_1145,N_1944);
and U2745 (N_2745,N_1009,N_1338);
nor U2746 (N_2746,N_1831,N_1811);
and U2747 (N_2747,N_1994,N_1643);
xnor U2748 (N_2748,N_1744,N_1778);
or U2749 (N_2749,N_1484,N_1056);
or U2750 (N_2750,N_1059,N_1154);
or U2751 (N_2751,N_1667,N_1502);
or U2752 (N_2752,N_1846,N_1067);
nor U2753 (N_2753,N_1130,N_1900);
nand U2754 (N_2754,N_1121,N_1404);
xnor U2755 (N_2755,N_1588,N_1813);
and U2756 (N_2756,N_1887,N_1700);
nor U2757 (N_2757,N_1151,N_1928);
xor U2758 (N_2758,N_1801,N_1441);
nand U2759 (N_2759,N_1117,N_1129);
nor U2760 (N_2760,N_1153,N_1986);
nand U2761 (N_2761,N_1791,N_1886);
or U2762 (N_2762,N_1409,N_1661);
nor U2763 (N_2763,N_1013,N_1913);
nor U2764 (N_2764,N_1675,N_1728);
or U2765 (N_2765,N_1621,N_1040);
or U2766 (N_2766,N_1475,N_1644);
or U2767 (N_2767,N_1940,N_1801);
or U2768 (N_2768,N_1926,N_1948);
nor U2769 (N_2769,N_1494,N_1094);
xor U2770 (N_2770,N_1651,N_1382);
or U2771 (N_2771,N_1628,N_1684);
and U2772 (N_2772,N_1105,N_1945);
or U2773 (N_2773,N_1299,N_1803);
nor U2774 (N_2774,N_1523,N_1544);
nor U2775 (N_2775,N_1202,N_1808);
nor U2776 (N_2776,N_1936,N_1371);
or U2777 (N_2777,N_1514,N_1587);
and U2778 (N_2778,N_1636,N_1253);
nor U2779 (N_2779,N_1501,N_1258);
or U2780 (N_2780,N_1102,N_1836);
and U2781 (N_2781,N_1663,N_1672);
nor U2782 (N_2782,N_1259,N_1647);
xor U2783 (N_2783,N_1982,N_1144);
and U2784 (N_2784,N_1204,N_1890);
and U2785 (N_2785,N_1136,N_1033);
and U2786 (N_2786,N_1709,N_1134);
or U2787 (N_2787,N_1270,N_1372);
xor U2788 (N_2788,N_1016,N_1524);
nand U2789 (N_2789,N_1449,N_1729);
xnor U2790 (N_2790,N_1977,N_1252);
nor U2791 (N_2791,N_1741,N_1845);
nor U2792 (N_2792,N_1202,N_1130);
and U2793 (N_2793,N_1210,N_1289);
nor U2794 (N_2794,N_1369,N_1184);
and U2795 (N_2795,N_1755,N_1415);
nor U2796 (N_2796,N_1499,N_1309);
and U2797 (N_2797,N_1171,N_1842);
nor U2798 (N_2798,N_1837,N_1749);
nand U2799 (N_2799,N_1406,N_1610);
or U2800 (N_2800,N_1219,N_1948);
and U2801 (N_2801,N_1400,N_1466);
or U2802 (N_2802,N_1425,N_1446);
or U2803 (N_2803,N_1467,N_1184);
nand U2804 (N_2804,N_1589,N_1581);
nor U2805 (N_2805,N_1787,N_1851);
nor U2806 (N_2806,N_1839,N_1955);
xor U2807 (N_2807,N_1827,N_1856);
and U2808 (N_2808,N_1537,N_1157);
nand U2809 (N_2809,N_1463,N_1911);
nand U2810 (N_2810,N_1627,N_1636);
nor U2811 (N_2811,N_1272,N_1504);
xor U2812 (N_2812,N_1895,N_1733);
nand U2813 (N_2813,N_1311,N_1770);
or U2814 (N_2814,N_1816,N_1726);
nand U2815 (N_2815,N_1453,N_1870);
and U2816 (N_2816,N_1252,N_1973);
or U2817 (N_2817,N_1799,N_1426);
nand U2818 (N_2818,N_1458,N_1675);
xnor U2819 (N_2819,N_1351,N_1062);
or U2820 (N_2820,N_1806,N_1344);
and U2821 (N_2821,N_1277,N_1370);
and U2822 (N_2822,N_1949,N_1534);
nor U2823 (N_2823,N_1129,N_1412);
and U2824 (N_2824,N_1013,N_1780);
nor U2825 (N_2825,N_1644,N_1902);
nand U2826 (N_2826,N_1215,N_1539);
nand U2827 (N_2827,N_1152,N_1883);
nand U2828 (N_2828,N_1578,N_1701);
nand U2829 (N_2829,N_1893,N_1675);
xor U2830 (N_2830,N_1815,N_1922);
or U2831 (N_2831,N_1117,N_1454);
xor U2832 (N_2832,N_1116,N_1486);
or U2833 (N_2833,N_1395,N_1291);
nor U2834 (N_2834,N_1791,N_1355);
nor U2835 (N_2835,N_1423,N_1822);
or U2836 (N_2836,N_1610,N_1376);
or U2837 (N_2837,N_1804,N_1147);
or U2838 (N_2838,N_1244,N_1412);
and U2839 (N_2839,N_1330,N_1399);
or U2840 (N_2840,N_1898,N_1955);
and U2841 (N_2841,N_1731,N_1719);
nand U2842 (N_2842,N_1059,N_1149);
or U2843 (N_2843,N_1361,N_1013);
nor U2844 (N_2844,N_1012,N_1633);
nand U2845 (N_2845,N_1877,N_1747);
nand U2846 (N_2846,N_1279,N_1679);
and U2847 (N_2847,N_1840,N_1635);
and U2848 (N_2848,N_1764,N_1194);
or U2849 (N_2849,N_1735,N_1426);
nor U2850 (N_2850,N_1014,N_1515);
nand U2851 (N_2851,N_1506,N_1040);
nand U2852 (N_2852,N_1713,N_1402);
nand U2853 (N_2853,N_1990,N_1496);
and U2854 (N_2854,N_1771,N_1921);
nand U2855 (N_2855,N_1842,N_1077);
and U2856 (N_2856,N_1196,N_1398);
and U2857 (N_2857,N_1480,N_1715);
and U2858 (N_2858,N_1023,N_1549);
nand U2859 (N_2859,N_1589,N_1349);
nand U2860 (N_2860,N_1186,N_1226);
nand U2861 (N_2861,N_1104,N_1112);
xnor U2862 (N_2862,N_1859,N_1228);
nor U2863 (N_2863,N_1753,N_1997);
nand U2864 (N_2864,N_1245,N_1226);
xor U2865 (N_2865,N_1394,N_1355);
or U2866 (N_2866,N_1601,N_1057);
nor U2867 (N_2867,N_1626,N_1432);
nor U2868 (N_2868,N_1144,N_1299);
and U2869 (N_2869,N_1009,N_1579);
and U2870 (N_2870,N_1632,N_1349);
nor U2871 (N_2871,N_1475,N_1442);
nor U2872 (N_2872,N_1048,N_1418);
or U2873 (N_2873,N_1003,N_1431);
or U2874 (N_2874,N_1687,N_1795);
nand U2875 (N_2875,N_1394,N_1372);
and U2876 (N_2876,N_1565,N_1486);
nor U2877 (N_2877,N_1709,N_1335);
and U2878 (N_2878,N_1206,N_1059);
nor U2879 (N_2879,N_1106,N_1703);
and U2880 (N_2880,N_1441,N_1008);
or U2881 (N_2881,N_1791,N_1670);
or U2882 (N_2882,N_1420,N_1865);
nand U2883 (N_2883,N_1485,N_1516);
nand U2884 (N_2884,N_1451,N_1529);
nor U2885 (N_2885,N_1165,N_1622);
and U2886 (N_2886,N_1935,N_1904);
xnor U2887 (N_2887,N_1594,N_1093);
or U2888 (N_2888,N_1319,N_1566);
nand U2889 (N_2889,N_1781,N_1010);
or U2890 (N_2890,N_1404,N_1043);
and U2891 (N_2891,N_1465,N_1517);
xor U2892 (N_2892,N_1364,N_1880);
and U2893 (N_2893,N_1781,N_1642);
and U2894 (N_2894,N_1719,N_1203);
nor U2895 (N_2895,N_1853,N_1590);
and U2896 (N_2896,N_1799,N_1963);
or U2897 (N_2897,N_1128,N_1315);
or U2898 (N_2898,N_1752,N_1550);
and U2899 (N_2899,N_1059,N_1130);
or U2900 (N_2900,N_1014,N_1500);
nor U2901 (N_2901,N_1361,N_1328);
nand U2902 (N_2902,N_1585,N_1418);
nor U2903 (N_2903,N_1373,N_1306);
and U2904 (N_2904,N_1256,N_1621);
nor U2905 (N_2905,N_1328,N_1260);
and U2906 (N_2906,N_1102,N_1828);
and U2907 (N_2907,N_1219,N_1421);
and U2908 (N_2908,N_1508,N_1327);
and U2909 (N_2909,N_1576,N_1121);
nor U2910 (N_2910,N_1904,N_1113);
xor U2911 (N_2911,N_1568,N_1107);
nand U2912 (N_2912,N_1208,N_1655);
nand U2913 (N_2913,N_1052,N_1818);
nor U2914 (N_2914,N_1016,N_1325);
or U2915 (N_2915,N_1654,N_1864);
or U2916 (N_2916,N_1766,N_1154);
nor U2917 (N_2917,N_1252,N_1231);
nor U2918 (N_2918,N_1117,N_1407);
nand U2919 (N_2919,N_1456,N_1624);
and U2920 (N_2920,N_1874,N_1317);
xnor U2921 (N_2921,N_1425,N_1129);
xor U2922 (N_2922,N_1770,N_1036);
or U2923 (N_2923,N_1230,N_1428);
or U2924 (N_2924,N_1691,N_1577);
nand U2925 (N_2925,N_1786,N_1420);
nand U2926 (N_2926,N_1926,N_1131);
nand U2927 (N_2927,N_1496,N_1697);
and U2928 (N_2928,N_1786,N_1645);
xor U2929 (N_2929,N_1503,N_1872);
or U2930 (N_2930,N_1106,N_1133);
or U2931 (N_2931,N_1984,N_1079);
xor U2932 (N_2932,N_1156,N_1593);
and U2933 (N_2933,N_1274,N_1990);
nor U2934 (N_2934,N_1411,N_1153);
or U2935 (N_2935,N_1393,N_1240);
xnor U2936 (N_2936,N_1204,N_1537);
nand U2937 (N_2937,N_1012,N_1723);
nor U2938 (N_2938,N_1561,N_1417);
nand U2939 (N_2939,N_1135,N_1202);
or U2940 (N_2940,N_1810,N_1152);
and U2941 (N_2941,N_1147,N_1200);
and U2942 (N_2942,N_1891,N_1000);
and U2943 (N_2943,N_1844,N_1089);
nand U2944 (N_2944,N_1190,N_1057);
nor U2945 (N_2945,N_1913,N_1360);
nor U2946 (N_2946,N_1085,N_1335);
and U2947 (N_2947,N_1282,N_1513);
and U2948 (N_2948,N_1600,N_1805);
nand U2949 (N_2949,N_1885,N_1939);
nor U2950 (N_2950,N_1980,N_1995);
and U2951 (N_2951,N_1616,N_1549);
and U2952 (N_2952,N_1479,N_1526);
and U2953 (N_2953,N_1751,N_1317);
or U2954 (N_2954,N_1208,N_1308);
nand U2955 (N_2955,N_1172,N_1096);
nor U2956 (N_2956,N_1093,N_1718);
and U2957 (N_2957,N_1900,N_1414);
and U2958 (N_2958,N_1989,N_1302);
nor U2959 (N_2959,N_1316,N_1270);
nor U2960 (N_2960,N_1240,N_1291);
xnor U2961 (N_2961,N_1993,N_1698);
or U2962 (N_2962,N_1357,N_1811);
and U2963 (N_2963,N_1256,N_1838);
xnor U2964 (N_2964,N_1543,N_1163);
xor U2965 (N_2965,N_1774,N_1046);
and U2966 (N_2966,N_1875,N_1271);
or U2967 (N_2967,N_1158,N_1496);
nand U2968 (N_2968,N_1142,N_1893);
nand U2969 (N_2969,N_1927,N_1212);
xnor U2970 (N_2970,N_1972,N_1498);
nor U2971 (N_2971,N_1804,N_1513);
xnor U2972 (N_2972,N_1078,N_1477);
or U2973 (N_2973,N_1404,N_1653);
or U2974 (N_2974,N_1357,N_1753);
nand U2975 (N_2975,N_1855,N_1106);
and U2976 (N_2976,N_1033,N_1376);
xnor U2977 (N_2977,N_1074,N_1780);
nor U2978 (N_2978,N_1265,N_1936);
and U2979 (N_2979,N_1329,N_1310);
or U2980 (N_2980,N_1404,N_1557);
and U2981 (N_2981,N_1763,N_1468);
nor U2982 (N_2982,N_1083,N_1132);
nand U2983 (N_2983,N_1091,N_1258);
nor U2984 (N_2984,N_1289,N_1116);
and U2985 (N_2985,N_1849,N_1705);
and U2986 (N_2986,N_1524,N_1324);
or U2987 (N_2987,N_1652,N_1381);
nand U2988 (N_2988,N_1137,N_1080);
xor U2989 (N_2989,N_1908,N_1601);
and U2990 (N_2990,N_1227,N_1352);
or U2991 (N_2991,N_1813,N_1443);
nor U2992 (N_2992,N_1490,N_1059);
nor U2993 (N_2993,N_1990,N_1704);
nand U2994 (N_2994,N_1605,N_1344);
nor U2995 (N_2995,N_1181,N_1085);
or U2996 (N_2996,N_1906,N_1329);
xor U2997 (N_2997,N_1290,N_1438);
nor U2998 (N_2998,N_1432,N_1149);
or U2999 (N_2999,N_1250,N_1393);
or U3000 (N_3000,N_2740,N_2142);
and U3001 (N_3001,N_2933,N_2160);
and U3002 (N_3002,N_2102,N_2758);
xor U3003 (N_3003,N_2387,N_2959);
nor U3004 (N_3004,N_2461,N_2477);
nand U3005 (N_3005,N_2549,N_2358);
nand U3006 (N_3006,N_2256,N_2576);
and U3007 (N_3007,N_2130,N_2333);
nand U3008 (N_3008,N_2242,N_2109);
and U3009 (N_3009,N_2071,N_2023);
nor U3010 (N_3010,N_2121,N_2619);
or U3011 (N_3011,N_2797,N_2480);
and U3012 (N_3012,N_2006,N_2575);
and U3013 (N_3013,N_2631,N_2572);
and U3014 (N_3014,N_2923,N_2170);
nor U3015 (N_3015,N_2562,N_2354);
and U3016 (N_3016,N_2326,N_2093);
xor U3017 (N_3017,N_2069,N_2731);
nor U3018 (N_3018,N_2329,N_2537);
or U3019 (N_3019,N_2310,N_2513);
or U3020 (N_3020,N_2807,N_2581);
nor U3021 (N_3021,N_2820,N_2827);
and U3022 (N_3022,N_2189,N_2486);
xor U3023 (N_3023,N_2272,N_2205);
or U3024 (N_3024,N_2482,N_2510);
nor U3025 (N_3025,N_2196,N_2384);
xnor U3026 (N_3026,N_2896,N_2120);
nand U3027 (N_3027,N_2678,N_2367);
nor U3028 (N_3028,N_2173,N_2290);
and U3029 (N_3029,N_2693,N_2249);
or U3030 (N_3030,N_2536,N_2532);
nor U3031 (N_3031,N_2008,N_2348);
nand U3032 (N_3032,N_2592,N_2941);
nand U3033 (N_3033,N_2202,N_2296);
and U3034 (N_3034,N_2190,N_2483);
nor U3035 (N_3035,N_2314,N_2541);
or U3036 (N_3036,N_2435,N_2110);
nand U3037 (N_3037,N_2894,N_2517);
nand U3038 (N_3038,N_2845,N_2889);
and U3039 (N_3039,N_2825,N_2369);
nor U3040 (N_3040,N_2129,N_2975);
and U3041 (N_3041,N_2945,N_2357);
nand U3042 (N_3042,N_2388,N_2317);
or U3043 (N_3043,N_2223,N_2735);
or U3044 (N_3044,N_2749,N_2640);
nand U3045 (N_3045,N_2706,N_2690);
nor U3046 (N_3046,N_2016,N_2607);
and U3047 (N_3047,N_2542,N_2049);
nand U3048 (N_3048,N_2606,N_2824);
xor U3049 (N_3049,N_2647,N_2504);
nand U3050 (N_3050,N_2495,N_2704);
xor U3051 (N_3051,N_2839,N_2065);
nor U3052 (N_3052,N_2230,N_2446);
or U3053 (N_3053,N_2765,N_2238);
nand U3054 (N_3054,N_2702,N_2382);
nor U3055 (N_3055,N_2309,N_2267);
and U3056 (N_3056,N_2083,N_2692);
and U3057 (N_3057,N_2087,N_2815);
or U3058 (N_3058,N_2750,N_2756);
and U3059 (N_3059,N_2315,N_2375);
nand U3060 (N_3060,N_2403,N_2588);
nand U3061 (N_3061,N_2208,N_2791);
and U3062 (N_3062,N_2641,N_2928);
nand U3063 (N_3063,N_2836,N_2224);
and U3064 (N_3064,N_2302,N_2970);
nand U3065 (N_3065,N_2359,N_2268);
or U3066 (N_3066,N_2343,N_2535);
nor U3067 (N_3067,N_2801,N_2968);
nand U3068 (N_3068,N_2991,N_2009);
and U3069 (N_3069,N_2436,N_2018);
nand U3070 (N_3070,N_2848,N_2940);
nor U3071 (N_3071,N_2241,N_2186);
nand U3072 (N_3072,N_2099,N_2442);
or U3073 (N_3073,N_2610,N_2322);
or U3074 (N_3074,N_2492,N_2448);
and U3075 (N_3075,N_2045,N_2644);
xor U3076 (N_3076,N_2728,N_2897);
and U3077 (N_3077,N_2283,N_2877);
or U3078 (N_3078,N_2462,N_2344);
nor U3079 (N_3079,N_2291,N_2155);
nor U3080 (N_3080,N_2299,N_2028);
nand U3081 (N_3081,N_2162,N_2490);
and U3082 (N_3082,N_2273,N_2425);
nor U3083 (N_3083,N_2307,N_2349);
nand U3084 (N_3084,N_2932,N_2404);
nand U3085 (N_3085,N_2761,N_2112);
and U3086 (N_3086,N_2324,N_2421);
nand U3087 (N_3087,N_2199,N_2091);
and U3088 (N_3088,N_2379,N_2034);
and U3089 (N_3089,N_2134,N_2040);
nand U3090 (N_3090,N_2946,N_2882);
nand U3091 (N_3091,N_2287,N_2598);
nor U3092 (N_3092,N_2488,N_2769);
nand U3093 (N_3093,N_2833,N_2188);
and U3094 (N_3094,N_2659,N_2271);
and U3095 (N_3095,N_2381,N_2440);
and U3096 (N_3096,N_2067,N_2548);
nor U3097 (N_3097,N_2392,N_2509);
or U3098 (N_3098,N_2989,N_2499);
and U3099 (N_3099,N_2340,N_2958);
nand U3100 (N_3100,N_2980,N_2987);
nor U3101 (N_3101,N_2696,N_2601);
and U3102 (N_3102,N_2543,N_2117);
or U3103 (N_3103,N_2507,N_2802);
nand U3104 (N_3104,N_2194,N_2540);
nor U3105 (N_3105,N_2497,N_2579);
nor U3106 (N_3106,N_2195,N_2954);
or U3107 (N_3107,N_2853,N_2675);
and U3108 (N_3108,N_2565,N_2926);
or U3109 (N_3109,N_2685,N_2417);
and U3110 (N_3110,N_2757,N_2676);
and U3111 (N_3111,N_2679,N_2491);
or U3112 (N_3112,N_2805,N_2337);
nand U3113 (N_3113,N_2145,N_2747);
nor U3114 (N_3114,N_2365,N_2856);
or U3115 (N_3115,N_2213,N_2452);
and U3116 (N_3116,N_2161,N_2526);
and U3117 (N_3117,N_2570,N_2867);
nor U3118 (N_3118,N_2220,N_2981);
and U3119 (N_3119,N_2364,N_2180);
nand U3120 (N_3120,N_2335,N_2064);
and U3121 (N_3121,N_2868,N_2808);
nand U3122 (N_3122,N_2870,N_2103);
nor U3123 (N_3123,N_2764,N_2128);
nand U3124 (N_3124,N_2261,N_2029);
nor U3125 (N_3125,N_2460,N_2264);
or U3126 (N_3126,N_2864,N_2396);
nor U3127 (N_3127,N_2438,N_2332);
and U3128 (N_3128,N_2687,N_2269);
and U3129 (N_3129,N_2245,N_2350);
nand U3130 (N_3130,N_2547,N_2809);
or U3131 (N_3131,N_2432,N_2092);
nor U3132 (N_3132,N_2754,N_2789);
or U3133 (N_3133,N_2445,N_2346);
nand U3134 (N_3134,N_2639,N_2783);
xnor U3135 (N_3135,N_2697,N_2304);
or U3136 (N_3136,N_2015,N_2829);
and U3137 (N_3137,N_2533,N_2921);
nor U3138 (N_3138,N_2101,N_2650);
nand U3139 (N_3139,N_2165,N_2823);
or U3140 (N_3140,N_2591,N_2605);
nand U3141 (N_3141,N_2026,N_2111);
nor U3142 (N_3142,N_2903,N_2506);
or U3143 (N_3143,N_2280,N_2297);
or U3144 (N_3144,N_2203,N_2984);
or U3145 (N_3145,N_2527,N_2722);
nand U3146 (N_3146,N_2686,N_2587);
xor U3147 (N_3147,N_2792,N_2669);
nor U3148 (N_3148,N_2390,N_2622);
nand U3149 (N_3149,N_2219,N_2412);
nor U3150 (N_3150,N_2760,N_2044);
nand U3151 (N_3151,N_2965,N_2100);
nor U3152 (N_3152,N_2885,N_2586);
nand U3153 (N_3153,N_2398,N_2990);
nor U3154 (N_3154,N_2455,N_2393);
nor U3155 (N_3155,N_2115,N_2996);
nand U3156 (N_3156,N_2881,N_2131);
nand U3157 (N_3157,N_2627,N_2567);
or U3158 (N_3158,N_2192,N_2185);
or U3159 (N_3159,N_2779,N_2342);
nor U3160 (N_3160,N_2955,N_2937);
and U3161 (N_3161,N_2226,N_2002);
nor U3162 (N_3162,N_2376,N_2454);
or U3163 (N_3163,N_2961,N_2846);
nand U3164 (N_3164,N_2236,N_2806);
and U3165 (N_3165,N_2739,N_2655);
xor U3166 (N_3166,N_2368,N_2905);
nor U3167 (N_3167,N_2027,N_2775);
or U3168 (N_3168,N_2469,N_2252);
nand U3169 (N_3169,N_2400,N_2555);
nand U3170 (N_3170,N_2988,N_2434);
or U3171 (N_3171,N_2431,N_2152);
and U3172 (N_3172,N_2553,N_2206);
nand U3173 (N_3173,N_2918,N_2457);
or U3174 (N_3174,N_2094,N_2193);
nor U3175 (N_3175,N_2227,N_2574);
nor U3176 (N_3176,N_2132,N_2840);
nor U3177 (N_3177,N_2578,N_2584);
and U3178 (N_3178,N_2695,N_2748);
or U3179 (N_3179,N_2682,N_2726);
or U3180 (N_3180,N_2951,N_2214);
nand U3181 (N_3181,N_2244,N_2943);
and U3182 (N_3182,N_2727,N_2013);
xnor U3183 (N_3183,N_2135,N_2851);
or U3184 (N_3184,N_2514,N_2184);
and U3185 (N_3185,N_2508,N_2914);
and U3186 (N_3186,N_2487,N_2850);
and U3187 (N_3187,N_2589,N_2604);
and U3188 (N_3188,N_2544,N_2920);
xor U3189 (N_3189,N_2922,N_2661);
nor U3190 (N_3190,N_2437,N_2246);
nand U3191 (N_3191,N_2830,N_2096);
xnor U3192 (N_3192,N_2843,N_2855);
or U3193 (N_3193,N_2966,N_2258);
nor U3194 (N_3194,N_2127,N_2600);
or U3195 (N_3195,N_2125,N_2568);
or U3196 (N_3196,N_2931,N_2355);
xnor U3197 (N_3197,N_2858,N_2871);
and U3198 (N_3198,N_2391,N_2123);
nand U3199 (N_3199,N_2175,N_2869);
or U3200 (N_3200,N_2628,N_2772);
xor U3201 (N_3201,N_2734,N_2904);
or U3202 (N_3202,N_2637,N_2608);
nor U3203 (N_3203,N_2472,N_2828);
and U3204 (N_3204,N_2612,N_2420);
nor U3205 (N_3205,N_2422,N_2439);
or U3206 (N_3206,N_2849,N_2416);
and U3207 (N_3207,N_2119,N_2077);
and U3208 (N_3208,N_2814,N_2153);
xor U3209 (N_3209,N_2992,N_2339);
and U3210 (N_3210,N_2876,N_2285);
and U3211 (N_3211,N_2642,N_2694);
xor U3212 (N_3212,N_2530,N_2620);
nand U3213 (N_3213,N_2072,N_2211);
nor U3214 (N_3214,N_2771,N_2260);
nor U3215 (N_3215,N_2038,N_2892);
and U3216 (N_3216,N_2090,N_2745);
nand U3217 (N_3217,N_2552,N_2182);
and U3218 (N_3218,N_2944,N_2863);
nor U3219 (N_3219,N_2832,N_2380);
or U3220 (N_3220,N_2137,N_2776);
or U3221 (N_3221,N_2278,N_2216);
nand U3222 (N_3222,N_2397,N_2086);
or U3223 (N_3223,N_2585,N_2079);
and U3224 (N_3224,N_2478,N_2113);
and U3225 (N_3225,N_2459,N_2172);
and U3226 (N_3226,N_2969,N_2232);
xor U3227 (N_3227,N_2738,N_2635);
nor U3228 (N_3228,N_2209,N_2037);
nor U3229 (N_3229,N_2239,N_2798);
or U3230 (N_3230,N_2473,N_2515);
and U3231 (N_3231,N_2962,N_2781);
or U3232 (N_3232,N_2908,N_2957);
nor U3233 (N_3233,N_2073,N_2468);
and U3234 (N_3234,N_2902,N_2330);
and U3235 (N_3235,N_2235,N_2124);
xnor U3236 (N_3236,N_2680,N_2947);
nand U3237 (N_3237,N_2875,N_2122);
nor U3238 (N_3238,N_2020,N_2952);
and U3239 (N_3239,N_2512,N_2777);
or U3240 (N_3240,N_2561,N_2025);
xor U3241 (N_3241,N_2429,N_2636);
and U3242 (N_3242,N_2934,N_2353);
and U3243 (N_3243,N_2237,N_2259);
nand U3244 (N_3244,N_2837,N_2383);
nand U3245 (N_3245,N_2816,N_2024);
or U3246 (N_3246,N_2658,N_2564);
and U3247 (N_3247,N_2838,N_2321);
or U3248 (N_3248,N_2709,N_2788);
and U3249 (N_3249,N_2156,N_2325);
nand U3250 (N_3250,N_2688,N_2463);
and U3251 (N_3251,N_2062,N_2187);
nand U3252 (N_3252,N_2010,N_2418);
and U3253 (N_3253,N_2590,N_2061);
nand U3254 (N_3254,N_2505,N_2058);
and U3255 (N_3255,N_2629,N_2812);
nor U3256 (N_3256,N_2138,N_2786);
nand U3257 (N_3257,N_2386,N_2394);
nor U3258 (N_3258,N_2281,N_2972);
nor U3259 (N_3259,N_2767,N_2942);
or U3260 (N_3260,N_2546,N_2233);
nand U3261 (N_3261,N_2274,N_2915);
nor U3262 (N_3262,N_2423,N_2810);
or U3263 (N_3263,N_2859,N_2645);
nor U3264 (N_3264,N_2030,N_2046);
nand U3265 (N_3265,N_2899,N_2179);
and U3266 (N_3266,N_2108,N_2372);
nor U3267 (N_3267,N_2146,N_2293);
or U3268 (N_3268,N_2303,N_2294);
or U3269 (N_3269,N_2060,N_2312);
or U3270 (N_3270,N_2430,N_2419);
or U3271 (N_3271,N_2973,N_2519);
or U3272 (N_3272,N_2768,N_2467);
xnor U3273 (N_3273,N_2566,N_2698);
nor U3274 (N_3274,N_2878,N_2668);
and U3275 (N_3275,N_2385,N_2649);
nor U3276 (N_3276,N_2593,N_2634);
and U3277 (N_3277,N_2427,N_2999);
nand U3278 (N_3278,N_2913,N_2068);
and U3279 (N_3279,N_2074,N_2912);
or U3280 (N_3280,N_2523,N_2036);
nand U3281 (N_3281,N_2720,N_2399);
or U3282 (N_3282,N_2596,N_2470);
or U3283 (N_3283,N_2983,N_2677);
xnor U3284 (N_3284,N_2318,N_2097);
and U3285 (N_3285,N_2662,N_2599);
nor U3286 (N_3286,N_2821,N_2774);
nand U3287 (N_3287,N_2450,N_2700);
nand U3288 (N_3288,N_2204,N_2818);
nor U3289 (N_3289,N_2770,N_2978);
nand U3290 (N_3290,N_2231,N_2361);
and U3291 (N_3291,N_2052,N_2377);
nand U3292 (N_3292,N_2893,N_2744);
nand U3293 (N_3293,N_2907,N_2550);
nand U3294 (N_3294,N_2316,N_2177);
or U3295 (N_3295,N_2901,N_2718);
nand U3296 (N_3296,N_2277,N_2674);
and U3297 (N_3297,N_2181,N_2313);
and U3298 (N_3298,N_2298,N_2545);
and U3299 (N_3299,N_2614,N_2755);
nand U3300 (N_3300,N_2736,N_2976);
xor U3301 (N_3301,N_2625,N_2331);
nand U3302 (N_3302,N_2887,N_2279);
and U3303 (N_3303,N_2813,N_2699);
or U3304 (N_3304,N_2844,N_2852);
and U3305 (N_3305,N_2166,N_2133);
xor U3306 (N_3306,N_2088,N_2880);
or U3307 (N_3307,N_2557,N_2105);
nor U3308 (N_3308,N_2993,N_2451);
and U3309 (N_3309,N_2306,N_2493);
nor U3310 (N_3310,N_2898,N_2270);
nor U3311 (N_3311,N_2534,N_2803);
xor U3312 (N_3312,N_2684,N_2939);
nand U3313 (N_3313,N_2822,N_2019);
and U3314 (N_3314,N_2248,N_2615);
nor U3315 (N_3315,N_2703,N_2705);
xnor U3316 (N_3316,N_2539,N_2656);
nor U3317 (N_3317,N_2319,N_2282);
and U3318 (N_3318,N_2667,N_2995);
or U3319 (N_3319,N_2672,N_2405);
nor U3320 (N_3320,N_2558,N_2070);
or U3321 (N_3321,N_2444,N_2638);
xor U3322 (N_3322,N_2571,N_2410);
or U3323 (N_3323,N_2466,N_2149);
or U3324 (N_3324,N_2106,N_2085);
or U3325 (N_3325,N_2831,N_2626);
or U3326 (N_3326,N_2401,N_2799);
nor U3327 (N_3327,N_2865,N_2778);
or U3328 (N_3328,N_2288,N_2496);
nor U3329 (N_3329,N_2114,N_2967);
or U3330 (N_3330,N_2300,N_2790);
xor U3331 (N_3331,N_2327,N_2743);
and U3332 (N_3332,N_2407,N_2582);
or U3333 (N_3333,N_2250,N_2043);
or U3334 (N_3334,N_2178,N_2652);
and U3335 (N_3335,N_2078,N_2465);
nor U3336 (N_3336,N_2243,N_2753);
and U3337 (N_3337,N_2580,N_2719);
nor U3338 (N_3338,N_2151,N_2633);
xor U3339 (N_3339,N_2042,N_2787);
nand U3340 (N_3340,N_2453,N_2144);
nor U3341 (N_3341,N_2721,N_2708);
nand U3342 (N_3342,N_2360,N_2900);
nand U3343 (N_3343,N_2929,N_2484);
and U3344 (N_3344,N_2408,N_2413);
nor U3345 (N_3345,N_2215,N_2167);
and U3346 (N_3346,N_2035,N_2653);
or U3347 (N_3347,N_2012,N_2075);
nand U3348 (N_3348,N_2500,N_2481);
or U3349 (N_3349,N_2081,N_2691);
nor U3350 (N_3350,N_2977,N_2597);
and U3351 (N_3351,N_2964,N_2240);
or U3352 (N_3352,N_2860,N_2059);
nand U3353 (N_3353,N_2559,N_2053);
and U3354 (N_3354,N_2784,N_2560);
or U3355 (N_3355,N_2169,N_2573);
or U3356 (N_3356,N_2143,N_2041);
and U3357 (N_3357,N_2657,N_2311);
and U3358 (N_3358,N_2971,N_2936);
nand U3359 (N_3359,N_2594,N_2371);
and U3360 (N_3360,N_2411,N_2356);
and U3361 (N_3361,N_2683,N_2363);
or U3362 (N_3362,N_2201,N_2854);
and U3363 (N_3363,N_2646,N_2011);
nand U3364 (N_3364,N_2842,N_2960);
nor U3365 (N_3365,N_2433,N_2681);
nor U3366 (N_3366,N_2005,N_2107);
nor U3367 (N_3367,N_2866,N_2456);
and U3368 (N_3368,N_2047,N_2773);
nor U3369 (N_3369,N_2336,N_2054);
or U3370 (N_3370,N_2800,N_2255);
or U3371 (N_3371,N_2927,N_2874);
and U3372 (N_3372,N_2819,N_2338);
xnor U3373 (N_3373,N_2489,N_2479);
or U3374 (N_3374,N_2056,N_2729);
nand U3375 (N_3375,N_2632,N_2001);
nor U3376 (N_3376,N_2328,N_2762);
or U3377 (N_3377,N_2714,N_2910);
and U3378 (N_3378,N_2847,N_2895);
nand U3379 (N_3379,N_2630,N_2014);
nor U3380 (N_3380,N_2183,N_2725);
and U3381 (N_3381,N_2221,N_2458);
and U3382 (N_3382,N_2395,N_2292);
or U3383 (N_3383,N_2136,N_2811);
or U3384 (N_3384,N_2524,N_2730);
xor U3385 (N_3385,N_2406,N_2516);
or U3386 (N_3386,N_2985,N_2664);
nor U3387 (N_3387,N_2474,N_2289);
nor U3388 (N_3388,N_2441,N_2569);
or U3389 (N_3389,N_2168,N_2424);
nor U3390 (N_3390,N_2263,N_2717);
nor U3391 (N_3391,N_2886,N_2148);
nor U3392 (N_3392,N_2554,N_2370);
or U3393 (N_3393,N_2449,N_2994);
nand U3394 (N_3394,N_2785,N_2766);
nor U3395 (N_3395,N_2159,N_2948);
or U3396 (N_3396,N_2911,N_2793);
or U3397 (N_3397,N_2826,N_2301);
or U3398 (N_3398,N_2225,N_2663);
nor U3399 (N_3399,N_2055,N_2022);
nor U3400 (N_3400,N_2207,N_2795);
nand U3401 (N_3401,N_2518,N_2949);
nand U3402 (N_3402,N_2118,N_2884);
nor U3403 (N_3403,N_2879,N_2341);
nor U3404 (N_3404,N_2538,N_2050);
nor U3405 (N_3405,N_2345,N_2198);
nor U3406 (N_3406,N_2141,N_2521);
nand U3407 (N_3407,N_2503,N_2613);
nand U3408 (N_3408,N_2498,N_2017);
nand U3409 (N_3409,N_2443,N_2021);
and U3410 (N_3410,N_2323,N_2935);
xor U3411 (N_3411,N_2715,N_2531);
nor U3412 (N_3412,N_2873,N_2835);
and U3413 (N_3413,N_2689,N_2909);
or U3414 (N_3414,N_2426,N_2212);
nor U3415 (N_3415,N_2611,N_2305);
and U3416 (N_3416,N_2295,N_2616);
nand U3417 (N_3417,N_2701,N_2098);
nor U3418 (N_3418,N_2095,N_2475);
nand U3419 (N_3419,N_2228,N_2670);
and U3420 (N_3420,N_2782,N_2872);
nor U3421 (N_3421,N_2522,N_2171);
nand U3422 (N_3422,N_2751,N_2660);
or U3423 (N_3423,N_2602,N_2716);
and U3424 (N_3424,N_2986,N_2039);
or U3425 (N_3425,N_2621,N_2033);
or U3426 (N_3426,N_2485,N_2862);
xnor U3427 (N_3427,N_2057,N_2247);
nand U3428 (N_3428,N_2953,N_2415);
or U3429 (N_3429,N_2150,N_2471);
nor U3430 (N_3430,N_2126,N_2950);
or U3431 (N_3431,N_2502,N_2603);
nand U3432 (N_3432,N_2724,N_2003);
or U3433 (N_3433,N_2841,N_2956);
and U3434 (N_3434,N_2082,N_2080);
nor U3435 (N_3435,N_2938,N_2076);
or U3436 (N_3436,N_2609,N_2643);
nand U3437 (N_3437,N_2906,N_2742);
or U3438 (N_3438,N_2262,N_2528);
nor U3439 (N_3439,N_2711,N_2997);
nor U3440 (N_3440,N_2229,N_2266);
nor U3441 (N_3441,N_2378,N_2671);
nor U3442 (N_3442,N_2556,N_2191);
nand U3443 (N_3443,N_2409,N_2917);
xnor U3444 (N_3444,N_2891,N_2116);
nor U3445 (N_3445,N_2217,N_2804);
nor U3446 (N_3446,N_2362,N_2998);
nor U3447 (N_3447,N_2710,N_2374);
or U3448 (N_3448,N_2234,N_2031);
or U3449 (N_3449,N_2919,N_2794);
nand U3450 (N_3450,N_2796,N_2780);
nand U3451 (N_3451,N_2210,N_2032);
nand U3452 (N_3452,N_2000,N_2218);
or U3453 (N_3453,N_2551,N_2347);
nand U3454 (N_3454,N_2834,N_2974);
or U3455 (N_3455,N_2200,N_2737);
and U3456 (N_3456,N_2925,N_2732);
and U3457 (N_3457,N_2595,N_2617);
and U3458 (N_3458,N_2857,N_2254);
nand U3459 (N_3459,N_2174,N_2494);
and U3460 (N_3460,N_2624,N_2618);
or U3461 (N_3461,N_2366,N_2276);
nor U3462 (N_3462,N_2066,N_2648);
nor U3463 (N_3463,N_2890,N_2265);
and U3464 (N_3464,N_2577,N_2197);
nand U3465 (N_3465,N_2476,N_2651);
nor U3466 (N_3466,N_2752,N_2286);
and U3467 (N_3467,N_2712,N_2673);
nand U3468 (N_3468,N_2176,N_2089);
and U3469 (N_3469,N_2251,N_2414);
xnor U3470 (N_3470,N_2373,N_2979);
nor U3471 (N_3471,N_2147,N_2759);
nor U3472 (N_3472,N_2447,N_2352);
and U3473 (N_3473,N_2051,N_2520);
and U3474 (N_3474,N_2930,N_2275);
or U3475 (N_3475,N_2723,N_2746);
nor U3476 (N_3476,N_2861,N_2284);
nand U3477 (N_3477,N_2253,N_2164);
or U3478 (N_3478,N_2525,N_2916);
and U3479 (N_3479,N_2501,N_2707);
or U3480 (N_3480,N_2888,N_2763);
nor U3481 (N_3481,N_2817,N_2741);
and U3482 (N_3482,N_2428,N_2139);
and U3483 (N_3483,N_2048,N_2623);
xnor U3484 (N_3484,N_2154,N_2666);
nor U3485 (N_3485,N_2389,N_2464);
and U3486 (N_3486,N_2158,N_2257);
nand U3487 (N_3487,N_2654,N_2104);
nand U3488 (N_3488,N_2334,N_2163);
and U3489 (N_3489,N_2924,N_2733);
xor U3490 (N_3490,N_2222,N_2402);
nand U3491 (N_3491,N_2084,N_2320);
or U3492 (N_3492,N_2351,N_2563);
and U3493 (N_3493,N_2511,N_2963);
or U3494 (N_3494,N_2883,N_2529);
nor U3495 (N_3495,N_2308,N_2713);
and U3496 (N_3496,N_2665,N_2982);
nand U3497 (N_3497,N_2583,N_2004);
xor U3498 (N_3498,N_2157,N_2140);
and U3499 (N_3499,N_2063,N_2007);
and U3500 (N_3500,N_2100,N_2932);
or U3501 (N_3501,N_2759,N_2239);
nor U3502 (N_3502,N_2321,N_2228);
nand U3503 (N_3503,N_2614,N_2373);
or U3504 (N_3504,N_2938,N_2212);
nor U3505 (N_3505,N_2353,N_2443);
and U3506 (N_3506,N_2290,N_2818);
nand U3507 (N_3507,N_2799,N_2813);
nand U3508 (N_3508,N_2972,N_2938);
nand U3509 (N_3509,N_2763,N_2772);
and U3510 (N_3510,N_2352,N_2158);
and U3511 (N_3511,N_2851,N_2984);
or U3512 (N_3512,N_2702,N_2447);
and U3513 (N_3513,N_2134,N_2933);
or U3514 (N_3514,N_2302,N_2182);
nand U3515 (N_3515,N_2637,N_2656);
or U3516 (N_3516,N_2518,N_2761);
nor U3517 (N_3517,N_2751,N_2267);
nor U3518 (N_3518,N_2301,N_2516);
or U3519 (N_3519,N_2708,N_2354);
and U3520 (N_3520,N_2777,N_2275);
nor U3521 (N_3521,N_2616,N_2932);
or U3522 (N_3522,N_2299,N_2478);
xor U3523 (N_3523,N_2995,N_2732);
nand U3524 (N_3524,N_2933,N_2039);
nand U3525 (N_3525,N_2477,N_2271);
nor U3526 (N_3526,N_2473,N_2076);
nand U3527 (N_3527,N_2642,N_2175);
or U3528 (N_3528,N_2363,N_2314);
and U3529 (N_3529,N_2143,N_2049);
nand U3530 (N_3530,N_2241,N_2009);
and U3531 (N_3531,N_2887,N_2694);
or U3532 (N_3532,N_2455,N_2982);
nand U3533 (N_3533,N_2586,N_2578);
nand U3534 (N_3534,N_2702,N_2280);
nand U3535 (N_3535,N_2249,N_2922);
xor U3536 (N_3536,N_2881,N_2165);
nor U3537 (N_3537,N_2120,N_2854);
nand U3538 (N_3538,N_2827,N_2767);
xnor U3539 (N_3539,N_2748,N_2131);
or U3540 (N_3540,N_2024,N_2562);
nand U3541 (N_3541,N_2718,N_2700);
nor U3542 (N_3542,N_2091,N_2421);
or U3543 (N_3543,N_2432,N_2969);
xor U3544 (N_3544,N_2280,N_2011);
nand U3545 (N_3545,N_2018,N_2543);
or U3546 (N_3546,N_2588,N_2969);
and U3547 (N_3547,N_2639,N_2440);
xor U3548 (N_3548,N_2325,N_2181);
and U3549 (N_3549,N_2911,N_2031);
nor U3550 (N_3550,N_2539,N_2439);
nand U3551 (N_3551,N_2576,N_2859);
nor U3552 (N_3552,N_2788,N_2392);
or U3553 (N_3553,N_2962,N_2610);
and U3554 (N_3554,N_2372,N_2843);
and U3555 (N_3555,N_2916,N_2262);
and U3556 (N_3556,N_2849,N_2379);
nand U3557 (N_3557,N_2728,N_2144);
nand U3558 (N_3558,N_2639,N_2958);
and U3559 (N_3559,N_2923,N_2647);
or U3560 (N_3560,N_2141,N_2079);
nor U3561 (N_3561,N_2362,N_2723);
or U3562 (N_3562,N_2277,N_2844);
and U3563 (N_3563,N_2039,N_2446);
nor U3564 (N_3564,N_2156,N_2159);
nand U3565 (N_3565,N_2705,N_2437);
nand U3566 (N_3566,N_2644,N_2968);
or U3567 (N_3567,N_2041,N_2213);
and U3568 (N_3568,N_2270,N_2248);
nor U3569 (N_3569,N_2494,N_2048);
nor U3570 (N_3570,N_2740,N_2563);
nor U3571 (N_3571,N_2462,N_2157);
or U3572 (N_3572,N_2796,N_2349);
nor U3573 (N_3573,N_2785,N_2349);
nand U3574 (N_3574,N_2492,N_2895);
nor U3575 (N_3575,N_2460,N_2921);
or U3576 (N_3576,N_2495,N_2824);
xnor U3577 (N_3577,N_2189,N_2983);
nand U3578 (N_3578,N_2807,N_2959);
or U3579 (N_3579,N_2613,N_2248);
xnor U3580 (N_3580,N_2388,N_2500);
and U3581 (N_3581,N_2989,N_2310);
or U3582 (N_3582,N_2315,N_2101);
nor U3583 (N_3583,N_2904,N_2742);
nor U3584 (N_3584,N_2641,N_2008);
nand U3585 (N_3585,N_2802,N_2657);
nor U3586 (N_3586,N_2113,N_2766);
or U3587 (N_3587,N_2280,N_2068);
and U3588 (N_3588,N_2642,N_2132);
nand U3589 (N_3589,N_2710,N_2365);
and U3590 (N_3590,N_2841,N_2470);
nor U3591 (N_3591,N_2694,N_2428);
nand U3592 (N_3592,N_2704,N_2390);
or U3593 (N_3593,N_2721,N_2014);
and U3594 (N_3594,N_2874,N_2845);
and U3595 (N_3595,N_2379,N_2622);
or U3596 (N_3596,N_2324,N_2346);
and U3597 (N_3597,N_2070,N_2199);
and U3598 (N_3598,N_2881,N_2054);
nor U3599 (N_3599,N_2201,N_2678);
or U3600 (N_3600,N_2628,N_2970);
or U3601 (N_3601,N_2941,N_2638);
or U3602 (N_3602,N_2711,N_2797);
or U3603 (N_3603,N_2773,N_2376);
nand U3604 (N_3604,N_2111,N_2650);
and U3605 (N_3605,N_2494,N_2180);
nor U3606 (N_3606,N_2079,N_2286);
nand U3607 (N_3607,N_2675,N_2349);
and U3608 (N_3608,N_2331,N_2296);
nand U3609 (N_3609,N_2543,N_2682);
or U3610 (N_3610,N_2528,N_2236);
nor U3611 (N_3611,N_2273,N_2172);
and U3612 (N_3612,N_2885,N_2937);
and U3613 (N_3613,N_2389,N_2747);
and U3614 (N_3614,N_2504,N_2468);
xnor U3615 (N_3615,N_2377,N_2281);
nand U3616 (N_3616,N_2287,N_2678);
and U3617 (N_3617,N_2946,N_2413);
nor U3618 (N_3618,N_2715,N_2089);
nand U3619 (N_3619,N_2591,N_2066);
and U3620 (N_3620,N_2779,N_2858);
nor U3621 (N_3621,N_2450,N_2675);
and U3622 (N_3622,N_2916,N_2820);
nand U3623 (N_3623,N_2915,N_2909);
or U3624 (N_3624,N_2957,N_2796);
and U3625 (N_3625,N_2486,N_2873);
xnor U3626 (N_3626,N_2794,N_2588);
nand U3627 (N_3627,N_2556,N_2376);
nand U3628 (N_3628,N_2702,N_2957);
nand U3629 (N_3629,N_2687,N_2014);
and U3630 (N_3630,N_2761,N_2916);
or U3631 (N_3631,N_2905,N_2746);
and U3632 (N_3632,N_2104,N_2682);
nand U3633 (N_3633,N_2531,N_2616);
and U3634 (N_3634,N_2203,N_2040);
nor U3635 (N_3635,N_2661,N_2299);
and U3636 (N_3636,N_2246,N_2311);
and U3637 (N_3637,N_2015,N_2136);
nand U3638 (N_3638,N_2562,N_2998);
or U3639 (N_3639,N_2298,N_2581);
nand U3640 (N_3640,N_2877,N_2862);
or U3641 (N_3641,N_2532,N_2457);
nand U3642 (N_3642,N_2138,N_2048);
nor U3643 (N_3643,N_2474,N_2122);
nor U3644 (N_3644,N_2391,N_2775);
or U3645 (N_3645,N_2231,N_2738);
or U3646 (N_3646,N_2178,N_2670);
nand U3647 (N_3647,N_2576,N_2564);
xnor U3648 (N_3648,N_2072,N_2014);
nand U3649 (N_3649,N_2881,N_2760);
and U3650 (N_3650,N_2664,N_2695);
and U3651 (N_3651,N_2330,N_2767);
nor U3652 (N_3652,N_2902,N_2629);
nand U3653 (N_3653,N_2203,N_2233);
and U3654 (N_3654,N_2229,N_2141);
nor U3655 (N_3655,N_2859,N_2246);
nand U3656 (N_3656,N_2157,N_2521);
xnor U3657 (N_3657,N_2342,N_2699);
nor U3658 (N_3658,N_2674,N_2253);
and U3659 (N_3659,N_2817,N_2246);
or U3660 (N_3660,N_2084,N_2542);
nor U3661 (N_3661,N_2005,N_2364);
nand U3662 (N_3662,N_2585,N_2892);
or U3663 (N_3663,N_2092,N_2043);
nor U3664 (N_3664,N_2642,N_2044);
nor U3665 (N_3665,N_2020,N_2395);
xor U3666 (N_3666,N_2082,N_2862);
nand U3667 (N_3667,N_2742,N_2666);
nor U3668 (N_3668,N_2358,N_2087);
xor U3669 (N_3669,N_2760,N_2370);
nand U3670 (N_3670,N_2688,N_2109);
nor U3671 (N_3671,N_2015,N_2265);
nor U3672 (N_3672,N_2301,N_2080);
xor U3673 (N_3673,N_2515,N_2915);
and U3674 (N_3674,N_2722,N_2011);
and U3675 (N_3675,N_2026,N_2977);
or U3676 (N_3676,N_2904,N_2716);
nor U3677 (N_3677,N_2433,N_2321);
nand U3678 (N_3678,N_2476,N_2994);
nand U3679 (N_3679,N_2825,N_2575);
or U3680 (N_3680,N_2060,N_2285);
and U3681 (N_3681,N_2692,N_2319);
nand U3682 (N_3682,N_2548,N_2444);
nand U3683 (N_3683,N_2594,N_2287);
nand U3684 (N_3684,N_2797,N_2769);
nor U3685 (N_3685,N_2821,N_2347);
nand U3686 (N_3686,N_2293,N_2916);
or U3687 (N_3687,N_2781,N_2946);
or U3688 (N_3688,N_2230,N_2586);
nand U3689 (N_3689,N_2393,N_2672);
nor U3690 (N_3690,N_2564,N_2139);
and U3691 (N_3691,N_2726,N_2318);
and U3692 (N_3692,N_2885,N_2654);
xor U3693 (N_3693,N_2517,N_2553);
and U3694 (N_3694,N_2840,N_2214);
and U3695 (N_3695,N_2198,N_2740);
and U3696 (N_3696,N_2252,N_2534);
or U3697 (N_3697,N_2807,N_2545);
nor U3698 (N_3698,N_2213,N_2143);
nand U3699 (N_3699,N_2218,N_2471);
nor U3700 (N_3700,N_2873,N_2379);
or U3701 (N_3701,N_2829,N_2534);
or U3702 (N_3702,N_2978,N_2675);
and U3703 (N_3703,N_2156,N_2783);
nand U3704 (N_3704,N_2758,N_2310);
and U3705 (N_3705,N_2075,N_2510);
and U3706 (N_3706,N_2293,N_2447);
nor U3707 (N_3707,N_2525,N_2668);
nand U3708 (N_3708,N_2083,N_2384);
xor U3709 (N_3709,N_2257,N_2119);
xnor U3710 (N_3710,N_2893,N_2971);
nand U3711 (N_3711,N_2842,N_2066);
and U3712 (N_3712,N_2798,N_2500);
nor U3713 (N_3713,N_2679,N_2994);
nand U3714 (N_3714,N_2969,N_2853);
and U3715 (N_3715,N_2541,N_2224);
and U3716 (N_3716,N_2619,N_2316);
or U3717 (N_3717,N_2889,N_2225);
or U3718 (N_3718,N_2118,N_2166);
nor U3719 (N_3719,N_2840,N_2808);
nand U3720 (N_3720,N_2025,N_2856);
xor U3721 (N_3721,N_2478,N_2823);
nand U3722 (N_3722,N_2176,N_2978);
or U3723 (N_3723,N_2058,N_2053);
nand U3724 (N_3724,N_2552,N_2232);
nor U3725 (N_3725,N_2559,N_2401);
and U3726 (N_3726,N_2552,N_2611);
nand U3727 (N_3727,N_2733,N_2358);
nor U3728 (N_3728,N_2583,N_2477);
nor U3729 (N_3729,N_2520,N_2420);
nor U3730 (N_3730,N_2107,N_2583);
xnor U3731 (N_3731,N_2322,N_2024);
or U3732 (N_3732,N_2045,N_2757);
nor U3733 (N_3733,N_2733,N_2740);
nor U3734 (N_3734,N_2577,N_2462);
nor U3735 (N_3735,N_2974,N_2003);
xnor U3736 (N_3736,N_2951,N_2694);
or U3737 (N_3737,N_2334,N_2409);
nor U3738 (N_3738,N_2952,N_2588);
and U3739 (N_3739,N_2190,N_2923);
nand U3740 (N_3740,N_2800,N_2631);
nor U3741 (N_3741,N_2415,N_2276);
nand U3742 (N_3742,N_2725,N_2674);
nand U3743 (N_3743,N_2531,N_2472);
nor U3744 (N_3744,N_2936,N_2715);
xnor U3745 (N_3745,N_2715,N_2004);
nand U3746 (N_3746,N_2420,N_2316);
nand U3747 (N_3747,N_2327,N_2285);
xnor U3748 (N_3748,N_2985,N_2108);
xnor U3749 (N_3749,N_2379,N_2446);
nor U3750 (N_3750,N_2025,N_2271);
and U3751 (N_3751,N_2769,N_2333);
nor U3752 (N_3752,N_2941,N_2337);
xor U3753 (N_3753,N_2495,N_2864);
or U3754 (N_3754,N_2100,N_2840);
or U3755 (N_3755,N_2368,N_2766);
xor U3756 (N_3756,N_2238,N_2886);
xnor U3757 (N_3757,N_2821,N_2460);
nand U3758 (N_3758,N_2073,N_2727);
or U3759 (N_3759,N_2355,N_2781);
or U3760 (N_3760,N_2276,N_2801);
nand U3761 (N_3761,N_2732,N_2551);
nor U3762 (N_3762,N_2076,N_2096);
nand U3763 (N_3763,N_2893,N_2072);
nand U3764 (N_3764,N_2307,N_2075);
and U3765 (N_3765,N_2137,N_2643);
or U3766 (N_3766,N_2453,N_2913);
or U3767 (N_3767,N_2483,N_2979);
nand U3768 (N_3768,N_2505,N_2322);
nor U3769 (N_3769,N_2213,N_2979);
nor U3770 (N_3770,N_2170,N_2011);
nand U3771 (N_3771,N_2873,N_2523);
nand U3772 (N_3772,N_2473,N_2141);
nor U3773 (N_3773,N_2490,N_2280);
nand U3774 (N_3774,N_2936,N_2011);
nor U3775 (N_3775,N_2801,N_2095);
nor U3776 (N_3776,N_2943,N_2872);
xor U3777 (N_3777,N_2270,N_2189);
nor U3778 (N_3778,N_2772,N_2306);
or U3779 (N_3779,N_2067,N_2102);
or U3780 (N_3780,N_2328,N_2306);
nand U3781 (N_3781,N_2030,N_2584);
or U3782 (N_3782,N_2663,N_2570);
xor U3783 (N_3783,N_2338,N_2908);
nor U3784 (N_3784,N_2576,N_2639);
nor U3785 (N_3785,N_2165,N_2216);
nor U3786 (N_3786,N_2956,N_2567);
and U3787 (N_3787,N_2133,N_2460);
nor U3788 (N_3788,N_2872,N_2842);
nand U3789 (N_3789,N_2346,N_2734);
xor U3790 (N_3790,N_2932,N_2542);
and U3791 (N_3791,N_2301,N_2458);
and U3792 (N_3792,N_2521,N_2656);
nand U3793 (N_3793,N_2853,N_2236);
and U3794 (N_3794,N_2985,N_2609);
and U3795 (N_3795,N_2204,N_2142);
xor U3796 (N_3796,N_2898,N_2029);
nor U3797 (N_3797,N_2716,N_2271);
nor U3798 (N_3798,N_2668,N_2812);
nor U3799 (N_3799,N_2571,N_2354);
nand U3800 (N_3800,N_2190,N_2379);
nand U3801 (N_3801,N_2277,N_2170);
nor U3802 (N_3802,N_2394,N_2607);
xor U3803 (N_3803,N_2461,N_2339);
nor U3804 (N_3804,N_2199,N_2348);
or U3805 (N_3805,N_2527,N_2027);
xnor U3806 (N_3806,N_2831,N_2740);
nand U3807 (N_3807,N_2578,N_2594);
and U3808 (N_3808,N_2793,N_2317);
or U3809 (N_3809,N_2645,N_2229);
nor U3810 (N_3810,N_2776,N_2836);
and U3811 (N_3811,N_2996,N_2894);
and U3812 (N_3812,N_2604,N_2768);
nor U3813 (N_3813,N_2188,N_2904);
or U3814 (N_3814,N_2343,N_2622);
or U3815 (N_3815,N_2290,N_2033);
and U3816 (N_3816,N_2777,N_2390);
and U3817 (N_3817,N_2382,N_2707);
nand U3818 (N_3818,N_2871,N_2894);
xor U3819 (N_3819,N_2312,N_2656);
or U3820 (N_3820,N_2933,N_2294);
or U3821 (N_3821,N_2737,N_2566);
and U3822 (N_3822,N_2130,N_2163);
nand U3823 (N_3823,N_2706,N_2496);
nand U3824 (N_3824,N_2098,N_2579);
and U3825 (N_3825,N_2736,N_2051);
or U3826 (N_3826,N_2935,N_2664);
or U3827 (N_3827,N_2223,N_2340);
or U3828 (N_3828,N_2277,N_2125);
or U3829 (N_3829,N_2201,N_2316);
nand U3830 (N_3830,N_2787,N_2346);
xor U3831 (N_3831,N_2159,N_2909);
nor U3832 (N_3832,N_2258,N_2247);
or U3833 (N_3833,N_2176,N_2433);
or U3834 (N_3834,N_2388,N_2506);
nor U3835 (N_3835,N_2825,N_2076);
nand U3836 (N_3836,N_2902,N_2712);
nor U3837 (N_3837,N_2589,N_2829);
nand U3838 (N_3838,N_2409,N_2688);
nor U3839 (N_3839,N_2472,N_2488);
and U3840 (N_3840,N_2720,N_2151);
nand U3841 (N_3841,N_2481,N_2154);
nand U3842 (N_3842,N_2966,N_2552);
nand U3843 (N_3843,N_2402,N_2527);
nor U3844 (N_3844,N_2846,N_2313);
or U3845 (N_3845,N_2509,N_2895);
nor U3846 (N_3846,N_2841,N_2618);
or U3847 (N_3847,N_2910,N_2338);
or U3848 (N_3848,N_2248,N_2451);
nor U3849 (N_3849,N_2951,N_2178);
and U3850 (N_3850,N_2709,N_2166);
nor U3851 (N_3851,N_2976,N_2202);
or U3852 (N_3852,N_2294,N_2126);
nand U3853 (N_3853,N_2374,N_2183);
and U3854 (N_3854,N_2067,N_2896);
nand U3855 (N_3855,N_2979,N_2938);
xor U3856 (N_3856,N_2150,N_2966);
or U3857 (N_3857,N_2735,N_2551);
xnor U3858 (N_3858,N_2516,N_2057);
and U3859 (N_3859,N_2318,N_2051);
or U3860 (N_3860,N_2784,N_2612);
nand U3861 (N_3861,N_2169,N_2484);
nand U3862 (N_3862,N_2923,N_2575);
or U3863 (N_3863,N_2746,N_2193);
nor U3864 (N_3864,N_2418,N_2852);
xnor U3865 (N_3865,N_2109,N_2348);
or U3866 (N_3866,N_2301,N_2465);
or U3867 (N_3867,N_2158,N_2661);
nand U3868 (N_3868,N_2543,N_2688);
nor U3869 (N_3869,N_2235,N_2310);
and U3870 (N_3870,N_2808,N_2595);
or U3871 (N_3871,N_2744,N_2626);
nand U3872 (N_3872,N_2844,N_2364);
nand U3873 (N_3873,N_2585,N_2300);
nand U3874 (N_3874,N_2926,N_2770);
nand U3875 (N_3875,N_2267,N_2714);
nand U3876 (N_3876,N_2426,N_2552);
or U3877 (N_3877,N_2258,N_2121);
nand U3878 (N_3878,N_2123,N_2318);
nor U3879 (N_3879,N_2763,N_2169);
or U3880 (N_3880,N_2126,N_2230);
or U3881 (N_3881,N_2910,N_2036);
nor U3882 (N_3882,N_2551,N_2216);
or U3883 (N_3883,N_2200,N_2554);
and U3884 (N_3884,N_2679,N_2886);
or U3885 (N_3885,N_2283,N_2465);
or U3886 (N_3886,N_2831,N_2601);
and U3887 (N_3887,N_2919,N_2328);
xnor U3888 (N_3888,N_2817,N_2278);
and U3889 (N_3889,N_2306,N_2685);
and U3890 (N_3890,N_2928,N_2978);
or U3891 (N_3891,N_2100,N_2597);
and U3892 (N_3892,N_2619,N_2857);
nor U3893 (N_3893,N_2007,N_2614);
and U3894 (N_3894,N_2807,N_2773);
nand U3895 (N_3895,N_2596,N_2061);
nor U3896 (N_3896,N_2268,N_2965);
or U3897 (N_3897,N_2849,N_2236);
or U3898 (N_3898,N_2718,N_2816);
xor U3899 (N_3899,N_2740,N_2450);
and U3900 (N_3900,N_2967,N_2682);
xnor U3901 (N_3901,N_2656,N_2232);
and U3902 (N_3902,N_2789,N_2871);
xnor U3903 (N_3903,N_2468,N_2237);
and U3904 (N_3904,N_2467,N_2413);
or U3905 (N_3905,N_2951,N_2546);
xnor U3906 (N_3906,N_2576,N_2168);
or U3907 (N_3907,N_2532,N_2255);
and U3908 (N_3908,N_2651,N_2474);
nand U3909 (N_3909,N_2303,N_2851);
or U3910 (N_3910,N_2299,N_2503);
nand U3911 (N_3911,N_2049,N_2063);
or U3912 (N_3912,N_2815,N_2272);
or U3913 (N_3913,N_2769,N_2746);
or U3914 (N_3914,N_2122,N_2262);
or U3915 (N_3915,N_2814,N_2141);
nand U3916 (N_3916,N_2160,N_2955);
xnor U3917 (N_3917,N_2590,N_2694);
nand U3918 (N_3918,N_2882,N_2428);
and U3919 (N_3919,N_2497,N_2265);
or U3920 (N_3920,N_2840,N_2460);
xor U3921 (N_3921,N_2417,N_2941);
xnor U3922 (N_3922,N_2584,N_2827);
nor U3923 (N_3923,N_2152,N_2673);
xor U3924 (N_3924,N_2087,N_2337);
or U3925 (N_3925,N_2365,N_2057);
and U3926 (N_3926,N_2040,N_2161);
and U3927 (N_3927,N_2016,N_2141);
nor U3928 (N_3928,N_2834,N_2872);
nand U3929 (N_3929,N_2832,N_2883);
and U3930 (N_3930,N_2119,N_2851);
xor U3931 (N_3931,N_2613,N_2137);
and U3932 (N_3932,N_2801,N_2305);
or U3933 (N_3933,N_2779,N_2610);
nor U3934 (N_3934,N_2857,N_2135);
nor U3935 (N_3935,N_2168,N_2438);
nor U3936 (N_3936,N_2408,N_2968);
or U3937 (N_3937,N_2973,N_2214);
nand U3938 (N_3938,N_2038,N_2477);
xor U3939 (N_3939,N_2674,N_2631);
or U3940 (N_3940,N_2434,N_2377);
nand U3941 (N_3941,N_2243,N_2518);
nand U3942 (N_3942,N_2928,N_2478);
xor U3943 (N_3943,N_2653,N_2672);
and U3944 (N_3944,N_2175,N_2278);
and U3945 (N_3945,N_2742,N_2067);
nor U3946 (N_3946,N_2964,N_2372);
nand U3947 (N_3947,N_2500,N_2973);
nand U3948 (N_3948,N_2239,N_2998);
or U3949 (N_3949,N_2498,N_2101);
and U3950 (N_3950,N_2508,N_2959);
nand U3951 (N_3951,N_2617,N_2667);
nor U3952 (N_3952,N_2347,N_2169);
nor U3953 (N_3953,N_2322,N_2851);
or U3954 (N_3954,N_2464,N_2940);
nand U3955 (N_3955,N_2179,N_2365);
xor U3956 (N_3956,N_2260,N_2528);
nor U3957 (N_3957,N_2955,N_2921);
and U3958 (N_3958,N_2979,N_2032);
or U3959 (N_3959,N_2400,N_2102);
nand U3960 (N_3960,N_2595,N_2314);
or U3961 (N_3961,N_2335,N_2572);
nand U3962 (N_3962,N_2350,N_2290);
nor U3963 (N_3963,N_2630,N_2841);
nand U3964 (N_3964,N_2728,N_2131);
nand U3965 (N_3965,N_2082,N_2183);
nor U3966 (N_3966,N_2345,N_2852);
and U3967 (N_3967,N_2054,N_2159);
nor U3968 (N_3968,N_2860,N_2424);
and U3969 (N_3969,N_2974,N_2607);
nor U3970 (N_3970,N_2800,N_2303);
xnor U3971 (N_3971,N_2845,N_2346);
or U3972 (N_3972,N_2940,N_2449);
nor U3973 (N_3973,N_2068,N_2535);
and U3974 (N_3974,N_2655,N_2028);
and U3975 (N_3975,N_2576,N_2281);
or U3976 (N_3976,N_2099,N_2091);
nor U3977 (N_3977,N_2047,N_2758);
nand U3978 (N_3978,N_2721,N_2104);
and U3979 (N_3979,N_2748,N_2178);
xnor U3980 (N_3980,N_2070,N_2372);
nor U3981 (N_3981,N_2927,N_2570);
nand U3982 (N_3982,N_2627,N_2935);
nand U3983 (N_3983,N_2002,N_2847);
or U3984 (N_3984,N_2888,N_2854);
xnor U3985 (N_3985,N_2357,N_2229);
and U3986 (N_3986,N_2586,N_2489);
nand U3987 (N_3987,N_2122,N_2112);
or U3988 (N_3988,N_2931,N_2526);
xnor U3989 (N_3989,N_2159,N_2385);
or U3990 (N_3990,N_2138,N_2022);
nor U3991 (N_3991,N_2668,N_2828);
nand U3992 (N_3992,N_2861,N_2373);
nand U3993 (N_3993,N_2862,N_2456);
and U3994 (N_3994,N_2262,N_2684);
nand U3995 (N_3995,N_2311,N_2396);
xnor U3996 (N_3996,N_2440,N_2462);
xor U3997 (N_3997,N_2963,N_2844);
or U3998 (N_3998,N_2137,N_2297);
or U3999 (N_3999,N_2438,N_2018);
nor U4000 (N_4000,N_3577,N_3166);
or U4001 (N_4001,N_3034,N_3480);
or U4002 (N_4002,N_3689,N_3580);
nand U4003 (N_4003,N_3040,N_3054);
or U4004 (N_4004,N_3059,N_3615);
nand U4005 (N_4005,N_3135,N_3940);
nor U4006 (N_4006,N_3065,N_3531);
and U4007 (N_4007,N_3275,N_3724);
or U4008 (N_4008,N_3351,N_3937);
or U4009 (N_4009,N_3907,N_3290);
and U4010 (N_4010,N_3323,N_3790);
or U4011 (N_4011,N_3637,N_3174);
or U4012 (N_4012,N_3903,N_3421);
or U4013 (N_4013,N_3855,N_3253);
or U4014 (N_4014,N_3045,N_3908);
nand U4015 (N_4015,N_3526,N_3538);
nand U4016 (N_4016,N_3869,N_3079);
nand U4017 (N_4017,N_3023,N_3212);
xor U4018 (N_4018,N_3634,N_3737);
and U4019 (N_4019,N_3407,N_3303);
or U4020 (N_4020,N_3990,N_3794);
or U4021 (N_4021,N_3168,N_3931);
and U4022 (N_4022,N_3177,N_3556);
or U4023 (N_4023,N_3611,N_3337);
or U4024 (N_4024,N_3194,N_3941);
or U4025 (N_4025,N_3492,N_3600);
or U4026 (N_4026,N_3491,N_3242);
and U4027 (N_4027,N_3442,N_3682);
and U4028 (N_4028,N_3785,N_3630);
nor U4029 (N_4029,N_3211,N_3613);
or U4030 (N_4030,N_3922,N_3128);
nor U4031 (N_4031,N_3277,N_3341);
or U4032 (N_4032,N_3245,N_3692);
and U4033 (N_4033,N_3821,N_3278);
nor U4034 (N_4034,N_3752,N_3878);
and U4035 (N_4035,N_3427,N_3814);
nand U4036 (N_4036,N_3149,N_3033);
xor U4037 (N_4037,N_3701,N_3688);
nand U4038 (N_4038,N_3781,N_3244);
xnor U4039 (N_4039,N_3017,N_3058);
or U4040 (N_4040,N_3266,N_3532);
and U4041 (N_4041,N_3552,N_3331);
and U4042 (N_4042,N_3932,N_3384);
and U4043 (N_4043,N_3909,N_3228);
or U4044 (N_4044,N_3731,N_3178);
or U4045 (N_4045,N_3569,N_3632);
nor U4046 (N_4046,N_3036,N_3896);
nand U4047 (N_4047,N_3025,N_3226);
nand U4048 (N_4048,N_3606,N_3155);
nand U4049 (N_4049,N_3392,N_3010);
and U4050 (N_4050,N_3276,N_3404);
nand U4051 (N_4051,N_3772,N_3215);
or U4052 (N_4052,N_3111,N_3496);
nor U4053 (N_4053,N_3679,N_3798);
and U4054 (N_4054,N_3476,N_3339);
nor U4055 (N_4055,N_3957,N_3830);
nand U4056 (N_4056,N_3271,N_3874);
or U4057 (N_4057,N_3140,N_3816);
nand U4058 (N_4058,N_3070,N_3340);
and U4059 (N_4059,N_3102,N_3915);
or U4060 (N_4060,N_3515,N_3343);
nor U4061 (N_4061,N_3997,N_3097);
or U4062 (N_4062,N_3839,N_3346);
nand U4063 (N_4063,N_3396,N_3857);
and U4064 (N_4064,N_3428,N_3049);
or U4065 (N_4065,N_3224,N_3365);
nor U4066 (N_4066,N_3248,N_3527);
and U4067 (N_4067,N_3848,N_3119);
xor U4068 (N_4068,N_3802,N_3176);
xor U4069 (N_4069,N_3638,N_3449);
or U4070 (N_4070,N_3456,N_3192);
nor U4071 (N_4071,N_3674,N_3465);
nor U4072 (N_4072,N_3451,N_3550);
nor U4073 (N_4073,N_3963,N_3944);
or U4074 (N_4074,N_3482,N_3769);
nand U4075 (N_4075,N_3188,N_3046);
or U4076 (N_4076,N_3359,N_3640);
nor U4077 (N_4077,N_3804,N_3795);
nand U4078 (N_4078,N_3060,N_3305);
and U4079 (N_4079,N_3240,N_3317);
and U4080 (N_4080,N_3865,N_3230);
or U4081 (N_4081,N_3601,N_3705);
nor U4082 (N_4082,N_3051,N_3858);
nand U4083 (N_4083,N_3513,N_3318);
xnor U4084 (N_4084,N_3229,N_3838);
or U4085 (N_4085,N_3555,N_3412);
nand U4086 (N_4086,N_3923,N_3622);
nand U4087 (N_4087,N_3257,N_3645);
nor U4088 (N_4088,N_3464,N_3787);
xor U4089 (N_4089,N_3319,N_3121);
and U4090 (N_4090,N_3489,N_3703);
nand U4091 (N_4091,N_3844,N_3993);
nor U4092 (N_4092,N_3545,N_3395);
nor U4093 (N_4093,N_3072,N_3131);
or U4094 (N_4094,N_3648,N_3180);
or U4095 (N_4095,N_3543,N_3946);
nor U4096 (N_4096,N_3831,N_3383);
or U4097 (N_4097,N_3547,N_3684);
xor U4098 (N_4098,N_3366,N_3508);
xor U4099 (N_4099,N_3676,N_3849);
nor U4100 (N_4100,N_3891,N_3759);
nor U4101 (N_4101,N_3742,N_3503);
xor U4102 (N_4102,N_3467,N_3165);
nand U4103 (N_4103,N_3726,N_3882);
and U4104 (N_4104,N_3163,N_3235);
and U4105 (N_4105,N_3595,N_3541);
or U4106 (N_4106,N_3069,N_3900);
or U4107 (N_4107,N_3660,N_3586);
or U4108 (N_4108,N_3976,N_3933);
nor U4109 (N_4109,N_3884,N_3610);
nor U4110 (N_4110,N_3446,N_3353);
nor U4111 (N_4111,N_3144,N_3517);
and U4112 (N_4112,N_3514,N_3700);
nor U4113 (N_4113,N_3588,N_3087);
or U4114 (N_4114,N_3336,N_3342);
xor U4115 (N_4115,N_3707,N_3860);
nor U4116 (N_4116,N_3950,N_3528);
or U4117 (N_4117,N_3916,N_3347);
or U4118 (N_4118,N_3362,N_3280);
xnor U4119 (N_4119,N_3284,N_3520);
xor U4120 (N_4120,N_3090,N_3551);
nor U4121 (N_4121,N_3071,N_3789);
nor U4122 (N_4122,N_3161,N_3107);
and U4123 (N_4123,N_3487,N_3559);
and U4124 (N_4124,N_3995,N_3263);
xnor U4125 (N_4125,N_3238,N_3420);
or U4126 (N_4126,N_3740,N_3589);
nand U4127 (N_4127,N_3231,N_3208);
nor U4128 (N_4128,N_3669,N_3098);
nor U4129 (N_4129,N_3246,N_3668);
nor U4130 (N_4130,N_3425,N_3289);
nand U4131 (N_4131,N_3698,N_3502);
xnor U4132 (N_4132,N_3554,N_3394);
and U4133 (N_4133,N_3416,N_3022);
or U4134 (N_4134,N_3762,N_3778);
nor U4135 (N_4135,N_3112,N_3979);
nor U4136 (N_4136,N_3130,N_3743);
nor U4137 (N_4137,N_3965,N_3234);
or U4138 (N_4138,N_3094,N_3003);
nor U4139 (N_4139,N_3695,N_3454);
xnor U4140 (N_4140,N_3475,N_3880);
and U4141 (N_4141,N_3445,N_3607);
and U4142 (N_4142,N_3481,N_3747);
nand U4143 (N_4143,N_3160,N_3977);
or U4144 (N_4144,N_3633,N_3067);
and U4145 (N_4145,N_3897,N_3564);
xor U4146 (N_4146,N_3443,N_3162);
nand U4147 (N_4147,N_3126,N_3297);
or U4148 (N_4148,N_3616,N_3409);
nor U4149 (N_4149,N_3103,N_3581);
and U4150 (N_4150,N_3530,N_3222);
and U4151 (N_4151,N_3856,N_3936);
and U4152 (N_4152,N_3593,N_3056);
or U4153 (N_4153,N_3175,N_3328);
nor U4154 (N_4154,N_3643,N_3618);
nor U4155 (N_4155,N_3375,N_3851);
nand U4156 (N_4156,N_3507,N_3115);
and U4157 (N_4157,N_3823,N_3237);
nor U4158 (N_4158,N_3068,N_3084);
nand U4159 (N_4159,N_3009,N_3898);
nand U4160 (N_4160,N_3085,N_3959);
and U4161 (N_4161,N_3599,N_3501);
and U4162 (N_4162,N_3980,N_3935);
and U4163 (N_4163,N_3354,N_3619);
nand U4164 (N_4164,N_3125,N_3751);
nand U4165 (N_4165,N_3225,N_3078);
or U4166 (N_4166,N_3544,N_3516);
and U4167 (N_4167,N_3870,N_3764);
and U4168 (N_4168,N_3939,N_3183);
nand U4169 (N_4169,N_3938,N_3157);
nand U4170 (N_4170,N_3716,N_3984);
and U4171 (N_4171,N_3199,N_3788);
or U4172 (N_4172,N_3461,N_3195);
nor U4173 (N_4173,N_3560,N_3817);
nand U4174 (N_4174,N_3720,N_3139);
or U4175 (N_4175,N_3437,N_3267);
or U4176 (N_4176,N_3846,N_3397);
nor U4177 (N_4177,N_3757,N_3118);
nand U4178 (N_4178,N_3986,N_3966);
and U4179 (N_4179,N_3904,N_3888);
xnor U4180 (N_4180,N_3770,N_3082);
and U4181 (N_4181,N_3924,N_3345);
xor U4182 (N_4182,N_3748,N_3500);
nor U4183 (N_4183,N_3575,N_3053);
and U4184 (N_4184,N_3686,N_3974);
or U4185 (N_4185,N_3291,N_3447);
and U4186 (N_4186,N_3361,N_3138);
and U4187 (N_4187,N_3326,N_3929);
or U4188 (N_4188,N_3256,N_3463);
or U4189 (N_4189,N_3307,N_3232);
or U4190 (N_4190,N_3988,N_3408);
or U4191 (N_4191,N_3598,N_3441);
nand U4192 (N_4192,N_3697,N_3110);
xor U4193 (N_4193,N_3871,N_3647);
or U4194 (N_4194,N_3962,N_3076);
and U4195 (N_4195,N_3887,N_3808);
and U4196 (N_4196,N_3631,N_3358);
nor U4197 (N_4197,N_3523,N_3928);
or U4198 (N_4198,N_3709,N_3310);
and U4199 (N_4199,N_3730,N_3654);
and U4200 (N_4200,N_3573,N_3609);
or U4201 (N_4201,N_3723,N_3591);
nor U4202 (N_4202,N_3822,N_3173);
and U4203 (N_4203,N_3088,N_3548);
nor U4204 (N_4204,N_3875,N_3587);
and U4205 (N_4205,N_3357,N_3594);
or U4206 (N_4206,N_3419,N_3145);
nor U4207 (N_4207,N_3189,N_3702);
nand U4208 (N_4208,N_3745,N_3952);
and U4209 (N_4209,N_3038,N_3032);
nor U4210 (N_4210,N_3095,N_3827);
and U4211 (N_4211,N_3854,N_3836);
or U4212 (N_4212,N_3430,N_3910);
and U4213 (N_4213,N_3294,N_3063);
nor U4214 (N_4214,N_3868,N_3512);
or U4215 (N_4215,N_3471,N_3967);
and U4216 (N_4216,N_3998,N_3279);
nor U4217 (N_4217,N_3114,N_3380);
or U4218 (N_4218,N_3249,N_3227);
and U4219 (N_4219,N_3184,N_3704);
or U4220 (N_4220,N_3272,N_3185);
nor U4221 (N_4221,N_3953,N_3756);
nand U4222 (N_4222,N_3106,N_3382);
and U4223 (N_4223,N_3217,N_3494);
xnor U4224 (N_4224,N_3829,N_3044);
and U4225 (N_4225,N_3920,N_3735);
xor U4226 (N_4226,N_3363,N_3288);
or U4227 (N_4227,N_3876,N_3295);
and U4228 (N_4228,N_3432,N_3561);
or U4229 (N_4229,N_3608,N_3566);
or U4230 (N_4230,N_3540,N_3028);
and U4231 (N_4231,N_3300,N_3687);
nor U4232 (N_4232,N_3158,N_3287);
nor U4233 (N_4233,N_3434,N_3123);
and U4234 (N_4234,N_3859,N_3843);
and U4235 (N_4235,N_3867,N_3578);
xnor U4236 (N_4236,N_3945,N_3086);
nor U4237 (N_4237,N_3925,N_3251);
and U4238 (N_4238,N_3711,N_3522);
and U4239 (N_4239,N_3186,N_3265);
nor U4240 (N_4240,N_3727,N_3777);
nand U4241 (N_4241,N_3919,N_3298);
or U4242 (N_4242,N_3623,N_3218);
xnor U4243 (N_4243,N_3377,N_3152);
or U4244 (N_4244,N_3570,N_3582);
xor U4245 (N_4245,N_3406,N_3536);
nand U4246 (N_4246,N_3971,N_3338);
or U4247 (N_4247,N_3485,N_3768);
xor U4248 (N_4248,N_3498,N_3886);
nor U4249 (N_4249,N_3433,N_3429);
nor U4250 (N_4250,N_3733,N_3292);
or U4251 (N_4251,N_3493,N_3504);
or U4252 (N_4252,N_3863,N_3081);
and U4253 (N_4253,N_3565,N_3926);
or U4254 (N_4254,N_3220,N_3850);
nor U4255 (N_4255,N_3665,N_3982);
and U4256 (N_4256,N_3533,N_3005);
nand U4257 (N_4257,N_3490,N_3042);
and U4258 (N_4258,N_3243,N_3393);
or U4259 (N_4259,N_3385,N_3579);
and U4260 (N_4260,N_3656,N_3386);
or U4261 (N_4261,N_3191,N_3422);
nor U4262 (N_4262,N_3614,N_3975);
and U4263 (N_4263,N_3690,N_3864);
nor U4264 (N_4264,N_3260,N_3439);
nand U4265 (N_4265,N_3813,N_3329);
nand U4266 (N_4266,N_3311,N_3728);
nand U4267 (N_4267,N_3077,N_3400);
nor U4268 (N_4268,N_3373,N_3722);
and U4269 (N_4269,N_3378,N_3983);
xnor U4270 (N_4270,N_3806,N_3732);
and U4271 (N_4271,N_3511,N_3283);
xor U4272 (N_4272,N_3809,N_3129);
nand U4273 (N_4273,N_3478,N_3807);
and U4274 (N_4274,N_3779,N_3472);
nor U4275 (N_4275,N_3364,N_3193);
xnor U4276 (N_4276,N_3096,N_3281);
nor U4277 (N_4277,N_3468,N_3774);
and U4278 (N_4278,N_3027,N_3572);
nor U4279 (N_4279,N_3196,N_3101);
or U4280 (N_4280,N_3398,N_3801);
nand U4281 (N_4281,N_3602,N_3255);
nand U4282 (N_4282,N_3661,N_3996);
xnor U4283 (N_4283,N_3466,N_3655);
nor U4284 (N_4284,N_3948,N_3391);
nand U4285 (N_4285,N_3021,N_3273);
nor U4286 (N_4286,N_3842,N_3198);
nor U4287 (N_4287,N_3209,N_3847);
and U4288 (N_4288,N_3505,N_3902);
nand U4289 (N_4289,N_3987,N_3073);
or U4290 (N_4290,N_3368,N_3693);
or U4291 (N_4291,N_3803,N_3985);
nor U4292 (N_4292,N_3156,N_3074);
and U4293 (N_4293,N_3004,N_3308);
and U4294 (N_4294,N_3518,N_3141);
or U4295 (N_4295,N_3321,N_3435);
xnor U4296 (N_4296,N_3201,N_3438);
xor U4297 (N_4297,N_3956,N_3685);
nor U4298 (N_4298,N_3765,N_3969);
nor U4299 (N_4299,N_3426,N_3080);
nand U4300 (N_4300,N_3546,N_3892);
or U4301 (N_4301,N_3968,N_3122);
nor U4302 (N_4302,N_3455,N_3893);
or U4303 (N_4303,N_3549,N_3497);
or U4304 (N_4304,N_3453,N_3000);
xnor U4305 (N_4305,N_3644,N_3773);
nor U4306 (N_4306,N_3026,N_3458);
or U4307 (N_4307,N_3889,N_3642);
and U4308 (N_4308,N_3370,N_3066);
nand U4309 (N_4309,N_3011,N_3791);
xnor U4310 (N_4310,N_3890,N_3629);
or U4311 (N_4311,N_3050,N_3845);
and U4312 (N_4312,N_3143,N_3994);
and U4313 (N_4313,N_3031,N_3167);
nand U4314 (N_4314,N_3861,N_3372);
or U4315 (N_4315,N_3360,N_3499);
nand U4316 (N_4316,N_3350,N_3583);
nor U4317 (N_4317,N_3320,N_3403);
nand U4318 (N_4318,N_3895,N_3763);
nand U4319 (N_4319,N_3571,N_3169);
xnor U4320 (N_4320,N_3239,N_3954);
or U4321 (N_4321,N_3658,N_3413);
or U4322 (N_4322,N_3495,N_3596);
nand U4323 (N_4323,N_3349,N_3335);
nand U4324 (N_4324,N_3374,N_3746);
and U4325 (N_4325,N_3824,N_3092);
nor U4326 (N_4326,N_3127,N_3091);
nand U4327 (N_4327,N_3563,N_3673);
nand U4328 (N_4328,N_3799,N_3402);
and U4329 (N_4329,N_3782,N_3057);
and U4330 (N_4330,N_3930,N_3672);
and U4331 (N_4331,N_3474,N_3261);
or U4332 (N_4332,N_3109,N_3214);
nor U4333 (N_4333,N_3815,N_3285);
xor U4334 (N_4334,N_3411,N_3992);
xor U4335 (N_4335,N_3605,N_3268);
nor U4336 (N_4336,N_3269,N_3677);
nand U4337 (N_4337,N_3911,N_3043);
xor U4338 (N_4338,N_3436,N_3834);
and U4339 (N_4339,N_3410,N_3755);
or U4340 (N_4340,N_3424,N_3734);
nand U4341 (N_4341,N_3905,N_3213);
nand U4342 (N_4342,N_3016,N_3714);
nand U4343 (N_4343,N_3306,N_3171);
and U4344 (N_4344,N_3008,N_3901);
xnor U4345 (N_4345,N_3484,N_3356);
or U4346 (N_4346,N_3825,N_3534);
and U4347 (N_4347,N_3918,N_3749);
nand U4348 (N_4348,N_3262,N_3664);
nand U4349 (N_4349,N_3883,N_3894);
nand U4350 (N_4350,N_3694,N_3620);
and U4351 (N_4351,N_3835,N_3172);
or U4352 (N_4352,N_3147,N_3286);
nor U4353 (N_4353,N_3483,N_3628);
xor U4354 (N_4354,N_3585,N_3713);
nand U4355 (N_4355,N_3444,N_3783);
nand U4356 (N_4356,N_3666,N_3473);
nor U4357 (N_4357,N_3187,N_3797);
and U4358 (N_4358,N_3812,N_3678);
nand U4359 (N_4359,N_3719,N_3236);
and U4360 (N_4360,N_3099,N_3680);
and U4361 (N_4361,N_3542,N_3019);
and U4362 (N_4362,N_3061,N_3604);
or U4363 (N_4363,N_3052,N_3250);
nor U4364 (N_4364,N_3899,N_3576);
nor U4365 (N_4365,N_3667,N_3978);
or U4366 (N_4366,N_3047,N_3137);
nand U4367 (N_4367,N_3592,N_3352);
or U4368 (N_4368,N_3348,N_3776);
and U4369 (N_4369,N_3837,N_3786);
and U4370 (N_4370,N_3379,N_3367);
xor U4371 (N_4371,N_3780,N_3659);
and U4372 (N_4372,N_3683,N_3767);
or U4373 (N_4373,N_3691,N_3866);
and U4374 (N_4374,N_3729,N_3216);
nand U4375 (N_4375,N_3626,N_3029);
nor U4376 (N_4376,N_3334,N_3089);
and U4377 (N_4377,N_3116,N_3270);
and U4378 (N_4378,N_3826,N_3293);
and U4379 (N_4379,N_3037,N_3970);
and U4380 (N_4380,N_3706,N_3146);
xor U4381 (N_4381,N_3862,N_3991);
and U4382 (N_4382,N_3206,N_3521);
xnor U4383 (N_4383,N_3927,N_3274);
and U4384 (N_4384,N_3327,N_3190);
and U4385 (N_4385,N_3917,N_3590);
nand U4386 (N_4386,N_3639,N_3775);
or U4387 (N_4387,N_3553,N_3636);
nand U4388 (N_4388,N_3316,N_3197);
nand U4389 (N_4389,N_3325,N_3738);
and U4390 (N_4390,N_3388,N_3369);
or U4391 (N_4391,N_3584,N_3819);
nor U4392 (N_4392,N_3947,N_3148);
nor U4393 (N_4393,N_3041,N_3431);
xor U4394 (N_4394,N_3840,N_3558);
or U4395 (N_4395,N_3333,N_3539);
and U4396 (N_4396,N_3663,N_3381);
or U4397 (N_4397,N_3299,N_3535);
or U4398 (N_4398,N_3376,N_3170);
nor U4399 (N_4399,N_3964,N_3247);
nor U4400 (N_4400,N_3204,N_3007);
and U4401 (N_4401,N_3418,N_3750);
nor U4402 (N_4402,N_3440,N_3989);
nand U4403 (N_4403,N_3972,N_3179);
or U4404 (N_4404,N_3717,N_3828);
or U4405 (N_4405,N_3912,N_3399);
or U4406 (N_4406,N_3653,N_3133);
nor U4407 (N_4407,N_3083,N_3259);
nand U4408 (N_4408,N_3486,N_3557);
xor U4409 (N_4409,N_3784,N_3617);
and U4410 (N_4410,N_3387,N_3833);
nor U4411 (N_4411,N_3800,N_3671);
or U4412 (N_4412,N_3509,N_3696);
nor U4413 (N_4413,N_3048,N_3312);
xnor U4414 (N_4414,N_3766,N_3736);
nor U4415 (N_4415,N_3233,N_3405);
and U4416 (N_4416,N_3142,N_3675);
nor U4417 (N_4417,N_3150,N_3258);
xor U4418 (N_4418,N_3314,N_3039);
nor U4419 (N_4419,N_3020,N_3914);
or U4420 (N_4420,N_3670,N_3104);
nor U4421 (N_4421,N_3223,N_3567);
and U4422 (N_4422,N_3030,N_3221);
nor U4423 (N_4423,N_3818,N_3574);
or U4424 (N_4424,N_3524,N_3650);
nor U4425 (N_4425,N_3018,N_3792);
or U4426 (N_4426,N_3568,N_3417);
nand U4427 (N_4427,N_3753,N_3960);
nand U4428 (N_4428,N_3649,N_3452);
nand U4429 (N_4429,N_3124,N_3062);
xnor U4430 (N_4430,N_3662,N_3949);
nand U4431 (N_4431,N_3760,N_3793);
and U4432 (N_4432,N_3641,N_3510);
nand U4433 (N_4433,N_3771,N_3635);
or U4434 (N_4434,N_3652,N_3315);
nand U4435 (N_4435,N_3120,N_3055);
nand U4436 (N_4436,N_3537,N_3881);
xor U4437 (N_4437,N_3758,N_3304);
or U4438 (N_4438,N_3093,N_3014);
nor U4439 (N_4439,N_3462,N_3296);
and U4440 (N_4440,N_3885,N_3390);
nor U4441 (N_4441,N_3942,N_3739);
or U4442 (N_4442,N_3252,N_3282);
and U4443 (N_4443,N_3159,N_3906);
and U4444 (N_4444,N_3820,N_3708);
xnor U4445 (N_4445,N_3401,N_3488);
nor U4446 (N_4446,N_3627,N_3264);
nand U4447 (N_4447,N_3035,N_3612);
xor U4448 (N_4448,N_3132,N_3961);
and U4449 (N_4449,N_3075,N_3853);
xor U4450 (N_4450,N_3371,N_3457);
or U4451 (N_4451,N_3718,N_3415);
or U4452 (N_4452,N_3302,N_3448);
xnor U4453 (N_4453,N_3301,N_3205);
or U4454 (N_4454,N_3741,N_3460);
and U4455 (N_4455,N_3951,N_3872);
nor U4456 (N_4456,N_3744,N_3254);
or U4457 (N_4457,N_3108,N_3519);
xor U4458 (N_4458,N_3624,N_3879);
or U4459 (N_4459,N_3006,N_3913);
nor U4460 (N_4460,N_3151,N_3113);
nand U4461 (N_4461,N_3529,N_3210);
or U4462 (N_4462,N_3241,N_3117);
nor U4463 (N_4463,N_3506,N_3015);
nand U4464 (N_4464,N_3958,N_3651);
nor U4465 (N_4465,N_3715,N_3562);
nor U4466 (N_4466,N_3810,N_3330);
and U4467 (N_4467,N_3725,N_3761);
and U4468 (N_4468,N_3154,N_3332);
or U4469 (N_4469,N_3710,N_3999);
or U4470 (N_4470,N_3182,N_3841);
and U4471 (N_4471,N_3164,N_3681);
and U4472 (N_4472,N_3934,N_3621);
nand U4473 (N_4473,N_3832,N_3805);
nand U4474 (N_4474,N_3423,N_3852);
nor U4475 (N_4475,N_3479,N_3309);
nor U4476 (N_4476,N_3754,N_3219);
nor U4477 (N_4477,N_3796,N_3625);
nor U4478 (N_4478,N_3389,N_3603);
xor U4479 (N_4479,N_3646,N_3811);
nand U4480 (N_4480,N_3100,N_3450);
nor U4481 (N_4481,N_3414,N_3877);
nand U4482 (N_4482,N_3200,N_3921);
and U4483 (N_4483,N_3344,N_3469);
nor U4484 (N_4484,N_3134,N_3699);
and U4485 (N_4485,N_3313,N_3981);
or U4486 (N_4486,N_3024,N_3136);
xor U4487 (N_4487,N_3597,N_3470);
and U4488 (N_4488,N_3001,N_3712);
xor U4489 (N_4489,N_3657,N_3955);
or U4490 (N_4490,N_3105,N_3207);
xnor U4491 (N_4491,N_3202,N_3064);
nand U4492 (N_4492,N_3203,N_3012);
nand U4493 (N_4493,N_3013,N_3322);
nand U4494 (N_4494,N_3943,N_3525);
nor U4495 (N_4495,N_3721,N_3477);
or U4496 (N_4496,N_3002,N_3459);
and U4497 (N_4497,N_3355,N_3153);
or U4498 (N_4498,N_3181,N_3324);
nand U4499 (N_4499,N_3873,N_3973);
nor U4500 (N_4500,N_3531,N_3844);
nand U4501 (N_4501,N_3657,N_3514);
nand U4502 (N_4502,N_3040,N_3084);
nand U4503 (N_4503,N_3687,N_3530);
or U4504 (N_4504,N_3193,N_3371);
nand U4505 (N_4505,N_3079,N_3872);
nand U4506 (N_4506,N_3071,N_3521);
and U4507 (N_4507,N_3595,N_3563);
and U4508 (N_4508,N_3331,N_3834);
nor U4509 (N_4509,N_3753,N_3081);
nand U4510 (N_4510,N_3814,N_3478);
or U4511 (N_4511,N_3757,N_3774);
xor U4512 (N_4512,N_3582,N_3362);
nor U4513 (N_4513,N_3648,N_3225);
nor U4514 (N_4514,N_3078,N_3489);
and U4515 (N_4515,N_3979,N_3996);
nand U4516 (N_4516,N_3083,N_3227);
and U4517 (N_4517,N_3931,N_3994);
nand U4518 (N_4518,N_3785,N_3965);
and U4519 (N_4519,N_3732,N_3019);
and U4520 (N_4520,N_3327,N_3331);
nor U4521 (N_4521,N_3930,N_3628);
or U4522 (N_4522,N_3845,N_3855);
xnor U4523 (N_4523,N_3652,N_3818);
nor U4524 (N_4524,N_3767,N_3778);
and U4525 (N_4525,N_3937,N_3809);
nor U4526 (N_4526,N_3492,N_3626);
and U4527 (N_4527,N_3559,N_3963);
nand U4528 (N_4528,N_3455,N_3218);
and U4529 (N_4529,N_3358,N_3896);
nand U4530 (N_4530,N_3536,N_3421);
xnor U4531 (N_4531,N_3731,N_3575);
and U4532 (N_4532,N_3192,N_3495);
and U4533 (N_4533,N_3370,N_3089);
and U4534 (N_4534,N_3640,N_3688);
or U4535 (N_4535,N_3675,N_3615);
nor U4536 (N_4536,N_3846,N_3350);
nand U4537 (N_4537,N_3470,N_3187);
xnor U4538 (N_4538,N_3254,N_3990);
xnor U4539 (N_4539,N_3447,N_3220);
xor U4540 (N_4540,N_3461,N_3528);
or U4541 (N_4541,N_3926,N_3101);
or U4542 (N_4542,N_3836,N_3049);
and U4543 (N_4543,N_3184,N_3124);
nor U4544 (N_4544,N_3032,N_3174);
nor U4545 (N_4545,N_3191,N_3017);
or U4546 (N_4546,N_3596,N_3124);
nand U4547 (N_4547,N_3239,N_3149);
or U4548 (N_4548,N_3399,N_3158);
nor U4549 (N_4549,N_3101,N_3546);
or U4550 (N_4550,N_3234,N_3635);
and U4551 (N_4551,N_3536,N_3128);
or U4552 (N_4552,N_3980,N_3815);
and U4553 (N_4553,N_3905,N_3243);
and U4554 (N_4554,N_3584,N_3192);
xor U4555 (N_4555,N_3666,N_3367);
nor U4556 (N_4556,N_3575,N_3892);
nand U4557 (N_4557,N_3141,N_3247);
nor U4558 (N_4558,N_3063,N_3084);
nand U4559 (N_4559,N_3539,N_3819);
nand U4560 (N_4560,N_3377,N_3208);
or U4561 (N_4561,N_3759,N_3650);
nor U4562 (N_4562,N_3931,N_3399);
nor U4563 (N_4563,N_3517,N_3606);
and U4564 (N_4564,N_3225,N_3005);
nand U4565 (N_4565,N_3339,N_3882);
or U4566 (N_4566,N_3508,N_3518);
and U4567 (N_4567,N_3562,N_3658);
nor U4568 (N_4568,N_3717,N_3076);
and U4569 (N_4569,N_3087,N_3407);
nor U4570 (N_4570,N_3917,N_3083);
and U4571 (N_4571,N_3619,N_3597);
xnor U4572 (N_4572,N_3859,N_3082);
xor U4573 (N_4573,N_3938,N_3128);
nor U4574 (N_4574,N_3835,N_3722);
and U4575 (N_4575,N_3295,N_3719);
nand U4576 (N_4576,N_3074,N_3355);
xnor U4577 (N_4577,N_3150,N_3140);
and U4578 (N_4578,N_3454,N_3087);
or U4579 (N_4579,N_3993,N_3242);
xor U4580 (N_4580,N_3969,N_3389);
and U4581 (N_4581,N_3067,N_3640);
nand U4582 (N_4582,N_3889,N_3483);
nor U4583 (N_4583,N_3315,N_3906);
and U4584 (N_4584,N_3969,N_3223);
and U4585 (N_4585,N_3561,N_3248);
nor U4586 (N_4586,N_3445,N_3861);
xnor U4587 (N_4587,N_3215,N_3175);
nand U4588 (N_4588,N_3354,N_3216);
nand U4589 (N_4589,N_3327,N_3412);
or U4590 (N_4590,N_3858,N_3238);
or U4591 (N_4591,N_3301,N_3355);
or U4592 (N_4592,N_3985,N_3116);
and U4593 (N_4593,N_3222,N_3454);
and U4594 (N_4594,N_3724,N_3650);
nand U4595 (N_4595,N_3133,N_3954);
nand U4596 (N_4596,N_3170,N_3144);
or U4597 (N_4597,N_3306,N_3610);
nand U4598 (N_4598,N_3639,N_3168);
and U4599 (N_4599,N_3912,N_3495);
xnor U4600 (N_4600,N_3068,N_3983);
xnor U4601 (N_4601,N_3738,N_3771);
nor U4602 (N_4602,N_3164,N_3462);
or U4603 (N_4603,N_3447,N_3031);
nand U4604 (N_4604,N_3743,N_3793);
xor U4605 (N_4605,N_3987,N_3262);
nand U4606 (N_4606,N_3111,N_3480);
xnor U4607 (N_4607,N_3250,N_3499);
xor U4608 (N_4608,N_3947,N_3882);
nand U4609 (N_4609,N_3988,N_3766);
nand U4610 (N_4610,N_3184,N_3346);
xnor U4611 (N_4611,N_3121,N_3268);
or U4612 (N_4612,N_3956,N_3013);
nor U4613 (N_4613,N_3296,N_3188);
nand U4614 (N_4614,N_3374,N_3267);
or U4615 (N_4615,N_3200,N_3132);
nor U4616 (N_4616,N_3213,N_3518);
nor U4617 (N_4617,N_3727,N_3261);
and U4618 (N_4618,N_3829,N_3327);
xnor U4619 (N_4619,N_3042,N_3323);
or U4620 (N_4620,N_3333,N_3683);
or U4621 (N_4621,N_3231,N_3168);
nand U4622 (N_4622,N_3137,N_3744);
or U4623 (N_4623,N_3578,N_3893);
or U4624 (N_4624,N_3738,N_3510);
nand U4625 (N_4625,N_3531,N_3201);
nand U4626 (N_4626,N_3803,N_3936);
and U4627 (N_4627,N_3537,N_3954);
nor U4628 (N_4628,N_3441,N_3663);
and U4629 (N_4629,N_3587,N_3770);
or U4630 (N_4630,N_3936,N_3421);
nor U4631 (N_4631,N_3120,N_3324);
or U4632 (N_4632,N_3114,N_3203);
or U4633 (N_4633,N_3053,N_3637);
and U4634 (N_4634,N_3492,N_3900);
and U4635 (N_4635,N_3330,N_3340);
nor U4636 (N_4636,N_3176,N_3888);
nand U4637 (N_4637,N_3475,N_3102);
and U4638 (N_4638,N_3466,N_3664);
nor U4639 (N_4639,N_3886,N_3246);
nand U4640 (N_4640,N_3316,N_3234);
or U4641 (N_4641,N_3534,N_3393);
xor U4642 (N_4642,N_3437,N_3009);
and U4643 (N_4643,N_3880,N_3012);
xor U4644 (N_4644,N_3717,N_3688);
nand U4645 (N_4645,N_3661,N_3352);
or U4646 (N_4646,N_3122,N_3691);
nor U4647 (N_4647,N_3021,N_3622);
nor U4648 (N_4648,N_3945,N_3650);
or U4649 (N_4649,N_3956,N_3682);
nand U4650 (N_4650,N_3483,N_3854);
or U4651 (N_4651,N_3545,N_3143);
and U4652 (N_4652,N_3233,N_3513);
nor U4653 (N_4653,N_3733,N_3146);
nand U4654 (N_4654,N_3350,N_3054);
and U4655 (N_4655,N_3520,N_3526);
nand U4656 (N_4656,N_3979,N_3666);
xnor U4657 (N_4657,N_3355,N_3002);
and U4658 (N_4658,N_3471,N_3741);
nand U4659 (N_4659,N_3521,N_3139);
or U4660 (N_4660,N_3808,N_3286);
and U4661 (N_4661,N_3156,N_3991);
nor U4662 (N_4662,N_3057,N_3690);
nand U4663 (N_4663,N_3374,N_3318);
and U4664 (N_4664,N_3864,N_3252);
and U4665 (N_4665,N_3940,N_3657);
nand U4666 (N_4666,N_3212,N_3933);
or U4667 (N_4667,N_3324,N_3309);
xor U4668 (N_4668,N_3579,N_3092);
or U4669 (N_4669,N_3442,N_3704);
nand U4670 (N_4670,N_3948,N_3240);
or U4671 (N_4671,N_3536,N_3650);
nand U4672 (N_4672,N_3029,N_3874);
and U4673 (N_4673,N_3006,N_3905);
or U4674 (N_4674,N_3651,N_3664);
and U4675 (N_4675,N_3414,N_3171);
nand U4676 (N_4676,N_3182,N_3818);
nand U4677 (N_4677,N_3721,N_3470);
xor U4678 (N_4678,N_3500,N_3948);
nand U4679 (N_4679,N_3448,N_3241);
and U4680 (N_4680,N_3693,N_3395);
or U4681 (N_4681,N_3767,N_3013);
and U4682 (N_4682,N_3204,N_3991);
nor U4683 (N_4683,N_3078,N_3748);
and U4684 (N_4684,N_3123,N_3689);
nor U4685 (N_4685,N_3469,N_3769);
nand U4686 (N_4686,N_3841,N_3053);
xor U4687 (N_4687,N_3259,N_3117);
xnor U4688 (N_4688,N_3730,N_3618);
nand U4689 (N_4689,N_3583,N_3216);
or U4690 (N_4690,N_3837,N_3683);
nand U4691 (N_4691,N_3641,N_3874);
nor U4692 (N_4692,N_3974,N_3021);
nor U4693 (N_4693,N_3585,N_3913);
xnor U4694 (N_4694,N_3901,N_3066);
and U4695 (N_4695,N_3480,N_3729);
and U4696 (N_4696,N_3776,N_3460);
and U4697 (N_4697,N_3607,N_3466);
nor U4698 (N_4698,N_3176,N_3335);
xor U4699 (N_4699,N_3699,N_3147);
and U4700 (N_4700,N_3377,N_3111);
or U4701 (N_4701,N_3421,N_3579);
nor U4702 (N_4702,N_3106,N_3949);
nor U4703 (N_4703,N_3847,N_3600);
xnor U4704 (N_4704,N_3266,N_3292);
and U4705 (N_4705,N_3983,N_3809);
nor U4706 (N_4706,N_3363,N_3266);
xnor U4707 (N_4707,N_3384,N_3948);
xor U4708 (N_4708,N_3846,N_3095);
nand U4709 (N_4709,N_3278,N_3760);
nor U4710 (N_4710,N_3193,N_3286);
or U4711 (N_4711,N_3494,N_3187);
or U4712 (N_4712,N_3603,N_3893);
or U4713 (N_4713,N_3576,N_3793);
nand U4714 (N_4714,N_3636,N_3113);
and U4715 (N_4715,N_3983,N_3654);
xnor U4716 (N_4716,N_3882,N_3663);
or U4717 (N_4717,N_3472,N_3369);
nor U4718 (N_4718,N_3332,N_3276);
xnor U4719 (N_4719,N_3044,N_3384);
nand U4720 (N_4720,N_3670,N_3291);
and U4721 (N_4721,N_3232,N_3580);
or U4722 (N_4722,N_3603,N_3633);
or U4723 (N_4723,N_3679,N_3987);
and U4724 (N_4724,N_3556,N_3637);
xor U4725 (N_4725,N_3462,N_3501);
or U4726 (N_4726,N_3969,N_3743);
or U4727 (N_4727,N_3027,N_3067);
nor U4728 (N_4728,N_3566,N_3540);
and U4729 (N_4729,N_3884,N_3435);
xnor U4730 (N_4730,N_3196,N_3612);
nor U4731 (N_4731,N_3238,N_3568);
or U4732 (N_4732,N_3198,N_3664);
or U4733 (N_4733,N_3317,N_3140);
and U4734 (N_4734,N_3450,N_3187);
nor U4735 (N_4735,N_3945,N_3289);
or U4736 (N_4736,N_3538,N_3349);
nor U4737 (N_4737,N_3343,N_3598);
nor U4738 (N_4738,N_3394,N_3890);
or U4739 (N_4739,N_3640,N_3968);
nand U4740 (N_4740,N_3284,N_3772);
nor U4741 (N_4741,N_3520,N_3712);
or U4742 (N_4742,N_3000,N_3890);
xor U4743 (N_4743,N_3898,N_3094);
nor U4744 (N_4744,N_3339,N_3402);
xnor U4745 (N_4745,N_3165,N_3031);
nor U4746 (N_4746,N_3482,N_3472);
and U4747 (N_4747,N_3204,N_3702);
nand U4748 (N_4748,N_3116,N_3062);
and U4749 (N_4749,N_3178,N_3611);
xnor U4750 (N_4750,N_3527,N_3307);
nor U4751 (N_4751,N_3676,N_3537);
nor U4752 (N_4752,N_3915,N_3271);
and U4753 (N_4753,N_3134,N_3865);
xnor U4754 (N_4754,N_3455,N_3718);
xor U4755 (N_4755,N_3839,N_3329);
nand U4756 (N_4756,N_3203,N_3025);
or U4757 (N_4757,N_3333,N_3182);
nor U4758 (N_4758,N_3797,N_3708);
nand U4759 (N_4759,N_3070,N_3098);
and U4760 (N_4760,N_3998,N_3536);
xnor U4761 (N_4761,N_3157,N_3993);
or U4762 (N_4762,N_3128,N_3810);
nand U4763 (N_4763,N_3461,N_3324);
and U4764 (N_4764,N_3746,N_3790);
nand U4765 (N_4765,N_3219,N_3169);
nand U4766 (N_4766,N_3302,N_3549);
nor U4767 (N_4767,N_3389,N_3879);
nor U4768 (N_4768,N_3559,N_3465);
nand U4769 (N_4769,N_3912,N_3198);
nor U4770 (N_4770,N_3191,N_3915);
or U4771 (N_4771,N_3682,N_3676);
and U4772 (N_4772,N_3816,N_3753);
xor U4773 (N_4773,N_3207,N_3592);
nand U4774 (N_4774,N_3211,N_3737);
nor U4775 (N_4775,N_3570,N_3646);
or U4776 (N_4776,N_3867,N_3312);
nor U4777 (N_4777,N_3138,N_3672);
nor U4778 (N_4778,N_3760,N_3584);
or U4779 (N_4779,N_3835,N_3412);
nor U4780 (N_4780,N_3554,N_3211);
and U4781 (N_4781,N_3794,N_3401);
nor U4782 (N_4782,N_3943,N_3514);
nor U4783 (N_4783,N_3966,N_3418);
or U4784 (N_4784,N_3016,N_3418);
or U4785 (N_4785,N_3907,N_3645);
nor U4786 (N_4786,N_3339,N_3268);
or U4787 (N_4787,N_3681,N_3174);
nand U4788 (N_4788,N_3317,N_3979);
or U4789 (N_4789,N_3318,N_3028);
xnor U4790 (N_4790,N_3365,N_3458);
or U4791 (N_4791,N_3592,N_3883);
and U4792 (N_4792,N_3629,N_3740);
nand U4793 (N_4793,N_3669,N_3964);
nor U4794 (N_4794,N_3314,N_3471);
xnor U4795 (N_4795,N_3279,N_3428);
nand U4796 (N_4796,N_3847,N_3046);
and U4797 (N_4797,N_3496,N_3096);
nand U4798 (N_4798,N_3084,N_3671);
and U4799 (N_4799,N_3223,N_3832);
nor U4800 (N_4800,N_3705,N_3043);
xor U4801 (N_4801,N_3543,N_3268);
and U4802 (N_4802,N_3681,N_3732);
or U4803 (N_4803,N_3807,N_3100);
or U4804 (N_4804,N_3805,N_3423);
nand U4805 (N_4805,N_3082,N_3643);
nor U4806 (N_4806,N_3529,N_3612);
and U4807 (N_4807,N_3068,N_3855);
nand U4808 (N_4808,N_3341,N_3690);
nand U4809 (N_4809,N_3130,N_3616);
nand U4810 (N_4810,N_3573,N_3472);
nor U4811 (N_4811,N_3854,N_3219);
nand U4812 (N_4812,N_3721,N_3864);
nand U4813 (N_4813,N_3154,N_3144);
and U4814 (N_4814,N_3002,N_3793);
and U4815 (N_4815,N_3596,N_3808);
xor U4816 (N_4816,N_3239,N_3287);
nor U4817 (N_4817,N_3901,N_3623);
and U4818 (N_4818,N_3173,N_3969);
nand U4819 (N_4819,N_3514,N_3891);
and U4820 (N_4820,N_3026,N_3555);
and U4821 (N_4821,N_3841,N_3738);
nand U4822 (N_4822,N_3843,N_3473);
or U4823 (N_4823,N_3738,N_3962);
nor U4824 (N_4824,N_3447,N_3790);
xor U4825 (N_4825,N_3729,N_3185);
and U4826 (N_4826,N_3607,N_3477);
nand U4827 (N_4827,N_3968,N_3694);
nor U4828 (N_4828,N_3240,N_3097);
xor U4829 (N_4829,N_3726,N_3708);
or U4830 (N_4830,N_3698,N_3092);
nor U4831 (N_4831,N_3272,N_3192);
and U4832 (N_4832,N_3445,N_3987);
and U4833 (N_4833,N_3641,N_3769);
and U4834 (N_4834,N_3560,N_3005);
and U4835 (N_4835,N_3642,N_3774);
nand U4836 (N_4836,N_3738,N_3954);
and U4837 (N_4837,N_3349,N_3200);
xnor U4838 (N_4838,N_3388,N_3506);
nand U4839 (N_4839,N_3911,N_3582);
and U4840 (N_4840,N_3595,N_3737);
and U4841 (N_4841,N_3284,N_3142);
and U4842 (N_4842,N_3488,N_3485);
nand U4843 (N_4843,N_3256,N_3213);
and U4844 (N_4844,N_3599,N_3756);
nor U4845 (N_4845,N_3919,N_3688);
and U4846 (N_4846,N_3909,N_3042);
xor U4847 (N_4847,N_3336,N_3720);
xor U4848 (N_4848,N_3848,N_3097);
or U4849 (N_4849,N_3090,N_3661);
xnor U4850 (N_4850,N_3868,N_3188);
nand U4851 (N_4851,N_3901,N_3590);
nor U4852 (N_4852,N_3589,N_3057);
or U4853 (N_4853,N_3087,N_3559);
nor U4854 (N_4854,N_3196,N_3271);
or U4855 (N_4855,N_3281,N_3593);
and U4856 (N_4856,N_3585,N_3460);
nor U4857 (N_4857,N_3908,N_3145);
or U4858 (N_4858,N_3549,N_3253);
nand U4859 (N_4859,N_3210,N_3471);
or U4860 (N_4860,N_3798,N_3897);
or U4861 (N_4861,N_3508,N_3482);
nand U4862 (N_4862,N_3634,N_3240);
xnor U4863 (N_4863,N_3342,N_3295);
nor U4864 (N_4864,N_3563,N_3985);
nor U4865 (N_4865,N_3949,N_3244);
nor U4866 (N_4866,N_3827,N_3919);
nor U4867 (N_4867,N_3878,N_3271);
nor U4868 (N_4868,N_3287,N_3514);
nor U4869 (N_4869,N_3318,N_3998);
xor U4870 (N_4870,N_3986,N_3303);
nand U4871 (N_4871,N_3952,N_3974);
nor U4872 (N_4872,N_3491,N_3686);
xor U4873 (N_4873,N_3695,N_3933);
or U4874 (N_4874,N_3344,N_3366);
nand U4875 (N_4875,N_3041,N_3221);
or U4876 (N_4876,N_3892,N_3955);
xnor U4877 (N_4877,N_3300,N_3705);
nor U4878 (N_4878,N_3848,N_3943);
or U4879 (N_4879,N_3396,N_3225);
nand U4880 (N_4880,N_3964,N_3115);
and U4881 (N_4881,N_3386,N_3458);
nand U4882 (N_4882,N_3312,N_3440);
xor U4883 (N_4883,N_3622,N_3205);
nor U4884 (N_4884,N_3097,N_3271);
or U4885 (N_4885,N_3770,N_3752);
nor U4886 (N_4886,N_3349,N_3583);
and U4887 (N_4887,N_3371,N_3292);
or U4888 (N_4888,N_3475,N_3385);
nand U4889 (N_4889,N_3753,N_3260);
nand U4890 (N_4890,N_3752,N_3090);
and U4891 (N_4891,N_3928,N_3313);
xor U4892 (N_4892,N_3404,N_3362);
nand U4893 (N_4893,N_3410,N_3232);
xnor U4894 (N_4894,N_3705,N_3105);
nor U4895 (N_4895,N_3491,N_3765);
or U4896 (N_4896,N_3546,N_3659);
or U4897 (N_4897,N_3494,N_3139);
and U4898 (N_4898,N_3771,N_3405);
or U4899 (N_4899,N_3312,N_3092);
nand U4900 (N_4900,N_3458,N_3430);
nand U4901 (N_4901,N_3550,N_3042);
xor U4902 (N_4902,N_3703,N_3267);
xor U4903 (N_4903,N_3758,N_3633);
nor U4904 (N_4904,N_3469,N_3690);
or U4905 (N_4905,N_3063,N_3443);
or U4906 (N_4906,N_3169,N_3327);
or U4907 (N_4907,N_3003,N_3478);
xnor U4908 (N_4908,N_3561,N_3549);
nand U4909 (N_4909,N_3409,N_3265);
or U4910 (N_4910,N_3389,N_3266);
nor U4911 (N_4911,N_3097,N_3677);
nor U4912 (N_4912,N_3616,N_3526);
nor U4913 (N_4913,N_3933,N_3465);
nor U4914 (N_4914,N_3100,N_3896);
nand U4915 (N_4915,N_3258,N_3039);
and U4916 (N_4916,N_3635,N_3572);
or U4917 (N_4917,N_3529,N_3799);
or U4918 (N_4918,N_3893,N_3246);
nor U4919 (N_4919,N_3542,N_3046);
nor U4920 (N_4920,N_3817,N_3610);
and U4921 (N_4921,N_3765,N_3277);
nand U4922 (N_4922,N_3601,N_3140);
nand U4923 (N_4923,N_3095,N_3808);
nor U4924 (N_4924,N_3978,N_3252);
and U4925 (N_4925,N_3618,N_3825);
or U4926 (N_4926,N_3244,N_3409);
nand U4927 (N_4927,N_3511,N_3417);
nand U4928 (N_4928,N_3995,N_3664);
and U4929 (N_4929,N_3206,N_3352);
nor U4930 (N_4930,N_3095,N_3207);
xor U4931 (N_4931,N_3378,N_3331);
nor U4932 (N_4932,N_3185,N_3700);
and U4933 (N_4933,N_3636,N_3037);
xor U4934 (N_4934,N_3175,N_3577);
nand U4935 (N_4935,N_3759,N_3128);
nor U4936 (N_4936,N_3706,N_3921);
nand U4937 (N_4937,N_3973,N_3447);
nand U4938 (N_4938,N_3820,N_3558);
and U4939 (N_4939,N_3374,N_3579);
and U4940 (N_4940,N_3110,N_3819);
and U4941 (N_4941,N_3462,N_3763);
nand U4942 (N_4942,N_3938,N_3208);
nor U4943 (N_4943,N_3392,N_3574);
nor U4944 (N_4944,N_3089,N_3320);
nand U4945 (N_4945,N_3600,N_3469);
xor U4946 (N_4946,N_3761,N_3615);
nor U4947 (N_4947,N_3214,N_3824);
and U4948 (N_4948,N_3525,N_3101);
nor U4949 (N_4949,N_3515,N_3719);
nand U4950 (N_4950,N_3511,N_3817);
nor U4951 (N_4951,N_3358,N_3235);
and U4952 (N_4952,N_3464,N_3098);
or U4953 (N_4953,N_3663,N_3371);
or U4954 (N_4954,N_3059,N_3720);
or U4955 (N_4955,N_3621,N_3133);
or U4956 (N_4956,N_3300,N_3809);
and U4957 (N_4957,N_3986,N_3707);
and U4958 (N_4958,N_3377,N_3688);
xnor U4959 (N_4959,N_3751,N_3232);
nand U4960 (N_4960,N_3774,N_3766);
nand U4961 (N_4961,N_3405,N_3470);
and U4962 (N_4962,N_3805,N_3752);
nand U4963 (N_4963,N_3126,N_3255);
or U4964 (N_4964,N_3222,N_3025);
and U4965 (N_4965,N_3501,N_3813);
and U4966 (N_4966,N_3964,N_3246);
or U4967 (N_4967,N_3819,N_3502);
and U4968 (N_4968,N_3123,N_3518);
xor U4969 (N_4969,N_3031,N_3888);
and U4970 (N_4970,N_3828,N_3869);
nand U4971 (N_4971,N_3206,N_3719);
or U4972 (N_4972,N_3716,N_3928);
nand U4973 (N_4973,N_3695,N_3246);
nor U4974 (N_4974,N_3896,N_3641);
xnor U4975 (N_4975,N_3933,N_3525);
and U4976 (N_4976,N_3570,N_3712);
nand U4977 (N_4977,N_3220,N_3068);
and U4978 (N_4978,N_3400,N_3524);
nor U4979 (N_4979,N_3012,N_3380);
and U4980 (N_4980,N_3335,N_3315);
or U4981 (N_4981,N_3823,N_3122);
nand U4982 (N_4982,N_3995,N_3295);
nor U4983 (N_4983,N_3264,N_3447);
nand U4984 (N_4984,N_3817,N_3409);
nand U4985 (N_4985,N_3612,N_3806);
or U4986 (N_4986,N_3996,N_3700);
or U4987 (N_4987,N_3788,N_3371);
and U4988 (N_4988,N_3868,N_3525);
or U4989 (N_4989,N_3705,N_3196);
nand U4990 (N_4990,N_3554,N_3873);
or U4991 (N_4991,N_3583,N_3228);
xor U4992 (N_4992,N_3598,N_3523);
xor U4993 (N_4993,N_3676,N_3465);
xnor U4994 (N_4994,N_3007,N_3617);
or U4995 (N_4995,N_3511,N_3789);
nor U4996 (N_4996,N_3268,N_3129);
nor U4997 (N_4997,N_3514,N_3328);
xor U4998 (N_4998,N_3407,N_3480);
nor U4999 (N_4999,N_3923,N_3370);
nor UO_0 (O_0,N_4809,N_4810);
xnor UO_1 (O_1,N_4413,N_4394);
nor UO_2 (O_2,N_4309,N_4705);
or UO_3 (O_3,N_4340,N_4134);
or UO_4 (O_4,N_4310,N_4876);
nand UO_5 (O_5,N_4797,N_4068);
nand UO_6 (O_6,N_4019,N_4192);
xnor UO_7 (O_7,N_4636,N_4556);
xnor UO_8 (O_8,N_4204,N_4040);
nor UO_9 (O_9,N_4376,N_4073);
xnor UO_10 (O_10,N_4072,N_4950);
nor UO_11 (O_11,N_4571,N_4238);
xor UO_12 (O_12,N_4869,N_4364);
and UO_13 (O_13,N_4349,N_4721);
xnor UO_14 (O_14,N_4841,N_4464);
nand UO_15 (O_15,N_4777,N_4021);
nand UO_16 (O_16,N_4664,N_4400);
and UO_17 (O_17,N_4739,N_4406);
nor UO_18 (O_18,N_4512,N_4768);
nor UO_19 (O_19,N_4829,N_4509);
nor UO_20 (O_20,N_4346,N_4493);
nand UO_21 (O_21,N_4297,N_4775);
and UO_22 (O_22,N_4578,N_4279);
nor UO_23 (O_23,N_4037,N_4295);
xor UO_24 (O_24,N_4332,N_4641);
and UO_25 (O_25,N_4685,N_4022);
and UO_26 (O_26,N_4202,N_4736);
xnor UO_27 (O_27,N_4363,N_4652);
and UO_28 (O_28,N_4534,N_4438);
nor UO_29 (O_29,N_4224,N_4890);
nand UO_30 (O_30,N_4393,N_4316);
or UO_31 (O_31,N_4947,N_4469);
and UO_32 (O_32,N_4697,N_4270);
nand UO_33 (O_33,N_4730,N_4712);
xnor UO_34 (O_34,N_4560,N_4563);
nand UO_35 (O_35,N_4517,N_4870);
or UO_36 (O_36,N_4350,N_4100);
or UO_37 (O_37,N_4344,N_4181);
xor UO_38 (O_38,N_4071,N_4503);
xor UO_39 (O_39,N_4672,N_4468);
nand UO_40 (O_40,N_4710,N_4959);
nor UO_41 (O_41,N_4137,N_4632);
and UO_42 (O_42,N_4006,N_4488);
or UO_43 (O_43,N_4035,N_4457);
nor UO_44 (O_44,N_4589,N_4814);
nand UO_45 (O_45,N_4616,N_4069);
xnor UO_46 (O_46,N_4348,N_4045);
and UO_47 (O_47,N_4405,N_4458);
and UO_48 (O_48,N_4859,N_4872);
nand UO_49 (O_49,N_4842,N_4601);
and UO_50 (O_50,N_4743,N_4253);
nor UO_51 (O_51,N_4545,N_4833);
and UO_52 (O_52,N_4983,N_4924);
nand UO_53 (O_53,N_4897,N_4764);
or UO_54 (O_54,N_4448,N_4934);
xnor UO_55 (O_55,N_4794,N_4081);
and UO_56 (O_56,N_4908,N_4343);
nand UO_57 (O_57,N_4276,N_4210);
xnor UO_58 (O_58,N_4803,N_4286);
or UO_59 (O_59,N_4533,N_4319);
or UO_60 (O_60,N_4709,N_4518);
xor UO_61 (O_61,N_4156,N_4133);
nand UO_62 (O_62,N_4942,N_4683);
and UO_63 (O_63,N_4757,N_4246);
or UO_64 (O_64,N_4805,N_4874);
nand UO_65 (O_65,N_4178,N_4886);
nor UO_66 (O_66,N_4956,N_4135);
nor UO_67 (O_67,N_4290,N_4561);
nand UO_68 (O_68,N_4419,N_4744);
or UO_69 (O_69,N_4409,N_4158);
nor UO_70 (O_70,N_4486,N_4108);
and UO_71 (O_71,N_4631,N_4226);
nand UO_72 (O_72,N_4639,N_4943);
nor UO_73 (O_73,N_4626,N_4701);
nand UO_74 (O_74,N_4434,N_4970);
or UO_75 (O_75,N_4583,N_4806);
and UO_76 (O_76,N_4926,N_4915);
nand UO_77 (O_77,N_4989,N_4369);
and UO_78 (O_78,N_4026,N_4440);
and UO_79 (O_79,N_4152,N_4746);
or UO_80 (O_80,N_4526,N_4304);
nand UO_81 (O_81,N_4058,N_4537);
nand UO_82 (O_82,N_4786,N_4592);
nor UO_83 (O_83,N_4665,N_4507);
and UO_84 (O_84,N_4816,N_4951);
nand UO_85 (O_85,N_4784,N_4031);
xor UO_86 (O_86,N_4716,N_4050);
or UO_87 (O_87,N_4195,N_4919);
and UO_88 (O_88,N_4427,N_4614);
xor UO_89 (O_89,N_4971,N_4234);
xnor UO_90 (O_90,N_4495,N_4769);
nand UO_91 (O_91,N_4837,N_4770);
or UO_92 (O_92,N_4048,N_4179);
nor UO_93 (O_93,N_4243,N_4149);
nor UO_94 (O_94,N_4525,N_4985);
nand UO_95 (O_95,N_4804,N_4162);
or UO_96 (O_96,N_4454,N_4142);
nand UO_97 (O_97,N_4387,N_4642);
nand UO_98 (O_98,N_4269,N_4686);
and UO_99 (O_99,N_4439,N_4548);
nor UO_100 (O_100,N_4868,N_4726);
and UO_101 (O_101,N_4939,N_4249);
or UO_102 (O_102,N_4496,N_4917);
or UO_103 (O_103,N_4096,N_4028);
and UO_104 (O_104,N_4586,N_4622);
nor UO_105 (O_105,N_4085,N_4873);
or UO_106 (O_106,N_4186,N_4030);
nor UO_107 (O_107,N_4783,N_4266);
nor UO_108 (O_108,N_4718,N_4000);
nor UO_109 (O_109,N_4264,N_4843);
nor UO_110 (O_110,N_4090,N_4717);
or UO_111 (O_111,N_4511,N_4161);
or UO_112 (O_112,N_4729,N_4492);
or UO_113 (O_113,N_4103,N_4542);
nor UO_114 (O_114,N_4954,N_4354);
nand UO_115 (O_115,N_4018,N_4447);
nor UO_116 (O_116,N_4044,N_4758);
nand UO_117 (O_117,N_4347,N_4127);
nor UO_118 (O_118,N_4884,N_4339);
nand UO_119 (O_119,N_4235,N_4504);
nand UO_120 (O_120,N_4274,N_4682);
or UO_121 (O_121,N_4898,N_4748);
nand UO_122 (O_122,N_4046,N_4587);
and UO_123 (O_123,N_4728,N_4909);
xor UO_124 (O_124,N_4061,N_4039);
nor UO_125 (O_125,N_4255,N_4719);
nor UO_126 (O_126,N_4042,N_4452);
nand UO_127 (O_127,N_4793,N_4017);
or UO_128 (O_128,N_4139,N_4341);
nor UO_129 (O_129,N_4706,N_4153);
or UO_130 (O_130,N_4315,N_4836);
and UO_131 (O_131,N_4593,N_4596);
xnor UO_132 (O_132,N_4602,N_4301);
nand UO_133 (O_133,N_4386,N_4051);
nand UO_134 (O_134,N_4351,N_4568);
or UO_135 (O_135,N_4015,N_4569);
or UO_136 (O_136,N_4429,N_4375);
nor UO_137 (O_137,N_4254,N_4145);
and UO_138 (O_138,N_4661,N_4215);
nor UO_139 (O_139,N_4272,N_4043);
and UO_140 (O_140,N_4328,N_4656);
and UO_141 (O_141,N_4407,N_4207);
and UO_142 (O_142,N_4727,N_4013);
nand UO_143 (O_143,N_4117,N_4763);
nand UO_144 (O_144,N_4443,N_4107);
nor UO_145 (O_145,N_4092,N_4180);
or UO_146 (O_146,N_4994,N_4595);
or UO_147 (O_147,N_4062,N_4978);
or UO_148 (O_148,N_4907,N_4016);
nor UO_149 (O_149,N_4654,N_4681);
nand UO_150 (O_150,N_4047,N_4307);
xor UO_151 (O_151,N_4846,N_4505);
xor UO_152 (O_152,N_4412,N_4223);
nand UO_153 (O_153,N_4766,N_4535);
nor UO_154 (O_154,N_4649,N_4080);
nor UO_155 (O_155,N_4337,N_4508);
and UO_156 (O_156,N_4009,N_4968);
nor UO_157 (O_157,N_4183,N_4762);
and UO_158 (O_158,N_4388,N_4314);
or UO_159 (O_159,N_4840,N_4300);
or UO_160 (O_160,N_4360,N_4657);
nand UO_161 (O_161,N_4860,N_4482);
nand UO_162 (O_162,N_4818,N_4123);
or UO_163 (O_163,N_4361,N_4263);
and UO_164 (O_164,N_4609,N_4577);
nor UO_165 (O_165,N_4737,N_4640);
or UO_166 (O_166,N_4077,N_4871);
xor UO_167 (O_167,N_4572,N_4828);
nand UO_168 (O_168,N_4421,N_4402);
and UO_169 (O_169,N_4713,N_4695);
and UO_170 (O_170,N_4693,N_4932);
nand UO_171 (O_171,N_4455,N_4168);
nand UO_172 (O_172,N_4115,N_4335);
nor UO_173 (O_173,N_4410,N_4403);
nor UO_174 (O_174,N_4952,N_4197);
nand UO_175 (O_175,N_4506,N_4397);
nor UO_176 (O_176,N_4064,N_4558);
nand UO_177 (O_177,N_4703,N_4617);
xor UO_178 (O_178,N_4381,N_4536);
nand UO_179 (O_179,N_4054,N_4882);
and UO_180 (O_180,N_4355,N_4819);
or UO_181 (O_181,N_4240,N_4753);
xor UO_182 (O_182,N_4895,N_4430);
or UO_183 (O_183,N_4707,N_4383);
nand UO_184 (O_184,N_4555,N_4257);
and UO_185 (O_185,N_4441,N_4544);
or UO_186 (O_186,N_4480,N_4415);
or UO_187 (O_187,N_4052,N_4151);
or UO_188 (O_188,N_4591,N_4754);
nor UO_189 (O_189,N_4620,N_4327);
and UO_190 (O_190,N_4305,N_4832);
nand UO_191 (O_191,N_4750,N_4060);
or UO_192 (O_192,N_4524,N_4476);
and UO_193 (O_193,N_4459,N_4838);
nand UO_194 (O_194,N_4651,N_4792);
nor UO_195 (O_195,N_4673,N_4170);
nor UO_196 (O_196,N_4949,N_4174);
and UO_197 (O_197,N_4093,N_4352);
or UO_198 (O_198,N_4193,N_4288);
nor UO_199 (O_199,N_4883,N_4755);
or UO_200 (O_200,N_4724,N_4416);
nand UO_201 (O_201,N_4998,N_4600);
nor UO_202 (O_202,N_4230,N_4513);
nand UO_203 (O_203,N_4848,N_4365);
and UO_204 (O_204,N_4236,N_4975);
nor UO_205 (O_205,N_4723,N_4888);
nand UO_206 (O_206,N_4114,N_4936);
xnor UO_207 (O_207,N_4188,N_4138);
and UO_208 (O_208,N_4611,N_4689);
nand UO_209 (O_209,N_4277,N_4958);
nand UO_210 (O_210,N_4191,N_4782);
nor UO_211 (O_211,N_4390,N_4258);
or UO_212 (O_212,N_4708,N_4466);
nand UO_213 (O_213,N_4324,N_4678);
and UO_214 (O_214,N_4920,N_4527);
or UO_215 (O_215,N_4112,N_4911);
nor UO_216 (O_216,N_4899,N_4219);
nand UO_217 (O_217,N_4567,N_4646);
and UO_218 (O_218,N_4231,N_4465);
or UO_219 (O_219,N_4627,N_4916);
or UO_220 (O_220,N_4399,N_4481);
and UO_221 (O_221,N_4218,N_4696);
nand UO_222 (O_222,N_4008,N_4095);
nand UO_223 (O_223,N_4576,N_4863);
nand UO_224 (O_224,N_4906,N_4529);
nor UO_225 (O_225,N_4357,N_4359);
nand UO_226 (O_226,N_4182,N_4725);
or UO_227 (O_227,N_4342,N_4613);
nand UO_228 (O_228,N_4580,N_4931);
nor UO_229 (O_229,N_4960,N_4785);
and UO_230 (O_230,N_4171,N_4029);
or UO_231 (O_231,N_4323,N_4756);
nor UO_232 (O_232,N_4554,N_4515);
nand UO_233 (O_233,N_4918,N_4281);
or UO_234 (O_234,N_4902,N_4293);
and UO_235 (O_235,N_4292,N_4317);
and UO_236 (O_236,N_4540,N_4519);
nand UO_237 (O_237,N_4878,N_4821);
or UO_238 (O_238,N_4087,N_4634);
or UO_239 (O_239,N_4606,N_4699);
nor UO_240 (O_240,N_4165,N_4528);
nand UO_241 (O_241,N_4088,N_4287);
xor UO_242 (O_242,N_4126,N_4865);
nand UO_243 (O_243,N_4904,N_4166);
nor UO_244 (O_244,N_4221,N_4996);
nand UO_245 (O_245,N_4033,N_4857);
xnor UO_246 (O_246,N_4391,N_4638);
nor UO_247 (O_247,N_4885,N_4067);
nand UO_248 (O_248,N_4745,N_4167);
or UO_249 (O_249,N_4377,N_4720);
nand UO_250 (O_250,N_4209,N_4834);
nand UO_251 (O_251,N_4928,N_4624);
and UO_252 (O_252,N_4698,N_4581);
nor UO_253 (O_253,N_4608,N_4575);
or UO_254 (O_254,N_4296,N_4120);
xor UO_255 (O_255,N_4371,N_4680);
nand UO_256 (O_256,N_4946,N_4500);
or UO_257 (O_257,N_4494,N_4423);
nor UO_258 (O_258,N_4237,N_4099);
xnor UO_259 (O_259,N_4861,N_4847);
or UO_260 (O_260,N_4278,N_4366);
and UO_261 (O_261,N_4590,N_4539);
nand UO_262 (O_262,N_4131,N_4815);
nand UO_263 (O_263,N_4795,N_4345);
xor UO_264 (O_264,N_4972,N_4749);
and UO_265 (O_265,N_4128,N_4944);
nand UO_266 (O_266,N_4232,N_4222);
nand UO_267 (O_267,N_4245,N_4294);
nand UO_268 (O_268,N_4176,N_4914);
nand UO_269 (O_269,N_4905,N_4903);
and UO_270 (O_270,N_4483,N_4227);
or UO_271 (O_271,N_4303,N_4066);
xor UO_272 (O_272,N_4273,N_4368);
or UO_273 (O_273,N_4005,N_4957);
nand UO_274 (O_274,N_4082,N_4160);
nand UO_275 (O_275,N_4489,N_4267);
and UO_276 (O_276,N_4014,N_4940);
or UO_277 (O_277,N_4825,N_4499);
nand UO_278 (O_278,N_4731,N_4658);
and UO_279 (O_279,N_4389,N_4420);
nor UO_280 (O_280,N_4562,N_4585);
nor UO_281 (O_281,N_4200,N_4738);
and UO_282 (O_282,N_4433,N_4676);
and UO_283 (O_283,N_4850,N_4852);
or UO_284 (O_284,N_4933,N_4119);
nand UO_285 (O_285,N_4262,N_4598);
nand UO_286 (O_286,N_4648,N_4930);
or UO_287 (O_287,N_4311,N_4086);
or UO_288 (O_288,N_4011,N_4485);
and UO_289 (O_289,N_4788,N_4291);
or UO_290 (O_290,N_4491,N_4650);
and UO_291 (O_291,N_4362,N_4663);
nand UO_292 (O_292,N_4955,N_4751);
nor UO_293 (O_293,N_4333,N_4426);
or UO_294 (O_294,N_4104,N_4655);
and UO_295 (O_295,N_4514,N_4189);
nand UO_296 (O_296,N_4472,N_4887);
nand UO_297 (O_297,N_4789,N_4004);
or UO_298 (O_298,N_4625,N_4945);
or UO_299 (O_299,N_4981,N_4835);
and UO_300 (O_300,N_4704,N_4523);
nand UO_301 (O_301,N_4025,N_4564);
nor UO_302 (O_302,N_4845,N_4306);
nand UO_303 (O_303,N_4367,N_4557);
nor UO_304 (O_304,N_4194,N_4284);
nand UO_305 (O_305,N_4089,N_4445);
nand UO_306 (O_306,N_4830,N_4125);
nand UO_307 (O_307,N_4164,N_4147);
or UO_308 (O_308,N_4338,N_4831);
and UO_309 (O_309,N_4817,N_4356);
nand UO_310 (O_310,N_4358,N_4570);
or UO_311 (O_311,N_4594,N_4501);
or UO_312 (O_312,N_4490,N_4922);
nand UO_313 (O_313,N_4057,N_4864);
and UO_314 (O_314,N_4644,N_4732);
and UO_315 (O_315,N_4444,N_4618);
nand UO_316 (O_316,N_4002,N_4690);
nor UO_317 (O_317,N_4453,N_4032);
nor UO_318 (O_318,N_4879,N_4599);
nor UO_319 (O_319,N_4964,N_4113);
or UO_320 (O_320,N_4110,N_4118);
and UO_321 (O_321,N_4612,N_4036);
xnor UO_322 (O_322,N_4479,N_4662);
nor UO_323 (O_323,N_4551,N_4992);
and UO_324 (O_324,N_4984,N_4948);
xor UO_325 (O_325,N_4844,N_4007);
and UO_326 (O_326,N_4659,N_4605);
and UO_327 (O_327,N_4761,N_4619);
xnor UO_328 (O_328,N_4382,N_4097);
or UO_329 (O_329,N_4823,N_4549);
and UO_330 (O_330,N_4299,N_4318);
nand UO_331 (O_331,N_4122,N_4734);
or UO_332 (O_332,N_4900,N_4408);
nand UO_333 (O_333,N_4079,N_4778);
nand UO_334 (O_334,N_4385,N_4552);
nand UO_335 (O_335,N_4893,N_4531);
and UO_336 (O_336,N_4866,N_4855);
or UO_337 (O_337,N_4321,N_4623);
and UO_338 (O_338,N_4302,N_4993);
nand UO_339 (O_339,N_4628,N_4203);
or UO_340 (O_340,N_4779,N_4858);
nor UO_341 (O_341,N_4688,N_4177);
nor UO_342 (O_342,N_4839,N_4941);
xnor UO_343 (O_343,N_4694,N_4330);
or UO_344 (O_344,N_4812,N_4742);
and UO_345 (O_345,N_4056,N_4473);
nand UO_346 (O_346,N_4208,N_4228);
xnor UO_347 (O_347,N_4670,N_4320);
nor UO_348 (O_348,N_4937,N_4083);
nand UO_349 (O_349,N_4862,N_4607);
or UO_350 (O_350,N_4132,N_4313);
and UO_351 (O_351,N_4038,N_4251);
and UO_352 (O_352,N_4669,N_4691);
and UO_353 (O_353,N_4331,N_4312);
or UO_354 (O_354,N_4935,N_4070);
and UO_355 (O_355,N_4962,N_4653);
xnor UO_356 (O_356,N_4881,N_4961);
and UO_357 (O_357,N_4484,N_4813);
or UO_358 (O_358,N_4379,N_4065);
and UO_359 (O_359,N_4787,N_4411);
nand UO_360 (O_360,N_4102,N_4275);
and UO_361 (O_361,N_4880,N_4715);
or UO_362 (O_362,N_4965,N_4449);
and UO_363 (O_363,N_4425,N_4169);
nand UO_364 (O_364,N_4635,N_4136);
nor UO_365 (O_365,N_4790,N_4807);
xnor UO_366 (O_366,N_4395,N_4767);
or UO_367 (O_367,N_4521,N_4001);
and UO_368 (O_368,N_4213,N_4667);
and UO_369 (O_369,N_4773,N_4925);
xnor UO_370 (O_370,N_4559,N_4820);
or UO_371 (O_371,N_4435,N_4211);
nor UO_372 (O_372,N_4326,N_4111);
and UO_373 (O_373,N_4280,N_4700);
xnor UO_374 (O_374,N_4666,N_4159);
nor UO_375 (O_375,N_4353,N_4239);
nor UO_376 (O_376,N_4765,N_4094);
xor UO_377 (O_377,N_4173,N_4024);
nor UO_378 (O_378,N_4442,N_4010);
or UO_379 (O_379,N_4760,N_4157);
and UO_380 (O_380,N_4702,N_4546);
nor UO_381 (O_381,N_4692,N_4212);
nand UO_382 (O_382,N_4621,N_4146);
nor UO_383 (O_383,N_4629,N_4078);
or UO_384 (O_384,N_4241,N_4822);
nand UO_385 (O_385,N_4285,N_4252);
xor UO_386 (O_386,N_4630,N_4982);
xnor UO_387 (O_387,N_4660,N_4380);
or UO_388 (O_388,N_4023,N_4053);
nand UO_389 (O_389,N_4225,N_4428);
xnor UO_390 (O_390,N_4198,N_4986);
and UO_391 (O_391,N_4901,N_4456);
nand UO_392 (O_392,N_4049,N_4205);
and UO_393 (O_393,N_4913,N_4076);
nor UO_394 (O_394,N_4130,N_4808);
nand UO_395 (O_395,N_4796,N_4196);
nand UO_396 (O_396,N_4260,N_4896);
nand UO_397 (O_397,N_4877,N_4547);
and UO_398 (O_398,N_4974,N_4637);
or UO_399 (O_399,N_4853,N_4741);
and UO_400 (O_400,N_4261,N_4522);
xor UO_401 (O_401,N_4436,N_4163);
nand UO_402 (O_402,N_4991,N_4584);
nor UO_403 (O_403,N_4470,N_4990);
and UO_404 (O_404,N_4398,N_4265);
and UO_405 (O_405,N_4217,N_4214);
nand UO_406 (O_406,N_4530,N_4668);
nand UO_407 (O_407,N_4116,N_4184);
nor UO_408 (O_408,N_4322,N_4516);
nor UO_409 (O_409,N_4502,N_4573);
or UO_410 (O_410,N_4610,N_4541);
and UO_411 (O_411,N_4474,N_4334);
and UO_412 (O_412,N_4802,N_4124);
and UO_413 (O_413,N_4098,N_4677);
nand UO_414 (O_414,N_4074,N_4461);
nand UO_415 (O_415,N_4109,N_4256);
nor UO_416 (O_416,N_4140,N_4520);
and UO_417 (O_417,N_4774,N_4929);
or UO_418 (O_418,N_4772,N_4336);
or UO_419 (O_419,N_4759,N_4675);
and UO_420 (O_420,N_4432,N_4910);
and UO_421 (O_421,N_4271,N_4477);
or UO_422 (O_422,N_4953,N_4150);
and UO_423 (O_423,N_4875,N_4997);
nand UO_424 (O_424,N_4565,N_4671);
and UO_425 (O_425,N_4121,N_4987);
or UO_426 (O_426,N_4771,N_4988);
nor UO_427 (O_427,N_4892,N_4851);
and UO_428 (O_428,N_4967,N_4976);
and UO_429 (O_429,N_4282,N_4973);
or UO_430 (O_430,N_4129,N_4063);
and UO_431 (O_431,N_4034,N_4467);
or UO_432 (O_432,N_4687,N_4475);
or UO_433 (O_433,N_4424,N_4041);
nand UO_434 (O_434,N_4615,N_4201);
nand UO_435 (O_435,N_4417,N_4259);
nor UO_436 (O_436,N_4824,N_4604);
or UO_437 (O_437,N_4776,N_4487);
nand UO_438 (O_438,N_4020,N_4370);
nor UO_439 (O_439,N_4141,N_4781);
and UO_440 (O_440,N_4206,N_4172);
nand UO_441 (O_441,N_4921,N_4233);
and UO_442 (O_442,N_4220,N_4867);
nand UO_443 (O_443,N_4229,N_4396);
nand UO_444 (O_444,N_4055,N_4498);
or UO_445 (O_445,N_4999,N_4553);
and UO_446 (O_446,N_4392,N_4298);
or UO_447 (O_447,N_4801,N_4827);
nor UO_448 (O_448,N_4977,N_4923);
nor UO_449 (O_449,N_4187,N_4579);
nand UO_450 (O_450,N_4574,N_4268);
or UO_451 (O_451,N_4144,N_4714);
or UO_452 (O_452,N_4437,N_4404);
nor UO_453 (O_453,N_4752,N_4374);
and UO_454 (O_454,N_4711,N_4105);
and UO_455 (O_455,N_4740,N_4422);
and UO_456 (O_456,N_4603,N_4643);
nand UO_457 (O_457,N_4154,N_4543);
and UO_458 (O_458,N_4927,N_4283);
nor UO_459 (O_459,N_4969,N_4849);
and UO_460 (O_460,N_4460,N_4471);
nor UO_461 (O_461,N_4532,N_4247);
and UO_462 (O_462,N_4155,N_4373);
nand UO_463 (O_463,N_4003,N_4735);
nand UO_464 (O_464,N_4431,N_4566);
or UO_465 (O_465,N_4582,N_4185);
nor UO_466 (O_466,N_4633,N_4550);
xnor UO_467 (O_467,N_4242,N_4679);
nor UO_468 (O_468,N_4084,N_4647);
xnor UO_469 (O_469,N_4106,N_4012);
and UO_470 (O_470,N_4497,N_4175);
or UO_471 (O_471,N_4384,N_4462);
nor UO_472 (O_472,N_4889,N_4190);
and UO_473 (O_473,N_4478,N_4463);
nor UO_474 (O_474,N_4091,N_4588);
or UO_475 (O_475,N_4101,N_4811);
or UO_476 (O_476,N_4966,N_4674);
nor UO_477 (O_477,N_4645,N_4289);
or UO_478 (O_478,N_4059,N_4826);
nor UO_479 (O_479,N_4722,N_4378);
nor UO_480 (O_480,N_4250,N_4372);
nand UO_481 (O_481,N_4148,N_4248);
nor UO_482 (O_482,N_4894,N_4510);
or UO_483 (O_483,N_4199,N_4938);
nor UO_484 (O_484,N_4747,N_4798);
and UO_485 (O_485,N_4980,N_4597);
or UO_486 (O_486,N_4244,N_4780);
and UO_487 (O_487,N_4684,N_4143);
or UO_488 (O_488,N_4414,N_4401);
nor UO_489 (O_489,N_4451,N_4733);
nand UO_490 (O_490,N_4891,N_4799);
nand UO_491 (O_491,N_4963,N_4791);
xor UO_492 (O_492,N_4854,N_4329);
and UO_493 (O_493,N_4325,N_4538);
and UO_494 (O_494,N_4216,N_4995);
and UO_495 (O_495,N_4912,N_4418);
or UO_496 (O_496,N_4450,N_4800);
or UO_497 (O_497,N_4979,N_4308);
or UO_498 (O_498,N_4856,N_4075);
nor UO_499 (O_499,N_4027,N_4446);
xnor UO_500 (O_500,N_4800,N_4296);
and UO_501 (O_501,N_4836,N_4612);
or UO_502 (O_502,N_4987,N_4626);
or UO_503 (O_503,N_4666,N_4417);
and UO_504 (O_504,N_4485,N_4389);
or UO_505 (O_505,N_4327,N_4953);
xor UO_506 (O_506,N_4717,N_4378);
nor UO_507 (O_507,N_4522,N_4211);
nor UO_508 (O_508,N_4595,N_4300);
and UO_509 (O_509,N_4069,N_4204);
nand UO_510 (O_510,N_4325,N_4037);
or UO_511 (O_511,N_4964,N_4485);
or UO_512 (O_512,N_4057,N_4373);
xor UO_513 (O_513,N_4194,N_4962);
and UO_514 (O_514,N_4022,N_4593);
nor UO_515 (O_515,N_4618,N_4039);
and UO_516 (O_516,N_4729,N_4066);
nand UO_517 (O_517,N_4852,N_4835);
nand UO_518 (O_518,N_4488,N_4651);
xnor UO_519 (O_519,N_4195,N_4390);
nor UO_520 (O_520,N_4272,N_4566);
xnor UO_521 (O_521,N_4758,N_4753);
nor UO_522 (O_522,N_4413,N_4030);
or UO_523 (O_523,N_4553,N_4902);
nand UO_524 (O_524,N_4529,N_4467);
or UO_525 (O_525,N_4889,N_4159);
and UO_526 (O_526,N_4282,N_4019);
nand UO_527 (O_527,N_4346,N_4516);
nand UO_528 (O_528,N_4287,N_4933);
or UO_529 (O_529,N_4448,N_4127);
nor UO_530 (O_530,N_4781,N_4519);
nand UO_531 (O_531,N_4625,N_4853);
nand UO_532 (O_532,N_4826,N_4270);
nand UO_533 (O_533,N_4160,N_4642);
or UO_534 (O_534,N_4353,N_4776);
nor UO_535 (O_535,N_4708,N_4040);
or UO_536 (O_536,N_4983,N_4075);
or UO_537 (O_537,N_4642,N_4831);
or UO_538 (O_538,N_4239,N_4527);
xnor UO_539 (O_539,N_4469,N_4020);
nand UO_540 (O_540,N_4803,N_4556);
and UO_541 (O_541,N_4126,N_4798);
and UO_542 (O_542,N_4536,N_4950);
nor UO_543 (O_543,N_4376,N_4602);
xnor UO_544 (O_544,N_4402,N_4432);
nand UO_545 (O_545,N_4754,N_4549);
nand UO_546 (O_546,N_4670,N_4286);
and UO_547 (O_547,N_4643,N_4997);
or UO_548 (O_548,N_4049,N_4587);
nand UO_549 (O_549,N_4528,N_4949);
and UO_550 (O_550,N_4709,N_4306);
nand UO_551 (O_551,N_4086,N_4194);
nand UO_552 (O_552,N_4114,N_4338);
nand UO_553 (O_553,N_4151,N_4390);
nor UO_554 (O_554,N_4750,N_4986);
or UO_555 (O_555,N_4733,N_4962);
nand UO_556 (O_556,N_4318,N_4968);
nand UO_557 (O_557,N_4938,N_4371);
and UO_558 (O_558,N_4632,N_4866);
and UO_559 (O_559,N_4660,N_4457);
and UO_560 (O_560,N_4478,N_4584);
xnor UO_561 (O_561,N_4223,N_4673);
xnor UO_562 (O_562,N_4388,N_4746);
nand UO_563 (O_563,N_4509,N_4790);
and UO_564 (O_564,N_4918,N_4502);
nor UO_565 (O_565,N_4257,N_4263);
and UO_566 (O_566,N_4895,N_4321);
nand UO_567 (O_567,N_4024,N_4434);
and UO_568 (O_568,N_4689,N_4161);
nor UO_569 (O_569,N_4495,N_4878);
or UO_570 (O_570,N_4119,N_4804);
and UO_571 (O_571,N_4631,N_4213);
or UO_572 (O_572,N_4347,N_4134);
nor UO_573 (O_573,N_4387,N_4234);
xor UO_574 (O_574,N_4162,N_4925);
xor UO_575 (O_575,N_4259,N_4822);
nand UO_576 (O_576,N_4133,N_4382);
nand UO_577 (O_577,N_4972,N_4127);
and UO_578 (O_578,N_4568,N_4359);
or UO_579 (O_579,N_4190,N_4007);
nor UO_580 (O_580,N_4543,N_4736);
xor UO_581 (O_581,N_4358,N_4517);
or UO_582 (O_582,N_4539,N_4531);
or UO_583 (O_583,N_4256,N_4448);
nand UO_584 (O_584,N_4696,N_4268);
nand UO_585 (O_585,N_4539,N_4158);
nand UO_586 (O_586,N_4483,N_4342);
and UO_587 (O_587,N_4131,N_4631);
or UO_588 (O_588,N_4370,N_4210);
or UO_589 (O_589,N_4958,N_4454);
nor UO_590 (O_590,N_4157,N_4064);
or UO_591 (O_591,N_4591,N_4054);
and UO_592 (O_592,N_4577,N_4087);
nor UO_593 (O_593,N_4984,N_4344);
xnor UO_594 (O_594,N_4472,N_4310);
or UO_595 (O_595,N_4778,N_4665);
nand UO_596 (O_596,N_4451,N_4293);
nor UO_597 (O_597,N_4525,N_4341);
and UO_598 (O_598,N_4633,N_4987);
xnor UO_599 (O_599,N_4636,N_4689);
and UO_600 (O_600,N_4351,N_4471);
or UO_601 (O_601,N_4528,N_4088);
and UO_602 (O_602,N_4052,N_4559);
xnor UO_603 (O_603,N_4405,N_4795);
and UO_604 (O_604,N_4778,N_4794);
and UO_605 (O_605,N_4149,N_4170);
nor UO_606 (O_606,N_4278,N_4828);
and UO_607 (O_607,N_4901,N_4084);
nor UO_608 (O_608,N_4520,N_4538);
and UO_609 (O_609,N_4928,N_4367);
nor UO_610 (O_610,N_4959,N_4015);
xor UO_611 (O_611,N_4545,N_4476);
or UO_612 (O_612,N_4383,N_4441);
and UO_613 (O_613,N_4146,N_4524);
nor UO_614 (O_614,N_4662,N_4752);
nand UO_615 (O_615,N_4584,N_4792);
nor UO_616 (O_616,N_4951,N_4691);
and UO_617 (O_617,N_4133,N_4735);
xor UO_618 (O_618,N_4933,N_4498);
nor UO_619 (O_619,N_4163,N_4440);
and UO_620 (O_620,N_4905,N_4818);
nand UO_621 (O_621,N_4495,N_4872);
xnor UO_622 (O_622,N_4062,N_4423);
and UO_623 (O_623,N_4412,N_4395);
nand UO_624 (O_624,N_4545,N_4255);
and UO_625 (O_625,N_4246,N_4417);
or UO_626 (O_626,N_4211,N_4322);
and UO_627 (O_627,N_4264,N_4778);
nand UO_628 (O_628,N_4087,N_4662);
xor UO_629 (O_629,N_4863,N_4403);
nand UO_630 (O_630,N_4755,N_4307);
or UO_631 (O_631,N_4965,N_4591);
nand UO_632 (O_632,N_4060,N_4204);
nor UO_633 (O_633,N_4087,N_4393);
and UO_634 (O_634,N_4644,N_4401);
or UO_635 (O_635,N_4038,N_4233);
and UO_636 (O_636,N_4925,N_4758);
xnor UO_637 (O_637,N_4788,N_4572);
or UO_638 (O_638,N_4838,N_4371);
and UO_639 (O_639,N_4484,N_4427);
nand UO_640 (O_640,N_4363,N_4163);
or UO_641 (O_641,N_4976,N_4496);
and UO_642 (O_642,N_4683,N_4336);
and UO_643 (O_643,N_4266,N_4516);
or UO_644 (O_644,N_4398,N_4823);
or UO_645 (O_645,N_4439,N_4905);
nand UO_646 (O_646,N_4485,N_4531);
nand UO_647 (O_647,N_4050,N_4003);
or UO_648 (O_648,N_4945,N_4947);
xnor UO_649 (O_649,N_4524,N_4279);
nor UO_650 (O_650,N_4999,N_4425);
and UO_651 (O_651,N_4795,N_4431);
and UO_652 (O_652,N_4408,N_4809);
or UO_653 (O_653,N_4817,N_4202);
or UO_654 (O_654,N_4511,N_4367);
nand UO_655 (O_655,N_4205,N_4553);
nor UO_656 (O_656,N_4446,N_4881);
nor UO_657 (O_657,N_4009,N_4054);
and UO_658 (O_658,N_4169,N_4392);
xnor UO_659 (O_659,N_4221,N_4236);
or UO_660 (O_660,N_4917,N_4467);
nand UO_661 (O_661,N_4270,N_4096);
nand UO_662 (O_662,N_4366,N_4177);
and UO_663 (O_663,N_4805,N_4516);
xor UO_664 (O_664,N_4981,N_4654);
and UO_665 (O_665,N_4117,N_4904);
nand UO_666 (O_666,N_4338,N_4415);
nand UO_667 (O_667,N_4090,N_4102);
xnor UO_668 (O_668,N_4364,N_4555);
nor UO_669 (O_669,N_4208,N_4365);
and UO_670 (O_670,N_4584,N_4580);
nor UO_671 (O_671,N_4088,N_4514);
or UO_672 (O_672,N_4884,N_4105);
and UO_673 (O_673,N_4230,N_4730);
nor UO_674 (O_674,N_4909,N_4089);
or UO_675 (O_675,N_4816,N_4658);
and UO_676 (O_676,N_4373,N_4018);
nor UO_677 (O_677,N_4369,N_4828);
nor UO_678 (O_678,N_4542,N_4001);
nand UO_679 (O_679,N_4947,N_4214);
nor UO_680 (O_680,N_4466,N_4350);
nor UO_681 (O_681,N_4292,N_4372);
nor UO_682 (O_682,N_4675,N_4761);
and UO_683 (O_683,N_4342,N_4335);
and UO_684 (O_684,N_4351,N_4763);
nor UO_685 (O_685,N_4959,N_4519);
nor UO_686 (O_686,N_4727,N_4907);
nor UO_687 (O_687,N_4963,N_4458);
or UO_688 (O_688,N_4609,N_4830);
and UO_689 (O_689,N_4065,N_4206);
nand UO_690 (O_690,N_4616,N_4527);
or UO_691 (O_691,N_4588,N_4906);
and UO_692 (O_692,N_4786,N_4132);
or UO_693 (O_693,N_4946,N_4236);
nand UO_694 (O_694,N_4590,N_4534);
and UO_695 (O_695,N_4947,N_4794);
nand UO_696 (O_696,N_4531,N_4721);
nand UO_697 (O_697,N_4729,N_4705);
nor UO_698 (O_698,N_4332,N_4669);
and UO_699 (O_699,N_4378,N_4069);
or UO_700 (O_700,N_4118,N_4952);
nor UO_701 (O_701,N_4653,N_4235);
nand UO_702 (O_702,N_4012,N_4265);
and UO_703 (O_703,N_4621,N_4228);
nand UO_704 (O_704,N_4446,N_4667);
nor UO_705 (O_705,N_4085,N_4134);
nor UO_706 (O_706,N_4657,N_4252);
or UO_707 (O_707,N_4359,N_4165);
nand UO_708 (O_708,N_4294,N_4187);
nor UO_709 (O_709,N_4993,N_4751);
nand UO_710 (O_710,N_4572,N_4700);
and UO_711 (O_711,N_4835,N_4815);
nor UO_712 (O_712,N_4648,N_4378);
nor UO_713 (O_713,N_4590,N_4470);
or UO_714 (O_714,N_4899,N_4374);
xnor UO_715 (O_715,N_4776,N_4367);
or UO_716 (O_716,N_4671,N_4211);
or UO_717 (O_717,N_4211,N_4950);
nor UO_718 (O_718,N_4737,N_4481);
nor UO_719 (O_719,N_4948,N_4869);
nor UO_720 (O_720,N_4042,N_4783);
or UO_721 (O_721,N_4761,N_4098);
and UO_722 (O_722,N_4100,N_4482);
nand UO_723 (O_723,N_4528,N_4890);
or UO_724 (O_724,N_4579,N_4982);
and UO_725 (O_725,N_4780,N_4097);
nand UO_726 (O_726,N_4420,N_4654);
nand UO_727 (O_727,N_4421,N_4878);
or UO_728 (O_728,N_4006,N_4027);
nor UO_729 (O_729,N_4831,N_4128);
xor UO_730 (O_730,N_4528,N_4197);
or UO_731 (O_731,N_4092,N_4192);
nor UO_732 (O_732,N_4069,N_4647);
xor UO_733 (O_733,N_4733,N_4331);
xnor UO_734 (O_734,N_4689,N_4041);
nor UO_735 (O_735,N_4248,N_4386);
and UO_736 (O_736,N_4640,N_4418);
nand UO_737 (O_737,N_4575,N_4700);
nor UO_738 (O_738,N_4632,N_4371);
and UO_739 (O_739,N_4206,N_4416);
nor UO_740 (O_740,N_4157,N_4879);
xor UO_741 (O_741,N_4190,N_4821);
nor UO_742 (O_742,N_4471,N_4727);
and UO_743 (O_743,N_4013,N_4987);
or UO_744 (O_744,N_4120,N_4582);
and UO_745 (O_745,N_4684,N_4079);
nand UO_746 (O_746,N_4132,N_4767);
or UO_747 (O_747,N_4353,N_4127);
or UO_748 (O_748,N_4156,N_4582);
and UO_749 (O_749,N_4058,N_4118);
and UO_750 (O_750,N_4415,N_4178);
nand UO_751 (O_751,N_4853,N_4395);
or UO_752 (O_752,N_4545,N_4242);
nor UO_753 (O_753,N_4199,N_4846);
nor UO_754 (O_754,N_4336,N_4997);
nand UO_755 (O_755,N_4963,N_4687);
nand UO_756 (O_756,N_4220,N_4065);
and UO_757 (O_757,N_4704,N_4767);
nor UO_758 (O_758,N_4815,N_4888);
nand UO_759 (O_759,N_4049,N_4982);
nor UO_760 (O_760,N_4770,N_4954);
nor UO_761 (O_761,N_4060,N_4651);
and UO_762 (O_762,N_4864,N_4423);
and UO_763 (O_763,N_4507,N_4611);
or UO_764 (O_764,N_4366,N_4179);
or UO_765 (O_765,N_4964,N_4401);
nand UO_766 (O_766,N_4501,N_4529);
nand UO_767 (O_767,N_4811,N_4278);
and UO_768 (O_768,N_4135,N_4286);
or UO_769 (O_769,N_4129,N_4226);
xnor UO_770 (O_770,N_4523,N_4768);
nor UO_771 (O_771,N_4169,N_4615);
and UO_772 (O_772,N_4853,N_4342);
nand UO_773 (O_773,N_4487,N_4609);
xor UO_774 (O_774,N_4116,N_4874);
or UO_775 (O_775,N_4831,N_4960);
xnor UO_776 (O_776,N_4964,N_4634);
xor UO_777 (O_777,N_4109,N_4864);
nand UO_778 (O_778,N_4217,N_4032);
xnor UO_779 (O_779,N_4325,N_4408);
nor UO_780 (O_780,N_4648,N_4491);
nand UO_781 (O_781,N_4564,N_4606);
nor UO_782 (O_782,N_4356,N_4828);
nand UO_783 (O_783,N_4668,N_4712);
and UO_784 (O_784,N_4903,N_4548);
and UO_785 (O_785,N_4982,N_4257);
or UO_786 (O_786,N_4542,N_4167);
nand UO_787 (O_787,N_4567,N_4617);
and UO_788 (O_788,N_4806,N_4503);
or UO_789 (O_789,N_4760,N_4979);
nor UO_790 (O_790,N_4496,N_4268);
and UO_791 (O_791,N_4513,N_4523);
xnor UO_792 (O_792,N_4753,N_4520);
or UO_793 (O_793,N_4711,N_4184);
or UO_794 (O_794,N_4508,N_4365);
nand UO_795 (O_795,N_4495,N_4767);
and UO_796 (O_796,N_4552,N_4686);
nand UO_797 (O_797,N_4191,N_4698);
and UO_798 (O_798,N_4851,N_4228);
and UO_799 (O_799,N_4016,N_4807);
nand UO_800 (O_800,N_4401,N_4768);
nor UO_801 (O_801,N_4093,N_4542);
xnor UO_802 (O_802,N_4034,N_4978);
nor UO_803 (O_803,N_4136,N_4554);
nor UO_804 (O_804,N_4483,N_4881);
nand UO_805 (O_805,N_4642,N_4834);
nand UO_806 (O_806,N_4161,N_4708);
and UO_807 (O_807,N_4440,N_4588);
nor UO_808 (O_808,N_4275,N_4852);
and UO_809 (O_809,N_4579,N_4989);
nand UO_810 (O_810,N_4134,N_4667);
or UO_811 (O_811,N_4837,N_4636);
xnor UO_812 (O_812,N_4688,N_4819);
nor UO_813 (O_813,N_4430,N_4327);
nand UO_814 (O_814,N_4034,N_4731);
nand UO_815 (O_815,N_4276,N_4483);
and UO_816 (O_816,N_4268,N_4324);
nand UO_817 (O_817,N_4792,N_4707);
nand UO_818 (O_818,N_4076,N_4148);
and UO_819 (O_819,N_4805,N_4138);
and UO_820 (O_820,N_4102,N_4009);
or UO_821 (O_821,N_4872,N_4252);
nor UO_822 (O_822,N_4095,N_4205);
nor UO_823 (O_823,N_4766,N_4528);
or UO_824 (O_824,N_4166,N_4496);
nand UO_825 (O_825,N_4517,N_4868);
nand UO_826 (O_826,N_4883,N_4511);
nand UO_827 (O_827,N_4163,N_4785);
nand UO_828 (O_828,N_4484,N_4581);
xor UO_829 (O_829,N_4585,N_4358);
or UO_830 (O_830,N_4837,N_4044);
and UO_831 (O_831,N_4444,N_4979);
nor UO_832 (O_832,N_4640,N_4649);
or UO_833 (O_833,N_4641,N_4043);
or UO_834 (O_834,N_4355,N_4016);
nand UO_835 (O_835,N_4948,N_4193);
nand UO_836 (O_836,N_4655,N_4677);
nor UO_837 (O_837,N_4360,N_4572);
nor UO_838 (O_838,N_4299,N_4352);
or UO_839 (O_839,N_4216,N_4929);
and UO_840 (O_840,N_4068,N_4279);
xnor UO_841 (O_841,N_4658,N_4960);
and UO_842 (O_842,N_4115,N_4834);
nor UO_843 (O_843,N_4296,N_4032);
nand UO_844 (O_844,N_4206,N_4476);
nand UO_845 (O_845,N_4146,N_4774);
and UO_846 (O_846,N_4353,N_4916);
and UO_847 (O_847,N_4730,N_4422);
or UO_848 (O_848,N_4580,N_4037);
and UO_849 (O_849,N_4517,N_4668);
or UO_850 (O_850,N_4196,N_4509);
nand UO_851 (O_851,N_4875,N_4196);
nand UO_852 (O_852,N_4816,N_4172);
nand UO_853 (O_853,N_4694,N_4666);
and UO_854 (O_854,N_4783,N_4499);
nor UO_855 (O_855,N_4113,N_4904);
or UO_856 (O_856,N_4571,N_4015);
nor UO_857 (O_857,N_4470,N_4592);
and UO_858 (O_858,N_4462,N_4228);
nor UO_859 (O_859,N_4841,N_4483);
and UO_860 (O_860,N_4169,N_4129);
or UO_861 (O_861,N_4117,N_4969);
or UO_862 (O_862,N_4585,N_4015);
and UO_863 (O_863,N_4447,N_4095);
nand UO_864 (O_864,N_4895,N_4097);
nand UO_865 (O_865,N_4595,N_4230);
nor UO_866 (O_866,N_4726,N_4511);
and UO_867 (O_867,N_4960,N_4917);
or UO_868 (O_868,N_4283,N_4477);
nand UO_869 (O_869,N_4800,N_4644);
or UO_870 (O_870,N_4882,N_4431);
or UO_871 (O_871,N_4037,N_4108);
or UO_872 (O_872,N_4465,N_4275);
and UO_873 (O_873,N_4245,N_4326);
nand UO_874 (O_874,N_4191,N_4514);
or UO_875 (O_875,N_4627,N_4660);
or UO_876 (O_876,N_4251,N_4000);
and UO_877 (O_877,N_4858,N_4033);
xnor UO_878 (O_878,N_4208,N_4589);
nor UO_879 (O_879,N_4564,N_4170);
nor UO_880 (O_880,N_4435,N_4655);
nor UO_881 (O_881,N_4190,N_4930);
and UO_882 (O_882,N_4969,N_4522);
or UO_883 (O_883,N_4796,N_4483);
or UO_884 (O_884,N_4543,N_4298);
nor UO_885 (O_885,N_4681,N_4853);
and UO_886 (O_886,N_4124,N_4765);
nand UO_887 (O_887,N_4700,N_4191);
and UO_888 (O_888,N_4763,N_4289);
nor UO_889 (O_889,N_4862,N_4441);
nand UO_890 (O_890,N_4760,N_4545);
nor UO_891 (O_891,N_4269,N_4354);
nand UO_892 (O_892,N_4362,N_4867);
nor UO_893 (O_893,N_4661,N_4354);
nor UO_894 (O_894,N_4714,N_4688);
nand UO_895 (O_895,N_4919,N_4441);
xor UO_896 (O_896,N_4032,N_4973);
and UO_897 (O_897,N_4925,N_4115);
nand UO_898 (O_898,N_4225,N_4760);
and UO_899 (O_899,N_4009,N_4353);
and UO_900 (O_900,N_4849,N_4903);
nand UO_901 (O_901,N_4346,N_4246);
nand UO_902 (O_902,N_4248,N_4935);
nor UO_903 (O_903,N_4562,N_4266);
nor UO_904 (O_904,N_4876,N_4526);
nor UO_905 (O_905,N_4385,N_4967);
and UO_906 (O_906,N_4884,N_4900);
nand UO_907 (O_907,N_4604,N_4749);
nand UO_908 (O_908,N_4209,N_4590);
and UO_909 (O_909,N_4958,N_4784);
nand UO_910 (O_910,N_4492,N_4224);
and UO_911 (O_911,N_4769,N_4370);
nand UO_912 (O_912,N_4377,N_4357);
and UO_913 (O_913,N_4439,N_4470);
nand UO_914 (O_914,N_4633,N_4861);
and UO_915 (O_915,N_4783,N_4151);
or UO_916 (O_916,N_4056,N_4415);
nand UO_917 (O_917,N_4596,N_4569);
and UO_918 (O_918,N_4073,N_4850);
nand UO_919 (O_919,N_4657,N_4102);
or UO_920 (O_920,N_4645,N_4391);
nor UO_921 (O_921,N_4407,N_4399);
xor UO_922 (O_922,N_4644,N_4625);
and UO_923 (O_923,N_4955,N_4011);
and UO_924 (O_924,N_4009,N_4879);
nor UO_925 (O_925,N_4653,N_4079);
nor UO_926 (O_926,N_4981,N_4929);
or UO_927 (O_927,N_4869,N_4491);
or UO_928 (O_928,N_4359,N_4877);
nand UO_929 (O_929,N_4870,N_4384);
nor UO_930 (O_930,N_4878,N_4817);
and UO_931 (O_931,N_4835,N_4364);
or UO_932 (O_932,N_4490,N_4503);
nor UO_933 (O_933,N_4881,N_4561);
nor UO_934 (O_934,N_4529,N_4738);
nor UO_935 (O_935,N_4785,N_4968);
nand UO_936 (O_936,N_4896,N_4963);
and UO_937 (O_937,N_4876,N_4762);
or UO_938 (O_938,N_4949,N_4618);
or UO_939 (O_939,N_4702,N_4334);
nand UO_940 (O_940,N_4112,N_4156);
or UO_941 (O_941,N_4306,N_4278);
or UO_942 (O_942,N_4850,N_4000);
or UO_943 (O_943,N_4749,N_4443);
and UO_944 (O_944,N_4928,N_4516);
and UO_945 (O_945,N_4386,N_4529);
nor UO_946 (O_946,N_4524,N_4495);
and UO_947 (O_947,N_4758,N_4211);
and UO_948 (O_948,N_4608,N_4254);
and UO_949 (O_949,N_4345,N_4352);
and UO_950 (O_950,N_4428,N_4369);
nand UO_951 (O_951,N_4352,N_4108);
and UO_952 (O_952,N_4080,N_4930);
or UO_953 (O_953,N_4236,N_4938);
nor UO_954 (O_954,N_4501,N_4208);
or UO_955 (O_955,N_4369,N_4351);
nand UO_956 (O_956,N_4592,N_4610);
nand UO_957 (O_957,N_4579,N_4460);
xnor UO_958 (O_958,N_4441,N_4818);
nor UO_959 (O_959,N_4649,N_4880);
and UO_960 (O_960,N_4487,N_4981);
and UO_961 (O_961,N_4492,N_4065);
and UO_962 (O_962,N_4667,N_4099);
and UO_963 (O_963,N_4059,N_4596);
and UO_964 (O_964,N_4534,N_4985);
or UO_965 (O_965,N_4879,N_4033);
nand UO_966 (O_966,N_4588,N_4999);
nand UO_967 (O_967,N_4023,N_4237);
nor UO_968 (O_968,N_4587,N_4044);
or UO_969 (O_969,N_4215,N_4325);
nand UO_970 (O_970,N_4247,N_4006);
or UO_971 (O_971,N_4195,N_4463);
nor UO_972 (O_972,N_4936,N_4933);
nand UO_973 (O_973,N_4765,N_4802);
and UO_974 (O_974,N_4284,N_4427);
nor UO_975 (O_975,N_4303,N_4230);
or UO_976 (O_976,N_4931,N_4763);
and UO_977 (O_977,N_4041,N_4728);
nand UO_978 (O_978,N_4106,N_4619);
or UO_979 (O_979,N_4489,N_4211);
nor UO_980 (O_980,N_4062,N_4421);
and UO_981 (O_981,N_4375,N_4175);
xor UO_982 (O_982,N_4851,N_4386);
xor UO_983 (O_983,N_4588,N_4997);
or UO_984 (O_984,N_4718,N_4866);
and UO_985 (O_985,N_4284,N_4800);
and UO_986 (O_986,N_4147,N_4939);
and UO_987 (O_987,N_4632,N_4279);
or UO_988 (O_988,N_4655,N_4883);
nand UO_989 (O_989,N_4539,N_4432);
nand UO_990 (O_990,N_4973,N_4048);
or UO_991 (O_991,N_4038,N_4175);
nand UO_992 (O_992,N_4001,N_4437);
nand UO_993 (O_993,N_4351,N_4498);
and UO_994 (O_994,N_4898,N_4769);
xnor UO_995 (O_995,N_4311,N_4147);
or UO_996 (O_996,N_4636,N_4127);
or UO_997 (O_997,N_4583,N_4307);
or UO_998 (O_998,N_4070,N_4012);
or UO_999 (O_999,N_4954,N_4913);
endmodule