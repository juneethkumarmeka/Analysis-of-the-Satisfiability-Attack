module basic_1500_15000_2000_5_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_401,In_854);
or U1 (N_1,In_1255,In_1261);
nor U2 (N_2,In_823,In_964);
nand U3 (N_3,In_1229,In_273);
nor U4 (N_4,In_10,In_951);
nand U5 (N_5,In_695,In_610);
nor U6 (N_6,In_1160,In_531);
nand U7 (N_7,In_1441,In_346);
nand U8 (N_8,In_563,In_659);
xor U9 (N_9,In_989,In_935);
nor U10 (N_10,In_1148,In_441);
and U11 (N_11,In_694,In_647);
and U12 (N_12,In_184,In_1082);
nand U13 (N_13,In_634,In_179);
and U14 (N_14,In_1205,In_163);
or U15 (N_15,In_551,In_491);
or U16 (N_16,In_1314,In_1245);
and U17 (N_17,In_1175,In_864);
nor U18 (N_18,In_845,In_1386);
or U19 (N_19,In_1480,In_1051);
or U20 (N_20,In_664,In_1005);
nor U21 (N_21,In_457,In_743);
nand U22 (N_22,In_379,In_192);
nor U23 (N_23,In_1010,In_1103);
nor U24 (N_24,In_389,In_586);
nand U25 (N_25,In_1418,In_1471);
nand U26 (N_26,In_1199,In_1495);
or U27 (N_27,In_1358,In_1341);
nand U28 (N_28,In_288,In_779);
or U29 (N_29,In_484,In_1004);
or U30 (N_30,In_1432,In_153);
nor U31 (N_31,In_166,In_337);
or U32 (N_32,In_640,In_1477);
xor U33 (N_33,In_573,In_482);
nand U34 (N_34,In_1047,In_617);
nor U35 (N_35,In_1489,In_203);
nor U36 (N_36,In_934,In_1074);
and U37 (N_37,In_592,In_17);
nand U38 (N_38,In_1254,In_1331);
nor U39 (N_39,In_519,In_1387);
nor U40 (N_40,In_675,In_858);
and U41 (N_41,In_649,In_644);
nand U42 (N_42,In_357,In_576);
nor U43 (N_43,In_927,In_15);
or U44 (N_44,In_663,In_528);
nand U45 (N_45,In_802,In_691);
nor U46 (N_46,In_585,In_1174);
and U47 (N_47,In_105,In_118);
nor U48 (N_48,In_134,In_777);
or U49 (N_49,In_997,In_186);
nand U50 (N_50,In_838,In_387);
or U51 (N_51,In_772,In_61);
and U52 (N_52,In_1252,In_1392);
or U53 (N_53,In_1034,In_570);
nor U54 (N_54,In_36,In_1421);
and U55 (N_55,In_1278,In_692);
or U56 (N_56,In_770,In_5);
nor U57 (N_57,In_1318,In_1285);
nor U58 (N_58,In_1135,In_417);
nand U59 (N_59,In_569,In_686);
and U60 (N_60,In_172,In_781);
nand U61 (N_61,In_521,In_1189);
nand U62 (N_62,In_653,In_413);
xor U63 (N_63,In_86,In_575);
and U64 (N_64,In_289,In_840);
nor U65 (N_65,In_810,In_1101);
nand U66 (N_66,In_1062,In_596);
nor U67 (N_67,In_1320,In_400);
or U68 (N_68,In_1420,In_1363);
nor U69 (N_69,In_1270,In_504);
nand U70 (N_70,In_44,In_236);
and U71 (N_71,In_104,In_442);
and U72 (N_72,In_499,In_247);
and U73 (N_73,In_1017,In_244);
or U74 (N_74,In_1227,In_9);
or U75 (N_75,In_533,In_587);
nand U76 (N_76,In_59,In_561);
nand U77 (N_77,In_322,In_656);
and U78 (N_78,In_875,In_385);
nand U79 (N_79,In_643,In_1413);
nor U80 (N_80,In_980,In_775);
nand U81 (N_81,In_77,In_588);
nand U82 (N_82,In_1059,In_751);
and U83 (N_83,In_809,In_125);
or U84 (N_84,In_886,In_96);
nand U85 (N_85,In_873,In_262);
nor U86 (N_86,In_308,In_1258);
and U87 (N_87,In_328,In_728);
nor U88 (N_88,In_992,In_43);
and U89 (N_89,In_880,In_1231);
xnor U90 (N_90,In_1066,In_1339);
nor U91 (N_91,In_568,In_48);
and U92 (N_92,In_269,In_277);
and U93 (N_93,In_591,In_967);
nor U94 (N_94,In_705,In_1086);
nor U95 (N_95,In_1228,In_267);
or U96 (N_96,In_386,In_45);
nor U97 (N_97,In_900,In_8);
and U98 (N_98,In_892,In_1294);
nor U99 (N_99,In_611,In_1403);
or U100 (N_100,In_536,In_366);
nor U101 (N_101,In_1451,In_853);
nor U102 (N_102,In_330,In_768);
nor U103 (N_103,In_1183,In_911);
nand U104 (N_104,In_919,In_1375);
nor U105 (N_105,In_776,In_1416);
nor U106 (N_106,In_537,In_693);
nor U107 (N_107,In_1207,In_928);
nand U108 (N_108,In_1394,In_317);
and U109 (N_109,In_508,In_762);
nor U110 (N_110,In_672,In_489);
nor U111 (N_111,In_954,In_1373);
nor U112 (N_112,In_807,In_766);
nand U113 (N_113,In_1242,In_1493);
and U114 (N_114,In_383,In_1498);
nor U115 (N_115,In_973,In_1043);
nand U116 (N_116,In_488,In_1406);
and U117 (N_117,In_517,In_32);
and U118 (N_118,In_174,In_314);
nor U119 (N_119,In_494,In_416);
and U120 (N_120,In_1049,In_365);
nand U121 (N_121,In_72,In_1192);
or U122 (N_122,In_1486,In_1391);
nor U123 (N_123,In_908,In_1385);
and U124 (N_124,In_1203,In_729);
nor U125 (N_125,In_1407,In_941);
xnor U126 (N_126,In_437,In_196);
nand U127 (N_127,In_1295,In_1152);
nor U128 (N_128,In_47,In_354);
nand U129 (N_129,In_189,In_683);
nand U130 (N_130,In_744,In_414);
nand U131 (N_131,In_1351,In_641);
and U132 (N_132,In_635,In_1388);
nand U133 (N_133,In_108,In_791);
nand U134 (N_134,In_783,In_456);
nor U135 (N_135,In_1447,In_520);
and U136 (N_136,In_627,In_1263);
nand U137 (N_137,In_996,In_1225);
or U138 (N_138,In_201,In_213);
and U139 (N_139,In_359,In_95);
or U140 (N_140,In_233,In_107);
nand U141 (N_141,In_657,In_897);
or U142 (N_142,In_771,In_861);
and U143 (N_143,In_191,In_1170);
and U144 (N_144,In_970,In_205);
nand U145 (N_145,In_297,In_1208);
and U146 (N_146,In_870,In_803);
and U147 (N_147,In_741,In_1052);
nand U148 (N_148,In_857,In_1326);
nor U149 (N_149,In_290,In_953);
nand U150 (N_150,In_30,In_968);
nor U151 (N_151,In_422,In_352);
nand U152 (N_152,In_122,In_439);
or U153 (N_153,In_320,In_90);
or U154 (N_154,In_1,In_206);
xnor U155 (N_155,In_376,In_1076);
or U156 (N_156,In_197,In_360);
nand U157 (N_157,In_390,In_1310);
nand U158 (N_158,In_1401,In_187);
nor U159 (N_159,In_374,In_1438);
and U160 (N_160,In_1464,In_1473);
and U161 (N_161,In_633,In_119);
and U162 (N_162,In_1313,In_620);
nor U163 (N_163,In_567,In_217);
or U164 (N_164,In_1130,In_79);
nand U165 (N_165,In_1277,In_1301);
or U166 (N_166,In_790,In_805);
or U167 (N_167,In_1281,In_235);
nor U168 (N_168,In_1377,In_1444);
nor U169 (N_169,In_1303,In_21);
nor U170 (N_170,In_181,In_27);
xor U171 (N_171,In_285,In_168);
or U172 (N_172,In_1134,In_1131);
and U173 (N_173,In_1382,In_1354);
nand U174 (N_174,In_625,In_532);
or U175 (N_175,In_1319,In_1172);
nand U176 (N_176,In_738,In_1380);
and U177 (N_177,In_1031,In_665);
nand U178 (N_178,In_527,In_1057);
nand U179 (N_179,In_176,In_1117);
or U180 (N_180,In_377,In_1023);
nand U181 (N_181,In_847,In_444);
or U182 (N_182,In_1223,In_1024);
nand U183 (N_183,In_68,In_923);
and U184 (N_184,In_883,In_1309);
and U185 (N_185,In_1342,In_507);
and U186 (N_186,In_19,In_654);
and U187 (N_187,In_605,In_291);
nand U188 (N_188,In_714,In_937);
xor U189 (N_189,In_995,In_792);
nand U190 (N_190,In_602,In_836);
nand U191 (N_191,In_324,In_849);
nor U192 (N_192,In_1122,In_1452);
nor U193 (N_193,In_81,In_501);
and U194 (N_194,In_500,In_740);
nand U195 (N_195,In_1497,In_326);
or U196 (N_196,In_1093,In_600);
nor U197 (N_197,In_966,In_1218);
or U198 (N_198,In_303,In_228);
or U199 (N_199,In_868,In_577);
and U200 (N_200,In_566,In_1132);
nand U201 (N_201,In_1012,In_1247);
nand U202 (N_202,In_938,In_851);
or U203 (N_203,In_804,In_188);
and U204 (N_204,In_433,In_550);
nor U205 (N_205,In_667,In_917);
nor U206 (N_206,In_1224,In_1325);
nand U207 (N_207,In_1197,In_340);
and U208 (N_208,In_475,In_425);
and U209 (N_209,In_645,In_986);
or U210 (N_210,In_1039,In_1081);
and U211 (N_211,In_755,In_394);
nor U212 (N_212,In_1143,In_699);
or U213 (N_213,In_929,In_582);
and U214 (N_214,In_406,In_100);
nand U215 (N_215,In_82,In_147);
nand U216 (N_216,In_372,In_1356);
nand U217 (N_217,In_231,In_1346);
or U218 (N_218,In_298,In_1013);
and U219 (N_219,In_974,In_204);
and U220 (N_220,In_1150,In_1063);
and U221 (N_221,In_432,In_60);
xor U222 (N_222,In_1204,In_1381);
nor U223 (N_223,In_1032,In_246);
or U224 (N_224,In_276,In_869);
or U225 (N_225,In_338,In_1352);
nor U226 (N_226,In_841,In_73);
or U227 (N_227,In_815,In_467);
or U228 (N_228,In_1332,In_256);
nand U229 (N_229,In_881,In_89);
nand U230 (N_230,In_944,In_129);
nand U231 (N_231,In_702,In_57);
and U232 (N_232,In_959,In_632);
or U233 (N_233,In_1417,In_801);
and U234 (N_234,In_396,In_302);
or U235 (N_235,In_343,In_1186);
and U236 (N_236,In_4,In_218);
and U237 (N_237,In_785,In_240);
nor U238 (N_238,In_157,In_274);
nand U239 (N_239,In_1129,In_170);
nor U240 (N_240,In_724,In_183);
and U241 (N_241,In_711,In_265);
nor U242 (N_242,In_1064,In_1304);
and U243 (N_243,In_637,In_50);
nand U244 (N_244,In_315,In_1410);
or U245 (N_245,In_239,In_286);
nor U246 (N_246,In_133,In_846);
nor U247 (N_247,In_872,In_1119);
nand U248 (N_248,In_306,In_393);
nand U249 (N_249,In_882,In_219);
or U250 (N_250,In_392,In_1379);
nand U251 (N_251,In_1250,In_1350);
and U252 (N_252,In_1334,In_34);
xnor U253 (N_253,In_327,In_301);
or U254 (N_254,In_956,In_144);
or U255 (N_255,In_1488,In_215);
nand U256 (N_256,In_1465,In_292);
nor U257 (N_257,In_1126,In_375);
nand U258 (N_258,In_926,In_347);
nand U259 (N_259,In_930,In_1196);
and U260 (N_260,In_1458,In_737);
and U261 (N_261,In_173,In_1287);
nand U262 (N_262,In_1469,In_1167);
nor U263 (N_263,In_1234,In_713);
nand U264 (N_264,In_1427,In_75);
or U265 (N_265,In_543,In_0);
and U266 (N_266,In_1436,In_651);
or U267 (N_267,In_689,In_227);
and U268 (N_268,In_150,In_1091);
nand U269 (N_269,In_595,In_789);
and U270 (N_270,In_545,In_947);
and U271 (N_271,In_1376,In_242);
and U272 (N_272,In_557,In_1163);
or U273 (N_273,In_492,In_1496);
and U274 (N_274,In_171,In_1299);
or U275 (N_275,In_1290,In_1366);
nor U276 (N_276,In_866,In_760);
and U277 (N_277,In_1022,In_1009);
nand U278 (N_278,In_1405,In_420);
or U279 (N_279,In_808,In_162);
xor U280 (N_280,In_80,In_158);
nor U281 (N_281,In_1328,In_37);
and U282 (N_282,In_1165,In_1302);
nor U283 (N_283,In_590,In_412);
and U284 (N_284,In_373,In_248);
xor U285 (N_285,In_842,In_1279);
or U286 (N_286,In_932,In_316);
nand U287 (N_287,In_283,In_712);
or U288 (N_288,In_598,In_1070);
nor U289 (N_289,In_421,In_1397);
nand U290 (N_290,In_1219,In_294);
xnor U291 (N_291,In_754,In_831);
xnor U292 (N_292,In_1158,In_31);
nand U293 (N_293,In_24,In_341);
and U294 (N_294,In_812,In_109);
xor U295 (N_295,In_1355,In_548);
xnor U296 (N_296,In_87,In_707);
or U297 (N_297,In_1045,In_39);
and U298 (N_298,In_668,In_1274);
nor U299 (N_299,In_1275,In_382);
or U300 (N_300,In_1124,In_924);
xor U301 (N_301,In_1054,In_731);
nor U302 (N_302,In_1232,In_621);
and U303 (N_303,In_395,In_669);
or U304 (N_304,In_296,In_1353);
nor U305 (N_305,In_111,In_350);
or U306 (N_306,In_516,In_304);
nand U307 (N_307,In_369,In_185);
nand U308 (N_308,In_180,In_493);
or U309 (N_309,In_1000,In_1137);
nand U310 (N_310,In_1036,In_701);
nand U311 (N_311,In_684,In_722);
nor U312 (N_312,In_1109,In_1359);
and U313 (N_313,In_121,In_349);
nor U314 (N_314,In_1075,In_402);
or U315 (N_315,In_1187,In_1067);
nor U316 (N_316,In_553,In_293);
nor U317 (N_317,In_850,In_1142);
nor U318 (N_318,In_468,In_1466);
nand U319 (N_319,In_795,In_601);
nor U320 (N_320,In_912,In_1144);
nand U321 (N_321,In_942,In_814);
nand U322 (N_322,In_1335,In_112);
or U323 (N_323,In_901,In_1033);
nand U324 (N_324,In_364,In_1195);
and U325 (N_325,In_1105,In_540);
or U326 (N_326,In_680,In_752);
or U327 (N_327,In_1425,In_1282);
or U328 (N_328,In_142,In_312);
or U329 (N_329,In_280,In_604);
or U330 (N_330,In_1389,In_1206);
nand U331 (N_331,In_11,In_1409);
or U332 (N_332,In_631,In_1111);
and U333 (N_333,In_1316,In_1372);
nor U334 (N_334,In_140,In_859);
nand U335 (N_335,In_918,In_979);
and U336 (N_336,In_607,In_1190);
nor U337 (N_337,In_1378,In_1085);
nor U338 (N_338,In_638,In_888);
or U339 (N_339,In_156,In_1198);
or U340 (N_340,In_313,In_137);
or U341 (N_341,In_909,In_1293);
nor U342 (N_342,In_1404,In_555);
or U343 (N_343,In_1073,In_593);
or U344 (N_344,In_198,In_1222);
or U345 (N_345,In_697,In_1237);
and U346 (N_346,In_1096,In_608);
nor U347 (N_347,In_817,In_1337);
or U348 (N_348,In_409,In_1315);
xnor U349 (N_349,In_703,In_523);
nand U350 (N_350,In_93,In_753);
and U351 (N_351,In_1030,In_1433);
nand U352 (N_352,In_844,In_397);
nand U353 (N_353,In_455,In_819);
and U354 (N_354,In_138,In_902);
or U355 (N_355,In_794,In_117);
nor U356 (N_356,In_787,In_1181);
nand U357 (N_357,In_348,In_258);
or U358 (N_358,In_56,In_54);
or U359 (N_359,In_483,In_1138);
nor U360 (N_360,In_939,In_1272);
nand U361 (N_361,In_1114,In_1180);
nor U362 (N_362,In_1151,In_678);
nor U363 (N_363,In_1323,In_83);
nor U364 (N_364,In_299,In_175);
nor U365 (N_365,In_130,In_534);
or U366 (N_366,In_445,In_435);
or U367 (N_367,In_1016,In_271);
or U368 (N_368,In_18,In_52);
or U369 (N_369,In_148,In_1360);
or U370 (N_370,In_1347,In_813);
or U371 (N_371,In_1253,In_55);
nand U372 (N_372,In_384,In_1089);
or U373 (N_373,In_746,In_613);
and U374 (N_374,In_1308,In_497);
nand U375 (N_375,In_358,In_355);
or U376 (N_376,In_42,In_35);
nand U377 (N_377,In_700,In_629);
and U378 (N_378,In_730,In_458);
nand U379 (N_379,In_1448,In_473);
nand U380 (N_380,In_6,In_899);
or U381 (N_381,In_898,In_132);
nor U382 (N_382,In_983,In_1133);
nor U383 (N_383,In_773,In_1149);
nor U384 (N_384,In_1393,In_676);
or U385 (N_385,In_1455,In_910);
or U386 (N_386,In_487,In_1490);
nor U387 (N_387,In_1145,In_933);
and U388 (N_388,In_750,In_202);
xnor U389 (N_389,In_245,In_490);
nand U390 (N_390,In_987,In_1044);
or U391 (N_391,In_1435,In_839);
nand U392 (N_392,In_380,In_399);
or U393 (N_393,In_65,In_20);
nor U394 (N_394,In_1140,In_1021);
or U395 (N_395,In_459,In_110);
nor U396 (N_396,In_1078,In_98);
nand U397 (N_397,In_440,In_169);
and U398 (N_398,In_426,In_542);
nand U399 (N_399,In_530,In_234);
nand U400 (N_400,In_1291,In_509);
xor U401 (N_401,In_1364,In_541);
nor U402 (N_402,In_1399,In_99);
or U403 (N_403,In_200,In_463);
nand U404 (N_404,In_12,In_67);
nor U405 (N_405,In_250,In_1159);
or U406 (N_406,In_834,In_1235);
or U407 (N_407,In_1450,In_1256);
and U408 (N_408,In_415,In_211);
and U409 (N_409,In_131,In_742);
or U410 (N_410,In_615,In_1209);
or U411 (N_411,In_411,In_720);
nand U412 (N_412,In_614,In_1147);
nand U413 (N_413,In_1305,In_757);
and U414 (N_414,In_261,In_1079);
nand U415 (N_415,In_786,In_749);
and U416 (N_416,In_1408,In_1214);
nor U417 (N_417,In_856,In_1061);
nand U418 (N_418,In_154,In_626);
or U419 (N_419,In_1348,In_477);
nand U420 (N_420,In_670,In_225);
nor U421 (N_421,In_1156,In_325);
nor U422 (N_422,In_706,In_74);
nor U423 (N_423,In_1440,In_165);
and U424 (N_424,In_1007,In_423);
nand U425 (N_425,In_1479,In_1468);
nor U426 (N_426,In_70,In_718);
nor U427 (N_427,In_1369,In_1179);
nor U428 (N_428,In_388,In_1296);
nand U429 (N_429,In_113,In_761);
and U430 (N_430,In_1475,In_1443);
xnor U431 (N_431,In_472,In_64);
nor U432 (N_432,In_774,In_13);
and U433 (N_433,In_1090,In_1188);
or U434 (N_434,In_3,In_616);
and U435 (N_435,In_102,In_565);
and U436 (N_436,In_1400,In_1260);
and U437 (N_437,In_685,In_332);
nand U438 (N_438,In_319,In_920);
or U439 (N_439,In_758,In_1095);
or U440 (N_440,In_619,In_403);
and U441 (N_441,In_91,In_1402);
nand U442 (N_442,In_1098,In_1414);
nor U443 (N_443,In_921,In_123);
and U444 (N_444,In_1239,In_1236);
or U445 (N_445,In_1484,In_465);
and U446 (N_446,In_1155,In_195);
nand U447 (N_447,In_903,In_1437);
nor U448 (N_448,In_427,In_287);
and U449 (N_449,In_251,In_958);
xor U450 (N_450,In_1002,In_811);
nand U451 (N_451,In_1454,In_1202);
nand U452 (N_452,In_571,In_1268);
nor U453 (N_453,In_253,In_574);
or U454 (N_454,In_1003,In_1077);
or U455 (N_455,In_345,In_960);
nor U456 (N_456,In_606,In_1494);
nand U457 (N_457,In_1390,In_1211);
nor U458 (N_458,In_915,In_1434);
and U459 (N_459,In_1461,In_1271);
and U460 (N_460,In_429,In_609);
or U461 (N_461,In_982,In_716);
and U462 (N_462,In_1446,In_1177);
and U463 (N_463,In_579,In_1395);
or U464 (N_464,In_554,In_85);
or U465 (N_465,In_241,In_1422);
nand U466 (N_466,In_896,In_450);
nor U467 (N_467,In_835,In_279);
nor U468 (N_468,In_522,In_1104);
or U469 (N_469,In_126,In_904);
nor U470 (N_470,In_1029,In_594);
or U471 (N_471,In_1345,In_511);
and U472 (N_472,In_1123,In_476);
and U473 (N_473,In_1362,In_661);
or U474 (N_474,In_1384,In_763);
or U475 (N_475,In_430,In_232);
or U476 (N_476,In_1474,In_275);
nor U477 (N_477,In_985,In_735);
nor U478 (N_478,In_905,In_136);
and U479 (N_479,In_146,In_1298);
or U480 (N_480,In_1141,In_650);
nand U481 (N_481,In_949,In_1194);
nor U482 (N_482,In_1419,In_1108);
or U483 (N_483,In_1248,In_318);
or U484 (N_484,In_481,In_1191);
and U485 (N_485,In_470,In_103);
nor U486 (N_486,In_282,In_270);
nand U487 (N_487,In_1262,In_529);
or U488 (N_488,In_822,In_922);
nor U489 (N_489,In_539,In_837);
nor U490 (N_490,In_69,In_224);
nand U491 (N_491,In_141,In_263);
nor U492 (N_492,In_658,In_978);
nand U493 (N_493,In_549,In_145);
or U494 (N_494,In_1481,In_370);
and U495 (N_495,In_1240,In_1128);
nand U496 (N_496,In_436,In_405);
and U497 (N_497,In_1284,In_793);
nand U498 (N_498,In_538,In_988);
xnor U499 (N_499,In_1307,In_193);
nor U500 (N_500,In_1026,In_581);
nand U501 (N_501,In_1338,In_14);
nor U502 (N_502,In_748,In_1491);
or U503 (N_503,In_268,In_1019);
nor U504 (N_504,In_1040,In_1110);
nor U505 (N_505,In_698,In_1439);
or U506 (N_506,In_462,In_1321);
nand U507 (N_507,In_344,In_562);
nand U508 (N_508,In_310,In_1058);
nor U509 (N_509,In_723,In_739);
or U510 (N_510,In_747,In_704);
or U511 (N_511,In_128,In_818);
or U512 (N_512,In_1415,In_1324);
and U513 (N_513,In_945,In_1115);
nand U514 (N_514,In_1042,In_871);
or U515 (N_515,In_480,In_1327);
or U516 (N_516,In_971,In_478);
or U517 (N_517,In_552,In_278);
or U518 (N_518,In_92,In_952);
nand U519 (N_519,In_190,In_116);
nor U520 (N_520,In_252,In_560);
nand U521 (N_521,In_623,In_696);
nor U522 (N_522,In_865,In_950);
nor U523 (N_523,In_510,In_1371);
nor U524 (N_524,In_1210,In_1084);
or U525 (N_525,In_1423,In_199);
and U526 (N_526,In_767,In_525);
nor U527 (N_527,In_438,In_1312);
nor U528 (N_528,In_732,In_769);
or U529 (N_529,In_1244,In_1046);
and U530 (N_530,In_1241,In_564);
nand U531 (N_531,In_1453,In_874);
nor U532 (N_532,In_194,In_449);
nand U533 (N_533,In_1015,In_361);
and U534 (N_534,In_305,In_367);
and U535 (N_535,In_662,In_1367);
nand U536 (N_536,In_404,In_784);
nand U537 (N_537,In_782,In_1449);
nand U538 (N_538,In_597,In_1457);
nor U539 (N_539,In_1038,In_71);
nand U540 (N_540,In_1472,In_257);
nand U541 (N_541,In_1092,In_471);
and U542 (N_542,In_1154,In_1340);
nor U543 (N_543,In_284,In_41);
nand U544 (N_544,In_214,In_599);
nand U545 (N_545,In_1283,In_1168);
nor U546 (N_546,In_321,In_957);
and U547 (N_547,In_419,In_852);
and U548 (N_548,In_646,In_78);
and U549 (N_549,In_991,In_106);
and U550 (N_550,In_486,In_1035);
nand U551 (N_551,In_84,In_725);
or U552 (N_552,In_727,In_862);
nand U553 (N_553,In_222,In_1317);
and U554 (N_554,In_1127,In_832);
nor U555 (N_555,In_688,In_977);
or U556 (N_556,In_124,In_120);
nor U557 (N_557,In_40,In_879);
and U558 (N_558,In_1336,In_1171);
or U559 (N_559,In_914,In_311);
or U560 (N_560,In_1161,In_572);
nor U561 (N_561,In_88,In_1146);
nor U562 (N_562,In_1273,In_464);
nand U563 (N_563,In_1153,In_1330);
and U564 (N_564,In_167,In_636);
nand U565 (N_565,In_940,In_1184);
or U566 (N_566,In_816,In_1056);
xnor U567 (N_567,In_894,In_446);
nor U568 (N_568,In_1221,In_1333);
and U569 (N_569,In_558,In_351);
nor U570 (N_570,In_1467,In_1001);
or U571 (N_571,In_479,In_407);
nor U572 (N_572,In_877,In_1396);
or U573 (N_573,In_1349,In_580);
nand U574 (N_574,In_963,In_855);
nor U575 (N_575,In_356,In_381);
and U576 (N_576,In_1257,In_1106);
nor U577 (N_577,In_825,In_101);
or U578 (N_578,In_466,In_1025);
nor U579 (N_579,In_447,In_876);
or U580 (N_580,In_495,In_962);
nor U581 (N_581,In_1456,In_916);
and U582 (N_582,In_1169,In_1011);
nor U583 (N_583,In_1487,In_1118);
nand U584 (N_584,In_906,In_1083);
nor U585 (N_585,In_1322,In_1125);
nand U586 (N_586,In_502,In_1162);
and U587 (N_587,In_1292,In_1459);
nand U588 (N_588,In_1041,In_434);
nand U589 (N_589,In_1424,In_1311);
nand U590 (N_590,In_1139,In_719);
or U591 (N_591,In_512,In_671);
nor U592 (N_592,In_143,In_734);
nand U593 (N_593,In_38,In_1099);
and U594 (N_594,In_893,In_1398);
or U595 (N_595,In_677,In_221);
nand U596 (N_596,In_160,In_965);
nand U597 (N_597,In_254,In_1200);
or U598 (N_598,In_589,In_708);
nor U599 (N_599,In_682,In_1088);
nor U600 (N_600,In_135,In_765);
and U601 (N_601,In_556,In_513);
and U602 (N_602,In_1220,In_583);
and U603 (N_603,In_612,In_797);
or U604 (N_604,In_1037,In_1176);
and U605 (N_605,In_1344,In_339);
nor U606 (N_606,In_152,In_1266);
or U607 (N_607,In_334,In_1499);
nor U608 (N_608,In_300,In_485);
nor U609 (N_609,In_584,In_806);
or U610 (N_610,In_544,In_955);
nand U611 (N_611,In_1178,In_46);
nor U612 (N_612,In_925,In_884);
or U613 (N_613,In_26,In_1068);
nor U614 (N_614,In_207,In_715);
or U615 (N_615,In_526,In_1121);
nor U616 (N_616,In_1112,In_690);
or U617 (N_617,In_1276,In_76);
nand U618 (N_618,In_159,In_51);
or U619 (N_619,In_535,In_1264);
nor U620 (N_620,In_281,In_547);
and U621 (N_621,In_1173,In_642);
nor U622 (N_622,In_460,In_418);
nand U623 (N_623,In_498,In_887);
or U624 (N_624,In_624,In_948);
or U625 (N_625,In_1470,In_1286);
and U626 (N_626,In_1217,In_1482);
nor U627 (N_627,In_260,In_1216);
nand U628 (N_628,In_333,In_890);
or U629 (N_629,In_295,In_114);
nand U630 (N_630,In_378,In_209);
and U631 (N_631,In_16,In_1476);
xor U632 (N_632,In_1343,In_1297);
nand U633 (N_633,In_1411,In_503);
or U634 (N_634,In_1102,In_1157);
nor U635 (N_635,In_681,In_1050);
or U636 (N_636,In_1071,In_94);
nor U637 (N_637,In_1368,In_1463);
or U638 (N_638,In_151,In_266);
nor U639 (N_639,In_721,In_223);
or U640 (N_640,In_1259,In_1060);
nand U641 (N_641,In_264,In_559);
nor U642 (N_642,In_878,In_474);
nand U643 (N_643,In_1269,In_335);
nor U644 (N_644,In_630,In_885);
nor U645 (N_645,In_639,In_216);
and U646 (N_646,In_1215,In_1249);
nor U647 (N_647,In_820,In_1370);
nor U648 (N_648,In_1120,In_946);
nand U649 (N_649,In_1430,In_149);
and U650 (N_650,In_28,In_424);
or U651 (N_651,In_687,In_1097);
and U652 (N_652,In_603,In_943);
nand U653 (N_653,In_1300,In_453);
and U654 (N_654,In_759,In_1226);
nand U655 (N_655,In_398,In_981);
nand U656 (N_656,In_1055,In_1442);
nand U657 (N_657,In_798,In_1374);
xnor U658 (N_658,In_628,In_238);
or U659 (N_659,In_1027,In_1014);
and U660 (N_660,In_726,In_1028);
or U661 (N_661,In_679,In_1265);
nor U662 (N_662,In_1329,In_1238);
nor U663 (N_663,In_307,In_824);
or U664 (N_664,In_1020,In_1065);
nor U665 (N_665,In_23,In_829);
and U666 (N_666,In_984,In_1087);
nor U667 (N_667,In_961,In_309);
and U668 (N_668,In_1429,In_655);
nor U669 (N_669,In_1018,In_226);
nand U670 (N_670,In_342,In_237);
or U671 (N_671,In_1460,In_229);
xnor U672 (N_672,In_709,In_329);
nand U673 (N_673,In_1478,In_975);
nand U674 (N_674,In_155,In_863);
nor U675 (N_675,In_249,In_127);
nand U676 (N_676,In_212,In_431);
nand U677 (N_677,In_1048,In_518);
nor U678 (N_678,In_999,In_1483);
nand U679 (N_679,In_7,In_660);
nand U680 (N_680,In_49,In_323);
and U681 (N_681,In_1069,In_506);
and U682 (N_682,In_177,In_1246);
or U683 (N_683,In_1185,In_391);
nor U684 (N_684,In_272,In_448);
and U685 (N_685,In_1462,In_827);
and U686 (N_686,In_733,In_461);
nor U687 (N_687,In_972,In_29);
nand U688 (N_688,In_58,In_1383);
and U689 (N_689,In_336,In_1251);
or U690 (N_690,In_1212,In_764);
or U691 (N_691,In_259,In_710);
nor U692 (N_692,In_826,In_208);
or U693 (N_693,In_408,In_799);
nand U694 (N_694,In_578,In_780);
xnor U695 (N_695,In_524,In_994);
nor U696 (N_696,In_454,In_452);
nand U697 (N_697,In_1233,In_1113);
nand U698 (N_698,In_833,In_889);
or U699 (N_699,In_2,In_652);
and U700 (N_700,In_410,In_788);
and U701 (N_701,In_66,In_1193);
nand U702 (N_702,In_496,In_990);
and U703 (N_703,In_778,In_164);
nand U704 (N_704,In_25,In_230);
nor U705 (N_705,In_1201,In_220);
or U706 (N_706,In_843,In_891);
and U707 (N_707,In_931,In_62);
and U708 (N_708,In_1492,In_830);
xor U709 (N_709,In_182,In_210);
nand U710 (N_710,In_1230,In_895);
or U711 (N_711,In_505,In_161);
nor U712 (N_712,In_1431,In_821);
and U713 (N_713,In_736,In_848);
and U714 (N_714,In_515,In_622);
or U715 (N_715,In_469,In_115);
and U716 (N_716,In_756,In_1072);
xnor U717 (N_717,In_717,In_800);
and U718 (N_718,In_428,In_1008);
and U719 (N_719,In_936,In_1094);
and U720 (N_720,In_243,In_867);
xnor U721 (N_721,In_546,In_443);
and U722 (N_722,In_1306,In_1080);
nand U723 (N_723,In_1365,In_1280);
nor U724 (N_724,In_828,In_1166);
or U725 (N_725,In_1428,In_255);
or U726 (N_726,In_33,In_1485);
and U727 (N_727,In_1426,In_1288);
or U728 (N_728,In_363,In_648);
nor U729 (N_729,In_1164,In_353);
nor U730 (N_730,In_993,In_998);
nand U731 (N_731,In_63,In_1182);
nand U732 (N_732,In_514,In_860);
and U733 (N_733,In_1361,In_1100);
nor U734 (N_734,In_371,In_1053);
and U735 (N_735,In_451,In_1136);
or U736 (N_736,In_1267,In_97);
or U737 (N_737,In_1243,In_1213);
or U738 (N_738,In_796,In_1116);
nor U739 (N_739,In_976,In_745);
or U740 (N_740,In_362,In_139);
nand U741 (N_741,In_969,In_618);
nor U742 (N_742,In_674,In_1357);
or U743 (N_743,In_1006,In_178);
nor U744 (N_744,In_53,In_907);
or U745 (N_745,In_331,In_1107);
nor U746 (N_746,In_913,In_666);
nor U747 (N_747,In_22,In_673);
nor U748 (N_748,In_1412,In_1445);
nand U749 (N_749,In_1289,In_368);
nand U750 (N_750,In_524,In_153);
and U751 (N_751,In_226,In_829);
or U752 (N_752,In_227,In_192);
and U753 (N_753,In_561,In_1091);
nand U754 (N_754,In_167,In_1481);
and U755 (N_755,In_548,In_501);
and U756 (N_756,In_161,In_1173);
and U757 (N_757,In_1100,In_593);
and U758 (N_758,In_312,In_458);
or U759 (N_759,In_894,In_1322);
or U760 (N_760,In_860,In_897);
nor U761 (N_761,In_1012,In_1489);
or U762 (N_762,In_140,In_1263);
nor U763 (N_763,In_37,In_1352);
nand U764 (N_764,In_1326,In_669);
nand U765 (N_765,In_628,In_643);
nor U766 (N_766,In_1482,In_1137);
or U767 (N_767,In_500,In_1040);
nor U768 (N_768,In_42,In_237);
nor U769 (N_769,In_789,In_652);
or U770 (N_770,In_178,In_787);
nand U771 (N_771,In_74,In_1197);
nor U772 (N_772,In_1052,In_928);
or U773 (N_773,In_93,In_491);
and U774 (N_774,In_1195,In_1206);
or U775 (N_775,In_1490,In_450);
nand U776 (N_776,In_212,In_1303);
nand U777 (N_777,In_53,In_1489);
or U778 (N_778,In_468,In_1086);
and U779 (N_779,In_1155,In_974);
or U780 (N_780,In_1324,In_1470);
nand U781 (N_781,In_1183,In_1482);
nor U782 (N_782,In_1091,In_1349);
and U783 (N_783,In_1178,In_865);
nor U784 (N_784,In_109,In_437);
and U785 (N_785,In_1287,In_1435);
nand U786 (N_786,In_226,In_1263);
or U787 (N_787,In_1336,In_1229);
nor U788 (N_788,In_458,In_1014);
nor U789 (N_789,In_93,In_1463);
nand U790 (N_790,In_119,In_851);
or U791 (N_791,In_570,In_394);
or U792 (N_792,In_818,In_1342);
and U793 (N_793,In_1224,In_177);
nor U794 (N_794,In_116,In_416);
nor U795 (N_795,In_1141,In_523);
nand U796 (N_796,In_1321,In_1238);
and U797 (N_797,In_834,In_792);
nand U798 (N_798,In_518,In_115);
xor U799 (N_799,In_1190,In_922);
nand U800 (N_800,In_1221,In_506);
nor U801 (N_801,In_1234,In_111);
nor U802 (N_802,In_1187,In_1155);
nor U803 (N_803,In_386,In_52);
and U804 (N_804,In_204,In_1326);
or U805 (N_805,In_131,In_1287);
or U806 (N_806,In_732,In_371);
and U807 (N_807,In_1436,In_400);
nand U808 (N_808,In_818,In_1018);
nand U809 (N_809,In_1006,In_1444);
or U810 (N_810,In_146,In_1249);
or U811 (N_811,In_621,In_1339);
nor U812 (N_812,In_370,In_232);
nor U813 (N_813,In_460,In_824);
or U814 (N_814,In_1292,In_524);
and U815 (N_815,In_105,In_35);
nor U816 (N_816,In_27,In_800);
nand U817 (N_817,In_744,In_1038);
nor U818 (N_818,In_1323,In_921);
nor U819 (N_819,In_1087,In_1322);
nor U820 (N_820,In_1347,In_1154);
nor U821 (N_821,In_1440,In_86);
and U822 (N_822,In_690,In_20);
nor U823 (N_823,In_293,In_1174);
nor U824 (N_824,In_512,In_928);
nor U825 (N_825,In_1158,In_826);
and U826 (N_826,In_686,In_1198);
or U827 (N_827,In_412,In_333);
nand U828 (N_828,In_391,In_22);
or U829 (N_829,In_310,In_879);
xor U830 (N_830,In_785,In_1353);
nor U831 (N_831,In_215,In_95);
or U832 (N_832,In_1289,In_1413);
and U833 (N_833,In_599,In_719);
or U834 (N_834,In_576,In_139);
and U835 (N_835,In_326,In_155);
nor U836 (N_836,In_1395,In_174);
nor U837 (N_837,In_920,In_1489);
or U838 (N_838,In_752,In_1404);
and U839 (N_839,In_703,In_495);
or U840 (N_840,In_467,In_685);
nand U841 (N_841,In_515,In_1393);
nand U842 (N_842,In_1264,In_792);
nand U843 (N_843,In_450,In_1071);
nor U844 (N_844,In_360,In_1234);
or U845 (N_845,In_749,In_673);
and U846 (N_846,In_453,In_1207);
nor U847 (N_847,In_359,In_884);
or U848 (N_848,In_561,In_1457);
and U849 (N_849,In_273,In_1027);
and U850 (N_850,In_1211,In_110);
and U851 (N_851,In_528,In_503);
and U852 (N_852,In_1180,In_1308);
and U853 (N_853,In_977,In_1260);
or U854 (N_854,In_335,In_142);
nor U855 (N_855,In_1410,In_1455);
nor U856 (N_856,In_1344,In_162);
nor U857 (N_857,In_1296,In_297);
nor U858 (N_858,In_729,In_939);
nand U859 (N_859,In_757,In_171);
nor U860 (N_860,In_187,In_242);
nand U861 (N_861,In_1332,In_809);
nor U862 (N_862,In_924,In_314);
or U863 (N_863,In_688,In_96);
and U864 (N_864,In_263,In_280);
and U865 (N_865,In_1488,In_419);
nand U866 (N_866,In_374,In_1288);
nor U867 (N_867,In_902,In_813);
nand U868 (N_868,In_734,In_1233);
or U869 (N_869,In_342,In_87);
or U870 (N_870,In_1220,In_250);
nor U871 (N_871,In_1170,In_447);
nor U872 (N_872,In_775,In_100);
or U873 (N_873,In_108,In_1109);
and U874 (N_874,In_900,In_269);
or U875 (N_875,In_1439,In_904);
xor U876 (N_876,In_968,In_403);
and U877 (N_877,In_802,In_1450);
or U878 (N_878,In_1112,In_811);
nand U879 (N_879,In_1326,In_216);
and U880 (N_880,In_1176,In_154);
nand U881 (N_881,In_468,In_594);
and U882 (N_882,In_771,In_208);
nor U883 (N_883,In_236,In_289);
or U884 (N_884,In_795,In_910);
nor U885 (N_885,In_1399,In_149);
nand U886 (N_886,In_796,In_1079);
or U887 (N_887,In_1152,In_29);
and U888 (N_888,In_198,In_381);
nor U889 (N_889,In_1356,In_523);
nand U890 (N_890,In_1063,In_270);
and U891 (N_891,In_950,In_648);
and U892 (N_892,In_1195,In_375);
nor U893 (N_893,In_1297,In_496);
and U894 (N_894,In_200,In_659);
nor U895 (N_895,In_664,In_1433);
nand U896 (N_896,In_644,In_888);
nand U897 (N_897,In_266,In_880);
or U898 (N_898,In_304,In_932);
nand U899 (N_899,In_434,In_530);
or U900 (N_900,In_14,In_887);
or U901 (N_901,In_1446,In_731);
nor U902 (N_902,In_827,In_990);
nand U903 (N_903,In_67,In_800);
xnor U904 (N_904,In_949,In_26);
and U905 (N_905,In_830,In_1252);
nor U906 (N_906,In_1011,In_748);
nand U907 (N_907,In_175,In_118);
or U908 (N_908,In_224,In_1146);
or U909 (N_909,In_9,In_1367);
or U910 (N_910,In_185,In_706);
nand U911 (N_911,In_329,In_292);
nand U912 (N_912,In_711,In_679);
or U913 (N_913,In_705,In_837);
or U914 (N_914,In_20,In_1215);
nand U915 (N_915,In_363,In_252);
and U916 (N_916,In_863,In_139);
or U917 (N_917,In_1250,In_0);
nor U918 (N_918,In_132,In_1301);
nor U919 (N_919,In_83,In_1364);
nor U920 (N_920,In_1093,In_1079);
nor U921 (N_921,In_40,In_28);
and U922 (N_922,In_349,In_504);
nor U923 (N_923,In_104,In_397);
or U924 (N_924,In_1372,In_611);
nor U925 (N_925,In_10,In_581);
nor U926 (N_926,In_1017,In_8);
nor U927 (N_927,In_21,In_310);
nor U928 (N_928,In_36,In_205);
or U929 (N_929,In_395,In_1064);
or U930 (N_930,In_1096,In_770);
nand U931 (N_931,In_1476,In_102);
nor U932 (N_932,In_936,In_424);
and U933 (N_933,In_738,In_537);
nor U934 (N_934,In_458,In_1383);
and U935 (N_935,In_975,In_1281);
nor U936 (N_936,In_882,In_1315);
nor U937 (N_937,In_1199,In_1095);
nor U938 (N_938,In_1018,In_526);
nand U939 (N_939,In_521,In_577);
nor U940 (N_940,In_591,In_722);
and U941 (N_941,In_432,In_1270);
nor U942 (N_942,In_68,In_1285);
and U943 (N_943,In_822,In_1383);
and U944 (N_944,In_418,In_1493);
and U945 (N_945,In_599,In_1473);
nor U946 (N_946,In_390,In_243);
nand U947 (N_947,In_984,In_1129);
xnor U948 (N_948,In_1226,In_1492);
and U949 (N_949,In_449,In_679);
nand U950 (N_950,In_972,In_745);
xnor U951 (N_951,In_530,In_1218);
nor U952 (N_952,In_400,In_1497);
nand U953 (N_953,In_747,In_33);
or U954 (N_954,In_33,In_182);
and U955 (N_955,In_817,In_306);
or U956 (N_956,In_836,In_1239);
nand U957 (N_957,In_692,In_26);
and U958 (N_958,In_375,In_151);
xor U959 (N_959,In_1394,In_559);
and U960 (N_960,In_1448,In_636);
nor U961 (N_961,In_552,In_774);
or U962 (N_962,In_310,In_280);
nand U963 (N_963,In_32,In_1264);
and U964 (N_964,In_1091,In_1371);
nor U965 (N_965,In_1322,In_989);
and U966 (N_966,In_762,In_1166);
nand U967 (N_967,In_98,In_2);
and U968 (N_968,In_973,In_113);
or U969 (N_969,In_184,In_1042);
and U970 (N_970,In_225,In_1375);
or U971 (N_971,In_209,In_543);
nor U972 (N_972,In_814,In_1218);
nor U973 (N_973,In_1451,In_1376);
and U974 (N_974,In_1143,In_487);
xnor U975 (N_975,In_1016,In_34);
nor U976 (N_976,In_233,In_1389);
nor U977 (N_977,In_99,In_1290);
nand U978 (N_978,In_989,In_150);
and U979 (N_979,In_691,In_514);
nand U980 (N_980,In_955,In_565);
and U981 (N_981,In_488,In_776);
nor U982 (N_982,In_1061,In_1426);
and U983 (N_983,In_570,In_168);
nand U984 (N_984,In_533,In_311);
nand U985 (N_985,In_1213,In_761);
nand U986 (N_986,In_757,In_426);
nor U987 (N_987,In_616,In_320);
nand U988 (N_988,In_786,In_1191);
and U989 (N_989,In_778,In_466);
and U990 (N_990,In_1153,In_172);
nor U991 (N_991,In_474,In_1108);
nand U992 (N_992,In_1394,In_703);
or U993 (N_993,In_788,In_303);
nor U994 (N_994,In_694,In_1055);
nand U995 (N_995,In_1304,In_334);
nor U996 (N_996,In_440,In_1460);
nor U997 (N_997,In_1460,In_38);
or U998 (N_998,In_930,In_1333);
and U999 (N_999,In_1080,In_805);
nand U1000 (N_1000,In_95,In_1325);
and U1001 (N_1001,In_1162,In_1029);
or U1002 (N_1002,In_854,In_1096);
nand U1003 (N_1003,In_1044,In_15);
or U1004 (N_1004,In_890,In_280);
or U1005 (N_1005,In_1225,In_1151);
or U1006 (N_1006,In_1364,In_87);
nor U1007 (N_1007,In_1060,In_860);
or U1008 (N_1008,In_841,In_1291);
nor U1009 (N_1009,In_1212,In_437);
or U1010 (N_1010,In_823,In_245);
xor U1011 (N_1011,In_476,In_117);
nor U1012 (N_1012,In_1276,In_1250);
and U1013 (N_1013,In_458,In_494);
nand U1014 (N_1014,In_635,In_858);
or U1015 (N_1015,In_951,In_1339);
nor U1016 (N_1016,In_690,In_177);
and U1017 (N_1017,In_1333,In_1237);
and U1018 (N_1018,In_1129,In_373);
nand U1019 (N_1019,In_1201,In_970);
nor U1020 (N_1020,In_1380,In_996);
nand U1021 (N_1021,In_375,In_662);
nand U1022 (N_1022,In_1034,In_705);
nor U1023 (N_1023,In_1448,In_707);
xnor U1024 (N_1024,In_90,In_1152);
and U1025 (N_1025,In_361,In_178);
nand U1026 (N_1026,In_1398,In_19);
or U1027 (N_1027,In_620,In_261);
or U1028 (N_1028,In_1141,In_264);
and U1029 (N_1029,In_1311,In_1165);
and U1030 (N_1030,In_316,In_508);
nor U1031 (N_1031,In_670,In_1363);
nand U1032 (N_1032,In_569,In_885);
and U1033 (N_1033,In_955,In_195);
nand U1034 (N_1034,In_1125,In_1280);
nor U1035 (N_1035,In_936,In_207);
and U1036 (N_1036,In_878,In_667);
nand U1037 (N_1037,In_1362,In_1160);
or U1038 (N_1038,In_247,In_268);
nor U1039 (N_1039,In_915,In_1462);
nand U1040 (N_1040,In_66,In_1258);
and U1041 (N_1041,In_1193,In_678);
nand U1042 (N_1042,In_702,In_334);
or U1043 (N_1043,In_341,In_106);
or U1044 (N_1044,In_73,In_1310);
or U1045 (N_1045,In_797,In_607);
and U1046 (N_1046,In_364,In_247);
or U1047 (N_1047,In_1474,In_364);
nand U1048 (N_1048,In_1121,In_12);
and U1049 (N_1049,In_61,In_1327);
and U1050 (N_1050,In_1182,In_246);
nor U1051 (N_1051,In_1287,In_35);
and U1052 (N_1052,In_203,In_1158);
nand U1053 (N_1053,In_1027,In_1486);
nor U1054 (N_1054,In_157,In_823);
and U1055 (N_1055,In_1235,In_497);
or U1056 (N_1056,In_277,In_525);
and U1057 (N_1057,In_164,In_1364);
or U1058 (N_1058,In_1104,In_919);
or U1059 (N_1059,In_601,In_914);
and U1060 (N_1060,In_479,In_992);
and U1061 (N_1061,In_510,In_867);
nand U1062 (N_1062,In_647,In_285);
nand U1063 (N_1063,In_597,In_1319);
nor U1064 (N_1064,In_1367,In_706);
or U1065 (N_1065,In_776,In_1298);
and U1066 (N_1066,In_627,In_567);
or U1067 (N_1067,In_1208,In_782);
nand U1068 (N_1068,In_188,In_211);
and U1069 (N_1069,In_1262,In_1461);
or U1070 (N_1070,In_100,In_752);
or U1071 (N_1071,In_53,In_89);
nand U1072 (N_1072,In_603,In_43);
nor U1073 (N_1073,In_925,In_149);
nand U1074 (N_1074,In_517,In_149);
or U1075 (N_1075,In_715,In_805);
and U1076 (N_1076,In_1201,In_86);
nand U1077 (N_1077,In_1364,In_209);
or U1078 (N_1078,In_1328,In_815);
nor U1079 (N_1079,In_1238,In_1345);
or U1080 (N_1080,In_234,In_1032);
and U1081 (N_1081,In_102,In_949);
nor U1082 (N_1082,In_624,In_928);
or U1083 (N_1083,In_731,In_510);
and U1084 (N_1084,In_1376,In_490);
and U1085 (N_1085,In_775,In_818);
or U1086 (N_1086,In_15,In_580);
or U1087 (N_1087,In_1479,In_341);
nor U1088 (N_1088,In_956,In_1458);
or U1089 (N_1089,In_1359,In_1036);
nor U1090 (N_1090,In_863,In_555);
xnor U1091 (N_1091,In_1351,In_82);
and U1092 (N_1092,In_1052,In_1421);
or U1093 (N_1093,In_1324,In_467);
and U1094 (N_1094,In_1064,In_430);
nor U1095 (N_1095,In_65,In_266);
and U1096 (N_1096,In_252,In_295);
nor U1097 (N_1097,In_774,In_670);
or U1098 (N_1098,In_1164,In_1321);
nand U1099 (N_1099,In_380,In_52);
nand U1100 (N_1100,In_445,In_111);
nand U1101 (N_1101,In_1060,In_573);
nand U1102 (N_1102,In_947,In_1042);
nor U1103 (N_1103,In_668,In_289);
nand U1104 (N_1104,In_556,In_109);
and U1105 (N_1105,In_168,In_129);
or U1106 (N_1106,In_1173,In_682);
nor U1107 (N_1107,In_573,In_386);
xor U1108 (N_1108,In_850,In_744);
nor U1109 (N_1109,In_644,In_105);
nand U1110 (N_1110,In_1257,In_313);
nand U1111 (N_1111,In_41,In_748);
or U1112 (N_1112,In_378,In_921);
or U1113 (N_1113,In_956,In_1205);
nand U1114 (N_1114,In_659,In_774);
or U1115 (N_1115,In_1353,In_395);
nor U1116 (N_1116,In_1454,In_775);
and U1117 (N_1117,In_1388,In_1054);
nand U1118 (N_1118,In_1068,In_687);
and U1119 (N_1119,In_1444,In_964);
or U1120 (N_1120,In_1221,In_856);
or U1121 (N_1121,In_406,In_1107);
and U1122 (N_1122,In_1308,In_882);
and U1123 (N_1123,In_1046,In_1442);
nand U1124 (N_1124,In_1387,In_933);
or U1125 (N_1125,In_761,In_805);
nand U1126 (N_1126,In_1141,In_1069);
or U1127 (N_1127,In_309,In_1061);
nor U1128 (N_1128,In_1417,In_1307);
nand U1129 (N_1129,In_1360,In_931);
and U1130 (N_1130,In_507,In_709);
or U1131 (N_1131,In_395,In_420);
and U1132 (N_1132,In_970,In_1436);
or U1133 (N_1133,In_768,In_580);
nand U1134 (N_1134,In_328,In_751);
and U1135 (N_1135,In_1035,In_1120);
and U1136 (N_1136,In_150,In_1469);
nor U1137 (N_1137,In_255,In_611);
and U1138 (N_1138,In_284,In_273);
and U1139 (N_1139,In_1400,In_1053);
nand U1140 (N_1140,In_1476,In_733);
and U1141 (N_1141,In_625,In_759);
or U1142 (N_1142,In_1164,In_275);
and U1143 (N_1143,In_528,In_1142);
or U1144 (N_1144,In_1193,In_1318);
and U1145 (N_1145,In_151,In_1083);
nand U1146 (N_1146,In_277,In_252);
and U1147 (N_1147,In_349,In_767);
or U1148 (N_1148,In_1156,In_1338);
nand U1149 (N_1149,In_3,In_476);
or U1150 (N_1150,In_8,In_881);
or U1151 (N_1151,In_594,In_193);
nor U1152 (N_1152,In_880,In_501);
and U1153 (N_1153,In_1303,In_165);
nor U1154 (N_1154,In_1449,In_747);
nand U1155 (N_1155,In_11,In_18);
and U1156 (N_1156,In_777,In_1093);
or U1157 (N_1157,In_1199,In_450);
or U1158 (N_1158,In_744,In_1083);
nor U1159 (N_1159,In_809,In_1240);
or U1160 (N_1160,In_860,In_877);
and U1161 (N_1161,In_227,In_29);
and U1162 (N_1162,In_1352,In_1159);
nand U1163 (N_1163,In_883,In_457);
xor U1164 (N_1164,In_801,In_716);
and U1165 (N_1165,In_1148,In_672);
and U1166 (N_1166,In_373,In_715);
or U1167 (N_1167,In_200,In_676);
and U1168 (N_1168,In_894,In_1269);
nor U1169 (N_1169,In_1114,In_728);
nand U1170 (N_1170,In_750,In_16);
or U1171 (N_1171,In_373,In_328);
xor U1172 (N_1172,In_666,In_1067);
and U1173 (N_1173,In_673,In_467);
nand U1174 (N_1174,In_864,In_965);
or U1175 (N_1175,In_777,In_360);
nor U1176 (N_1176,In_761,In_889);
nor U1177 (N_1177,In_524,In_1167);
nor U1178 (N_1178,In_1248,In_983);
or U1179 (N_1179,In_524,In_1481);
nor U1180 (N_1180,In_140,In_366);
and U1181 (N_1181,In_1081,In_125);
or U1182 (N_1182,In_83,In_323);
nand U1183 (N_1183,In_199,In_166);
xor U1184 (N_1184,In_180,In_568);
nor U1185 (N_1185,In_1105,In_1172);
or U1186 (N_1186,In_431,In_822);
nor U1187 (N_1187,In_719,In_136);
nor U1188 (N_1188,In_1166,In_373);
and U1189 (N_1189,In_1433,In_631);
and U1190 (N_1190,In_1168,In_1063);
and U1191 (N_1191,In_897,In_1409);
nand U1192 (N_1192,In_138,In_483);
nand U1193 (N_1193,In_1485,In_912);
or U1194 (N_1194,In_55,In_1320);
nor U1195 (N_1195,In_449,In_560);
and U1196 (N_1196,In_199,In_512);
xnor U1197 (N_1197,In_1187,In_1102);
or U1198 (N_1198,In_731,In_518);
or U1199 (N_1199,In_886,In_320);
and U1200 (N_1200,In_241,In_1258);
nand U1201 (N_1201,In_1008,In_808);
or U1202 (N_1202,In_1133,In_1388);
or U1203 (N_1203,In_918,In_362);
nand U1204 (N_1204,In_584,In_888);
nand U1205 (N_1205,In_420,In_939);
or U1206 (N_1206,In_734,In_647);
nor U1207 (N_1207,In_141,In_159);
nor U1208 (N_1208,In_100,In_1038);
nor U1209 (N_1209,In_934,In_705);
or U1210 (N_1210,In_914,In_449);
nor U1211 (N_1211,In_701,In_646);
nand U1212 (N_1212,In_794,In_1021);
nor U1213 (N_1213,In_791,In_1089);
and U1214 (N_1214,In_983,In_410);
or U1215 (N_1215,In_214,In_975);
and U1216 (N_1216,In_77,In_533);
nor U1217 (N_1217,In_414,In_1132);
and U1218 (N_1218,In_502,In_1149);
and U1219 (N_1219,In_1142,In_587);
xor U1220 (N_1220,In_313,In_647);
or U1221 (N_1221,In_996,In_877);
and U1222 (N_1222,In_997,In_227);
and U1223 (N_1223,In_1326,In_940);
or U1224 (N_1224,In_727,In_1482);
nand U1225 (N_1225,In_167,In_656);
and U1226 (N_1226,In_62,In_208);
and U1227 (N_1227,In_334,In_1101);
nor U1228 (N_1228,In_1376,In_712);
nand U1229 (N_1229,In_495,In_837);
and U1230 (N_1230,In_1002,In_11);
nand U1231 (N_1231,In_1151,In_506);
nor U1232 (N_1232,In_447,In_1493);
nor U1233 (N_1233,In_879,In_377);
nand U1234 (N_1234,In_149,In_827);
or U1235 (N_1235,In_1386,In_1311);
nand U1236 (N_1236,In_1468,In_366);
nor U1237 (N_1237,In_1329,In_731);
nor U1238 (N_1238,In_1087,In_1462);
and U1239 (N_1239,In_104,In_458);
and U1240 (N_1240,In_532,In_679);
and U1241 (N_1241,In_855,In_838);
nor U1242 (N_1242,In_1475,In_1484);
nand U1243 (N_1243,In_980,In_626);
nand U1244 (N_1244,In_1302,In_1100);
or U1245 (N_1245,In_276,In_825);
and U1246 (N_1246,In_725,In_365);
and U1247 (N_1247,In_52,In_459);
and U1248 (N_1248,In_458,In_1445);
and U1249 (N_1249,In_1088,In_324);
or U1250 (N_1250,In_1324,In_762);
and U1251 (N_1251,In_768,In_270);
or U1252 (N_1252,In_9,In_148);
and U1253 (N_1253,In_1062,In_988);
and U1254 (N_1254,In_283,In_879);
or U1255 (N_1255,In_781,In_1239);
nand U1256 (N_1256,In_163,In_1307);
nor U1257 (N_1257,In_653,In_960);
and U1258 (N_1258,In_165,In_810);
nor U1259 (N_1259,In_1251,In_384);
nor U1260 (N_1260,In_1362,In_352);
or U1261 (N_1261,In_642,In_322);
nor U1262 (N_1262,In_1421,In_191);
or U1263 (N_1263,In_1088,In_830);
or U1264 (N_1264,In_170,In_936);
nor U1265 (N_1265,In_1456,In_782);
nand U1266 (N_1266,In_337,In_846);
or U1267 (N_1267,In_560,In_21);
nor U1268 (N_1268,In_1140,In_16);
and U1269 (N_1269,In_962,In_544);
or U1270 (N_1270,In_1286,In_897);
and U1271 (N_1271,In_336,In_930);
and U1272 (N_1272,In_705,In_719);
nor U1273 (N_1273,In_1290,In_915);
nor U1274 (N_1274,In_538,In_701);
and U1275 (N_1275,In_273,In_238);
and U1276 (N_1276,In_636,In_273);
nand U1277 (N_1277,In_692,In_400);
and U1278 (N_1278,In_1128,In_1251);
and U1279 (N_1279,In_379,In_1276);
nand U1280 (N_1280,In_609,In_50);
and U1281 (N_1281,In_1320,In_1439);
and U1282 (N_1282,In_268,In_853);
xor U1283 (N_1283,In_1198,In_1392);
or U1284 (N_1284,In_362,In_1267);
nor U1285 (N_1285,In_612,In_155);
and U1286 (N_1286,In_256,In_1122);
and U1287 (N_1287,In_1218,In_524);
and U1288 (N_1288,In_156,In_423);
nor U1289 (N_1289,In_1082,In_653);
or U1290 (N_1290,In_556,In_1369);
nor U1291 (N_1291,In_1136,In_849);
or U1292 (N_1292,In_170,In_1203);
or U1293 (N_1293,In_1256,In_250);
nor U1294 (N_1294,In_553,In_390);
xor U1295 (N_1295,In_261,In_1136);
or U1296 (N_1296,In_62,In_280);
nor U1297 (N_1297,In_1428,In_749);
or U1298 (N_1298,In_843,In_1471);
or U1299 (N_1299,In_1013,In_312);
nor U1300 (N_1300,In_793,In_1418);
nand U1301 (N_1301,In_1295,In_991);
and U1302 (N_1302,In_787,In_935);
and U1303 (N_1303,In_804,In_630);
nor U1304 (N_1304,In_920,In_941);
and U1305 (N_1305,In_122,In_504);
nand U1306 (N_1306,In_871,In_560);
nor U1307 (N_1307,In_1212,In_803);
nand U1308 (N_1308,In_67,In_675);
and U1309 (N_1309,In_358,In_695);
and U1310 (N_1310,In_195,In_741);
or U1311 (N_1311,In_185,In_241);
and U1312 (N_1312,In_562,In_1074);
or U1313 (N_1313,In_354,In_169);
xor U1314 (N_1314,In_913,In_615);
nor U1315 (N_1315,In_1136,In_1395);
nor U1316 (N_1316,In_874,In_887);
nand U1317 (N_1317,In_683,In_1323);
or U1318 (N_1318,In_696,In_1374);
and U1319 (N_1319,In_39,In_519);
and U1320 (N_1320,In_128,In_1436);
and U1321 (N_1321,In_1182,In_1119);
nor U1322 (N_1322,In_152,In_200);
and U1323 (N_1323,In_991,In_148);
nand U1324 (N_1324,In_218,In_635);
nand U1325 (N_1325,In_385,In_172);
nand U1326 (N_1326,In_731,In_757);
nor U1327 (N_1327,In_360,In_901);
or U1328 (N_1328,In_1293,In_77);
or U1329 (N_1329,In_877,In_81);
and U1330 (N_1330,In_1499,In_221);
nor U1331 (N_1331,In_1250,In_1113);
nand U1332 (N_1332,In_1039,In_555);
nand U1333 (N_1333,In_736,In_683);
and U1334 (N_1334,In_919,In_495);
and U1335 (N_1335,In_356,In_511);
or U1336 (N_1336,In_969,In_1242);
nand U1337 (N_1337,In_672,In_676);
nand U1338 (N_1338,In_1334,In_584);
or U1339 (N_1339,In_296,In_1240);
nor U1340 (N_1340,In_835,In_269);
or U1341 (N_1341,In_702,In_1265);
nor U1342 (N_1342,In_930,In_978);
nand U1343 (N_1343,In_934,In_350);
nand U1344 (N_1344,In_1440,In_1192);
or U1345 (N_1345,In_1345,In_656);
or U1346 (N_1346,In_538,In_629);
or U1347 (N_1347,In_50,In_545);
or U1348 (N_1348,In_129,In_188);
and U1349 (N_1349,In_896,In_323);
and U1350 (N_1350,In_114,In_557);
nor U1351 (N_1351,In_248,In_962);
or U1352 (N_1352,In_887,In_1282);
nor U1353 (N_1353,In_1215,In_1396);
or U1354 (N_1354,In_304,In_1445);
or U1355 (N_1355,In_285,In_967);
and U1356 (N_1356,In_236,In_973);
nand U1357 (N_1357,In_182,In_885);
and U1358 (N_1358,In_1247,In_1484);
nor U1359 (N_1359,In_1017,In_669);
and U1360 (N_1360,In_117,In_1448);
and U1361 (N_1361,In_86,In_621);
or U1362 (N_1362,In_475,In_1490);
nor U1363 (N_1363,In_770,In_1276);
nor U1364 (N_1364,In_592,In_1296);
nand U1365 (N_1365,In_597,In_27);
nand U1366 (N_1366,In_295,In_828);
nand U1367 (N_1367,In_1121,In_698);
or U1368 (N_1368,In_799,In_1087);
nand U1369 (N_1369,In_806,In_835);
xnor U1370 (N_1370,In_475,In_400);
nand U1371 (N_1371,In_1020,In_1470);
nand U1372 (N_1372,In_468,In_425);
nand U1373 (N_1373,In_809,In_233);
and U1374 (N_1374,In_135,In_385);
nor U1375 (N_1375,In_199,In_1155);
or U1376 (N_1376,In_507,In_197);
nand U1377 (N_1377,In_385,In_961);
nand U1378 (N_1378,In_1101,In_964);
and U1379 (N_1379,In_865,In_995);
nand U1380 (N_1380,In_585,In_755);
or U1381 (N_1381,In_589,In_458);
nor U1382 (N_1382,In_516,In_935);
nor U1383 (N_1383,In_1444,In_1083);
and U1384 (N_1384,In_89,In_1467);
nand U1385 (N_1385,In_269,In_796);
or U1386 (N_1386,In_525,In_311);
nor U1387 (N_1387,In_533,In_534);
nand U1388 (N_1388,In_871,In_683);
nand U1389 (N_1389,In_321,In_17);
and U1390 (N_1390,In_175,In_850);
nor U1391 (N_1391,In_613,In_498);
nand U1392 (N_1392,In_742,In_370);
and U1393 (N_1393,In_1145,In_1206);
nand U1394 (N_1394,In_87,In_1401);
or U1395 (N_1395,In_840,In_335);
nor U1396 (N_1396,In_837,In_1371);
and U1397 (N_1397,In_1062,In_1138);
nor U1398 (N_1398,In_979,In_673);
and U1399 (N_1399,In_346,In_121);
xor U1400 (N_1400,In_117,In_917);
nand U1401 (N_1401,In_839,In_1075);
and U1402 (N_1402,In_281,In_501);
nor U1403 (N_1403,In_1103,In_476);
nand U1404 (N_1404,In_1424,In_1484);
and U1405 (N_1405,In_1149,In_249);
nor U1406 (N_1406,In_1389,In_96);
nand U1407 (N_1407,In_1080,In_653);
xor U1408 (N_1408,In_1463,In_240);
or U1409 (N_1409,In_644,In_179);
and U1410 (N_1410,In_620,In_1446);
or U1411 (N_1411,In_923,In_238);
or U1412 (N_1412,In_1266,In_1001);
or U1413 (N_1413,In_924,In_409);
nand U1414 (N_1414,In_1432,In_1068);
or U1415 (N_1415,In_765,In_1351);
or U1416 (N_1416,In_1012,In_958);
or U1417 (N_1417,In_37,In_1128);
and U1418 (N_1418,In_611,In_1312);
and U1419 (N_1419,In_189,In_955);
nor U1420 (N_1420,In_773,In_226);
and U1421 (N_1421,In_1452,In_160);
or U1422 (N_1422,In_76,In_399);
nand U1423 (N_1423,In_1192,In_638);
xnor U1424 (N_1424,In_297,In_899);
nor U1425 (N_1425,In_335,In_202);
and U1426 (N_1426,In_726,In_1300);
or U1427 (N_1427,In_1496,In_310);
and U1428 (N_1428,In_691,In_1029);
and U1429 (N_1429,In_134,In_1128);
nand U1430 (N_1430,In_495,In_16);
nand U1431 (N_1431,In_895,In_258);
nor U1432 (N_1432,In_1129,In_168);
nor U1433 (N_1433,In_489,In_463);
or U1434 (N_1434,In_1053,In_985);
nand U1435 (N_1435,In_37,In_392);
and U1436 (N_1436,In_251,In_553);
and U1437 (N_1437,In_727,In_1045);
or U1438 (N_1438,In_25,In_1404);
and U1439 (N_1439,In_289,In_957);
nor U1440 (N_1440,In_908,In_706);
nor U1441 (N_1441,In_163,In_471);
nor U1442 (N_1442,In_1011,In_1235);
nand U1443 (N_1443,In_203,In_374);
nand U1444 (N_1444,In_263,In_534);
or U1445 (N_1445,In_658,In_766);
nand U1446 (N_1446,In_648,In_1192);
nand U1447 (N_1447,In_39,In_205);
xnor U1448 (N_1448,In_1119,In_149);
nand U1449 (N_1449,In_135,In_277);
or U1450 (N_1450,In_1133,In_1248);
or U1451 (N_1451,In_22,In_216);
nor U1452 (N_1452,In_180,In_614);
nand U1453 (N_1453,In_225,In_178);
and U1454 (N_1454,In_416,In_1009);
and U1455 (N_1455,In_424,In_1490);
nand U1456 (N_1456,In_47,In_946);
or U1457 (N_1457,In_311,In_1032);
or U1458 (N_1458,In_709,In_1421);
or U1459 (N_1459,In_314,In_1369);
or U1460 (N_1460,In_793,In_849);
and U1461 (N_1461,In_545,In_524);
nand U1462 (N_1462,In_177,In_523);
or U1463 (N_1463,In_1015,In_695);
and U1464 (N_1464,In_1286,In_1028);
and U1465 (N_1465,In_615,In_816);
nand U1466 (N_1466,In_572,In_957);
nor U1467 (N_1467,In_167,In_869);
nor U1468 (N_1468,In_138,In_470);
and U1469 (N_1469,In_631,In_1181);
nor U1470 (N_1470,In_886,In_888);
or U1471 (N_1471,In_551,In_904);
or U1472 (N_1472,In_188,In_163);
or U1473 (N_1473,In_484,In_499);
nand U1474 (N_1474,In_1006,In_1400);
nor U1475 (N_1475,In_1045,In_1240);
xnor U1476 (N_1476,In_467,In_18);
nand U1477 (N_1477,In_4,In_6);
or U1478 (N_1478,In_1076,In_1045);
and U1479 (N_1479,In_1296,In_625);
and U1480 (N_1480,In_426,In_889);
xnor U1481 (N_1481,In_1114,In_368);
or U1482 (N_1482,In_503,In_1156);
nor U1483 (N_1483,In_926,In_66);
nor U1484 (N_1484,In_462,In_804);
and U1485 (N_1485,In_311,In_223);
xor U1486 (N_1486,In_603,In_1125);
or U1487 (N_1487,In_845,In_1225);
and U1488 (N_1488,In_77,In_239);
and U1489 (N_1489,In_663,In_784);
and U1490 (N_1490,In_1161,In_15);
nor U1491 (N_1491,In_574,In_1129);
or U1492 (N_1492,In_892,In_1194);
and U1493 (N_1493,In_888,In_1136);
or U1494 (N_1494,In_761,In_363);
or U1495 (N_1495,In_1148,In_576);
nand U1496 (N_1496,In_1066,In_1454);
and U1497 (N_1497,In_1171,In_1439);
nand U1498 (N_1498,In_764,In_964);
nand U1499 (N_1499,In_507,In_612);
and U1500 (N_1500,In_206,In_96);
nor U1501 (N_1501,In_646,In_950);
nand U1502 (N_1502,In_1427,In_189);
nand U1503 (N_1503,In_759,In_521);
and U1504 (N_1504,In_442,In_248);
and U1505 (N_1505,In_1075,In_285);
nand U1506 (N_1506,In_1437,In_136);
and U1507 (N_1507,In_473,In_1189);
nand U1508 (N_1508,In_261,In_409);
nor U1509 (N_1509,In_1023,In_708);
nor U1510 (N_1510,In_1384,In_701);
nor U1511 (N_1511,In_423,In_428);
xnor U1512 (N_1512,In_178,In_1219);
and U1513 (N_1513,In_181,In_865);
nor U1514 (N_1514,In_1482,In_1491);
xor U1515 (N_1515,In_19,In_354);
nand U1516 (N_1516,In_98,In_1406);
and U1517 (N_1517,In_758,In_225);
nand U1518 (N_1518,In_920,In_20);
nand U1519 (N_1519,In_878,In_77);
nand U1520 (N_1520,In_102,In_383);
nand U1521 (N_1521,In_334,In_576);
and U1522 (N_1522,In_941,In_1475);
nor U1523 (N_1523,In_211,In_969);
nand U1524 (N_1524,In_1097,In_1196);
and U1525 (N_1525,In_1014,In_432);
or U1526 (N_1526,In_620,In_535);
or U1527 (N_1527,In_347,In_1255);
or U1528 (N_1528,In_1136,In_1470);
xnor U1529 (N_1529,In_479,In_601);
or U1530 (N_1530,In_46,In_366);
nor U1531 (N_1531,In_859,In_420);
nor U1532 (N_1532,In_1085,In_1399);
xor U1533 (N_1533,In_1077,In_131);
nor U1534 (N_1534,In_1312,In_24);
nor U1535 (N_1535,In_1131,In_985);
nor U1536 (N_1536,In_1412,In_1499);
nor U1537 (N_1537,In_221,In_541);
and U1538 (N_1538,In_139,In_1168);
nor U1539 (N_1539,In_257,In_1461);
nor U1540 (N_1540,In_1498,In_1110);
nor U1541 (N_1541,In_708,In_12);
nor U1542 (N_1542,In_87,In_566);
or U1543 (N_1543,In_487,In_1122);
and U1544 (N_1544,In_1289,In_544);
nand U1545 (N_1545,In_266,In_1113);
nor U1546 (N_1546,In_787,In_452);
nor U1547 (N_1547,In_636,In_405);
xor U1548 (N_1548,In_563,In_243);
nor U1549 (N_1549,In_1267,In_163);
and U1550 (N_1550,In_780,In_1305);
nor U1551 (N_1551,In_447,In_1413);
and U1552 (N_1552,In_614,In_469);
nand U1553 (N_1553,In_919,In_1467);
and U1554 (N_1554,In_444,In_879);
and U1555 (N_1555,In_1273,In_1358);
or U1556 (N_1556,In_563,In_1120);
and U1557 (N_1557,In_76,In_956);
nor U1558 (N_1558,In_35,In_800);
or U1559 (N_1559,In_1450,In_1237);
and U1560 (N_1560,In_1194,In_869);
nand U1561 (N_1561,In_515,In_932);
or U1562 (N_1562,In_825,In_57);
or U1563 (N_1563,In_426,In_488);
nor U1564 (N_1564,In_737,In_1157);
nor U1565 (N_1565,In_836,In_603);
and U1566 (N_1566,In_1023,In_395);
or U1567 (N_1567,In_631,In_811);
nand U1568 (N_1568,In_1309,In_1088);
nand U1569 (N_1569,In_630,In_731);
or U1570 (N_1570,In_575,In_200);
and U1571 (N_1571,In_622,In_1375);
and U1572 (N_1572,In_603,In_251);
and U1573 (N_1573,In_272,In_769);
nor U1574 (N_1574,In_18,In_940);
or U1575 (N_1575,In_1326,In_558);
or U1576 (N_1576,In_950,In_383);
nor U1577 (N_1577,In_505,In_1209);
nor U1578 (N_1578,In_42,In_971);
xnor U1579 (N_1579,In_95,In_433);
nor U1580 (N_1580,In_694,In_180);
nor U1581 (N_1581,In_1456,In_968);
nor U1582 (N_1582,In_1267,In_1019);
and U1583 (N_1583,In_375,In_837);
xnor U1584 (N_1584,In_754,In_540);
nand U1585 (N_1585,In_69,In_648);
nand U1586 (N_1586,In_428,In_1184);
and U1587 (N_1587,In_1453,In_255);
nand U1588 (N_1588,In_1029,In_847);
nor U1589 (N_1589,In_460,In_235);
nor U1590 (N_1590,In_548,In_795);
nand U1591 (N_1591,In_1353,In_869);
or U1592 (N_1592,In_1169,In_99);
or U1593 (N_1593,In_1041,In_271);
nand U1594 (N_1594,In_943,In_651);
nor U1595 (N_1595,In_949,In_893);
nor U1596 (N_1596,In_1085,In_424);
nor U1597 (N_1597,In_127,In_612);
and U1598 (N_1598,In_1132,In_1037);
or U1599 (N_1599,In_267,In_101);
or U1600 (N_1600,In_702,In_453);
nand U1601 (N_1601,In_175,In_646);
and U1602 (N_1602,In_1062,In_917);
and U1603 (N_1603,In_1400,In_1240);
nand U1604 (N_1604,In_590,In_857);
or U1605 (N_1605,In_272,In_1487);
nand U1606 (N_1606,In_302,In_1482);
nor U1607 (N_1607,In_537,In_1117);
and U1608 (N_1608,In_302,In_1362);
nand U1609 (N_1609,In_951,In_234);
nor U1610 (N_1610,In_1411,In_455);
nand U1611 (N_1611,In_752,In_162);
nor U1612 (N_1612,In_476,In_1054);
nand U1613 (N_1613,In_578,In_1490);
nand U1614 (N_1614,In_834,In_1398);
nor U1615 (N_1615,In_527,In_1170);
nand U1616 (N_1616,In_676,In_685);
xnor U1617 (N_1617,In_1404,In_154);
nand U1618 (N_1618,In_863,In_1473);
or U1619 (N_1619,In_1063,In_1481);
or U1620 (N_1620,In_1435,In_146);
nor U1621 (N_1621,In_295,In_1413);
xnor U1622 (N_1622,In_108,In_804);
and U1623 (N_1623,In_931,In_806);
nor U1624 (N_1624,In_822,In_458);
or U1625 (N_1625,In_637,In_691);
nand U1626 (N_1626,In_297,In_1415);
or U1627 (N_1627,In_1030,In_1199);
and U1628 (N_1628,In_807,In_585);
nor U1629 (N_1629,In_97,In_1456);
nor U1630 (N_1630,In_774,In_268);
nor U1631 (N_1631,In_245,In_1427);
and U1632 (N_1632,In_394,In_468);
nor U1633 (N_1633,In_496,In_287);
nand U1634 (N_1634,In_852,In_522);
and U1635 (N_1635,In_467,In_16);
and U1636 (N_1636,In_436,In_1125);
or U1637 (N_1637,In_3,In_614);
nor U1638 (N_1638,In_1006,In_951);
and U1639 (N_1639,In_1015,In_192);
or U1640 (N_1640,In_299,In_997);
nand U1641 (N_1641,In_647,In_2);
or U1642 (N_1642,In_423,In_458);
nor U1643 (N_1643,In_964,In_203);
nand U1644 (N_1644,In_845,In_751);
or U1645 (N_1645,In_87,In_1461);
or U1646 (N_1646,In_87,In_822);
and U1647 (N_1647,In_180,In_213);
nand U1648 (N_1648,In_937,In_1060);
nor U1649 (N_1649,In_750,In_29);
nand U1650 (N_1650,In_1169,In_852);
and U1651 (N_1651,In_114,In_1291);
nor U1652 (N_1652,In_532,In_357);
or U1653 (N_1653,In_1031,In_426);
and U1654 (N_1654,In_584,In_21);
or U1655 (N_1655,In_406,In_179);
and U1656 (N_1656,In_1210,In_962);
or U1657 (N_1657,In_496,In_278);
and U1658 (N_1658,In_1483,In_963);
nor U1659 (N_1659,In_569,In_201);
and U1660 (N_1660,In_362,In_577);
nand U1661 (N_1661,In_1188,In_1422);
nor U1662 (N_1662,In_821,In_1031);
nand U1663 (N_1663,In_182,In_10);
and U1664 (N_1664,In_784,In_1465);
nand U1665 (N_1665,In_791,In_888);
nor U1666 (N_1666,In_1103,In_1168);
nand U1667 (N_1667,In_404,In_1429);
or U1668 (N_1668,In_458,In_693);
and U1669 (N_1669,In_1386,In_831);
or U1670 (N_1670,In_407,In_596);
or U1671 (N_1671,In_1169,In_954);
nand U1672 (N_1672,In_1105,In_430);
and U1673 (N_1673,In_57,In_553);
nor U1674 (N_1674,In_867,In_1153);
nand U1675 (N_1675,In_113,In_438);
nor U1676 (N_1676,In_885,In_1246);
nand U1677 (N_1677,In_672,In_182);
nor U1678 (N_1678,In_1088,In_949);
or U1679 (N_1679,In_858,In_1150);
or U1680 (N_1680,In_342,In_1183);
nor U1681 (N_1681,In_427,In_556);
nand U1682 (N_1682,In_1476,In_738);
or U1683 (N_1683,In_1361,In_754);
nor U1684 (N_1684,In_346,In_1273);
nand U1685 (N_1685,In_1487,In_1427);
nor U1686 (N_1686,In_204,In_1144);
and U1687 (N_1687,In_1378,In_894);
and U1688 (N_1688,In_800,In_348);
and U1689 (N_1689,In_1425,In_1072);
and U1690 (N_1690,In_1312,In_155);
or U1691 (N_1691,In_1204,In_1216);
nand U1692 (N_1692,In_973,In_1156);
and U1693 (N_1693,In_527,In_197);
or U1694 (N_1694,In_192,In_1204);
nor U1695 (N_1695,In_365,In_533);
nand U1696 (N_1696,In_873,In_850);
nand U1697 (N_1697,In_890,In_1318);
nand U1698 (N_1698,In_208,In_919);
nand U1699 (N_1699,In_1223,In_920);
and U1700 (N_1700,In_805,In_504);
and U1701 (N_1701,In_712,In_894);
nor U1702 (N_1702,In_43,In_1237);
nand U1703 (N_1703,In_237,In_1305);
nor U1704 (N_1704,In_587,In_1348);
or U1705 (N_1705,In_223,In_559);
and U1706 (N_1706,In_1249,In_1202);
nand U1707 (N_1707,In_333,In_343);
or U1708 (N_1708,In_486,In_1324);
nor U1709 (N_1709,In_1369,In_763);
nand U1710 (N_1710,In_887,In_845);
nor U1711 (N_1711,In_791,In_419);
nor U1712 (N_1712,In_1073,In_123);
nand U1713 (N_1713,In_1374,In_1245);
nor U1714 (N_1714,In_1206,In_139);
nor U1715 (N_1715,In_673,In_478);
nand U1716 (N_1716,In_796,In_919);
or U1717 (N_1717,In_1008,In_904);
nor U1718 (N_1718,In_1194,In_1063);
and U1719 (N_1719,In_156,In_574);
and U1720 (N_1720,In_178,In_8);
nor U1721 (N_1721,In_956,In_743);
nor U1722 (N_1722,In_274,In_922);
nor U1723 (N_1723,In_676,In_28);
nor U1724 (N_1724,In_443,In_1122);
and U1725 (N_1725,In_671,In_35);
nand U1726 (N_1726,In_859,In_1103);
xnor U1727 (N_1727,In_796,In_1266);
nand U1728 (N_1728,In_1061,In_1121);
or U1729 (N_1729,In_685,In_1160);
nor U1730 (N_1730,In_248,In_966);
and U1731 (N_1731,In_227,In_97);
and U1732 (N_1732,In_416,In_747);
nor U1733 (N_1733,In_1098,In_1466);
nor U1734 (N_1734,In_820,In_1443);
and U1735 (N_1735,In_682,In_943);
and U1736 (N_1736,In_150,In_503);
or U1737 (N_1737,In_524,In_225);
nand U1738 (N_1738,In_234,In_1215);
nor U1739 (N_1739,In_256,In_1444);
or U1740 (N_1740,In_580,In_1124);
and U1741 (N_1741,In_974,In_967);
or U1742 (N_1742,In_345,In_557);
or U1743 (N_1743,In_617,In_411);
nor U1744 (N_1744,In_816,In_966);
xnor U1745 (N_1745,In_1406,In_810);
nor U1746 (N_1746,In_436,In_406);
nand U1747 (N_1747,In_1202,In_1218);
and U1748 (N_1748,In_463,In_1188);
nand U1749 (N_1749,In_455,In_255);
nor U1750 (N_1750,In_1044,In_919);
nand U1751 (N_1751,In_603,In_983);
nor U1752 (N_1752,In_142,In_1007);
and U1753 (N_1753,In_1211,In_1276);
nand U1754 (N_1754,In_1120,In_467);
and U1755 (N_1755,In_1051,In_820);
or U1756 (N_1756,In_475,In_209);
and U1757 (N_1757,In_1228,In_1316);
nand U1758 (N_1758,In_1358,In_846);
nand U1759 (N_1759,In_1078,In_351);
or U1760 (N_1760,In_390,In_15);
nor U1761 (N_1761,In_165,In_820);
and U1762 (N_1762,In_992,In_332);
or U1763 (N_1763,In_1036,In_1224);
and U1764 (N_1764,In_327,In_405);
or U1765 (N_1765,In_256,In_827);
and U1766 (N_1766,In_69,In_247);
nor U1767 (N_1767,In_1235,In_1152);
and U1768 (N_1768,In_1286,In_394);
and U1769 (N_1769,In_334,In_946);
nor U1770 (N_1770,In_105,In_403);
and U1771 (N_1771,In_977,In_380);
nand U1772 (N_1772,In_1159,In_1036);
nand U1773 (N_1773,In_51,In_668);
or U1774 (N_1774,In_966,In_359);
nand U1775 (N_1775,In_1401,In_1422);
or U1776 (N_1776,In_1265,In_1186);
nor U1777 (N_1777,In_1474,In_11);
nor U1778 (N_1778,In_377,In_443);
nor U1779 (N_1779,In_1459,In_1026);
or U1780 (N_1780,In_938,In_565);
xnor U1781 (N_1781,In_1051,In_1251);
nand U1782 (N_1782,In_1004,In_104);
nor U1783 (N_1783,In_712,In_425);
nor U1784 (N_1784,In_1419,In_516);
and U1785 (N_1785,In_18,In_611);
and U1786 (N_1786,In_565,In_371);
and U1787 (N_1787,In_1488,In_1135);
nand U1788 (N_1788,In_623,In_359);
nor U1789 (N_1789,In_1333,In_876);
nand U1790 (N_1790,In_740,In_876);
or U1791 (N_1791,In_886,In_363);
nor U1792 (N_1792,In_174,In_428);
or U1793 (N_1793,In_150,In_370);
nor U1794 (N_1794,In_217,In_439);
nor U1795 (N_1795,In_907,In_363);
and U1796 (N_1796,In_51,In_252);
nor U1797 (N_1797,In_961,In_1051);
or U1798 (N_1798,In_288,In_880);
or U1799 (N_1799,In_218,In_1194);
nand U1800 (N_1800,In_451,In_270);
and U1801 (N_1801,In_1252,In_1027);
and U1802 (N_1802,In_831,In_1025);
and U1803 (N_1803,In_1448,In_84);
nor U1804 (N_1804,In_1014,In_111);
and U1805 (N_1805,In_929,In_436);
nor U1806 (N_1806,In_1002,In_32);
and U1807 (N_1807,In_175,In_208);
and U1808 (N_1808,In_113,In_1370);
and U1809 (N_1809,In_611,In_1348);
nor U1810 (N_1810,In_445,In_1244);
and U1811 (N_1811,In_741,In_1379);
or U1812 (N_1812,In_1068,In_650);
or U1813 (N_1813,In_214,In_807);
nand U1814 (N_1814,In_580,In_76);
xnor U1815 (N_1815,In_1117,In_1447);
and U1816 (N_1816,In_680,In_640);
nor U1817 (N_1817,In_61,In_1447);
nand U1818 (N_1818,In_79,In_1160);
or U1819 (N_1819,In_856,In_361);
nor U1820 (N_1820,In_1388,In_304);
nor U1821 (N_1821,In_848,In_175);
or U1822 (N_1822,In_673,In_804);
xor U1823 (N_1823,In_27,In_211);
nor U1824 (N_1824,In_235,In_335);
or U1825 (N_1825,In_1113,In_606);
nand U1826 (N_1826,In_207,In_1005);
or U1827 (N_1827,In_400,In_450);
or U1828 (N_1828,In_659,In_288);
nand U1829 (N_1829,In_156,In_350);
nor U1830 (N_1830,In_338,In_679);
nand U1831 (N_1831,In_1474,In_1258);
nand U1832 (N_1832,In_360,In_965);
or U1833 (N_1833,In_496,In_467);
or U1834 (N_1834,In_632,In_1325);
nor U1835 (N_1835,In_1035,In_1341);
or U1836 (N_1836,In_117,In_322);
nor U1837 (N_1837,In_345,In_53);
or U1838 (N_1838,In_1157,In_1152);
and U1839 (N_1839,In_711,In_1186);
nor U1840 (N_1840,In_418,In_1144);
nand U1841 (N_1841,In_281,In_1338);
or U1842 (N_1842,In_443,In_937);
and U1843 (N_1843,In_156,In_1457);
nor U1844 (N_1844,In_748,In_1448);
or U1845 (N_1845,In_307,In_332);
and U1846 (N_1846,In_1012,In_123);
nor U1847 (N_1847,In_1278,In_125);
or U1848 (N_1848,In_819,In_1230);
nor U1849 (N_1849,In_971,In_349);
nor U1850 (N_1850,In_1034,In_7);
nand U1851 (N_1851,In_1086,In_1491);
xor U1852 (N_1852,In_280,In_1477);
nand U1853 (N_1853,In_947,In_1373);
or U1854 (N_1854,In_426,In_1083);
and U1855 (N_1855,In_296,In_122);
and U1856 (N_1856,In_1302,In_1451);
or U1857 (N_1857,In_129,In_1049);
nand U1858 (N_1858,In_1102,In_1310);
nor U1859 (N_1859,In_602,In_878);
and U1860 (N_1860,In_779,In_1402);
nor U1861 (N_1861,In_401,In_1433);
nand U1862 (N_1862,In_683,In_1241);
nand U1863 (N_1863,In_338,In_929);
nand U1864 (N_1864,In_55,In_180);
or U1865 (N_1865,In_1257,In_766);
or U1866 (N_1866,In_618,In_442);
nand U1867 (N_1867,In_541,In_722);
xnor U1868 (N_1868,In_362,In_324);
and U1869 (N_1869,In_252,In_1371);
nor U1870 (N_1870,In_777,In_479);
or U1871 (N_1871,In_1262,In_404);
nand U1872 (N_1872,In_355,In_612);
or U1873 (N_1873,In_471,In_1101);
nor U1874 (N_1874,In_607,In_117);
or U1875 (N_1875,In_1107,In_603);
nor U1876 (N_1876,In_474,In_1478);
xnor U1877 (N_1877,In_1268,In_425);
nor U1878 (N_1878,In_397,In_856);
and U1879 (N_1879,In_542,In_727);
and U1880 (N_1880,In_480,In_840);
and U1881 (N_1881,In_1135,In_681);
nand U1882 (N_1882,In_684,In_1229);
nand U1883 (N_1883,In_151,In_1393);
and U1884 (N_1884,In_177,In_974);
nand U1885 (N_1885,In_509,In_227);
nand U1886 (N_1886,In_605,In_68);
nor U1887 (N_1887,In_124,In_919);
and U1888 (N_1888,In_1262,In_1209);
or U1889 (N_1889,In_27,In_1422);
nand U1890 (N_1890,In_935,In_416);
nor U1891 (N_1891,In_495,In_1306);
and U1892 (N_1892,In_859,In_768);
or U1893 (N_1893,In_338,In_1258);
or U1894 (N_1894,In_106,In_246);
or U1895 (N_1895,In_782,In_364);
or U1896 (N_1896,In_57,In_629);
or U1897 (N_1897,In_538,In_586);
or U1898 (N_1898,In_570,In_1497);
and U1899 (N_1899,In_293,In_193);
nor U1900 (N_1900,In_1026,In_484);
or U1901 (N_1901,In_1001,In_565);
nand U1902 (N_1902,In_1213,In_468);
and U1903 (N_1903,In_516,In_873);
or U1904 (N_1904,In_341,In_222);
and U1905 (N_1905,In_679,In_1096);
or U1906 (N_1906,In_663,In_535);
and U1907 (N_1907,In_432,In_535);
or U1908 (N_1908,In_833,In_1126);
nor U1909 (N_1909,In_933,In_1154);
nand U1910 (N_1910,In_1181,In_122);
nand U1911 (N_1911,In_567,In_712);
nor U1912 (N_1912,In_1414,In_1229);
nor U1913 (N_1913,In_676,In_1333);
nor U1914 (N_1914,In_507,In_906);
nand U1915 (N_1915,In_1413,In_203);
nor U1916 (N_1916,In_284,In_907);
nor U1917 (N_1917,In_433,In_1482);
nor U1918 (N_1918,In_761,In_614);
or U1919 (N_1919,In_740,In_752);
and U1920 (N_1920,In_1199,In_597);
nand U1921 (N_1921,In_2,In_295);
nor U1922 (N_1922,In_583,In_61);
or U1923 (N_1923,In_726,In_650);
nor U1924 (N_1924,In_1273,In_799);
nor U1925 (N_1925,In_1223,In_253);
nor U1926 (N_1926,In_806,In_632);
nand U1927 (N_1927,In_1356,In_462);
or U1928 (N_1928,In_565,In_194);
nand U1929 (N_1929,In_459,In_359);
nand U1930 (N_1930,In_1011,In_866);
or U1931 (N_1931,In_1185,In_1113);
or U1932 (N_1932,In_573,In_505);
nor U1933 (N_1933,In_1326,In_914);
or U1934 (N_1934,In_989,In_1459);
nor U1935 (N_1935,In_1300,In_770);
nand U1936 (N_1936,In_852,In_850);
or U1937 (N_1937,In_1041,In_1154);
nand U1938 (N_1938,In_56,In_316);
or U1939 (N_1939,In_192,In_1478);
nand U1940 (N_1940,In_561,In_726);
or U1941 (N_1941,In_1091,In_1401);
or U1942 (N_1942,In_923,In_909);
nand U1943 (N_1943,In_1191,In_463);
nand U1944 (N_1944,In_324,In_740);
and U1945 (N_1945,In_1254,In_675);
nand U1946 (N_1946,In_269,In_288);
and U1947 (N_1947,In_1062,In_746);
or U1948 (N_1948,In_91,In_551);
or U1949 (N_1949,In_421,In_1480);
or U1950 (N_1950,In_749,In_309);
nand U1951 (N_1951,In_1468,In_41);
nor U1952 (N_1952,In_363,In_889);
and U1953 (N_1953,In_254,In_529);
and U1954 (N_1954,In_1307,In_499);
nor U1955 (N_1955,In_1494,In_1066);
and U1956 (N_1956,In_508,In_506);
nor U1957 (N_1957,In_726,In_140);
or U1958 (N_1958,In_629,In_1104);
or U1959 (N_1959,In_1435,In_1413);
xor U1960 (N_1960,In_1099,In_428);
or U1961 (N_1961,In_80,In_313);
nor U1962 (N_1962,In_591,In_1092);
or U1963 (N_1963,In_850,In_644);
and U1964 (N_1964,In_156,In_1188);
nand U1965 (N_1965,In_905,In_344);
and U1966 (N_1966,In_338,In_359);
or U1967 (N_1967,In_595,In_1467);
and U1968 (N_1968,In_429,In_119);
or U1969 (N_1969,In_917,In_255);
nor U1970 (N_1970,In_1487,In_1156);
or U1971 (N_1971,In_360,In_1490);
and U1972 (N_1972,In_879,In_1119);
nor U1973 (N_1973,In_191,In_1297);
or U1974 (N_1974,In_873,In_685);
or U1975 (N_1975,In_583,In_479);
and U1976 (N_1976,In_203,In_1461);
xnor U1977 (N_1977,In_12,In_1163);
nor U1978 (N_1978,In_1274,In_582);
nand U1979 (N_1979,In_1141,In_976);
nor U1980 (N_1980,In_865,In_236);
and U1981 (N_1981,In_689,In_925);
xor U1982 (N_1982,In_1253,In_302);
nor U1983 (N_1983,In_836,In_37);
and U1984 (N_1984,In_1438,In_456);
and U1985 (N_1985,In_605,In_831);
nand U1986 (N_1986,In_1467,In_685);
or U1987 (N_1987,In_287,In_173);
or U1988 (N_1988,In_1038,In_618);
nand U1989 (N_1989,In_1339,In_1242);
nor U1990 (N_1990,In_192,In_1415);
and U1991 (N_1991,In_718,In_338);
nand U1992 (N_1992,In_270,In_235);
nand U1993 (N_1993,In_361,In_1140);
or U1994 (N_1994,In_1367,In_907);
or U1995 (N_1995,In_360,In_955);
nand U1996 (N_1996,In_380,In_720);
and U1997 (N_1997,In_465,In_778);
or U1998 (N_1998,In_14,In_470);
nand U1999 (N_1999,In_1413,In_392);
or U2000 (N_2000,In_1327,In_445);
nor U2001 (N_2001,In_1192,In_1269);
nor U2002 (N_2002,In_1002,In_1452);
nand U2003 (N_2003,In_973,In_176);
nor U2004 (N_2004,In_483,In_1070);
and U2005 (N_2005,In_795,In_797);
or U2006 (N_2006,In_379,In_1110);
or U2007 (N_2007,In_711,In_946);
and U2008 (N_2008,In_1197,In_198);
nand U2009 (N_2009,In_387,In_608);
and U2010 (N_2010,In_296,In_830);
or U2011 (N_2011,In_777,In_769);
and U2012 (N_2012,In_701,In_741);
nor U2013 (N_2013,In_513,In_1282);
or U2014 (N_2014,In_1336,In_1317);
or U2015 (N_2015,In_1096,In_839);
nor U2016 (N_2016,In_1490,In_101);
and U2017 (N_2017,In_199,In_1288);
nor U2018 (N_2018,In_689,In_146);
and U2019 (N_2019,In_485,In_1430);
nor U2020 (N_2020,In_71,In_1436);
or U2021 (N_2021,In_151,In_842);
or U2022 (N_2022,In_898,In_1251);
xnor U2023 (N_2023,In_372,In_436);
and U2024 (N_2024,In_163,In_755);
nor U2025 (N_2025,In_569,In_967);
or U2026 (N_2026,In_232,In_1486);
or U2027 (N_2027,In_801,In_485);
or U2028 (N_2028,In_778,In_55);
nand U2029 (N_2029,In_673,In_734);
and U2030 (N_2030,In_815,In_1285);
nand U2031 (N_2031,In_875,In_1372);
nor U2032 (N_2032,In_1312,In_1121);
or U2033 (N_2033,In_521,In_342);
and U2034 (N_2034,In_152,In_419);
or U2035 (N_2035,In_1463,In_1445);
or U2036 (N_2036,In_1048,In_613);
and U2037 (N_2037,In_425,In_364);
nor U2038 (N_2038,In_646,In_843);
or U2039 (N_2039,In_755,In_423);
or U2040 (N_2040,In_1085,In_1370);
or U2041 (N_2041,In_1099,In_679);
nor U2042 (N_2042,In_779,In_491);
and U2043 (N_2043,In_21,In_955);
and U2044 (N_2044,In_431,In_1210);
or U2045 (N_2045,In_233,In_1034);
nor U2046 (N_2046,In_109,In_477);
or U2047 (N_2047,In_777,In_78);
nor U2048 (N_2048,In_1339,In_1341);
nand U2049 (N_2049,In_880,In_1274);
and U2050 (N_2050,In_552,In_615);
nor U2051 (N_2051,In_1407,In_1183);
nand U2052 (N_2052,In_590,In_280);
and U2053 (N_2053,In_591,In_995);
nand U2054 (N_2054,In_772,In_501);
and U2055 (N_2055,In_666,In_1122);
and U2056 (N_2056,In_213,In_1081);
nand U2057 (N_2057,In_376,In_205);
nand U2058 (N_2058,In_1043,In_1442);
or U2059 (N_2059,In_1112,In_698);
nand U2060 (N_2060,In_717,In_944);
and U2061 (N_2061,In_870,In_1439);
nor U2062 (N_2062,In_1253,In_136);
or U2063 (N_2063,In_1278,In_1149);
or U2064 (N_2064,In_805,In_1287);
nor U2065 (N_2065,In_1458,In_1385);
and U2066 (N_2066,In_1064,In_282);
or U2067 (N_2067,In_426,In_1252);
nand U2068 (N_2068,In_47,In_625);
nor U2069 (N_2069,In_446,In_795);
nand U2070 (N_2070,In_436,In_784);
nand U2071 (N_2071,In_1447,In_994);
or U2072 (N_2072,In_1327,In_1028);
and U2073 (N_2073,In_1439,In_723);
and U2074 (N_2074,In_75,In_984);
nor U2075 (N_2075,In_1067,In_251);
nand U2076 (N_2076,In_1338,In_1311);
nand U2077 (N_2077,In_1210,In_487);
and U2078 (N_2078,In_1323,In_362);
nor U2079 (N_2079,In_1384,In_1119);
and U2080 (N_2080,In_855,In_1331);
nand U2081 (N_2081,In_6,In_733);
xnor U2082 (N_2082,In_989,In_1182);
or U2083 (N_2083,In_736,In_1331);
nand U2084 (N_2084,In_1142,In_721);
and U2085 (N_2085,In_675,In_987);
or U2086 (N_2086,In_598,In_1195);
nand U2087 (N_2087,In_320,In_512);
and U2088 (N_2088,In_483,In_565);
xor U2089 (N_2089,In_118,In_838);
and U2090 (N_2090,In_1121,In_1182);
nor U2091 (N_2091,In_1172,In_331);
or U2092 (N_2092,In_376,In_653);
or U2093 (N_2093,In_662,In_1179);
or U2094 (N_2094,In_650,In_340);
nor U2095 (N_2095,In_523,In_1194);
nand U2096 (N_2096,In_758,In_1241);
nor U2097 (N_2097,In_807,In_1227);
or U2098 (N_2098,In_57,In_1237);
or U2099 (N_2099,In_771,In_1458);
and U2100 (N_2100,In_794,In_582);
nor U2101 (N_2101,In_1263,In_774);
nand U2102 (N_2102,In_563,In_244);
or U2103 (N_2103,In_1361,In_363);
or U2104 (N_2104,In_653,In_1037);
and U2105 (N_2105,In_1437,In_623);
or U2106 (N_2106,In_134,In_368);
and U2107 (N_2107,In_890,In_89);
or U2108 (N_2108,In_1361,In_1068);
nor U2109 (N_2109,In_1442,In_1021);
nand U2110 (N_2110,In_1374,In_201);
nor U2111 (N_2111,In_595,In_451);
nor U2112 (N_2112,In_603,In_505);
or U2113 (N_2113,In_1133,In_228);
and U2114 (N_2114,In_949,In_738);
and U2115 (N_2115,In_716,In_298);
and U2116 (N_2116,In_508,In_846);
or U2117 (N_2117,In_1438,In_1410);
or U2118 (N_2118,In_38,In_223);
or U2119 (N_2119,In_1021,In_1016);
and U2120 (N_2120,In_798,In_1085);
xnor U2121 (N_2121,In_1352,In_184);
nand U2122 (N_2122,In_1164,In_75);
nor U2123 (N_2123,In_45,In_918);
or U2124 (N_2124,In_472,In_1165);
nand U2125 (N_2125,In_583,In_532);
nand U2126 (N_2126,In_1195,In_838);
or U2127 (N_2127,In_1184,In_1053);
nand U2128 (N_2128,In_1061,In_229);
nand U2129 (N_2129,In_1028,In_1062);
nor U2130 (N_2130,In_790,In_699);
or U2131 (N_2131,In_833,In_1259);
nor U2132 (N_2132,In_581,In_9);
nand U2133 (N_2133,In_867,In_917);
nand U2134 (N_2134,In_1225,In_146);
and U2135 (N_2135,In_1099,In_897);
or U2136 (N_2136,In_1297,In_852);
or U2137 (N_2137,In_1382,In_1287);
and U2138 (N_2138,In_222,In_75);
nor U2139 (N_2139,In_82,In_1212);
and U2140 (N_2140,In_1082,In_1379);
and U2141 (N_2141,In_1307,In_898);
nor U2142 (N_2142,In_467,In_469);
nor U2143 (N_2143,In_26,In_553);
nand U2144 (N_2144,In_1,In_1122);
nor U2145 (N_2145,In_1087,In_1331);
nand U2146 (N_2146,In_427,In_1206);
xnor U2147 (N_2147,In_187,In_1325);
and U2148 (N_2148,In_1308,In_129);
nand U2149 (N_2149,In_136,In_1430);
xor U2150 (N_2150,In_110,In_128);
nor U2151 (N_2151,In_1268,In_30);
nand U2152 (N_2152,In_1122,In_76);
nand U2153 (N_2153,In_503,In_1495);
nor U2154 (N_2154,In_104,In_1093);
nor U2155 (N_2155,In_1312,In_157);
nor U2156 (N_2156,In_87,In_699);
or U2157 (N_2157,In_493,In_1334);
nand U2158 (N_2158,In_801,In_1193);
and U2159 (N_2159,In_935,In_1365);
nand U2160 (N_2160,In_1215,In_817);
or U2161 (N_2161,In_351,In_98);
nand U2162 (N_2162,In_317,In_351);
nor U2163 (N_2163,In_822,In_1182);
and U2164 (N_2164,In_87,In_1140);
or U2165 (N_2165,In_488,In_147);
or U2166 (N_2166,In_425,In_161);
or U2167 (N_2167,In_866,In_826);
nand U2168 (N_2168,In_1494,In_387);
nand U2169 (N_2169,In_887,In_1068);
nand U2170 (N_2170,In_983,In_946);
nand U2171 (N_2171,In_871,In_628);
and U2172 (N_2172,In_1271,In_569);
nor U2173 (N_2173,In_953,In_1380);
nand U2174 (N_2174,In_1243,In_118);
or U2175 (N_2175,In_1348,In_1155);
nor U2176 (N_2176,In_225,In_250);
nand U2177 (N_2177,In_724,In_220);
nor U2178 (N_2178,In_1381,In_942);
and U2179 (N_2179,In_270,In_749);
or U2180 (N_2180,In_300,In_1453);
nand U2181 (N_2181,In_1394,In_308);
and U2182 (N_2182,In_1392,In_169);
nor U2183 (N_2183,In_402,In_766);
or U2184 (N_2184,In_862,In_522);
nand U2185 (N_2185,In_97,In_342);
and U2186 (N_2186,In_20,In_967);
xor U2187 (N_2187,In_307,In_821);
or U2188 (N_2188,In_1446,In_1474);
or U2189 (N_2189,In_701,In_1223);
nor U2190 (N_2190,In_594,In_568);
nand U2191 (N_2191,In_1087,In_51);
and U2192 (N_2192,In_626,In_559);
or U2193 (N_2193,In_713,In_1163);
or U2194 (N_2194,In_1259,In_1218);
nor U2195 (N_2195,In_21,In_1231);
nor U2196 (N_2196,In_88,In_62);
nor U2197 (N_2197,In_610,In_87);
nand U2198 (N_2198,In_419,In_1355);
or U2199 (N_2199,In_477,In_1367);
nor U2200 (N_2200,In_1188,In_1288);
or U2201 (N_2201,In_846,In_1006);
nand U2202 (N_2202,In_289,In_1058);
nor U2203 (N_2203,In_1224,In_1142);
nand U2204 (N_2204,In_654,In_841);
or U2205 (N_2205,In_1269,In_194);
or U2206 (N_2206,In_394,In_429);
and U2207 (N_2207,In_1479,In_49);
or U2208 (N_2208,In_1348,In_1252);
nor U2209 (N_2209,In_249,In_417);
nand U2210 (N_2210,In_475,In_98);
nor U2211 (N_2211,In_1423,In_1005);
nor U2212 (N_2212,In_218,In_657);
and U2213 (N_2213,In_1176,In_550);
and U2214 (N_2214,In_843,In_128);
nand U2215 (N_2215,In_200,In_1145);
nor U2216 (N_2216,In_430,In_42);
and U2217 (N_2217,In_1419,In_1262);
nor U2218 (N_2218,In_990,In_1197);
and U2219 (N_2219,In_1493,In_236);
nor U2220 (N_2220,In_773,In_532);
nor U2221 (N_2221,In_508,In_299);
and U2222 (N_2222,In_463,In_1097);
and U2223 (N_2223,In_297,In_791);
nand U2224 (N_2224,In_1340,In_770);
nand U2225 (N_2225,In_563,In_972);
or U2226 (N_2226,In_159,In_995);
or U2227 (N_2227,In_519,In_1300);
or U2228 (N_2228,In_893,In_594);
nor U2229 (N_2229,In_972,In_500);
and U2230 (N_2230,In_1464,In_1312);
or U2231 (N_2231,In_576,In_48);
or U2232 (N_2232,In_346,In_370);
nor U2233 (N_2233,In_1157,In_1441);
and U2234 (N_2234,In_918,In_705);
nor U2235 (N_2235,In_1229,In_1361);
or U2236 (N_2236,In_636,In_1273);
or U2237 (N_2237,In_813,In_608);
or U2238 (N_2238,In_520,In_67);
and U2239 (N_2239,In_1337,In_307);
nor U2240 (N_2240,In_685,In_989);
and U2241 (N_2241,In_50,In_314);
and U2242 (N_2242,In_192,In_1468);
xnor U2243 (N_2243,In_165,In_673);
and U2244 (N_2244,In_1392,In_1323);
and U2245 (N_2245,In_1461,In_1426);
nor U2246 (N_2246,In_1429,In_917);
and U2247 (N_2247,In_970,In_864);
nor U2248 (N_2248,In_947,In_1445);
and U2249 (N_2249,In_653,In_1056);
and U2250 (N_2250,In_458,In_1311);
nor U2251 (N_2251,In_198,In_1443);
nor U2252 (N_2252,In_4,In_613);
or U2253 (N_2253,In_1107,In_1349);
or U2254 (N_2254,In_1353,In_1371);
and U2255 (N_2255,In_1069,In_783);
xor U2256 (N_2256,In_839,In_1315);
or U2257 (N_2257,In_1164,In_623);
and U2258 (N_2258,In_816,In_513);
nand U2259 (N_2259,In_139,In_616);
or U2260 (N_2260,In_1082,In_1137);
nand U2261 (N_2261,In_569,In_598);
nor U2262 (N_2262,In_1007,In_692);
nand U2263 (N_2263,In_449,In_170);
and U2264 (N_2264,In_1342,In_1035);
and U2265 (N_2265,In_1385,In_437);
nor U2266 (N_2266,In_16,In_1454);
nor U2267 (N_2267,In_79,In_101);
nor U2268 (N_2268,In_1224,In_830);
xor U2269 (N_2269,In_1126,In_439);
nor U2270 (N_2270,In_851,In_1001);
nand U2271 (N_2271,In_987,In_1244);
nor U2272 (N_2272,In_982,In_1078);
nand U2273 (N_2273,In_793,In_780);
nor U2274 (N_2274,In_357,In_1198);
nand U2275 (N_2275,In_361,In_109);
or U2276 (N_2276,In_434,In_627);
or U2277 (N_2277,In_241,In_729);
nand U2278 (N_2278,In_966,In_373);
nand U2279 (N_2279,In_1207,In_1167);
nor U2280 (N_2280,In_1209,In_614);
or U2281 (N_2281,In_129,In_1369);
and U2282 (N_2282,In_1267,In_868);
and U2283 (N_2283,In_1230,In_20);
nand U2284 (N_2284,In_230,In_1323);
or U2285 (N_2285,In_617,In_217);
nand U2286 (N_2286,In_990,In_31);
or U2287 (N_2287,In_395,In_9);
nor U2288 (N_2288,In_1025,In_677);
nor U2289 (N_2289,In_653,In_305);
nand U2290 (N_2290,In_938,In_373);
nor U2291 (N_2291,In_905,In_853);
or U2292 (N_2292,In_851,In_1244);
and U2293 (N_2293,In_856,In_1232);
xnor U2294 (N_2294,In_992,In_754);
and U2295 (N_2295,In_256,In_292);
nor U2296 (N_2296,In_1203,In_1084);
nor U2297 (N_2297,In_265,In_1395);
nand U2298 (N_2298,In_1118,In_219);
nor U2299 (N_2299,In_1261,In_183);
nor U2300 (N_2300,In_854,In_679);
nand U2301 (N_2301,In_1321,In_98);
nand U2302 (N_2302,In_603,In_427);
nor U2303 (N_2303,In_493,In_1118);
or U2304 (N_2304,In_199,In_1276);
nor U2305 (N_2305,In_801,In_1374);
or U2306 (N_2306,In_807,In_612);
nand U2307 (N_2307,In_1066,In_98);
nor U2308 (N_2308,In_932,In_1407);
and U2309 (N_2309,In_861,In_875);
nor U2310 (N_2310,In_1193,In_1407);
and U2311 (N_2311,In_393,In_750);
nand U2312 (N_2312,In_1138,In_196);
or U2313 (N_2313,In_174,In_12);
or U2314 (N_2314,In_1001,In_1498);
nor U2315 (N_2315,In_734,In_701);
or U2316 (N_2316,In_204,In_838);
and U2317 (N_2317,In_1358,In_509);
nand U2318 (N_2318,In_1145,In_616);
nor U2319 (N_2319,In_421,In_687);
or U2320 (N_2320,In_1035,In_537);
nand U2321 (N_2321,In_733,In_811);
nand U2322 (N_2322,In_705,In_1470);
nor U2323 (N_2323,In_700,In_860);
nor U2324 (N_2324,In_789,In_331);
and U2325 (N_2325,In_1447,In_356);
or U2326 (N_2326,In_335,In_789);
or U2327 (N_2327,In_1228,In_3);
nand U2328 (N_2328,In_141,In_563);
and U2329 (N_2329,In_1005,In_1297);
nor U2330 (N_2330,In_604,In_625);
nor U2331 (N_2331,In_190,In_1152);
nor U2332 (N_2332,In_1137,In_1374);
or U2333 (N_2333,In_1075,In_169);
or U2334 (N_2334,In_208,In_1480);
nand U2335 (N_2335,In_1349,In_1252);
nor U2336 (N_2336,In_1,In_335);
or U2337 (N_2337,In_236,In_1013);
or U2338 (N_2338,In_1480,In_291);
and U2339 (N_2339,In_348,In_786);
or U2340 (N_2340,In_118,In_1118);
and U2341 (N_2341,In_386,In_669);
or U2342 (N_2342,In_717,In_658);
nand U2343 (N_2343,In_1400,In_1394);
nand U2344 (N_2344,In_508,In_1329);
nor U2345 (N_2345,In_897,In_745);
and U2346 (N_2346,In_1464,In_1150);
nor U2347 (N_2347,In_931,In_220);
nor U2348 (N_2348,In_916,In_1421);
and U2349 (N_2349,In_1244,In_626);
nand U2350 (N_2350,In_113,In_475);
and U2351 (N_2351,In_1006,In_578);
and U2352 (N_2352,In_960,In_1023);
and U2353 (N_2353,In_26,In_207);
or U2354 (N_2354,In_611,In_300);
xor U2355 (N_2355,In_834,In_1317);
and U2356 (N_2356,In_143,In_667);
nand U2357 (N_2357,In_1481,In_597);
nand U2358 (N_2358,In_1348,In_18);
and U2359 (N_2359,In_949,In_1103);
nand U2360 (N_2360,In_1283,In_117);
and U2361 (N_2361,In_654,In_372);
nand U2362 (N_2362,In_393,In_1181);
or U2363 (N_2363,In_756,In_644);
nor U2364 (N_2364,In_955,In_786);
nor U2365 (N_2365,In_657,In_1341);
nand U2366 (N_2366,In_1438,In_1021);
nor U2367 (N_2367,In_144,In_1282);
and U2368 (N_2368,In_412,In_95);
nand U2369 (N_2369,In_458,In_1145);
and U2370 (N_2370,In_45,In_681);
nand U2371 (N_2371,In_820,In_643);
nor U2372 (N_2372,In_72,In_393);
or U2373 (N_2373,In_740,In_144);
or U2374 (N_2374,In_300,In_1126);
nor U2375 (N_2375,In_95,In_1054);
nand U2376 (N_2376,In_89,In_1139);
or U2377 (N_2377,In_969,In_1121);
nand U2378 (N_2378,In_1465,In_951);
nand U2379 (N_2379,In_440,In_78);
and U2380 (N_2380,In_164,In_309);
and U2381 (N_2381,In_36,In_1192);
nand U2382 (N_2382,In_539,In_999);
nand U2383 (N_2383,In_578,In_889);
xnor U2384 (N_2384,In_1064,In_1089);
and U2385 (N_2385,In_798,In_799);
and U2386 (N_2386,In_227,In_1054);
or U2387 (N_2387,In_1254,In_641);
nand U2388 (N_2388,In_1018,In_1271);
nor U2389 (N_2389,In_949,In_331);
nor U2390 (N_2390,In_15,In_1371);
xor U2391 (N_2391,In_189,In_166);
or U2392 (N_2392,In_1207,In_1071);
or U2393 (N_2393,In_1478,In_636);
nor U2394 (N_2394,In_1320,In_1256);
nand U2395 (N_2395,In_744,In_110);
or U2396 (N_2396,In_67,In_1393);
nor U2397 (N_2397,In_405,In_563);
nor U2398 (N_2398,In_365,In_911);
and U2399 (N_2399,In_1351,In_599);
or U2400 (N_2400,In_1019,In_191);
and U2401 (N_2401,In_819,In_1101);
and U2402 (N_2402,In_241,In_250);
nand U2403 (N_2403,In_1191,In_415);
nor U2404 (N_2404,In_122,In_1253);
or U2405 (N_2405,In_742,In_267);
nor U2406 (N_2406,In_904,In_334);
or U2407 (N_2407,In_417,In_361);
nand U2408 (N_2408,In_540,In_1107);
nor U2409 (N_2409,In_725,In_672);
nor U2410 (N_2410,In_1077,In_105);
nor U2411 (N_2411,In_36,In_1288);
nand U2412 (N_2412,In_1221,In_1002);
xor U2413 (N_2413,In_268,In_1281);
nor U2414 (N_2414,In_738,In_5);
or U2415 (N_2415,In_1188,In_952);
nand U2416 (N_2416,In_1302,In_1288);
or U2417 (N_2417,In_738,In_1108);
and U2418 (N_2418,In_503,In_110);
and U2419 (N_2419,In_161,In_25);
and U2420 (N_2420,In_596,In_1058);
nand U2421 (N_2421,In_1234,In_891);
and U2422 (N_2422,In_1190,In_1192);
or U2423 (N_2423,In_248,In_590);
or U2424 (N_2424,In_99,In_180);
or U2425 (N_2425,In_1436,In_561);
xor U2426 (N_2426,In_609,In_1486);
nand U2427 (N_2427,In_1059,In_44);
or U2428 (N_2428,In_905,In_1091);
or U2429 (N_2429,In_1252,In_562);
or U2430 (N_2430,In_706,In_1388);
and U2431 (N_2431,In_577,In_783);
or U2432 (N_2432,In_365,In_840);
or U2433 (N_2433,In_462,In_326);
or U2434 (N_2434,In_51,In_1073);
nor U2435 (N_2435,In_1169,In_1297);
or U2436 (N_2436,In_574,In_99);
and U2437 (N_2437,In_1328,In_1013);
nor U2438 (N_2438,In_491,In_380);
or U2439 (N_2439,In_263,In_1291);
or U2440 (N_2440,In_202,In_1262);
nand U2441 (N_2441,In_1061,In_402);
or U2442 (N_2442,In_578,In_1148);
nor U2443 (N_2443,In_239,In_978);
or U2444 (N_2444,In_4,In_202);
or U2445 (N_2445,In_554,In_914);
or U2446 (N_2446,In_359,In_296);
nand U2447 (N_2447,In_469,In_1173);
nor U2448 (N_2448,In_1303,In_333);
nand U2449 (N_2449,In_951,In_947);
or U2450 (N_2450,In_1002,In_586);
or U2451 (N_2451,In_1496,In_183);
and U2452 (N_2452,In_1282,In_199);
nand U2453 (N_2453,In_29,In_976);
nand U2454 (N_2454,In_621,In_1303);
nand U2455 (N_2455,In_322,In_463);
and U2456 (N_2456,In_29,In_1357);
xnor U2457 (N_2457,In_1318,In_838);
xnor U2458 (N_2458,In_882,In_911);
nand U2459 (N_2459,In_137,In_828);
and U2460 (N_2460,In_127,In_210);
and U2461 (N_2461,In_60,In_1016);
nor U2462 (N_2462,In_1392,In_1411);
nor U2463 (N_2463,In_634,In_1332);
nand U2464 (N_2464,In_469,In_622);
or U2465 (N_2465,In_1432,In_703);
nand U2466 (N_2466,In_650,In_1368);
nor U2467 (N_2467,In_369,In_814);
or U2468 (N_2468,In_306,In_1420);
nand U2469 (N_2469,In_79,In_1263);
nand U2470 (N_2470,In_974,In_1350);
or U2471 (N_2471,In_427,In_542);
and U2472 (N_2472,In_1113,In_1184);
and U2473 (N_2473,In_73,In_1182);
nor U2474 (N_2474,In_473,In_126);
or U2475 (N_2475,In_90,In_1113);
nor U2476 (N_2476,In_1304,In_1322);
or U2477 (N_2477,In_926,In_1325);
and U2478 (N_2478,In_1048,In_267);
nor U2479 (N_2479,In_1383,In_1220);
nor U2480 (N_2480,In_1108,In_497);
nand U2481 (N_2481,In_1186,In_95);
or U2482 (N_2482,In_1269,In_819);
and U2483 (N_2483,In_382,In_491);
nor U2484 (N_2484,In_10,In_643);
xnor U2485 (N_2485,In_1459,In_235);
nor U2486 (N_2486,In_877,In_503);
xor U2487 (N_2487,In_607,In_1371);
or U2488 (N_2488,In_1253,In_327);
nor U2489 (N_2489,In_934,In_6);
nand U2490 (N_2490,In_77,In_283);
nor U2491 (N_2491,In_729,In_1452);
nor U2492 (N_2492,In_748,In_93);
nand U2493 (N_2493,In_1484,In_925);
or U2494 (N_2494,In_1170,In_3);
and U2495 (N_2495,In_714,In_1059);
nand U2496 (N_2496,In_1154,In_1478);
nand U2497 (N_2497,In_704,In_888);
and U2498 (N_2498,In_497,In_771);
nand U2499 (N_2499,In_755,In_140);
or U2500 (N_2500,In_325,In_357);
or U2501 (N_2501,In_278,In_533);
nor U2502 (N_2502,In_1456,In_1439);
and U2503 (N_2503,In_98,In_1128);
and U2504 (N_2504,In_311,In_1176);
or U2505 (N_2505,In_889,In_1468);
and U2506 (N_2506,In_1331,In_1069);
nor U2507 (N_2507,In_939,In_823);
and U2508 (N_2508,In_820,In_783);
nand U2509 (N_2509,In_905,In_1474);
or U2510 (N_2510,In_1227,In_52);
and U2511 (N_2511,In_733,In_114);
nand U2512 (N_2512,In_1130,In_649);
nand U2513 (N_2513,In_723,In_829);
or U2514 (N_2514,In_639,In_262);
nor U2515 (N_2515,In_766,In_318);
and U2516 (N_2516,In_545,In_89);
or U2517 (N_2517,In_1321,In_22);
nor U2518 (N_2518,In_632,In_1258);
or U2519 (N_2519,In_482,In_262);
or U2520 (N_2520,In_927,In_333);
and U2521 (N_2521,In_535,In_1311);
xnor U2522 (N_2522,In_395,In_1035);
or U2523 (N_2523,In_804,In_1154);
nor U2524 (N_2524,In_1054,In_120);
or U2525 (N_2525,In_133,In_952);
nor U2526 (N_2526,In_492,In_689);
nor U2527 (N_2527,In_1028,In_515);
nand U2528 (N_2528,In_391,In_660);
or U2529 (N_2529,In_327,In_196);
or U2530 (N_2530,In_13,In_72);
or U2531 (N_2531,In_759,In_854);
nor U2532 (N_2532,In_307,In_1106);
nand U2533 (N_2533,In_775,In_791);
and U2534 (N_2534,In_546,In_921);
nand U2535 (N_2535,In_90,In_391);
nor U2536 (N_2536,In_1175,In_802);
nor U2537 (N_2537,In_164,In_1436);
nor U2538 (N_2538,In_798,In_1369);
or U2539 (N_2539,In_1350,In_548);
nor U2540 (N_2540,In_485,In_1379);
xor U2541 (N_2541,In_373,In_1004);
xnor U2542 (N_2542,In_1039,In_322);
and U2543 (N_2543,In_1041,In_149);
or U2544 (N_2544,In_389,In_1251);
and U2545 (N_2545,In_728,In_1479);
or U2546 (N_2546,In_1403,In_695);
nand U2547 (N_2547,In_1244,In_1324);
and U2548 (N_2548,In_329,In_1363);
nor U2549 (N_2549,In_1180,In_8);
and U2550 (N_2550,In_244,In_1308);
nand U2551 (N_2551,In_1072,In_515);
and U2552 (N_2552,In_713,In_250);
and U2553 (N_2553,In_669,In_857);
nand U2554 (N_2554,In_1408,In_798);
and U2555 (N_2555,In_357,In_713);
or U2556 (N_2556,In_1271,In_606);
nand U2557 (N_2557,In_832,In_1046);
and U2558 (N_2558,In_1258,In_1177);
nor U2559 (N_2559,In_580,In_1366);
nor U2560 (N_2560,In_892,In_1295);
or U2561 (N_2561,In_123,In_875);
nor U2562 (N_2562,In_288,In_676);
nand U2563 (N_2563,In_199,In_518);
and U2564 (N_2564,In_794,In_697);
nand U2565 (N_2565,In_916,In_1443);
or U2566 (N_2566,In_381,In_1053);
and U2567 (N_2567,In_1382,In_764);
nand U2568 (N_2568,In_1079,In_320);
or U2569 (N_2569,In_453,In_780);
nor U2570 (N_2570,In_226,In_1445);
nand U2571 (N_2571,In_847,In_694);
and U2572 (N_2572,In_611,In_1094);
or U2573 (N_2573,In_1010,In_313);
and U2574 (N_2574,In_559,In_229);
nor U2575 (N_2575,In_701,In_1370);
nor U2576 (N_2576,In_262,In_313);
nand U2577 (N_2577,In_454,In_1039);
nor U2578 (N_2578,In_21,In_954);
and U2579 (N_2579,In_1015,In_782);
or U2580 (N_2580,In_1032,In_1212);
and U2581 (N_2581,In_465,In_1274);
and U2582 (N_2582,In_1213,In_1123);
nor U2583 (N_2583,In_445,In_1170);
nor U2584 (N_2584,In_169,In_1070);
nor U2585 (N_2585,In_83,In_30);
nor U2586 (N_2586,In_1117,In_1091);
nand U2587 (N_2587,In_866,In_634);
nand U2588 (N_2588,In_178,In_1169);
or U2589 (N_2589,In_75,In_1367);
nand U2590 (N_2590,In_703,In_552);
or U2591 (N_2591,In_546,In_764);
and U2592 (N_2592,In_1124,In_1028);
nand U2593 (N_2593,In_1233,In_1317);
nor U2594 (N_2594,In_650,In_1128);
nor U2595 (N_2595,In_387,In_569);
nand U2596 (N_2596,In_821,In_1416);
nor U2597 (N_2597,In_542,In_338);
and U2598 (N_2598,In_26,In_719);
nand U2599 (N_2599,In_207,In_599);
and U2600 (N_2600,In_548,In_1482);
and U2601 (N_2601,In_200,In_1430);
nor U2602 (N_2602,In_425,In_588);
nand U2603 (N_2603,In_908,In_1037);
nor U2604 (N_2604,In_585,In_635);
or U2605 (N_2605,In_1294,In_929);
and U2606 (N_2606,In_699,In_777);
nor U2607 (N_2607,In_832,In_495);
nand U2608 (N_2608,In_366,In_1273);
and U2609 (N_2609,In_950,In_576);
or U2610 (N_2610,In_635,In_1018);
and U2611 (N_2611,In_220,In_325);
xnor U2612 (N_2612,In_1447,In_251);
or U2613 (N_2613,In_1340,In_312);
or U2614 (N_2614,In_1141,In_1234);
nand U2615 (N_2615,In_1194,In_1292);
nand U2616 (N_2616,In_468,In_45);
xnor U2617 (N_2617,In_964,In_872);
and U2618 (N_2618,In_1178,In_1408);
and U2619 (N_2619,In_316,In_718);
nand U2620 (N_2620,In_960,In_115);
and U2621 (N_2621,In_642,In_793);
xor U2622 (N_2622,In_1359,In_38);
xnor U2623 (N_2623,In_1393,In_159);
nand U2624 (N_2624,In_1339,In_318);
nor U2625 (N_2625,In_724,In_149);
nand U2626 (N_2626,In_1397,In_787);
nor U2627 (N_2627,In_397,In_1274);
or U2628 (N_2628,In_451,In_635);
or U2629 (N_2629,In_212,In_205);
or U2630 (N_2630,In_184,In_501);
and U2631 (N_2631,In_1203,In_1343);
nand U2632 (N_2632,In_593,In_490);
nor U2633 (N_2633,In_1497,In_368);
nand U2634 (N_2634,In_1061,In_931);
nor U2635 (N_2635,In_1112,In_129);
nor U2636 (N_2636,In_956,In_154);
and U2637 (N_2637,In_791,In_1479);
nor U2638 (N_2638,In_851,In_594);
or U2639 (N_2639,In_965,In_670);
nand U2640 (N_2640,In_437,In_793);
nor U2641 (N_2641,In_133,In_957);
nor U2642 (N_2642,In_52,In_286);
nand U2643 (N_2643,In_1042,In_1453);
nand U2644 (N_2644,In_1134,In_817);
or U2645 (N_2645,In_905,In_1235);
nor U2646 (N_2646,In_1463,In_1315);
or U2647 (N_2647,In_151,In_1467);
nor U2648 (N_2648,In_1213,In_1357);
nor U2649 (N_2649,In_1349,In_380);
nand U2650 (N_2650,In_236,In_717);
and U2651 (N_2651,In_258,In_544);
nand U2652 (N_2652,In_929,In_475);
nand U2653 (N_2653,In_357,In_491);
nand U2654 (N_2654,In_199,In_461);
or U2655 (N_2655,In_346,In_492);
or U2656 (N_2656,In_370,In_1089);
and U2657 (N_2657,In_870,In_886);
xor U2658 (N_2658,In_1133,In_231);
or U2659 (N_2659,In_1454,In_1274);
nor U2660 (N_2660,In_748,In_659);
nor U2661 (N_2661,In_32,In_803);
nand U2662 (N_2662,In_328,In_348);
nand U2663 (N_2663,In_1455,In_1013);
nand U2664 (N_2664,In_570,In_247);
nor U2665 (N_2665,In_676,In_383);
and U2666 (N_2666,In_284,In_393);
and U2667 (N_2667,In_1113,In_716);
or U2668 (N_2668,In_531,In_126);
or U2669 (N_2669,In_1188,In_202);
or U2670 (N_2670,In_938,In_936);
nand U2671 (N_2671,In_562,In_95);
nand U2672 (N_2672,In_1124,In_1316);
nand U2673 (N_2673,In_639,In_1404);
nand U2674 (N_2674,In_129,In_1341);
and U2675 (N_2675,In_636,In_722);
or U2676 (N_2676,In_953,In_482);
or U2677 (N_2677,In_902,In_1436);
and U2678 (N_2678,In_258,In_916);
nor U2679 (N_2679,In_236,In_1133);
or U2680 (N_2680,In_988,In_823);
nand U2681 (N_2681,In_872,In_734);
nand U2682 (N_2682,In_713,In_222);
xnor U2683 (N_2683,In_334,In_338);
and U2684 (N_2684,In_659,In_105);
nor U2685 (N_2685,In_196,In_634);
nor U2686 (N_2686,In_305,In_287);
nor U2687 (N_2687,In_914,In_536);
nor U2688 (N_2688,In_1170,In_39);
and U2689 (N_2689,In_75,In_1227);
or U2690 (N_2690,In_618,In_498);
and U2691 (N_2691,In_872,In_647);
or U2692 (N_2692,In_971,In_183);
and U2693 (N_2693,In_479,In_336);
and U2694 (N_2694,In_500,In_332);
nand U2695 (N_2695,In_1259,In_637);
nor U2696 (N_2696,In_598,In_377);
xor U2697 (N_2697,In_115,In_119);
and U2698 (N_2698,In_399,In_431);
and U2699 (N_2699,In_272,In_1199);
and U2700 (N_2700,In_443,In_403);
and U2701 (N_2701,In_1477,In_1411);
nand U2702 (N_2702,In_302,In_1026);
nand U2703 (N_2703,In_845,In_388);
and U2704 (N_2704,In_51,In_1313);
or U2705 (N_2705,In_1280,In_1274);
and U2706 (N_2706,In_1358,In_686);
and U2707 (N_2707,In_500,In_1172);
nand U2708 (N_2708,In_1287,In_1334);
nand U2709 (N_2709,In_183,In_714);
or U2710 (N_2710,In_289,In_318);
nand U2711 (N_2711,In_1160,In_338);
and U2712 (N_2712,In_659,In_1061);
nand U2713 (N_2713,In_418,In_920);
or U2714 (N_2714,In_397,In_1453);
nor U2715 (N_2715,In_949,In_642);
nor U2716 (N_2716,In_158,In_481);
nor U2717 (N_2717,In_183,In_999);
or U2718 (N_2718,In_720,In_12);
or U2719 (N_2719,In_159,In_1194);
nor U2720 (N_2720,In_256,In_1241);
nand U2721 (N_2721,In_561,In_1151);
and U2722 (N_2722,In_1348,In_1246);
and U2723 (N_2723,In_1015,In_874);
nor U2724 (N_2724,In_1178,In_92);
and U2725 (N_2725,In_870,In_977);
xnor U2726 (N_2726,In_707,In_670);
nand U2727 (N_2727,In_779,In_1418);
nand U2728 (N_2728,In_1174,In_701);
nor U2729 (N_2729,In_519,In_171);
nand U2730 (N_2730,In_591,In_3);
nand U2731 (N_2731,In_1430,In_666);
and U2732 (N_2732,In_1288,In_176);
nand U2733 (N_2733,In_1223,In_1091);
nand U2734 (N_2734,In_1054,In_1097);
nand U2735 (N_2735,In_290,In_1297);
xor U2736 (N_2736,In_1281,In_799);
and U2737 (N_2737,In_880,In_9);
and U2738 (N_2738,In_472,In_330);
and U2739 (N_2739,In_485,In_121);
and U2740 (N_2740,In_494,In_805);
nor U2741 (N_2741,In_1187,In_1004);
nor U2742 (N_2742,In_1235,In_1481);
and U2743 (N_2743,In_1077,In_1122);
nor U2744 (N_2744,In_269,In_921);
nand U2745 (N_2745,In_237,In_1424);
xor U2746 (N_2746,In_1044,In_684);
and U2747 (N_2747,In_826,In_197);
xor U2748 (N_2748,In_36,In_1411);
and U2749 (N_2749,In_375,In_1388);
and U2750 (N_2750,In_242,In_129);
nand U2751 (N_2751,In_1385,In_95);
and U2752 (N_2752,In_702,In_959);
nand U2753 (N_2753,In_1179,In_1268);
nand U2754 (N_2754,In_413,In_496);
nor U2755 (N_2755,In_1014,In_422);
nand U2756 (N_2756,In_800,In_1453);
or U2757 (N_2757,In_358,In_413);
nor U2758 (N_2758,In_1383,In_6);
or U2759 (N_2759,In_305,In_547);
or U2760 (N_2760,In_296,In_433);
nand U2761 (N_2761,In_522,In_411);
nor U2762 (N_2762,In_834,In_318);
xor U2763 (N_2763,In_1228,In_1450);
and U2764 (N_2764,In_90,In_1126);
and U2765 (N_2765,In_288,In_1018);
or U2766 (N_2766,In_1137,In_337);
nor U2767 (N_2767,In_1237,In_260);
nand U2768 (N_2768,In_999,In_973);
nor U2769 (N_2769,In_1120,In_740);
or U2770 (N_2770,In_1425,In_955);
nand U2771 (N_2771,In_113,In_682);
or U2772 (N_2772,In_772,In_1454);
nand U2773 (N_2773,In_158,In_323);
nand U2774 (N_2774,In_1291,In_1158);
nand U2775 (N_2775,In_617,In_1183);
and U2776 (N_2776,In_1123,In_330);
nand U2777 (N_2777,In_675,In_978);
nand U2778 (N_2778,In_176,In_790);
nor U2779 (N_2779,In_436,In_1463);
or U2780 (N_2780,In_572,In_845);
and U2781 (N_2781,In_86,In_870);
nor U2782 (N_2782,In_1475,In_1215);
nand U2783 (N_2783,In_340,In_1202);
and U2784 (N_2784,In_1402,In_411);
or U2785 (N_2785,In_890,In_1159);
nand U2786 (N_2786,In_1313,In_571);
and U2787 (N_2787,In_1020,In_305);
and U2788 (N_2788,In_291,In_549);
nor U2789 (N_2789,In_1272,In_1261);
or U2790 (N_2790,In_1198,In_460);
nor U2791 (N_2791,In_752,In_252);
nor U2792 (N_2792,In_1062,In_391);
or U2793 (N_2793,In_1013,In_994);
nor U2794 (N_2794,In_1485,In_48);
nand U2795 (N_2795,In_707,In_773);
nand U2796 (N_2796,In_712,In_834);
nor U2797 (N_2797,In_396,In_765);
and U2798 (N_2798,In_956,In_359);
nor U2799 (N_2799,In_356,In_114);
nand U2800 (N_2800,In_425,In_1001);
and U2801 (N_2801,In_36,In_1086);
and U2802 (N_2802,In_704,In_1194);
and U2803 (N_2803,In_14,In_844);
and U2804 (N_2804,In_1287,In_1121);
nand U2805 (N_2805,In_37,In_481);
nor U2806 (N_2806,In_1400,In_1033);
or U2807 (N_2807,In_575,In_890);
or U2808 (N_2808,In_253,In_220);
or U2809 (N_2809,In_380,In_1092);
xor U2810 (N_2810,In_201,In_993);
nand U2811 (N_2811,In_380,In_691);
nand U2812 (N_2812,In_103,In_765);
nand U2813 (N_2813,In_42,In_9);
or U2814 (N_2814,In_579,In_957);
nor U2815 (N_2815,In_510,In_405);
xnor U2816 (N_2816,In_361,In_934);
or U2817 (N_2817,In_972,In_364);
nor U2818 (N_2818,In_1064,In_773);
or U2819 (N_2819,In_987,In_349);
nand U2820 (N_2820,In_485,In_1417);
or U2821 (N_2821,In_1062,In_134);
and U2822 (N_2822,In_663,In_163);
and U2823 (N_2823,In_1415,In_8);
nand U2824 (N_2824,In_685,In_13);
nand U2825 (N_2825,In_180,In_1162);
nor U2826 (N_2826,In_226,In_1493);
or U2827 (N_2827,In_1199,In_914);
xor U2828 (N_2828,In_1217,In_866);
and U2829 (N_2829,In_1446,In_459);
nand U2830 (N_2830,In_1415,In_667);
or U2831 (N_2831,In_1276,In_846);
and U2832 (N_2832,In_1077,In_496);
nand U2833 (N_2833,In_1128,In_496);
nand U2834 (N_2834,In_214,In_458);
nor U2835 (N_2835,In_787,In_174);
or U2836 (N_2836,In_869,In_425);
or U2837 (N_2837,In_58,In_549);
and U2838 (N_2838,In_308,In_25);
nand U2839 (N_2839,In_345,In_1315);
and U2840 (N_2840,In_1282,In_1192);
nor U2841 (N_2841,In_1309,In_468);
and U2842 (N_2842,In_1012,In_922);
nor U2843 (N_2843,In_897,In_347);
or U2844 (N_2844,In_42,In_1498);
nand U2845 (N_2845,In_523,In_716);
or U2846 (N_2846,In_119,In_1452);
and U2847 (N_2847,In_1126,In_1085);
and U2848 (N_2848,In_1443,In_1081);
or U2849 (N_2849,In_893,In_401);
nand U2850 (N_2850,In_18,In_922);
nor U2851 (N_2851,In_1000,In_1160);
nand U2852 (N_2852,In_1408,In_527);
nand U2853 (N_2853,In_817,In_576);
or U2854 (N_2854,In_1411,In_444);
or U2855 (N_2855,In_521,In_619);
and U2856 (N_2856,In_658,In_125);
and U2857 (N_2857,In_1299,In_1210);
nor U2858 (N_2858,In_659,In_277);
or U2859 (N_2859,In_1465,In_877);
nand U2860 (N_2860,In_288,In_794);
or U2861 (N_2861,In_956,In_725);
and U2862 (N_2862,In_1336,In_79);
and U2863 (N_2863,In_903,In_266);
or U2864 (N_2864,In_1308,In_1191);
nor U2865 (N_2865,In_275,In_535);
nor U2866 (N_2866,In_197,In_519);
nor U2867 (N_2867,In_1390,In_94);
and U2868 (N_2868,In_143,In_596);
nor U2869 (N_2869,In_733,In_1225);
and U2870 (N_2870,In_696,In_413);
nor U2871 (N_2871,In_1356,In_1284);
or U2872 (N_2872,In_241,In_293);
or U2873 (N_2873,In_653,In_221);
nor U2874 (N_2874,In_423,In_636);
nor U2875 (N_2875,In_1243,In_1283);
nand U2876 (N_2876,In_40,In_801);
nor U2877 (N_2877,In_548,In_601);
nand U2878 (N_2878,In_1202,In_1173);
and U2879 (N_2879,In_413,In_574);
xnor U2880 (N_2880,In_633,In_1086);
or U2881 (N_2881,In_171,In_708);
or U2882 (N_2882,In_649,In_263);
or U2883 (N_2883,In_838,In_949);
nand U2884 (N_2884,In_1375,In_559);
and U2885 (N_2885,In_951,In_246);
or U2886 (N_2886,In_352,In_299);
or U2887 (N_2887,In_1064,In_39);
or U2888 (N_2888,In_713,In_1111);
nor U2889 (N_2889,In_425,In_1426);
nor U2890 (N_2890,In_1055,In_1258);
or U2891 (N_2891,In_109,In_1318);
nor U2892 (N_2892,In_33,In_564);
or U2893 (N_2893,In_757,In_1342);
nand U2894 (N_2894,In_624,In_1445);
or U2895 (N_2895,In_634,In_487);
or U2896 (N_2896,In_1022,In_554);
nor U2897 (N_2897,In_540,In_1315);
nor U2898 (N_2898,In_561,In_95);
and U2899 (N_2899,In_1364,In_800);
nand U2900 (N_2900,In_774,In_1325);
and U2901 (N_2901,In_207,In_1273);
nand U2902 (N_2902,In_785,In_1456);
and U2903 (N_2903,In_638,In_1378);
xnor U2904 (N_2904,In_303,In_1065);
or U2905 (N_2905,In_1405,In_1312);
and U2906 (N_2906,In_1011,In_1380);
nor U2907 (N_2907,In_972,In_324);
or U2908 (N_2908,In_1274,In_50);
nand U2909 (N_2909,In_743,In_234);
and U2910 (N_2910,In_170,In_960);
nand U2911 (N_2911,In_638,In_1438);
xor U2912 (N_2912,In_1179,In_223);
or U2913 (N_2913,In_1482,In_811);
or U2914 (N_2914,In_645,In_22);
nor U2915 (N_2915,In_485,In_1163);
nand U2916 (N_2916,In_440,In_368);
and U2917 (N_2917,In_1361,In_563);
or U2918 (N_2918,In_1252,In_392);
or U2919 (N_2919,In_1370,In_1129);
and U2920 (N_2920,In_3,In_927);
and U2921 (N_2921,In_707,In_370);
and U2922 (N_2922,In_247,In_524);
nand U2923 (N_2923,In_1319,In_77);
or U2924 (N_2924,In_922,In_1457);
and U2925 (N_2925,In_1142,In_557);
and U2926 (N_2926,In_411,In_611);
nor U2927 (N_2927,In_318,In_650);
or U2928 (N_2928,In_229,In_867);
nand U2929 (N_2929,In_1166,In_1077);
or U2930 (N_2930,In_72,In_578);
or U2931 (N_2931,In_1479,In_1465);
nand U2932 (N_2932,In_896,In_995);
nor U2933 (N_2933,In_1236,In_1266);
or U2934 (N_2934,In_979,In_657);
or U2935 (N_2935,In_1488,In_801);
nor U2936 (N_2936,In_229,In_1188);
nor U2937 (N_2937,In_173,In_516);
nor U2938 (N_2938,In_682,In_908);
and U2939 (N_2939,In_425,In_1300);
and U2940 (N_2940,In_244,In_443);
nand U2941 (N_2941,In_714,In_562);
or U2942 (N_2942,In_355,In_1032);
nand U2943 (N_2943,In_1048,In_1010);
or U2944 (N_2944,In_473,In_1069);
nand U2945 (N_2945,In_1174,In_462);
or U2946 (N_2946,In_88,In_574);
or U2947 (N_2947,In_1400,In_12);
nand U2948 (N_2948,In_1257,In_547);
and U2949 (N_2949,In_855,In_1192);
nand U2950 (N_2950,In_299,In_1027);
or U2951 (N_2951,In_3,In_954);
nor U2952 (N_2952,In_702,In_214);
nor U2953 (N_2953,In_1339,In_600);
nor U2954 (N_2954,In_683,In_111);
and U2955 (N_2955,In_399,In_1253);
or U2956 (N_2956,In_1236,In_353);
nor U2957 (N_2957,In_1384,In_268);
or U2958 (N_2958,In_135,In_656);
or U2959 (N_2959,In_107,In_1441);
nor U2960 (N_2960,In_609,In_485);
and U2961 (N_2961,In_625,In_613);
nor U2962 (N_2962,In_80,In_542);
or U2963 (N_2963,In_449,In_1495);
and U2964 (N_2964,In_206,In_330);
or U2965 (N_2965,In_1347,In_624);
nor U2966 (N_2966,In_1041,In_812);
nor U2967 (N_2967,In_908,In_270);
nand U2968 (N_2968,In_1329,In_378);
or U2969 (N_2969,In_209,In_469);
nor U2970 (N_2970,In_1314,In_611);
or U2971 (N_2971,In_1429,In_1225);
or U2972 (N_2972,In_1398,In_1453);
nor U2973 (N_2973,In_247,In_1238);
nand U2974 (N_2974,In_1298,In_24);
and U2975 (N_2975,In_1472,In_538);
or U2976 (N_2976,In_248,In_252);
and U2977 (N_2977,In_647,In_817);
nor U2978 (N_2978,In_700,In_1318);
or U2979 (N_2979,In_325,In_884);
nor U2980 (N_2980,In_1415,In_386);
nand U2981 (N_2981,In_596,In_417);
nor U2982 (N_2982,In_738,In_1375);
and U2983 (N_2983,In_139,In_1174);
nor U2984 (N_2984,In_398,In_1126);
or U2985 (N_2985,In_1083,In_976);
nand U2986 (N_2986,In_952,In_269);
or U2987 (N_2987,In_299,In_1226);
and U2988 (N_2988,In_1359,In_273);
nor U2989 (N_2989,In_947,In_264);
or U2990 (N_2990,In_794,In_594);
and U2991 (N_2991,In_218,In_314);
nor U2992 (N_2992,In_601,In_1254);
and U2993 (N_2993,In_470,In_360);
nor U2994 (N_2994,In_1424,In_1380);
nand U2995 (N_2995,In_276,In_231);
nand U2996 (N_2996,In_413,In_26);
and U2997 (N_2997,In_263,In_239);
nor U2998 (N_2998,In_1457,In_1171);
or U2999 (N_2999,In_337,In_570);
nand U3000 (N_3000,N_670,N_736);
nand U3001 (N_3001,N_2139,N_2539);
and U3002 (N_3002,N_1908,N_1168);
nor U3003 (N_3003,N_50,N_1712);
nand U3004 (N_3004,N_744,N_1213);
or U3005 (N_3005,N_133,N_415);
or U3006 (N_3006,N_709,N_363);
nand U3007 (N_3007,N_2870,N_353);
or U3008 (N_3008,N_1534,N_1063);
and U3009 (N_3009,N_1246,N_2512);
or U3010 (N_3010,N_494,N_2902);
and U3011 (N_3011,N_636,N_889);
nand U3012 (N_3012,N_137,N_90);
or U3013 (N_3013,N_2538,N_1957);
nand U3014 (N_3014,N_1748,N_1634);
and U3015 (N_3015,N_796,N_2829);
and U3016 (N_3016,N_210,N_2848);
nand U3017 (N_3017,N_354,N_1357);
nand U3018 (N_3018,N_109,N_2570);
nor U3019 (N_3019,N_2561,N_2391);
nor U3020 (N_3020,N_1121,N_1846);
or U3021 (N_3021,N_2238,N_1726);
nand U3022 (N_3022,N_2114,N_706);
nand U3023 (N_3023,N_1149,N_1385);
or U3024 (N_3024,N_2579,N_1216);
and U3025 (N_3025,N_1010,N_162);
and U3026 (N_3026,N_1513,N_1218);
and U3027 (N_3027,N_2367,N_387);
nor U3028 (N_3028,N_1612,N_2595);
nand U3029 (N_3029,N_1450,N_1483);
or U3030 (N_3030,N_521,N_682);
or U3031 (N_3031,N_2261,N_1166);
nand U3032 (N_3032,N_1599,N_1167);
or U3033 (N_3033,N_1834,N_2287);
nand U3034 (N_3034,N_952,N_729);
and U3035 (N_3035,N_1425,N_1332);
nor U3036 (N_3036,N_2953,N_569);
nor U3037 (N_3037,N_452,N_245);
and U3038 (N_3038,N_1873,N_761);
and U3039 (N_3039,N_2656,N_1485);
and U3040 (N_3040,N_346,N_1869);
and U3041 (N_3041,N_1369,N_1864);
nor U3042 (N_3042,N_1071,N_1894);
nor U3043 (N_3043,N_2423,N_1404);
nand U3044 (N_3044,N_2153,N_1630);
nor U3045 (N_3045,N_1274,N_170);
or U3046 (N_3046,N_1230,N_2523);
nor U3047 (N_3047,N_1878,N_142);
or U3048 (N_3048,N_823,N_983);
nor U3049 (N_3049,N_2294,N_2142);
and U3050 (N_3050,N_186,N_620);
nand U3051 (N_3051,N_2684,N_2118);
nand U3052 (N_3052,N_990,N_720);
and U3053 (N_3053,N_2224,N_1366);
nand U3054 (N_3054,N_2044,N_442);
nor U3055 (N_3055,N_2792,N_2018);
nand U3056 (N_3056,N_1505,N_2651);
nand U3057 (N_3057,N_1284,N_984);
nor U3058 (N_3058,N_1028,N_1740);
and U3059 (N_3059,N_1234,N_322);
xor U3060 (N_3060,N_181,N_2981);
and U3061 (N_3061,N_759,N_2970);
nand U3062 (N_3062,N_1448,N_1103);
and U3063 (N_3063,N_503,N_1333);
and U3064 (N_3064,N_2425,N_614);
nor U3065 (N_3065,N_1855,N_1527);
and U3066 (N_3066,N_2794,N_2136);
nor U3067 (N_3067,N_1879,N_1470);
nor U3068 (N_3068,N_2757,N_2589);
nand U3069 (N_3069,N_1428,N_2184);
or U3070 (N_3070,N_1866,N_2083);
xor U3071 (N_3071,N_2747,N_1271);
and U3072 (N_3072,N_2341,N_1889);
and U3073 (N_3073,N_965,N_373);
and U3074 (N_3074,N_2664,N_660);
nand U3075 (N_3075,N_1229,N_2925);
nand U3076 (N_3076,N_2368,N_1750);
nor U3077 (N_3077,N_253,N_159);
nand U3078 (N_3078,N_479,N_2440);
or U3079 (N_3079,N_334,N_1443);
nand U3080 (N_3080,N_718,N_1567);
nor U3081 (N_3081,N_949,N_687);
nor U3082 (N_3082,N_207,N_2766);
or U3083 (N_3083,N_2063,N_2340);
nand U3084 (N_3084,N_2861,N_1638);
and U3085 (N_3085,N_1992,N_1890);
and U3086 (N_3086,N_1952,N_1938);
and U3087 (N_3087,N_1558,N_1858);
or U3088 (N_3088,N_2031,N_1411);
nand U3089 (N_3089,N_212,N_907);
nor U3090 (N_3090,N_1742,N_2042);
nor U3091 (N_3091,N_1144,N_93);
nor U3092 (N_3092,N_531,N_888);
or U3093 (N_3093,N_1391,N_2007);
nor U3094 (N_3094,N_751,N_2326);
or U3095 (N_3095,N_627,N_2160);
and U3096 (N_3096,N_1590,N_2827);
or U3097 (N_3097,N_2991,N_2453);
and U3098 (N_3098,N_944,N_675);
or U3099 (N_3099,N_992,N_2845);
nor U3100 (N_3100,N_1387,N_691);
nor U3101 (N_3101,N_1456,N_669);
nand U3102 (N_3102,N_1833,N_2895);
nor U3103 (N_3103,N_1845,N_1407);
and U3104 (N_3104,N_1731,N_2662);
nand U3105 (N_3105,N_2610,N_1588);
nor U3106 (N_3106,N_1023,N_2898);
xnor U3107 (N_3107,N_1549,N_1329);
nand U3108 (N_3108,N_1530,N_2374);
and U3109 (N_3109,N_2641,N_189);
and U3110 (N_3110,N_2020,N_2501);
or U3111 (N_3111,N_609,N_355);
nand U3112 (N_3112,N_2727,N_509);
or U3113 (N_3113,N_804,N_192);
xor U3114 (N_3114,N_1482,N_2030);
nor U3115 (N_3115,N_824,N_161);
or U3116 (N_3116,N_2145,N_1086);
or U3117 (N_3117,N_1123,N_844);
nand U3118 (N_3118,N_229,N_1943);
nor U3119 (N_3119,N_1337,N_1054);
nor U3120 (N_3120,N_790,N_2585);
nor U3121 (N_3121,N_2858,N_243);
or U3122 (N_3122,N_668,N_632);
nand U3123 (N_3123,N_1143,N_2249);
or U3124 (N_3124,N_2108,N_1209);
nand U3125 (N_3125,N_1705,N_197);
or U3126 (N_3126,N_356,N_2574);
nor U3127 (N_3127,N_2093,N_2856);
and U3128 (N_3128,N_1165,N_1999);
and U3129 (N_3129,N_277,N_85);
nand U3130 (N_3130,N_1586,N_2413);
nand U3131 (N_3131,N_2596,N_2404);
and U3132 (N_3132,N_1629,N_612);
xor U3133 (N_3133,N_2303,N_1001);
nor U3134 (N_3134,N_1316,N_1733);
nand U3135 (N_3135,N_2759,N_2069);
and U3136 (N_3136,N_385,N_1545);
nor U3137 (N_3137,N_1370,N_2935);
xor U3138 (N_3138,N_2163,N_1679);
xnor U3139 (N_3139,N_834,N_2572);
nor U3140 (N_3140,N_1120,N_541);
or U3141 (N_3141,N_2985,N_1698);
and U3142 (N_3142,N_2079,N_550);
and U3143 (N_3143,N_2939,N_2584);
and U3144 (N_3144,N_1159,N_1270);
nor U3145 (N_3145,N_1049,N_421);
or U3146 (N_3146,N_953,N_2693);
or U3147 (N_3147,N_445,N_1793);
or U3148 (N_3148,N_1072,N_1512);
and U3149 (N_3149,N_1675,N_1185);
and U3150 (N_3150,N_1900,N_484);
nand U3151 (N_3151,N_1635,N_1918);
nand U3152 (N_3152,N_1281,N_409);
nand U3153 (N_3153,N_1220,N_1202);
xnor U3154 (N_3154,N_1319,N_105);
and U3155 (N_3155,N_1499,N_2254);
nor U3156 (N_3156,N_321,N_1783);
xor U3157 (N_3157,N_427,N_1575);
nand U3158 (N_3158,N_516,N_1324);
and U3159 (N_3159,N_383,N_2147);
or U3160 (N_3160,N_2522,N_2458);
or U3161 (N_3161,N_505,N_848);
nand U3162 (N_3162,N_2677,N_2011);
nand U3163 (N_3163,N_359,N_2557);
or U3164 (N_3164,N_1860,N_1475);
nor U3165 (N_3165,N_2164,N_585);
and U3166 (N_3166,N_1597,N_513);
and U3167 (N_3167,N_1109,N_1183);
nor U3168 (N_3168,N_2000,N_95);
and U3169 (N_3169,N_87,N_1901);
and U3170 (N_3170,N_1160,N_2524);
nand U3171 (N_3171,N_868,N_1497);
or U3172 (N_3172,N_119,N_255);
or U3173 (N_3173,N_961,N_1665);
nand U3174 (N_3174,N_2484,N_1042);
nor U3175 (N_3175,N_815,N_1080);
nor U3176 (N_3176,N_2810,N_141);
nand U3177 (N_3177,N_361,N_1722);
and U3178 (N_3178,N_2377,N_589);
nor U3179 (N_3179,N_2571,N_2806);
nor U3180 (N_3180,N_135,N_778);
or U3181 (N_3181,N_2888,N_2882);
nand U3182 (N_3182,N_854,N_1829);
or U3183 (N_3183,N_2014,N_753);
nand U3184 (N_3184,N_2434,N_1169);
or U3185 (N_3185,N_534,N_1419);
or U3186 (N_3186,N_1707,N_2361);
and U3187 (N_3187,N_1719,N_1467);
nand U3188 (N_3188,N_637,N_615);
and U3189 (N_3189,N_573,N_1155);
and U3190 (N_3190,N_746,N_2299);
nor U3191 (N_3191,N_1529,N_572);
nand U3192 (N_3192,N_2243,N_145);
or U3193 (N_3193,N_2753,N_279);
and U3194 (N_3194,N_1442,N_114);
and U3195 (N_3195,N_1418,N_1591);
nand U3196 (N_3196,N_1771,N_969);
nand U3197 (N_3197,N_1294,N_2847);
nand U3198 (N_3198,N_1314,N_1613);
nor U3199 (N_3199,N_847,N_2466);
nor U3200 (N_3200,N_1173,N_743);
nand U3201 (N_3201,N_1382,N_846);
nand U3202 (N_3202,N_113,N_317);
or U3203 (N_3203,N_1636,N_2071);
nor U3204 (N_3204,N_74,N_2887);
nor U3205 (N_3205,N_560,N_1417);
or U3206 (N_3206,N_2725,N_2609);
or U3207 (N_3207,N_2526,N_947);
nor U3208 (N_3208,N_1709,N_324);
nor U3209 (N_3209,N_1269,N_118);
or U3210 (N_3210,N_1827,N_511);
or U3211 (N_3211,N_2611,N_2566);
nand U3212 (N_3212,N_1596,N_1353);
and U3213 (N_3213,N_291,N_1227);
or U3214 (N_3214,N_1728,N_196);
nand U3215 (N_3215,N_2172,N_108);
and U3216 (N_3216,N_2003,N_677);
nand U3217 (N_3217,N_2120,N_2293);
nor U3218 (N_3218,N_2032,N_443);
or U3219 (N_3219,N_2039,N_2883);
and U3220 (N_3220,N_2781,N_268);
xnor U3221 (N_3221,N_2102,N_987);
or U3222 (N_3222,N_1649,N_1201);
xnor U3223 (N_3223,N_2124,N_1255);
nor U3224 (N_3224,N_1318,N_2036);
and U3225 (N_3225,N_2080,N_2868);
nor U3226 (N_3226,N_2786,N_597);
or U3227 (N_3227,N_1487,N_14);
nand U3228 (N_3228,N_1395,N_2715);
nor U3229 (N_3229,N_775,N_1790);
nor U3230 (N_3230,N_293,N_993);
or U3231 (N_3231,N_481,N_1376);
nor U3232 (N_3232,N_1538,N_958);
nand U3233 (N_3233,N_314,N_507);
and U3234 (N_3234,N_2351,N_1122);
and U3235 (N_3235,N_2699,N_2756);
nand U3236 (N_3236,N_1666,N_2698);
or U3237 (N_3237,N_1661,N_2182);
or U3238 (N_3238,N_1498,N_2265);
nor U3239 (N_3239,N_1096,N_1960);
nand U3240 (N_3240,N_1163,N_1701);
nand U3241 (N_3241,N_2625,N_110);
nor U3242 (N_3242,N_802,N_126);
or U3243 (N_3243,N_2737,N_727);
or U3244 (N_3244,N_1189,N_1533);
and U3245 (N_3245,N_2438,N_914);
or U3246 (N_3246,N_859,N_2089);
and U3247 (N_3247,N_547,N_1018);
or U3248 (N_3248,N_2795,N_2683);
or U3249 (N_3249,N_428,N_203);
nand U3250 (N_3250,N_1643,N_1587);
nor U3251 (N_3251,N_2754,N_1090);
and U3252 (N_3252,N_719,N_806);
or U3253 (N_3253,N_856,N_1039);
nand U3254 (N_3254,N_1432,N_67);
nor U3255 (N_3255,N_1204,N_1364);
nor U3256 (N_3256,N_716,N_2387);
and U3257 (N_3257,N_2734,N_368);
xnor U3258 (N_3258,N_2646,N_1823);
and U3259 (N_3259,N_1126,N_1552);
or U3260 (N_3260,N_1133,N_880);
nand U3261 (N_3261,N_1258,N_2494);
and U3262 (N_3262,N_2969,N_730);
nand U3263 (N_3263,N_1044,N_1261);
and U3264 (N_3264,N_2209,N_881);
or U3265 (N_3265,N_2323,N_2594);
and U3266 (N_3266,N_1776,N_2949);
nand U3267 (N_3267,N_357,N_1152);
nand U3268 (N_3268,N_741,N_1013);
and U3269 (N_3269,N_595,N_2195);
and U3270 (N_3270,N_2964,N_2608);
xor U3271 (N_3271,N_728,N_1251);
or U3272 (N_3272,N_1979,N_2285);
or U3273 (N_3273,N_2697,N_2170);
nor U3274 (N_3274,N_2733,N_2782);
nor U3275 (N_3275,N_257,N_171);
nor U3276 (N_3276,N_1891,N_1);
xor U3277 (N_3277,N_1279,N_2614);
nor U3278 (N_3278,N_1190,N_799);
or U3279 (N_3279,N_2426,N_2808);
nor U3280 (N_3280,N_475,N_1430);
or U3281 (N_3281,N_2360,N_2783);
or U3282 (N_3282,N_2167,N_2101);
and U3283 (N_3283,N_1998,N_2132);
nor U3284 (N_3284,N_1885,N_470);
xor U3285 (N_3285,N_578,N_616);
nand U3286 (N_3286,N_2119,N_1494);
and U3287 (N_3287,N_1600,N_28);
nand U3288 (N_3288,N_2098,N_1799);
or U3289 (N_3289,N_1566,N_593);
nand U3290 (N_3290,N_447,N_1170);
and U3291 (N_3291,N_1621,N_285);
nor U3292 (N_3292,N_2331,N_226);
and U3293 (N_3293,N_1029,N_598);
or U3294 (N_3294,N_2722,N_1438);
nand U3295 (N_3295,N_1875,N_2223);
nand U3296 (N_3296,N_750,N_2175);
or U3297 (N_3297,N_1589,N_588);
nor U3298 (N_3298,N_2633,N_1784);
or U3299 (N_3299,N_2463,N_1219);
nand U3300 (N_3300,N_2680,N_1871);
or U3301 (N_3301,N_2022,N_332);
or U3302 (N_3302,N_490,N_1046);
and U3303 (N_3303,N_2780,N_954);
nand U3304 (N_3304,N_89,N_905);
and U3305 (N_3305,N_301,N_2834);
nor U3306 (N_3306,N_2073,N_2705);
or U3307 (N_3307,N_178,N_2380);
and U3308 (N_3308,N_111,N_629);
or U3309 (N_3309,N_584,N_2517);
and U3310 (N_3310,N_643,N_2230);
nor U3311 (N_3311,N_2359,N_1349);
and U3312 (N_3312,N_2672,N_2393);
and U3313 (N_3313,N_1727,N_173);
nor U3314 (N_3314,N_2710,N_2140);
nand U3315 (N_3315,N_400,N_1259);
or U3316 (N_3316,N_496,N_2258);
or U3317 (N_3317,N_1064,N_2886);
or U3318 (N_3318,N_2558,N_734);
nor U3319 (N_3319,N_98,N_1604);
nor U3320 (N_3320,N_2822,N_1618);
and U3321 (N_3321,N_1786,N_11);
nand U3322 (N_3322,N_2112,N_685);
or U3323 (N_3323,N_2338,N_97);
nand U3324 (N_3324,N_388,N_244);
and U3325 (N_3325,N_2605,N_1897);
nand U3326 (N_3326,N_195,N_619);
nand U3327 (N_3327,N_2122,N_367);
nor U3328 (N_3328,N_239,N_2681);
and U3329 (N_3329,N_2666,N_2905);
nor U3330 (N_3330,N_2502,N_681);
or U3331 (N_3331,N_1902,N_1058);
nand U3332 (N_3332,N_2477,N_1045);
and U3333 (N_3333,N_250,N_2926);
and U3334 (N_3334,N_347,N_1555);
nor U3335 (N_3335,N_331,N_2505);
nor U3336 (N_3336,N_749,N_403);
nor U3337 (N_3337,N_2527,N_956);
nand U3338 (N_3338,N_1304,N_1933);
nor U3339 (N_3339,N_1547,N_1822);
or U3340 (N_3340,N_2247,N_1704);
nor U3341 (N_3341,N_1610,N_2910);
and U3342 (N_3342,N_1124,N_2573);
nor U3343 (N_3343,N_840,N_1321);
nor U3344 (N_3344,N_1373,N_2156);
or U3345 (N_3345,N_164,N_1343);
or U3346 (N_3346,N_1789,N_1848);
nor U3347 (N_3347,N_875,N_2049);
nor U3348 (N_3348,N_2062,N_2474);
nand U3349 (N_3349,N_2017,N_939);
nand U3350 (N_3350,N_2966,N_1754);
and U3351 (N_3351,N_29,N_2383);
nor U3352 (N_3352,N_134,N_2053);
nand U3353 (N_3353,N_1753,N_1509);
nand U3354 (N_3354,N_2240,N_704);
nand U3355 (N_3355,N_2729,N_527);
nor U3356 (N_3356,N_39,N_2736);
or U3357 (N_3357,N_957,N_813);
or U3358 (N_3358,N_2429,N_2612);
nand U3359 (N_3359,N_2028,N_432);
nand U3360 (N_3360,N_913,N_2242);
or U3361 (N_3361,N_2791,N_57);
nand U3362 (N_3362,N_248,N_1562);
and U3363 (N_3363,N_890,N_1300);
nor U3364 (N_3364,N_1836,N_2128);
xnor U3365 (N_3365,N_2913,N_2961);
and U3366 (N_3366,N_885,N_1747);
nand U3367 (N_3367,N_468,N_2298);
or U3368 (N_3368,N_2998,N_1863);
or U3369 (N_3369,N_2983,N_2823);
nand U3370 (N_3370,N_2047,N_2567);
or U3371 (N_3371,N_1479,N_252);
nor U3372 (N_3372,N_2437,N_2520);
nand U3373 (N_3373,N_1496,N_665);
and U3374 (N_3374,N_84,N_2016);
or U3375 (N_3375,N_2492,N_1296);
and U3376 (N_3376,N_1852,N_167);
or U3377 (N_3377,N_107,N_1415);
and U3378 (N_3378,N_2357,N_1454);
or U3379 (N_3379,N_1557,N_1951);
nand U3380 (N_3380,N_1367,N_571);
nor U3381 (N_3381,N_940,N_1288);
or U3382 (N_3382,N_1995,N_842);
nand U3383 (N_3383,N_2916,N_1068);
and U3384 (N_3384,N_146,N_1581);
and U3385 (N_3385,N_459,N_92);
nor U3386 (N_3386,N_1535,N_254);
nor U3387 (N_3387,N_283,N_2933);
nand U3388 (N_3388,N_2691,N_61);
and U3389 (N_3389,N_2545,N_1328);
xor U3390 (N_3390,N_2192,N_821);
or U3391 (N_3391,N_492,N_1221);
and U3392 (N_3392,N_1702,N_2850);
nor U3393 (N_3393,N_2838,N_2473);
nor U3394 (N_3394,N_1921,N_1652);
nand U3395 (N_3395,N_973,N_1940);
nor U3396 (N_3396,N_2457,N_2256);
nand U3397 (N_3397,N_32,N_1473);
and U3398 (N_3398,N_59,N_2407);
and U3399 (N_3399,N_1762,N_2282);
and U3400 (N_3400,N_2655,N_1350);
nand U3401 (N_3401,N_1544,N_1317);
nor U3402 (N_3402,N_2078,N_1162);
nand U3403 (N_3403,N_1977,N_2577);
or U3404 (N_3404,N_2645,N_233);
and U3405 (N_3405,N_2601,N_2931);
nand U3406 (N_3406,N_1135,N_2695);
or U3407 (N_3407,N_58,N_2021);
nand U3408 (N_3408,N_2944,N_1856);
and U3409 (N_3409,N_2009,N_828);
or U3410 (N_3410,N_912,N_2730);
and U3411 (N_3411,N_1476,N_853);
nand U3412 (N_3412,N_2410,N_683);
nor U3413 (N_3413,N_49,N_62);
or U3414 (N_3414,N_2619,N_1208);
or U3415 (N_3415,N_1292,N_917);
nor U3416 (N_3416,N_316,N_274);
xor U3417 (N_3417,N_2864,N_2065);
nand U3418 (N_3418,N_2771,N_2312);
nand U3419 (N_3419,N_1368,N_16);
and U3420 (N_3420,N_2744,N_696);
and U3421 (N_3421,N_1660,N_2694);
nand U3422 (N_3422,N_345,N_2620);
and U3423 (N_3423,N_2726,N_1434);
and U3424 (N_3424,N_2309,N_1775);
nand U3425 (N_3425,N_482,N_2513);
and U3426 (N_3426,N_2951,N_1912);
nand U3427 (N_3427,N_1093,N_722);
nand U3428 (N_3428,N_1254,N_44);
or U3429 (N_3429,N_765,N_1560);
xnor U3430 (N_3430,N_1516,N_319);
and U3431 (N_3431,N_262,N_2201);
or U3432 (N_3432,N_2547,N_287);
and U3433 (N_3433,N_418,N_525);
and U3434 (N_3434,N_485,N_5);
nor U3435 (N_3435,N_517,N_1232);
nor U3436 (N_3436,N_1813,N_671);
or U3437 (N_3437,N_2804,N_486);
nand U3438 (N_3438,N_1027,N_2334);
nor U3439 (N_3439,N_1101,N_1346);
and U3440 (N_3440,N_2352,N_610);
and U3441 (N_3441,N_2421,N_2131);
nand U3442 (N_3442,N_2061,N_1272);
and U3443 (N_3443,N_1928,N_1131);
and U3444 (N_3444,N_2511,N_1031);
and U3445 (N_3445,N_2389,N_2464);
or U3446 (N_3446,N_2129,N_1510);
and U3447 (N_3447,N_2920,N_2642);
or U3448 (N_3448,N_874,N_2234);
nand U3449 (N_3449,N_613,N_312);
and U3450 (N_3450,N_349,N_152);
nor U3451 (N_3451,N_561,N_182);
nor U3452 (N_3452,N_2321,N_2909);
and U3453 (N_3453,N_1989,N_1524);
and U3454 (N_3454,N_1214,N_713);
nor U3455 (N_3455,N_2973,N_1186);
and U3456 (N_3456,N_1097,N_100);
and U3457 (N_3457,N_893,N_2470);
or U3458 (N_3458,N_60,N_776);
nor U3459 (N_3459,N_2322,N_2554);
or U3460 (N_3460,N_1307,N_2603);
and U3461 (N_3461,N_908,N_1615);
or U3462 (N_3462,N_2213,N_2319);
xor U3463 (N_3463,N_223,N_2491);
or U3464 (N_3464,N_389,N_2496);
nor U3465 (N_3465,N_607,N_1913);
nor U3466 (N_3466,N_1215,N_2365);
and U3467 (N_3467,N_748,N_2154);
nand U3468 (N_3468,N_576,N_2994);
and U3469 (N_3469,N_333,N_767);
nand U3470 (N_3470,N_1386,N_756);
or U3471 (N_3471,N_2005,N_1797);
nand U3472 (N_3472,N_872,N_472);
and U3473 (N_3473,N_975,N_1686);
or U3474 (N_3474,N_2957,N_787);
and U3475 (N_3475,N_2659,N_551);
nor U3476 (N_3476,N_2207,N_272);
nand U3477 (N_3477,N_2235,N_2354);
or U3478 (N_3478,N_2187,N_2210);
nand U3479 (N_3479,N_315,N_1840);
or U3480 (N_3480,N_394,N_1355);
nor U3481 (N_3481,N_583,N_2890);
nand U3482 (N_3482,N_2863,N_762);
and U3483 (N_3483,N_2023,N_1495);
or U3484 (N_3484,N_1584,N_2576);
nor U3485 (N_3485,N_27,N_2873);
and U3486 (N_3486,N_1462,N_1238);
or U3487 (N_3487,N_672,N_360);
nand U3488 (N_3488,N_2125,N_1689);
or U3489 (N_3489,N_305,N_537);
nor U3490 (N_3490,N_735,N_608);
and U3491 (N_3491,N_2741,N_1950);
or U3492 (N_3492,N_1464,N_2095);
or U3493 (N_3493,N_1503,N_2064);
nand U3494 (N_3494,N_1816,N_1260);
nor U3495 (N_3495,N_1769,N_2904);
and U3496 (N_3496,N_1005,N_267);
and U3497 (N_3497,N_402,N_733);
xor U3498 (N_3498,N_1670,N_2819);
nor U3499 (N_3499,N_2402,N_1542);
and U3500 (N_3500,N_2586,N_1298);
nand U3501 (N_3501,N_2504,N_2435);
or U3502 (N_3502,N_1198,N_1257);
and U3503 (N_3503,N_260,N_2692);
and U3504 (N_3504,N_1658,N_902);
or U3505 (N_3505,N_858,N_1128);
or U3506 (N_3506,N_1306,N_1465);
nor U3507 (N_3507,N_2489,N_117);
nand U3508 (N_3508,N_2872,N_2165);
or U3509 (N_3509,N_1819,N_144);
nor U3510 (N_3510,N_2486,N_798);
nand U3511 (N_3511,N_2701,N_694);
nor U3512 (N_3512,N_180,N_1550);
nor U3513 (N_3513,N_1708,N_2013);
or U3514 (N_3514,N_1655,N_667);
and U3515 (N_3515,N_221,N_2855);
or U3516 (N_3516,N_24,N_772);
or U3517 (N_3517,N_884,N_344);
and U3518 (N_3518,N_702,N_2599);
or U3519 (N_3519,N_967,N_2498);
nand U3520 (N_3520,N_441,N_1972);
nand U3521 (N_3521,N_2467,N_1752);
nor U3522 (N_3522,N_231,N_2001);
nand U3523 (N_3523,N_469,N_835);
nand U3524 (N_3524,N_2840,N_1887);
nor U3525 (N_3525,N_1818,N_1745);
nor U3526 (N_3526,N_392,N_1569);
nand U3527 (N_3527,N_1773,N_2649);
nand U3528 (N_3528,N_1026,N_2943);
nor U3529 (N_3529,N_1312,N_931);
nor U3530 (N_3530,N_1807,N_1037);
xor U3531 (N_3531,N_1853,N_80);
nor U3532 (N_3532,N_2493,N_2738);
or U3533 (N_3533,N_1910,N_370);
nand U3534 (N_3534,N_860,N_2211);
nor U3535 (N_3535,N_1377,N_1014);
nand U3536 (N_3536,N_792,N_997);
or U3537 (N_3537,N_797,N_1975);
or U3538 (N_3538,N_1573,N_2428);
or U3539 (N_3539,N_586,N_999);
nand U3540 (N_3540,N_2743,N_456);
and U3541 (N_3541,N_2244,N_717);
and U3542 (N_3542,N_1765,N_1617);
nor U3543 (N_3543,N_474,N_147);
nand U3544 (N_3544,N_2188,N_2653);
nand U3545 (N_3545,N_2392,N_1782);
nand U3546 (N_3546,N_2451,N_1132);
or U3547 (N_3547,N_2345,N_2639);
nor U3548 (N_3548,N_2475,N_1595);
nand U3549 (N_3549,N_1691,N_1110);
nand U3550 (N_3550,N_6,N_1158);
or U3551 (N_3551,N_298,N_2789);
and U3552 (N_3552,N_1446,N_700);
nor U3553 (N_3553,N_2449,N_2516);
nand U3554 (N_3554,N_1142,N_870);
and U3555 (N_3555,N_106,N_227);
nor U3556 (N_3556,N_2982,N_1250);
nor U3557 (N_3557,N_1330,N_2236);
or U3558 (N_3558,N_2521,N_904);
or U3559 (N_3559,N_125,N_2086);
nor U3560 (N_3560,N_937,N_1956);
or U3561 (N_3561,N_590,N_364);
or U3562 (N_3562,N_630,N_928);
nand U3563 (N_3563,N_2837,N_1511);
or U3564 (N_3564,N_2055,N_2816);
or U3565 (N_3565,N_2194,N_2682);
or U3566 (N_3566,N_215,N_396);
nor U3567 (N_3567,N_2885,N_862);
or U3568 (N_3568,N_2372,N_1015);
or U3569 (N_3569,N_366,N_1187);
or U3570 (N_3570,N_1690,N_1118);
or U3571 (N_3571,N_544,N_1463);
nor U3572 (N_3572,N_261,N_1396);
or U3573 (N_3573,N_2569,N_241);
and U3574 (N_3574,N_514,N_628);
or U3575 (N_3575,N_2562,N_124);
nand U3576 (N_3576,N_2186,N_929);
or U3577 (N_3577,N_891,N_1631);
nor U3578 (N_3578,N_935,N_656);
or U3579 (N_3579,N_692,N_165);
nand U3580 (N_3580,N_1011,N_2836);
and U3581 (N_3581,N_810,N_883);
or U3582 (N_3582,N_2665,N_430);
or U3583 (N_3583,N_2615,N_1849);
nand U3584 (N_3584,N_1694,N_1117);
nand U3585 (N_3585,N_1099,N_2094);
nor U3586 (N_3586,N_2739,N_1414);
and U3587 (N_3587,N_453,N_83);
nor U3588 (N_3588,N_2713,N_1310);
nor U3589 (N_3589,N_1094,N_2109);
nor U3590 (N_3590,N_563,N_1032);
and U3591 (N_3591,N_1401,N_2424);
or U3592 (N_3592,N_275,N_467);
nor U3593 (N_3593,N_601,N_457);
nor U3594 (N_3594,N_1749,N_379);
nor U3595 (N_3595,N_1627,N_960);
or U3596 (N_3596,N_296,N_47);
nand U3597 (N_3597,N_1757,N_3);
and U3598 (N_3598,N_362,N_666);
nor U3599 (N_3599,N_1423,N_1303);
nor U3600 (N_3600,N_809,N_2168);
nand U3601 (N_3601,N_2852,N_2183);
nor U3602 (N_3602,N_2563,N_2476);
and U3603 (N_3603,N_2082,N_603);
or U3604 (N_3604,N_1226,N_782);
nand U3605 (N_3605,N_2912,N_1883);
nand U3606 (N_3606,N_130,N_1968);
xnor U3607 (N_3607,N_2214,N_2185);
nor U3608 (N_3608,N_313,N_249);
nor U3609 (N_3609,N_2150,N_104);
and U3610 (N_3610,N_1282,N_410);
and U3611 (N_3611,N_1523,N_2769);
or U3612 (N_3612,N_966,N_434);
nor U3613 (N_3613,N_2825,N_1253);
and U3614 (N_3614,N_1870,N_2272);
nand U3615 (N_3615,N_808,N_318);
or U3616 (N_3616,N_2661,N_26);
nor U3617 (N_3617,N_1127,N_1920);
or U3618 (N_3618,N_655,N_1399);
or U3619 (N_3619,N_2518,N_2897);
nand U3620 (N_3620,N_894,N_1336);
or U3621 (N_3621,N_1682,N_2010);
nand U3622 (N_3622,N_2499,N_783);
or U3623 (N_3623,N_1939,N_2500);
or U3624 (N_3624,N_2394,N_1084);
nand U3625 (N_3625,N_1177,N_2388);
and U3626 (N_3626,N_1565,N_2252);
or U3627 (N_3627,N_581,N_2483);
nand U3628 (N_3628,N_2137,N_2654);
and U3629 (N_3629,N_1315,N_2050);
and U3630 (N_3630,N_2941,N_661);
or U3631 (N_3631,N_1664,N_2329);
nand U3632 (N_3632,N_755,N_1426);
or U3633 (N_3633,N_1400,N_1800);
and U3634 (N_3634,N_2918,N_1334);
nor U3635 (N_3635,N_426,N_2849);
nand U3636 (N_3636,N_214,N_1985);
nand U3637 (N_3637,N_822,N_1299);
nor U3638 (N_3638,N_54,N_766);
xnor U3639 (N_3639,N_715,N_2465);
nor U3640 (N_3640,N_1515,N_689);
nor U3641 (N_3641,N_1138,N_2141);
nor U3642 (N_3642,N_1077,N_1508);
nor U3643 (N_3643,N_1559,N_1233);
or U3644 (N_3644,N_2347,N_1895);
nand U3645 (N_3645,N_2024,N_1263);
and U3646 (N_3646,N_2975,N_2509);
and U3647 (N_3647,N_1331,N_555);
and U3648 (N_3648,N_185,N_451);
and U3649 (N_3649,N_292,N_1320);
nand U3650 (N_3650,N_827,N_2278);
nor U3651 (N_3651,N_830,N_2647);
nand U3652 (N_3652,N_2763,N_2503);
and U3653 (N_3653,N_1632,N_2604);
nor U3654 (N_3654,N_1130,N_1452);
and U3655 (N_3655,N_1688,N_1983);
or U3656 (N_3656,N_1025,N_2056);
nand U3657 (N_3657,N_2900,N_2675);
and U3658 (N_3658,N_1898,N_1801);
nand U3659 (N_3659,N_1228,N_1625);
nor U3660 (N_3660,N_2399,N_72);
or U3661 (N_3661,N_1469,N_2958);
and U3662 (N_3662,N_81,N_150);
or U3663 (N_3663,N_22,N_1265);
xor U3664 (N_3664,N_1075,N_236);
or U3665 (N_3665,N_723,N_2839);
and U3666 (N_3666,N_1129,N_2990);
and U3667 (N_3667,N_1876,N_166);
nand U3668 (N_3668,N_596,N_1019);
nand U3669 (N_3669,N_2087,N_2433);
nor U3670 (N_3670,N_529,N_458);
nand U3671 (N_3671,N_1344,N_2130);
or U3672 (N_3672,N_781,N_906);
or U3673 (N_3673,N_1814,N_2406);
nor U3674 (N_3674,N_417,N_1824);
and U3675 (N_3675,N_1948,N_295);
or U3676 (N_3676,N_2917,N_446);
and U3677 (N_3677,N_2613,N_2671);
nor U3678 (N_3678,N_160,N_500);
xor U3679 (N_3679,N_1838,N_566);
nand U3680 (N_3680,N_2706,N_1582);
and U3681 (N_3681,N_1008,N_30);
nor U3682 (N_3682,N_384,N_1358);
xor U3683 (N_3683,N_2105,N_971);
or U3684 (N_3684,N_565,N_579);
nor U3685 (N_3685,N_1175,N_391);
and U3686 (N_3686,N_602,N_2487);
nor U3687 (N_3687,N_2412,N_570);
or U3688 (N_3688,N_2914,N_1179);
nand U3689 (N_3689,N_1057,N_568);
nand U3690 (N_3690,N_1390,N_2507);
or U3691 (N_3691,N_641,N_155);
or U3692 (N_3692,N_1609,N_2307);
xnor U3693 (N_3693,N_230,N_1844);
nor U3694 (N_3694,N_1164,N_1427);
nor U3695 (N_3695,N_1699,N_2418);
nand U3696 (N_3696,N_836,N_1449);
and U3697 (N_3697,N_63,N_512);
and U3698 (N_3698,N_86,N_1153);
nor U3699 (N_3699,N_1051,N_1861);
and U3700 (N_3700,N_763,N_921);
nand U3701 (N_3701,N_2922,N_995);
nor U3702 (N_3702,N_1791,N_2761);
and U3703 (N_3703,N_1460,N_2276);
nor U3704 (N_3704,N_2099,N_270);
nor U3705 (N_3705,N_2788,N_1341);
xor U3706 (N_3706,N_592,N_951);
and U3707 (N_3707,N_404,N_1506);
or U3708 (N_3708,N_2621,N_2405);
nand U3709 (N_3709,N_2369,N_991);
nor U3710 (N_3710,N_1904,N_365);
or U3711 (N_3711,N_1195,N_228);
or U3712 (N_3712,N_1821,N_1035);
nor U3713 (N_3713,N_2748,N_710);
or U3714 (N_3714,N_40,N_397);
nor U3715 (N_3715,N_2229,N_649);
nand U3716 (N_3716,N_538,N_2088);
nand U3717 (N_3717,N_2790,N_1974);
or U3718 (N_3718,N_1107,N_1285);
and U3719 (N_3719,N_2004,N_1717);
or U3720 (N_3720,N_638,N_2266);
or U3721 (N_3721,N_2714,N_2490);
nand U3722 (N_3722,N_1720,N_2395);
and U3723 (N_3723,N_1381,N_695);
or U3724 (N_3724,N_536,N_2422);
xnor U3725 (N_3725,N_1137,N_1338);
nor U3726 (N_3726,N_339,N_9);
and U3727 (N_3727,N_2987,N_2901);
nor U3728 (N_3728,N_724,N_1809);
and U3729 (N_3729,N_1012,N_923);
nand U3730 (N_3730,N_2928,N_183);
nand U3731 (N_3731,N_2638,N_1896);
or U3732 (N_3732,N_1540,N_1907);
xnor U3733 (N_3733,N_2301,N_673);
and U3734 (N_3734,N_1624,N_1398);
nor U3735 (N_3735,N_372,N_290);
or U3736 (N_3736,N_1422,N_2950);
nand U3737 (N_3737,N_1546,N_1991);
nand U3738 (N_3738,N_2408,N_1614);
or U3739 (N_3739,N_1236,N_623);
and U3740 (N_3740,N_1961,N_2191);
or U3741 (N_3741,N_1095,N_2600);
and U3742 (N_3742,N_2844,N_2411);
nand U3743 (N_3743,N_1283,N_2776);
nor U3744 (N_3744,N_2963,N_1881);
nor U3745 (N_3745,N_1106,N_2535);
or U3746 (N_3746,N_1191,N_2295);
nand U3747 (N_3747,N_2543,N_2813);
nand U3748 (N_3748,N_805,N_1803);
nor U3749 (N_3749,N_2197,N_1360);
nand U3750 (N_3750,N_1772,N_68);
nand U3751 (N_3751,N_269,N_2817);
and U3752 (N_3752,N_1681,N_1157);
nand U3753 (N_3753,N_2658,N_419);
and U3754 (N_3754,N_1949,N_99);
nor U3755 (N_3755,N_855,N_2348);
nor U3756 (N_3756,N_2959,N_959);
or U3757 (N_3757,N_2072,N_2262);
nand U3758 (N_3758,N_1929,N_1273);
nor U3759 (N_3759,N_1804,N_676);
nor U3760 (N_3760,N_1859,N_2828);
and U3761 (N_3761,N_2720,N_941);
nor U3762 (N_3762,N_247,N_2860);
nand U3763 (N_3763,N_1758,N_1222);
and U3764 (N_3764,N_148,N_1504);
or U3765 (N_3765,N_2181,N_1802);
nand U3766 (N_3766,N_769,N_1847);
or U3767 (N_3767,N_2690,N_1016);
and U3768 (N_3768,N_1112,N_1841);
nor U3769 (N_3769,N_1919,N_2673);
and U3770 (N_3770,N_1725,N_2765);
and U3771 (N_3771,N_2704,N_2986);
or U3772 (N_3772,N_2454,N_1436);
nor U3773 (N_3773,N_2259,N_2934);
nand U3774 (N_3774,N_1593,N_2034);
nand U3775 (N_3775,N_2667,N_120);
nand U3776 (N_3776,N_886,N_879);
nor U3777 (N_3777,N_101,N_2923);
nand U3778 (N_3778,N_2376,N_175);
nor U3779 (N_3779,N_174,N_140);
and U3780 (N_3780,N_803,N_962);
nand U3781 (N_3781,N_1888,N_742);
or U3782 (N_3782,N_193,N_1990);
or U3783 (N_3783,N_542,N_721);
or U3784 (N_3784,N_1926,N_1212);
nand U3785 (N_3785,N_2927,N_1501);
or U3786 (N_3786,N_708,N_1656);
nor U3787 (N_3787,N_2315,N_1851);
and U3788 (N_3788,N_1811,N_737);
and U3789 (N_3789,N_2552,N_2519);
or U3790 (N_3790,N_1047,N_1993);
nand U3791 (N_3791,N_2104,N_2565);
or U3792 (N_3792,N_2157,N_498);
or U3793 (N_3793,N_2723,N_1252);
or U3794 (N_3794,N_1351,N_1578);
nand U3795 (N_3795,N_1323,N_1410);
nor U3796 (N_3796,N_1606,N_645);
and U3797 (N_3797,N_477,N_892);
and U3798 (N_3798,N_955,N_1732);
and U3799 (N_3799,N_1140,N_1459);
nor U3800 (N_3800,N_1911,N_1718);
or U3801 (N_3801,N_1447,N_784);
and U3802 (N_3802,N_2143,N_2952);
nor U3803 (N_3803,N_1493,N_2344);
nor U3804 (N_3804,N_2286,N_1245);
nor U3805 (N_3805,N_2070,N_1551);
nand U3806 (N_3806,N_2891,N_518);
nor U3807 (N_3807,N_435,N_1672);
nor U3808 (N_3808,N_878,N_1739);
or U3809 (N_3809,N_217,N_1205);
nand U3810 (N_3810,N_1104,N_2173);
or U3811 (N_3811,N_2472,N_1941);
or U3812 (N_3812,N_422,N_745);
or U3813 (N_3813,N_2008,N_1628);
nor U3814 (N_3814,N_399,N_1440);
nand U3815 (N_3815,N_2356,N_789);
nand U3816 (N_3816,N_2040,N_2239);
and U3817 (N_3817,N_1302,N_213);
nor U3818 (N_3818,N_739,N_1211);
and U3819 (N_3819,N_2248,N_2506);
nor U3820 (N_3820,N_625,N_1743);
and U3821 (N_3821,N_535,N_2046);
or U3822 (N_3822,N_1713,N_401);
nand U3823 (N_3823,N_495,N_752);
nor U3824 (N_3824,N_841,N_2274);
nor U3825 (N_3825,N_1677,N_300);
and U3826 (N_3826,N_2712,N_2936);
or U3827 (N_3827,N_2110,N_2814);
or U3828 (N_3828,N_1004,N_2218);
and U3829 (N_3829,N_218,N_1893);
and U3830 (N_3830,N_2208,N_168);
or U3831 (N_3831,N_1715,N_2871);
nor U3832 (N_3832,N_688,N_77);
nor U3833 (N_3833,N_2401,N_712);
nor U3834 (N_3834,N_1207,N_1024);
xor U3835 (N_3835,N_1478,N_259);
or U3836 (N_3836,N_2432,N_2038);
or U3837 (N_3837,N_2090,N_2179);
or U3838 (N_3838,N_2478,N_2495);
nor U3839 (N_3839,N_553,N_172);
xnor U3840 (N_3840,N_2750,N_556);
and U3841 (N_3841,N_1361,N_838);
and U3842 (N_3842,N_2962,N_2279);
or U3843 (N_3843,N_2196,N_1022);
or U3844 (N_3844,N_819,N_1755);
and U3845 (N_3845,N_1729,N_1603);
nor U3846 (N_3846,N_66,N_96);
nand U3847 (N_3847,N_1340,N_1520);
nor U3848 (N_3848,N_2320,N_43);
xnor U3849 (N_3849,N_2398,N_2755);
and U3850 (N_3850,N_528,N_1468);
and U3851 (N_3851,N_646,N_1491);
or U3852 (N_3852,N_2346,N_2116);
nor U3853 (N_3853,N_626,N_2189);
nor U3854 (N_3854,N_1402,N_1197);
nand U3855 (N_3855,N_1842,N_2385);
nor U3856 (N_3856,N_1379,N_2960);
nor U3857 (N_3857,N_18,N_574);
xnor U3858 (N_3858,N_502,N_2059);
or U3859 (N_3859,N_179,N_2859);
or U3860 (N_3860,N_52,N_2821);
and U3861 (N_3861,N_2296,N_1692);
nand U3862 (N_3862,N_1295,N_2350);
and U3863 (N_3863,N_2430,N_2989);
nor U3864 (N_3864,N_2233,N_2025);
or U3865 (N_3865,N_2289,N_190);
nand U3866 (N_3866,N_1151,N_644);
and U3867 (N_3867,N_1714,N_2803);
nor U3868 (N_3868,N_240,N_533);
and U3869 (N_3869,N_2339,N_348);
or U3870 (N_3870,N_2674,N_2637);
and U3871 (N_3871,N_504,N_194);
or U3872 (N_3872,N_2865,N_1079);
and U3873 (N_3873,N_2937,N_1532);
nand U3874 (N_3874,N_1892,N_1378);
nand U3875 (N_3875,N_2283,N_1150);
nand U3876 (N_3876,N_1647,N_1243);
nor U3877 (N_3877,N_678,N_903);
or U3878 (N_3878,N_2251,N_1036);
or U3879 (N_3879,N_1561,N_1654);
or U3880 (N_3880,N_71,N_216);
nor U3881 (N_3881,N_2749,N_1695);
nor U3882 (N_3882,N_246,N_2327);
and U3883 (N_3883,N_2308,N_1805);
or U3884 (N_3884,N_91,N_1526);
and U3885 (N_3885,N_690,N_909);
or U3886 (N_3886,N_2171,N_2908);
or U3887 (N_3887,N_1081,N_220);
xor U3888 (N_3888,N_863,N_31);
or U3889 (N_3889,N_1067,N_869);
nor U3890 (N_3890,N_2807,N_2002);
or U3891 (N_3891,N_2420,N_1971);
and U3892 (N_3892,N_46,N_1787);
nor U3893 (N_3893,N_1059,N_251);
and U3894 (N_3894,N_1266,N_2809);
nand U3895 (N_3895,N_604,N_851);
or U3896 (N_3896,N_1017,N_1953);
nand U3897 (N_3897,N_2436,N_2174);
and U3898 (N_3898,N_2060,N_2811);
nand U3899 (N_3899,N_2445,N_698);
and U3900 (N_3900,N_1125,N_1038);
nand U3901 (N_3901,N_922,N_20);
nand U3902 (N_3902,N_811,N_816);
or U3903 (N_3903,N_2833,N_2728);
or U3904 (N_3904,N_340,N_2027);
nand U3905 (N_3905,N_1611,N_2006);
nor U3906 (N_3906,N_697,N_757);
nand U3907 (N_3907,N_557,N_1113);
or U3908 (N_3908,N_1835,N_812);
or U3909 (N_3909,N_338,N_53);
nand U3910 (N_3910,N_2940,N_2996);
or U3911 (N_3911,N_978,N_1461);
or U3912 (N_3912,N_2390,N_2735);
nand U3913 (N_3913,N_777,N_1623);
and U3914 (N_3914,N_429,N_1034);
nand U3915 (N_3915,N_770,N_1413);
nand U3916 (N_3916,N_1305,N_1241);
xor U3917 (N_3917,N_900,N_1180);
nand U3918 (N_3918,N_1564,N_69);
nor U3919 (N_3919,N_2169,N_1997);
and U3920 (N_3920,N_1223,N_2231);
nor U3921 (N_3921,N_2787,N_374);
and U3922 (N_3922,N_2978,N_994);
and U3923 (N_3923,N_1100,N_1988);
nand U3924 (N_3924,N_2660,N_2835);
nand U3925 (N_3925,N_1056,N_2052);
nand U3926 (N_3926,N_2956,N_2419);
and U3927 (N_3927,N_1916,N_837);
nor U3928 (N_3928,N_591,N_1669);
nand U3929 (N_3929,N_1706,N_408);
nor U3930 (N_3930,N_1942,N_1644);
and U3931 (N_3931,N_302,N_480);
nor U3932 (N_3932,N_1724,N_2134);
or U3933 (N_3933,N_1592,N_2724);
nor U3934 (N_3934,N_725,N_788);
and U3935 (N_3935,N_785,N_2550);
or U3936 (N_3936,N_1224,N_121);
and U3937 (N_3937,N_2220,N_2700);
nor U3938 (N_3938,N_2469,N_294);
nor U3939 (N_3939,N_2881,N_2275);
and U3940 (N_3940,N_2531,N_1696);
nor U3941 (N_3941,N_2302,N_2455);
or U3942 (N_3942,N_1837,N_658);
and U3943 (N_3943,N_1832,N_599);
nor U3944 (N_3944,N_375,N_1882);
nor U3945 (N_3945,N_1268,N_2598);
nand U3946 (N_3946,N_1810,N_2636);
nand U3947 (N_3947,N_1925,N_234);
nor U3948 (N_3948,N_2288,N_2903);
xor U3949 (N_3949,N_996,N_2624);
or U3950 (N_3950,N_2878,N_1980);
xor U3951 (N_3951,N_2077,N_310);
and U3952 (N_3952,N_263,N_242);
and U3953 (N_3953,N_1392,N_932);
and U3954 (N_3954,N_1311,N_2892);
or U3955 (N_3955,N_2199,N_924);
or U3956 (N_3956,N_138,N_554);
and U3957 (N_3957,N_2212,N_1231);
or U3958 (N_3958,N_437,N_703);
or U3959 (N_3959,N_1488,N_23);
or U3960 (N_3960,N_2075,N_1291);
nor U3961 (N_3961,N_1721,N_1363);
nand U3962 (N_3962,N_13,N_2826);
or U3963 (N_3963,N_25,N_2616);
nor U3964 (N_3964,N_462,N_1808);
and U3965 (N_3965,N_2232,N_1536);
nor U3966 (N_3966,N_2702,N_1798);
nand U3967 (N_3967,N_2919,N_2648);
nor U3968 (N_3968,N_1171,N_652);
xor U3969 (N_3969,N_1030,N_559);
nor U3970 (N_3970,N_2227,N_2267);
and U3971 (N_3971,N_2111,N_515);
or U3972 (N_3972,N_483,N_2403);
nor U3973 (N_3973,N_2284,N_2530);
and U3974 (N_3974,N_1667,N_549);
nor U3975 (N_3975,N_639,N_128);
nand U3976 (N_3976,N_1862,N_936);
nor U3977 (N_3977,N_2439,N_1339);
and U3978 (N_3978,N_2880,N_1437);
xor U3979 (N_3979,N_1978,N_2824);
nand U3980 (N_3980,N_2045,N_577);
and U3981 (N_3981,N_2622,N_2442);
nand U3982 (N_3982,N_1405,N_1830);
and U3983 (N_3983,N_2330,N_2764);
nor U3984 (N_3984,N_2379,N_1553);
and U3985 (N_3985,N_487,N_1406);
nand U3986 (N_3986,N_1471,N_2198);
or U3987 (N_3987,N_2607,N_1930);
nor U3988 (N_3988,N_1781,N_2618);
nor U3989 (N_3989,N_2029,N_64);
nor U3990 (N_3990,N_2371,N_524);
nor U3991 (N_3991,N_2427,N_2687);
or U3992 (N_3992,N_1619,N_1571);
xor U3993 (N_3993,N_1676,N_1884);
and U3994 (N_3994,N_82,N_303);
or U3995 (N_3995,N_1352,N_2542);
or U3996 (N_3996,N_1777,N_2226);
or U3997 (N_3997,N_2556,N_2773);
nor U3998 (N_3998,N_382,N_2532);
nor U3999 (N_3999,N_1453,N_1048);
nor U4000 (N_4000,N_2623,N_2107);
nor U4001 (N_4001,N_1648,N_1568);
or U4002 (N_4002,N_2057,N_201);
or U4003 (N_4003,N_281,N_1981);
nor U4004 (N_4004,N_2938,N_2084);
nand U4005 (N_4005,N_2271,N_1225);
and U4006 (N_4006,N_919,N_440);
or U4007 (N_4007,N_1066,N_1936);
or U4008 (N_4008,N_2929,N_818);
nor U4009 (N_4009,N_831,N_1286);
nor U4010 (N_4010,N_2222,N_2541);
and U4011 (N_4011,N_2580,N_575);
nand U4012 (N_4012,N_15,N_2297);
and U4013 (N_4013,N_1115,N_1206);
nor U4014 (N_4014,N_1982,N_1308);
nand U4015 (N_4015,N_38,N_1716);
and U4016 (N_4016,N_1070,N_55);
nand U4017 (N_4017,N_1737,N_2884);
and U4018 (N_4018,N_2796,N_369);
and U4019 (N_4019,N_1277,N_2597);
nand U4020 (N_4020,N_2415,N_845);
nor U4021 (N_4021,N_501,N_1640);
nor U4022 (N_4022,N_1959,N_116);
and U4023 (N_4023,N_2896,N_674);
or U4024 (N_4024,N_942,N_659);
or U4025 (N_4025,N_423,N_2257);
nand U4026 (N_4026,N_1537,N_2311);
and U4027 (N_4027,N_266,N_41);
nand U4028 (N_4028,N_2479,N_1147);
or U4029 (N_4029,N_896,N_2762);
nand U4030 (N_4030,N_1040,N_2043);
nor U4031 (N_4031,N_2135,N_2688);
and U4032 (N_4032,N_2471,N_657);
or U4033 (N_4033,N_1309,N_2054);
nand U4034 (N_4034,N_2159,N_1680);
xnor U4035 (N_4035,N_2752,N_2869);
and U4036 (N_4036,N_103,N_2644);
and U4037 (N_4037,N_2370,N_284);
xnor U4038 (N_4038,N_1763,N_2510);
nand U4039 (N_4039,N_1903,N_520);
and U4040 (N_4040,N_1192,N_2689);
and U4041 (N_4041,N_634,N_1148);
nor U4042 (N_4042,N_2777,N_945);
or U4043 (N_4043,N_297,N_2268);
and U4044 (N_4044,N_2155,N_1293);
and U4045 (N_4045,N_1345,N_1774);
and U4046 (N_4046,N_1043,N_2732);
nand U4047 (N_4047,N_2606,N_654);
or U4048 (N_4048,N_1362,N_2012);
or U4049 (N_4049,N_662,N_1641);
and U4050 (N_4050,N_1146,N_506);
nor U4051 (N_4051,N_865,N_307);
nand U4052 (N_4052,N_2820,N_2992);
nor U4053 (N_4053,N_1089,N_934);
or U4054 (N_4054,N_1290,N_1178);
or U4055 (N_4055,N_1326,N_2544);
nand U4056 (N_4056,N_1909,N_950);
nand U4057 (N_4057,N_1480,N_2246);
and U4058 (N_4058,N_1235,N_1424);
nor U4059 (N_4059,N_2528,N_817);
or U4060 (N_4060,N_1583,N_1539);
or U4061 (N_4061,N_1703,N_814);
or U4062 (N_4062,N_2602,N_336);
and U4063 (N_4063,N_2657,N_1934);
and U4064 (N_4064,N_758,N_850);
nor U4065 (N_4065,N_2066,N_1088);
and U4066 (N_4066,N_2583,N_1210);
nor U4067 (N_4067,N_1007,N_2533);
and U4068 (N_4068,N_222,N_2397);
or U4069 (N_4069,N_1780,N_930);
and U4070 (N_4070,N_464,N_1517);
nand U4071 (N_4071,N_1659,N_1806);
or U4072 (N_4072,N_2366,N_2076);
or U4073 (N_4073,N_311,N_2889);
nand U4074 (N_4074,N_1388,N_1356);
and U4075 (N_4075,N_1525,N_663);
nor U4076 (N_4076,N_407,N_1607);
and U4077 (N_4077,N_2133,N_1421);
or U4078 (N_4078,N_1060,N_19);
nor U4079 (N_4079,N_2767,N_2219);
nor U4080 (N_4080,N_1932,N_901);
nand U4081 (N_4081,N_1193,N_151);
nor U4082 (N_4082,N_1217,N_176);
nor U4083 (N_4083,N_2635,N_2915);
or U4084 (N_4084,N_37,N_2617);
and U4085 (N_4085,N_2906,N_1196);
nor U4086 (N_4086,N_2942,N_2485);
nand U4087 (N_4087,N_491,N_986);
nand U4088 (N_4088,N_2663,N_1917);
nor U4089 (N_4089,N_1455,N_773);
or U4090 (N_4090,N_0,N_1994);
nand U4091 (N_4091,N_1616,N_2333);
and U4092 (N_4092,N_2846,N_2091);
nand U4093 (N_4093,N_471,N_2793);
nor U4094 (N_4094,N_1145,N_264);
nor U4095 (N_4095,N_2841,N_1576);
nand U4096 (N_4096,N_2081,N_2707);
nor U4097 (N_4097,N_594,N_2206);
nor U4098 (N_4098,N_406,N_2709);
or U4099 (N_4099,N_460,N_2310);
nand U4100 (N_4100,N_2678,N_754);
nor U4101 (N_4101,N_2332,N_977);
and U4102 (N_4102,N_2797,N_1521);
nand U4103 (N_4103,N_580,N_2292);
nand U4104 (N_4104,N_330,N_2685);
nand U4105 (N_4105,N_2630,N_2843);
nand U4106 (N_4106,N_927,N_76);
nand U4107 (N_4107,N_2481,N_1500);
nor U4108 (N_4108,N_1857,N_2593);
nand U4109 (N_4109,N_1033,N_2151);
or U4110 (N_4110,N_2802,N_2260);
nor U4111 (N_4111,N_2974,N_1770);
or U4112 (N_4112,N_1069,N_998);
nor U4113 (N_4113,N_605,N_2138);
nor U4114 (N_4114,N_280,N_1416);
nand U4115 (N_4115,N_237,N_1700);
and U4116 (N_4116,N_2525,N_2245);
and U4117 (N_4117,N_2314,N_12);
or U4118 (N_4118,N_530,N_1601);
nand U4119 (N_4119,N_358,N_843);
or U4120 (N_4120,N_1828,N_1812);
nand U4121 (N_4121,N_473,N_2161);
or U4122 (N_4122,N_562,N_2893);
and U4123 (N_4123,N_1906,N_849);
or U4124 (N_4124,N_45,N_143);
or U4125 (N_4125,N_1342,N_416);
or U4126 (N_4126,N_2358,N_2930);
or U4127 (N_4127,N_2431,N_1445);
xnor U4128 (N_4128,N_1139,N_795);
nand U4129 (N_4129,N_2444,N_651);
or U4130 (N_4130,N_1531,N_2676);
or U4131 (N_4131,N_1322,N_177);
and U4132 (N_4132,N_1200,N_2113);
nor U4133 (N_4133,N_2984,N_1002);
and U4134 (N_4134,N_1947,N_1785);
and U4135 (N_4135,N_1668,N_1474);
and U4136 (N_4136,N_807,N_1955);
nor U4137 (N_4137,N_2988,N_1176);
and U4138 (N_4138,N_153,N_320);
and U4139 (N_4139,N_2955,N_2924);
xor U4140 (N_4140,N_2546,N_2058);
or U4141 (N_4141,N_488,N_1945);
and U4142 (N_4142,N_1868,N_1055);
or U4143 (N_4143,N_306,N_1826);
nor U4144 (N_4144,N_325,N_35);
nor U4145 (N_4145,N_448,N_343);
nor U4146 (N_4146,N_232,N_976);
nor U4147 (N_4147,N_2997,N_395);
nand U4148 (N_4148,N_1244,N_1973);
or U4149 (N_4149,N_154,N_1958);
nand U4150 (N_4150,N_1964,N_1741);
or U4151 (N_4151,N_2874,N_2237);
nor U4152 (N_4152,N_1091,N_1996);
nor U4153 (N_4153,N_679,N_650);
nor U4154 (N_4154,N_1779,N_915);
and U4155 (N_4155,N_2103,N_2152);
or U4156 (N_4156,N_867,N_2176);
nor U4157 (N_4157,N_793,N_2652);
and U4158 (N_4158,N_1746,N_1579);
nor U4159 (N_4159,N_2770,N_2634);
or U4160 (N_4160,N_1000,N_1673);
nand U4161 (N_4161,N_461,N_948);
nand U4162 (N_4162,N_1767,N_918);
nor U4163 (N_4163,N_2193,N_1987);
or U4164 (N_4164,N_2993,N_747);
and U4165 (N_4165,N_897,N_1734);
and U4166 (N_4166,N_943,N_398);
nand U4167 (N_4167,N_1085,N_1663);
or U4168 (N_4168,N_390,N_2097);
nor U4169 (N_4169,N_2277,N_34);
nand U4170 (N_4170,N_1761,N_2336);
nand U4171 (N_4171,N_764,N_323);
nand U4172 (N_4172,N_2721,N_132);
or U4173 (N_4173,N_779,N_1602);
nand U4174 (N_4174,N_1116,N_1009);
nand U4175 (N_4175,N_532,N_1924);
nand U4176 (N_4176,N_635,N_2041);
nor U4177 (N_4177,N_1626,N_895);
and U4178 (N_4178,N_2830,N_2460);
or U4179 (N_4179,N_271,N_1441);
and U4180 (N_4180,N_1825,N_1671);
nor U4181 (N_4181,N_970,N_465);
nand U4182 (N_4182,N_979,N_664);
or U4183 (N_4183,N_582,N_225);
nor U4184 (N_4184,N_1678,N_926);
or U4185 (N_4185,N_1502,N_1693);
nand U4186 (N_4186,N_1585,N_1519);
and U4187 (N_4187,N_286,N_1622);
or U4188 (N_4188,N_1944,N_1735);
and U4189 (N_4189,N_2177,N_2669);
nor U4190 (N_4190,N_829,N_1062);
nor U4191 (N_4191,N_414,N_51);
or U4192 (N_4192,N_2560,N_711);
and U4193 (N_4193,N_79,N_2719);
nand U4194 (N_4194,N_2971,N_1966);
or U4195 (N_4195,N_1194,N_455);
nand U4196 (N_4196,N_265,N_94);
nand U4197 (N_4197,N_1371,N_1794);
nand U4198 (N_4198,N_1248,N_1050);
and U4199 (N_4199,N_1518,N_887);
nor U4200 (N_4200,N_2946,N_2217);
and U4201 (N_4201,N_1374,N_7);
nor U4202 (N_4202,N_611,N_1041);
and U4203 (N_4203,N_617,N_1633);
nor U4204 (N_4204,N_139,N_65);
nor U4205 (N_4205,N_2253,N_1393);
nand U4206 (N_4206,N_499,N_1674);
nor U4207 (N_4207,N_622,N_2180);
or U4208 (N_4208,N_1969,N_2559);
and U4209 (N_4209,N_2337,N_350);
xor U4210 (N_4210,N_56,N_539);
nor U4211 (N_4211,N_2355,N_740);
nand U4212 (N_4212,N_1289,N_2631);
and U4213 (N_4213,N_378,N_618);
or U4214 (N_4214,N_2204,N_2300);
and U4215 (N_4215,N_1102,N_2441);
and U4216 (N_4216,N_2643,N_1489);
xnor U4217 (N_4217,N_988,N_273);
and U4218 (N_4218,N_439,N_1161);
nor U4219 (N_4219,N_17,N_2263);
nor U4220 (N_4220,N_1970,N_1154);
or U4221 (N_4221,N_2106,N_2416);
or U4222 (N_4222,N_278,N_1817);
or U4223 (N_4223,N_1639,N_1136);
nor U4224 (N_4224,N_497,N_335);
and U4225 (N_4225,N_1935,N_123);
nand U4226 (N_4226,N_873,N_2158);
nand U4227 (N_4227,N_2772,N_129);
or U4228 (N_4228,N_564,N_1365);
and U4229 (N_4229,N_2215,N_2149);
nand U4230 (N_4230,N_2386,N_2378);
nor U4231 (N_4231,N_2588,N_1105);
and U4232 (N_4232,N_1570,N_2857);
or U4233 (N_4233,N_1444,N_2146);
and U4234 (N_4234,N_2650,N_1199);
or U4235 (N_4235,N_1347,N_2854);
or U4236 (N_4236,N_519,N_508);
nand U4237 (N_4237,N_1760,N_714);
or U4238 (N_4238,N_1256,N_1937);
nand U4239 (N_4239,N_2255,N_288);
xor U4240 (N_4240,N_1646,N_2048);
or U4241 (N_4241,N_624,N_1484);
and U4242 (N_4242,N_2488,N_938);
nand U4243 (N_4243,N_1092,N_1394);
and U4244 (N_4244,N_2205,N_2591);
and U4245 (N_4245,N_2443,N_1420);
nor U4246 (N_4246,N_2742,N_1788);
and U4247 (N_4247,N_2778,N_731);
or U4248 (N_4248,N_1946,N_791);
or U4249 (N_4249,N_1736,N_376);
and U4250 (N_4250,N_1354,N_1697);
nor U4251 (N_4251,N_985,N_567);
or U4252 (N_4252,N_380,N_1458);
nand U4253 (N_4253,N_774,N_1327);
and U4254 (N_4254,N_2968,N_2948);
nor U4255 (N_4255,N_1962,N_377);
xnor U4256 (N_4256,N_1409,N_1477);
nor U4257 (N_4257,N_1237,N_1408);
and U4258 (N_4258,N_2587,N_552);
and U4259 (N_4259,N_705,N_1156);
and U4260 (N_4260,N_436,N_1429);
nor U4261 (N_4261,N_2758,N_1839);
nor U4262 (N_4262,N_1389,N_42);
or U4263 (N_4263,N_2529,N_256);
nand U4264 (N_4264,N_686,N_1608);
or U4265 (N_4265,N_2328,N_2775);
or U4266 (N_4266,N_2216,N_2015);
and U4267 (N_4267,N_2051,N_1683);
and U4268 (N_4268,N_2364,N_115);
nor U4269 (N_4269,N_2117,N_876);
nand U4270 (N_4270,N_2540,N_2452);
or U4271 (N_4271,N_1886,N_642);
and U4272 (N_4272,N_1278,N_1792);
nor U4273 (N_4273,N_2166,N_2921);
nand U4274 (N_4274,N_2067,N_2508);
or U4275 (N_4275,N_2190,N_882);
and U4276 (N_4276,N_653,N_2740);
or U4277 (N_4277,N_2273,N_1466);
and U4278 (N_4278,N_526,N_558);
or U4279 (N_4279,N_21,N_208);
and U4280 (N_4280,N_1439,N_127);
and U4281 (N_4281,N_600,N_2815);
nand U4282 (N_4282,N_431,N_1335);
nand U4283 (N_4283,N_1653,N_1915);
or U4284 (N_4284,N_826,N_1188);
or U4285 (N_4285,N_2768,N_258);
or U4286 (N_4286,N_188,N_1684);
or U4287 (N_4287,N_701,N_2575);
nor U4288 (N_4288,N_2318,N_933);
nand U4289 (N_4289,N_621,N_1098);
or U4290 (N_4290,N_2894,N_946);
or U4291 (N_4291,N_680,N_1433);
or U4292 (N_4292,N_202,N_546);
and U4293 (N_4293,N_1247,N_209);
or U4294 (N_4294,N_2115,N_2801);
and U4295 (N_4295,N_866,N_2324);
nand U4296 (N_4296,N_981,N_1372);
nand U4297 (N_4297,N_1711,N_489);
and U4298 (N_4298,N_2995,N_1778);
nor U4299 (N_4299,N_425,N_1061);
nand U4300 (N_4300,N_2450,N_801);
or U4301 (N_4301,N_2534,N_1751);
nand U4302 (N_4302,N_780,N_631);
nand U4303 (N_4303,N_199,N_2026);
and U4304 (N_4304,N_200,N_2862);
nand U4305 (N_4305,N_1472,N_707);
nor U4306 (N_4306,N_122,N_1073);
and U4307 (N_4307,N_326,N_2640);
or U4308 (N_4308,N_1574,N_2373);
nor U4309 (N_4309,N_2751,N_1820);
nand U4310 (N_4310,N_2711,N_693);
nor U4311 (N_4311,N_1563,N_1637);
nor U4312 (N_4312,N_1759,N_1768);
nor U4313 (N_4313,N_1240,N_1239);
nor U4314 (N_4314,N_219,N_205);
nand U4315 (N_4315,N_861,N_543);
nand U4316 (N_4316,N_732,N_2851);
xnor U4317 (N_4317,N_2696,N_2590);
and U4318 (N_4318,N_1877,N_2280);
nand U4319 (N_4319,N_633,N_1764);
or U4320 (N_4320,N_852,N_2774);
or U4321 (N_4321,N_1172,N_463);
and U4322 (N_4322,N_2564,N_450);
nor U4323 (N_4323,N_466,N_1931);
nor U4324 (N_4324,N_1325,N_36);
nand U4325 (N_4325,N_898,N_2447);
and U4326 (N_4326,N_1431,N_1457);
or U4327 (N_4327,N_2121,N_299);
and U4328 (N_4328,N_2907,N_2304);
nor U4329 (N_4329,N_412,N_1403);
nand U4330 (N_4330,N_1756,N_1087);
and U4331 (N_4331,N_2362,N_1280);
or U4332 (N_4332,N_911,N_2400);
and U4333 (N_4333,N_871,N_1867);
nand U4334 (N_4334,N_910,N_309);
or U4335 (N_4335,N_2375,N_1594);
nand U4336 (N_4336,N_2514,N_2899);
and U4337 (N_4337,N_1528,N_1065);
or U4338 (N_4338,N_2798,N_648);
nand U4339 (N_4339,N_393,N_1598);
or U4340 (N_4340,N_1297,N_1710);
or U4341 (N_4341,N_1451,N_2555);
or U4342 (N_4342,N_925,N_351);
and U4343 (N_4343,N_2911,N_2342);
nand U4344 (N_4344,N_833,N_1662);
nand U4345 (N_4345,N_1738,N_2779);
nand U4346 (N_4346,N_2162,N_2876);
or U4347 (N_4347,N_493,N_2203);
nor U4348 (N_4348,N_1850,N_1874);
nor U4349 (N_4349,N_2264,N_794);
nand U4350 (N_4350,N_2250,N_2035);
nand U4351 (N_4351,N_825,N_211);
nand U4352 (N_4352,N_2515,N_149);
xnor U4353 (N_4353,N_2703,N_198);
nor U4354 (N_4354,N_158,N_1620);
and U4355 (N_4355,N_352,N_433);
nor U4356 (N_4356,N_820,N_916);
or U4357 (N_4357,N_1657,N_2947);
nand U4358 (N_4358,N_1865,N_328);
and U4359 (N_4359,N_1730,N_10);
nor U4360 (N_4360,N_2627,N_877);
or U4361 (N_4361,N_1481,N_768);
or U4362 (N_4362,N_1348,N_2468);
nor U4363 (N_4363,N_102,N_2325);
or U4364 (N_4364,N_2877,N_522);
nand U4365 (N_4365,N_454,N_1003);
and U4366 (N_4366,N_136,N_2144);
and U4367 (N_4367,N_1815,N_1249);
or U4368 (N_4368,N_2,N_2100);
nor U4369 (N_4369,N_2462,N_1119);
nand U4370 (N_4370,N_2092,N_70);
nor U4371 (N_4371,N_587,N_206);
or U4372 (N_4372,N_1053,N_1976);
nor U4373 (N_4373,N_2972,N_2746);
or U4374 (N_4374,N_1795,N_420);
and U4375 (N_4375,N_2148,N_2343);
xnor U4376 (N_4376,N_1965,N_235);
nand U4377 (N_4377,N_411,N_2967);
nor U4378 (N_4378,N_337,N_327);
and U4379 (N_4379,N_282,N_2668);
xnor U4380 (N_4380,N_2202,N_2417);
and U4381 (N_4381,N_2718,N_972);
or U4382 (N_4382,N_2800,N_88);
and U4383 (N_4383,N_1831,N_2551);
nor U4384 (N_4384,N_2306,N_2784);
and U4385 (N_4385,N_156,N_606);
and U4386 (N_4386,N_2037,N_2999);
nand U4387 (N_4387,N_1899,N_2785);
nand U4388 (N_4388,N_1397,N_2832);
nor U4389 (N_4389,N_449,N_131);
or U4390 (N_4390,N_2316,N_2979);
or U4391 (N_4391,N_2875,N_2799);
nor U4392 (N_4392,N_1541,N_2632);
or U4393 (N_4393,N_1986,N_1301);
nor U4394 (N_4394,N_1082,N_238);
nand U4395 (N_4395,N_2313,N_1923);
and U4396 (N_4396,N_1843,N_1522);
and U4397 (N_4397,N_857,N_1174);
nor U4398 (N_4398,N_2626,N_1490);
nor U4399 (N_4399,N_2290,N_1134);
nor U4400 (N_4400,N_2123,N_2805);
and U4401 (N_4401,N_800,N_1967);
and U4402 (N_4402,N_1262,N_2932);
and U4403 (N_4403,N_2553,N_1006);
or U4404 (N_4404,N_2068,N_1914);
nand U4405 (N_4405,N_2629,N_1287);
nand U4406 (N_4406,N_2353,N_640);
nor U4407 (N_4407,N_48,N_2446);
and U4408 (N_4408,N_2578,N_2592);
nand U4409 (N_4409,N_163,N_839);
or U4410 (N_4410,N_371,N_1203);
xnor U4411 (N_4411,N_276,N_1111);
or U4412 (N_4412,N_760,N_2980);
and U4413 (N_4413,N_1984,N_2977);
and U4414 (N_4414,N_1880,N_2461);
and U4415 (N_4415,N_1963,N_2686);
xor U4416 (N_4416,N_2270,N_2549);
and U4417 (N_4417,N_545,N_2568);
or U4418 (N_4418,N_444,N_1076);
xor U4419 (N_4419,N_2945,N_1114);
and U4420 (N_4420,N_1383,N_2760);
nor U4421 (N_4421,N_308,N_169);
and U4422 (N_4422,N_1375,N_963);
nor U4423 (N_4423,N_684,N_2536);
and U4424 (N_4424,N_2221,N_2096);
and U4425 (N_4425,N_1083,N_478);
and U4426 (N_4426,N_2414,N_386);
nand U4427 (N_4427,N_1723,N_2482);
nand U4428 (N_4428,N_2537,N_224);
and U4429 (N_4429,N_405,N_2548);
nor U4430 (N_4430,N_2269,N_2241);
and U4431 (N_4431,N_75,N_2965);
and U4432 (N_4432,N_112,N_1905);
or U4433 (N_4433,N_2670,N_540);
nand U4434 (N_4434,N_2225,N_342);
nand U4435 (N_4435,N_2456,N_786);
or U4436 (N_4436,N_2842,N_2708);
nor U4437 (N_4437,N_1543,N_2335);
nor U4438 (N_4438,N_1267,N_1275);
nand U4439 (N_4439,N_1744,N_647);
nor U4440 (N_4440,N_523,N_2396);
and U4441 (N_4441,N_2178,N_381);
or U4442 (N_4442,N_191,N_413);
nor U4443 (N_4443,N_2459,N_2085);
nor U4444 (N_4444,N_2866,N_8);
nand U4445 (N_4445,N_2409,N_1572);
and U4446 (N_4446,N_1313,N_1359);
xor U4447 (N_4447,N_1642,N_1184);
nand U4448 (N_4448,N_329,N_2812);
nor U4449 (N_4449,N_1021,N_832);
or U4450 (N_4450,N_2033,N_2717);
nor U4451 (N_4451,N_1651,N_2497);
and U4452 (N_4452,N_738,N_1264);
or U4453 (N_4453,N_1796,N_2853);
or U4454 (N_4454,N_157,N_1954);
nand U4455 (N_4455,N_726,N_968);
nand U4456 (N_4456,N_1242,N_2628);
or U4457 (N_4457,N_2291,N_1922);
and U4458 (N_4458,N_2448,N_424);
nand U4459 (N_4459,N_1554,N_920);
or U4460 (N_4460,N_2867,N_2019);
nor U4461 (N_4461,N_2716,N_899);
nand U4462 (N_4462,N_438,N_33);
nor U4463 (N_4463,N_2126,N_2381);
or U4464 (N_4464,N_2879,N_1052);
nand U4465 (N_4465,N_1927,N_476);
nor U4466 (N_4466,N_510,N_1577);
nor U4467 (N_4467,N_1492,N_2127);
nor U4468 (N_4468,N_980,N_771);
or U4469 (N_4469,N_1108,N_2281);
and U4470 (N_4470,N_1074,N_1078);
nor U4471 (N_4471,N_989,N_1685);
nor U4472 (N_4472,N_289,N_1020);
or U4473 (N_4473,N_78,N_1514);
nand U4474 (N_4474,N_1412,N_1766);
and U4475 (N_4475,N_1605,N_2480);
or U4476 (N_4476,N_2200,N_187);
nand U4477 (N_4477,N_2679,N_2582);
nor U4478 (N_4478,N_2831,N_964);
or U4479 (N_4479,N_184,N_1435);
and U4480 (N_4480,N_2384,N_1380);
nand U4481 (N_4481,N_2228,N_2731);
and U4482 (N_4482,N_4,N_2349);
nand U4483 (N_4483,N_1486,N_1650);
and U4484 (N_4484,N_2363,N_2382);
or U4485 (N_4485,N_699,N_1580);
nor U4486 (N_4486,N_1507,N_982);
nand U4487 (N_4487,N_2745,N_341);
or U4488 (N_4488,N_1141,N_1645);
nand U4489 (N_4489,N_1182,N_2074);
and U4490 (N_4490,N_304,N_974);
nand U4491 (N_4491,N_1687,N_1548);
nor U4492 (N_4492,N_2954,N_1872);
and U4493 (N_4493,N_2818,N_1556);
nand U4494 (N_4494,N_1181,N_204);
or U4495 (N_4495,N_2581,N_1276);
nand U4496 (N_4496,N_73,N_548);
nand U4497 (N_4497,N_1384,N_2305);
nand U4498 (N_4498,N_1854,N_2976);
and U4499 (N_4499,N_864,N_2317);
and U4500 (N_4500,N_23,N_815);
and U4501 (N_4501,N_547,N_2779);
or U4502 (N_4502,N_1862,N_1851);
nor U4503 (N_4503,N_2449,N_459);
or U4504 (N_4504,N_1147,N_1451);
and U4505 (N_4505,N_2400,N_1518);
xnor U4506 (N_4506,N_1273,N_1275);
nor U4507 (N_4507,N_2607,N_1144);
and U4508 (N_4508,N_1025,N_1380);
nand U4509 (N_4509,N_408,N_765);
and U4510 (N_4510,N_1323,N_952);
or U4511 (N_4511,N_1332,N_2311);
and U4512 (N_4512,N_173,N_1780);
nand U4513 (N_4513,N_1717,N_1427);
or U4514 (N_4514,N_545,N_2319);
and U4515 (N_4515,N_1712,N_88);
nor U4516 (N_4516,N_2873,N_2165);
nor U4517 (N_4517,N_2978,N_2877);
nor U4518 (N_4518,N_2832,N_907);
and U4519 (N_4519,N_1620,N_2023);
nand U4520 (N_4520,N_2079,N_2945);
or U4521 (N_4521,N_338,N_1038);
nor U4522 (N_4522,N_2209,N_70);
nand U4523 (N_4523,N_2627,N_2748);
or U4524 (N_4524,N_1413,N_2590);
nor U4525 (N_4525,N_602,N_2176);
or U4526 (N_4526,N_526,N_1591);
nor U4527 (N_4527,N_181,N_1969);
nand U4528 (N_4528,N_2401,N_2605);
nor U4529 (N_4529,N_615,N_2711);
and U4530 (N_4530,N_2212,N_192);
and U4531 (N_4531,N_1227,N_27);
nor U4532 (N_4532,N_1831,N_2699);
nand U4533 (N_4533,N_1105,N_1061);
nand U4534 (N_4534,N_2946,N_1892);
or U4535 (N_4535,N_242,N_308);
nand U4536 (N_4536,N_2239,N_491);
or U4537 (N_4537,N_124,N_1621);
or U4538 (N_4538,N_1073,N_555);
and U4539 (N_4539,N_900,N_637);
and U4540 (N_4540,N_594,N_1569);
or U4541 (N_4541,N_1318,N_801);
or U4542 (N_4542,N_2727,N_386);
nand U4543 (N_4543,N_1280,N_2023);
and U4544 (N_4544,N_309,N_548);
nor U4545 (N_4545,N_2193,N_151);
nand U4546 (N_4546,N_61,N_366);
nand U4547 (N_4547,N_2182,N_1855);
or U4548 (N_4548,N_2277,N_1313);
nand U4549 (N_4549,N_1656,N_1736);
nor U4550 (N_4550,N_209,N_168);
nor U4551 (N_4551,N_2199,N_2249);
nor U4552 (N_4552,N_2594,N_2445);
nor U4553 (N_4553,N_650,N_2057);
nor U4554 (N_4554,N_376,N_644);
nor U4555 (N_4555,N_698,N_2457);
nor U4556 (N_4556,N_1463,N_1442);
or U4557 (N_4557,N_705,N_1844);
or U4558 (N_4558,N_1571,N_23);
or U4559 (N_4559,N_2064,N_952);
nand U4560 (N_4560,N_2486,N_554);
nor U4561 (N_4561,N_1419,N_1015);
and U4562 (N_4562,N_697,N_2908);
or U4563 (N_4563,N_2084,N_1296);
nand U4564 (N_4564,N_2526,N_651);
nand U4565 (N_4565,N_2571,N_1069);
nand U4566 (N_4566,N_2610,N_1362);
or U4567 (N_4567,N_483,N_2375);
and U4568 (N_4568,N_363,N_1145);
and U4569 (N_4569,N_807,N_1879);
nand U4570 (N_4570,N_1324,N_2561);
or U4571 (N_4571,N_2950,N_2656);
or U4572 (N_4572,N_293,N_1624);
and U4573 (N_4573,N_1385,N_2116);
and U4574 (N_4574,N_2175,N_1025);
or U4575 (N_4575,N_1061,N_1519);
xnor U4576 (N_4576,N_62,N_2673);
or U4577 (N_4577,N_2526,N_489);
and U4578 (N_4578,N_2237,N_1780);
or U4579 (N_4579,N_1955,N_1966);
nor U4580 (N_4580,N_1443,N_1676);
nor U4581 (N_4581,N_566,N_470);
or U4582 (N_4582,N_1092,N_724);
nor U4583 (N_4583,N_2981,N_717);
and U4584 (N_4584,N_262,N_751);
nand U4585 (N_4585,N_695,N_157);
and U4586 (N_4586,N_1832,N_362);
and U4587 (N_4587,N_1160,N_2125);
and U4588 (N_4588,N_9,N_1931);
nor U4589 (N_4589,N_1506,N_838);
or U4590 (N_4590,N_1483,N_2486);
and U4591 (N_4591,N_877,N_1407);
nor U4592 (N_4592,N_1511,N_1694);
nand U4593 (N_4593,N_2174,N_678);
or U4594 (N_4594,N_1637,N_2918);
or U4595 (N_4595,N_2142,N_2746);
or U4596 (N_4596,N_369,N_1434);
or U4597 (N_4597,N_2630,N_1083);
nor U4598 (N_4598,N_2859,N_587);
nand U4599 (N_4599,N_100,N_2426);
nor U4600 (N_4600,N_443,N_820);
nand U4601 (N_4601,N_2717,N_1981);
nand U4602 (N_4602,N_53,N_2166);
nor U4603 (N_4603,N_2615,N_822);
or U4604 (N_4604,N_1135,N_1917);
nand U4605 (N_4605,N_1963,N_1983);
and U4606 (N_4606,N_41,N_2540);
or U4607 (N_4607,N_1188,N_87);
nor U4608 (N_4608,N_836,N_1061);
and U4609 (N_4609,N_2136,N_1879);
or U4610 (N_4610,N_2375,N_211);
or U4611 (N_4611,N_868,N_962);
nand U4612 (N_4612,N_1423,N_1440);
nor U4613 (N_4613,N_1814,N_887);
and U4614 (N_4614,N_668,N_1898);
or U4615 (N_4615,N_1127,N_2669);
or U4616 (N_4616,N_1959,N_1110);
and U4617 (N_4617,N_2628,N_241);
or U4618 (N_4618,N_1962,N_1489);
or U4619 (N_4619,N_588,N_519);
nand U4620 (N_4620,N_175,N_2888);
xor U4621 (N_4621,N_185,N_1155);
and U4622 (N_4622,N_1457,N_291);
and U4623 (N_4623,N_1139,N_2968);
xor U4624 (N_4624,N_1646,N_255);
or U4625 (N_4625,N_1417,N_44);
and U4626 (N_4626,N_230,N_1556);
nor U4627 (N_4627,N_1023,N_1224);
and U4628 (N_4628,N_2668,N_1384);
nor U4629 (N_4629,N_68,N_1827);
and U4630 (N_4630,N_2185,N_304);
nor U4631 (N_4631,N_1961,N_366);
nand U4632 (N_4632,N_75,N_2453);
nand U4633 (N_4633,N_1636,N_1557);
and U4634 (N_4634,N_863,N_72);
nor U4635 (N_4635,N_891,N_2710);
nor U4636 (N_4636,N_297,N_2945);
or U4637 (N_4637,N_2553,N_2372);
nor U4638 (N_4638,N_1899,N_238);
or U4639 (N_4639,N_2519,N_303);
nand U4640 (N_4640,N_720,N_1797);
or U4641 (N_4641,N_1437,N_2019);
and U4642 (N_4642,N_14,N_2628);
nor U4643 (N_4643,N_2549,N_2908);
or U4644 (N_4644,N_2860,N_2761);
xor U4645 (N_4645,N_2348,N_2719);
and U4646 (N_4646,N_253,N_378);
or U4647 (N_4647,N_206,N_114);
nand U4648 (N_4648,N_1899,N_1141);
or U4649 (N_4649,N_1693,N_610);
and U4650 (N_4650,N_786,N_680);
or U4651 (N_4651,N_92,N_2353);
and U4652 (N_4652,N_1642,N_642);
nand U4653 (N_4653,N_988,N_771);
nand U4654 (N_4654,N_2764,N_2518);
nor U4655 (N_4655,N_887,N_2644);
nand U4656 (N_4656,N_799,N_2821);
nor U4657 (N_4657,N_2025,N_2351);
nor U4658 (N_4658,N_1386,N_62);
and U4659 (N_4659,N_2494,N_149);
nor U4660 (N_4660,N_2542,N_1948);
nand U4661 (N_4661,N_2748,N_2927);
nor U4662 (N_4662,N_601,N_1763);
or U4663 (N_4663,N_1560,N_730);
or U4664 (N_4664,N_2127,N_2553);
nor U4665 (N_4665,N_1397,N_2289);
nand U4666 (N_4666,N_1318,N_1257);
nor U4667 (N_4667,N_712,N_532);
nand U4668 (N_4668,N_816,N_2121);
and U4669 (N_4669,N_2,N_743);
nand U4670 (N_4670,N_1249,N_2320);
nand U4671 (N_4671,N_2548,N_1968);
nor U4672 (N_4672,N_280,N_810);
nand U4673 (N_4673,N_1863,N_1241);
nor U4674 (N_4674,N_471,N_1924);
or U4675 (N_4675,N_73,N_2830);
xor U4676 (N_4676,N_1515,N_2041);
and U4677 (N_4677,N_2598,N_207);
and U4678 (N_4678,N_1234,N_114);
or U4679 (N_4679,N_787,N_770);
nor U4680 (N_4680,N_1094,N_2009);
and U4681 (N_4681,N_2727,N_2431);
nand U4682 (N_4682,N_56,N_572);
or U4683 (N_4683,N_400,N_1848);
nor U4684 (N_4684,N_454,N_1851);
and U4685 (N_4685,N_2931,N_514);
or U4686 (N_4686,N_821,N_712);
or U4687 (N_4687,N_2779,N_871);
or U4688 (N_4688,N_233,N_531);
nand U4689 (N_4689,N_2568,N_101);
nor U4690 (N_4690,N_1143,N_2125);
and U4691 (N_4691,N_2046,N_2925);
or U4692 (N_4692,N_991,N_2392);
nand U4693 (N_4693,N_169,N_323);
or U4694 (N_4694,N_879,N_2802);
nand U4695 (N_4695,N_1134,N_531);
nor U4696 (N_4696,N_1059,N_341);
or U4697 (N_4697,N_1679,N_619);
and U4698 (N_4698,N_1184,N_2229);
nor U4699 (N_4699,N_697,N_172);
nand U4700 (N_4700,N_1675,N_867);
nand U4701 (N_4701,N_1727,N_352);
and U4702 (N_4702,N_332,N_1118);
nor U4703 (N_4703,N_1279,N_64);
nor U4704 (N_4704,N_397,N_1339);
nand U4705 (N_4705,N_424,N_2101);
nor U4706 (N_4706,N_1354,N_1897);
and U4707 (N_4707,N_802,N_582);
nand U4708 (N_4708,N_1010,N_2835);
nand U4709 (N_4709,N_828,N_1639);
nand U4710 (N_4710,N_2278,N_1353);
and U4711 (N_4711,N_2296,N_2153);
nor U4712 (N_4712,N_2172,N_552);
nand U4713 (N_4713,N_2144,N_1905);
or U4714 (N_4714,N_269,N_1389);
xor U4715 (N_4715,N_2345,N_577);
or U4716 (N_4716,N_1989,N_1586);
nand U4717 (N_4717,N_1430,N_1074);
and U4718 (N_4718,N_2156,N_1493);
nand U4719 (N_4719,N_511,N_840);
nand U4720 (N_4720,N_2491,N_1245);
or U4721 (N_4721,N_2714,N_2127);
nand U4722 (N_4722,N_2324,N_1099);
and U4723 (N_4723,N_327,N_2393);
or U4724 (N_4724,N_1677,N_2593);
and U4725 (N_4725,N_1358,N_2224);
nor U4726 (N_4726,N_1123,N_594);
or U4727 (N_4727,N_874,N_1610);
nor U4728 (N_4728,N_1857,N_2321);
nor U4729 (N_4729,N_767,N_1592);
nor U4730 (N_4730,N_2115,N_999);
nor U4731 (N_4731,N_2608,N_867);
and U4732 (N_4732,N_1758,N_142);
nor U4733 (N_4733,N_2155,N_177);
or U4734 (N_4734,N_1762,N_2655);
or U4735 (N_4735,N_1093,N_741);
nand U4736 (N_4736,N_121,N_2662);
nor U4737 (N_4737,N_1261,N_2672);
nor U4738 (N_4738,N_2125,N_1251);
nand U4739 (N_4739,N_1061,N_2579);
or U4740 (N_4740,N_1235,N_2300);
and U4741 (N_4741,N_1951,N_1488);
nand U4742 (N_4742,N_1404,N_739);
or U4743 (N_4743,N_931,N_2750);
nor U4744 (N_4744,N_2331,N_62);
and U4745 (N_4745,N_1269,N_2509);
xnor U4746 (N_4746,N_140,N_72);
and U4747 (N_4747,N_970,N_1199);
and U4748 (N_4748,N_1234,N_2724);
nand U4749 (N_4749,N_658,N_1839);
nor U4750 (N_4750,N_2300,N_2920);
nand U4751 (N_4751,N_561,N_882);
nand U4752 (N_4752,N_785,N_1456);
or U4753 (N_4753,N_167,N_720);
nor U4754 (N_4754,N_1089,N_2967);
or U4755 (N_4755,N_2437,N_488);
or U4756 (N_4756,N_922,N_873);
and U4757 (N_4757,N_662,N_2172);
nand U4758 (N_4758,N_1612,N_58);
or U4759 (N_4759,N_2872,N_1899);
and U4760 (N_4760,N_915,N_235);
nand U4761 (N_4761,N_2854,N_222);
nand U4762 (N_4762,N_917,N_225);
and U4763 (N_4763,N_1321,N_2709);
or U4764 (N_4764,N_876,N_2034);
nor U4765 (N_4765,N_2262,N_1180);
nand U4766 (N_4766,N_1063,N_159);
or U4767 (N_4767,N_2520,N_2313);
and U4768 (N_4768,N_1558,N_267);
xor U4769 (N_4769,N_1807,N_1790);
and U4770 (N_4770,N_846,N_2550);
nand U4771 (N_4771,N_2316,N_1132);
nand U4772 (N_4772,N_638,N_1716);
or U4773 (N_4773,N_1191,N_130);
or U4774 (N_4774,N_2992,N_1603);
nor U4775 (N_4775,N_785,N_767);
nand U4776 (N_4776,N_1444,N_92);
or U4777 (N_4777,N_169,N_586);
and U4778 (N_4778,N_83,N_2176);
and U4779 (N_4779,N_1113,N_2770);
or U4780 (N_4780,N_479,N_113);
nand U4781 (N_4781,N_116,N_1631);
nand U4782 (N_4782,N_2202,N_1003);
nand U4783 (N_4783,N_1801,N_2624);
nand U4784 (N_4784,N_649,N_1663);
xor U4785 (N_4785,N_1505,N_1673);
and U4786 (N_4786,N_2205,N_1383);
or U4787 (N_4787,N_1251,N_987);
or U4788 (N_4788,N_303,N_2311);
nand U4789 (N_4789,N_2061,N_2724);
and U4790 (N_4790,N_1576,N_2865);
nand U4791 (N_4791,N_1770,N_1519);
or U4792 (N_4792,N_354,N_1612);
nand U4793 (N_4793,N_553,N_1653);
nand U4794 (N_4794,N_1853,N_607);
nor U4795 (N_4795,N_1220,N_2652);
and U4796 (N_4796,N_779,N_2969);
nand U4797 (N_4797,N_1034,N_1135);
and U4798 (N_4798,N_1712,N_886);
nor U4799 (N_4799,N_654,N_2262);
nor U4800 (N_4800,N_1862,N_2715);
nor U4801 (N_4801,N_2986,N_682);
nor U4802 (N_4802,N_2261,N_1321);
nor U4803 (N_4803,N_2864,N_492);
nand U4804 (N_4804,N_1505,N_338);
or U4805 (N_4805,N_396,N_1815);
or U4806 (N_4806,N_441,N_718);
nor U4807 (N_4807,N_2338,N_2330);
nor U4808 (N_4808,N_1226,N_1715);
or U4809 (N_4809,N_1424,N_500);
and U4810 (N_4810,N_2864,N_2370);
nor U4811 (N_4811,N_2801,N_2356);
or U4812 (N_4812,N_1415,N_849);
and U4813 (N_4813,N_2558,N_1018);
nor U4814 (N_4814,N_1911,N_2801);
nand U4815 (N_4815,N_997,N_2399);
nor U4816 (N_4816,N_104,N_30);
nor U4817 (N_4817,N_1952,N_134);
and U4818 (N_4818,N_85,N_376);
or U4819 (N_4819,N_2748,N_489);
or U4820 (N_4820,N_476,N_330);
nor U4821 (N_4821,N_30,N_929);
nor U4822 (N_4822,N_1484,N_371);
or U4823 (N_4823,N_1166,N_2649);
or U4824 (N_4824,N_1363,N_1015);
and U4825 (N_4825,N_2417,N_2159);
nand U4826 (N_4826,N_155,N_2688);
and U4827 (N_4827,N_969,N_687);
nor U4828 (N_4828,N_519,N_1231);
and U4829 (N_4829,N_2313,N_1239);
or U4830 (N_4830,N_2800,N_2998);
xnor U4831 (N_4831,N_754,N_2596);
and U4832 (N_4832,N_2767,N_2294);
nand U4833 (N_4833,N_2929,N_472);
or U4834 (N_4834,N_2427,N_379);
or U4835 (N_4835,N_2516,N_2966);
or U4836 (N_4836,N_2976,N_338);
nand U4837 (N_4837,N_1402,N_1415);
nor U4838 (N_4838,N_636,N_235);
and U4839 (N_4839,N_724,N_34);
nand U4840 (N_4840,N_2855,N_2023);
or U4841 (N_4841,N_1714,N_2029);
and U4842 (N_4842,N_2362,N_495);
nor U4843 (N_4843,N_353,N_1403);
and U4844 (N_4844,N_1573,N_1896);
nor U4845 (N_4845,N_405,N_2926);
or U4846 (N_4846,N_1951,N_179);
nor U4847 (N_4847,N_1542,N_2973);
nand U4848 (N_4848,N_65,N_1382);
and U4849 (N_4849,N_2602,N_1034);
or U4850 (N_4850,N_240,N_1498);
or U4851 (N_4851,N_2842,N_2031);
nor U4852 (N_4852,N_1470,N_2697);
nand U4853 (N_4853,N_2119,N_270);
nor U4854 (N_4854,N_669,N_2404);
nand U4855 (N_4855,N_2388,N_2800);
nand U4856 (N_4856,N_2516,N_1533);
nor U4857 (N_4857,N_2804,N_759);
nand U4858 (N_4858,N_2123,N_730);
nand U4859 (N_4859,N_1963,N_34);
nor U4860 (N_4860,N_718,N_1511);
nand U4861 (N_4861,N_932,N_981);
and U4862 (N_4862,N_2387,N_1302);
or U4863 (N_4863,N_1949,N_2690);
nor U4864 (N_4864,N_2743,N_2426);
and U4865 (N_4865,N_816,N_1564);
and U4866 (N_4866,N_1870,N_388);
nor U4867 (N_4867,N_2731,N_1081);
nor U4868 (N_4868,N_60,N_2515);
nor U4869 (N_4869,N_2597,N_534);
nor U4870 (N_4870,N_388,N_2837);
nand U4871 (N_4871,N_2352,N_966);
nand U4872 (N_4872,N_2870,N_1783);
nor U4873 (N_4873,N_438,N_2776);
nor U4874 (N_4874,N_220,N_2826);
nand U4875 (N_4875,N_1828,N_1516);
nor U4876 (N_4876,N_2560,N_854);
or U4877 (N_4877,N_1651,N_120);
nor U4878 (N_4878,N_2130,N_1526);
nand U4879 (N_4879,N_2461,N_1442);
nand U4880 (N_4880,N_1392,N_1597);
or U4881 (N_4881,N_963,N_1975);
and U4882 (N_4882,N_1539,N_2177);
nand U4883 (N_4883,N_2687,N_2552);
or U4884 (N_4884,N_1636,N_652);
nand U4885 (N_4885,N_173,N_818);
or U4886 (N_4886,N_1840,N_2469);
nand U4887 (N_4887,N_2749,N_2793);
xnor U4888 (N_4888,N_1031,N_1513);
nand U4889 (N_4889,N_2899,N_1419);
or U4890 (N_4890,N_491,N_964);
and U4891 (N_4891,N_1878,N_317);
or U4892 (N_4892,N_531,N_1816);
nand U4893 (N_4893,N_2524,N_642);
nor U4894 (N_4894,N_2867,N_1481);
and U4895 (N_4895,N_2418,N_17);
or U4896 (N_4896,N_1248,N_1322);
nand U4897 (N_4897,N_2908,N_2135);
and U4898 (N_4898,N_1799,N_2481);
nand U4899 (N_4899,N_2046,N_2225);
xnor U4900 (N_4900,N_86,N_1835);
nor U4901 (N_4901,N_2425,N_1640);
or U4902 (N_4902,N_2805,N_1873);
nand U4903 (N_4903,N_552,N_2416);
or U4904 (N_4904,N_1664,N_721);
and U4905 (N_4905,N_335,N_1701);
nor U4906 (N_4906,N_317,N_2358);
or U4907 (N_4907,N_2513,N_555);
nand U4908 (N_4908,N_2356,N_2075);
or U4909 (N_4909,N_875,N_2913);
and U4910 (N_4910,N_2363,N_2786);
nor U4911 (N_4911,N_2647,N_264);
nor U4912 (N_4912,N_1960,N_1523);
nand U4913 (N_4913,N_1392,N_213);
nand U4914 (N_4914,N_1369,N_2122);
and U4915 (N_4915,N_1893,N_2712);
nor U4916 (N_4916,N_2487,N_523);
nand U4917 (N_4917,N_2370,N_1615);
nand U4918 (N_4918,N_1455,N_2599);
and U4919 (N_4919,N_2891,N_1795);
or U4920 (N_4920,N_2084,N_2);
nor U4921 (N_4921,N_210,N_2154);
and U4922 (N_4922,N_748,N_2478);
nor U4923 (N_4923,N_597,N_2515);
nand U4924 (N_4924,N_959,N_2636);
nor U4925 (N_4925,N_1182,N_36);
and U4926 (N_4926,N_793,N_1914);
and U4927 (N_4927,N_515,N_205);
and U4928 (N_4928,N_2972,N_2031);
and U4929 (N_4929,N_1472,N_1777);
nor U4930 (N_4930,N_2846,N_1569);
nor U4931 (N_4931,N_420,N_1506);
and U4932 (N_4932,N_838,N_234);
nor U4933 (N_4933,N_2278,N_1955);
and U4934 (N_4934,N_2316,N_2732);
nor U4935 (N_4935,N_2805,N_2377);
or U4936 (N_4936,N_2201,N_1122);
and U4937 (N_4937,N_2188,N_1083);
nand U4938 (N_4938,N_2221,N_2201);
and U4939 (N_4939,N_631,N_1259);
nor U4940 (N_4940,N_2955,N_380);
or U4941 (N_4941,N_530,N_393);
nand U4942 (N_4942,N_360,N_2087);
and U4943 (N_4943,N_2130,N_1551);
or U4944 (N_4944,N_1948,N_2233);
or U4945 (N_4945,N_2236,N_206);
or U4946 (N_4946,N_2295,N_1496);
or U4947 (N_4947,N_648,N_1226);
nor U4948 (N_4948,N_1070,N_1399);
and U4949 (N_4949,N_933,N_2508);
xnor U4950 (N_4950,N_1168,N_2182);
nor U4951 (N_4951,N_2820,N_2996);
and U4952 (N_4952,N_2140,N_211);
or U4953 (N_4953,N_376,N_766);
nand U4954 (N_4954,N_649,N_2056);
nor U4955 (N_4955,N_626,N_103);
and U4956 (N_4956,N_744,N_546);
nand U4957 (N_4957,N_1497,N_875);
nand U4958 (N_4958,N_751,N_2620);
nor U4959 (N_4959,N_292,N_1132);
and U4960 (N_4960,N_1640,N_1921);
nand U4961 (N_4961,N_791,N_355);
nor U4962 (N_4962,N_736,N_1407);
nor U4963 (N_4963,N_2303,N_2396);
nor U4964 (N_4964,N_233,N_2677);
nor U4965 (N_4965,N_307,N_1196);
and U4966 (N_4966,N_765,N_2383);
nor U4967 (N_4967,N_1353,N_2311);
or U4968 (N_4968,N_1867,N_2485);
or U4969 (N_4969,N_1217,N_2064);
nor U4970 (N_4970,N_567,N_1495);
or U4971 (N_4971,N_669,N_926);
or U4972 (N_4972,N_394,N_551);
or U4973 (N_4973,N_2025,N_2236);
or U4974 (N_4974,N_31,N_2262);
and U4975 (N_4975,N_2809,N_2061);
or U4976 (N_4976,N_2449,N_1929);
nand U4977 (N_4977,N_2522,N_2749);
nor U4978 (N_4978,N_448,N_853);
nor U4979 (N_4979,N_1993,N_224);
nand U4980 (N_4980,N_1435,N_2354);
nor U4981 (N_4981,N_2468,N_721);
and U4982 (N_4982,N_1074,N_1482);
or U4983 (N_4983,N_130,N_837);
nand U4984 (N_4984,N_2502,N_2008);
and U4985 (N_4985,N_1518,N_2937);
or U4986 (N_4986,N_1594,N_1790);
nor U4987 (N_4987,N_7,N_2553);
or U4988 (N_4988,N_1370,N_2913);
nand U4989 (N_4989,N_1384,N_2218);
nor U4990 (N_4990,N_1244,N_1825);
and U4991 (N_4991,N_108,N_323);
and U4992 (N_4992,N_827,N_180);
or U4993 (N_4993,N_776,N_1853);
or U4994 (N_4994,N_2973,N_1208);
nand U4995 (N_4995,N_2029,N_2711);
nand U4996 (N_4996,N_1041,N_2486);
nor U4997 (N_4997,N_1502,N_1600);
nand U4998 (N_4998,N_2278,N_2625);
or U4999 (N_4999,N_2227,N_1113);
and U5000 (N_5000,N_2371,N_2212);
and U5001 (N_5001,N_581,N_2048);
nand U5002 (N_5002,N_1031,N_671);
nand U5003 (N_5003,N_1014,N_672);
or U5004 (N_5004,N_2290,N_2961);
nand U5005 (N_5005,N_141,N_1339);
nor U5006 (N_5006,N_1313,N_2290);
nand U5007 (N_5007,N_2797,N_1930);
and U5008 (N_5008,N_354,N_1054);
xor U5009 (N_5009,N_2556,N_2220);
and U5010 (N_5010,N_2402,N_107);
nor U5011 (N_5011,N_1567,N_1378);
nand U5012 (N_5012,N_2078,N_576);
nor U5013 (N_5013,N_2446,N_2224);
or U5014 (N_5014,N_1299,N_1242);
nor U5015 (N_5015,N_498,N_1760);
and U5016 (N_5016,N_26,N_1192);
nand U5017 (N_5017,N_1184,N_263);
or U5018 (N_5018,N_2911,N_1560);
nor U5019 (N_5019,N_295,N_2569);
nor U5020 (N_5020,N_2924,N_2773);
nand U5021 (N_5021,N_2373,N_410);
or U5022 (N_5022,N_941,N_764);
and U5023 (N_5023,N_1981,N_9);
nor U5024 (N_5024,N_2775,N_2112);
and U5025 (N_5025,N_2118,N_2317);
nand U5026 (N_5026,N_1319,N_1432);
nand U5027 (N_5027,N_175,N_1277);
xnor U5028 (N_5028,N_605,N_2079);
nor U5029 (N_5029,N_2187,N_2998);
nand U5030 (N_5030,N_1465,N_626);
or U5031 (N_5031,N_2142,N_325);
nand U5032 (N_5032,N_1084,N_2260);
and U5033 (N_5033,N_773,N_2255);
nor U5034 (N_5034,N_1658,N_2630);
xor U5035 (N_5035,N_1023,N_1795);
nor U5036 (N_5036,N_1087,N_1489);
nand U5037 (N_5037,N_2825,N_2782);
nand U5038 (N_5038,N_2480,N_1337);
and U5039 (N_5039,N_1945,N_1248);
and U5040 (N_5040,N_2233,N_84);
nand U5041 (N_5041,N_1082,N_1157);
or U5042 (N_5042,N_1117,N_1433);
or U5043 (N_5043,N_1899,N_1409);
nor U5044 (N_5044,N_1424,N_1134);
nand U5045 (N_5045,N_644,N_2459);
or U5046 (N_5046,N_1646,N_2188);
nor U5047 (N_5047,N_2243,N_178);
nand U5048 (N_5048,N_2102,N_1563);
nor U5049 (N_5049,N_2020,N_819);
or U5050 (N_5050,N_2669,N_75);
and U5051 (N_5051,N_1227,N_1870);
nand U5052 (N_5052,N_391,N_467);
and U5053 (N_5053,N_31,N_1915);
nand U5054 (N_5054,N_1393,N_1964);
nand U5055 (N_5055,N_460,N_2550);
nor U5056 (N_5056,N_798,N_1621);
xnor U5057 (N_5057,N_1,N_2007);
nor U5058 (N_5058,N_2657,N_467);
and U5059 (N_5059,N_2597,N_578);
nor U5060 (N_5060,N_2462,N_3);
nor U5061 (N_5061,N_1238,N_769);
nand U5062 (N_5062,N_1746,N_809);
and U5063 (N_5063,N_1871,N_1085);
nand U5064 (N_5064,N_132,N_2112);
nand U5065 (N_5065,N_2051,N_133);
nand U5066 (N_5066,N_1758,N_2457);
nor U5067 (N_5067,N_1,N_2844);
nor U5068 (N_5068,N_502,N_1449);
nor U5069 (N_5069,N_276,N_2894);
and U5070 (N_5070,N_2937,N_1711);
nand U5071 (N_5071,N_1819,N_638);
nand U5072 (N_5072,N_978,N_2684);
nand U5073 (N_5073,N_141,N_449);
nor U5074 (N_5074,N_651,N_2098);
and U5075 (N_5075,N_865,N_1411);
nor U5076 (N_5076,N_615,N_384);
nand U5077 (N_5077,N_1326,N_1671);
and U5078 (N_5078,N_211,N_1961);
nor U5079 (N_5079,N_1096,N_1215);
nand U5080 (N_5080,N_1913,N_277);
nor U5081 (N_5081,N_82,N_2010);
nor U5082 (N_5082,N_2581,N_335);
nor U5083 (N_5083,N_2173,N_772);
nor U5084 (N_5084,N_1287,N_1793);
nand U5085 (N_5085,N_1276,N_1422);
nand U5086 (N_5086,N_887,N_2434);
nor U5087 (N_5087,N_1899,N_125);
or U5088 (N_5088,N_1161,N_276);
nor U5089 (N_5089,N_103,N_2627);
or U5090 (N_5090,N_200,N_1858);
nand U5091 (N_5091,N_1792,N_812);
nand U5092 (N_5092,N_1751,N_2042);
and U5093 (N_5093,N_1441,N_111);
or U5094 (N_5094,N_1221,N_1209);
or U5095 (N_5095,N_1687,N_341);
and U5096 (N_5096,N_2341,N_132);
nand U5097 (N_5097,N_1126,N_1338);
and U5098 (N_5098,N_42,N_2875);
xnor U5099 (N_5099,N_982,N_143);
nor U5100 (N_5100,N_716,N_827);
or U5101 (N_5101,N_1504,N_1206);
and U5102 (N_5102,N_947,N_569);
or U5103 (N_5103,N_53,N_2705);
or U5104 (N_5104,N_1997,N_2930);
nand U5105 (N_5105,N_1705,N_1314);
or U5106 (N_5106,N_1598,N_144);
and U5107 (N_5107,N_2766,N_2102);
or U5108 (N_5108,N_2175,N_195);
nor U5109 (N_5109,N_97,N_2325);
nand U5110 (N_5110,N_811,N_2920);
nand U5111 (N_5111,N_1176,N_2368);
and U5112 (N_5112,N_2560,N_103);
nand U5113 (N_5113,N_935,N_2335);
nand U5114 (N_5114,N_2846,N_2348);
or U5115 (N_5115,N_216,N_2144);
nand U5116 (N_5116,N_491,N_185);
or U5117 (N_5117,N_397,N_771);
and U5118 (N_5118,N_1740,N_1150);
nand U5119 (N_5119,N_2713,N_1200);
nand U5120 (N_5120,N_1535,N_2947);
or U5121 (N_5121,N_599,N_1791);
and U5122 (N_5122,N_2689,N_2528);
nand U5123 (N_5123,N_2750,N_1199);
nor U5124 (N_5124,N_795,N_2067);
and U5125 (N_5125,N_2148,N_1672);
nand U5126 (N_5126,N_2197,N_1071);
and U5127 (N_5127,N_767,N_2514);
or U5128 (N_5128,N_2020,N_2550);
nand U5129 (N_5129,N_128,N_1394);
and U5130 (N_5130,N_1280,N_173);
and U5131 (N_5131,N_1402,N_509);
or U5132 (N_5132,N_1001,N_951);
xor U5133 (N_5133,N_2367,N_1070);
nor U5134 (N_5134,N_1992,N_2809);
and U5135 (N_5135,N_1030,N_1541);
or U5136 (N_5136,N_386,N_2168);
nor U5137 (N_5137,N_2900,N_1492);
or U5138 (N_5138,N_2035,N_2955);
or U5139 (N_5139,N_713,N_362);
nand U5140 (N_5140,N_50,N_2617);
nand U5141 (N_5141,N_2677,N_1090);
xor U5142 (N_5142,N_1495,N_254);
nand U5143 (N_5143,N_1839,N_1541);
nand U5144 (N_5144,N_571,N_677);
nor U5145 (N_5145,N_188,N_2529);
xnor U5146 (N_5146,N_1493,N_2036);
nand U5147 (N_5147,N_2251,N_2992);
xor U5148 (N_5148,N_280,N_1198);
nor U5149 (N_5149,N_2438,N_46);
or U5150 (N_5150,N_355,N_212);
nor U5151 (N_5151,N_180,N_1729);
nand U5152 (N_5152,N_1989,N_99);
xnor U5153 (N_5153,N_574,N_1569);
and U5154 (N_5154,N_998,N_393);
or U5155 (N_5155,N_2958,N_1820);
nor U5156 (N_5156,N_2074,N_486);
nor U5157 (N_5157,N_106,N_2878);
or U5158 (N_5158,N_2359,N_574);
nor U5159 (N_5159,N_2593,N_2696);
and U5160 (N_5160,N_2221,N_182);
nand U5161 (N_5161,N_1544,N_2147);
nand U5162 (N_5162,N_797,N_2107);
nand U5163 (N_5163,N_1534,N_2991);
and U5164 (N_5164,N_2929,N_752);
nand U5165 (N_5165,N_436,N_1071);
or U5166 (N_5166,N_345,N_2884);
or U5167 (N_5167,N_1798,N_1746);
nor U5168 (N_5168,N_2590,N_2215);
and U5169 (N_5169,N_2429,N_1398);
nor U5170 (N_5170,N_2422,N_1378);
nor U5171 (N_5171,N_87,N_1069);
nand U5172 (N_5172,N_2481,N_2490);
xor U5173 (N_5173,N_2366,N_124);
nor U5174 (N_5174,N_1469,N_84);
nor U5175 (N_5175,N_369,N_55);
or U5176 (N_5176,N_2445,N_2364);
or U5177 (N_5177,N_344,N_2145);
and U5178 (N_5178,N_2215,N_212);
nand U5179 (N_5179,N_1737,N_2299);
or U5180 (N_5180,N_1195,N_2295);
nand U5181 (N_5181,N_2277,N_969);
or U5182 (N_5182,N_2972,N_1813);
or U5183 (N_5183,N_1874,N_1284);
nand U5184 (N_5184,N_665,N_286);
or U5185 (N_5185,N_2082,N_1690);
xnor U5186 (N_5186,N_561,N_2003);
nand U5187 (N_5187,N_44,N_296);
or U5188 (N_5188,N_690,N_619);
nor U5189 (N_5189,N_2160,N_2986);
and U5190 (N_5190,N_1024,N_422);
nor U5191 (N_5191,N_181,N_449);
nor U5192 (N_5192,N_295,N_2529);
nand U5193 (N_5193,N_2772,N_241);
or U5194 (N_5194,N_240,N_2684);
nor U5195 (N_5195,N_1175,N_2500);
nand U5196 (N_5196,N_2344,N_2423);
or U5197 (N_5197,N_2599,N_459);
nor U5198 (N_5198,N_215,N_2837);
or U5199 (N_5199,N_2237,N_502);
and U5200 (N_5200,N_2861,N_764);
or U5201 (N_5201,N_1097,N_475);
nor U5202 (N_5202,N_1334,N_97);
nor U5203 (N_5203,N_2346,N_437);
and U5204 (N_5204,N_1195,N_2740);
and U5205 (N_5205,N_1203,N_789);
or U5206 (N_5206,N_437,N_1474);
or U5207 (N_5207,N_555,N_1328);
nand U5208 (N_5208,N_2666,N_2814);
nor U5209 (N_5209,N_415,N_1307);
nor U5210 (N_5210,N_1963,N_641);
nor U5211 (N_5211,N_1769,N_564);
nand U5212 (N_5212,N_2953,N_2453);
or U5213 (N_5213,N_2662,N_237);
nor U5214 (N_5214,N_1501,N_270);
or U5215 (N_5215,N_1655,N_2334);
and U5216 (N_5216,N_1592,N_1945);
nor U5217 (N_5217,N_1474,N_1934);
or U5218 (N_5218,N_1260,N_2087);
or U5219 (N_5219,N_1331,N_375);
nor U5220 (N_5220,N_1225,N_2462);
and U5221 (N_5221,N_644,N_278);
and U5222 (N_5222,N_1109,N_46);
nor U5223 (N_5223,N_1090,N_2618);
nor U5224 (N_5224,N_2121,N_2612);
nand U5225 (N_5225,N_2433,N_832);
or U5226 (N_5226,N_996,N_2405);
nand U5227 (N_5227,N_716,N_687);
nor U5228 (N_5228,N_2375,N_1082);
nor U5229 (N_5229,N_1784,N_121);
nand U5230 (N_5230,N_592,N_638);
nand U5231 (N_5231,N_57,N_1170);
or U5232 (N_5232,N_43,N_2892);
or U5233 (N_5233,N_2727,N_2902);
and U5234 (N_5234,N_2053,N_91);
nand U5235 (N_5235,N_875,N_1061);
nor U5236 (N_5236,N_70,N_293);
nor U5237 (N_5237,N_747,N_1460);
and U5238 (N_5238,N_419,N_2435);
or U5239 (N_5239,N_137,N_2960);
and U5240 (N_5240,N_2256,N_305);
and U5241 (N_5241,N_1878,N_2413);
nor U5242 (N_5242,N_1456,N_341);
and U5243 (N_5243,N_1628,N_293);
and U5244 (N_5244,N_2028,N_1153);
and U5245 (N_5245,N_473,N_295);
or U5246 (N_5246,N_2547,N_186);
xor U5247 (N_5247,N_2349,N_1002);
nor U5248 (N_5248,N_2922,N_1938);
nor U5249 (N_5249,N_1173,N_1775);
and U5250 (N_5250,N_2327,N_2248);
or U5251 (N_5251,N_1537,N_1142);
nor U5252 (N_5252,N_923,N_918);
and U5253 (N_5253,N_554,N_2753);
nand U5254 (N_5254,N_331,N_52);
and U5255 (N_5255,N_393,N_2599);
nor U5256 (N_5256,N_685,N_1077);
or U5257 (N_5257,N_2591,N_607);
or U5258 (N_5258,N_4,N_25);
nor U5259 (N_5259,N_1882,N_745);
and U5260 (N_5260,N_2988,N_49);
or U5261 (N_5261,N_19,N_258);
and U5262 (N_5262,N_920,N_2371);
nand U5263 (N_5263,N_903,N_229);
nor U5264 (N_5264,N_961,N_51);
nand U5265 (N_5265,N_960,N_1578);
or U5266 (N_5266,N_618,N_1981);
or U5267 (N_5267,N_2572,N_1370);
nand U5268 (N_5268,N_2758,N_2822);
or U5269 (N_5269,N_2828,N_2515);
and U5270 (N_5270,N_142,N_69);
or U5271 (N_5271,N_2945,N_246);
nor U5272 (N_5272,N_837,N_16);
nor U5273 (N_5273,N_1424,N_543);
or U5274 (N_5274,N_2520,N_1644);
xor U5275 (N_5275,N_2996,N_605);
nor U5276 (N_5276,N_1368,N_2303);
nand U5277 (N_5277,N_1290,N_1346);
nor U5278 (N_5278,N_906,N_504);
and U5279 (N_5279,N_924,N_1665);
nand U5280 (N_5280,N_1044,N_2738);
or U5281 (N_5281,N_2875,N_2173);
nor U5282 (N_5282,N_2540,N_1559);
and U5283 (N_5283,N_2924,N_2523);
and U5284 (N_5284,N_2661,N_556);
or U5285 (N_5285,N_120,N_1658);
nor U5286 (N_5286,N_464,N_1240);
or U5287 (N_5287,N_1698,N_936);
and U5288 (N_5288,N_1239,N_2614);
or U5289 (N_5289,N_1972,N_2754);
nor U5290 (N_5290,N_2191,N_1809);
or U5291 (N_5291,N_119,N_853);
and U5292 (N_5292,N_1698,N_492);
nand U5293 (N_5293,N_2708,N_2989);
or U5294 (N_5294,N_2853,N_788);
nor U5295 (N_5295,N_799,N_2180);
and U5296 (N_5296,N_2152,N_893);
or U5297 (N_5297,N_275,N_2269);
and U5298 (N_5298,N_187,N_293);
and U5299 (N_5299,N_1689,N_1467);
nand U5300 (N_5300,N_155,N_531);
nor U5301 (N_5301,N_2736,N_123);
nor U5302 (N_5302,N_2984,N_1170);
nand U5303 (N_5303,N_2290,N_1849);
nand U5304 (N_5304,N_2302,N_1216);
or U5305 (N_5305,N_1715,N_2515);
or U5306 (N_5306,N_1716,N_474);
nor U5307 (N_5307,N_2766,N_2918);
nor U5308 (N_5308,N_1922,N_2966);
or U5309 (N_5309,N_279,N_2366);
or U5310 (N_5310,N_1829,N_2103);
nand U5311 (N_5311,N_1299,N_394);
nor U5312 (N_5312,N_2926,N_380);
and U5313 (N_5313,N_2945,N_1240);
nand U5314 (N_5314,N_1402,N_1753);
nand U5315 (N_5315,N_2548,N_411);
nor U5316 (N_5316,N_1112,N_2580);
nand U5317 (N_5317,N_1410,N_104);
and U5318 (N_5318,N_721,N_1174);
nor U5319 (N_5319,N_299,N_377);
and U5320 (N_5320,N_2094,N_2821);
nand U5321 (N_5321,N_1654,N_539);
nand U5322 (N_5322,N_2999,N_602);
and U5323 (N_5323,N_2147,N_500);
nand U5324 (N_5324,N_2201,N_1128);
xor U5325 (N_5325,N_2036,N_2708);
and U5326 (N_5326,N_846,N_2757);
or U5327 (N_5327,N_525,N_181);
nand U5328 (N_5328,N_801,N_766);
or U5329 (N_5329,N_1499,N_694);
and U5330 (N_5330,N_594,N_415);
or U5331 (N_5331,N_1406,N_889);
nand U5332 (N_5332,N_1556,N_2134);
nand U5333 (N_5333,N_702,N_932);
and U5334 (N_5334,N_666,N_1517);
or U5335 (N_5335,N_516,N_2891);
and U5336 (N_5336,N_202,N_371);
or U5337 (N_5337,N_2634,N_1614);
nand U5338 (N_5338,N_1539,N_1495);
and U5339 (N_5339,N_873,N_696);
nand U5340 (N_5340,N_2624,N_2031);
and U5341 (N_5341,N_2001,N_1586);
and U5342 (N_5342,N_823,N_711);
nor U5343 (N_5343,N_1865,N_1151);
nor U5344 (N_5344,N_2437,N_2219);
and U5345 (N_5345,N_1426,N_2480);
and U5346 (N_5346,N_2411,N_1970);
and U5347 (N_5347,N_1718,N_2997);
nand U5348 (N_5348,N_1027,N_1388);
or U5349 (N_5349,N_2412,N_1720);
nand U5350 (N_5350,N_1355,N_416);
or U5351 (N_5351,N_1420,N_27);
or U5352 (N_5352,N_1703,N_2598);
nor U5353 (N_5353,N_2412,N_2084);
or U5354 (N_5354,N_1920,N_1766);
nor U5355 (N_5355,N_1067,N_2739);
nor U5356 (N_5356,N_1410,N_2834);
xnor U5357 (N_5357,N_851,N_2638);
or U5358 (N_5358,N_14,N_323);
nand U5359 (N_5359,N_2856,N_2483);
nand U5360 (N_5360,N_1987,N_2998);
and U5361 (N_5361,N_1821,N_2526);
nor U5362 (N_5362,N_1547,N_2379);
nor U5363 (N_5363,N_1785,N_2855);
nand U5364 (N_5364,N_1387,N_2305);
and U5365 (N_5365,N_1745,N_2907);
nor U5366 (N_5366,N_800,N_1567);
or U5367 (N_5367,N_1447,N_2243);
and U5368 (N_5368,N_990,N_204);
nand U5369 (N_5369,N_2537,N_401);
or U5370 (N_5370,N_37,N_206);
or U5371 (N_5371,N_61,N_239);
or U5372 (N_5372,N_1583,N_1212);
or U5373 (N_5373,N_2506,N_2726);
nor U5374 (N_5374,N_1453,N_32);
nand U5375 (N_5375,N_1300,N_477);
nor U5376 (N_5376,N_2795,N_2218);
or U5377 (N_5377,N_2294,N_2473);
or U5378 (N_5378,N_882,N_2398);
nor U5379 (N_5379,N_1543,N_1644);
xnor U5380 (N_5380,N_1577,N_852);
or U5381 (N_5381,N_640,N_2076);
or U5382 (N_5382,N_1677,N_2619);
nand U5383 (N_5383,N_1161,N_328);
or U5384 (N_5384,N_1190,N_2866);
and U5385 (N_5385,N_2126,N_2464);
or U5386 (N_5386,N_209,N_2097);
and U5387 (N_5387,N_1976,N_2928);
xor U5388 (N_5388,N_2239,N_1361);
or U5389 (N_5389,N_1064,N_526);
or U5390 (N_5390,N_719,N_103);
nand U5391 (N_5391,N_2450,N_187);
and U5392 (N_5392,N_1353,N_592);
nand U5393 (N_5393,N_252,N_1516);
or U5394 (N_5394,N_2072,N_1610);
xor U5395 (N_5395,N_925,N_1193);
or U5396 (N_5396,N_1629,N_787);
nand U5397 (N_5397,N_891,N_1192);
and U5398 (N_5398,N_1592,N_1191);
nor U5399 (N_5399,N_553,N_47);
nor U5400 (N_5400,N_622,N_2400);
nor U5401 (N_5401,N_2659,N_2574);
and U5402 (N_5402,N_2491,N_2099);
nand U5403 (N_5403,N_2687,N_1083);
and U5404 (N_5404,N_703,N_1261);
nor U5405 (N_5405,N_1884,N_1400);
and U5406 (N_5406,N_2302,N_305);
or U5407 (N_5407,N_996,N_302);
and U5408 (N_5408,N_472,N_646);
or U5409 (N_5409,N_259,N_543);
nor U5410 (N_5410,N_1716,N_2771);
or U5411 (N_5411,N_664,N_1562);
or U5412 (N_5412,N_712,N_1963);
and U5413 (N_5413,N_223,N_31);
or U5414 (N_5414,N_1019,N_1104);
and U5415 (N_5415,N_325,N_2621);
or U5416 (N_5416,N_2149,N_33);
or U5417 (N_5417,N_2833,N_552);
nor U5418 (N_5418,N_1552,N_1325);
nor U5419 (N_5419,N_1361,N_1182);
nor U5420 (N_5420,N_1245,N_1981);
nand U5421 (N_5421,N_242,N_1489);
nand U5422 (N_5422,N_2767,N_2180);
nor U5423 (N_5423,N_2696,N_2887);
nand U5424 (N_5424,N_621,N_166);
and U5425 (N_5425,N_2965,N_96);
or U5426 (N_5426,N_847,N_673);
and U5427 (N_5427,N_1380,N_1558);
nand U5428 (N_5428,N_2165,N_2693);
or U5429 (N_5429,N_2559,N_2355);
or U5430 (N_5430,N_1472,N_1008);
and U5431 (N_5431,N_2549,N_2903);
or U5432 (N_5432,N_2748,N_257);
nor U5433 (N_5433,N_1384,N_65);
nand U5434 (N_5434,N_2313,N_2476);
nor U5435 (N_5435,N_2983,N_446);
or U5436 (N_5436,N_2081,N_2447);
and U5437 (N_5437,N_1764,N_1237);
and U5438 (N_5438,N_1407,N_1628);
and U5439 (N_5439,N_2347,N_543);
xor U5440 (N_5440,N_2824,N_1640);
and U5441 (N_5441,N_490,N_2430);
nand U5442 (N_5442,N_2443,N_1483);
nand U5443 (N_5443,N_2440,N_349);
or U5444 (N_5444,N_2991,N_2401);
nor U5445 (N_5445,N_900,N_2557);
and U5446 (N_5446,N_164,N_1874);
and U5447 (N_5447,N_2047,N_1887);
nor U5448 (N_5448,N_1711,N_2735);
or U5449 (N_5449,N_437,N_2094);
nor U5450 (N_5450,N_825,N_850);
nand U5451 (N_5451,N_596,N_1930);
nor U5452 (N_5452,N_666,N_2147);
or U5453 (N_5453,N_2658,N_1478);
nand U5454 (N_5454,N_2652,N_1202);
or U5455 (N_5455,N_1220,N_2563);
and U5456 (N_5456,N_2221,N_1997);
nor U5457 (N_5457,N_221,N_2314);
and U5458 (N_5458,N_439,N_1850);
nand U5459 (N_5459,N_871,N_2457);
or U5460 (N_5460,N_2797,N_856);
and U5461 (N_5461,N_162,N_1522);
nor U5462 (N_5462,N_2391,N_421);
nor U5463 (N_5463,N_1011,N_1651);
nor U5464 (N_5464,N_129,N_1962);
and U5465 (N_5465,N_2023,N_2576);
nand U5466 (N_5466,N_1623,N_2415);
or U5467 (N_5467,N_2516,N_1422);
nor U5468 (N_5468,N_2333,N_1821);
or U5469 (N_5469,N_640,N_60);
nand U5470 (N_5470,N_1050,N_358);
nand U5471 (N_5471,N_2773,N_2181);
nor U5472 (N_5472,N_107,N_2777);
xnor U5473 (N_5473,N_533,N_678);
nor U5474 (N_5474,N_1383,N_2587);
or U5475 (N_5475,N_805,N_1642);
nor U5476 (N_5476,N_979,N_1404);
and U5477 (N_5477,N_1387,N_2858);
or U5478 (N_5478,N_2168,N_1432);
and U5479 (N_5479,N_2800,N_798);
and U5480 (N_5480,N_674,N_2216);
nor U5481 (N_5481,N_927,N_2402);
nor U5482 (N_5482,N_2253,N_265);
nor U5483 (N_5483,N_791,N_2434);
or U5484 (N_5484,N_1178,N_627);
and U5485 (N_5485,N_1328,N_31);
and U5486 (N_5486,N_1517,N_1004);
xnor U5487 (N_5487,N_29,N_2728);
and U5488 (N_5488,N_145,N_2451);
nand U5489 (N_5489,N_724,N_169);
nand U5490 (N_5490,N_1460,N_2400);
nor U5491 (N_5491,N_1730,N_131);
nand U5492 (N_5492,N_752,N_2242);
and U5493 (N_5493,N_1940,N_2513);
nand U5494 (N_5494,N_334,N_2505);
xnor U5495 (N_5495,N_681,N_2935);
or U5496 (N_5496,N_530,N_2589);
and U5497 (N_5497,N_46,N_215);
and U5498 (N_5498,N_158,N_383);
nor U5499 (N_5499,N_1982,N_1382);
nand U5500 (N_5500,N_2640,N_1452);
nand U5501 (N_5501,N_2710,N_1780);
and U5502 (N_5502,N_595,N_2135);
or U5503 (N_5503,N_2533,N_104);
nor U5504 (N_5504,N_45,N_1784);
nand U5505 (N_5505,N_1115,N_2179);
nor U5506 (N_5506,N_2378,N_882);
nand U5507 (N_5507,N_1641,N_1411);
or U5508 (N_5508,N_2499,N_1667);
nand U5509 (N_5509,N_271,N_2829);
nand U5510 (N_5510,N_276,N_248);
nor U5511 (N_5511,N_1446,N_1707);
or U5512 (N_5512,N_524,N_350);
and U5513 (N_5513,N_249,N_2154);
and U5514 (N_5514,N_1768,N_2727);
and U5515 (N_5515,N_1552,N_420);
and U5516 (N_5516,N_498,N_1639);
nand U5517 (N_5517,N_111,N_2117);
and U5518 (N_5518,N_1295,N_104);
nor U5519 (N_5519,N_2972,N_144);
xor U5520 (N_5520,N_2175,N_2337);
or U5521 (N_5521,N_1265,N_496);
nand U5522 (N_5522,N_2424,N_1101);
nor U5523 (N_5523,N_800,N_1853);
nor U5524 (N_5524,N_955,N_399);
or U5525 (N_5525,N_59,N_2571);
nand U5526 (N_5526,N_1157,N_2350);
nand U5527 (N_5527,N_1168,N_1310);
xor U5528 (N_5528,N_1743,N_2966);
nand U5529 (N_5529,N_1747,N_2740);
nor U5530 (N_5530,N_703,N_656);
and U5531 (N_5531,N_2577,N_1814);
or U5532 (N_5532,N_2560,N_1140);
nor U5533 (N_5533,N_819,N_94);
nor U5534 (N_5534,N_280,N_1608);
or U5535 (N_5535,N_2275,N_789);
nand U5536 (N_5536,N_24,N_1574);
and U5537 (N_5537,N_1108,N_258);
or U5538 (N_5538,N_2730,N_2165);
nand U5539 (N_5539,N_1471,N_1432);
nand U5540 (N_5540,N_798,N_235);
nor U5541 (N_5541,N_2517,N_2574);
or U5542 (N_5542,N_1311,N_818);
or U5543 (N_5543,N_443,N_2322);
nand U5544 (N_5544,N_1349,N_118);
and U5545 (N_5545,N_1886,N_170);
and U5546 (N_5546,N_1697,N_1418);
nand U5547 (N_5547,N_2284,N_2465);
and U5548 (N_5548,N_636,N_127);
nor U5549 (N_5549,N_103,N_221);
or U5550 (N_5550,N_2608,N_1947);
nor U5551 (N_5551,N_2615,N_1501);
nor U5552 (N_5552,N_452,N_2073);
nand U5553 (N_5553,N_2261,N_1021);
and U5554 (N_5554,N_1544,N_2878);
or U5555 (N_5555,N_2375,N_194);
and U5556 (N_5556,N_1694,N_789);
nand U5557 (N_5557,N_2824,N_1833);
or U5558 (N_5558,N_116,N_1761);
or U5559 (N_5559,N_1430,N_193);
nand U5560 (N_5560,N_2153,N_2213);
nand U5561 (N_5561,N_1934,N_2537);
and U5562 (N_5562,N_2342,N_1779);
or U5563 (N_5563,N_2704,N_1120);
nor U5564 (N_5564,N_865,N_1874);
nand U5565 (N_5565,N_201,N_2683);
or U5566 (N_5566,N_1350,N_1079);
nand U5567 (N_5567,N_1079,N_1038);
nand U5568 (N_5568,N_1983,N_2376);
and U5569 (N_5569,N_1337,N_2706);
nand U5570 (N_5570,N_481,N_2079);
nand U5571 (N_5571,N_480,N_624);
nor U5572 (N_5572,N_1009,N_2579);
nand U5573 (N_5573,N_242,N_813);
and U5574 (N_5574,N_2697,N_460);
or U5575 (N_5575,N_667,N_828);
nand U5576 (N_5576,N_2284,N_475);
and U5577 (N_5577,N_1684,N_1739);
nor U5578 (N_5578,N_2285,N_2693);
and U5579 (N_5579,N_1015,N_744);
and U5580 (N_5580,N_2564,N_1766);
nand U5581 (N_5581,N_822,N_1690);
nor U5582 (N_5582,N_1191,N_80);
and U5583 (N_5583,N_896,N_708);
nand U5584 (N_5584,N_1174,N_2695);
nor U5585 (N_5585,N_796,N_1381);
or U5586 (N_5586,N_352,N_596);
nand U5587 (N_5587,N_1168,N_2080);
and U5588 (N_5588,N_1367,N_1511);
or U5589 (N_5589,N_1322,N_2033);
nand U5590 (N_5590,N_2453,N_1522);
or U5591 (N_5591,N_1910,N_1479);
nand U5592 (N_5592,N_475,N_1338);
nor U5593 (N_5593,N_2059,N_1594);
or U5594 (N_5594,N_171,N_1876);
and U5595 (N_5595,N_1198,N_2606);
and U5596 (N_5596,N_1439,N_2051);
and U5597 (N_5597,N_1664,N_1970);
nor U5598 (N_5598,N_1004,N_584);
nor U5599 (N_5599,N_2781,N_2515);
nor U5600 (N_5600,N_68,N_735);
or U5601 (N_5601,N_1043,N_192);
nand U5602 (N_5602,N_2559,N_1271);
xor U5603 (N_5603,N_313,N_1152);
or U5604 (N_5604,N_1076,N_1319);
or U5605 (N_5605,N_674,N_1273);
nand U5606 (N_5606,N_1628,N_273);
nor U5607 (N_5607,N_2657,N_2623);
nor U5608 (N_5608,N_2911,N_1670);
and U5609 (N_5609,N_295,N_2658);
nand U5610 (N_5610,N_2585,N_660);
and U5611 (N_5611,N_2356,N_2405);
or U5612 (N_5612,N_1697,N_1268);
or U5613 (N_5613,N_2847,N_2741);
and U5614 (N_5614,N_154,N_780);
and U5615 (N_5615,N_1441,N_2851);
nor U5616 (N_5616,N_2155,N_2114);
nand U5617 (N_5617,N_299,N_953);
nand U5618 (N_5618,N_716,N_1532);
nor U5619 (N_5619,N_2581,N_2965);
and U5620 (N_5620,N_975,N_910);
nor U5621 (N_5621,N_2751,N_2095);
nand U5622 (N_5622,N_2699,N_396);
xor U5623 (N_5623,N_1539,N_422);
nand U5624 (N_5624,N_220,N_1508);
nor U5625 (N_5625,N_444,N_301);
and U5626 (N_5626,N_2143,N_2265);
nor U5627 (N_5627,N_2122,N_76);
and U5628 (N_5628,N_1300,N_197);
and U5629 (N_5629,N_1758,N_2125);
or U5630 (N_5630,N_2176,N_1911);
nand U5631 (N_5631,N_2942,N_1727);
or U5632 (N_5632,N_2146,N_1230);
and U5633 (N_5633,N_372,N_2240);
nand U5634 (N_5634,N_2574,N_1757);
nand U5635 (N_5635,N_2570,N_2795);
and U5636 (N_5636,N_594,N_435);
or U5637 (N_5637,N_2348,N_2418);
nor U5638 (N_5638,N_1408,N_1798);
nor U5639 (N_5639,N_1877,N_2304);
and U5640 (N_5640,N_1847,N_589);
and U5641 (N_5641,N_1612,N_1480);
or U5642 (N_5642,N_1998,N_1279);
nand U5643 (N_5643,N_913,N_1470);
or U5644 (N_5644,N_1092,N_125);
nand U5645 (N_5645,N_1504,N_1084);
nand U5646 (N_5646,N_2221,N_2799);
xor U5647 (N_5647,N_1732,N_1662);
nor U5648 (N_5648,N_535,N_2293);
or U5649 (N_5649,N_420,N_160);
or U5650 (N_5650,N_1636,N_2511);
and U5651 (N_5651,N_340,N_490);
and U5652 (N_5652,N_2497,N_774);
nand U5653 (N_5653,N_1382,N_2313);
nor U5654 (N_5654,N_499,N_2041);
nor U5655 (N_5655,N_2670,N_2958);
or U5656 (N_5656,N_1904,N_2705);
xor U5657 (N_5657,N_170,N_1258);
or U5658 (N_5658,N_829,N_1646);
or U5659 (N_5659,N_253,N_533);
and U5660 (N_5660,N_867,N_2686);
nor U5661 (N_5661,N_2787,N_598);
nor U5662 (N_5662,N_1006,N_2792);
or U5663 (N_5663,N_1821,N_499);
or U5664 (N_5664,N_2257,N_915);
or U5665 (N_5665,N_2971,N_2246);
or U5666 (N_5666,N_2309,N_476);
nor U5667 (N_5667,N_1827,N_1145);
or U5668 (N_5668,N_1567,N_2830);
xor U5669 (N_5669,N_370,N_837);
nand U5670 (N_5670,N_2789,N_699);
nand U5671 (N_5671,N_2609,N_2848);
nor U5672 (N_5672,N_1844,N_779);
and U5673 (N_5673,N_1252,N_251);
or U5674 (N_5674,N_2331,N_881);
nand U5675 (N_5675,N_2426,N_504);
or U5676 (N_5676,N_1477,N_850);
and U5677 (N_5677,N_2977,N_1430);
or U5678 (N_5678,N_748,N_2316);
or U5679 (N_5679,N_1818,N_1310);
nor U5680 (N_5680,N_1851,N_1562);
or U5681 (N_5681,N_1881,N_1565);
nor U5682 (N_5682,N_2553,N_361);
and U5683 (N_5683,N_229,N_1649);
or U5684 (N_5684,N_2868,N_1786);
nand U5685 (N_5685,N_1460,N_1164);
or U5686 (N_5686,N_399,N_259);
and U5687 (N_5687,N_1382,N_81);
or U5688 (N_5688,N_2583,N_326);
xnor U5689 (N_5689,N_2825,N_710);
or U5690 (N_5690,N_1830,N_149);
and U5691 (N_5691,N_349,N_2814);
and U5692 (N_5692,N_1075,N_1449);
and U5693 (N_5693,N_2712,N_1171);
and U5694 (N_5694,N_105,N_819);
nor U5695 (N_5695,N_688,N_433);
nand U5696 (N_5696,N_571,N_1593);
and U5697 (N_5697,N_1938,N_2587);
nand U5698 (N_5698,N_1880,N_730);
nand U5699 (N_5699,N_1952,N_520);
and U5700 (N_5700,N_1552,N_1000);
and U5701 (N_5701,N_995,N_2034);
and U5702 (N_5702,N_633,N_1079);
nand U5703 (N_5703,N_1,N_1500);
nor U5704 (N_5704,N_2924,N_1392);
nor U5705 (N_5705,N_2727,N_1243);
nor U5706 (N_5706,N_2840,N_1424);
nor U5707 (N_5707,N_1758,N_1701);
or U5708 (N_5708,N_1147,N_520);
and U5709 (N_5709,N_1089,N_1241);
nand U5710 (N_5710,N_2647,N_2127);
and U5711 (N_5711,N_1516,N_250);
and U5712 (N_5712,N_1026,N_1139);
and U5713 (N_5713,N_708,N_1664);
nand U5714 (N_5714,N_2633,N_1408);
nor U5715 (N_5715,N_1045,N_1765);
or U5716 (N_5716,N_2554,N_2697);
or U5717 (N_5717,N_1739,N_2220);
nand U5718 (N_5718,N_203,N_2123);
nor U5719 (N_5719,N_2607,N_772);
xor U5720 (N_5720,N_297,N_2618);
nand U5721 (N_5721,N_1033,N_2320);
xnor U5722 (N_5722,N_2270,N_1855);
nor U5723 (N_5723,N_352,N_655);
or U5724 (N_5724,N_1425,N_2952);
or U5725 (N_5725,N_300,N_2948);
and U5726 (N_5726,N_142,N_2688);
or U5727 (N_5727,N_1218,N_1657);
nand U5728 (N_5728,N_2329,N_1591);
nor U5729 (N_5729,N_2117,N_2434);
nor U5730 (N_5730,N_1503,N_1486);
and U5731 (N_5731,N_1850,N_735);
nand U5732 (N_5732,N_2054,N_2838);
and U5733 (N_5733,N_1053,N_2234);
or U5734 (N_5734,N_1146,N_1495);
and U5735 (N_5735,N_2689,N_2517);
and U5736 (N_5736,N_1166,N_54);
nand U5737 (N_5737,N_2531,N_2367);
nand U5738 (N_5738,N_382,N_2712);
nand U5739 (N_5739,N_938,N_166);
nor U5740 (N_5740,N_294,N_1246);
nor U5741 (N_5741,N_261,N_756);
nand U5742 (N_5742,N_706,N_312);
or U5743 (N_5743,N_2098,N_1991);
nor U5744 (N_5744,N_384,N_324);
and U5745 (N_5745,N_2902,N_193);
or U5746 (N_5746,N_2773,N_708);
and U5747 (N_5747,N_2870,N_2037);
nor U5748 (N_5748,N_2490,N_1449);
nand U5749 (N_5749,N_1387,N_1781);
or U5750 (N_5750,N_1214,N_987);
or U5751 (N_5751,N_746,N_1487);
or U5752 (N_5752,N_1083,N_2309);
nor U5753 (N_5753,N_15,N_1798);
nor U5754 (N_5754,N_2631,N_1950);
or U5755 (N_5755,N_1345,N_191);
and U5756 (N_5756,N_913,N_486);
nor U5757 (N_5757,N_2195,N_468);
or U5758 (N_5758,N_2411,N_2985);
xor U5759 (N_5759,N_1132,N_1660);
and U5760 (N_5760,N_2309,N_1114);
or U5761 (N_5761,N_2804,N_811);
or U5762 (N_5762,N_1975,N_18);
and U5763 (N_5763,N_1258,N_449);
or U5764 (N_5764,N_30,N_1349);
nor U5765 (N_5765,N_2628,N_1547);
nand U5766 (N_5766,N_1451,N_1482);
nand U5767 (N_5767,N_836,N_901);
and U5768 (N_5768,N_462,N_1504);
or U5769 (N_5769,N_1041,N_1181);
or U5770 (N_5770,N_1235,N_2427);
or U5771 (N_5771,N_787,N_2197);
and U5772 (N_5772,N_452,N_877);
nor U5773 (N_5773,N_1646,N_2182);
nand U5774 (N_5774,N_1570,N_1150);
nor U5775 (N_5775,N_885,N_1573);
nor U5776 (N_5776,N_1061,N_718);
nor U5777 (N_5777,N_1,N_392);
and U5778 (N_5778,N_954,N_616);
and U5779 (N_5779,N_734,N_2929);
nor U5780 (N_5780,N_484,N_235);
or U5781 (N_5781,N_1275,N_2152);
nor U5782 (N_5782,N_1637,N_2443);
nor U5783 (N_5783,N_241,N_1063);
nor U5784 (N_5784,N_2339,N_2769);
nor U5785 (N_5785,N_1856,N_2417);
or U5786 (N_5786,N_183,N_2744);
nor U5787 (N_5787,N_2600,N_1163);
and U5788 (N_5788,N_1200,N_1905);
xnor U5789 (N_5789,N_1537,N_1748);
nor U5790 (N_5790,N_2560,N_1847);
nor U5791 (N_5791,N_1045,N_1663);
nand U5792 (N_5792,N_1556,N_1860);
nand U5793 (N_5793,N_1335,N_374);
or U5794 (N_5794,N_1452,N_2381);
or U5795 (N_5795,N_2552,N_2840);
or U5796 (N_5796,N_830,N_158);
xor U5797 (N_5797,N_2790,N_1299);
nor U5798 (N_5798,N_2771,N_2069);
or U5799 (N_5799,N_2594,N_2460);
and U5800 (N_5800,N_1908,N_2863);
or U5801 (N_5801,N_1219,N_2552);
or U5802 (N_5802,N_1543,N_2186);
nand U5803 (N_5803,N_1808,N_1865);
nor U5804 (N_5804,N_929,N_2837);
nor U5805 (N_5805,N_2510,N_1054);
nand U5806 (N_5806,N_1050,N_1509);
nor U5807 (N_5807,N_1764,N_2323);
nor U5808 (N_5808,N_934,N_395);
and U5809 (N_5809,N_942,N_2293);
or U5810 (N_5810,N_1106,N_1314);
and U5811 (N_5811,N_1995,N_1464);
or U5812 (N_5812,N_1772,N_437);
or U5813 (N_5813,N_1236,N_2620);
and U5814 (N_5814,N_1414,N_1694);
nand U5815 (N_5815,N_627,N_111);
and U5816 (N_5816,N_772,N_1708);
or U5817 (N_5817,N_1323,N_762);
nand U5818 (N_5818,N_2239,N_1211);
nand U5819 (N_5819,N_60,N_1530);
nand U5820 (N_5820,N_2719,N_2215);
nor U5821 (N_5821,N_1757,N_1289);
or U5822 (N_5822,N_1623,N_1178);
and U5823 (N_5823,N_1862,N_1673);
or U5824 (N_5824,N_1792,N_2054);
nor U5825 (N_5825,N_1479,N_1659);
nor U5826 (N_5826,N_1953,N_2337);
nand U5827 (N_5827,N_1472,N_2503);
nor U5828 (N_5828,N_215,N_22);
and U5829 (N_5829,N_1697,N_992);
and U5830 (N_5830,N_2445,N_1655);
nand U5831 (N_5831,N_2292,N_1894);
and U5832 (N_5832,N_2250,N_2220);
or U5833 (N_5833,N_2191,N_1621);
or U5834 (N_5834,N_1842,N_1209);
and U5835 (N_5835,N_2952,N_2773);
nor U5836 (N_5836,N_2720,N_2710);
and U5837 (N_5837,N_1667,N_1363);
and U5838 (N_5838,N_495,N_859);
or U5839 (N_5839,N_827,N_1237);
and U5840 (N_5840,N_1954,N_1904);
and U5841 (N_5841,N_596,N_1562);
and U5842 (N_5842,N_1097,N_340);
and U5843 (N_5843,N_677,N_1514);
nor U5844 (N_5844,N_687,N_2205);
xor U5845 (N_5845,N_2613,N_2235);
nor U5846 (N_5846,N_2948,N_843);
and U5847 (N_5847,N_493,N_2543);
or U5848 (N_5848,N_2952,N_2379);
or U5849 (N_5849,N_1651,N_1682);
nor U5850 (N_5850,N_2194,N_2495);
or U5851 (N_5851,N_540,N_1746);
nand U5852 (N_5852,N_2756,N_732);
and U5853 (N_5853,N_537,N_1473);
nand U5854 (N_5854,N_2901,N_1033);
or U5855 (N_5855,N_2546,N_1155);
nor U5856 (N_5856,N_1801,N_2412);
nand U5857 (N_5857,N_636,N_1512);
nor U5858 (N_5858,N_344,N_1979);
and U5859 (N_5859,N_2984,N_2257);
nand U5860 (N_5860,N_1866,N_1539);
or U5861 (N_5861,N_2226,N_2720);
and U5862 (N_5862,N_2168,N_252);
nor U5863 (N_5863,N_1932,N_2226);
nor U5864 (N_5864,N_1815,N_722);
and U5865 (N_5865,N_2382,N_2417);
and U5866 (N_5866,N_32,N_2417);
xor U5867 (N_5867,N_318,N_368);
xor U5868 (N_5868,N_478,N_613);
and U5869 (N_5869,N_1638,N_1804);
nand U5870 (N_5870,N_1117,N_2676);
or U5871 (N_5871,N_2154,N_2633);
and U5872 (N_5872,N_1444,N_1719);
nand U5873 (N_5873,N_1128,N_2128);
or U5874 (N_5874,N_1020,N_2853);
or U5875 (N_5875,N_2759,N_2108);
and U5876 (N_5876,N_2905,N_1237);
nor U5877 (N_5877,N_2139,N_227);
nor U5878 (N_5878,N_983,N_2473);
nand U5879 (N_5879,N_637,N_1725);
and U5880 (N_5880,N_448,N_926);
or U5881 (N_5881,N_2944,N_2433);
or U5882 (N_5882,N_2790,N_2397);
nor U5883 (N_5883,N_2944,N_616);
nor U5884 (N_5884,N_1648,N_2335);
or U5885 (N_5885,N_687,N_539);
nand U5886 (N_5886,N_1308,N_2632);
and U5887 (N_5887,N_1394,N_2208);
nor U5888 (N_5888,N_632,N_1340);
or U5889 (N_5889,N_1370,N_646);
nand U5890 (N_5890,N_1278,N_530);
nor U5891 (N_5891,N_1083,N_2804);
nand U5892 (N_5892,N_2786,N_2522);
or U5893 (N_5893,N_1891,N_1271);
nor U5894 (N_5894,N_2349,N_1999);
or U5895 (N_5895,N_1065,N_393);
or U5896 (N_5896,N_128,N_721);
nand U5897 (N_5897,N_2546,N_2749);
nand U5898 (N_5898,N_362,N_917);
or U5899 (N_5899,N_214,N_975);
or U5900 (N_5900,N_1754,N_2148);
and U5901 (N_5901,N_2337,N_1064);
and U5902 (N_5902,N_2681,N_1787);
xor U5903 (N_5903,N_674,N_1591);
or U5904 (N_5904,N_1920,N_1448);
and U5905 (N_5905,N_2683,N_1410);
and U5906 (N_5906,N_333,N_1813);
or U5907 (N_5907,N_575,N_1264);
nand U5908 (N_5908,N_2002,N_424);
and U5909 (N_5909,N_131,N_1509);
and U5910 (N_5910,N_2955,N_2513);
nor U5911 (N_5911,N_2290,N_1083);
and U5912 (N_5912,N_2880,N_1306);
nand U5913 (N_5913,N_1599,N_2866);
or U5914 (N_5914,N_82,N_1332);
and U5915 (N_5915,N_1873,N_2157);
nor U5916 (N_5916,N_1323,N_2662);
nor U5917 (N_5917,N_1104,N_1130);
nor U5918 (N_5918,N_1645,N_2760);
nand U5919 (N_5919,N_2169,N_311);
nor U5920 (N_5920,N_637,N_2250);
nor U5921 (N_5921,N_1597,N_2170);
nor U5922 (N_5922,N_1646,N_2040);
and U5923 (N_5923,N_107,N_751);
nor U5924 (N_5924,N_2241,N_216);
nor U5925 (N_5925,N_74,N_2380);
and U5926 (N_5926,N_1788,N_2528);
or U5927 (N_5927,N_2032,N_2831);
or U5928 (N_5928,N_1211,N_1548);
nor U5929 (N_5929,N_378,N_2042);
or U5930 (N_5930,N_2212,N_2189);
and U5931 (N_5931,N_2713,N_1351);
and U5932 (N_5932,N_1855,N_2848);
and U5933 (N_5933,N_699,N_1659);
nor U5934 (N_5934,N_1011,N_922);
and U5935 (N_5935,N_1138,N_199);
nand U5936 (N_5936,N_2295,N_1393);
nor U5937 (N_5937,N_907,N_587);
xnor U5938 (N_5938,N_846,N_2367);
and U5939 (N_5939,N_7,N_1959);
or U5940 (N_5940,N_2143,N_161);
nor U5941 (N_5941,N_783,N_1789);
and U5942 (N_5942,N_135,N_1000);
or U5943 (N_5943,N_2565,N_2496);
nor U5944 (N_5944,N_244,N_2747);
or U5945 (N_5945,N_742,N_1408);
nor U5946 (N_5946,N_854,N_385);
nor U5947 (N_5947,N_1690,N_174);
and U5948 (N_5948,N_1496,N_392);
nand U5949 (N_5949,N_350,N_2453);
or U5950 (N_5950,N_632,N_1954);
and U5951 (N_5951,N_1499,N_2660);
or U5952 (N_5952,N_273,N_645);
nor U5953 (N_5953,N_2144,N_1523);
nor U5954 (N_5954,N_2437,N_2841);
nor U5955 (N_5955,N_432,N_2063);
and U5956 (N_5956,N_507,N_294);
nand U5957 (N_5957,N_2585,N_85);
and U5958 (N_5958,N_2454,N_230);
and U5959 (N_5959,N_360,N_480);
nor U5960 (N_5960,N_1042,N_1209);
nand U5961 (N_5961,N_2838,N_175);
and U5962 (N_5962,N_678,N_1167);
nand U5963 (N_5963,N_1293,N_2638);
or U5964 (N_5964,N_916,N_129);
and U5965 (N_5965,N_2863,N_1932);
nand U5966 (N_5966,N_1072,N_164);
nand U5967 (N_5967,N_745,N_2880);
or U5968 (N_5968,N_953,N_2215);
or U5969 (N_5969,N_506,N_1825);
or U5970 (N_5970,N_1893,N_1031);
and U5971 (N_5971,N_238,N_2724);
nand U5972 (N_5972,N_1604,N_261);
nand U5973 (N_5973,N_2828,N_95);
and U5974 (N_5974,N_2343,N_1447);
nor U5975 (N_5975,N_263,N_1557);
nor U5976 (N_5976,N_1640,N_1613);
or U5977 (N_5977,N_2732,N_809);
nor U5978 (N_5978,N_1741,N_929);
nor U5979 (N_5979,N_181,N_1933);
or U5980 (N_5980,N_2911,N_289);
nor U5981 (N_5981,N_2661,N_756);
nor U5982 (N_5982,N_895,N_1909);
nand U5983 (N_5983,N_278,N_2215);
or U5984 (N_5984,N_2552,N_584);
nor U5985 (N_5985,N_1844,N_439);
nor U5986 (N_5986,N_493,N_178);
nor U5987 (N_5987,N_1658,N_1003);
nand U5988 (N_5988,N_2434,N_189);
and U5989 (N_5989,N_2665,N_35);
and U5990 (N_5990,N_1198,N_1977);
and U5991 (N_5991,N_58,N_2998);
and U5992 (N_5992,N_1138,N_437);
nand U5993 (N_5993,N_1248,N_2080);
nand U5994 (N_5994,N_1441,N_390);
or U5995 (N_5995,N_1879,N_1086);
nor U5996 (N_5996,N_1072,N_305);
or U5997 (N_5997,N_1517,N_1593);
or U5998 (N_5998,N_877,N_2623);
and U5999 (N_5999,N_997,N_339);
xor U6000 (N_6000,N_5079,N_3157);
and U6001 (N_6001,N_3238,N_5413);
nand U6002 (N_6002,N_3277,N_5613);
or U6003 (N_6003,N_3441,N_3496);
and U6004 (N_6004,N_4619,N_4422);
or U6005 (N_6005,N_5431,N_4686);
and U6006 (N_6006,N_3226,N_4902);
nand U6007 (N_6007,N_3819,N_4814);
nor U6008 (N_6008,N_4205,N_5879);
or U6009 (N_6009,N_3674,N_3993);
and U6010 (N_6010,N_3721,N_4250);
nand U6011 (N_6011,N_4363,N_5816);
and U6012 (N_6012,N_5632,N_3672);
or U6013 (N_6013,N_3710,N_4696);
and U6014 (N_6014,N_3874,N_3654);
nand U6015 (N_6015,N_3352,N_5030);
nor U6016 (N_6016,N_4770,N_5611);
nand U6017 (N_6017,N_5484,N_4340);
or U6018 (N_6018,N_4586,N_5565);
and U6019 (N_6019,N_4090,N_4197);
nand U6020 (N_6020,N_3377,N_4753);
nor U6021 (N_6021,N_3093,N_5767);
or U6022 (N_6022,N_4269,N_3535);
nor U6023 (N_6023,N_3625,N_3965);
nand U6024 (N_6024,N_3029,N_3776);
nor U6025 (N_6025,N_5150,N_3921);
nor U6026 (N_6026,N_4656,N_4628);
xnor U6027 (N_6027,N_4674,N_4783);
nor U6028 (N_6028,N_3188,N_3778);
xor U6029 (N_6029,N_3574,N_3709);
and U6030 (N_6030,N_3018,N_3459);
nor U6031 (N_6031,N_5369,N_5218);
or U6032 (N_6032,N_3952,N_3135);
nor U6033 (N_6033,N_5552,N_5324);
or U6034 (N_6034,N_4719,N_3065);
nor U6035 (N_6035,N_4798,N_3418);
nor U6036 (N_6036,N_4597,N_3026);
and U6037 (N_6037,N_4713,N_5537);
nor U6038 (N_6038,N_5846,N_5612);
xnor U6039 (N_6039,N_3376,N_3255);
nand U6040 (N_6040,N_3012,N_5931);
xor U6041 (N_6041,N_5837,N_5509);
or U6042 (N_6042,N_4987,N_4041);
nand U6043 (N_6043,N_5425,N_4716);
or U6044 (N_6044,N_5270,N_5661);
or U6045 (N_6045,N_3167,N_3390);
and U6046 (N_6046,N_3842,N_4694);
and U6047 (N_6047,N_5185,N_4795);
xor U6048 (N_6048,N_4106,N_3225);
or U6049 (N_6049,N_3798,N_4915);
nand U6050 (N_6050,N_4213,N_3306);
or U6051 (N_6051,N_4638,N_5576);
and U6052 (N_6052,N_5823,N_5800);
nand U6053 (N_6053,N_3683,N_5629);
nor U6054 (N_6054,N_4991,N_3178);
or U6055 (N_6055,N_4542,N_5455);
nor U6056 (N_6056,N_4605,N_5312);
or U6057 (N_6057,N_3967,N_4731);
and U6058 (N_6058,N_3177,N_5309);
or U6059 (N_6059,N_5551,N_5591);
or U6060 (N_6060,N_5797,N_3671);
or U6061 (N_6061,N_4048,N_5262);
nand U6062 (N_6062,N_5199,N_4938);
nand U6063 (N_6063,N_5464,N_4612);
nand U6064 (N_6064,N_3364,N_4773);
and U6065 (N_6065,N_5906,N_5119);
nor U6066 (N_6066,N_5021,N_5553);
or U6067 (N_6067,N_4979,N_3963);
or U6068 (N_6068,N_3885,N_3310);
nor U6069 (N_6069,N_3518,N_4644);
nand U6070 (N_6070,N_4543,N_3665);
nor U6071 (N_6071,N_3244,N_5922);
nand U6072 (N_6072,N_5014,N_3427);
or U6073 (N_6073,N_3525,N_4399);
or U6074 (N_6074,N_5265,N_3270);
nand U6075 (N_6075,N_4837,N_5794);
nand U6076 (N_6076,N_5725,N_3544);
nor U6077 (N_6077,N_5192,N_4920);
or U6078 (N_6078,N_3581,N_5409);
or U6079 (N_6079,N_4050,N_3969);
or U6080 (N_6080,N_4194,N_3351);
or U6081 (N_6081,N_3582,N_4917);
and U6082 (N_6082,N_4424,N_5514);
or U6083 (N_6083,N_4517,N_5515);
nand U6084 (N_6084,N_4342,N_3751);
or U6085 (N_6085,N_4116,N_5229);
and U6086 (N_6086,N_5886,N_5663);
and U6087 (N_6087,N_5709,N_4055);
nand U6088 (N_6088,N_5226,N_4409);
and U6089 (N_6089,N_5863,N_4959);
and U6090 (N_6090,N_3136,N_5257);
or U6091 (N_6091,N_4463,N_4956);
nand U6092 (N_6092,N_5224,N_3460);
nor U6093 (N_6093,N_5433,N_5850);
or U6094 (N_6094,N_3098,N_3328);
nor U6095 (N_6095,N_4357,N_3566);
nor U6096 (N_6096,N_4198,N_3103);
or U6097 (N_6097,N_3733,N_3162);
nor U6098 (N_6098,N_3901,N_3458);
nor U6099 (N_6099,N_4157,N_5996);
or U6100 (N_6100,N_4162,N_3298);
nand U6101 (N_6101,N_3747,N_4166);
xnor U6102 (N_6102,N_3023,N_5173);
or U6103 (N_6103,N_3895,N_3999);
and U6104 (N_6104,N_3402,N_5077);
xnor U6105 (N_6105,N_3449,N_4123);
or U6106 (N_6106,N_3595,N_4334);
xor U6107 (N_6107,N_3447,N_4602);
and U6108 (N_6108,N_5956,N_5743);
nor U6109 (N_6109,N_3156,N_5458);
nor U6110 (N_6110,N_4774,N_3773);
or U6111 (N_6111,N_4675,N_4679);
or U6112 (N_6112,N_5950,N_5750);
and U6113 (N_6113,N_5590,N_4436);
or U6114 (N_6114,N_3510,N_4385);
or U6115 (N_6115,N_4867,N_5721);
and U6116 (N_6116,N_4668,N_3913);
nor U6117 (N_6117,N_5081,N_5019);
nor U6118 (N_6118,N_4320,N_4819);
nand U6119 (N_6119,N_3176,N_4370);
and U6120 (N_6120,N_4152,N_5798);
nand U6121 (N_6121,N_3243,N_5035);
or U6122 (N_6122,N_5066,N_3825);
nor U6123 (N_6123,N_3196,N_3828);
nand U6124 (N_6124,N_3860,N_4038);
or U6125 (N_6125,N_5838,N_4164);
nor U6126 (N_6126,N_3557,N_4892);
or U6127 (N_6127,N_4231,N_3164);
nor U6128 (N_6128,N_4066,N_4986);
nor U6129 (N_6129,N_3658,N_3327);
and U6130 (N_6130,N_5404,N_4810);
or U6131 (N_6131,N_3320,N_4667);
nand U6132 (N_6132,N_3133,N_3884);
or U6133 (N_6133,N_5527,N_4144);
xor U6134 (N_6134,N_3573,N_4497);
and U6135 (N_6135,N_3900,N_4448);
nand U6136 (N_6136,N_4440,N_3384);
and U6137 (N_6137,N_5714,N_4715);
nand U6138 (N_6138,N_3618,N_3546);
or U6139 (N_6139,N_3565,N_4997);
nor U6140 (N_6140,N_4728,N_3564);
nor U6141 (N_6141,N_5271,N_4035);
nand U6142 (N_6142,N_4786,N_5008);
or U6143 (N_6143,N_3989,N_4528);
nand U6144 (N_6144,N_3934,N_4763);
and U6145 (N_6145,N_3732,N_3263);
nand U6146 (N_6146,N_5340,N_5542);
nand U6147 (N_6147,N_3251,N_4909);
nor U6148 (N_6148,N_3818,N_5386);
or U6149 (N_6149,N_5584,N_5341);
or U6150 (N_6150,N_5364,N_4598);
nor U6151 (N_6151,N_5116,N_5653);
nor U6152 (N_6152,N_4812,N_5272);
or U6153 (N_6153,N_3676,N_3533);
nor U6154 (N_6154,N_3631,N_4148);
nor U6155 (N_6155,N_5997,N_5052);
or U6156 (N_6156,N_5761,N_3219);
and U6157 (N_6157,N_3089,N_5827);
or U6158 (N_6158,N_5456,N_4530);
xor U6159 (N_6159,N_3706,N_5450);
or U6160 (N_6160,N_4913,N_4421);
and U6161 (N_6161,N_3511,N_5323);
nand U6162 (N_6162,N_4594,N_3448);
nand U6163 (N_6163,N_3583,N_3772);
and U6164 (N_6164,N_3703,N_4898);
and U6165 (N_6165,N_3001,N_3260);
and U6166 (N_6166,N_3570,N_5532);
nor U6167 (N_6167,N_3221,N_5697);
and U6168 (N_6168,N_3105,N_3222);
nor U6169 (N_6169,N_5964,N_4744);
nand U6170 (N_6170,N_5604,N_4985);
and U6171 (N_6171,N_4373,N_5546);
or U6172 (N_6172,N_5525,N_3757);
nor U6173 (N_6173,N_4304,N_4172);
nor U6174 (N_6174,N_5040,N_4721);
and U6175 (N_6175,N_5786,N_4631);
nor U6176 (N_6176,N_4725,N_4151);
and U6177 (N_6177,N_4040,N_5680);
and U6178 (N_6178,N_4627,N_3047);
nand U6179 (N_6179,N_5111,N_4435);
and U6180 (N_6180,N_5062,N_4473);
nor U6181 (N_6181,N_4397,N_4047);
and U6182 (N_6182,N_5094,N_3370);
and U6183 (N_6183,N_3291,N_4647);
nand U6184 (N_6184,N_3727,N_3561);
or U6185 (N_6185,N_3958,N_5275);
nor U6186 (N_6186,N_5910,N_4345);
nor U6187 (N_6187,N_4268,N_3633);
and U6188 (N_6188,N_4792,N_3062);
nor U6189 (N_6189,N_4838,N_5160);
or U6190 (N_6190,N_5004,N_3144);
nor U6191 (N_6191,N_4722,N_4886);
or U6192 (N_6192,N_3037,N_4097);
and U6193 (N_6193,N_3899,N_3229);
and U6194 (N_6194,N_5089,N_4811);
and U6195 (N_6195,N_3013,N_4200);
and U6196 (N_6196,N_5740,N_3610);
or U6197 (N_6197,N_3455,N_4236);
nor U6198 (N_6198,N_4365,N_5999);
and U6199 (N_6199,N_3630,N_4566);
nand U6200 (N_6200,N_5822,N_3181);
or U6201 (N_6201,N_4177,N_4489);
nand U6202 (N_6202,N_5874,N_4564);
and U6203 (N_6203,N_3354,N_3638);
and U6204 (N_6204,N_4141,N_4953);
or U6205 (N_6205,N_4962,N_5443);
nand U6206 (N_6206,N_4046,N_5320);
and U6207 (N_6207,N_5943,N_4622);
and U6208 (N_6208,N_3278,N_3262);
or U6209 (N_6209,N_4547,N_4687);
and U6210 (N_6210,N_5353,N_3962);
and U6211 (N_6211,N_5934,N_5766);
or U6212 (N_6212,N_3143,N_3560);
and U6213 (N_6213,N_4681,N_4544);
nor U6214 (N_6214,N_3168,N_4709);
and U6215 (N_6215,N_4673,N_5292);
and U6216 (N_6216,N_3669,N_3163);
nand U6217 (N_6217,N_5238,N_3623);
nor U6218 (N_6218,N_3466,N_3141);
nor U6219 (N_6219,N_3695,N_4394);
and U6220 (N_6220,N_5967,N_4242);
nor U6221 (N_6221,N_4636,N_5621);
and U6222 (N_6222,N_4036,N_3571);
nor U6223 (N_6223,N_5673,N_5523);
nor U6224 (N_6224,N_5401,N_5940);
nor U6225 (N_6225,N_5361,N_3737);
or U6226 (N_6226,N_3759,N_4367);
and U6227 (N_6227,N_5311,N_5316);
nor U6228 (N_6228,N_3073,N_3283);
nand U6229 (N_6229,N_3128,N_3827);
nand U6230 (N_6230,N_5083,N_5881);
nand U6231 (N_6231,N_5171,N_5009);
or U6232 (N_6232,N_4767,N_4910);
and U6233 (N_6233,N_4764,N_3381);
nand U6234 (N_6234,N_5826,N_4623);
nand U6235 (N_6235,N_5255,N_5435);
and U6236 (N_6236,N_5451,N_4477);
nor U6237 (N_6237,N_3649,N_5109);
and U6238 (N_6238,N_5903,N_3102);
xor U6239 (N_6239,N_4456,N_3451);
nand U6240 (N_6240,N_3894,N_4119);
and U6241 (N_6241,N_5560,N_3010);
or U6242 (N_6242,N_4387,N_3517);
and U6243 (N_6243,N_5503,N_4089);
nor U6244 (N_6244,N_5318,N_3567);
xnor U6245 (N_6245,N_4330,N_5500);
nor U6246 (N_6246,N_5860,N_3300);
and U6247 (N_6247,N_5317,N_4759);
or U6248 (N_6248,N_3982,N_3304);
nand U6249 (N_6249,N_4691,N_4318);
and U6250 (N_6250,N_4347,N_3534);
and U6251 (N_6251,N_5246,N_5832);
nand U6252 (N_6252,N_5402,N_4068);
nor U6253 (N_6253,N_3216,N_5923);
nand U6254 (N_6254,N_5988,N_5396);
nor U6255 (N_6255,N_3456,N_4850);
or U6256 (N_6256,N_3104,N_5876);
nand U6257 (N_6257,N_4768,N_4961);
and U6258 (N_6258,N_4740,N_3284);
nor U6259 (N_6259,N_3175,N_5908);
nor U6260 (N_6260,N_3584,N_3323);
and U6261 (N_6261,N_5828,N_3948);
nand U6262 (N_6262,N_4265,N_5681);
or U6263 (N_6263,N_4897,N_3598);
and U6264 (N_6264,N_4929,N_4806);
nor U6265 (N_6265,N_5189,N_5958);
and U6266 (N_6266,N_3285,N_5985);
nor U6267 (N_6267,N_4896,N_4008);
and U6268 (N_6268,N_3033,N_4610);
or U6269 (N_6269,N_5266,N_5424);
or U6270 (N_6270,N_5061,N_4014);
and U6271 (N_6271,N_4800,N_3097);
and U6272 (N_6272,N_4158,N_4229);
or U6273 (N_6273,N_4255,N_3954);
or U6274 (N_6274,N_5533,N_3562);
nand U6275 (N_6275,N_4939,N_4076);
or U6276 (N_6276,N_4498,N_4491);
nor U6277 (N_6277,N_3522,N_3042);
nand U6278 (N_6278,N_4053,N_4904);
and U6279 (N_6279,N_3739,N_4429);
or U6280 (N_6280,N_5907,N_3927);
nor U6281 (N_6281,N_3760,N_3212);
and U6282 (N_6282,N_3118,N_5891);
and U6283 (N_6283,N_5344,N_5268);
nor U6284 (N_6284,N_4824,N_3987);
nand U6285 (N_6285,N_5148,N_5734);
and U6286 (N_6286,N_4259,N_5780);
and U6287 (N_6287,N_4003,N_4678);
xnor U6288 (N_6288,N_5479,N_5519);
nor U6289 (N_6289,N_5279,N_5407);
nand U6290 (N_6290,N_3789,N_4510);
nor U6291 (N_6291,N_4879,N_5904);
or U6292 (N_6292,N_4572,N_4512);
and U6293 (N_6293,N_4181,N_3258);
or U6294 (N_6294,N_4227,N_4741);
nor U6295 (N_6295,N_4472,N_3980);
nor U6296 (N_6296,N_4327,N_4112);
nor U6297 (N_6297,N_4126,N_5785);
and U6298 (N_6298,N_5890,N_4735);
nand U6299 (N_6299,N_3101,N_3691);
nor U6300 (N_6300,N_3984,N_4595);
xnor U6301 (N_6301,N_3811,N_5788);
nand U6302 (N_6302,N_4273,N_3768);
or U6303 (N_6303,N_4883,N_3990);
and U6304 (N_6304,N_4964,N_5773);
nand U6305 (N_6305,N_5383,N_4588);
and U6306 (N_6306,N_3752,N_5921);
and U6307 (N_6307,N_5625,N_4955);
and U6308 (N_6308,N_5650,N_3675);
nand U6309 (N_6309,N_3485,N_4377);
xor U6310 (N_6310,N_4529,N_5884);
xnor U6311 (N_6311,N_3765,N_4178);
or U6312 (N_6312,N_3315,N_5535);
nor U6313 (N_6313,N_4880,N_3646);
or U6314 (N_6314,N_4493,N_5772);
and U6315 (N_6315,N_5472,N_3854);
nor U6316 (N_6316,N_5713,N_4091);
nand U6317 (N_6317,N_5656,N_5108);
or U6318 (N_6318,N_3594,N_4682);
nor U6319 (N_6319,N_3408,N_3746);
nor U6320 (N_6320,N_4305,N_4616);
nor U6321 (N_6321,N_3079,N_5962);
or U6322 (N_6322,N_4190,N_5712);
nor U6323 (N_6323,N_5841,N_3410);
or U6324 (N_6324,N_5616,N_5559);
or U6325 (N_6325,N_5372,N_4858);
or U6326 (N_6326,N_5412,N_5952);
nand U6327 (N_6327,N_4195,N_5840);
nand U6328 (N_6328,N_4965,N_4807);
or U6329 (N_6329,N_4717,N_4996);
and U6330 (N_6330,N_5360,N_5038);
nand U6331 (N_6331,N_3530,N_3849);
or U6332 (N_6332,N_4012,N_3488);
or U6333 (N_6333,N_4534,N_3876);
nand U6334 (N_6334,N_3555,N_3605);
and U6335 (N_6335,N_4051,N_5454);
nand U6336 (N_6336,N_4702,N_5287);
nor U6337 (N_6337,N_5313,N_5668);
or U6338 (N_6338,N_3689,N_4835);
nor U6339 (N_6339,N_4065,N_3856);
and U6340 (N_6340,N_5134,N_3422);
and U6341 (N_6341,N_5034,N_3115);
nand U6342 (N_6342,N_4462,N_5099);
or U6343 (N_6343,N_3426,N_4300);
or U6344 (N_6344,N_4058,N_5015);
nand U6345 (N_6345,N_5677,N_3325);
and U6346 (N_6346,N_3777,N_5544);
nor U6347 (N_6347,N_4587,N_3545);
nor U6348 (N_6348,N_5593,N_4270);
xor U6349 (N_6349,N_3763,N_5504);
nand U6350 (N_6350,N_5487,N_3066);
and U6351 (N_6351,N_4211,N_3099);
nand U6352 (N_6352,N_3119,N_5894);
and U6353 (N_6353,N_5184,N_4614);
and U6354 (N_6354,N_4427,N_4700);
and U6355 (N_6355,N_5288,N_3558);
or U6356 (N_6356,N_3968,N_4998);
nand U6357 (N_6357,N_5736,N_5441);
and U6358 (N_6358,N_3694,N_4108);
or U6359 (N_6359,N_4176,N_5421);
or U6360 (N_6360,N_4568,N_3592);
or U6361 (N_6361,N_3724,N_3000);
or U6362 (N_6362,N_3614,N_3180);
nand U6363 (N_6363,N_3866,N_3959);
nand U6364 (N_6364,N_4626,N_5483);
nand U6365 (N_6365,N_3486,N_5623);
nand U6366 (N_6366,N_4930,N_3915);
nand U6367 (N_6367,N_5687,N_5346);
nand U6368 (N_6368,N_4787,N_5252);
or U6369 (N_6369,N_4086,N_5334);
xor U6370 (N_6370,N_3941,N_3750);
nor U6371 (N_6371,N_3392,N_4083);
and U6372 (N_6372,N_3344,N_4978);
and U6373 (N_6373,N_4620,N_5147);
or U6374 (N_6374,N_5011,N_5058);
nand U6375 (N_6375,N_3085,N_3740);
or U6376 (N_6376,N_3813,N_4856);
nor U6377 (N_6377,N_4027,N_3815);
or U6378 (N_6378,N_4400,N_4968);
and U6379 (N_6379,N_4125,N_3312);
and U6380 (N_6380,N_5332,N_5852);
and U6381 (N_6381,N_4074,N_5641);
nor U6382 (N_6382,N_5810,N_4201);
nor U6383 (N_6383,N_3139,N_3621);
and U6384 (N_6384,N_5044,N_4037);
and U6385 (N_6385,N_5831,N_3906);
and U6386 (N_6386,N_5135,N_5573);
and U6387 (N_6387,N_3972,N_5654);
nor U6388 (N_6388,N_5121,N_4481);
and U6389 (N_6389,N_4827,N_3076);
xor U6390 (N_6390,N_3052,N_4437);
nand U6391 (N_6391,N_4779,N_5662);
or U6392 (N_6392,N_4445,N_5902);
nand U6393 (N_6393,N_4079,N_5315);
and U6394 (N_6394,N_3870,N_3231);
and U6395 (N_6395,N_4004,N_3109);
or U6396 (N_6396,N_3536,N_4360);
nor U6397 (N_6397,N_3563,N_3853);
nor U6398 (N_6398,N_4718,N_5337);
or U6399 (N_6399,N_5209,N_3786);
or U6400 (N_6400,N_3539,N_3430);
nand U6401 (N_6401,N_5351,N_3235);
nor U6402 (N_6402,N_5737,N_4624);
nor U6403 (N_6403,N_5665,N_4852);
nor U6404 (N_6404,N_5670,N_3892);
and U6405 (N_6405,N_5133,N_3577);
nand U6406 (N_6406,N_5374,N_3607);
and U6407 (N_6407,N_3356,N_3494);
or U6408 (N_6408,N_4532,N_5578);
or U6409 (N_6409,N_5060,N_3753);
or U6410 (N_6410,N_5363,N_5541);
xor U6411 (N_6411,N_5664,N_5088);
nand U6412 (N_6412,N_5003,N_5319);
or U6413 (N_6413,N_3034,N_3788);
or U6414 (N_6414,N_5177,N_4967);
nand U6415 (N_6415,N_4020,N_5580);
and U6416 (N_6416,N_5124,N_5103);
nor U6417 (N_6417,N_4271,N_5093);
and U6418 (N_6418,N_4441,N_5195);
or U6419 (N_6419,N_5954,N_4969);
nand U6420 (N_6420,N_4911,N_5774);
and U6421 (N_6421,N_4793,N_5916);
nand U6422 (N_6422,N_3730,N_3891);
nand U6423 (N_6423,N_5779,N_4414);
and U6424 (N_6424,N_3249,N_3396);
nor U6425 (N_6425,N_4482,N_4567);
nand U6426 (N_6426,N_4748,N_3161);
and U6427 (N_6427,N_4220,N_3795);
or U6428 (N_6428,N_4021,N_4524);
nor U6429 (N_6429,N_4278,N_5624);
nand U6430 (N_6430,N_5408,N_4903);
and U6431 (N_6431,N_3922,N_3311);
and U6432 (N_6432,N_3083,N_4285);
or U6433 (N_6433,N_5100,N_4546);
nor U6434 (N_6434,N_4193,N_5990);
nand U6435 (N_6435,N_3933,N_4557);
or U6436 (N_6436,N_5204,N_4840);
nand U6437 (N_6437,N_3925,N_3121);
nor U6438 (N_6438,N_3480,N_5101);
nor U6439 (N_6439,N_4695,N_5684);
and U6440 (N_6440,N_5130,N_4444);
nand U6441 (N_6441,N_4488,N_5178);
nor U6442 (N_6442,N_3883,N_4196);
nor U6443 (N_6443,N_4833,N_5814);
nand U6444 (N_6444,N_5545,N_4452);
and U6445 (N_6445,N_3829,N_3991);
nor U6446 (N_6446,N_3888,N_3366);
and U6447 (N_6447,N_5889,N_5227);
nor U6448 (N_6448,N_3762,N_5154);
nor U6449 (N_6449,N_3971,N_3679);
nor U6450 (N_6450,N_5742,N_4309);
or U6451 (N_6451,N_4379,N_3322);
nor U6452 (N_6452,N_5595,N_4140);
nor U6453 (N_6453,N_5300,N_4752);
or U6454 (N_6454,N_4854,N_4573);
nand U6455 (N_6455,N_4013,N_5352);
nand U6456 (N_6456,N_3148,N_4705);
and U6457 (N_6457,N_3371,N_3514);
nand U6458 (N_6458,N_3650,N_3401);
and U6459 (N_6459,N_3158,N_3660);
and U6460 (N_6460,N_4789,N_5187);
or U6461 (N_6461,N_3008,N_4077);
or U6462 (N_6462,N_3857,N_3443);
and U6463 (N_6463,N_3245,N_5702);
nor U6464 (N_6464,N_4611,N_5834);
or U6465 (N_6465,N_4104,N_5260);
or U6466 (N_6466,N_5550,N_3149);
or U6467 (N_6467,N_5068,N_4933);
and U6468 (N_6468,N_3345,N_4416);
nor U6469 (N_6469,N_5070,N_3326);
nor U6470 (N_6470,N_5603,N_4168);
nor U6471 (N_6471,N_5717,N_4353);
nor U6472 (N_6472,N_4252,N_3420);
and U6473 (N_6473,N_3836,N_4299);
nand U6474 (N_6474,N_5864,N_5302);
nand U6475 (N_6475,N_3930,N_4266);
xnor U6476 (N_6476,N_5636,N_5280);
or U6477 (N_6477,N_3412,N_5770);
or U6478 (N_6478,N_5416,N_3804);
nand U6479 (N_6479,N_5769,N_3334);
and U6480 (N_6480,N_4492,N_5065);
nand U6481 (N_6481,N_4290,N_5293);
and U6482 (N_6482,N_3796,N_5283);
nor U6483 (N_6483,N_3682,N_5887);
nand U6484 (N_6484,N_5146,N_4672);
and U6485 (N_6485,N_4582,N_4727);
or U6486 (N_6486,N_5866,N_5120);
nand U6487 (N_6487,N_4160,N_5201);
or U6488 (N_6488,N_5858,N_4212);
nor U6489 (N_6489,N_4433,N_4683);
and U6490 (N_6490,N_4857,N_4254);
and U6491 (N_6491,N_3230,N_4350);
and U6492 (N_6492,N_3191,N_5675);
and U6493 (N_6493,N_5805,N_4155);
nand U6494 (N_6494,N_5149,N_4889);
nor U6495 (N_6495,N_3194,N_4135);
nand U6496 (N_6496,N_5434,N_5251);
or U6497 (N_6497,N_4006,N_4960);
nand U6498 (N_6498,N_4335,N_5781);
nor U6499 (N_6499,N_5029,N_5753);
or U6500 (N_6500,N_4453,N_3280);
nand U6501 (N_6501,N_5543,N_4584);
or U6502 (N_6502,N_3692,N_5426);
nor U6503 (N_6503,N_3021,N_3006);
nor U6504 (N_6504,N_4082,N_4388);
or U6505 (N_6505,N_3523,N_4408);
nand U6506 (N_6506,N_5505,N_3908);
nand U6507 (N_6507,N_4561,N_4559);
nand U6508 (N_6508,N_3252,N_4571);
or U6509 (N_6509,N_4670,N_4368);
xnor U6510 (N_6510,N_3718,N_3869);
and U6511 (N_6511,N_3032,N_3716);
nor U6512 (N_6512,N_3951,N_3516);
nor U6513 (N_6513,N_4025,N_5107);
nand U6514 (N_6514,N_4689,N_3587);
xnor U6515 (N_6515,N_3423,N_5801);
nor U6516 (N_6516,N_3602,N_5222);
or U6517 (N_6517,N_5127,N_5754);
and U6518 (N_6518,N_5200,N_3187);
and U6519 (N_6519,N_5521,N_5465);
nand U6520 (N_6520,N_5606,N_4832);
or U6521 (N_6521,N_5699,N_4846);
nor U6522 (N_6522,N_3970,N_3182);
nand U6523 (N_6523,N_4224,N_5411);
and U6524 (N_6524,N_4519,N_3205);
and U6525 (N_6525,N_5017,N_4156);
or U6526 (N_6526,N_4465,N_4049);
nor U6527 (N_6527,N_3484,N_3785);
nand U6528 (N_6528,N_5295,N_5870);
or U6529 (N_6529,N_4071,N_4099);
nand U6530 (N_6530,N_3299,N_3040);
or U6531 (N_6531,N_5626,N_3465);
nor U6532 (N_6532,N_5914,N_5759);
and U6533 (N_6533,N_4118,N_3996);
or U6534 (N_6534,N_3388,N_4147);
or U6535 (N_6535,N_5583,N_3506);
and U6536 (N_6536,N_5165,N_5979);
nand U6537 (N_6537,N_5691,N_4355);
or U6538 (N_6538,N_5384,N_5984);
nor U6539 (N_6539,N_3368,N_4260);
nand U6540 (N_6540,N_3549,N_4336);
and U6541 (N_6541,N_4502,N_5232);
and U6542 (N_6542,N_3792,N_5269);
or U6543 (N_6543,N_4217,N_5473);
nor U6544 (N_6544,N_3513,N_4230);
or U6545 (N_6545,N_5562,N_4927);
nand U6546 (N_6546,N_3347,N_4684);
and U6547 (N_6547,N_4790,N_4874);
and U6548 (N_6548,N_5649,N_4218);
and U6549 (N_6549,N_5137,N_3078);
nand U6550 (N_6550,N_4894,N_3080);
nand U6551 (N_6551,N_5857,N_4576);
nor U6552 (N_6552,N_5186,N_4639);
nand U6553 (N_6553,N_3835,N_4699);
or U6554 (N_6554,N_4096,N_3190);
and U6555 (N_6555,N_4851,N_3521);
nand U6556 (N_6556,N_4383,N_5694);
or U6557 (N_6557,N_5470,N_3379);
or U6558 (N_6558,N_3024,N_4301);
nor U6559 (N_6559,N_3628,N_5811);
nand U6560 (N_6560,N_5291,N_5256);
and U6561 (N_6561,N_5610,N_5516);
nand U6562 (N_6562,N_5428,N_5955);
and U6563 (N_6563,N_4081,N_4966);
or U6564 (N_6564,N_5878,N_3454);
nand U6565 (N_6565,N_3005,N_4295);
nand U6566 (N_6566,N_5486,N_3246);
or U6567 (N_6567,N_3002,N_5276);
or U6568 (N_6568,N_5946,N_4420);
nand U6569 (N_6569,N_5506,N_3250);
nor U6570 (N_6570,N_4362,N_5928);
and U6571 (N_6571,N_5719,N_4591);
and U6572 (N_6572,N_3684,N_5607);
xor U6573 (N_6573,N_5924,N_4474);
or U6574 (N_6574,N_5157,N_3738);
and U6575 (N_6575,N_5259,N_4188);
and U6576 (N_6576,N_4232,N_3593);
or U6577 (N_6577,N_5775,N_4593);
or U6578 (N_6578,N_5410,N_3914);
and U6579 (N_6579,N_3613,N_4483);
and U6580 (N_6580,N_3220,N_3247);
or U6581 (N_6581,N_3949,N_5651);
nor U6582 (N_6582,N_5873,N_4450);
or U6583 (N_6583,N_5882,N_3224);
nand U6584 (N_6584,N_4797,N_5748);
or U6585 (N_6585,N_3697,N_3049);
or U6586 (N_6586,N_5203,N_4554);
and U6587 (N_6587,N_4940,N_4971);
and U6588 (N_6588,N_5480,N_4815);
and U6589 (N_6589,N_5056,N_5110);
xor U6590 (N_6590,N_3011,N_5143);
nor U6591 (N_6591,N_3604,N_5972);
or U6592 (N_6592,N_5809,N_3140);
and U6593 (N_6593,N_3569,N_5715);
or U6594 (N_6594,N_3124,N_3112);
and U6595 (N_6595,N_4901,N_4043);
nor U6596 (N_6596,N_3767,N_5652);
nor U6597 (N_6597,N_3897,N_3729);
nor U6598 (N_6598,N_5478,N_4803);
and U6599 (N_6599,N_5983,N_5485);
nor U6600 (N_6600,N_5631,N_3917);
nand U6601 (N_6601,N_5329,N_5420);
nand U6602 (N_6602,N_5290,N_3286);
and U6603 (N_6603,N_5114,N_4022);
or U6604 (N_6604,N_5898,N_3663);
nor U6605 (N_6605,N_3039,N_3482);
nand U6606 (N_6606,N_4402,N_4992);
and U6607 (N_6607,N_3383,N_3976);
or U6608 (N_6608,N_3463,N_5937);
nor U6609 (N_6609,N_5151,N_5893);
nand U6610 (N_6610,N_4257,N_5824);
and U6611 (N_6611,N_5328,N_4887);
nor U6612 (N_6612,N_3348,N_3554);
and U6613 (N_6613,N_4957,N_5461);
or U6614 (N_6614,N_3071,N_5020);
nor U6615 (N_6615,N_5273,N_4495);
and U6616 (N_6616,N_4742,N_3816);
and U6617 (N_6617,N_4671,N_3872);
and U6618 (N_6618,N_4146,N_5024);
nand U6619 (N_6619,N_4931,N_4629);
or U6620 (N_6620,N_3830,N_5529);
or U6621 (N_6621,N_3515,N_5138);
and U6622 (N_6622,N_4319,N_5929);
xor U6623 (N_6623,N_4475,N_5998);
xnor U6624 (N_6624,N_4977,N_5342);
or U6625 (N_6625,N_3468,N_4539);
and U6626 (N_6626,N_5054,N_5987);
nor U6627 (N_6627,N_3537,N_5236);
nand U6628 (N_6628,N_3077,N_4507);
nand U6629 (N_6629,N_3425,N_5045);
nand U6630 (N_6630,N_4520,N_5724);
nor U6631 (N_6631,N_4186,N_5571);
nand U6632 (N_6632,N_4199,N_4221);
nor U6633 (N_6633,N_4248,N_5414);
or U6634 (N_6634,N_5234,N_4853);
nand U6635 (N_6635,N_3453,N_4970);
or U6636 (N_6636,N_4828,N_5063);
or U6637 (N_6637,N_3450,N_5856);
nand U6638 (N_6638,N_4413,N_3321);
nor U6639 (N_6639,N_5885,N_3084);
or U6640 (N_6640,N_3068,N_5370);
nor U6641 (N_6641,N_5791,N_5638);
and U6642 (N_6642,N_3781,N_3169);
and U6643 (N_6643,N_5043,N_5690);
nor U6644 (N_6644,N_5371,N_4263);
nand U6645 (N_6645,N_4757,N_5513);
nand U6646 (N_6646,N_5572,N_4258);
nand U6647 (N_6647,N_4348,N_3945);
or U6648 (N_6648,N_4117,N_3265);
nand U6649 (N_6649,N_3009,N_4167);
nand U6650 (N_6650,N_5917,N_3146);
or U6651 (N_6651,N_5689,N_4974);
and U6652 (N_6652,N_5655,N_4608);
nor U6653 (N_6653,N_3058,N_4447);
or U6654 (N_6654,N_4805,N_3501);
nand U6655 (N_6655,N_3117,N_3597);
nor U6656 (N_6656,N_4249,N_4664);
or U6657 (N_6657,N_3154,N_4105);
or U6658 (N_6658,N_3038,N_5216);
or U6659 (N_6659,N_3414,N_3957);
nor U6660 (N_6660,N_4877,N_4378);
nand U6661 (N_6661,N_3395,N_4237);
nor U6662 (N_6662,N_5577,N_5327);
or U6663 (N_6663,N_3210,N_3269);
xnor U6664 (N_6664,N_4150,N_4338);
nor U6665 (N_6665,N_5193,N_5096);
nor U6666 (N_6666,N_3467,N_5074);
or U6667 (N_6667,N_4948,N_3608);
nand U6668 (N_6668,N_5264,N_4688);
nor U6669 (N_6669,N_3030,N_3807);
and U6670 (N_6670,N_5225,N_4100);
nand U6671 (N_6671,N_3868,N_3391);
nand U6672 (N_6672,N_3590,N_3992);
and U6673 (N_6673,N_3926,N_4372);
or U6674 (N_6674,N_5395,N_5392);
or U6675 (N_6675,N_5326,N_3775);
and U6676 (N_6676,N_3475,N_5672);
nor U6677 (N_6677,N_3997,N_5037);
or U6678 (N_6678,N_4129,N_5862);
nand U6679 (N_6679,N_4802,N_4359);
nor U6680 (N_6680,N_5385,N_4458);
nor U6681 (N_6681,N_5499,N_5530);
and U6682 (N_6682,N_5139,N_5618);
nand U6683 (N_6683,N_3601,N_5422);
and U6684 (N_6684,N_3407,N_5711);
nor U6685 (N_6685,N_4294,N_4486);
nor U6686 (N_6686,N_5049,N_3020);
or U6687 (N_6687,N_4663,N_3708);
nor U6688 (N_6688,N_4459,N_4891);
nand U6689 (N_6689,N_3611,N_4692);
nor U6690 (N_6690,N_4669,N_5498);
or U6691 (N_6691,N_5048,N_3147);
nor U6692 (N_6692,N_3406,N_5977);
or U6693 (N_6693,N_5930,N_5016);
nor U6694 (N_6694,N_4120,N_5732);
or U6695 (N_6695,N_3203,N_5892);
nand U6696 (N_6696,N_5883,N_4093);
nand U6697 (N_6697,N_3288,N_5208);
and U6698 (N_6698,N_3036,N_3626);
and U6699 (N_6699,N_5911,N_5175);
or U6700 (N_6700,N_5253,N_3208);
nor U6701 (N_6701,N_4000,N_5796);
nand U6702 (N_6702,N_3677,N_4207);
nand U6703 (N_6703,N_5131,N_4711);
and U6704 (N_6704,N_5627,N_5566);
and U6705 (N_6705,N_3821,N_5646);
and U6706 (N_6706,N_5469,N_3699);
nand U6707 (N_6707,N_5102,N_3844);
or U6708 (N_6708,N_5783,N_4311);
and U6709 (N_6709,N_4697,N_4386);
nand U6710 (N_6710,N_5118,N_4829);
nand U6711 (N_6711,N_4778,N_5637);
nand U6712 (N_6712,N_3940,N_3960);
or U6713 (N_6713,N_3882,N_4039);
or U6714 (N_6714,N_3896,N_4743);
or U6715 (N_6715,N_5071,N_5555);
and U6716 (N_6716,N_4973,N_4023);
and U6717 (N_6717,N_5818,N_3127);
nor U6718 (N_6718,N_4600,N_4822);
nand U6719 (N_6719,N_3054,N_5695);
nand U6720 (N_6720,N_4240,N_4900);
nand U6721 (N_6721,N_4575,N_3275);
nor U6722 (N_6722,N_4698,N_5104);
nand U6723 (N_6723,N_4907,N_3832);
nand U6724 (N_6724,N_3648,N_3134);
or U6725 (N_6725,N_5419,N_3031);
and U6726 (N_6726,N_3859,N_4316);
nand U6727 (N_6727,N_5741,N_5475);
or U6728 (N_6728,N_3108,N_3074);
and U6729 (N_6729,N_3509,N_4754);
nand U6730 (N_6730,N_4823,N_4426);
xor U6731 (N_6731,N_4411,N_4331);
and U6732 (N_6732,N_3159,N_3839);
or U6733 (N_6733,N_4860,N_3579);
nor U6734 (N_6734,N_3698,N_5678);
or U6735 (N_6735,N_5871,N_3340);
and U6736 (N_6736,N_3110,N_4756);
or U6737 (N_6737,N_5156,N_3749);
and U6738 (N_6738,N_3680,N_5880);
nand U6739 (N_6739,N_5900,N_5284);
nor U6740 (N_6740,N_4549,N_5161);
nor U6741 (N_6741,N_3655,N_4975);
and U6742 (N_6742,N_5706,N_4558);
nor U6743 (N_6743,N_4134,N_5949);
nand U6744 (N_6744,N_3918,N_5586);
and U6745 (N_6745,N_4603,N_5875);
nand U6746 (N_6746,N_4073,N_5112);
or U6747 (N_6747,N_4113,N_3861);
nor U6748 (N_6748,N_5526,N_3589);
nand U6749 (N_6749,N_4932,N_4026);
nand U6750 (N_6750,N_3666,N_5909);
and U6751 (N_6751,N_3981,N_3685);
nor U6752 (N_6752,N_5918,N_5554);
and U6753 (N_6753,N_3600,N_5989);
or U6754 (N_6754,N_3389,N_4659);
nand U6755 (N_6755,N_3090,N_4655);
and U6756 (N_6756,N_5405,N_4601);
nand U6757 (N_6757,N_4281,N_5596);
nand U6758 (N_6758,N_3254,N_3342);
and U6759 (N_6759,N_3490,N_4375);
or U6760 (N_6760,N_3428,N_3637);
or U6761 (N_6761,N_5481,N_5688);
nor U6762 (N_6762,N_5582,N_3817);
nor U6763 (N_6763,N_5338,N_3553);
and U6764 (N_6764,N_4505,N_4951);
nand U6765 (N_6765,N_3919,N_3820);
nand U6766 (N_6766,N_4982,N_4439);
nand U6767 (N_6767,N_5540,N_5659);
and U6768 (N_6768,N_5982,N_3845);
nand U6769 (N_6769,N_5219,N_3100);
nor U6770 (N_6770,N_5033,N_3358);
and U6771 (N_6771,N_5387,N_5467);
nor U6772 (N_6772,N_4471,N_4862);
nor U6773 (N_6773,N_4253,N_3838);
xnor U6774 (N_6774,N_5764,N_5833);
or U6775 (N_6775,N_5230,N_4428);
nand U6776 (N_6776,N_4346,N_5927);
or U6777 (N_6777,N_4132,N_5855);
or U6778 (N_6778,N_3580,N_5073);
or U6779 (N_6779,N_4138,N_4243);
and U6780 (N_6780,N_3802,N_5807);
nor U6781 (N_6781,N_4830,N_3924);
or U6782 (N_6782,N_5176,N_4949);
or U6783 (N_6783,N_3120,N_5491);
xor U6784 (N_6784,N_4127,N_5084);
or U6785 (N_6785,N_5630,N_4816);
nor U6786 (N_6786,N_3887,N_4264);
nor U6787 (N_6787,N_5459,N_4490);
and U6788 (N_6788,N_4288,N_5600);
and U6789 (N_6789,N_4485,N_4054);
nor U6790 (N_6790,N_4369,N_4358);
nand U6791 (N_6791,N_4890,N_5602);
nand U6792 (N_6792,N_4925,N_4443);
nand U6793 (N_6793,N_3378,N_4599);
nand U6794 (N_6794,N_4749,N_4553);
nor U6795 (N_6795,N_5538,N_4511);
xor U6796 (N_6796,N_3153,N_3619);
nand U6797 (N_6797,N_4454,N_3242);
nand U6798 (N_6798,N_3979,N_5399);
or U6799 (N_6799,N_3943,N_5365);
or U6800 (N_6800,N_4596,N_4914);
and U6801 (N_6801,N_4449,N_4396);
and U6802 (N_6802,N_3297,N_4583);
nand U6803 (N_6803,N_3442,N_5676);
nand U6804 (N_6804,N_5298,N_5683);
or U6805 (N_6805,N_4761,N_5836);
xor U6806 (N_6806,N_4522,N_3130);
and U6807 (N_6807,N_4746,N_3022);
nor U6808 (N_6808,N_4562,N_5128);
nor U6809 (N_6809,N_5418,N_4494);
nand U6810 (N_6810,N_4801,N_3664);
nand U6811 (N_6811,N_5403,N_4680);
nor U6812 (N_6812,N_3335,N_3476);
and U6813 (N_6813,N_4315,N_3902);
nor U6814 (N_6814,N_3847,N_5053);
nor U6815 (N_6815,N_5777,N_3556);
nor U6816 (N_6816,N_5793,N_3893);
and U6817 (N_6817,N_4314,N_5944);
nor U6818 (N_6818,N_5406,N_5547);
nor U6819 (N_6819,N_5397,N_4908);
nor U6820 (N_6820,N_4349,N_4095);
nor U6821 (N_6821,N_4934,N_3744);
or U6822 (N_6822,N_4460,N_3923);
or U6823 (N_6823,N_5155,N_4337);
nor U6824 (N_6824,N_4092,N_3881);
and U6825 (N_6825,N_3662,N_5640);
nand U6826 (N_6826,N_3462,N_4070);
nor U6827 (N_6827,N_4825,N_3469);
and U6828 (N_6828,N_4780,N_4208);
nand U6829 (N_6829,N_4556,N_5164);
nand U6830 (N_6830,N_4665,N_3701);
or U6831 (N_6831,N_3171,N_5245);
or U6832 (N_6832,N_3578,N_5430);
nand U6833 (N_6833,N_5758,N_3309);
nor U6834 (N_6834,N_5938,N_3303);
nor U6835 (N_6835,N_4936,N_4352);
nand U6836 (N_6836,N_5041,N_4589);
nor U6837 (N_6837,N_5919,N_4989);
nand U6838 (N_6838,N_5432,N_4988);
or U6839 (N_6839,N_3316,N_4225);
or U6840 (N_6840,N_4541,N_3186);
nand U6841 (N_6841,N_5620,N_5281);
nor U6842 (N_6842,N_3512,N_3741);
nand U6843 (N_6843,N_4645,N_3145);
xnor U6844 (N_6844,N_4521,N_5415);
nand U6845 (N_6845,N_3784,N_3764);
and U6846 (N_6846,N_3532,N_3519);
nor U6847 (N_6847,N_4760,N_4464);
and U6848 (N_6848,N_4782,N_4457);
nand U6849 (N_6849,N_3508,N_5965);
and U6850 (N_6850,N_5394,N_3173);
or U6851 (N_6851,N_5589,N_5771);
and U6852 (N_6852,N_3007,N_3053);
or U6853 (N_6853,N_4818,N_5237);
or U6854 (N_6854,N_3806,N_4537);
or U6855 (N_6855,N_4214,N_4609);
nand U6856 (N_6856,N_3296,N_5211);
nand U6857 (N_6857,N_4203,N_4234);
nor U6858 (N_6858,N_5250,N_4843);
or U6859 (N_6859,N_4540,N_5808);
nor U6860 (N_6860,N_4376,N_3713);
or U6861 (N_6861,N_4809,N_5446);
nor U6862 (N_6862,N_4223,N_5159);
nor U6863 (N_6863,N_5848,N_5598);
nor U6864 (N_6864,N_3061,N_4859);
nand U6865 (N_6865,N_4019,N_5915);
nor U6866 (N_6866,N_4130,N_4389);
nand U6867 (N_6867,N_3964,N_4650);
and U6868 (N_6868,N_4533,N_3722);
nand U6869 (N_6869,N_3051,N_3111);
nor U6870 (N_6870,N_5817,N_4209);
nor U6871 (N_6871,N_4999,N_5140);
nor U6872 (N_6872,N_3043,N_4310);
and U6873 (N_6873,N_3172,N_4662);
nand U6874 (N_6874,N_3107,N_3223);
nand U6875 (N_6875,N_3787,N_5267);
nor U6876 (N_6876,N_3290,N_3909);
xnor U6877 (N_6877,N_4308,N_3461);
and U6878 (N_6878,N_3491,N_5980);
nor U6879 (N_6879,N_5400,N_5975);
nor U6880 (N_6880,N_4841,N_4766);
and U6881 (N_6881,N_3201,N_3833);
or U6882 (N_6882,N_4775,N_3014);
and U6883 (N_6883,N_3686,N_5679);
and U6884 (N_6884,N_3367,N_5162);
nand U6885 (N_6885,N_5013,N_3432);
and U6886 (N_6886,N_5179,N_4241);
nand U6887 (N_6887,N_4937,N_3627);
and U6888 (N_6888,N_3748,N_5933);
nor U6889 (N_6889,N_4115,N_3129);
or U6890 (N_6890,N_5492,N_3704);
nand U6891 (N_6891,N_4075,N_5970);
xnor U6892 (N_6892,N_5723,N_4206);
or U6893 (N_6893,N_4555,N_4057);
or U6894 (N_6894,N_4730,N_5445);
or U6895 (N_6895,N_3409,N_3616);
nor U6896 (N_6896,N_4648,N_4002);
xor U6897 (N_6897,N_5738,N_5214);
or U6898 (N_6898,N_4855,N_4312);
and U6899 (N_6899,N_3308,N_5969);
nor U6900 (N_6900,N_5493,N_5888);
or U6901 (N_6901,N_3936,N_5768);
nor U6902 (N_6902,N_3487,N_3259);
and U6903 (N_6903,N_3374,N_5839);
or U6904 (N_6904,N_4280,N_5896);
nor U6905 (N_6905,N_5763,N_4865);
nand U6906 (N_6906,N_5355,N_4216);
nand U6907 (N_6907,N_5289,N_5978);
nand U6908 (N_6908,N_4882,N_4788);
or U6909 (N_6909,N_5751,N_3477);
nor U6910 (N_6910,N_4771,N_5597);
nand U6911 (N_6911,N_3705,N_4478);
nor U6912 (N_6912,N_3282,N_5854);
nor U6913 (N_6913,N_3687,N_5031);
nand U6914 (N_6914,N_4947,N_3667);
or U6915 (N_6915,N_4729,N_5579);
nor U6916 (N_6916,N_3551,N_3137);
nor U6917 (N_6917,N_4114,N_5032);
nand U6918 (N_6918,N_5601,N_5376);
and U6919 (N_6919,N_4183,N_5951);
or U6920 (N_6920,N_5117,N_4298);
nor U6921 (N_6921,N_3911,N_5028);
and U6922 (N_6922,N_3879,N_3294);
nand U6923 (N_6923,N_4785,N_4313);
and U6924 (N_6924,N_4406,N_5968);
and U6925 (N_6925,N_3274,N_5122);
nor U6926 (N_6926,N_4765,N_5587);
or U6927 (N_6927,N_5039,N_3095);
nand U6928 (N_6928,N_4581,N_4432);
nor U6929 (N_6929,N_4876,N_4064);
and U6930 (N_6930,N_5247,N_4499);
nand U6931 (N_6931,N_4287,N_5776);
nand U6932 (N_6932,N_4087,N_5123);
and U6933 (N_6933,N_5722,N_5105);
or U6934 (N_6934,N_4303,N_4747);
nand U6935 (N_6935,N_5466,N_3228);
nor U6936 (N_6936,N_3234,N_5845);
and U6937 (N_6937,N_4750,N_5556);
xnor U6938 (N_6938,N_4703,N_3405);
nand U6939 (N_6939,N_5813,N_4958);
nor U6940 (N_6940,N_3782,N_3576);
and U6941 (N_6941,N_4905,N_4548);
or U6942 (N_6942,N_4590,N_4552);
xor U6943 (N_6943,N_5789,N_3779);
nand U6944 (N_6944,N_4523,N_5703);
nand U6945 (N_6945,N_5153,N_4233);
or U6946 (N_6946,N_3520,N_4560);
nor U6947 (N_6947,N_3069,N_5539);
and U6948 (N_6948,N_4366,N_5806);
or U6949 (N_6949,N_3387,N_4354);
nand U6950 (N_6950,N_3670,N_5981);
or U6951 (N_6951,N_3361,N_5901);
and U6952 (N_6952,N_3657,N_5784);
nor U6953 (N_6953,N_5460,N_3985);
and U6954 (N_6954,N_5744,N_4279);
nor U6955 (N_6955,N_3855,N_5440);
and U6956 (N_6956,N_5169,N_4098);
and U6957 (N_6957,N_3808,N_5438);
nand U6958 (N_6958,N_3239,N_4080);
and U6959 (N_6959,N_5321,N_4496);
nor U6960 (N_6960,N_3505,N_5574);
nand U6961 (N_6961,N_3653,N_5221);
and U6962 (N_6962,N_3735,N_3843);
nand U6963 (N_6963,N_5599,N_5992);
or U6964 (N_6964,N_5941,N_4418);
nand U6965 (N_6965,N_4110,N_4235);
nand U6966 (N_6966,N_3526,N_5842);
and U6967 (N_6967,N_5843,N_4912);
nand U6968 (N_6968,N_3452,N_5142);
nand U6969 (N_6969,N_3812,N_5132);
and U6970 (N_6970,N_3028,N_5145);
and U6971 (N_6971,N_3651,N_4161);
or U6972 (N_6972,N_3527,N_5804);
or U6973 (N_6973,N_5973,N_4215);
nand U6974 (N_6974,N_3678,N_4101);
or U6975 (N_6975,N_5897,N_5347);
and U6976 (N_6976,N_4769,N_3193);
and U6977 (N_6977,N_3780,N_4466);
and U6978 (N_6978,N_4451,N_5704);
or U6979 (N_6979,N_3793,N_4356);
and U6980 (N_6980,N_5212,N_5243);
or U6981 (N_6981,N_5558,N_4173);
or U6982 (N_6982,N_5036,N_5905);
nor U6983 (N_6983,N_4044,N_3266);
nand U6984 (N_6984,N_5635,N_5393);
or U6985 (N_6985,N_3823,N_3369);
nand U6986 (N_6986,N_5936,N_3096);
and U6987 (N_6987,N_5803,N_4412);
nor U6988 (N_6988,N_5072,N_3492);
or U6989 (N_6989,N_5844,N_5091);
or U6990 (N_6990,N_4580,N_3338);
nor U6991 (N_6991,N_4062,N_4712);
and U6992 (N_6992,N_4009,N_4094);
nor U6993 (N_6993,N_3248,N_3440);
nor U6994 (N_6994,N_5235,N_4005);
or U6995 (N_6995,N_4332,N_4029);
and U6996 (N_6996,N_5254,N_5144);
or U6997 (N_6997,N_4923,N_5242);
or U6998 (N_6998,N_3599,N_4306);
and U6999 (N_6999,N_4165,N_3048);
and U7000 (N_7000,N_4404,N_3720);
nand U7001 (N_7001,N_4726,N_5815);
or U7002 (N_7002,N_4606,N_3862);
or U7003 (N_7003,N_5368,N_5345);
or U7004 (N_7004,N_4391,N_5359);
and U7005 (N_7005,N_5025,N_4646);
nand U7006 (N_7006,N_3045,N_4535);
and U7007 (N_7007,N_4323,N_5141);
nand U7008 (N_7008,N_3307,N_5948);
nand U7009 (N_7009,N_3360,N_5076);
nand U7010 (N_7010,N_4024,N_3907);
and U7011 (N_7011,N_4210,N_5358);
nand U7012 (N_7012,N_4693,N_5974);
nor U7013 (N_7013,N_3419,N_5296);
nand U7014 (N_7014,N_3185,N_4189);
nor U7015 (N_7015,N_3474,N_5867);
nor U7016 (N_7016,N_4487,N_3399);
or U7017 (N_7017,N_3652,N_3292);
and U7018 (N_7018,N_3966,N_3814);
nand U7019 (N_7019,N_5026,N_4734);
or U7020 (N_7020,N_4720,N_4875);
and U7021 (N_7021,N_3151,N_4267);
and U7022 (N_7022,N_3961,N_5524);
nand U7023 (N_7023,N_3629,N_4238);
nand U7024 (N_7024,N_4550,N_4906);
nor U7025 (N_7025,N_4292,N_5692);
nand U7026 (N_7026,N_5305,N_4924);
or U7027 (N_7027,N_3603,N_5308);
nand U7028 (N_7028,N_3871,N_3035);
or U7029 (N_7029,N_5442,N_3213);
and U7030 (N_7030,N_5248,N_3497);
nand U7031 (N_7031,N_4899,N_4072);
and U7032 (N_7032,N_3198,N_3905);
nand U7033 (N_7033,N_5086,N_5536);
nor U7034 (N_7034,N_4102,N_4228);
nand U7035 (N_7035,N_5622,N_4781);
nand U7036 (N_7036,N_3799,N_5707);
or U7037 (N_7037,N_5756,N_3445);
or U7038 (N_7038,N_4724,N_3774);
or U7039 (N_7039,N_4739,N_4570);
nand U7040 (N_7040,N_4171,N_3541);
nor U7041 (N_7041,N_3800,N_5055);
nand U7042 (N_7042,N_4122,N_3267);
nand U7043 (N_7043,N_4469,N_5080);
and U7044 (N_7044,N_3415,N_4307);
nor U7045 (N_7045,N_4643,N_3542);
or U7046 (N_7046,N_3271,N_3264);
and U7047 (N_7047,N_3500,N_3944);
and U7048 (N_7048,N_4410,N_4946);
nand U7049 (N_7049,N_3240,N_5729);
nand U7050 (N_7050,N_5398,N_4455);
or U7051 (N_7051,N_5935,N_3070);
and U7052 (N_7052,N_5939,N_3438);
and U7053 (N_7053,N_4676,N_5310);
or U7054 (N_7054,N_5027,N_5322);
nand U7055 (N_7055,N_3003,N_5233);
nor U7056 (N_7056,N_5877,N_3436);
nor U7057 (N_7057,N_4839,N_5925);
nand U7058 (N_7058,N_4618,N_3417);
or U7059 (N_7059,N_3673,N_4284);
nand U7060 (N_7060,N_5382,N_5304);
xor U7061 (N_7061,N_3431,N_3912);
nand U7062 (N_7062,N_4755,N_5731);
and U7063 (N_7063,N_4604,N_5564);
nor U7064 (N_7064,N_3060,N_4732);
nand U7065 (N_7065,N_3801,N_3123);
and U7066 (N_7066,N_5188,N_5531);
nand U7067 (N_7067,N_3165,N_4617);
nor U7068 (N_7068,N_3942,N_5439);
nor U7069 (N_7069,N_5647,N_4078);
nor U7070 (N_7070,N_4419,N_3202);
or U7071 (N_7071,N_3995,N_3920);
or U7072 (N_7072,N_4329,N_3403);
and U7073 (N_7073,N_5569,N_3797);
nor U7074 (N_7074,N_3125,N_4943);
nor U7075 (N_7075,N_3375,N_5067);
xor U7076 (N_7076,N_5633,N_4526);
nor U7077 (N_7077,N_5082,N_3938);
nor U7078 (N_7078,N_5427,N_4170);
or U7079 (N_7079,N_3215,N_4710);
and U7080 (N_7080,N_3736,N_3197);
nand U7081 (N_7081,N_5339,N_3082);
nand U7082 (N_7082,N_5747,N_5180);
or U7083 (N_7083,N_5174,N_5126);
and U7084 (N_7084,N_3081,N_4289);
or U7085 (N_7085,N_3831,N_5047);
nor U7086 (N_7086,N_3635,N_5658);
nand U7087 (N_7087,N_3809,N_3336);
and U7088 (N_7088,N_4895,N_5861);
or U7089 (N_7089,N_5125,N_3617);
and U7090 (N_7090,N_5085,N_4461);
nand U7091 (N_7091,N_5436,N_3330);
nand U7092 (N_7092,N_3540,N_5899);
or U7093 (N_7093,N_3647,N_5762);
nor U7094 (N_7094,N_4159,N_3446);
or U7095 (N_7095,N_3931,N_4762);
or U7096 (N_7096,N_5388,N_5196);
nand U7097 (N_7097,N_3434,N_5693);
or U7098 (N_7098,N_3067,N_4637);
nor U7099 (N_7099,N_5534,N_3712);
and U7100 (N_7100,N_4706,N_4515);
and U7101 (N_7101,N_3088,N_4187);
nor U7102 (N_7102,N_5830,N_3464);
or U7103 (N_7103,N_5097,N_3114);
nand U7104 (N_7104,N_4630,N_4994);
nor U7105 (N_7105,N_4247,N_3852);
nand U7106 (N_7106,N_3301,N_4028);
nand U7107 (N_7107,N_5202,N_5932);
or U7108 (N_7108,N_3363,N_4060);
or U7109 (N_7109,N_5752,N_4063);
and U7110 (N_7110,N_3019,N_5568);
nand U7111 (N_7111,N_4001,N_4504);
nor U7112 (N_7112,N_5494,N_5001);
nand U7113 (N_7113,N_3769,N_5674);
or U7114 (N_7114,N_3725,N_5274);
nand U7115 (N_7115,N_5380,N_5727);
and U7116 (N_7116,N_4425,N_3837);
nand U7117 (N_7117,N_4341,N_3950);
xnor U7118 (N_7118,N_4791,N_3411);
nand U7119 (N_7119,N_4607,N_3661);
and U7120 (N_7120,N_3848,N_3696);
nor U7121 (N_7121,N_5136,N_4714);
nor U7122 (N_7122,N_4500,N_4708);
and U7123 (N_7123,N_5733,N_4192);
nand U7124 (N_7124,N_3273,N_3552);
or U7125 (N_7125,N_4632,N_5391);
and U7126 (N_7126,N_5657,N_3160);
and U7127 (N_7127,N_5423,N_3642);
and U7128 (N_7128,N_4136,N_3559);
or U7129 (N_7129,N_4633,N_4952);
nand U7130 (N_7130,N_3087,N_5306);
xor U7131 (N_7131,N_5645,N_5152);
nor U7132 (N_7132,N_5182,N_5608);
and U7133 (N_7133,N_5644,N_3622);
nor U7134 (N_7134,N_3416,N_4942);
nor U7135 (N_7135,N_3524,N_4344);
nand U7136 (N_7136,N_3217,N_4972);
xor U7137 (N_7137,N_4222,N_4861);
nand U7138 (N_7138,N_5765,N_3152);
or U7139 (N_7139,N_5615,N_4976);
and U7140 (N_7140,N_5957,N_5820);
nand U7141 (N_7141,N_3404,N_3261);
nand U7142 (N_7142,N_5437,N_4291);
or U7143 (N_7143,N_5113,N_3717);
or U7144 (N_7144,N_5920,N_4653);
nor U7145 (N_7145,N_4246,N_4103);
nor U7146 (N_7146,N_3386,N_4143);
nor U7147 (N_7147,N_5463,N_3863);
nand U7148 (N_7148,N_5686,N_4251);
or U7149 (N_7149,N_3719,N_5417);
nand U7150 (N_7150,N_3903,N_4509);
or U7151 (N_7151,N_3639,N_3236);
and U7152 (N_7152,N_3606,N_3400);
nor U7153 (N_7153,N_5517,N_3783);
or U7154 (N_7154,N_5942,N_3645);
and U7155 (N_7155,N_5489,N_5285);
nor U7156 (N_7156,N_5511,N_3106);
nor U7157 (N_7157,N_4796,N_4518);
or U7158 (N_7158,N_3174,N_5718);
nor U7159 (N_7159,N_5163,N_4921);
and U7160 (N_7160,N_4045,N_4834);
nor U7161 (N_7161,N_5023,N_4407);
nand U7162 (N_7162,N_5335,N_3794);
nor U7163 (N_7163,N_4390,N_3056);
and U7164 (N_7164,N_5594,N_3318);
nand U7165 (N_7165,N_3805,N_4677);
nand U7166 (N_7166,N_3253,N_3745);
nor U7167 (N_7167,N_5087,N_5617);
nor U7168 (N_7168,N_3493,N_4944);
nor U7169 (N_7169,N_3846,N_4842);
nor U7170 (N_7170,N_4926,N_5367);
nor U7171 (N_7171,N_5895,N_5476);
and U7172 (N_7172,N_3142,N_3091);
or U7173 (N_7173,N_4324,N_5314);
or U7174 (N_7174,N_3332,N_3041);
or U7175 (N_7175,N_5851,N_5746);
and U7176 (N_7176,N_4034,N_3346);
nand U7177 (N_7177,N_3199,N_4873);
and U7178 (N_7178,N_5307,N_4403);
nor U7179 (N_7179,N_3575,N_3044);
nor U7180 (N_7180,N_5614,N_5343);
nor U7181 (N_7181,N_4015,N_5705);
and U7182 (N_7182,N_4030,N_4685);
or U7183 (N_7183,N_3025,N_5757);
or U7184 (N_7184,N_5592,N_3470);
xnor U7185 (N_7185,N_5167,N_3873);
or U7186 (N_7186,N_3362,N_3317);
nor U7187 (N_7187,N_3382,N_5634);
nand U7188 (N_7188,N_3932,N_3189);
or U7189 (N_7189,N_3543,N_4484);
nor U7190 (N_7190,N_3946,N_5228);
nand U7191 (N_7191,N_5474,N_3064);
nand U7192 (N_7192,N_4033,N_4326);
nand U7193 (N_7193,N_4007,N_4826);
xor U7194 (N_7194,N_5194,N_3489);
and U7195 (N_7195,N_4871,N_4343);
or U7196 (N_7196,N_5301,N_5299);
and U7197 (N_7197,N_3528,N_3293);
nand U7198 (N_7198,N_3538,N_5172);
xnor U7199 (N_7199,N_3904,N_5648);
and U7200 (N_7200,N_5294,N_5945);
and U7201 (N_7201,N_3075,N_4737);
and U7202 (N_7202,N_5348,N_4398);
nor U7203 (N_7203,N_4613,N_4538);
nor U7204 (N_7204,N_4430,N_5277);
nor U7205 (N_7205,N_3585,N_5567);
nor U7206 (N_7206,N_4866,N_4578);
or U7207 (N_7207,N_3429,N_5913);
nor U7208 (N_7208,N_4885,N_5522);
or U7209 (N_7209,N_3531,N_3166);
xnor U7210 (N_7210,N_5502,N_3302);
or U7211 (N_7211,N_5282,N_3726);
nor U7212 (N_7212,N_3668,N_5682);
or U7213 (N_7213,N_3851,N_3393);
nand U7214 (N_7214,N_5448,N_3055);
nand U7215 (N_7215,N_4864,N_4772);
nor U7216 (N_7216,N_5297,N_5947);
or U7217 (N_7217,N_4661,N_4274);
nand U7218 (N_7218,N_5168,N_3495);
nand U7219 (N_7219,N_4503,N_4634);
and U7220 (N_7220,N_5390,N_5961);
or U7221 (N_7221,N_5755,N_3479);
or U7222 (N_7222,N_4061,N_3329);
or U7223 (N_7223,N_5373,N_4179);
nand U7224 (N_7224,N_3688,N_4508);
and U7225 (N_7225,N_3170,N_5963);
or U7226 (N_7226,N_4283,N_5106);
nand U7227 (N_7227,N_5231,N_3394);
nand U7228 (N_7228,N_3755,N_5660);
and U7229 (N_7229,N_3016,N_4881);
nand U7230 (N_7230,N_5778,N_5497);
xor U7231 (N_7231,N_4516,N_4423);
or U7232 (N_7232,N_4738,N_5452);
nor U7233 (N_7233,N_5639,N_3113);
nand U7234 (N_7234,N_5790,N_3596);
nor U7235 (N_7235,N_5050,N_5496);
and U7236 (N_7236,N_4945,N_3204);
or U7237 (N_7237,N_4651,N_5429);
and U7238 (N_7238,N_5575,N_3295);
nand U7239 (N_7239,N_3331,N_3357);
and U7240 (N_7240,N_5728,N_4836);
and U7241 (N_7241,N_4084,N_4954);
xor U7242 (N_7242,N_4275,N_5792);
nor U7243 (N_7243,N_4990,N_3257);
nand U7244 (N_7244,N_4733,N_3372);
and U7245 (N_7245,N_4182,N_3268);
nand U7246 (N_7246,N_4128,N_4690);
and U7247 (N_7247,N_5468,N_3890);
and U7248 (N_7248,N_4272,N_3353);
or U7249 (N_7249,N_4276,N_5286);
and U7250 (N_7250,N_3397,N_3502);
nor U7251 (N_7251,N_5170,N_4981);
and U7252 (N_7252,N_4393,N_3435);
nor U7253 (N_7253,N_5609,N_3155);
and U7254 (N_7254,N_4869,N_5561);
and U7255 (N_7255,N_3693,N_5381);
nor U7256 (N_7256,N_5356,N_4983);
nand U7257 (N_7257,N_5477,N_5349);
xor U7258 (N_7258,N_3385,N_3421);
xor U7259 (N_7259,N_3929,N_4468);
or U7260 (N_7260,N_5241,N_3227);
nand U7261 (N_7261,N_4817,N_3232);
and U7262 (N_7262,N_5462,N_4657);
and U7263 (N_7263,N_4145,N_5528);
nor U7264 (N_7264,N_5971,N_3355);
or U7265 (N_7265,N_5022,N_5872);
nor U7266 (N_7266,N_5057,N_4916);
and U7267 (N_7267,N_3898,N_3350);
and U7268 (N_7268,N_3214,N_5191);
or U7269 (N_7269,N_5059,N_4654);
nand U7270 (N_7270,N_5859,N_3743);
nand U7271 (N_7271,N_5018,N_5994);
nor U7272 (N_7272,N_4364,N_5507);
nand U7273 (N_7273,N_4069,N_5198);
or U7274 (N_7274,N_5490,N_4847);
nand U7275 (N_7275,N_3507,N_5158);
nand U7276 (N_7276,N_4577,N_4625);
nor U7277 (N_7277,N_4574,N_4017);
and U7278 (N_7278,N_4950,N_5508);
nand U7279 (N_7279,N_5698,N_5993);
nand U7280 (N_7280,N_4088,N_3690);
nor U7281 (N_7281,N_3761,N_3643);
nor U7282 (N_7282,N_3218,N_3313);
nor U7283 (N_7283,N_3644,N_4565);
or U7284 (N_7284,N_3439,N_3850);
nor U7285 (N_7285,N_5628,N_4984);
nor U7286 (N_7286,N_4863,N_3758);
nand U7287 (N_7287,N_3568,N_4479);
or U7288 (N_7288,N_3015,N_3790);
and U7289 (N_7289,N_4282,N_4701);
nand U7290 (N_7290,N_3504,N_5518);
and U7291 (N_7291,N_3728,N_4922);
nand U7292 (N_7292,N_3548,N_3841);
or U7293 (N_7293,N_4615,N_4226);
nand U7294 (N_7294,N_5976,N_5853);
nor U7295 (N_7295,N_4149,N_4794);
and U7296 (N_7296,N_4758,N_4514);
nor U7297 (N_7297,N_4480,N_3373);
nand U7298 (N_7298,N_4415,N_4056);
and U7299 (N_7299,N_4995,N_4893);
xor U7300 (N_7300,N_5051,N_3770);
and U7301 (N_7301,N_5002,N_4382);
or U7302 (N_7302,N_4277,N_3192);
or U7303 (N_7303,N_5730,N_4328);
nor U7304 (N_7304,N_4131,N_4640);
and U7305 (N_7305,N_5912,N_3150);
nand U7306 (N_7306,N_4361,N_3365);
or U7307 (N_7307,N_3499,N_5444);
nor U7308 (N_7308,N_3636,N_4339);
nand U7309 (N_7309,N_3572,N_3059);
or U7310 (N_7310,N_4777,N_3947);
and U7311 (N_7311,N_5006,N_4296);
and U7312 (N_7312,N_5449,N_5495);
or U7313 (N_7313,N_5350,N_4262);
and U7314 (N_7314,N_3233,N_5239);
and U7315 (N_7315,N_5366,N_3473);
and U7316 (N_7316,N_3977,N_5549);
nand U7317 (N_7317,N_3659,N_3398);
nor U7318 (N_7318,N_4380,N_4434);
nor U7319 (N_7319,N_4579,N_4935);
nor U7320 (N_7320,N_4153,N_3324);
or U7321 (N_7321,N_3756,N_4405);
nand U7322 (N_7322,N_3138,N_5336);
nor U7323 (N_7323,N_3437,N_3004);
nor U7324 (N_7324,N_3988,N_3834);
and U7325 (N_7325,N_5249,N_4844);
nor U7326 (N_7326,N_4239,N_5557);
or U7327 (N_7327,N_5207,N_4642);
xnor U7328 (N_7328,N_4032,N_4293);
or U7329 (N_7329,N_5520,N_5667);
nor U7330 (N_7330,N_4351,N_5995);
or U7331 (N_7331,N_3211,N_3207);
nor U7332 (N_7332,N_4501,N_4180);
xnor U7333 (N_7333,N_4139,N_4928);
nor U7334 (N_7334,N_3928,N_4635);
nand U7335 (N_7335,N_5046,N_3256);
or U7336 (N_7336,N_4784,N_3723);
nand U7337 (N_7337,N_3822,N_5303);
and U7338 (N_7338,N_4745,N_4621);
and U7339 (N_7339,N_3116,N_5605);
nand U7340 (N_7340,N_3333,N_5278);
or U7341 (N_7341,N_4666,N_5749);
xor U7342 (N_7342,N_4868,N_3281);
nor U7343 (N_7343,N_3063,N_4506);
nand U7344 (N_7344,N_4831,N_3824);
and U7345 (N_7345,N_5005,N_3771);
or U7346 (N_7346,N_5825,N_4219);
nor U7347 (N_7347,N_3791,N_5183);
nand U7348 (N_7348,N_4317,N_3529);
or U7349 (N_7349,N_4321,N_5696);
nand U7350 (N_7350,N_5453,N_4820);
nand U7351 (N_7351,N_4371,N_4381);
nor U7352 (N_7352,N_4175,N_5330);
and U7353 (N_7353,N_3734,N_5716);
and U7354 (N_7354,N_3339,N_5966);
nor U7355 (N_7355,N_5959,N_4384);
and U7356 (N_7356,N_5642,N_3289);
and U7357 (N_7357,N_5471,N_3702);
nor U7358 (N_7358,N_4442,N_4585);
or U7359 (N_7359,N_5217,N_3731);
nor U7360 (N_7360,N_3126,N_4704);
or U7361 (N_7361,N_3132,N_3122);
or U7362 (N_7362,N_3742,N_5377);
nor U7363 (N_7363,N_3444,N_5671);
nor U7364 (N_7364,N_5669,N_4202);
and U7365 (N_7365,N_3094,N_5835);
nand U7366 (N_7366,N_5739,N_4918);
nor U7367 (N_7367,N_4551,N_5787);
nor U7368 (N_7368,N_4446,N_3343);
or U7369 (N_7369,N_3072,N_3975);
or U7370 (N_7370,N_5069,N_4919);
or U7371 (N_7371,N_3714,N_4884);
or U7372 (N_7372,N_4649,N_4191);
or U7373 (N_7373,N_4563,N_5357);
nor U7374 (N_7374,N_3483,N_5223);
nor U7375 (N_7375,N_3046,N_4723);
nand U7376 (N_7376,N_3359,N_3131);
or U7377 (N_7377,N_3715,N_3050);
or U7378 (N_7378,N_4322,N_3241);
or U7379 (N_7379,N_3974,N_5735);
and U7380 (N_7380,N_3803,N_5078);
nor U7381 (N_7381,N_5488,N_3632);
and U7382 (N_7382,N_3314,N_5953);
xor U7383 (N_7383,N_4286,N_3057);
and U7384 (N_7384,N_3337,N_3086);
nor U7385 (N_7385,N_4174,N_5666);
or U7386 (N_7386,N_5007,N_5205);
nand U7387 (N_7387,N_5581,N_4963);
xnor U7388 (N_7388,N_5720,N_4169);
nor U7389 (N_7389,N_5213,N_4993);
and U7390 (N_7390,N_3017,N_3953);
nand U7391 (N_7391,N_3935,N_5181);
nor U7392 (N_7392,N_3886,N_5115);
xor U7393 (N_7393,N_5512,N_3878);
or U7394 (N_7394,N_4569,N_3916);
xnor U7395 (N_7395,N_4401,N_4067);
nor U7396 (N_7396,N_3457,N_3978);
nor U7397 (N_7397,N_5095,N_3865);
or U7398 (N_7398,N_5220,N_4107);
nor U7399 (N_7399,N_5457,N_3424);
xnor U7400 (N_7400,N_4204,N_5482);
nand U7401 (N_7401,N_4256,N_4736);
or U7402 (N_7402,N_3200,N_3766);
nand U7403 (N_7403,N_4052,N_3305);
and U7404 (N_7404,N_5090,N_3413);
or U7405 (N_7405,N_3640,N_4808);
and U7406 (N_7406,N_3826,N_4154);
or U7407 (N_7407,N_3471,N_5795);
nand U7408 (N_7408,N_4374,N_4333);
nand U7409 (N_7409,N_3754,N_3641);
or U7410 (N_7410,N_3656,N_5821);
nand U7411 (N_7411,N_4476,N_5258);
nand U7412 (N_7412,N_4848,N_3880);
and U7413 (N_7413,N_5510,N_3711);
or U7414 (N_7414,N_4878,N_4870);
or U7415 (N_7415,N_4124,N_3591);
nor U7416 (N_7416,N_4660,N_4776);
or U7417 (N_7417,N_4185,N_4392);
or U7418 (N_7418,N_5325,N_4010);
nand U7419 (N_7419,N_5869,N_4109);
or U7420 (N_7420,N_5760,N_5868);
and U7421 (N_7421,N_5619,N_4163);
or U7422 (N_7422,N_3612,N_3889);
nor U7423 (N_7423,N_3547,N_3503);
and U7424 (N_7424,N_5190,N_3875);
nor U7425 (N_7425,N_4395,N_5389);
and U7426 (N_7426,N_5331,N_4470);
nor U7427 (N_7427,N_5010,N_3858);
xor U7428 (N_7428,N_3184,N_3840);
nand U7429 (N_7429,N_3810,N_4085);
nand U7430 (N_7430,N_4325,N_4799);
or U7431 (N_7431,N_3973,N_3027);
xor U7432 (N_7432,N_4018,N_3588);
nand U7433 (N_7433,N_4525,N_4804);
nor U7434 (N_7434,N_4536,N_5263);
or U7435 (N_7435,N_4011,N_5261);
or U7436 (N_7436,N_5782,N_3349);
or U7437 (N_7437,N_4059,N_3707);
nand U7438 (N_7438,N_5064,N_5700);
nor U7439 (N_7439,N_4245,N_3939);
nor U7440 (N_7440,N_5098,N_5991);
or U7441 (N_7441,N_3209,N_4431);
nand U7442 (N_7442,N_5585,N_3615);
or U7443 (N_7443,N_4821,N_5379);
nand U7444 (N_7444,N_4707,N_4244);
nand U7445 (N_7445,N_4137,N_3380);
nand U7446 (N_7446,N_3994,N_5215);
nand U7447 (N_7447,N_4527,N_5819);
xnor U7448 (N_7448,N_4417,N_3498);
nor U7449 (N_7449,N_5129,N_4031);
nor U7450 (N_7450,N_3620,N_3986);
and U7451 (N_7451,N_4641,N_3472);
and U7452 (N_7452,N_5092,N_3864);
nor U7453 (N_7453,N_4872,N_4592);
and U7454 (N_7454,N_3183,N_4467);
nor U7455 (N_7455,N_5865,N_5362);
nor U7456 (N_7456,N_5333,N_4941);
nand U7457 (N_7457,N_5240,N_3279);
and U7458 (N_7458,N_5710,N_5960);
nand U7459 (N_7459,N_3983,N_5685);
nand U7460 (N_7460,N_3910,N_5548);
nand U7461 (N_7461,N_5643,N_4849);
nand U7462 (N_7462,N_4658,N_3956);
nor U7463 (N_7463,N_3681,N_3481);
nand U7464 (N_7464,N_5829,N_5726);
and U7465 (N_7465,N_5745,N_3955);
and U7466 (N_7466,N_3700,N_4302);
nand U7467 (N_7467,N_5812,N_3586);
nand U7468 (N_7468,N_5802,N_4813);
nand U7469 (N_7469,N_4121,N_5000);
and U7470 (N_7470,N_5378,N_5701);
nand U7471 (N_7471,N_3237,N_5197);
nor U7472 (N_7472,N_3867,N_5375);
and U7473 (N_7473,N_3634,N_4531);
or U7474 (N_7474,N_4261,N_5012);
nor U7475 (N_7475,N_3877,N_4184);
nand U7476 (N_7476,N_3624,N_4652);
nor U7477 (N_7477,N_3433,N_3195);
and U7478 (N_7478,N_5570,N_3276);
and U7479 (N_7479,N_5588,N_3287);
nand U7480 (N_7480,N_4545,N_3609);
nand U7481 (N_7481,N_4111,N_3550);
nand U7482 (N_7482,N_5447,N_5042);
nand U7483 (N_7483,N_5501,N_4297);
or U7484 (N_7484,N_5206,N_4980);
or U7485 (N_7485,N_3341,N_4042);
and U7486 (N_7486,N_3478,N_3206);
nand U7487 (N_7487,N_4133,N_5563);
and U7488 (N_7488,N_5926,N_3272);
and U7489 (N_7489,N_5799,N_5075);
nor U7490 (N_7490,N_5847,N_3998);
and U7491 (N_7491,N_5849,N_5244);
nand U7492 (N_7492,N_4888,N_3092);
nand U7493 (N_7493,N_4513,N_4845);
or U7494 (N_7494,N_4438,N_3319);
nor U7495 (N_7495,N_5166,N_3937);
nand U7496 (N_7496,N_4142,N_4016);
and U7497 (N_7497,N_5986,N_5708);
and U7498 (N_7498,N_3179,N_4751);
and U7499 (N_7499,N_5210,N_5354);
or U7500 (N_7500,N_4996,N_5166);
nand U7501 (N_7501,N_3474,N_5783);
and U7502 (N_7502,N_3264,N_4276);
nor U7503 (N_7503,N_3529,N_4871);
nor U7504 (N_7504,N_3124,N_3506);
and U7505 (N_7505,N_4368,N_5530);
xor U7506 (N_7506,N_4768,N_5361);
nor U7507 (N_7507,N_4065,N_3070);
and U7508 (N_7508,N_5919,N_5531);
nand U7509 (N_7509,N_5589,N_4532);
and U7510 (N_7510,N_3684,N_3689);
or U7511 (N_7511,N_4476,N_3726);
and U7512 (N_7512,N_3382,N_3035);
xor U7513 (N_7513,N_4379,N_5189);
and U7514 (N_7514,N_3044,N_4721);
nor U7515 (N_7515,N_4386,N_4073);
and U7516 (N_7516,N_5130,N_4957);
or U7517 (N_7517,N_5610,N_3164);
nand U7518 (N_7518,N_3808,N_5655);
nor U7519 (N_7519,N_3961,N_5329);
nand U7520 (N_7520,N_3624,N_4290);
or U7521 (N_7521,N_3938,N_3160);
and U7522 (N_7522,N_5912,N_4565);
nand U7523 (N_7523,N_5475,N_3295);
nand U7524 (N_7524,N_4287,N_4954);
and U7525 (N_7525,N_3412,N_5627);
nand U7526 (N_7526,N_3154,N_3795);
or U7527 (N_7527,N_4750,N_4964);
nor U7528 (N_7528,N_3605,N_5107);
and U7529 (N_7529,N_4216,N_3371);
or U7530 (N_7530,N_4435,N_4512);
or U7531 (N_7531,N_5568,N_3972);
or U7532 (N_7532,N_3101,N_5870);
xor U7533 (N_7533,N_5209,N_3844);
or U7534 (N_7534,N_4798,N_3855);
and U7535 (N_7535,N_4488,N_3237);
nand U7536 (N_7536,N_3598,N_3190);
nor U7537 (N_7537,N_5071,N_3671);
nand U7538 (N_7538,N_3263,N_5865);
nor U7539 (N_7539,N_4301,N_4089);
nor U7540 (N_7540,N_5393,N_5791);
xor U7541 (N_7541,N_5144,N_4386);
nor U7542 (N_7542,N_3052,N_5744);
and U7543 (N_7543,N_3454,N_5887);
nor U7544 (N_7544,N_4891,N_3627);
or U7545 (N_7545,N_4245,N_4200);
or U7546 (N_7546,N_3968,N_4317);
and U7547 (N_7547,N_5480,N_3849);
xnor U7548 (N_7548,N_3654,N_5448);
nand U7549 (N_7549,N_3380,N_5724);
nand U7550 (N_7550,N_4851,N_5647);
nor U7551 (N_7551,N_4094,N_4832);
nor U7552 (N_7552,N_3272,N_5297);
xor U7553 (N_7553,N_3253,N_3357);
and U7554 (N_7554,N_3466,N_4257);
nand U7555 (N_7555,N_5209,N_3302);
or U7556 (N_7556,N_5638,N_4390);
or U7557 (N_7557,N_3444,N_5361);
nand U7558 (N_7558,N_3425,N_3673);
nor U7559 (N_7559,N_3759,N_3550);
and U7560 (N_7560,N_3072,N_5733);
nand U7561 (N_7561,N_4208,N_5814);
nand U7562 (N_7562,N_3989,N_4380);
nand U7563 (N_7563,N_5292,N_5721);
or U7564 (N_7564,N_5190,N_4358);
nand U7565 (N_7565,N_5032,N_4029);
or U7566 (N_7566,N_3394,N_4804);
or U7567 (N_7567,N_4843,N_4622);
and U7568 (N_7568,N_4831,N_5840);
and U7569 (N_7569,N_3224,N_5580);
or U7570 (N_7570,N_4576,N_4639);
and U7571 (N_7571,N_4699,N_4214);
nor U7572 (N_7572,N_3936,N_4972);
nand U7573 (N_7573,N_5452,N_3478);
nor U7574 (N_7574,N_3694,N_5874);
nand U7575 (N_7575,N_4496,N_5799);
nor U7576 (N_7576,N_4300,N_4368);
or U7577 (N_7577,N_3378,N_3384);
nor U7578 (N_7578,N_5864,N_3592);
nand U7579 (N_7579,N_3127,N_3495);
or U7580 (N_7580,N_4675,N_3518);
or U7581 (N_7581,N_5754,N_4364);
nand U7582 (N_7582,N_5697,N_4513);
nand U7583 (N_7583,N_3279,N_5930);
nand U7584 (N_7584,N_4591,N_3123);
or U7585 (N_7585,N_5699,N_5380);
or U7586 (N_7586,N_5459,N_4292);
and U7587 (N_7587,N_3313,N_5201);
nand U7588 (N_7588,N_5245,N_4022);
nand U7589 (N_7589,N_4676,N_3878);
nor U7590 (N_7590,N_4258,N_5086);
nand U7591 (N_7591,N_5397,N_3995);
nor U7592 (N_7592,N_5488,N_3183);
nand U7593 (N_7593,N_3450,N_5599);
nor U7594 (N_7594,N_4905,N_4951);
and U7595 (N_7595,N_5249,N_5555);
nand U7596 (N_7596,N_5535,N_5235);
or U7597 (N_7597,N_4378,N_5754);
nand U7598 (N_7598,N_4313,N_5925);
or U7599 (N_7599,N_4221,N_4570);
or U7600 (N_7600,N_3846,N_5430);
nand U7601 (N_7601,N_3603,N_3867);
nor U7602 (N_7602,N_4360,N_3413);
nor U7603 (N_7603,N_4375,N_5596);
nand U7604 (N_7604,N_3391,N_3455);
or U7605 (N_7605,N_3313,N_3347);
nor U7606 (N_7606,N_5681,N_4120);
xnor U7607 (N_7607,N_4514,N_4566);
xnor U7608 (N_7608,N_5222,N_3201);
nand U7609 (N_7609,N_3275,N_4279);
and U7610 (N_7610,N_3431,N_3778);
nor U7611 (N_7611,N_4006,N_3190);
and U7612 (N_7612,N_4870,N_4807);
xor U7613 (N_7613,N_5750,N_3577);
and U7614 (N_7614,N_4561,N_4380);
or U7615 (N_7615,N_5159,N_4952);
or U7616 (N_7616,N_5555,N_5699);
and U7617 (N_7617,N_5393,N_4216);
nand U7618 (N_7618,N_4038,N_5866);
or U7619 (N_7619,N_4303,N_5223);
nand U7620 (N_7620,N_3525,N_4859);
or U7621 (N_7621,N_3480,N_4758);
xnor U7622 (N_7622,N_3084,N_3500);
or U7623 (N_7623,N_3134,N_5806);
nand U7624 (N_7624,N_3705,N_3087);
nor U7625 (N_7625,N_5542,N_4115);
and U7626 (N_7626,N_3489,N_4578);
nor U7627 (N_7627,N_4892,N_5000);
and U7628 (N_7628,N_3502,N_5085);
xnor U7629 (N_7629,N_4130,N_5076);
nor U7630 (N_7630,N_5743,N_4506);
nor U7631 (N_7631,N_3237,N_5126);
nand U7632 (N_7632,N_4037,N_3827);
and U7633 (N_7633,N_3009,N_5912);
nor U7634 (N_7634,N_3291,N_3729);
nor U7635 (N_7635,N_4985,N_4928);
or U7636 (N_7636,N_3016,N_4170);
nand U7637 (N_7637,N_5185,N_4590);
nand U7638 (N_7638,N_5931,N_5878);
xor U7639 (N_7639,N_3172,N_5130);
or U7640 (N_7640,N_3640,N_5825);
nand U7641 (N_7641,N_3337,N_3360);
or U7642 (N_7642,N_5464,N_4805);
nor U7643 (N_7643,N_3254,N_5807);
nand U7644 (N_7644,N_3312,N_4140);
and U7645 (N_7645,N_4073,N_3981);
nand U7646 (N_7646,N_3247,N_5641);
or U7647 (N_7647,N_4322,N_4712);
or U7648 (N_7648,N_5380,N_5434);
nand U7649 (N_7649,N_3609,N_4351);
nand U7650 (N_7650,N_4871,N_4903);
or U7651 (N_7651,N_3292,N_5710);
or U7652 (N_7652,N_5838,N_5864);
nand U7653 (N_7653,N_4937,N_5795);
and U7654 (N_7654,N_3909,N_4170);
xor U7655 (N_7655,N_4626,N_4618);
xor U7656 (N_7656,N_5496,N_4805);
nand U7657 (N_7657,N_3179,N_4051);
nand U7658 (N_7658,N_3816,N_4109);
and U7659 (N_7659,N_4368,N_4595);
nor U7660 (N_7660,N_5437,N_5453);
nand U7661 (N_7661,N_4002,N_3785);
nor U7662 (N_7662,N_5593,N_5449);
xor U7663 (N_7663,N_4721,N_5738);
or U7664 (N_7664,N_4332,N_3053);
or U7665 (N_7665,N_3180,N_4323);
nand U7666 (N_7666,N_5259,N_3333);
nand U7667 (N_7667,N_3231,N_3413);
and U7668 (N_7668,N_3305,N_4330);
nor U7669 (N_7669,N_5772,N_3853);
nor U7670 (N_7670,N_4618,N_4902);
nor U7671 (N_7671,N_4365,N_5683);
and U7672 (N_7672,N_4938,N_3284);
nor U7673 (N_7673,N_5784,N_3348);
nor U7674 (N_7674,N_3676,N_3613);
and U7675 (N_7675,N_4176,N_4481);
and U7676 (N_7676,N_4917,N_3728);
or U7677 (N_7677,N_3272,N_3594);
or U7678 (N_7678,N_5905,N_4492);
and U7679 (N_7679,N_4995,N_5659);
nand U7680 (N_7680,N_4814,N_3629);
and U7681 (N_7681,N_5954,N_5443);
or U7682 (N_7682,N_3292,N_5543);
nand U7683 (N_7683,N_4689,N_4207);
nand U7684 (N_7684,N_5111,N_4336);
or U7685 (N_7685,N_5959,N_4049);
nor U7686 (N_7686,N_5334,N_5846);
and U7687 (N_7687,N_5255,N_4369);
and U7688 (N_7688,N_4437,N_4132);
nor U7689 (N_7689,N_4499,N_3040);
nand U7690 (N_7690,N_5984,N_4519);
or U7691 (N_7691,N_5458,N_4693);
nor U7692 (N_7692,N_4195,N_5681);
or U7693 (N_7693,N_3442,N_4743);
nand U7694 (N_7694,N_4194,N_5846);
or U7695 (N_7695,N_4951,N_3970);
nor U7696 (N_7696,N_4724,N_5347);
nand U7697 (N_7697,N_3312,N_3706);
or U7698 (N_7698,N_5920,N_3729);
nor U7699 (N_7699,N_4641,N_5837);
nor U7700 (N_7700,N_3322,N_3566);
or U7701 (N_7701,N_3935,N_5727);
or U7702 (N_7702,N_3396,N_3932);
or U7703 (N_7703,N_5166,N_5505);
or U7704 (N_7704,N_3418,N_5198);
and U7705 (N_7705,N_4691,N_3916);
nand U7706 (N_7706,N_4777,N_5653);
nand U7707 (N_7707,N_4362,N_5283);
nand U7708 (N_7708,N_5919,N_3241);
nor U7709 (N_7709,N_4495,N_5732);
nor U7710 (N_7710,N_3206,N_4578);
and U7711 (N_7711,N_5587,N_4246);
nand U7712 (N_7712,N_5396,N_4462);
nor U7713 (N_7713,N_5508,N_4783);
nor U7714 (N_7714,N_5916,N_5233);
or U7715 (N_7715,N_3260,N_4187);
and U7716 (N_7716,N_5826,N_5017);
or U7717 (N_7717,N_4854,N_4475);
nor U7718 (N_7718,N_4458,N_5414);
nand U7719 (N_7719,N_3990,N_3142);
nor U7720 (N_7720,N_5278,N_3268);
nor U7721 (N_7721,N_5439,N_5850);
and U7722 (N_7722,N_5976,N_5070);
nor U7723 (N_7723,N_4001,N_3436);
or U7724 (N_7724,N_3823,N_5200);
nand U7725 (N_7725,N_4469,N_4344);
and U7726 (N_7726,N_5804,N_3295);
or U7727 (N_7727,N_3832,N_3500);
or U7728 (N_7728,N_4060,N_4932);
nor U7729 (N_7729,N_4324,N_3757);
nor U7730 (N_7730,N_5083,N_4591);
and U7731 (N_7731,N_3705,N_5868);
and U7732 (N_7732,N_4869,N_5768);
nor U7733 (N_7733,N_3680,N_5258);
xor U7734 (N_7734,N_4840,N_3027);
or U7735 (N_7735,N_5830,N_5367);
or U7736 (N_7736,N_4933,N_5402);
nand U7737 (N_7737,N_3485,N_4036);
or U7738 (N_7738,N_5118,N_5200);
nand U7739 (N_7739,N_3480,N_5428);
and U7740 (N_7740,N_3102,N_4167);
xor U7741 (N_7741,N_4732,N_5250);
or U7742 (N_7742,N_3465,N_5843);
nand U7743 (N_7743,N_5065,N_3295);
nand U7744 (N_7744,N_5603,N_3970);
nand U7745 (N_7745,N_5217,N_3608);
and U7746 (N_7746,N_4908,N_4110);
xnor U7747 (N_7747,N_4039,N_3567);
and U7748 (N_7748,N_4659,N_5799);
nand U7749 (N_7749,N_5388,N_4675);
and U7750 (N_7750,N_3596,N_5125);
or U7751 (N_7751,N_5072,N_4571);
nand U7752 (N_7752,N_5114,N_3617);
or U7753 (N_7753,N_4724,N_4039);
nand U7754 (N_7754,N_3090,N_5136);
nand U7755 (N_7755,N_3707,N_5854);
nor U7756 (N_7756,N_4578,N_5370);
and U7757 (N_7757,N_3790,N_4078);
nor U7758 (N_7758,N_5969,N_4798);
and U7759 (N_7759,N_4372,N_3468);
xor U7760 (N_7760,N_4253,N_3372);
nor U7761 (N_7761,N_4172,N_5304);
nand U7762 (N_7762,N_4793,N_4525);
nor U7763 (N_7763,N_4311,N_4964);
nor U7764 (N_7764,N_4330,N_3180);
and U7765 (N_7765,N_3773,N_3853);
and U7766 (N_7766,N_5616,N_3974);
or U7767 (N_7767,N_4051,N_4762);
or U7768 (N_7768,N_4904,N_4881);
nand U7769 (N_7769,N_5957,N_4659);
or U7770 (N_7770,N_3383,N_5074);
nand U7771 (N_7771,N_4554,N_3045);
or U7772 (N_7772,N_5022,N_4934);
or U7773 (N_7773,N_4688,N_4313);
nor U7774 (N_7774,N_5281,N_5546);
and U7775 (N_7775,N_3320,N_3946);
nand U7776 (N_7776,N_4293,N_4646);
nor U7777 (N_7777,N_5029,N_3522);
or U7778 (N_7778,N_3422,N_3838);
nand U7779 (N_7779,N_3034,N_5710);
nand U7780 (N_7780,N_5320,N_5961);
nand U7781 (N_7781,N_3871,N_3419);
nand U7782 (N_7782,N_4768,N_4329);
nand U7783 (N_7783,N_5146,N_3401);
or U7784 (N_7784,N_5090,N_3915);
and U7785 (N_7785,N_4947,N_3389);
nand U7786 (N_7786,N_3585,N_3351);
or U7787 (N_7787,N_5422,N_5602);
nand U7788 (N_7788,N_5801,N_4851);
xor U7789 (N_7789,N_3487,N_4294);
nor U7790 (N_7790,N_3721,N_3942);
nand U7791 (N_7791,N_3859,N_5685);
nand U7792 (N_7792,N_4680,N_5770);
and U7793 (N_7793,N_5193,N_5117);
or U7794 (N_7794,N_4323,N_5491);
nor U7795 (N_7795,N_5071,N_3636);
and U7796 (N_7796,N_3192,N_3563);
nand U7797 (N_7797,N_3254,N_4973);
nor U7798 (N_7798,N_5453,N_4807);
or U7799 (N_7799,N_4934,N_3758);
nand U7800 (N_7800,N_3721,N_4383);
and U7801 (N_7801,N_4284,N_3407);
and U7802 (N_7802,N_3980,N_4049);
nand U7803 (N_7803,N_3989,N_4698);
or U7804 (N_7804,N_4726,N_5291);
nor U7805 (N_7805,N_5417,N_5178);
or U7806 (N_7806,N_5077,N_4334);
nand U7807 (N_7807,N_5446,N_5089);
nor U7808 (N_7808,N_4089,N_3330);
nand U7809 (N_7809,N_4278,N_5149);
nand U7810 (N_7810,N_3460,N_5024);
and U7811 (N_7811,N_4604,N_5458);
nand U7812 (N_7812,N_5918,N_3181);
nand U7813 (N_7813,N_5472,N_4009);
and U7814 (N_7814,N_5180,N_3694);
and U7815 (N_7815,N_5291,N_5969);
nand U7816 (N_7816,N_5049,N_5778);
and U7817 (N_7817,N_4611,N_3719);
nor U7818 (N_7818,N_3949,N_4134);
nor U7819 (N_7819,N_4591,N_5875);
and U7820 (N_7820,N_5857,N_5097);
or U7821 (N_7821,N_3687,N_5118);
nand U7822 (N_7822,N_5177,N_5505);
nand U7823 (N_7823,N_5350,N_5546);
or U7824 (N_7824,N_3949,N_3730);
nand U7825 (N_7825,N_3533,N_4315);
nand U7826 (N_7826,N_4573,N_5193);
xor U7827 (N_7827,N_4528,N_5210);
or U7828 (N_7828,N_4633,N_3470);
nor U7829 (N_7829,N_5919,N_5179);
and U7830 (N_7830,N_3128,N_4730);
or U7831 (N_7831,N_3322,N_5164);
xor U7832 (N_7832,N_3084,N_5346);
nor U7833 (N_7833,N_4962,N_5327);
and U7834 (N_7834,N_4151,N_3429);
nor U7835 (N_7835,N_4234,N_3780);
and U7836 (N_7836,N_3793,N_5967);
or U7837 (N_7837,N_5416,N_4954);
or U7838 (N_7838,N_5578,N_4620);
nor U7839 (N_7839,N_4017,N_3849);
nand U7840 (N_7840,N_3785,N_5807);
xor U7841 (N_7841,N_5814,N_3820);
nand U7842 (N_7842,N_4754,N_5723);
or U7843 (N_7843,N_5217,N_3853);
xor U7844 (N_7844,N_4704,N_3632);
nand U7845 (N_7845,N_5069,N_5357);
nand U7846 (N_7846,N_5982,N_4313);
nand U7847 (N_7847,N_3453,N_5818);
xnor U7848 (N_7848,N_4391,N_3744);
nand U7849 (N_7849,N_5592,N_3954);
and U7850 (N_7850,N_5152,N_5185);
nand U7851 (N_7851,N_4257,N_5965);
and U7852 (N_7852,N_3204,N_4859);
or U7853 (N_7853,N_4893,N_3808);
or U7854 (N_7854,N_5491,N_3839);
and U7855 (N_7855,N_5202,N_3042);
nand U7856 (N_7856,N_5580,N_4276);
nor U7857 (N_7857,N_4722,N_4741);
and U7858 (N_7858,N_3134,N_3480);
nand U7859 (N_7859,N_5338,N_3393);
nand U7860 (N_7860,N_3449,N_3229);
nor U7861 (N_7861,N_4200,N_3578);
nand U7862 (N_7862,N_4785,N_5444);
or U7863 (N_7863,N_5596,N_5350);
or U7864 (N_7864,N_5484,N_5860);
nor U7865 (N_7865,N_4876,N_4419);
nand U7866 (N_7866,N_4135,N_5388);
and U7867 (N_7867,N_4029,N_4883);
or U7868 (N_7868,N_3930,N_3415);
and U7869 (N_7869,N_4821,N_4964);
nor U7870 (N_7870,N_4269,N_4924);
xnor U7871 (N_7871,N_3940,N_4066);
or U7872 (N_7872,N_5456,N_4639);
nand U7873 (N_7873,N_3616,N_5309);
nand U7874 (N_7874,N_4737,N_4740);
nor U7875 (N_7875,N_3293,N_4841);
or U7876 (N_7876,N_3527,N_5225);
and U7877 (N_7877,N_5964,N_5552);
nand U7878 (N_7878,N_3744,N_3221);
nand U7879 (N_7879,N_3415,N_5624);
or U7880 (N_7880,N_4350,N_5457);
nand U7881 (N_7881,N_4198,N_5950);
nand U7882 (N_7882,N_5583,N_4082);
and U7883 (N_7883,N_4086,N_3166);
or U7884 (N_7884,N_4822,N_4392);
nor U7885 (N_7885,N_3009,N_3027);
and U7886 (N_7886,N_5588,N_4644);
and U7887 (N_7887,N_3102,N_5056);
or U7888 (N_7888,N_5330,N_5810);
or U7889 (N_7889,N_4905,N_4674);
or U7890 (N_7890,N_3316,N_3027);
and U7891 (N_7891,N_3830,N_4560);
nand U7892 (N_7892,N_3155,N_3610);
nor U7893 (N_7893,N_4785,N_5939);
and U7894 (N_7894,N_3419,N_3810);
and U7895 (N_7895,N_3036,N_5233);
or U7896 (N_7896,N_3723,N_3986);
or U7897 (N_7897,N_3935,N_5715);
nor U7898 (N_7898,N_3065,N_5810);
nor U7899 (N_7899,N_3759,N_5528);
or U7900 (N_7900,N_3665,N_3817);
xor U7901 (N_7901,N_4113,N_5753);
or U7902 (N_7902,N_5857,N_5460);
nor U7903 (N_7903,N_4293,N_3845);
nand U7904 (N_7904,N_4606,N_3446);
or U7905 (N_7905,N_5647,N_4345);
nor U7906 (N_7906,N_3216,N_5871);
or U7907 (N_7907,N_4071,N_4281);
xnor U7908 (N_7908,N_3294,N_5046);
nor U7909 (N_7909,N_4159,N_4226);
nand U7910 (N_7910,N_3695,N_5143);
or U7911 (N_7911,N_5333,N_3852);
or U7912 (N_7912,N_5207,N_5758);
or U7913 (N_7913,N_5055,N_3230);
nor U7914 (N_7914,N_4412,N_5370);
or U7915 (N_7915,N_5560,N_5584);
nand U7916 (N_7916,N_3412,N_4719);
or U7917 (N_7917,N_5489,N_3715);
or U7918 (N_7918,N_4403,N_3386);
and U7919 (N_7919,N_3979,N_4291);
nand U7920 (N_7920,N_5460,N_5121);
and U7921 (N_7921,N_3724,N_4000);
nor U7922 (N_7922,N_5397,N_5531);
or U7923 (N_7923,N_4277,N_5546);
and U7924 (N_7924,N_4474,N_5242);
or U7925 (N_7925,N_3761,N_5913);
nand U7926 (N_7926,N_5663,N_4063);
nand U7927 (N_7927,N_5869,N_3740);
and U7928 (N_7928,N_3506,N_5252);
or U7929 (N_7929,N_4510,N_5234);
nand U7930 (N_7930,N_4165,N_5065);
and U7931 (N_7931,N_5259,N_5150);
nor U7932 (N_7932,N_5433,N_5665);
nand U7933 (N_7933,N_3502,N_4098);
nand U7934 (N_7934,N_3622,N_5550);
or U7935 (N_7935,N_3334,N_5620);
and U7936 (N_7936,N_4746,N_3988);
nand U7937 (N_7937,N_3023,N_4989);
nand U7938 (N_7938,N_3105,N_3760);
and U7939 (N_7939,N_5870,N_5378);
and U7940 (N_7940,N_5262,N_4449);
or U7941 (N_7941,N_5176,N_5074);
nor U7942 (N_7942,N_3766,N_3325);
and U7943 (N_7943,N_5315,N_5942);
nand U7944 (N_7944,N_5030,N_4921);
nand U7945 (N_7945,N_3406,N_5511);
nand U7946 (N_7946,N_4949,N_3352);
nor U7947 (N_7947,N_3071,N_3823);
nand U7948 (N_7948,N_4041,N_3365);
nor U7949 (N_7949,N_4980,N_4088);
or U7950 (N_7950,N_3990,N_5736);
and U7951 (N_7951,N_5718,N_5900);
or U7952 (N_7952,N_3481,N_4646);
xor U7953 (N_7953,N_3850,N_4867);
nor U7954 (N_7954,N_3989,N_5233);
nor U7955 (N_7955,N_4545,N_3664);
nand U7956 (N_7956,N_3968,N_4145);
nand U7957 (N_7957,N_3789,N_5877);
or U7958 (N_7958,N_3343,N_5024);
or U7959 (N_7959,N_4736,N_5018);
or U7960 (N_7960,N_5516,N_3957);
nand U7961 (N_7961,N_5228,N_5872);
or U7962 (N_7962,N_5126,N_5829);
nor U7963 (N_7963,N_4147,N_5143);
nor U7964 (N_7964,N_5770,N_4060);
xnor U7965 (N_7965,N_3147,N_4389);
and U7966 (N_7966,N_4073,N_4422);
nor U7967 (N_7967,N_3690,N_3928);
nor U7968 (N_7968,N_5604,N_5485);
nand U7969 (N_7969,N_3512,N_4752);
nand U7970 (N_7970,N_4103,N_5986);
nor U7971 (N_7971,N_4223,N_5881);
and U7972 (N_7972,N_3996,N_4299);
nand U7973 (N_7973,N_3955,N_4642);
and U7974 (N_7974,N_3598,N_3379);
and U7975 (N_7975,N_3005,N_4179);
or U7976 (N_7976,N_4595,N_3351);
and U7977 (N_7977,N_5312,N_3969);
nor U7978 (N_7978,N_4022,N_4714);
nor U7979 (N_7979,N_4651,N_5529);
nand U7980 (N_7980,N_5990,N_3968);
nand U7981 (N_7981,N_5751,N_5904);
nor U7982 (N_7982,N_4038,N_4545);
nand U7983 (N_7983,N_4681,N_5904);
nor U7984 (N_7984,N_5795,N_3582);
xor U7985 (N_7985,N_5783,N_5905);
and U7986 (N_7986,N_4882,N_3341);
and U7987 (N_7987,N_5915,N_4251);
and U7988 (N_7988,N_4537,N_5704);
nand U7989 (N_7989,N_4191,N_3935);
and U7990 (N_7990,N_5555,N_4354);
and U7991 (N_7991,N_5054,N_4726);
nor U7992 (N_7992,N_5827,N_4974);
and U7993 (N_7993,N_4609,N_4206);
nor U7994 (N_7994,N_3844,N_4832);
nand U7995 (N_7995,N_4770,N_5151);
or U7996 (N_7996,N_5130,N_5999);
nand U7997 (N_7997,N_3239,N_5813);
and U7998 (N_7998,N_5670,N_5174);
nor U7999 (N_7999,N_4231,N_5856);
or U8000 (N_8000,N_4818,N_4066);
nor U8001 (N_8001,N_4142,N_5471);
nand U8002 (N_8002,N_5589,N_3789);
and U8003 (N_8003,N_3405,N_5814);
nor U8004 (N_8004,N_3605,N_3708);
or U8005 (N_8005,N_3853,N_3389);
or U8006 (N_8006,N_3120,N_5384);
and U8007 (N_8007,N_3005,N_4270);
nand U8008 (N_8008,N_3653,N_3744);
nor U8009 (N_8009,N_4184,N_3605);
xnor U8010 (N_8010,N_5293,N_3570);
nand U8011 (N_8011,N_3906,N_5306);
and U8012 (N_8012,N_3533,N_4129);
and U8013 (N_8013,N_4563,N_4076);
nor U8014 (N_8014,N_4377,N_5601);
and U8015 (N_8015,N_5687,N_3819);
or U8016 (N_8016,N_3204,N_3667);
nand U8017 (N_8017,N_4834,N_5946);
nand U8018 (N_8018,N_5300,N_5040);
or U8019 (N_8019,N_5368,N_3771);
and U8020 (N_8020,N_5866,N_3968);
or U8021 (N_8021,N_4520,N_3000);
nor U8022 (N_8022,N_4403,N_4451);
nand U8023 (N_8023,N_5305,N_4267);
or U8024 (N_8024,N_3042,N_5879);
xnor U8025 (N_8025,N_3836,N_4735);
nor U8026 (N_8026,N_3360,N_5361);
and U8027 (N_8027,N_4259,N_5701);
nand U8028 (N_8028,N_5016,N_5201);
nand U8029 (N_8029,N_3272,N_4694);
and U8030 (N_8030,N_3331,N_4468);
or U8031 (N_8031,N_3699,N_4870);
nand U8032 (N_8032,N_5945,N_4617);
and U8033 (N_8033,N_5802,N_3673);
and U8034 (N_8034,N_4232,N_3404);
nor U8035 (N_8035,N_4343,N_3338);
xor U8036 (N_8036,N_3082,N_4583);
and U8037 (N_8037,N_4856,N_3642);
or U8038 (N_8038,N_5415,N_5954);
and U8039 (N_8039,N_5179,N_4797);
or U8040 (N_8040,N_3002,N_5685);
and U8041 (N_8041,N_4749,N_4721);
and U8042 (N_8042,N_5831,N_3191);
nand U8043 (N_8043,N_4908,N_4953);
and U8044 (N_8044,N_3675,N_3078);
and U8045 (N_8045,N_5757,N_5382);
and U8046 (N_8046,N_5832,N_5627);
or U8047 (N_8047,N_3568,N_3510);
nand U8048 (N_8048,N_4172,N_5613);
and U8049 (N_8049,N_4656,N_4180);
nor U8050 (N_8050,N_4802,N_3637);
and U8051 (N_8051,N_5445,N_4554);
nand U8052 (N_8052,N_5672,N_5138);
or U8053 (N_8053,N_3667,N_4871);
and U8054 (N_8054,N_4489,N_4001);
nand U8055 (N_8055,N_3110,N_3100);
and U8056 (N_8056,N_3227,N_5242);
and U8057 (N_8057,N_4725,N_3047);
and U8058 (N_8058,N_3770,N_3558);
nor U8059 (N_8059,N_3357,N_5769);
nand U8060 (N_8060,N_5516,N_4280);
and U8061 (N_8061,N_3349,N_5907);
nor U8062 (N_8062,N_4359,N_3112);
nand U8063 (N_8063,N_5785,N_3064);
nor U8064 (N_8064,N_4559,N_3092);
nor U8065 (N_8065,N_5692,N_3481);
and U8066 (N_8066,N_3170,N_3668);
nand U8067 (N_8067,N_3232,N_4568);
nand U8068 (N_8068,N_3949,N_4593);
or U8069 (N_8069,N_4480,N_5246);
nand U8070 (N_8070,N_4515,N_3742);
and U8071 (N_8071,N_3070,N_4121);
or U8072 (N_8072,N_4713,N_3668);
and U8073 (N_8073,N_4515,N_4112);
and U8074 (N_8074,N_3740,N_3777);
nor U8075 (N_8075,N_5764,N_5843);
or U8076 (N_8076,N_4008,N_4042);
and U8077 (N_8077,N_3307,N_4950);
nand U8078 (N_8078,N_5284,N_3614);
nand U8079 (N_8079,N_4144,N_5145);
or U8080 (N_8080,N_5269,N_3170);
and U8081 (N_8081,N_4245,N_3818);
nor U8082 (N_8082,N_4309,N_3623);
nand U8083 (N_8083,N_5747,N_4313);
or U8084 (N_8084,N_5640,N_4091);
and U8085 (N_8085,N_5920,N_3508);
or U8086 (N_8086,N_3115,N_5409);
or U8087 (N_8087,N_5109,N_5192);
or U8088 (N_8088,N_3531,N_4984);
or U8089 (N_8089,N_5868,N_4312);
nand U8090 (N_8090,N_4135,N_3735);
and U8091 (N_8091,N_3682,N_3189);
nand U8092 (N_8092,N_4567,N_5867);
nand U8093 (N_8093,N_4561,N_4431);
and U8094 (N_8094,N_4501,N_5824);
nand U8095 (N_8095,N_5780,N_3681);
nand U8096 (N_8096,N_3469,N_5038);
or U8097 (N_8097,N_5449,N_4164);
nor U8098 (N_8098,N_5029,N_4344);
or U8099 (N_8099,N_3050,N_5703);
nor U8100 (N_8100,N_4524,N_3396);
or U8101 (N_8101,N_3685,N_5239);
or U8102 (N_8102,N_4880,N_3888);
nand U8103 (N_8103,N_5339,N_5682);
nand U8104 (N_8104,N_4552,N_4614);
nor U8105 (N_8105,N_4390,N_4554);
and U8106 (N_8106,N_4975,N_4867);
nand U8107 (N_8107,N_5649,N_5705);
and U8108 (N_8108,N_4002,N_4373);
and U8109 (N_8109,N_5694,N_3331);
nand U8110 (N_8110,N_5911,N_4870);
and U8111 (N_8111,N_3428,N_3939);
or U8112 (N_8112,N_4114,N_3656);
and U8113 (N_8113,N_5260,N_3108);
nor U8114 (N_8114,N_4161,N_4752);
or U8115 (N_8115,N_5781,N_5317);
xor U8116 (N_8116,N_4623,N_5156);
nor U8117 (N_8117,N_3383,N_4162);
nor U8118 (N_8118,N_3387,N_4394);
and U8119 (N_8119,N_5012,N_5903);
xor U8120 (N_8120,N_3740,N_3243);
nand U8121 (N_8121,N_4046,N_5363);
and U8122 (N_8122,N_5126,N_5677);
or U8123 (N_8123,N_5619,N_3559);
and U8124 (N_8124,N_4460,N_5598);
and U8125 (N_8125,N_5264,N_5583);
and U8126 (N_8126,N_5262,N_4259);
or U8127 (N_8127,N_3295,N_5296);
nor U8128 (N_8128,N_4449,N_4086);
nor U8129 (N_8129,N_5470,N_5232);
or U8130 (N_8130,N_4710,N_3524);
nor U8131 (N_8131,N_5239,N_4149);
or U8132 (N_8132,N_3721,N_4694);
and U8133 (N_8133,N_5098,N_3120);
and U8134 (N_8134,N_3766,N_3619);
or U8135 (N_8135,N_5301,N_5435);
nand U8136 (N_8136,N_3003,N_5119);
nor U8137 (N_8137,N_5117,N_3482);
nor U8138 (N_8138,N_4587,N_4087);
nor U8139 (N_8139,N_4644,N_5350);
and U8140 (N_8140,N_3977,N_3092);
nand U8141 (N_8141,N_5791,N_3874);
xnor U8142 (N_8142,N_4925,N_5173);
nand U8143 (N_8143,N_4793,N_5066);
and U8144 (N_8144,N_5517,N_5626);
xor U8145 (N_8145,N_5998,N_5900);
nor U8146 (N_8146,N_4112,N_3579);
nand U8147 (N_8147,N_3890,N_5248);
or U8148 (N_8148,N_4338,N_5458);
nand U8149 (N_8149,N_4121,N_4839);
or U8150 (N_8150,N_4779,N_4472);
or U8151 (N_8151,N_3617,N_4666);
nor U8152 (N_8152,N_4651,N_5637);
and U8153 (N_8153,N_3374,N_5565);
nand U8154 (N_8154,N_3342,N_3813);
or U8155 (N_8155,N_4853,N_3331);
and U8156 (N_8156,N_3481,N_4649);
and U8157 (N_8157,N_3701,N_5684);
or U8158 (N_8158,N_3818,N_5826);
nand U8159 (N_8159,N_5990,N_4779);
and U8160 (N_8160,N_3880,N_5299);
nand U8161 (N_8161,N_5369,N_5153);
nor U8162 (N_8162,N_5386,N_5109);
or U8163 (N_8163,N_3869,N_3046);
or U8164 (N_8164,N_3198,N_3255);
nor U8165 (N_8165,N_4120,N_3851);
nor U8166 (N_8166,N_4049,N_5133);
and U8167 (N_8167,N_3479,N_4982);
or U8168 (N_8168,N_3065,N_4429);
nor U8169 (N_8169,N_3437,N_3606);
nand U8170 (N_8170,N_5681,N_3828);
and U8171 (N_8171,N_5374,N_5267);
nand U8172 (N_8172,N_4113,N_5369);
and U8173 (N_8173,N_5376,N_5680);
nand U8174 (N_8174,N_4449,N_5899);
nand U8175 (N_8175,N_3491,N_5817);
and U8176 (N_8176,N_5078,N_4453);
nor U8177 (N_8177,N_5685,N_4969);
and U8178 (N_8178,N_4406,N_4312);
nor U8179 (N_8179,N_5219,N_3104);
nand U8180 (N_8180,N_5839,N_5082);
and U8181 (N_8181,N_4631,N_4399);
nor U8182 (N_8182,N_5050,N_4237);
and U8183 (N_8183,N_3020,N_3059);
nor U8184 (N_8184,N_4144,N_3888);
nand U8185 (N_8185,N_4118,N_5604);
xnor U8186 (N_8186,N_5438,N_5834);
or U8187 (N_8187,N_3323,N_3999);
nand U8188 (N_8188,N_3925,N_5204);
nor U8189 (N_8189,N_3701,N_4012);
nand U8190 (N_8190,N_5278,N_4286);
nand U8191 (N_8191,N_5520,N_5743);
nor U8192 (N_8192,N_3999,N_3641);
and U8193 (N_8193,N_3927,N_3562);
nand U8194 (N_8194,N_4125,N_4877);
or U8195 (N_8195,N_5303,N_3295);
or U8196 (N_8196,N_5430,N_4547);
xnor U8197 (N_8197,N_3753,N_4041);
and U8198 (N_8198,N_5971,N_5856);
nand U8199 (N_8199,N_4685,N_3752);
xor U8200 (N_8200,N_4308,N_3235);
and U8201 (N_8201,N_5688,N_4621);
nor U8202 (N_8202,N_4640,N_4966);
and U8203 (N_8203,N_4895,N_5372);
or U8204 (N_8204,N_4743,N_5930);
nand U8205 (N_8205,N_3417,N_3430);
or U8206 (N_8206,N_4246,N_4194);
or U8207 (N_8207,N_3128,N_5378);
and U8208 (N_8208,N_4975,N_4553);
nand U8209 (N_8209,N_3272,N_3398);
or U8210 (N_8210,N_5355,N_4106);
nor U8211 (N_8211,N_3794,N_3953);
or U8212 (N_8212,N_4741,N_4453);
nand U8213 (N_8213,N_3086,N_4291);
and U8214 (N_8214,N_5712,N_4032);
or U8215 (N_8215,N_4950,N_4572);
xnor U8216 (N_8216,N_5396,N_5783);
nand U8217 (N_8217,N_4198,N_3107);
or U8218 (N_8218,N_3790,N_5071);
or U8219 (N_8219,N_4023,N_3877);
or U8220 (N_8220,N_4025,N_4436);
and U8221 (N_8221,N_3149,N_5040);
or U8222 (N_8222,N_3490,N_5869);
nor U8223 (N_8223,N_5012,N_4896);
and U8224 (N_8224,N_3734,N_4506);
nor U8225 (N_8225,N_3401,N_5043);
nand U8226 (N_8226,N_4680,N_3045);
nand U8227 (N_8227,N_5520,N_4291);
and U8228 (N_8228,N_4014,N_4449);
nand U8229 (N_8229,N_5225,N_5199);
or U8230 (N_8230,N_5370,N_4486);
and U8231 (N_8231,N_5297,N_4491);
and U8232 (N_8232,N_4645,N_3914);
and U8233 (N_8233,N_4358,N_3258);
and U8234 (N_8234,N_5854,N_4566);
nor U8235 (N_8235,N_5468,N_5061);
nor U8236 (N_8236,N_3673,N_5740);
or U8237 (N_8237,N_3338,N_4804);
or U8238 (N_8238,N_5029,N_3744);
or U8239 (N_8239,N_4608,N_5896);
and U8240 (N_8240,N_4175,N_5805);
or U8241 (N_8241,N_5686,N_3129);
nand U8242 (N_8242,N_3249,N_3402);
or U8243 (N_8243,N_3562,N_5392);
nand U8244 (N_8244,N_3363,N_3051);
nand U8245 (N_8245,N_5130,N_5887);
nand U8246 (N_8246,N_4601,N_3894);
nand U8247 (N_8247,N_4505,N_3886);
nand U8248 (N_8248,N_4447,N_5124);
or U8249 (N_8249,N_3313,N_5225);
and U8250 (N_8250,N_5981,N_3994);
or U8251 (N_8251,N_3110,N_4763);
or U8252 (N_8252,N_4237,N_4047);
and U8253 (N_8253,N_5041,N_4306);
and U8254 (N_8254,N_3909,N_5459);
nor U8255 (N_8255,N_5908,N_4607);
nor U8256 (N_8256,N_4930,N_3271);
nand U8257 (N_8257,N_3320,N_4212);
or U8258 (N_8258,N_5275,N_3934);
and U8259 (N_8259,N_5722,N_3479);
or U8260 (N_8260,N_4355,N_5009);
nand U8261 (N_8261,N_4168,N_3966);
and U8262 (N_8262,N_5695,N_3210);
or U8263 (N_8263,N_4198,N_3499);
xor U8264 (N_8264,N_4019,N_4459);
and U8265 (N_8265,N_4612,N_5012);
or U8266 (N_8266,N_4414,N_4008);
and U8267 (N_8267,N_4597,N_5705);
and U8268 (N_8268,N_3761,N_4058);
nand U8269 (N_8269,N_5629,N_3968);
xnor U8270 (N_8270,N_4018,N_5252);
or U8271 (N_8271,N_3180,N_3942);
or U8272 (N_8272,N_5503,N_5538);
or U8273 (N_8273,N_5352,N_3873);
nor U8274 (N_8274,N_5547,N_3776);
or U8275 (N_8275,N_5428,N_3745);
nor U8276 (N_8276,N_4473,N_5326);
xor U8277 (N_8277,N_4724,N_3799);
or U8278 (N_8278,N_3779,N_5619);
or U8279 (N_8279,N_5187,N_5364);
nand U8280 (N_8280,N_3530,N_3380);
and U8281 (N_8281,N_3322,N_5819);
and U8282 (N_8282,N_5380,N_4184);
nor U8283 (N_8283,N_3975,N_4741);
nand U8284 (N_8284,N_4916,N_3379);
or U8285 (N_8285,N_3236,N_3257);
nand U8286 (N_8286,N_4559,N_5995);
nand U8287 (N_8287,N_3770,N_5863);
nor U8288 (N_8288,N_4345,N_3012);
and U8289 (N_8289,N_3164,N_3289);
nor U8290 (N_8290,N_4973,N_3891);
or U8291 (N_8291,N_5669,N_3053);
or U8292 (N_8292,N_3566,N_4836);
and U8293 (N_8293,N_4414,N_4708);
and U8294 (N_8294,N_3772,N_4039);
or U8295 (N_8295,N_5471,N_5119);
xor U8296 (N_8296,N_5203,N_4044);
and U8297 (N_8297,N_5921,N_4778);
nor U8298 (N_8298,N_5534,N_5660);
nor U8299 (N_8299,N_3208,N_5450);
or U8300 (N_8300,N_4212,N_4953);
nand U8301 (N_8301,N_3497,N_4096);
nor U8302 (N_8302,N_3549,N_4913);
nor U8303 (N_8303,N_4074,N_3141);
nor U8304 (N_8304,N_4678,N_3188);
or U8305 (N_8305,N_5746,N_5907);
and U8306 (N_8306,N_5738,N_4370);
or U8307 (N_8307,N_5113,N_4511);
or U8308 (N_8308,N_4288,N_4475);
or U8309 (N_8309,N_4162,N_4335);
or U8310 (N_8310,N_5275,N_3584);
or U8311 (N_8311,N_3782,N_4739);
and U8312 (N_8312,N_5583,N_4956);
and U8313 (N_8313,N_4884,N_3251);
nand U8314 (N_8314,N_3964,N_3297);
nand U8315 (N_8315,N_4024,N_3830);
nor U8316 (N_8316,N_3895,N_5936);
nor U8317 (N_8317,N_4137,N_3415);
xor U8318 (N_8318,N_5592,N_4293);
xor U8319 (N_8319,N_3999,N_3635);
or U8320 (N_8320,N_4427,N_5614);
nor U8321 (N_8321,N_3839,N_5363);
and U8322 (N_8322,N_3644,N_5068);
or U8323 (N_8323,N_5752,N_4798);
nor U8324 (N_8324,N_3502,N_3895);
nand U8325 (N_8325,N_3202,N_3649);
nor U8326 (N_8326,N_5079,N_4803);
and U8327 (N_8327,N_3345,N_4818);
and U8328 (N_8328,N_5586,N_5145);
and U8329 (N_8329,N_5840,N_4507);
nor U8330 (N_8330,N_3858,N_4289);
nor U8331 (N_8331,N_4653,N_3551);
and U8332 (N_8332,N_3949,N_4101);
nor U8333 (N_8333,N_4283,N_4133);
nor U8334 (N_8334,N_4892,N_3727);
nor U8335 (N_8335,N_5367,N_5335);
nand U8336 (N_8336,N_4968,N_5423);
xnor U8337 (N_8337,N_3885,N_4268);
and U8338 (N_8338,N_5838,N_4198);
nand U8339 (N_8339,N_3249,N_5884);
nand U8340 (N_8340,N_3027,N_4015);
or U8341 (N_8341,N_4268,N_3516);
nor U8342 (N_8342,N_3501,N_5870);
and U8343 (N_8343,N_4447,N_5469);
or U8344 (N_8344,N_5446,N_3950);
and U8345 (N_8345,N_5858,N_3374);
nor U8346 (N_8346,N_4209,N_4790);
nor U8347 (N_8347,N_3169,N_5511);
nand U8348 (N_8348,N_4487,N_4779);
xor U8349 (N_8349,N_4972,N_4221);
and U8350 (N_8350,N_3687,N_5542);
and U8351 (N_8351,N_3371,N_4228);
and U8352 (N_8352,N_5120,N_4137);
and U8353 (N_8353,N_3230,N_4824);
nor U8354 (N_8354,N_3251,N_5354);
and U8355 (N_8355,N_4648,N_5643);
nand U8356 (N_8356,N_4897,N_4377);
or U8357 (N_8357,N_3938,N_4655);
or U8358 (N_8358,N_3338,N_3292);
nor U8359 (N_8359,N_5348,N_3116);
and U8360 (N_8360,N_3088,N_5179);
or U8361 (N_8361,N_5024,N_4418);
nor U8362 (N_8362,N_3696,N_4398);
nand U8363 (N_8363,N_4993,N_5335);
and U8364 (N_8364,N_5886,N_3569);
nand U8365 (N_8365,N_4767,N_3123);
or U8366 (N_8366,N_3936,N_4587);
and U8367 (N_8367,N_5943,N_5097);
nand U8368 (N_8368,N_4259,N_5604);
nor U8369 (N_8369,N_4663,N_5925);
or U8370 (N_8370,N_5547,N_3497);
nand U8371 (N_8371,N_3640,N_5165);
or U8372 (N_8372,N_3205,N_5924);
and U8373 (N_8373,N_5071,N_4375);
or U8374 (N_8374,N_5168,N_3826);
and U8375 (N_8375,N_3635,N_4023);
nor U8376 (N_8376,N_5065,N_4322);
nand U8377 (N_8377,N_4200,N_4090);
nor U8378 (N_8378,N_4009,N_5323);
and U8379 (N_8379,N_3076,N_5602);
nand U8380 (N_8380,N_5428,N_3956);
and U8381 (N_8381,N_5561,N_4582);
xnor U8382 (N_8382,N_3808,N_5086);
nand U8383 (N_8383,N_4930,N_4546);
and U8384 (N_8384,N_5561,N_5580);
nor U8385 (N_8385,N_3034,N_4347);
and U8386 (N_8386,N_3010,N_4670);
nor U8387 (N_8387,N_4231,N_3931);
and U8388 (N_8388,N_5435,N_4221);
and U8389 (N_8389,N_4451,N_4446);
xor U8390 (N_8390,N_4743,N_3642);
and U8391 (N_8391,N_5666,N_5725);
or U8392 (N_8392,N_4013,N_4314);
and U8393 (N_8393,N_3775,N_4135);
and U8394 (N_8394,N_3373,N_4149);
and U8395 (N_8395,N_4886,N_4739);
or U8396 (N_8396,N_4572,N_4579);
and U8397 (N_8397,N_5956,N_4826);
or U8398 (N_8398,N_5821,N_5386);
or U8399 (N_8399,N_3353,N_3127);
or U8400 (N_8400,N_5646,N_4247);
nand U8401 (N_8401,N_5482,N_5818);
or U8402 (N_8402,N_3282,N_5494);
nand U8403 (N_8403,N_3686,N_5330);
nand U8404 (N_8404,N_4717,N_5434);
and U8405 (N_8405,N_5778,N_4916);
or U8406 (N_8406,N_3176,N_5413);
and U8407 (N_8407,N_5027,N_3869);
or U8408 (N_8408,N_5407,N_5221);
nor U8409 (N_8409,N_3726,N_4277);
or U8410 (N_8410,N_3690,N_3208);
nor U8411 (N_8411,N_3548,N_3971);
nand U8412 (N_8412,N_5881,N_4014);
and U8413 (N_8413,N_4166,N_4041);
nor U8414 (N_8414,N_3823,N_3335);
nand U8415 (N_8415,N_5664,N_5612);
nor U8416 (N_8416,N_3500,N_3068);
or U8417 (N_8417,N_4466,N_4128);
nand U8418 (N_8418,N_3478,N_3102);
nor U8419 (N_8419,N_5853,N_3648);
and U8420 (N_8420,N_3075,N_4849);
or U8421 (N_8421,N_5626,N_5013);
and U8422 (N_8422,N_3796,N_5281);
nor U8423 (N_8423,N_3546,N_5314);
nand U8424 (N_8424,N_4189,N_3580);
nand U8425 (N_8425,N_3086,N_3253);
or U8426 (N_8426,N_3690,N_3551);
nand U8427 (N_8427,N_4671,N_3504);
and U8428 (N_8428,N_3238,N_5690);
nand U8429 (N_8429,N_3289,N_3943);
nand U8430 (N_8430,N_3254,N_4506);
nor U8431 (N_8431,N_3910,N_3402);
nor U8432 (N_8432,N_3086,N_4835);
or U8433 (N_8433,N_3280,N_4654);
nand U8434 (N_8434,N_3877,N_3378);
or U8435 (N_8435,N_4501,N_4019);
nor U8436 (N_8436,N_4114,N_4500);
nor U8437 (N_8437,N_3131,N_3978);
or U8438 (N_8438,N_4841,N_4663);
or U8439 (N_8439,N_5702,N_5121);
and U8440 (N_8440,N_5267,N_5300);
nor U8441 (N_8441,N_5825,N_5237);
xnor U8442 (N_8442,N_4559,N_5745);
and U8443 (N_8443,N_3582,N_4317);
or U8444 (N_8444,N_5671,N_3917);
or U8445 (N_8445,N_4752,N_4949);
or U8446 (N_8446,N_3681,N_5231);
and U8447 (N_8447,N_3675,N_3417);
nand U8448 (N_8448,N_4170,N_5527);
and U8449 (N_8449,N_5383,N_3315);
nor U8450 (N_8450,N_5578,N_5706);
or U8451 (N_8451,N_4230,N_4243);
nand U8452 (N_8452,N_4611,N_4350);
nor U8453 (N_8453,N_5506,N_3746);
nand U8454 (N_8454,N_4912,N_4951);
nor U8455 (N_8455,N_3868,N_4215);
and U8456 (N_8456,N_4003,N_4840);
or U8457 (N_8457,N_5826,N_4717);
and U8458 (N_8458,N_3525,N_4983);
or U8459 (N_8459,N_5123,N_3566);
nor U8460 (N_8460,N_3499,N_3310);
or U8461 (N_8461,N_5524,N_3943);
nor U8462 (N_8462,N_5899,N_5895);
xnor U8463 (N_8463,N_5732,N_5159);
xor U8464 (N_8464,N_4148,N_4494);
nor U8465 (N_8465,N_4038,N_3221);
nand U8466 (N_8466,N_3196,N_4318);
nor U8467 (N_8467,N_5820,N_4514);
and U8468 (N_8468,N_4580,N_3496);
and U8469 (N_8469,N_5552,N_5535);
and U8470 (N_8470,N_3007,N_3159);
nand U8471 (N_8471,N_5504,N_5326);
or U8472 (N_8472,N_3469,N_5674);
or U8473 (N_8473,N_4255,N_4185);
nand U8474 (N_8474,N_3270,N_3853);
nand U8475 (N_8475,N_3037,N_3241);
nor U8476 (N_8476,N_5298,N_3737);
nor U8477 (N_8477,N_5528,N_5111);
nand U8478 (N_8478,N_4471,N_3168);
or U8479 (N_8479,N_3589,N_5898);
nand U8480 (N_8480,N_5545,N_4761);
nand U8481 (N_8481,N_4871,N_4533);
nand U8482 (N_8482,N_4899,N_4232);
and U8483 (N_8483,N_4949,N_5931);
nand U8484 (N_8484,N_5820,N_5932);
nand U8485 (N_8485,N_3955,N_4956);
or U8486 (N_8486,N_4925,N_5635);
xnor U8487 (N_8487,N_3229,N_5046);
nand U8488 (N_8488,N_3351,N_5136);
and U8489 (N_8489,N_4014,N_4686);
nor U8490 (N_8490,N_4071,N_3499);
or U8491 (N_8491,N_4845,N_3396);
nand U8492 (N_8492,N_5341,N_3114);
nor U8493 (N_8493,N_5979,N_3641);
nor U8494 (N_8494,N_4148,N_3116);
and U8495 (N_8495,N_5338,N_3731);
or U8496 (N_8496,N_4509,N_3541);
nand U8497 (N_8497,N_5179,N_4356);
nand U8498 (N_8498,N_5189,N_3312);
and U8499 (N_8499,N_5877,N_4917);
nor U8500 (N_8500,N_3168,N_4858);
nor U8501 (N_8501,N_4193,N_3828);
nor U8502 (N_8502,N_5439,N_3656);
nor U8503 (N_8503,N_3373,N_5927);
or U8504 (N_8504,N_3425,N_5002);
nor U8505 (N_8505,N_3729,N_3717);
nand U8506 (N_8506,N_3123,N_3607);
nor U8507 (N_8507,N_4281,N_5448);
and U8508 (N_8508,N_3906,N_3068);
and U8509 (N_8509,N_4546,N_5977);
nor U8510 (N_8510,N_3315,N_5081);
or U8511 (N_8511,N_4600,N_3855);
and U8512 (N_8512,N_3080,N_3519);
nand U8513 (N_8513,N_3593,N_4911);
nor U8514 (N_8514,N_3792,N_5270);
nand U8515 (N_8515,N_5453,N_3232);
nor U8516 (N_8516,N_4127,N_5286);
nand U8517 (N_8517,N_3996,N_4306);
and U8518 (N_8518,N_3752,N_4150);
nor U8519 (N_8519,N_5218,N_4368);
and U8520 (N_8520,N_4132,N_5293);
and U8521 (N_8521,N_5337,N_3763);
nand U8522 (N_8522,N_3397,N_5686);
and U8523 (N_8523,N_5336,N_5051);
nand U8524 (N_8524,N_5070,N_3148);
or U8525 (N_8525,N_4299,N_4716);
and U8526 (N_8526,N_3322,N_4496);
and U8527 (N_8527,N_5827,N_3895);
or U8528 (N_8528,N_3951,N_4777);
or U8529 (N_8529,N_4547,N_3000);
nor U8530 (N_8530,N_5960,N_4934);
and U8531 (N_8531,N_4323,N_5420);
xor U8532 (N_8532,N_3300,N_3366);
xor U8533 (N_8533,N_5812,N_3788);
or U8534 (N_8534,N_3339,N_5304);
or U8535 (N_8535,N_5923,N_4033);
and U8536 (N_8536,N_3776,N_4564);
or U8537 (N_8537,N_5220,N_3361);
nand U8538 (N_8538,N_5036,N_3509);
nor U8539 (N_8539,N_3982,N_4540);
xnor U8540 (N_8540,N_4024,N_3820);
xnor U8541 (N_8541,N_4963,N_4344);
xnor U8542 (N_8542,N_3843,N_3296);
or U8543 (N_8543,N_4358,N_5001);
or U8544 (N_8544,N_4406,N_5609);
nand U8545 (N_8545,N_5638,N_4935);
or U8546 (N_8546,N_3878,N_3033);
and U8547 (N_8547,N_3586,N_5655);
nor U8548 (N_8548,N_3018,N_4257);
or U8549 (N_8549,N_4279,N_3224);
nor U8550 (N_8550,N_5766,N_3756);
nand U8551 (N_8551,N_5547,N_3758);
nand U8552 (N_8552,N_5438,N_3079);
and U8553 (N_8553,N_4262,N_4728);
and U8554 (N_8554,N_3884,N_4040);
and U8555 (N_8555,N_5562,N_3140);
or U8556 (N_8556,N_3114,N_3991);
or U8557 (N_8557,N_4344,N_4766);
nor U8558 (N_8558,N_3149,N_4557);
or U8559 (N_8559,N_3900,N_5869);
nand U8560 (N_8560,N_5224,N_5227);
and U8561 (N_8561,N_3595,N_5771);
or U8562 (N_8562,N_3749,N_3940);
or U8563 (N_8563,N_4186,N_3521);
and U8564 (N_8564,N_4697,N_4221);
nor U8565 (N_8565,N_4146,N_4221);
and U8566 (N_8566,N_5186,N_4219);
or U8567 (N_8567,N_5605,N_4955);
nand U8568 (N_8568,N_4219,N_4532);
and U8569 (N_8569,N_5388,N_3969);
or U8570 (N_8570,N_4892,N_5223);
nor U8571 (N_8571,N_3008,N_4507);
or U8572 (N_8572,N_4804,N_3478);
nor U8573 (N_8573,N_5442,N_5585);
nor U8574 (N_8574,N_3909,N_3078);
nand U8575 (N_8575,N_5108,N_3552);
or U8576 (N_8576,N_4005,N_4028);
nor U8577 (N_8577,N_4758,N_5685);
xnor U8578 (N_8578,N_3058,N_3793);
nor U8579 (N_8579,N_3052,N_5031);
or U8580 (N_8580,N_3163,N_3263);
or U8581 (N_8581,N_4797,N_4285);
and U8582 (N_8582,N_3293,N_4321);
and U8583 (N_8583,N_4523,N_5438);
nand U8584 (N_8584,N_5392,N_4086);
nor U8585 (N_8585,N_3804,N_4388);
nor U8586 (N_8586,N_4471,N_3662);
and U8587 (N_8587,N_5827,N_3514);
nand U8588 (N_8588,N_3517,N_5548);
nand U8589 (N_8589,N_3297,N_4321);
nand U8590 (N_8590,N_4181,N_5158);
or U8591 (N_8591,N_5722,N_5056);
and U8592 (N_8592,N_3332,N_3861);
nand U8593 (N_8593,N_3919,N_3536);
nand U8594 (N_8594,N_4510,N_5733);
nand U8595 (N_8595,N_4925,N_4247);
or U8596 (N_8596,N_5505,N_3816);
or U8597 (N_8597,N_4795,N_5118);
and U8598 (N_8598,N_5487,N_3581);
or U8599 (N_8599,N_3455,N_3735);
xnor U8600 (N_8600,N_5465,N_5527);
and U8601 (N_8601,N_4657,N_3047);
and U8602 (N_8602,N_5267,N_3877);
and U8603 (N_8603,N_5117,N_3558);
or U8604 (N_8604,N_3632,N_4185);
nand U8605 (N_8605,N_3206,N_5652);
or U8606 (N_8606,N_3099,N_4702);
and U8607 (N_8607,N_4859,N_4351);
or U8608 (N_8608,N_5523,N_5827);
nor U8609 (N_8609,N_4239,N_5010);
nor U8610 (N_8610,N_5353,N_3566);
nand U8611 (N_8611,N_4348,N_4369);
nor U8612 (N_8612,N_3116,N_5908);
nand U8613 (N_8613,N_4173,N_5735);
nand U8614 (N_8614,N_3043,N_4725);
or U8615 (N_8615,N_3280,N_4196);
nand U8616 (N_8616,N_5675,N_3974);
or U8617 (N_8617,N_4381,N_4246);
nand U8618 (N_8618,N_5175,N_4780);
or U8619 (N_8619,N_5332,N_3406);
or U8620 (N_8620,N_5261,N_3515);
nand U8621 (N_8621,N_3067,N_4531);
nand U8622 (N_8622,N_3010,N_4995);
nand U8623 (N_8623,N_3782,N_3577);
nand U8624 (N_8624,N_3806,N_3134);
nand U8625 (N_8625,N_5479,N_5846);
nor U8626 (N_8626,N_3263,N_3085);
nand U8627 (N_8627,N_5638,N_5996);
or U8628 (N_8628,N_4044,N_5301);
nand U8629 (N_8629,N_4188,N_4505);
and U8630 (N_8630,N_5203,N_4591);
and U8631 (N_8631,N_5844,N_3614);
and U8632 (N_8632,N_5240,N_5359);
and U8633 (N_8633,N_3307,N_5067);
nor U8634 (N_8634,N_4293,N_3296);
or U8635 (N_8635,N_4919,N_5358);
nand U8636 (N_8636,N_5370,N_5561);
nand U8637 (N_8637,N_4176,N_3061);
and U8638 (N_8638,N_4871,N_4608);
nand U8639 (N_8639,N_5572,N_4634);
nand U8640 (N_8640,N_4583,N_5691);
nor U8641 (N_8641,N_3451,N_5985);
and U8642 (N_8642,N_4032,N_5285);
nor U8643 (N_8643,N_4545,N_3781);
nor U8644 (N_8644,N_3275,N_5062);
nand U8645 (N_8645,N_4105,N_4209);
and U8646 (N_8646,N_5282,N_3553);
and U8647 (N_8647,N_4097,N_3717);
nand U8648 (N_8648,N_5262,N_5209);
nand U8649 (N_8649,N_3221,N_4596);
and U8650 (N_8650,N_5301,N_4798);
and U8651 (N_8651,N_5470,N_5782);
nor U8652 (N_8652,N_5960,N_3507);
and U8653 (N_8653,N_4415,N_5778);
nand U8654 (N_8654,N_4400,N_4057);
or U8655 (N_8655,N_3829,N_5401);
nor U8656 (N_8656,N_3131,N_5360);
or U8657 (N_8657,N_3767,N_5899);
nor U8658 (N_8658,N_3588,N_3710);
nand U8659 (N_8659,N_3461,N_4079);
or U8660 (N_8660,N_3174,N_3085);
or U8661 (N_8661,N_4150,N_3597);
nor U8662 (N_8662,N_5030,N_4832);
nand U8663 (N_8663,N_4512,N_4288);
nand U8664 (N_8664,N_5189,N_5990);
and U8665 (N_8665,N_4388,N_5671);
or U8666 (N_8666,N_5973,N_4730);
nand U8667 (N_8667,N_5983,N_4143);
nand U8668 (N_8668,N_5244,N_3025);
or U8669 (N_8669,N_5846,N_4945);
nor U8670 (N_8670,N_3753,N_4536);
or U8671 (N_8671,N_3997,N_3008);
nand U8672 (N_8672,N_3648,N_5725);
nor U8673 (N_8673,N_4841,N_4464);
nand U8674 (N_8674,N_4857,N_3813);
nand U8675 (N_8675,N_3586,N_5542);
or U8676 (N_8676,N_3395,N_3889);
nand U8677 (N_8677,N_4370,N_4702);
nor U8678 (N_8678,N_3525,N_3282);
nand U8679 (N_8679,N_3397,N_5901);
or U8680 (N_8680,N_3859,N_5679);
and U8681 (N_8681,N_3599,N_3301);
nor U8682 (N_8682,N_5533,N_5034);
nand U8683 (N_8683,N_5409,N_3599);
nor U8684 (N_8684,N_4756,N_3757);
and U8685 (N_8685,N_3214,N_5963);
nand U8686 (N_8686,N_5894,N_5984);
nand U8687 (N_8687,N_4499,N_4200);
or U8688 (N_8688,N_4829,N_3731);
or U8689 (N_8689,N_3750,N_4972);
nor U8690 (N_8690,N_4050,N_4388);
and U8691 (N_8691,N_4942,N_4781);
nor U8692 (N_8692,N_4630,N_4458);
nor U8693 (N_8693,N_3244,N_4735);
nor U8694 (N_8694,N_4434,N_4679);
nor U8695 (N_8695,N_5006,N_4065);
or U8696 (N_8696,N_5522,N_3707);
nand U8697 (N_8697,N_4401,N_5264);
nand U8698 (N_8698,N_5434,N_5293);
and U8699 (N_8699,N_4405,N_5322);
xor U8700 (N_8700,N_5651,N_4935);
nand U8701 (N_8701,N_4696,N_5992);
and U8702 (N_8702,N_3430,N_3547);
and U8703 (N_8703,N_3800,N_3865);
or U8704 (N_8704,N_5355,N_5816);
and U8705 (N_8705,N_5844,N_3854);
nand U8706 (N_8706,N_3052,N_4010);
and U8707 (N_8707,N_3971,N_4039);
or U8708 (N_8708,N_5410,N_5953);
or U8709 (N_8709,N_4298,N_5718);
nor U8710 (N_8710,N_3653,N_3063);
or U8711 (N_8711,N_4127,N_3254);
or U8712 (N_8712,N_4010,N_4156);
or U8713 (N_8713,N_5931,N_5409);
and U8714 (N_8714,N_3003,N_5114);
and U8715 (N_8715,N_4635,N_5849);
or U8716 (N_8716,N_4923,N_3146);
nand U8717 (N_8717,N_3911,N_4689);
nor U8718 (N_8718,N_4413,N_4030);
nand U8719 (N_8719,N_5467,N_3765);
nor U8720 (N_8720,N_3818,N_3510);
nor U8721 (N_8721,N_5028,N_4367);
and U8722 (N_8722,N_4692,N_4685);
or U8723 (N_8723,N_3963,N_4813);
nor U8724 (N_8724,N_4665,N_3459);
nor U8725 (N_8725,N_5295,N_3143);
and U8726 (N_8726,N_5492,N_4583);
or U8727 (N_8727,N_3725,N_3310);
or U8728 (N_8728,N_3845,N_3026);
nand U8729 (N_8729,N_4239,N_4279);
nand U8730 (N_8730,N_5385,N_4565);
or U8731 (N_8731,N_4401,N_4114);
and U8732 (N_8732,N_5405,N_4602);
nor U8733 (N_8733,N_5348,N_4121);
or U8734 (N_8734,N_3539,N_5979);
and U8735 (N_8735,N_3206,N_4529);
nand U8736 (N_8736,N_3128,N_3855);
nor U8737 (N_8737,N_3425,N_5985);
nand U8738 (N_8738,N_5508,N_4358);
nand U8739 (N_8739,N_5055,N_3561);
and U8740 (N_8740,N_3042,N_5489);
nor U8741 (N_8741,N_5243,N_4395);
or U8742 (N_8742,N_5421,N_5427);
nand U8743 (N_8743,N_5013,N_3203);
nor U8744 (N_8744,N_4648,N_5860);
nor U8745 (N_8745,N_5198,N_5936);
nand U8746 (N_8746,N_5439,N_3987);
nor U8747 (N_8747,N_5641,N_3480);
and U8748 (N_8748,N_5017,N_3743);
or U8749 (N_8749,N_3007,N_5678);
or U8750 (N_8750,N_3225,N_3897);
or U8751 (N_8751,N_4999,N_5401);
or U8752 (N_8752,N_4223,N_4713);
or U8753 (N_8753,N_5846,N_3327);
or U8754 (N_8754,N_3483,N_3553);
nand U8755 (N_8755,N_5703,N_4825);
nor U8756 (N_8756,N_3296,N_5006);
or U8757 (N_8757,N_4418,N_3456);
and U8758 (N_8758,N_5832,N_3625);
nand U8759 (N_8759,N_4181,N_5972);
and U8760 (N_8760,N_3948,N_4825);
nand U8761 (N_8761,N_3597,N_4476);
or U8762 (N_8762,N_5458,N_5248);
or U8763 (N_8763,N_3433,N_3053);
or U8764 (N_8764,N_5869,N_5535);
nand U8765 (N_8765,N_3708,N_4833);
xor U8766 (N_8766,N_4789,N_4188);
nand U8767 (N_8767,N_3273,N_4979);
nor U8768 (N_8768,N_5381,N_3518);
nand U8769 (N_8769,N_5181,N_5146);
nand U8770 (N_8770,N_3733,N_4707);
nand U8771 (N_8771,N_4631,N_3757);
or U8772 (N_8772,N_4060,N_5120);
or U8773 (N_8773,N_4551,N_4381);
or U8774 (N_8774,N_4416,N_3896);
or U8775 (N_8775,N_4429,N_3680);
nor U8776 (N_8776,N_4560,N_5545);
nor U8777 (N_8777,N_4619,N_4161);
nand U8778 (N_8778,N_4944,N_4341);
or U8779 (N_8779,N_4843,N_3318);
and U8780 (N_8780,N_4163,N_5201);
and U8781 (N_8781,N_3063,N_4791);
nand U8782 (N_8782,N_3023,N_4979);
or U8783 (N_8783,N_3376,N_3346);
nand U8784 (N_8784,N_5416,N_3903);
or U8785 (N_8785,N_5554,N_4468);
nor U8786 (N_8786,N_4858,N_5326);
xnor U8787 (N_8787,N_5170,N_5209);
and U8788 (N_8788,N_5964,N_4363);
nand U8789 (N_8789,N_5480,N_3644);
nor U8790 (N_8790,N_5704,N_5682);
nor U8791 (N_8791,N_4945,N_3114);
or U8792 (N_8792,N_4591,N_4832);
nand U8793 (N_8793,N_5418,N_3927);
nand U8794 (N_8794,N_3716,N_5892);
and U8795 (N_8795,N_4310,N_4817);
and U8796 (N_8796,N_4479,N_5670);
nand U8797 (N_8797,N_3271,N_5285);
or U8798 (N_8798,N_5606,N_3844);
nor U8799 (N_8799,N_3337,N_3484);
or U8800 (N_8800,N_4714,N_4312);
or U8801 (N_8801,N_4128,N_4343);
or U8802 (N_8802,N_3659,N_5638);
or U8803 (N_8803,N_3312,N_3719);
nor U8804 (N_8804,N_4538,N_3086);
nor U8805 (N_8805,N_3890,N_3468);
nand U8806 (N_8806,N_3595,N_5327);
or U8807 (N_8807,N_5683,N_4768);
nand U8808 (N_8808,N_5231,N_3626);
nor U8809 (N_8809,N_3339,N_3448);
nand U8810 (N_8810,N_4319,N_4942);
or U8811 (N_8811,N_3646,N_3231);
nand U8812 (N_8812,N_3359,N_4692);
and U8813 (N_8813,N_4655,N_3679);
nor U8814 (N_8814,N_5368,N_5226);
or U8815 (N_8815,N_5790,N_3105);
nand U8816 (N_8816,N_5028,N_5040);
or U8817 (N_8817,N_3818,N_5338);
nor U8818 (N_8818,N_4630,N_4148);
and U8819 (N_8819,N_5819,N_3089);
xor U8820 (N_8820,N_4905,N_5765);
nor U8821 (N_8821,N_5274,N_3430);
nand U8822 (N_8822,N_4289,N_3446);
or U8823 (N_8823,N_3825,N_5607);
nand U8824 (N_8824,N_5599,N_3697);
and U8825 (N_8825,N_3052,N_5719);
or U8826 (N_8826,N_5663,N_3629);
nand U8827 (N_8827,N_4407,N_4309);
or U8828 (N_8828,N_4526,N_3325);
nand U8829 (N_8829,N_5516,N_4712);
nor U8830 (N_8830,N_4178,N_3384);
and U8831 (N_8831,N_5521,N_4613);
nor U8832 (N_8832,N_4920,N_3279);
or U8833 (N_8833,N_4550,N_4058);
nor U8834 (N_8834,N_5481,N_3083);
nor U8835 (N_8835,N_5618,N_4058);
nor U8836 (N_8836,N_3711,N_5599);
and U8837 (N_8837,N_3721,N_3690);
or U8838 (N_8838,N_5192,N_4793);
or U8839 (N_8839,N_4495,N_3856);
and U8840 (N_8840,N_4074,N_3010);
or U8841 (N_8841,N_5320,N_3073);
and U8842 (N_8842,N_4184,N_5126);
and U8843 (N_8843,N_4728,N_5792);
nor U8844 (N_8844,N_5253,N_5516);
or U8845 (N_8845,N_5123,N_4863);
or U8846 (N_8846,N_4373,N_5265);
nor U8847 (N_8847,N_4846,N_4848);
or U8848 (N_8848,N_3641,N_5045);
nor U8849 (N_8849,N_4586,N_3338);
and U8850 (N_8850,N_5067,N_3709);
or U8851 (N_8851,N_4254,N_5083);
and U8852 (N_8852,N_5168,N_5241);
nor U8853 (N_8853,N_5759,N_3986);
and U8854 (N_8854,N_4974,N_4146);
nand U8855 (N_8855,N_3078,N_5993);
and U8856 (N_8856,N_5390,N_3668);
or U8857 (N_8857,N_4238,N_4092);
or U8858 (N_8858,N_5985,N_5850);
nor U8859 (N_8859,N_3434,N_3868);
nor U8860 (N_8860,N_4790,N_4777);
or U8861 (N_8861,N_4168,N_3032);
and U8862 (N_8862,N_5181,N_3108);
nand U8863 (N_8863,N_5524,N_3877);
nand U8864 (N_8864,N_4833,N_4562);
nand U8865 (N_8865,N_5918,N_5188);
nor U8866 (N_8866,N_4055,N_4091);
or U8867 (N_8867,N_4588,N_3814);
or U8868 (N_8868,N_4693,N_5562);
nand U8869 (N_8869,N_3705,N_3266);
and U8870 (N_8870,N_4048,N_3021);
nand U8871 (N_8871,N_5986,N_3630);
and U8872 (N_8872,N_4058,N_3133);
nand U8873 (N_8873,N_3111,N_5542);
or U8874 (N_8874,N_5137,N_5262);
or U8875 (N_8875,N_4584,N_5940);
or U8876 (N_8876,N_5565,N_5013);
or U8877 (N_8877,N_3120,N_5012);
and U8878 (N_8878,N_5636,N_3228);
nand U8879 (N_8879,N_4980,N_4564);
and U8880 (N_8880,N_4372,N_3016);
xnor U8881 (N_8881,N_4286,N_4082);
nor U8882 (N_8882,N_4627,N_5786);
and U8883 (N_8883,N_3708,N_4208);
or U8884 (N_8884,N_5136,N_3376);
nand U8885 (N_8885,N_4791,N_4055);
nand U8886 (N_8886,N_3364,N_3366);
or U8887 (N_8887,N_5189,N_5896);
nand U8888 (N_8888,N_5635,N_4589);
nand U8889 (N_8889,N_3934,N_4726);
or U8890 (N_8890,N_3035,N_3461);
or U8891 (N_8891,N_4862,N_4594);
and U8892 (N_8892,N_5479,N_4886);
nor U8893 (N_8893,N_4749,N_3419);
nor U8894 (N_8894,N_4852,N_3326);
and U8895 (N_8895,N_5952,N_5820);
nand U8896 (N_8896,N_5855,N_4259);
nor U8897 (N_8897,N_5110,N_5712);
or U8898 (N_8898,N_3303,N_4869);
or U8899 (N_8899,N_5926,N_3666);
xnor U8900 (N_8900,N_3999,N_5815);
nor U8901 (N_8901,N_4890,N_4620);
nand U8902 (N_8902,N_5284,N_5533);
nand U8903 (N_8903,N_4486,N_4695);
nor U8904 (N_8904,N_3029,N_5078);
nand U8905 (N_8905,N_3391,N_4641);
or U8906 (N_8906,N_5863,N_4300);
nor U8907 (N_8907,N_4185,N_3323);
or U8908 (N_8908,N_4688,N_5880);
and U8909 (N_8909,N_3893,N_4381);
or U8910 (N_8910,N_3189,N_4898);
or U8911 (N_8911,N_4621,N_4354);
or U8912 (N_8912,N_3438,N_3536);
nor U8913 (N_8913,N_4514,N_5780);
or U8914 (N_8914,N_5440,N_5149);
or U8915 (N_8915,N_4617,N_4164);
or U8916 (N_8916,N_3759,N_3008);
nand U8917 (N_8917,N_4474,N_5175);
nand U8918 (N_8918,N_4997,N_5112);
nor U8919 (N_8919,N_3626,N_4576);
and U8920 (N_8920,N_5508,N_5891);
or U8921 (N_8921,N_4375,N_5763);
or U8922 (N_8922,N_4274,N_3113);
xnor U8923 (N_8923,N_4341,N_5249);
or U8924 (N_8924,N_4413,N_4869);
and U8925 (N_8925,N_4182,N_5908);
nor U8926 (N_8926,N_5555,N_5953);
and U8927 (N_8927,N_3194,N_3501);
nor U8928 (N_8928,N_5178,N_5836);
nor U8929 (N_8929,N_3600,N_4660);
nand U8930 (N_8930,N_4961,N_5811);
nand U8931 (N_8931,N_5627,N_4483);
and U8932 (N_8932,N_5935,N_3297);
nor U8933 (N_8933,N_3137,N_3139);
nand U8934 (N_8934,N_5079,N_5275);
nor U8935 (N_8935,N_4662,N_4481);
nor U8936 (N_8936,N_4075,N_4638);
and U8937 (N_8937,N_3939,N_4475);
or U8938 (N_8938,N_3046,N_3850);
or U8939 (N_8939,N_3466,N_5342);
and U8940 (N_8940,N_4114,N_4941);
or U8941 (N_8941,N_3581,N_4633);
or U8942 (N_8942,N_3312,N_3487);
nor U8943 (N_8943,N_4963,N_3585);
xnor U8944 (N_8944,N_3873,N_3788);
or U8945 (N_8945,N_5134,N_3306);
and U8946 (N_8946,N_4916,N_4316);
or U8947 (N_8947,N_3298,N_3815);
and U8948 (N_8948,N_4566,N_4255);
nand U8949 (N_8949,N_4137,N_3537);
and U8950 (N_8950,N_5279,N_3733);
nor U8951 (N_8951,N_3999,N_3038);
and U8952 (N_8952,N_3354,N_3973);
nor U8953 (N_8953,N_3560,N_3847);
xor U8954 (N_8954,N_3115,N_3238);
nor U8955 (N_8955,N_5568,N_4279);
and U8956 (N_8956,N_5554,N_5866);
nor U8957 (N_8957,N_3596,N_4990);
nor U8958 (N_8958,N_4252,N_4017);
and U8959 (N_8959,N_4330,N_3137);
and U8960 (N_8960,N_5410,N_4591);
or U8961 (N_8961,N_3633,N_3356);
nor U8962 (N_8962,N_3675,N_4296);
nor U8963 (N_8963,N_3395,N_3176);
and U8964 (N_8964,N_3008,N_4403);
nor U8965 (N_8965,N_5303,N_3049);
nor U8966 (N_8966,N_4911,N_3022);
or U8967 (N_8967,N_4378,N_3236);
xor U8968 (N_8968,N_4226,N_3060);
nand U8969 (N_8969,N_5399,N_5499);
or U8970 (N_8970,N_4051,N_3008);
nand U8971 (N_8971,N_4514,N_5153);
or U8972 (N_8972,N_3432,N_3642);
and U8973 (N_8973,N_4571,N_5307);
nor U8974 (N_8974,N_4671,N_3594);
nor U8975 (N_8975,N_3514,N_4069);
nor U8976 (N_8976,N_5404,N_5889);
and U8977 (N_8977,N_5025,N_4748);
nand U8978 (N_8978,N_4731,N_3635);
or U8979 (N_8979,N_5227,N_5137);
nor U8980 (N_8980,N_5139,N_4586);
nor U8981 (N_8981,N_5636,N_3464);
or U8982 (N_8982,N_4702,N_3247);
and U8983 (N_8983,N_3386,N_5337);
and U8984 (N_8984,N_5009,N_3884);
nand U8985 (N_8985,N_3334,N_5917);
nor U8986 (N_8986,N_3233,N_4510);
or U8987 (N_8987,N_4483,N_3438);
and U8988 (N_8988,N_4945,N_4082);
and U8989 (N_8989,N_4054,N_3667);
nand U8990 (N_8990,N_3564,N_4976);
nand U8991 (N_8991,N_5536,N_5416);
or U8992 (N_8992,N_3390,N_5899);
or U8993 (N_8993,N_3283,N_4031);
or U8994 (N_8994,N_4488,N_5480);
nor U8995 (N_8995,N_3459,N_5390);
or U8996 (N_8996,N_4902,N_3376);
nand U8997 (N_8997,N_3805,N_3131);
nor U8998 (N_8998,N_5416,N_3168);
nand U8999 (N_8999,N_5983,N_5985);
nor U9000 (N_9000,N_7553,N_7305);
and U9001 (N_9001,N_6062,N_8153);
nand U9002 (N_9002,N_8361,N_6936);
nand U9003 (N_9003,N_7357,N_7636);
or U9004 (N_9004,N_8898,N_6508);
or U9005 (N_9005,N_6781,N_6960);
nand U9006 (N_9006,N_6362,N_7383);
nor U9007 (N_9007,N_6877,N_6043);
and U9008 (N_9008,N_8467,N_6899);
or U9009 (N_9009,N_8779,N_7818);
or U9010 (N_9010,N_7143,N_6582);
nor U9011 (N_9011,N_8428,N_7466);
and U9012 (N_9012,N_8638,N_7049);
and U9013 (N_9013,N_6669,N_8941);
nor U9014 (N_9014,N_8372,N_8060);
xor U9015 (N_9015,N_6096,N_7483);
and U9016 (N_9016,N_8148,N_6600);
nand U9017 (N_9017,N_7887,N_7460);
and U9018 (N_9018,N_6882,N_8750);
or U9019 (N_9019,N_7931,N_7408);
nand U9020 (N_9020,N_6097,N_7214);
nand U9021 (N_9021,N_8554,N_6547);
nor U9022 (N_9022,N_8850,N_7212);
and U9023 (N_9023,N_6870,N_8838);
or U9024 (N_9024,N_8120,N_8589);
nor U9025 (N_9025,N_8393,N_6796);
or U9026 (N_9026,N_8913,N_7651);
nand U9027 (N_9027,N_6159,N_6701);
nand U9028 (N_9028,N_8548,N_6550);
or U9029 (N_9029,N_8522,N_8977);
and U9030 (N_9030,N_7325,N_6304);
nor U9031 (N_9031,N_7092,N_7421);
nand U9032 (N_9032,N_7938,N_8640);
nor U9033 (N_9033,N_8930,N_8403);
nor U9034 (N_9034,N_8788,N_8785);
and U9035 (N_9035,N_8727,N_7500);
or U9036 (N_9036,N_7086,N_6680);
nand U9037 (N_9037,N_6921,N_7004);
and U9038 (N_9038,N_6203,N_8461);
and U9039 (N_9039,N_8127,N_6045);
xor U9040 (N_9040,N_8248,N_6109);
nor U9041 (N_9041,N_8162,N_6447);
xor U9042 (N_9042,N_6070,N_7803);
and U9043 (N_9043,N_7504,N_8019);
nor U9044 (N_9044,N_6965,N_8365);
or U9045 (N_9045,N_6033,N_7259);
or U9046 (N_9046,N_6213,N_7193);
nand U9047 (N_9047,N_8689,N_6682);
nor U9048 (N_9048,N_6040,N_6923);
or U9049 (N_9049,N_6641,N_8831);
or U9050 (N_9050,N_6256,N_8613);
or U9051 (N_9051,N_8944,N_6349);
or U9052 (N_9052,N_7933,N_7414);
xor U9053 (N_9053,N_6355,N_8732);
nand U9054 (N_9054,N_7463,N_6080);
nand U9055 (N_9055,N_6453,N_7334);
nor U9056 (N_9056,N_6254,N_8796);
nand U9057 (N_9057,N_6897,N_6873);
nor U9058 (N_9058,N_7542,N_7409);
nand U9059 (N_9059,N_8111,N_8812);
or U9060 (N_9060,N_8581,N_7951);
nand U9061 (N_9061,N_8752,N_6719);
nand U9062 (N_9062,N_7566,N_6412);
xor U9063 (N_9063,N_6761,N_8423);
or U9064 (N_9064,N_8511,N_7210);
nor U9065 (N_9065,N_8299,N_6674);
or U9066 (N_9066,N_6335,N_8059);
or U9067 (N_9067,N_7755,N_6057);
or U9068 (N_9068,N_7665,N_7967);
xor U9069 (N_9069,N_7908,N_7101);
or U9070 (N_9070,N_6437,N_6200);
nor U9071 (N_9071,N_7100,N_7759);
or U9072 (N_9072,N_6857,N_7019);
nor U9073 (N_9073,N_8792,N_8506);
and U9074 (N_9074,N_7794,N_7679);
nor U9075 (N_9075,N_7142,N_7717);
or U9076 (N_9076,N_8904,N_7940);
and U9077 (N_9077,N_7944,N_6458);
nor U9078 (N_9078,N_6117,N_8591);
nand U9079 (N_9079,N_6121,N_6614);
nor U9080 (N_9080,N_8586,N_7351);
and U9081 (N_9081,N_8290,N_7688);
nor U9082 (N_9082,N_6445,N_8606);
nor U9083 (N_9083,N_6378,N_8495);
and U9084 (N_9084,N_8707,N_8834);
or U9085 (N_9085,N_8772,N_6177);
and U9086 (N_9086,N_6773,N_7986);
or U9087 (N_9087,N_7451,N_6691);
and U9088 (N_9088,N_7180,N_6481);
nand U9089 (N_9089,N_6717,N_6257);
or U9090 (N_9090,N_7691,N_8949);
and U9091 (N_9091,N_6367,N_6364);
xor U9092 (N_9092,N_7709,N_7001);
nor U9093 (N_9093,N_8966,N_6460);
nor U9094 (N_9094,N_8265,N_6132);
xnor U9095 (N_9095,N_8339,N_7878);
nand U9096 (N_9096,N_8442,N_6363);
xnor U9097 (N_9097,N_8194,N_6373);
nor U9098 (N_9098,N_6424,N_6498);
nand U9099 (N_9099,N_8722,N_7747);
and U9100 (N_9100,N_8536,N_6069);
or U9101 (N_9101,N_8616,N_8680);
nor U9102 (N_9102,N_7237,N_8252);
and U9103 (N_9103,N_8870,N_7309);
nand U9104 (N_9104,N_8644,N_8537);
and U9105 (N_9105,N_8446,N_8912);
nand U9106 (N_9106,N_8953,N_6459);
nor U9107 (N_9107,N_6598,N_6782);
xor U9108 (N_9108,N_7094,N_8603);
nand U9109 (N_9109,N_8106,N_6461);
nand U9110 (N_9110,N_8086,N_6210);
nor U9111 (N_9111,N_8380,N_8142);
xor U9112 (N_9112,N_6162,N_8227);
or U9113 (N_9113,N_6737,N_8013);
or U9114 (N_9114,N_8432,N_6654);
nor U9115 (N_9115,N_7563,N_7356);
and U9116 (N_9116,N_6065,N_6799);
or U9117 (N_9117,N_7645,N_6830);
and U9118 (N_9118,N_6837,N_6038);
or U9119 (N_9119,N_8183,N_8512);
or U9120 (N_9120,N_6934,N_8447);
xor U9121 (N_9121,N_6995,N_8806);
and U9122 (N_9122,N_8645,N_8824);
nor U9123 (N_9123,N_7576,N_6665);
and U9124 (N_9124,N_7946,N_8328);
or U9125 (N_9125,N_7216,N_8138);
nor U9126 (N_9126,N_7233,N_8196);
and U9127 (N_9127,N_6049,N_6146);
or U9128 (N_9128,N_7162,N_7958);
or U9129 (N_9129,N_8344,N_7410);
nand U9130 (N_9130,N_7798,N_7978);
and U9131 (N_9131,N_6432,N_6279);
nand U9132 (N_9132,N_7883,N_6945);
or U9133 (N_9133,N_8657,N_6968);
or U9134 (N_9134,N_8452,N_7917);
and U9135 (N_9135,N_7980,N_7033);
nand U9136 (N_9136,N_7664,N_6677);
or U9137 (N_9137,N_6115,N_8787);
and U9138 (N_9138,N_8297,N_6720);
nand U9139 (N_9139,N_6532,N_8542);
or U9140 (N_9140,N_6606,N_8139);
nor U9141 (N_9141,N_6118,N_8797);
and U9142 (N_9142,N_7849,N_6884);
or U9143 (N_9143,N_7150,N_7997);
and U9144 (N_9144,N_7468,N_6484);
or U9145 (N_9145,N_8291,N_8090);
and U9146 (N_9146,N_7670,N_7415);
and U9147 (N_9147,N_7718,N_7523);
nor U9148 (N_9148,N_7027,N_6535);
nor U9149 (N_9149,N_8652,N_6875);
or U9150 (N_9150,N_7526,N_7970);
nor U9151 (N_9151,N_7634,N_8596);
and U9152 (N_9152,N_7554,N_6134);
nand U9153 (N_9153,N_6000,N_8822);
or U9154 (N_9154,N_8763,N_6268);
or U9155 (N_9155,N_7559,N_6905);
nor U9156 (N_9156,N_6061,N_6091);
and U9157 (N_9157,N_7923,N_8879);
nor U9158 (N_9158,N_8818,N_7083);
and U9159 (N_9159,N_6433,N_7249);
nand U9160 (N_9160,N_6483,N_8778);
nor U9161 (N_9161,N_6170,N_8985);
and U9162 (N_9162,N_8597,N_8078);
nand U9163 (N_9163,N_8798,N_7771);
nand U9164 (N_9164,N_7624,N_6456);
or U9165 (N_9165,N_7400,N_7306);
and U9166 (N_9166,N_6812,N_6738);
or U9167 (N_9167,N_8015,N_7821);
and U9168 (N_9168,N_8206,N_6314);
and U9169 (N_9169,N_8696,N_7762);
nand U9170 (N_9170,N_7613,N_6077);
nand U9171 (N_9171,N_6151,N_7165);
nand U9172 (N_9172,N_6999,N_6730);
or U9173 (N_9173,N_6026,N_7630);
xnor U9174 (N_9174,N_8678,N_7112);
or U9175 (N_9175,N_7708,N_8523);
or U9176 (N_9176,N_6591,N_6551);
and U9177 (N_9177,N_8402,N_7437);
nand U9178 (N_9178,N_7653,N_7682);
or U9179 (N_9179,N_7797,N_6615);
and U9180 (N_9180,N_8832,N_6222);
nor U9181 (N_9181,N_6122,N_6495);
nand U9182 (N_9182,N_7328,N_6107);
and U9183 (N_9183,N_8909,N_6834);
or U9184 (N_9184,N_8287,N_6455);
nor U9185 (N_9185,N_8395,N_6332);
nand U9186 (N_9186,N_6369,N_8427);
and U9187 (N_9187,N_6711,N_6172);
or U9188 (N_9188,N_6813,N_7293);
nor U9189 (N_9189,N_8840,N_8802);
and U9190 (N_9190,N_6755,N_8864);
and U9191 (N_9191,N_7000,N_6180);
and U9192 (N_9192,N_7099,N_8045);
nor U9193 (N_9193,N_7612,N_8959);
and U9194 (N_9194,N_8373,N_6868);
or U9195 (N_9195,N_6129,N_7181);
and U9196 (N_9196,N_6793,N_7564);
and U9197 (N_9197,N_7174,N_7643);
xor U9198 (N_9198,N_7372,N_6404);
nand U9199 (N_9199,N_7315,N_7528);
nor U9200 (N_9200,N_6540,N_7584);
or U9201 (N_9201,N_8988,N_8410);
nand U9202 (N_9202,N_8226,N_8711);
nor U9203 (N_9203,N_8841,N_7109);
nor U9204 (N_9204,N_6305,N_8048);
and U9205 (N_9205,N_7657,N_7440);
xnor U9206 (N_9206,N_8209,N_8004);
or U9207 (N_9207,N_6165,N_7031);
nand U9208 (N_9208,N_8407,N_8418);
and U9209 (N_9209,N_6524,N_7072);
or U9210 (N_9210,N_6673,N_6021);
nand U9211 (N_9211,N_7623,N_8621);
nor U9212 (N_9212,N_8574,N_7711);
or U9213 (N_9213,N_6864,N_8530);
or U9214 (N_9214,N_8963,N_7188);
or U9215 (N_9215,N_8334,N_8992);
nand U9216 (N_9216,N_6291,N_7186);
nor U9217 (N_9217,N_8136,N_6734);
nand U9218 (N_9218,N_6729,N_7561);
nor U9219 (N_9219,N_8243,N_8939);
and U9220 (N_9220,N_7405,N_8911);
nand U9221 (N_9221,N_7605,N_6224);
and U9222 (N_9222,N_6478,N_7407);
nand U9223 (N_9223,N_6321,N_7458);
nand U9224 (N_9224,N_8774,N_7982);
and U9225 (N_9225,N_7920,N_7501);
or U9226 (N_9226,N_6164,N_7135);
nand U9227 (N_9227,N_7377,N_6209);
and U9228 (N_9228,N_8999,N_8814);
and U9229 (N_9229,N_6539,N_8490);
and U9230 (N_9230,N_6388,N_6329);
or U9231 (N_9231,N_7192,N_6991);
or U9232 (N_9232,N_7827,N_7453);
nor U9233 (N_9233,N_6643,N_6385);
nand U9234 (N_9234,N_7784,N_7834);
or U9235 (N_9235,N_6855,N_8240);
or U9236 (N_9236,N_7714,N_8076);
nor U9237 (N_9237,N_6687,N_6750);
nor U9238 (N_9238,N_8583,N_6892);
or U9239 (N_9239,N_8234,N_7161);
nor U9240 (N_9240,N_6860,N_7694);
and U9241 (N_9241,N_8389,N_6593);
or U9242 (N_9242,N_8066,N_7601);
nor U9243 (N_9243,N_8510,N_6940);
or U9244 (N_9244,N_8457,N_7469);
or U9245 (N_9245,N_8108,N_8768);
and U9246 (N_9246,N_6240,N_7993);
and U9247 (N_9247,N_8883,N_6377);
nor U9248 (N_9248,N_7117,N_8284);
nand U9249 (N_9249,N_8995,N_7716);
or U9250 (N_9250,N_7676,N_6490);
and U9251 (N_9251,N_6629,N_6264);
or U9252 (N_9252,N_7729,N_8493);
or U9253 (N_9253,N_6058,N_7168);
or U9254 (N_9254,N_7077,N_8965);
nand U9255 (N_9255,N_7011,N_7062);
nor U9256 (N_9256,N_8282,N_6604);
nor U9257 (N_9257,N_6572,N_8725);
and U9258 (N_9258,N_8320,N_7198);
and U9259 (N_9259,N_8466,N_6282);
and U9260 (N_9260,N_8804,N_7484);
nand U9261 (N_9261,N_8257,N_6048);
nor U9262 (N_9262,N_6772,N_6366);
nand U9263 (N_9263,N_7859,N_8502);
nor U9264 (N_9264,N_8653,N_7738);
nand U9265 (N_9265,N_7585,N_8665);
or U9266 (N_9266,N_6039,N_7391);
nor U9267 (N_9267,N_8417,N_7575);
nor U9268 (N_9268,N_6939,N_6683);
nand U9269 (N_9269,N_8642,N_8926);
xor U9270 (N_9270,N_7517,N_6866);
nand U9271 (N_9271,N_7530,N_8844);
nor U9272 (N_9272,N_8238,N_7422);
and U9273 (N_9273,N_6273,N_8193);
or U9274 (N_9274,N_8169,N_8026);
nor U9275 (N_9275,N_8156,N_8740);
nor U9276 (N_9276,N_6266,N_6098);
nand U9277 (N_9277,N_8181,N_8842);
nor U9278 (N_9278,N_6429,N_7366);
or U9279 (N_9279,N_7807,N_7071);
and U9280 (N_9280,N_8826,N_7477);
or U9281 (N_9281,N_6150,N_6148);
nand U9282 (N_9282,N_8945,N_7782);
nand U9283 (N_9283,N_8358,N_8274);
or U9284 (N_9284,N_8541,N_6742);
and U9285 (N_9285,N_8412,N_7173);
nand U9286 (N_9286,N_8314,N_7208);
nand U9287 (N_9287,N_7531,N_8783);
nor U9288 (N_9288,N_7488,N_7318);
and U9289 (N_9289,N_6578,N_7511);
and U9290 (N_9290,N_6698,N_8702);
or U9291 (N_9291,N_7301,N_6102);
or U9292 (N_9292,N_6569,N_8628);
nand U9293 (N_9293,N_7147,N_7856);
and U9294 (N_9294,N_8103,N_7361);
and U9295 (N_9295,N_8376,N_7543);
nand U9296 (N_9296,N_8764,N_7590);
nor U9297 (N_9297,N_6814,N_7635);
nor U9298 (N_9298,N_8400,N_7209);
nor U9299 (N_9299,N_8755,N_7218);
nand U9300 (N_9300,N_8242,N_6636);
and U9301 (N_9301,N_8917,N_8592);
or U9302 (N_9302,N_8914,N_8040);
and U9303 (N_9303,N_7822,N_8363);
and U9304 (N_9304,N_6880,N_7076);
or U9305 (N_9305,N_7600,N_7379);
and U9306 (N_9306,N_7698,N_7133);
or U9307 (N_9307,N_7829,N_7393);
nand U9308 (N_9308,N_8884,N_6630);
and U9309 (N_9309,N_6703,N_8599);
and U9310 (N_9310,N_8690,N_7290);
nand U9311 (N_9311,N_6056,N_6211);
nand U9312 (N_9312,N_8770,N_6700);
or U9313 (N_9313,N_8967,N_6356);
nor U9314 (N_9314,N_6339,N_6913);
nor U9315 (N_9315,N_6632,N_6619);
nand U9316 (N_9316,N_6405,N_8672);
and U9317 (N_9317,N_7901,N_7882);
nand U9318 (N_9318,N_7593,N_6617);
or U9319 (N_9319,N_6438,N_6189);
nand U9320 (N_9320,N_6451,N_7835);
nor U9321 (N_9321,N_8882,N_6794);
xor U9322 (N_9322,N_7229,N_8232);
xnor U9323 (N_9323,N_6980,N_7017);
or U9324 (N_9324,N_6399,N_6709);
nor U9325 (N_9325,N_8043,N_7296);
and U9326 (N_9326,N_6346,N_7654);
or U9327 (N_9327,N_6579,N_6950);
nor U9328 (N_9328,N_7028,N_8024);
nor U9329 (N_9329,N_6589,N_8073);
or U9330 (N_9330,N_7953,N_7539);
nor U9331 (N_9331,N_7874,N_6120);
nor U9332 (N_9332,N_8430,N_8267);
nor U9333 (N_9333,N_7943,N_8927);
nand U9334 (N_9334,N_8643,N_8097);
nand U9335 (N_9335,N_7727,N_7104);
nor U9336 (N_9336,N_7226,N_6086);
nand U9337 (N_9337,N_8590,N_6612);
nor U9338 (N_9338,N_6488,N_8919);
xor U9339 (N_9339,N_7111,N_7572);
nand U9340 (N_9340,N_8710,N_7146);
nor U9341 (N_9341,N_7236,N_6610);
nand U9342 (N_9342,N_7941,N_6798);
and U9343 (N_9343,N_7574,N_6956);
nor U9344 (N_9344,N_8901,N_7544);
nand U9345 (N_9345,N_7088,N_7129);
xnor U9346 (N_9346,N_8161,N_8067);
nand U9347 (N_9347,N_8937,N_7446);
nor U9348 (N_9348,N_6382,N_7425);
and U9349 (N_9349,N_7428,N_7847);
nand U9350 (N_9350,N_7702,N_7139);
nor U9351 (N_9351,N_6450,N_6368);
or U9352 (N_9352,N_7204,N_8113);
or U9353 (N_9353,N_8211,N_6771);
and U9354 (N_9354,N_6536,N_7308);
nor U9355 (N_9355,N_8731,N_6998);
or U9356 (N_9356,N_8070,N_8860);
nand U9357 (N_9357,N_8145,N_7474);
nor U9358 (N_9358,N_7090,N_6649);
and U9359 (N_9359,N_7044,N_8411);
or U9360 (N_9360,N_7341,N_8546);
nand U9361 (N_9361,N_8527,N_7270);
or U9362 (N_9362,N_6199,N_6660);
nor U9363 (N_9363,N_8253,N_7808);
or U9364 (N_9364,N_6853,N_7696);
and U9365 (N_9365,N_7051,N_6762);
or U9366 (N_9366,N_8610,N_6246);
or U9367 (N_9367,N_7787,N_7668);
or U9368 (N_9368,N_8155,N_7426);
or U9369 (N_9369,N_8164,N_6898);
nand U9370 (N_9370,N_6901,N_8994);
or U9371 (N_9371,N_6646,N_7141);
nand U9372 (N_9372,N_8688,N_6885);
nor U9373 (N_9373,N_7981,N_8098);
nand U9374 (N_9374,N_8283,N_8342);
or U9375 (N_9375,N_7343,N_8935);
nand U9376 (N_9376,N_7115,N_6081);
or U9377 (N_9377,N_6258,N_8387);
nor U9378 (N_9378,N_6252,N_7929);
or U9379 (N_9379,N_7178,N_8741);
nor U9380 (N_9380,N_8292,N_7040);
and U9381 (N_9381,N_6124,N_8126);
nand U9382 (N_9382,N_7744,N_7286);
or U9383 (N_9383,N_6477,N_8479);
and U9384 (N_9384,N_7470,N_6952);
and U9385 (N_9385,N_6419,N_8092);
nand U9386 (N_9386,N_8504,N_7969);
nand U9387 (N_9387,N_6126,N_6247);
nand U9388 (N_9388,N_7871,N_6214);
nor U9389 (N_9389,N_8135,N_8132);
nand U9390 (N_9390,N_6753,N_7687);
and U9391 (N_9391,N_7621,N_7438);
or U9392 (N_9392,N_6492,N_7235);
or U9393 (N_9393,N_7080,N_6336);
nor U9394 (N_9394,N_8371,N_7433);
nand U9395 (N_9395,N_6789,N_8396);
and U9396 (N_9396,N_8760,N_6108);
or U9397 (N_9397,N_6178,N_6975);
or U9398 (N_9398,N_8236,N_6149);
nor U9399 (N_9399,N_8484,N_7340);
or U9400 (N_9400,N_7331,N_8046);
nor U9401 (N_9401,N_7345,N_8575);
or U9402 (N_9402,N_6309,N_8654);
and U9403 (N_9403,N_8891,N_7007);
or U9404 (N_9404,N_6634,N_7804);
nor U9405 (N_9405,N_6347,N_8681);
or U9406 (N_9406,N_8202,N_8617);
nor U9407 (N_9407,N_7082,N_7965);
nor U9408 (N_9408,N_6290,N_7295);
or U9409 (N_9409,N_8037,N_7302);
and U9410 (N_9410,N_6095,N_8647);
nor U9411 (N_9411,N_6895,N_6425);
nor U9412 (N_9412,N_7862,N_7891);
nor U9413 (N_9413,N_8170,N_8398);
nor U9414 (N_9414,N_6760,N_7690);
nor U9415 (N_9415,N_6168,N_8140);
or U9416 (N_9416,N_6838,N_6401);
nor U9417 (N_9417,N_7906,N_6245);
nand U9418 (N_9418,N_7897,N_8295);
or U9419 (N_9419,N_7948,N_8134);
nor U9420 (N_9420,N_7371,N_7697);
or U9421 (N_9421,N_8191,N_7441);
and U9422 (N_9422,N_6645,N_8491);
and U9423 (N_9423,N_7840,N_8795);
nand U9424 (N_9424,N_7170,N_7321);
and U9425 (N_9425,N_7316,N_8154);
nor U9426 (N_9426,N_8852,N_8027);
nand U9427 (N_9427,N_7942,N_7105);
and U9428 (N_9428,N_8706,N_6743);
and U9429 (N_9429,N_8805,N_7754);
or U9430 (N_9430,N_7768,N_7277);
nand U9431 (N_9431,N_6025,N_8861);
nand U9432 (N_9432,N_7476,N_6766);
nand U9433 (N_9433,N_7546,N_7093);
nor U9434 (N_9434,N_7478,N_6911);
and U9435 (N_9435,N_7102,N_8679);
or U9436 (N_9436,N_7994,N_8958);
xnor U9437 (N_9437,N_7860,N_8399);
and U9438 (N_9438,N_6902,N_7486);
or U9439 (N_9439,N_6816,N_7573);
nor U9440 (N_9440,N_6662,N_6472);
or U9441 (N_9441,N_8099,N_6034);
or U9442 (N_9442,N_8986,N_7239);
nor U9443 (N_9443,N_8199,N_8925);
and U9444 (N_9444,N_6588,N_6325);
xnor U9445 (N_9445,N_8498,N_6411);
and U9446 (N_9446,N_8656,N_6667);
nor U9447 (N_9447,N_8499,N_8765);
and U9448 (N_9448,N_6713,N_6935);
nand U9449 (N_9449,N_8118,N_6690);
nor U9450 (N_9450,N_6153,N_8876);
and U9451 (N_9451,N_6644,N_8269);
nand U9452 (N_9452,N_8285,N_7527);
or U9453 (N_9453,N_7513,N_8359);
nand U9454 (N_9454,N_6575,N_8719);
and U9455 (N_9455,N_7403,N_7973);
nor U9456 (N_9456,N_8437,N_8748);
xor U9457 (N_9457,N_6847,N_7746);
nand U9458 (N_9458,N_8345,N_7786);
and U9459 (N_9459,N_7620,N_8503);
and U9460 (N_9460,N_8823,N_7597);
and U9461 (N_9461,N_8421,N_7018);
and U9462 (N_9462,N_7073,N_8893);
nand U9463 (N_9463,N_7227,N_7269);
or U9464 (N_9464,N_7869,N_6278);
nor U9465 (N_9465,N_6978,N_8188);
and U9466 (N_9466,N_8472,N_8668);
nand U9467 (N_9467,N_8375,N_7805);
and U9468 (N_9468,N_6616,N_7074);
or U9469 (N_9469,N_7963,N_6655);
and U9470 (N_9470,N_6613,N_7547);
nor U9471 (N_9471,N_8897,N_7230);
nand U9472 (N_9472,N_8262,N_7140);
nor U9473 (N_9473,N_6809,N_8367);
or U9474 (N_9474,N_7155,N_7335);
or U9475 (N_9475,N_6239,N_8956);
nand U9476 (N_9476,N_7138,N_6393);
nand U9477 (N_9477,N_6955,N_7386);
and U9478 (N_9478,N_6028,N_8746);
nor U9479 (N_9479,N_6127,N_6856);
nand U9480 (N_9480,N_7861,N_7926);
nor U9481 (N_9481,N_6193,N_6962);
nor U9482 (N_9482,N_7008,N_8619);
nor U9483 (N_9483,N_6696,N_6397);
nand U9484 (N_9484,N_8218,N_7934);
nor U9485 (N_9485,N_8789,N_6387);
or U9486 (N_9486,N_7482,N_7987);
nand U9487 (N_9487,N_7913,N_7995);
nor U9488 (N_9488,N_8793,N_6002);
or U9489 (N_9489,N_8223,N_8231);
or U9490 (N_9490,N_7626,N_8250);
nor U9491 (N_9491,N_8001,N_8381);
nand U9492 (N_9492,N_7063,N_6139);
or U9493 (N_9493,N_6989,N_8500);
or U9494 (N_9494,N_8996,N_7809);
or U9495 (N_9495,N_6922,N_7078);
nand U9496 (N_9496,N_8434,N_7519);
and U9497 (N_9497,N_6480,N_6560);
and U9498 (N_9498,N_8176,N_8386);
xor U9499 (N_9499,N_6534,N_7411);
nor U9500 (N_9500,N_6543,N_7516);
nor U9501 (N_9501,N_6681,N_6852);
nand U9502 (N_9502,N_7790,N_6352);
and U9503 (N_9503,N_6442,N_8872);
or U9504 (N_9504,N_8351,N_8185);
nand U9505 (N_9505,N_7156,N_6276);
nand U9506 (N_9506,N_8228,N_6850);
and U9507 (N_9507,N_8392,N_8057);
nor U9508 (N_9508,N_8029,N_6896);
nand U9509 (N_9509,N_6516,N_6476);
nand U9510 (N_9510,N_6749,N_8686);
nand U9511 (N_9511,N_7022,N_8743);
and U9512 (N_9512,N_7581,N_8947);
or U9513 (N_9513,N_6241,N_7456);
or U9514 (N_9514,N_7037,N_6993);
or U9515 (N_9515,N_8694,N_7659);
nand U9516 (N_9516,N_7646,N_6916);
nand U9517 (N_9517,N_7010,N_7510);
and U9518 (N_9518,N_8069,N_6196);
and U9519 (N_9519,N_7815,N_8924);
nor U9520 (N_9520,N_7503,N_8453);
nand U9521 (N_9521,N_6144,N_8331);
or U9522 (N_9522,N_6596,N_6027);
nor U9523 (N_9523,N_7256,N_6623);
nor U9524 (N_9524,N_7652,N_6573);
and U9525 (N_9525,N_7362,N_8470);
nand U9526 (N_9526,N_8666,N_8160);
nand U9527 (N_9527,N_6842,N_7024);
nand U9528 (N_9528,N_7841,N_7119);
and U9529 (N_9529,N_8286,N_7988);
nor U9530 (N_9530,N_6041,N_7592);
xnor U9531 (N_9531,N_8347,N_8296);
and U9532 (N_9532,N_7347,N_6076);
nor U9533 (N_9533,N_6759,N_6223);
and U9534 (N_9534,N_6828,N_7875);
and U9535 (N_9535,N_7359,N_6007);
nand U9536 (N_9536,N_6074,N_6887);
nand U9537 (N_9537,N_8327,N_8829);
nand U9538 (N_9538,N_6804,N_7179);
nand U9539 (N_9539,N_8189,N_8096);
or U9540 (N_9540,N_8708,N_6710);
and U9541 (N_9541,N_7413,N_6780);
nand U9542 (N_9542,N_7322,N_8254);
nand U9543 (N_9543,N_7800,N_8117);
nor U9544 (N_9544,N_8158,N_8055);
nor U9545 (N_9545,N_7002,N_6651);
nand U9546 (N_9546,N_8553,N_8125);
or U9547 (N_9547,N_6464,N_7536);
nor U9548 (N_9548,N_7644,N_7681);
nor U9549 (N_9549,N_8229,N_6267);
and U9550 (N_9550,N_7303,N_7114);
or U9551 (N_9551,N_6858,N_8508);
nand U9552 (N_9552,N_8114,N_7021);
and U9553 (N_9553,N_7169,N_7455);
nor U9554 (N_9554,N_7893,N_7672);
nor U9555 (N_9555,N_6972,N_6746);
or U9556 (N_9556,N_6071,N_7452);
nor U9557 (N_9557,N_6306,N_7991);
nand U9558 (N_9558,N_6340,N_7220);
and U9559 (N_9559,N_8890,N_6503);
nand U9560 (N_9560,N_6198,N_7392);
or U9561 (N_9561,N_6788,N_7642);
and U9562 (N_9562,N_8932,N_8350);
nand U9563 (N_9563,N_6867,N_6068);
nor U9564 (N_9564,N_8929,N_8195);
nor U9565 (N_9565,N_7655,N_6705);
nand U9566 (N_9566,N_6190,N_7436);
nor U9567 (N_9567,N_7338,N_8425);
and U9568 (N_9568,N_8121,N_7435);
or U9569 (N_9569,N_6658,N_8390);
xor U9570 (N_9570,N_8641,N_6554);
and U9571 (N_9571,N_8382,N_8810);
and U9572 (N_9572,N_8701,N_8715);
or U9573 (N_9573,N_8907,N_7016);
nor U9574 (N_9574,N_7937,N_7507);
xnor U9575 (N_9575,N_8649,N_6001);
nand U9576 (N_9576,N_8309,N_8718);
nor U9577 (N_9577,N_8179,N_7692);
or U9578 (N_9578,N_6063,N_8272);
nor U9579 (N_9579,N_8163,N_6920);
nor U9580 (N_9580,N_6281,N_7394);
nand U9581 (N_9581,N_8167,N_6402);
and U9582 (N_9582,N_6318,N_8888);
or U9583 (N_9583,N_8102,N_7916);
and U9584 (N_9584,N_7388,N_8624);
and U9585 (N_9585,N_8088,N_6625);
and U9586 (N_9586,N_8736,N_8699);
and U9587 (N_9587,N_8780,N_7225);
nor U9588 (N_9588,N_8462,N_7195);
or U9589 (N_9589,N_7118,N_7910);
nand U9590 (N_9590,N_8724,N_7113);
nor U9591 (N_9591,N_7288,N_8639);
and U9592 (N_9592,N_7757,N_7153);
nand U9593 (N_9593,N_6308,N_6602);
nand U9594 (N_9594,N_7683,N_8660);
and U9595 (N_9595,N_6790,N_6525);
or U9596 (N_9596,N_6119,N_6947);
nand U9597 (N_9597,N_7312,N_7381);
and U9598 (N_9598,N_8835,N_6664);
nor U9599 (N_9599,N_6015,N_6786);
or U9600 (N_9600,N_8082,N_7495);
or U9601 (N_9601,N_7720,N_8588);
nor U9602 (N_9602,N_6702,N_7812);
or U9603 (N_9603,N_7419,N_6471);
nand U9604 (N_9604,N_6207,N_6073);
nand U9605 (N_9605,N_6047,N_6277);
or U9606 (N_9606,N_7907,N_6383);
nand U9607 (N_9607,N_8487,N_8394);
or U9608 (N_9608,N_6269,N_7267);
and U9609 (N_9609,N_6631,N_8543);
and U9610 (N_9610,N_6529,N_6295);
nand U9611 (N_9611,N_7832,N_7903);
or U9612 (N_9612,N_6518,N_6092);
or U9613 (N_9613,N_6050,N_7693);
or U9614 (N_9614,N_7914,N_8889);
or U9615 (N_9615,N_7949,N_7412);
and U9616 (N_9616,N_6859,N_6778);
nand U9617 (N_9617,N_6800,N_7617);
xor U9618 (N_9618,N_7299,N_7203);
nand U9619 (N_9619,N_8036,N_8658);
nor U9620 (N_9620,N_8771,N_6128);
or U9621 (N_9621,N_8340,N_7013);
nand U9622 (N_9622,N_6250,N_6840);
nand U9623 (N_9623,N_6692,N_8915);
nor U9624 (N_9624,N_8565,N_8419);
nor U9625 (N_9625,N_8415,N_7712);
nand U9626 (N_9626,N_7313,N_7745);
or U9627 (N_9627,N_6087,N_7936);
nor U9628 (N_9628,N_7848,N_8815);
xnor U9629 (N_9629,N_8449,N_7776);
nor U9630 (N_9630,N_7493,N_6910);
and U9631 (N_9631,N_7721,N_6260);
nor U9632 (N_9632,N_8745,N_8168);
or U9633 (N_9633,N_6555,N_7339);
nor U9634 (N_9634,N_8635,N_7450);
nor U9635 (N_9635,N_7283,N_7125);
and U9636 (N_9636,N_6562,N_7972);
or U9637 (N_9637,N_7921,N_7996);
nand U9638 (N_9638,N_6334,N_6653);
or U9639 (N_9639,N_6155,N_8713);
or U9640 (N_9640,N_8362,N_7349);
xor U9641 (N_9641,N_7781,N_8951);
nor U9642 (N_9642,N_6526,N_7764);
nor U9643 (N_9643,N_7833,N_7320);
xor U9644 (N_9644,N_8021,N_6499);
nor U9645 (N_9645,N_7029,N_6237);
and U9646 (N_9646,N_8605,N_6869);
nand U9647 (N_9647,N_7496,N_7567);
nor U9648 (N_9648,N_7489,N_8549);
nor U9649 (N_9649,N_6821,N_7032);
or U9650 (N_9650,N_8845,N_8782);
and U9651 (N_9651,N_8791,N_6843);
nor U9652 (N_9652,N_8540,N_7079);
and U9653 (N_9653,N_7502,N_7990);
or U9654 (N_9654,N_7911,N_6927);
and U9655 (N_9655,N_6022,N_6310);
and U9656 (N_9656,N_7548,N_8875);
nor U9657 (N_9657,N_8825,N_7326);
nand U9658 (N_9658,N_6416,N_8662);
nor U9659 (N_9659,N_6275,N_6187);
or U9660 (N_9660,N_8518,N_7813);
and U9661 (N_9661,N_7675,N_7853);
nor U9662 (N_9662,N_7769,N_7999);
nor U9663 (N_9663,N_7609,N_6958);
xor U9664 (N_9664,N_7892,N_6448);
nor U9665 (N_9665,N_7549,N_7163);
or U9666 (N_9666,N_8182,N_6865);
nand U9667 (N_9667,N_8980,N_6933);
and U9668 (N_9668,N_6112,N_7310);
nor U9669 (N_9669,N_7166,N_7615);
and U9670 (N_9670,N_7602,N_7122);
and U9671 (N_9671,N_7323,N_7070);
and U9672 (N_9672,N_7667,N_6861);
and U9673 (N_9673,N_6925,N_6205);
nor U9674 (N_9674,N_8582,N_6417);
and U9675 (N_9675,N_7662,N_6089);
nand U9676 (N_9676,N_6741,N_7206);
and U9677 (N_9677,N_8180,N_7257);
or U9678 (N_9678,N_6906,N_6272);
nand U9679 (N_9679,N_7187,N_7047);
or U9680 (N_9680,N_6592,N_6191);
nor U9681 (N_9681,N_6408,N_8241);
nand U9682 (N_9682,N_6891,N_7157);
or U9683 (N_9683,N_8391,N_8928);
or U9684 (N_9684,N_6435,N_8514);
nand U9685 (N_9685,N_8225,N_8519);
nor U9686 (N_9686,N_7108,N_8352);
nor U9687 (N_9687,N_8714,N_6298);
and U9688 (N_9688,N_7292,N_6444);
nand U9689 (N_9689,N_6396,N_7087);
nand U9690 (N_9690,N_7836,N_7713);
nand U9691 (N_9691,N_7485,N_8733);
nand U9692 (N_9692,N_6576,N_6475);
nand U9693 (N_9693,N_8197,N_6194);
nor U9694 (N_9694,N_7726,N_6685);
nand U9695 (N_9695,N_7054,N_7684);
nor U9696 (N_9696,N_7618,N_6052);
and U9697 (N_9697,N_8955,N_7065);
nor U9698 (N_9698,N_7791,N_6285);
nand U9699 (N_9699,N_8942,N_8011);
or U9700 (N_9700,N_8261,N_6301);
nor U9701 (N_9701,N_8100,N_8186);
nor U9702 (N_9702,N_8408,N_8464);
and U9703 (N_9703,N_8233,N_7107);
and U9704 (N_9704,N_8049,N_6287);
nor U9705 (N_9705,N_8934,N_7404);
or U9706 (N_9706,N_8700,N_7067);
or U9707 (N_9707,N_7291,N_6341);
nand U9708 (N_9708,N_6583,N_6908);
or U9709 (N_9709,N_7278,N_6491);
or U9710 (N_9710,N_7137,N_6894);
nor U9711 (N_9711,N_7894,N_8330);
and U9712 (N_9712,N_7459,N_7959);
xor U9713 (N_9713,N_7445,N_7221);
nand U9714 (N_9714,N_8224,N_8611);
or U9715 (N_9715,N_8012,N_8212);
and U9716 (N_9716,N_7038,N_7607);
nor U9717 (N_9717,N_6179,N_7535);
or U9718 (N_9718,N_8501,N_7424);
nand U9719 (N_9719,N_8315,N_6767);
and U9720 (N_9720,N_8217,N_6215);
nor U9721 (N_9721,N_6066,N_8485);
nand U9722 (N_9722,N_8830,N_8157);
and U9723 (N_9723,N_7880,N_7380);
nand U9724 (N_9724,N_6594,N_8072);
or U9725 (N_9725,N_8307,N_7075);
and U9726 (N_9726,N_8042,N_7872);
nor U9727 (N_9727,N_8020,N_7244);
and U9728 (N_9728,N_6792,N_7748);
nor U9729 (N_9729,N_6621,N_7515);
nand U9730 (N_9730,N_8171,N_8458);
nor U9731 (N_9731,N_8397,N_7199);
nor U9732 (N_9732,N_6082,N_7238);
nor U9733 (N_9733,N_6167,N_8865);
or U9734 (N_9734,N_8239,N_6558);
nand U9735 (N_9735,N_8303,N_6351);
nor U9736 (N_9736,N_6835,N_8809);
nand U9737 (N_9737,N_6145,N_6517);
nand U9738 (N_9738,N_8207,N_8561);
xor U9739 (N_9739,N_6125,N_8294);
xor U9740 (N_9740,N_6977,N_7706);
nand U9741 (N_9741,N_8366,N_7172);
and U9742 (N_9742,N_6003,N_6521);
or U9743 (N_9743,N_7556,N_8521);
or U9744 (N_9744,N_6608,N_6083);
or U9745 (N_9745,N_6542,N_7015);
nor U9746 (N_9746,N_8459,N_8123);
nand U9747 (N_9747,N_6831,N_7327);
nor U9748 (N_9748,N_6359,N_8335);
or U9749 (N_9749,N_6111,N_8697);
and U9750 (N_9750,N_7246,N_6354);
and U9751 (N_9751,N_6443,N_6017);
and U9752 (N_9752,N_7541,N_6380);
nor U9753 (N_9753,N_6751,N_6917);
or U9754 (N_9754,N_8936,N_6953);
or U9755 (N_9755,N_7779,N_8646);
and U9756 (N_9756,N_8535,N_8878);
or U9757 (N_9757,N_7191,N_7509);
nand U9758 (N_9758,N_7159,N_8969);
and U9759 (N_9759,N_8489,N_8563);
nand U9760 (N_9760,N_7160,N_8584);
or U9761 (N_9761,N_6360,N_8216);
or U9762 (N_9762,N_8742,N_8280);
nor U9763 (N_9763,N_7035,N_7974);
xnor U9764 (N_9764,N_6020,N_7839);
nand U9765 (N_9765,N_8981,N_7545);
and U9766 (N_9766,N_7957,N_7843);
or U9767 (N_9767,N_8270,N_7068);
nand U9768 (N_9768,N_8273,N_8505);
or U9769 (N_9769,N_7979,N_7751);
nor U9770 (N_9770,N_8348,N_8165);
nand U9771 (N_9771,N_7205,N_7439);
nor U9772 (N_9772,N_6496,N_8520);
or U9773 (N_9773,N_8259,N_6889);
nand U9774 (N_9774,N_6757,N_7370);
or U9775 (N_9775,N_7614,N_7622);
and U9776 (N_9776,N_7057,N_6611);
nand U9777 (N_9777,N_7870,N_7578);
nor U9778 (N_9778,N_7604,N_6055);
nor U9779 (N_9779,N_8370,N_8978);
and U9780 (N_9780,N_8166,N_8931);
or U9781 (N_9781,N_8545,N_8817);
or U9782 (N_9782,N_6274,N_6487);
and U9783 (N_9783,N_7752,N_6836);
nand U9784 (N_9784,N_8579,N_7175);
or U9785 (N_9785,N_6507,N_7912);
nor U9786 (N_9786,N_6391,N_7215);
or U9787 (N_9787,N_7211,N_7631);
nor U9788 (N_9788,N_8047,N_7228);
and U9789 (N_9789,N_8856,N_6820);
and U9790 (N_9790,N_6370,N_7785);
or U9791 (N_9791,N_6964,N_8094);
nor U9792 (N_9792,N_8669,N_7263);
xor U9793 (N_9793,N_8762,N_7686);
nand U9794 (N_9794,N_7020,N_6745);
nand U9795 (N_9795,N_7562,N_7043);
nand U9796 (N_9796,N_6633,N_8143);
nor U9797 (N_9797,N_6262,N_6184);
or U9798 (N_9798,N_7660,N_6216);
and U9799 (N_9799,N_6470,N_8551);
nand U9800 (N_9800,N_7733,N_6728);
nand U9801 (N_9801,N_6514,N_7793);
nand U9802 (N_9802,N_8023,N_7873);
nand U9803 (N_9803,N_6023,N_8766);
nor U9804 (N_9804,N_8444,N_6659);
nand U9805 (N_9805,N_8077,N_7925);
or U9806 (N_9806,N_8263,N_7465);
or U9807 (N_9807,N_8208,N_6430);
and U9808 (N_9808,N_6202,N_8032);
or U9809 (N_9809,N_8326,N_7639);
nor U9810 (N_9810,N_6317,N_6783);
and U9811 (N_9811,N_7603,N_8058);
and U9812 (N_9812,N_7480,N_7778);
or U9813 (N_9813,N_7128,N_6265);
nor U9814 (N_9814,N_6338,N_7534);
and U9815 (N_9815,N_8028,N_6181);
nand U9816 (N_9816,N_8858,N_6722);
or U9817 (N_9817,N_7268,N_6486);
or U9818 (N_9818,N_8448,N_7758);
and U9819 (N_9819,N_7061,N_6157);
nor U9820 (N_9820,N_6548,N_8867);
xnor U9821 (N_9821,N_6987,N_8235);
nand U9822 (N_9822,N_6684,N_7888);
nor U9823 (N_9823,N_7336,N_8424);
nor U9824 (N_9824,N_6326,N_6494);
nor U9825 (N_9825,N_6942,N_7289);
nor U9826 (N_9826,N_8051,N_7780);
nand U9827 (N_9827,N_7265,N_8990);
or U9828 (N_9828,N_6986,N_6104);
nor U9829 (N_9829,N_7649,N_8488);
nor U9830 (N_9830,N_6642,N_8557);
and U9831 (N_9831,N_8562,N_8881);
and U9832 (N_9832,N_7739,N_7551);
and U9833 (N_9833,N_7552,N_6626);
and U9834 (N_9834,N_7704,N_8009);
and U9835 (N_9835,N_8035,N_7396);
nand U9836 (N_9836,N_6854,N_8712);
and U9837 (N_9837,N_8271,N_7149);
nand U9838 (N_9838,N_6890,N_6833);
and U9839 (N_9839,N_8482,N_7724);
and U9840 (N_9840,N_7900,N_7053);
nand U9841 (N_9841,N_8031,N_6874);
xor U9842 (N_9842,N_7324,N_7427);
xnor U9843 (N_9843,N_7276,N_8357);
nand U9844 (N_9844,N_8661,N_8671);
or U9845 (N_9845,N_6235,N_6079);
nor U9846 (N_9846,N_8895,N_7026);
or U9847 (N_9847,N_8455,N_8753);
nor U9848 (N_9848,N_7059,N_8730);
and U9849 (N_9849,N_7625,N_7971);
and U9850 (N_9850,N_8950,N_6726);
or U9851 (N_9851,N_7756,N_7311);
nor U9852 (N_9852,N_8065,N_7492);
or U9853 (N_9853,N_7741,N_6418);
nor U9854 (N_9854,N_7719,N_6754);
nand U9855 (N_9855,N_7879,N_8144);
or U9856 (N_9856,N_7648,N_6403);
nor U9857 (N_9857,N_7884,N_7964);
nor U9858 (N_9858,N_6661,N_8438);
and U9859 (N_9859,N_6785,N_6292);
nand U9860 (N_9860,N_7046,N_6032);
or U9861 (N_9861,N_7012,N_6863);
and U9862 (N_9862,N_6603,N_7423);
or U9863 (N_9863,N_7124,N_8483);
nor U9864 (N_9864,N_6903,N_6647);
nand U9865 (N_9865,N_6328,N_8738);
nor U9866 (N_9866,N_8056,N_7864);
nor U9867 (N_9867,N_6320,N_6454);
nor U9868 (N_9868,N_8629,N_6031);
and U9869 (N_9869,N_8608,N_7577);
nor U9870 (N_9870,N_6957,N_8150);
or U9871 (N_9871,N_8473,N_7763);
nand U9872 (N_9872,N_8476,N_6345);
nand U9873 (N_9873,N_6152,N_8534);
nand U9874 (N_9874,N_7650,N_8761);
and U9875 (N_9875,N_8323,N_7240);
or U9876 (N_9876,N_7589,N_7182);
and U9877 (N_9877,N_6818,N_6160);
xor U9878 (N_9878,N_7201,N_6100);
and U9879 (N_9879,N_8496,N_8757);
and U9880 (N_9880,N_6004,N_6302);
nor U9881 (N_9881,N_6966,N_8529);
and U9882 (N_9882,N_6769,N_8604);
xor U9883 (N_9883,N_8664,N_6231);
nand U9884 (N_9884,N_7148,N_6099);
nand U9885 (N_9885,N_8807,N_8851);
nor U9886 (N_9886,N_8552,N_7333);
nand U9887 (N_9887,N_7789,N_8989);
and U9888 (N_9888,N_7945,N_6313);
xnor U9889 (N_9889,N_6808,N_6929);
nor U9890 (N_9890,N_6465,N_6924);
nand U9891 (N_9891,N_6580,N_7594);
and U9892 (N_9892,N_6042,N_6883);
nand U9893 (N_9893,N_7825,N_6671);
and U9894 (N_9894,N_7479,N_8405);
nand U9895 (N_9895,N_8033,N_6259);
nand U9896 (N_9896,N_6176,N_8801);
nand U9897 (N_9897,N_6452,N_6764);
or U9898 (N_9898,N_8754,N_7304);
nand U9899 (N_9899,N_8068,N_7760);
and U9900 (N_9900,N_7003,N_8976);
nand U9901 (N_9901,N_8474,N_6815);
nor U9902 (N_9902,N_8799,N_8627);
nor U9903 (N_9903,N_6666,N_6331);
or U9904 (N_9904,N_8219,N_8887);
or U9905 (N_9905,N_8632,N_8877);
nor U9906 (N_9906,N_8308,N_8866);
nand U9907 (N_9907,N_6538,N_6395);
or U9908 (N_9908,N_8147,N_6571);
or U9909 (N_9909,N_7508,N_7927);
or U9910 (N_9910,N_7728,N_7890);
and U9911 (N_9911,N_6510,N_6420);
and U9912 (N_9912,N_8456,N_6672);
and U9913 (N_9913,N_6409,N_8533);
nor U9914 (N_9914,N_8281,N_6639);
or U9915 (N_9915,N_7255,N_6727);
nand U9916 (N_9916,N_8137,N_6441);
nor U9917 (N_9917,N_7036,N_7197);
or U9918 (N_9918,N_6565,N_6400);
or U9919 (N_9919,N_6044,N_6016);
and U9920 (N_9920,N_7264,N_6312);
nand U9921 (N_9921,N_8109,N_6497);
or U9922 (N_9922,N_8532,N_7641);
xnor U9923 (N_9923,N_8404,N_6776);
or U9924 (N_9924,N_6300,N_6221);
nand U9925 (N_9925,N_8703,N_8578);
nor U9926 (N_9926,N_6090,N_8625);
or U9927 (N_9927,N_7224,N_8200);
nor U9928 (N_9928,N_8721,N_7550);
nor U9929 (N_9929,N_6706,N_6289);
nor U9930 (N_9930,N_7599,N_6721);
nor U9931 (N_9931,N_8093,N_8346);
and U9932 (N_9932,N_7116,N_6217);
nand U9933 (N_9933,N_8726,N_6946);
or U9934 (N_9934,N_6154,N_6286);
nand U9935 (N_9935,N_6567,N_6195);
or U9936 (N_9936,N_6426,N_6718);
xor U9937 (N_9937,N_7770,N_7399);
and U9938 (N_9938,N_7242,N_6166);
and U9939 (N_9939,N_6131,N_7464);
and U9940 (N_9940,N_6981,N_8343);
and U9941 (N_9941,N_6143,N_6954);
or U9942 (N_9942,N_8744,N_6348);
and U9943 (N_9943,N_8441,N_6992);
or U9944 (N_9944,N_6389,N_6219);
or U9945 (N_9945,N_7583,N_7777);
and U9946 (N_9946,N_6141,N_7935);
xnor U9947 (N_9947,N_7703,N_7850);
or U9948 (N_9948,N_8091,N_6365);
or U9949 (N_9949,N_8833,N_8107);
nor U9950 (N_9950,N_8899,N_8920);
nand U9951 (N_9951,N_6014,N_8567);
or U9952 (N_9952,N_8550,N_8378);
nand U9953 (N_9953,N_6872,N_8383);
nand U9954 (N_9954,N_8626,N_6468);
and U9955 (N_9955,N_6415,N_6156);
nor U9956 (N_9956,N_7444,N_7084);
and U9957 (N_9957,N_8000,N_8313);
or U9958 (N_9958,N_8673,N_8513);
nor U9959 (N_9959,N_8431,N_8827);
nor U9960 (N_9960,N_7055,N_8311);
or U9961 (N_9961,N_7685,N_7886);
xor U9962 (N_9962,N_7432,N_7252);
nor U9963 (N_9963,N_8962,N_8293);
or U9964 (N_9964,N_7091,N_6574);
nand U9965 (N_9965,N_7828,N_7796);
nand U9966 (N_9966,N_6735,N_7337);
and U9967 (N_9967,N_7490,N_6697);
nor U9968 (N_9968,N_8214,N_7243);
nand U9969 (N_9969,N_6566,N_7632);
and U9970 (N_9970,N_7374,N_6037);
and U9971 (N_9971,N_8277,N_6009);
nand U9972 (N_9972,N_7332,N_8074);
or U9973 (N_9973,N_7783,N_8244);
and U9974 (N_9974,N_8316,N_6263);
or U9975 (N_9975,N_6676,N_8676);
nor U9976 (N_9976,N_6988,N_6515);
and U9977 (N_9977,N_7151,N_8175);
nand U9978 (N_9978,N_8213,N_7461);
nand U9979 (N_9979,N_6012,N_6133);
nor U9980 (N_9980,N_8993,N_6584);
or U9981 (N_9981,N_6585,N_8301);
nor U9982 (N_9982,N_8685,N_7154);
xnor U9983 (N_9983,N_7608,N_6707);
nor U9984 (N_9984,N_7637,N_6694);
nor U9985 (N_9985,N_7367,N_8321);
or U9986 (N_9986,N_7831,N_7171);
or U9987 (N_9987,N_6489,N_6983);
and U9988 (N_9988,N_8869,N_6876);
nor U9989 (N_9989,N_8190,N_6914);
nor U9990 (N_9990,N_7498,N_8910);
nand U9991 (N_9991,N_6549,N_8364);
nand U9992 (N_9992,N_7819,N_8422);
or U9993 (N_9993,N_7930,N_7097);
nor U9994 (N_9994,N_7968,N_7254);
nor U9995 (N_9995,N_8333,N_7799);
nor U9996 (N_9996,N_6053,N_8716);
nand U9997 (N_9997,N_6638,N_6182);
nand U9998 (N_9998,N_8615,N_6018);
or U9999 (N_9999,N_6595,N_7899);
or U10000 (N_10000,N_8784,N_8758);
or U10001 (N_10001,N_8811,N_8008);
nand U10002 (N_10002,N_7300,N_7961);
nand U10003 (N_10003,N_6620,N_7919);
nor U10004 (N_10004,N_8278,N_7457);
or U10005 (N_10005,N_8813,N_6294);
nand U10006 (N_10006,N_6206,N_8515);
or U10007 (N_10007,N_7669,N_7788);
nor U10008 (N_10008,N_6019,N_6088);
nand U10009 (N_10009,N_8325,N_7985);
or U10010 (N_10010,N_6376,N_8300);
nand U10011 (N_10011,N_8905,N_8674);
nor U10012 (N_10012,N_8354,N_6161);
and U10013 (N_10013,N_7342,N_6725);
and U10014 (N_10014,N_8528,N_7280);
nand U10015 (N_10015,N_8414,N_8683);
nand U10016 (N_10016,N_8837,N_6845);
xor U10017 (N_10017,N_8318,N_8922);
and U10018 (N_10018,N_6839,N_8420);
nor U10019 (N_10019,N_6982,N_8445);
nor U10020 (N_10020,N_7569,N_7127);
and U10021 (N_10021,N_7858,N_6271);
and U10022 (N_10022,N_7250,N_7647);
or U10023 (N_10023,N_7472,N_6765);
nor U10024 (N_10024,N_6140,N_8769);
and U10025 (N_10025,N_8564,N_6976);
and U10026 (N_10026,N_7854,N_6482);
nand U10027 (N_10027,N_6434,N_7628);
or U10028 (N_10028,N_6457,N_8756);
nor U10029 (N_10029,N_6590,N_8494);
and U10030 (N_10030,N_6824,N_7245);
or U10031 (N_10031,N_7885,N_8237);
or U10032 (N_10032,N_6469,N_8747);
xnor U10033 (N_10033,N_7557,N_7512);
nand U10034 (N_10034,N_7081,N_8110);
nor U10035 (N_10035,N_6926,N_7390);
or U10036 (N_10036,N_6072,N_7866);
or U10037 (N_10037,N_6581,N_8384);
nor U10038 (N_10038,N_6116,N_6627);
nand U10039 (N_10039,N_6142,N_8332);
nand U10040 (N_10040,N_6407,N_8602);
and U10041 (N_10041,N_7742,N_8538);
or U10042 (N_10042,N_6316,N_8480);
and U10043 (N_10043,N_7915,N_6846);
and U10044 (N_10044,N_8862,N_7876);
and U10045 (N_10045,N_6985,N_6775);
nand U10046 (N_10046,N_8083,N_8062);
nor U10047 (N_10047,N_7674,N_7294);
nor U10048 (N_10048,N_8918,N_6094);
or U10049 (N_10049,N_7830,N_8836);
or U10050 (N_10050,N_8987,N_6485);
and U10051 (N_10051,N_7164,N_8775);
or U10052 (N_10052,N_7740,N_6531);
and U10053 (N_10053,N_8614,N_6284);
or U10054 (N_10054,N_8317,N_8739);
nand U10055 (N_10055,N_6810,N_7810);
nand U10056 (N_10056,N_6670,N_7285);
and U10057 (N_10057,N_6825,N_7258);
or U10058 (N_10058,N_8061,N_6628);
or U10059 (N_10059,N_6648,N_7298);
or U10060 (N_10060,N_8693,N_7126);
nand U10061 (N_10061,N_8820,N_8374);
nor U10062 (N_10062,N_7473,N_7219);
or U10063 (N_10063,N_8005,N_6251);
nor U10064 (N_10064,N_7373,N_8982);
nand U10065 (N_10065,N_8289,N_6944);
or U10066 (N_10066,N_6114,N_8734);
nor U10067 (N_10067,N_6242,N_6381);
and U10068 (N_10068,N_8663,N_7006);
or U10069 (N_10069,N_8885,N_7924);
or U10070 (N_10070,N_7529,N_7792);
and U10071 (N_10071,N_8735,N_7217);
nor U10072 (N_10072,N_8709,N_6008);
nand U10073 (N_10073,N_8794,N_6723);
nor U10074 (N_10074,N_7023,N_6695);
nand U10075 (N_10075,N_7420,N_6806);
or U10076 (N_10076,N_7417,N_8486);
nor U10077 (N_10077,N_8174,N_8451);
or U10078 (N_10078,N_7801,N_7826);
or U10079 (N_10079,N_7434,N_7431);
nand U10080 (N_10080,N_7629,N_8204);
nand U10081 (N_10081,N_6421,N_6996);
nor U10082 (N_10082,N_6678,N_8436);
or U10083 (N_10083,N_8847,N_6036);
xor U10084 (N_10084,N_7085,N_6803);
and U10085 (N_10085,N_8997,N_8081);
xnor U10086 (N_10086,N_6656,N_7939);
nor U10087 (N_10087,N_6787,N_6293);
and U10088 (N_10088,N_8463,N_6570);
nor U10089 (N_10089,N_6462,N_8355);
nor U10090 (N_10090,N_8379,N_7656);
and U10091 (N_10091,N_7189,N_6948);
and U10092 (N_10092,N_6225,N_6135);
and U10093 (N_10093,N_6101,N_8577);
and U10094 (N_10094,N_8298,N_8720);
nor U10095 (N_10095,N_8492,N_6446);
nand U10096 (N_10096,N_7058,N_8215);
or U10097 (N_10097,N_6236,N_7384);
nor U10098 (N_10098,N_8622,N_7487);
or U10099 (N_10099,N_6640,N_6511);
nor U10100 (N_10100,N_6474,N_8247);
nor U10101 (N_10101,N_6974,N_8921);
nor U10102 (N_10102,N_8044,N_6288);
nor U10103 (N_10103,N_6030,N_6739);
or U10104 (N_10104,N_6563,N_6805);
nor U10105 (N_10105,N_7904,N_8695);
nor U10106 (N_10106,N_6777,N_6909);
or U10107 (N_10107,N_7753,N_6005);
nor U10108 (N_10108,N_6714,N_6493);
nand U10109 (N_10109,N_6708,N_6704);
nand U10110 (N_10110,N_6297,N_8675);
or U10111 (N_10111,N_8085,N_8593);
xor U10112 (N_10112,N_6597,N_8041);
nor U10113 (N_10113,N_8576,N_6663);
or U10114 (N_10114,N_8112,N_6106);
or U10115 (N_10115,N_6577,N_8555);
and U10116 (N_10116,N_7395,N_6748);
nor U10117 (N_10117,N_8570,N_7658);
nor U10118 (N_10118,N_8908,N_8433);
nor U10119 (N_10119,N_6059,N_7896);
and U10120 (N_10120,N_7120,N_6871);
or U10121 (N_10121,N_8440,N_8874);
nor U10122 (N_10122,N_6879,N_6105);
and U10123 (N_10123,N_7121,N_7816);
or U10124 (N_10124,N_8759,N_7905);
nand U10125 (N_10125,N_7723,N_8933);
nand U10126 (N_10126,N_8324,N_6568);
nor U10127 (N_10127,N_7176,N_7579);
nand U10128 (N_10128,N_7202,N_8790);
or U10129 (N_10129,N_6163,N_7677);
nand U10130 (N_10130,N_7273,N_7358);
or U10131 (N_10131,N_8038,N_8843);
and U10132 (N_10132,N_8903,N_8245);
nand U10133 (N_10133,N_8991,N_8469);
nor U10134 (N_10134,N_7385,N_7443);
or U10135 (N_10135,N_7772,N_7354);
or U10136 (N_10136,N_6844,N_8256);
or U10137 (N_10137,N_6587,N_8302);
or U10138 (N_10138,N_7663,N_8460);
nor U10139 (N_10139,N_6545,N_7382);
nand U10140 (N_10140,N_6797,N_7520);
or U10141 (N_10141,N_8173,N_8524);
nor U10142 (N_10142,N_8443,N_7881);
and U10143 (N_10143,N_8630,N_6463);
nor U10144 (N_10144,N_8159,N_6768);
or U10145 (N_10145,N_8264,N_8960);
and U10146 (N_10146,N_7368,N_6618);
nand U10147 (N_10147,N_7918,N_6949);
nor U10148 (N_10148,N_7253,N_8050);
nor U10149 (N_10149,N_8016,N_8863);
and U10150 (N_10150,N_8401,N_8205);
and U10151 (N_10151,N_7766,N_6315);
nor U10152 (N_10152,N_7598,N_6046);
nor U10153 (N_10153,N_7363,N_8819);
nor U10154 (N_10154,N_6829,N_8101);
and U10155 (N_10155,N_7152,N_8848);
xor U10156 (N_10156,N_6010,N_8481);
or U10157 (N_10157,N_8187,N_8525);
or U10158 (N_10158,N_7454,N_6959);
nor U10159 (N_10159,N_7802,N_7954);
and U10160 (N_10160,N_7989,N_6024);
or U10161 (N_10161,N_6900,N_8192);
and U10162 (N_10162,N_7518,N_6064);
nand U10163 (N_10163,N_6758,N_8846);
nor U10164 (N_10164,N_6997,N_6712);
or U10165 (N_10165,N_6862,N_6244);
or U10166 (N_10166,N_7369,N_6188);
nand U10167 (N_10167,N_7234,N_8053);
and U10168 (N_10168,N_7052,N_7889);
or U10169 (N_10169,N_7587,N_7845);
nand U10170 (N_10170,N_8305,N_7823);
or U10171 (N_10171,N_6371,N_8595);
and U10172 (N_10172,N_6756,N_6138);
and U10173 (N_10173,N_6979,N_7633);
nor U10174 (N_10174,N_6372,N_8007);
nand U10175 (N_10175,N_7045,N_7795);
nand U10176 (N_10176,N_8010,N_7375);
nor U10177 (N_10177,N_8571,N_7571);
nor U10178 (N_10178,N_6732,N_6556);
nor U10179 (N_10179,N_6984,N_7130);
nor U10180 (N_10180,N_7565,N_7998);
and U10181 (N_10181,N_8620,N_6937);
and U10182 (N_10182,N_6533,N_6973);
and U10183 (N_10183,N_7177,N_6186);
nand U10184 (N_10184,N_8539,N_6173);
nand U10185 (N_10185,N_6544,N_7271);
and U10186 (N_10186,N_8116,N_8821);
and U10187 (N_10187,N_7064,N_6599);
nand U10188 (N_10188,N_7588,N_8655);
nand U10189 (N_10189,N_7701,N_8923);
nand U10190 (N_10190,N_6795,N_7098);
nand U10191 (N_10191,N_6051,N_6410);
nor U10192 (N_10192,N_7525,N_8006);
and U10193 (N_10193,N_8507,N_6774);
nand U10194 (N_10194,N_6827,N_7532);
and U10195 (N_10195,N_6103,N_8478);
nand U10196 (N_10196,N_7134,N_7610);
nor U10197 (N_10197,N_6969,N_6527);
or U10198 (N_10198,N_6422,N_8587);
nor U10199 (N_10199,N_7475,N_8573);
nor U10200 (N_10200,N_8260,N_7611);
nor U10201 (N_10201,N_8249,N_7376);
and U10202 (N_10202,N_6384,N_8426);
and U10203 (N_10203,N_7279,N_8871);
or U10204 (N_10204,N_7570,N_6201);
nand U10205 (N_10205,N_8266,N_6324);
nand U10206 (N_10206,N_7966,N_7251);
nand U10207 (N_10207,N_7749,N_7136);
and U10208 (N_10208,N_8651,N_6505);
xor U10209 (N_10209,N_6650,N_6307);
or U10210 (N_10210,N_7962,N_7307);
nand U10211 (N_10211,N_6006,N_7775);
and U10212 (N_10212,N_7041,N_7491);
xnor U10213 (N_10213,N_7619,N_8178);
nor U10214 (N_10214,N_8022,N_7700);
nand U10215 (N_10215,N_7346,N_6668);
nor U10216 (N_10216,N_7522,N_8786);
nor U10217 (N_10217,N_7731,N_6928);
xor U10218 (N_10218,N_8601,N_7983);
and U10219 (N_10219,N_8572,N_8892);
nor U10220 (N_10220,N_7895,N_7606);
or U10221 (N_10221,N_6192,N_8360);
nor U10222 (N_10222,N_7481,N_7922);
nor U10223 (N_10223,N_7096,N_8222);
nand U10224 (N_10224,N_8691,N_6204);
nand U10225 (N_10225,N_7353,N_6183);
and U10226 (N_10226,N_8276,N_7131);
or U10227 (N_10227,N_6232,N_8268);
xor U10228 (N_10228,N_7582,N_7844);
or U10229 (N_10229,N_8556,N_6060);
and U10230 (N_10230,N_6392,N_6523);
nand U10231 (N_10231,N_6185,N_6414);
nor U10232 (N_10232,N_8975,N_6561);
nand U10233 (N_10233,N_7194,N_8634);
nor U10234 (N_10234,N_8636,N_6675);
nor U10235 (N_10235,N_7842,N_8648);
nor U10236 (N_10236,N_7952,N_8003);
and U10237 (N_10237,N_7992,N_6283);
nand U10238 (N_10238,N_7867,N_6234);
nand U10239 (N_10239,N_8201,N_7185);
nor U10240 (N_10240,N_6212,N_8475);
or U10241 (N_10241,N_8385,N_6961);
or U10242 (N_10242,N_7902,N_8704);
nand U10243 (N_10243,N_7514,N_7350);
nor U10244 (N_10244,N_7806,N_7272);
or U10245 (N_10245,N_8609,N_8279);
nand U10246 (N_10246,N_7167,N_7042);
nor U10247 (N_10247,N_6394,N_8310);
nand U10248 (N_10248,N_6374,N_6546);
nor U10249 (N_10249,N_6528,N_8454);
nor U10250 (N_10250,N_6280,N_7344);
nor U10251 (N_10251,N_8677,N_7442);
xnor U10252 (N_10252,N_8251,N_8416);
or U10253 (N_10253,N_7715,N_7009);
nor U10254 (N_10254,N_8319,N_8717);
or U10255 (N_10255,N_7183,N_6230);
nor U10256 (N_10256,N_8258,N_6208);
and U10257 (N_10257,N_8071,N_6175);
nand U10258 (N_10258,N_8938,N_8687);
nor U10259 (N_10259,N_6851,N_7223);
and U10260 (N_10260,N_6963,N_7868);
nand U10261 (N_10261,N_8853,N_6013);
and U10262 (N_10262,N_8130,N_8906);
or U10263 (N_10263,N_7030,N_6943);
or U10264 (N_10264,N_6428,N_7389);
xor U10265 (N_10265,N_7638,N_6147);
and U10266 (N_10266,N_8230,N_6171);
and U10267 (N_10267,N_8329,N_7857);
xnor U10268 (N_10268,N_8220,N_6822);
nand U10269 (N_10269,N_7735,N_8151);
nor U10270 (N_10270,N_8568,N_8337);
and U10271 (N_10271,N_6918,N_6819);
and U10272 (N_10272,N_8943,N_6784);
nand U10273 (N_10273,N_6035,N_8972);
or U10274 (N_10274,N_6971,N_8030);
nor U10275 (N_10275,N_8569,N_7110);
and U10276 (N_10276,N_7725,N_6689);
and U10277 (N_10277,N_7909,N_8246);
nor U10278 (N_10278,N_7266,N_8080);
xnor U10279 (N_10279,N_7095,N_7947);
nand U10280 (N_10280,N_8353,N_6512);
and U10281 (N_10281,N_8902,N_6740);
and U10282 (N_10282,N_6951,N_8816);
or U10283 (N_10283,N_8124,N_8377);
and U10284 (N_10284,N_8894,N_7448);
nor U10285 (N_10285,N_7722,N_6553);
and U10286 (N_10286,N_6255,N_7287);
nand U10287 (N_10287,N_8900,N_8002);
and U10288 (N_10288,N_6652,N_7730);
and U10289 (N_10289,N_8560,N_6311);
and U10290 (N_10290,N_8079,N_8737);
or U10291 (N_10291,N_6731,N_8558);
or U10292 (N_10292,N_7048,N_8306);
and U10293 (N_10293,N_7817,N_8526);
and U10294 (N_10294,N_6343,N_7132);
and U10295 (N_10295,N_8087,N_7591);
nor U10296 (N_10296,N_8129,N_8751);
or U10297 (N_10297,N_7282,N_7595);
and U10298 (N_10298,N_6930,N_6970);
or U10299 (N_10299,N_6522,N_6752);
and U10300 (N_10300,N_8970,N_8954);
nor U10301 (N_10301,N_7837,N_6220);
or U10302 (N_10302,N_6357,N_6436);
nor U10303 (N_10303,N_7932,N_8089);
nor U10304 (N_10304,N_8477,N_6327);
and U10305 (N_10305,N_6801,N_6113);
and U10306 (N_10306,N_6322,N_7196);
or U10307 (N_10307,N_6605,N_8998);
and U10308 (N_10308,N_8149,N_8896);
nor U10309 (N_10309,N_7863,N_6439);
and U10310 (N_10310,N_8517,N_6504);
nor U10311 (N_10311,N_8406,N_7710);
nor U10312 (N_10312,N_7329,N_6358);
nor U10313 (N_10313,N_8105,N_6541);
and U10314 (N_10314,N_8808,N_7533);
or U10315 (N_10315,N_6826,N_6375);
nor U10316 (N_10316,N_6848,N_7222);
or U10317 (N_10317,N_8255,N_8968);
or U10318 (N_10318,N_6832,N_8973);
nand U10319 (N_10319,N_7274,N_6067);
or U10320 (N_10320,N_7103,N_6423);
or U10321 (N_10321,N_6479,N_8946);
nor U10322 (N_10322,N_8839,N_8054);
and U10323 (N_10323,N_6686,N_7773);
and U10324 (N_10324,N_7401,N_6912);
nor U10325 (N_10325,N_8450,N_6337);
nand U10326 (N_10326,N_7960,N_6586);
nor U10327 (N_10327,N_6085,N_8667);
nor U10328 (N_10328,N_6537,N_8723);
nand U10329 (N_10329,N_6878,N_6635);
or U10330 (N_10330,N_8800,N_8063);
or U10331 (N_10331,N_8141,N_6075);
nor U10332 (N_10332,N_8052,N_7811);
and U10333 (N_10333,N_8172,N_7406);
or U10334 (N_10334,N_6248,N_7537);
or U10335 (N_10335,N_8670,N_7317);
and U10336 (N_10336,N_6688,N_8698);
nand U10337 (N_10337,N_8115,N_8516);
nand U10338 (N_10338,N_7737,N_7750);
nand U10339 (N_10339,N_8781,N_7429);
nand U10340 (N_10340,N_6226,N_8018);
nand U10341 (N_10341,N_8854,N_7743);
nor U10342 (N_10342,N_7184,N_8468);
or U10343 (N_10343,N_6238,N_8547);
and U10344 (N_10344,N_7213,N_7398);
nand U10345 (N_10345,N_6817,N_6888);
nor U10346 (N_10346,N_6379,N_7671);
or U10347 (N_10347,N_7689,N_8133);
nand U10348 (N_10348,N_6406,N_6509);
or U10349 (N_10349,N_8034,N_8855);
nor U10350 (N_10350,N_6249,N_7705);
or U10351 (N_10351,N_8435,N_6174);
and U10352 (N_10352,N_7666,N_6227);
nor U10353 (N_10353,N_7898,N_7089);
and U10354 (N_10354,N_6624,N_7039);
and U10355 (N_10355,N_6932,N_8859);
xor U10356 (N_10356,N_6299,N_8961);
nor U10357 (N_10357,N_6078,N_7397);
and U10358 (N_10358,N_7330,N_7319);
nor U10359 (N_10359,N_6323,N_7505);
nand U10360 (N_10360,N_6657,N_8388);
and U10361 (N_10361,N_6622,N_7497);
nand U10362 (N_10362,N_8095,N_8979);
nor U10363 (N_10363,N_8177,N_7416);
nand U10364 (N_10364,N_6770,N_6520);
nor U10365 (N_10365,N_6530,N_8749);
nand U10366 (N_10366,N_8146,N_6333);
nand U10367 (N_10367,N_7865,N_7014);
nor U10368 (N_10368,N_6552,N_6084);
or U10369 (N_10369,N_7260,N_7365);
nand U10370 (N_10370,N_8025,N_7560);
nor U10371 (N_10371,N_6319,N_7699);
nor U10372 (N_10372,N_7462,N_6938);
nor U10373 (N_10373,N_7506,N_7005);
or U10374 (N_10374,N_6413,N_8509);
nand U10375 (N_10375,N_7314,N_6350);
nor U10376 (N_10376,N_7761,N_8039);
nand U10377 (N_10377,N_7955,N_6609);
nor U10378 (N_10378,N_6228,N_7851);
nor U10379 (N_10379,N_8631,N_7838);
nand U10380 (N_10380,N_6811,N_7680);
nor U10381 (N_10381,N_8152,N_8600);
nand U10382 (N_10382,N_6440,N_7855);
and U10383 (N_10383,N_7846,N_8773);
nand U10384 (N_10384,N_6502,N_7596);
and U10385 (N_10385,N_6054,N_8338);
nand U10386 (N_10386,N_8288,N_7232);
nor U10387 (N_10387,N_6763,N_7734);
and U10388 (N_10388,N_8880,N_8684);
nand U10389 (N_10389,N_7387,N_8637);
and U10390 (N_10390,N_6990,N_8580);
or U10391 (N_10391,N_6967,N_8429);
nor U10392 (N_10392,N_8369,N_7352);
or U10393 (N_10393,N_7200,N_6386);
or U10394 (N_10394,N_8531,N_7123);
nor U10395 (N_10395,N_6715,N_6361);
and U10396 (N_10396,N_7580,N_7355);
nor U10397 (N_10397,N_6744,N_7418);
nand U10398 (N_10398,N_8612,N_6931);
nand U10399 (N_10399,N_8104,N_6466);
nand U10400 (N_10400,N_7106,N_6802);
and U10401 (N_10401,N_7066,N_8322);
nand U10402 (N_10402,N_6218,N_6342);
and U10403 (N_10403,N_6169,N_8275);
or U10404 (N_10404,N_6353,N_7231);
and U10405 (N_10405,N_7956,N_8566);
nand U10406 (N_10406,N_8940,N_7247);
and U10407 (N_10407,N_7616,N_7060);
nand U10408 (N_10408,N_7661,N_6733);
or U10409 (N_10409,N_6693,N_8948);
nand U10410 (N_10410,N_8349,N_7521);
and U10411 (N_10411,N_6501,N_8728);
nor U10412 (N_10412,N_6253,N_7540);
and U10413 (N_10413,N_8692,N_6158);
or U10414 (N_10414,N_7524,N_6303);
and U10415 (N_10415,N_8886,N_8471);
nor U10416 (N_10416,N_8075,N_6791);
or U10417 (N_10417,N_7281,N_8803);
nand U10418 (N_10418,N_8971,N_6467);
and U10419 (N_10419,N_8128,N_7824);
or U10420 (N_10420,N_7499,N_8413);
nor U10421 (N_10421,N_8964,N_6110);
nand U10422 (N_10422,N_7284,N_8409);
or U10423 (N_10423,N_6823,N_6513);
nor U10424 (N_10424,N_6011,N_6994);
nand U10425 (N_10425,N_7364,N_8916);
and U10426 (N_10426,N_8607,N_6881);
nor U10427 (N_10427,N_8210,N_6724);
nor U10428 (N_10428,N_6123,N_6679);
nor U10429 (N_10429,N_7467,N_7261);
or U10430 (N_10430,N_7430,N_6296);
and U10431 (N_10431,N_7707,N_8633);
and U10432 (N_10432,N_6473,N_8198);
nand U10433 (N_10433,N_6398,N_8767);
xnor U10434 (N_10434,N_8497,N_8184);
nand U10435 (N_10435,N_8777,N_7975);
nor U10436 (N_10436,N_7262,N_7555);
or U10437 (N_10437,N_8336,N_7774);
nand U10438 (N_10438,N_8857,N_7640);
or U10439 (N_10439,N_7558,N_6197);
or U10440 (N_10440,N_7275,N_6919);
nor U10441 (N_10441,N_7449,N_8849);
nor U10442 (N_10442,N_7025,N_8559);
and U10443 (N_10443,N_6716,N_6736);
or U10444 (N_10444,N_8705,N_7360);
and U10445 (N_10445,N_6243,N_8585);
nand U10446 (N_10446,N_7144,N_7241);
nor U10447 (N_10447,N_8983,N_8952);
nand U10448 (N_10448,N_7984,N_8659);
and U10449 (N_10449,N_7976,N_8868);
nand U10450 (N_10450,N_6344,N_7678);
nor U10451 (N_10451,N_8465,N_8828);
or U10452 (N_10452,N_8131,N_6130);
nor U10453 (N_10453,N_7950,N_7695);
nand U10454 (N_10454,N_8014,N_7977);
and U10455 (N_10455,N_8368,N_8776);
xnor U10456 (N_10456,N_8017,N_6557);
and U10457 (N_10457,N_8873,N_8957);
nor U10458 (N_10458,N_8084,N_6500);
nand U10459 (N_10459,N_7158,N_8544);
and U10460 (N_10460,N_7069,N_8623);
nor U10461 (N_10461,N_7494,N_6233);
and U10462 (N_10462,N_7207,N_6564);
or U10463 (N_10463,N_7568,N_8119);
or U10464 (N_10464,N_7736,N_7586);
nand U10465 (N_10465,N_7297,N_7378);
nor U10466 (N_10466,N_6841,N_6261);
nand U10467 (N_10467,N_8974,N_8312);
and U10468 (N_10468,N_8122,N_7814);
and U10469 (N_10469,N_8203,N_7820);
nor U10470 (N_10470,N_8729,N_8064);
nor U10471 (N_10471,N_6431,N_6137);
and U10472 (N_10472,N_6637,N_6699);
nor U10473 (N_10473,N_7034,N_6893);
nand U10474 (N_10474,N_6449,N_6807);
and U10475 (N_10475,N_8682,N_6607);
nor U10476 (N_10476,N_8439,N_7767);
xnor U10477 (N_10477,N_7732,N_7538);
xnor U10478 (N_10478,N_6941,N_8618);
and U10479 (N_10479,N_6915,N_8984);
nand U10480 (N_10480,N_6427,N_6747);
or U10481 (N_10481,N_7056,N_8650);
and U10482 (N_10482,N_6093,N_6519);
or U10483 (N_10483,N_8341,N_8598);
nor U10484 (N_10484,N_6886,N_7765);
or U10485 (N_10485,N_6849,N_8356);
nand U10486 (N_10486,N_6029,N_6601);
nand U10487 (N_10487,N_7673,N_7627);
and U10488 (N_10488,N_6907,N_6229);
or U10489 (N_10489,N_6904,N_6270);
or U10490 (N_10490,N_7852,N_7190);
and U10491 (N_10491,N_7348,N_7877);
and U10492 (N_10492,N_6559,N_6779);
nand U10493 (N_10493,N_7471,N_6136);
nand U10494 (N_10494,N_7145,N_6390);
nor U10495 (N_10495,N_7402,N_8304);
nand U10496 (N_10496,N_6330,N_8594);
nor U10497 (N_10497,N_8221,N_7928);
nand U10498 (N_10498,N_6506,N_7447);
nor U10499 (N_10499,N_7050,N_7248);
and U10500 (N_10500,N_6786,N_6191);
or U10501 (N_10501,N_7139,N_8255);
nand U10502 (N_10502,N_7619,N_8647);
xnor U10503 (N_10503,N_6304,N_7572);
nor U10504 (N_10504,N_6328,N_8095);
nand U10505 (N_10505,N_6387,N_7348);
nor U10506 (N_10506,N_6127,N_8781);
and U10507 (N_10507,N_6557,N_7163);
and U10508 (N_10508,N_8013,N_7097);
nor U10509 (N_10509,N_6562,N_7959);
nand U10510 (N_10510,N_7911,N_8895);
and U10511 (N_10511,N_6255,N_8686);
and U10512 (N_10512,N_8183,N_8481);
and U10513 (N_10513,N_6035,N_8629);
nand U10514 (N_10514,N_6313,N_7306);
and U10515 (N_10515,N_6506,N_8124);
or U10516 (N_10516,N_8916,N_6496);
or U10517 (N_10517,N_6503,N_8224);
nor U10518 (N_10518,N_6272,N_7835);
nor U10519 (N_10519,N_7612,N_8484);
nand U10520 (N_10520,N_6341,N_6597);
nand U10521 (N_10521,N_6259,N_6546);
and U10522 (N_10522,N_6831,N_6056);
nand U10523 (N_10523,N_6904,N_6071);
and U10524 (N_10524,N_6058,N_6375);
nor U10525 (N_10525,N_8422,N_7132);
nor U10526 (N_10526,N_8101,N_6981);
or U10527 (N_10527,N_6520,N_8498);
nor U10528 (N_10528,N_8143,N_8707);
or U10529 (N_10529,N_7255,N_8093);
and U10530 (N_10530,N_8612,N_7246);
or U10531 (N_10531,N_8295,N_7309);
and U10532 (N_10532,N_6787,N_8745);
or U10533 (N_10533,N_8625,N_8688);
and U10534 (N_10534,N_7675,N_7759);
and U10535 (N_10535,N_6436,N_8749);
and U10536 (N_10536,N_7961,N_7965);
nand U10537 (N_10537,N_6369,N_7303);
and U10538 (N_10538,N_6885,N_7675);
nor U10539 (N_10539,N_7856,N_6457);
nand U10540 (N_10540,N_6365,N_6585);
nand U10541 (N_10541,N_7599,N_7969);
nor U10542 (N_10542,N_7083,N_6903);
and U10543 (N_10543,N_8725,N_6730);
nor U10544 (N_10544,N_7749,N_6868);
and U10545 (N_10545,N_8532,N_7988);
nor U10546 (N_10546,N_6725,N_6848);
nor U10547 (N_10547,N_6306,N_7667);
or U10548 (N_10548,N_7866,N_8939);
nor U10549 (N_10549,N_7783,N_8871);
and U10550 (N_10550,N_7117,N_6051);
nand U10551 (N_10551,N_6915,N_8170);
nand U10552 (N_10552,N_7606,N_6539);
and U10553 (N_10553,N_8235,N_7106);
or U10554 (N_10554,N_6757,N_8631);
nor U10555 (N_10555,N_7219,N_7158);
nand U10556 (N_10556,N_8111,N_8417);
and U10557 (N_10557,N_8686,N_7795);
xor U10558 (N_10558,N_8792,N_8053);
nand U10559 (N_10559,N_6960,N_6823);
nor U10560 (N_10560,N_7734,N_7557);
and U10561 (N_10561,N_7036,N_7703);
nand U10562 (N_10562,N_6499,N_8141);
or U10563 (N_10563,N_6488,N_6264);
and U10564 (N_10564,N_6822,N_8583);
and U10565 (N_10565,N_7767,N_7627);
and U10566 (N_10566,N_8100,N_7157);
nand U10567 (N_10567,N_6936,N_6079);
and U10568 (N_10568,N_7875,N_6735);
nand U10569 (N_10569,N_6932,N_6661);
nor U10570 (N_10570,N_8786,N_6536);
nor U10571 (N_10571,N_7207,N_8904);
and U10572 (N_10572,N_6916,N_7279);
nand U10573 (N_10573,N_8255,N_7672);
nand U10574 (N_10574,N_7232,N_7036);
nor U10575 (N_10575,N_7835,N_6388);
and U10576 (N_10576,N_6299,N_6023);
xnor U10577 (N_10577,N_6883,N_6990);
nor U10578 (N_10578,N_6369,N_6871);
nand U10579 (N_10579,N_7202,N_7245);
and U10580 (N_10580,N_6591,N_8502);
xor U10581 (N_10581,N_7960,N_6387);
nor U10582 (N_10582,N_8649,N_6810);
or U10583 (N_10583,N_6064,N_8609);
or U10584 (N_10584,N_6552,N_7653);
nor U10585 (N_10585,N_7074,N_8382);
nor U10586 (N_10586,N_7484,N_6032);
nor U10587 (N_10587,N_6098,N_8927);
and U10588 (N_10588,N_7983,N_6689);
nor U10589 (N_10589,N_7839,N_7075);
and U10590 (N_10590,N_6964,N_8071);
or U10591 (N_10591,N_7322,N_7354);
and U10592 (N_10592,N_8950,N_6866);
or U10593 (N_10593,N_6690,N_6075);
nor U10594 (N_10594,N_7326,N_8045);
nor U10595 (N_10595,N_6403,N_8991);
and U10596 (N_10596,N_8157,N_7816);
nor U10597 (N_10597,N_7581,N_8445);
and U10598 (N_10598,N_8746,N_8536);
nand U10599 (N_10599,N_6723,N_6715);
or U10600 (N_10600,N_7969,N_6368);
nor U10601 (N_10601,N_8843,N_6333);
or U10602 (N_10602,N_8656,N_7002);
and U10603 (N_10603,N_8537,N_7906);
or U10604 (N_10604,N_8705,N_8922);
and U10605 (N_10605,N_8516,N_6764);
or U10606 (N_10606,N_6758,N_8487);
nor U10607 (N_10607,N_8439,N_7267);
nor U10608 (N_10608,N_6667,N_8979);
nand U10609 (N_10609,N_7381,N_8329);
and U10610 (N_10610,N_7766,N_6070);
nand U10611 (N_10611,N_8810,N_8581);
or U10612 (N_10612,N_6293,N_8034);
or U10613 (N_10613,N_6898,N_8261);
nand U10614 (N_10614,N_6027,N_8691);
nand U10615 (N_10615,N_7836,N_6435);
or U10616 (N_10616,N_8186,N_6841);
or U10617 (N_10617,N_8192,N_7310);
nand U10618 (N_10618,N_8724,N_8335);
or U10619 (N_10619,N_7960,N_7926);
and U10620 (N_10620,N_8873,N_8910);
nor U10621 (N_10621,N_7641,N_6709);
and U10622 (N_10622,N_6605,N_8572);
and U10623 (N_10623,N_6407,N_6568);
nor U10624 (N_10624,N_8007,N_6044);
nand U10625 (N_10625,N_8202,N_8792);
and U10626 (N_10626,N_6483,N_8123);
or U10627 (N_10627,N_7265,N_7984);
nor U10628 (N_10628,N_7960,N_6519);
nor U10629 (N_10629,N_7070,N_7485);
or U10630 (N_10630,N_6429,N_7829);
or U10631 (N_10631,N_7728,N_8293);
nor U10632 (N_10632,N_7964,N_8305);
or U10633 (N_10633,N_6428,N_8347);
nor U10634 (N_10634,N_6859,N_7472);
or U10635 (N_10635,N_8092,N_6410);
nor U10636 (N_10636,N_7805,N_8686);
and U10637 (N_10637,N_6083,N_8226);
and U10638 (N_10638,N_7052,N_8013);
nor U10639 (N_10639,N_6268,N_6282);
xor U10640 (N_10640,N_6179,N_7633);
and U10641 (N_10641,N_8029,N_8771);
nand U10642 (N_10642,N_7031,N_6445);
or U10643 (N_10643,N_8425,N_6043);
xnor U10644 (N_10644,N_8935,N_6349);
nor U10645 (N_10645,N_6601,N_7416);
or U10646 (N_10646,N_6595,N_8547);
xor U10647 (N_10647,N_7439,N_7428);
nor U10648 (N_10648,N_6723,N_7417);
nand U10649 (N_10649,N_7845,N_7021);
nor U10650 (N_10650,N_6162,N_7027);
nand U10651 (N_10651,N_8361,N_6074);
or U10652 (N_10652,N_6017,N_8912);
nor U10653 (N_10653,N_6487,N_7562);
nor U10654 (N_10654,N_8828,N_6091);
nand U10655 (N_10655,N_7640,N_7121);
nor U10656 (N_10656,N_8477,N_7846);
or U10657 (N_10657,N_6065,N_8151);
nor U10658 (N_10658,N_8988,N_8303);
nor U10659 (N_10659,N_7165,N_8860);
nor U10660 (N_10660,N_8803,N_6431);
and U10661 (N_10661,N_6857,N_7930);
or U10662 (N_10662,N_6979,N_6023);
nand U10663 (N_10663,N_8921,N_7267);
nand U10664 (N_10664,N_8491,N_7575);
nand U10665 (N_10665,N_7104,N_6772);
nor U10666 (N_10666,N_8520,N_6151);
or U10667 (N_10667,N_7128,N_7882);
nor U10668 (N_10668,N_8682,N_7902);
nand U10669 (N_10669,N_6685,N_8867);
and U10670 (N_10670,N_7345,N_7660);
or U10671 (N_10671,N_7077,N_7169);
nor U10672 (N_10672,N_7292,N_6996);
or U10673 (N_10673,N_7842,N_7462);
and U10674 (N_10674,N_6686,N_8738);
xnor U10675 (N_10675,N_7159,N_7071);
nand U10676 (N_10676,N_8198,N_8786);
and U10677 (N_10677,N_7923,N_6017);
nand U10678 (N_10678,N_8202,N_6025);
nor U10679 (N_10679,N_6513,N_7041);
or U10680 (N_10680,N_6070,N_6892);
nor U10681 (N_10681,N_8005,N_8614);
or U10682 (N_10682,N_7620,N_8611);
nor U10683 (N_10683,N_8560,N_7411);
or U10684 (N_10684,N_8725,N_7480);
nor U10685 (N_10685,N_6094,N_7597);
or U10686 (N_10686,N_7587,N_7617);
and U10687 (N_10687,N_7980,N_7121);
and U10688 (N_10688,N_7228,N_8963);
and U10689 (N_10689,N_7953,N_6753);
or U10690 (N_10690,N_8042,N_8155);
or U10691 (N_10691,N_6096,N_6176);
and U10692 (N_10692,N_6638,N_6216);
and U10693 (N_10693,N_7280,N_7649);
nor U10694 (N_10694,N_6749,N_7477);
or U10695 (N_10695,N_7591,N_6649);
nand U10696 (N_10696,N_7592,N_7157);
or U10697 (N_10697,N_6051,N_8208);
nor U10698 (N_10698,N_8141,N_8769);
and U10699 (N_10699,N_7554,N_7715);
and U10700 (N_10700,N_6963,N_7848);
nand U10701 (N_10701,N_6733,N_8545);
nand U10702 (N_10702,N_7469,N_6755);
and U10703 (N_10703,N_6260,N_8157);
or U10704 (N_10704,N_7338,N_7095);
nor U10705 (N_10705,N_8456,N_7472);
nor U10706 (N_10706,N_7090,N_7022);
nor U10707 (N_10707,N_6432,N_7462);
nor U10708 (N_10708,N_7904,N_8429);
nor U10709 (N_10709,N_8316,N_8480);
xnor U10710 (N_10710,N_6397,N_6289);
and U10711 (N_10711,N_7492,N_8368);
nor U10712 (N_10712,N_8028,N_6180);
or U10713 (N_10713,N_6694,N_8458);
nor U10714 (N_10714,N_6453,N_8437);
or U10715 (N_10715,N_6119,N_8292);
and U10716 (N_10716,N_7329,N_7587);
nor U10717 (N_10717,N_8560,N_7637);
nor U10718 (N_10718,N_8756,N_8773);
nor U10719 (N_10719,N_6142,N_6793);
xor U10720 (N_10720,N_6121,N_8764);
and U10721 (N_10721,N_8922,N_6535);
xor U10722 (N_10722,N_6489,N_7071);
or U10723 (N_10723,N_8351,N_6103);
or U10724 (N_10724,N_7178,N_6996);
or U10725 (N_10725,N_8579,N_8181);
and U10726 (N_10726,N_6594,N_8733);
nor U10727 (N_10727,N_8813,N_6342);
nand U10728 (N_10728,N_7896,N_8251);
nor U10729 (N_10729,N_7126,N_7205);
or U10730 (N_10730,N_8487,N_7366);
or U10731 (N_10731,N_8130,N_7166);
nand U10732 (N_10732,N_6480,N_8558);
or U10733 (N_10733,N_8777,N_7844);
or U10734 (N_10734,N_6067,N_7818);
and U10735 (N_10735,N_6028,N_6547);
and U10736 (N_10736,N_8437,N_6647);
nand U10737 (N_10737,N_7690,N_7349);
nand U10738 (N_10738,N_6137,N_8916);
nand U10739 (N_10739,N_8611,N_8920);
nor U10740 (N_10740,N_8191,N_8012);
xor U10741 (N_10741,N_8234,N_7905);
and U10742 (N_10742,N_7535,N_6501);
or U10743 (N_10743,N_7934,N_7448);
and U10744 (N_10744,N_7381,N_7147);
nand U10745 (N_10745,N_8161,N_8137);
or U10746 (N_10746,N_8600,N_8928);
or U10747 (N_10747,N_7549,N_7116);
nor U10748 (N_10748,N_7320,N_6970);
nand U10749 (N_10749,N_6686,N_7241);
and U10750 (N_10750,N_8832,N_7866);
nand U10751 (N_10751,N_6229,N_7326);
or U10752 (N_10752,N_6645,N_7153);
or U10753 (N_10753,N_7364,N_7499);
and U10754 (N_10754,N_6133,N_6307);
nor U10755 (N_10755,N_6594,N_7646);
nand U10756 (N_10756,N_8039,N_6900);
or U10757 (N_10757,N_6962,N_7216);
nand U10758 (N_10758,N_7934,N_6144);
or U10759 (N_10759,N_6713,N_7593);
nor U10760 (N_10760,N_8536,N_7013);
or U10761 (N_10761,N_7013,N_6820);
nand U10762 (N_10762,N_6060,N_7451);
and U10763 (N_10763,N_8207,N_7710);
and U10764 (N_10764,N_8267,N_7431);
or U10765 (N_10765,N_7335,N_7188);
nand U10766 (N_10766,N_7378,N_7996);
nand U10767 (N_10767,N_7469,N_8757);
or U10768 (N_10768,N_7101,N_7643);
and U10769 (N_10769,N_6088,N_6250);
and U10770 (N_10770,N_7808,N_6915);
xnor U10771 (N_10771,N_6507,N_8910);
nand U10772 (N_10772,N_7791,N_7363);
nand U10773 (N_10773,N_6752,N_6355);
xor U10774 (N_10774,N_8597,N_8098);
nand U10775 (N_10775,N_7171,N_8898);
or U10776 (N_10776,N_7847,N_7715);
nor U10777 (N_10777,N_8676,N_7629);
nand U10778 (N_10778,N_8754,N_8400);
nand U10779 (N_10779,N_6290,N_8501);
or U10780 (N_10780,N_6475,N_8691);
nor U10781 (N_10781,N_7080,N_8724);
nand U10782 (N_10782,N_8353,N_8926);
and U10783 (N_10783,N_6391,N_7197);
nor U10784 (N_10784,N_8570,N_6713);
nor U10785 (N_10785,N_6448,N_7803);
nor U10786 (N_10786,N_7115,N_7914);
nor U10787 (N_10787,N_7720,N_7719);
or U10788 (N_10788,N_8247,N_6732);
nand U10789 (N_10789,N_7955,N_6192);
and U10790 (N_10790,N_8985,N_6571);
nand U10791 (N_10791,N_7982,N_6780);
nand U10792 (N_10792,N_7207,N_6494);
nand U10793 (N_10793,N_8245,N_7520);
xor U10794 (N_10794,N_7959,N_7835);
or U10795 (N_10795,N_7918,N_8478);
nor U10796 (N_10796,N_7526,N_6355);
nor U10797 (N_10797,N_7967,N_6842);
and U10798 (N_10798,N_6112,N_8763);
or U10799 (N_10799,N_7438,N_8876);
nor U10800 (N_10800,N_6744,N_7673);
or U10801 (N_10801,N_7666,N_6077);
and U10802 (N_10802,N_8091,N_8960);
and U10803 (N_10803,N_7535,N_7126);
or U10804 (N_10804,N_8932,N_6489);
nand U10805 (N_10805,N_8305,N_8223);
nor U10806 (N_10806,N_8472,N_7662);
and U10807 (N_10807,N_8572,N_6206);
and U10808 (N_10808,N_8841,N_8303);
nor U10809 (N_10809,N_6261,N_7873);
nand U10810 (N_10810,N_7285,N_7367);
nand U10811 (N_10811,N_8133,N_7138);
or U10812 (N_10812,N_7845,N_8290);
nor U10813 (N_10813,N_6837,N_7047);
or U10814 (N_10814,N_7356,N_7789);
or U10815 (N_10815,N_8645,N_6025);
or U10816 (N_10816,N_7782,N_6198);
nor U10817 (N_10817,N_7304,N_6672);
nor U10818 (N_10818,N_8292,N_8995);
nor U10819 (N_10819,N_6099,N_7008);
nor U10820 (N_10820,N_6962,N_6632);
nand U10821 (N_10821,N_6513,N_8013);
nand U10822 (N_10822,N_7200,N_8775);
and U10823 (N_10823,N_7743,N_6897);
and U10824 (N_10824,N_7880,N_8537);
xnor U10825 (N_10825,N_8288,N_8581);
xnor U10826 (N_10826,N_7354,N_6767);
and U10827 (N_10827,N_6385,N_7572);
and U10828 (N_10828,N_8912,N_7861);
nor U10829 (N_10829,N_8354,N_8336);
nor U10830 (N_10830,N_7137,N_6272);
or U10831 (N_10831,N_6209,N_8164);
and U10832 (N_10832,N_7040,N_6600);
and U10833 (N_10833,N_7404,N_8387);
nor U10834 (N_10834,N_6618,N_6533);
nand U10835 (N_10835,N_7376,N_7329);
nor U10836 (N_10836,N_8845,N_7525);
or U10837 (N_10837,N_7947,N_6913);
nor U10838 (N_10838,N_7744,N_6875);
nor U10839 (N_10839,N_7859,N_6248);
xnor U10840 (N_10840,N_7443,N_7549);
xor U10841 (N_10841,N_8825,N_6815);
or U10842 (N_10842,N_6416,N_8308);
nand U10843 (N_10843,N_8272,N_8256);
nand U10844 (N_10844,N_6434,N_8299);
or U10845 (N_10845,N_6214,N_8749);
or U10846 (N_10846,N_6316,N_6916);
nand U10847 (N_10847,N_7004,N_8115);
and U10848 (N_10848,N_7650,N_8616);
nor U10849 (N_10849,N_8358,N_6220);
and U10850 (N_10850,N_8019,N_6577);
nand U10851 (N_10851,N_6681,N_7032);
nor U10852 (N_10852,N_7909,N_7847);
nor U10853 (N_10853,N_7931,N_6269);
nand U10854 (N_10854,N_6798,N_8421);
nor U10855 (N_10855,N_8716,N_6333);
nand U10856 (N_10856,N_8658,N_6935);
nor U10857 (N_10857,N_7576,N_8611);
nor U10858 (N_10858,N_6004,N_7750);
nor U10859 (N_10859,N_6818,N_6360);
nand U10860 (N_10860,N_8264,N_7978);
or U10861 (N_10861,N_8300,N_7826);
or U10862 (N_10862,N_8641,N_7010);
nand U10863 (N_10863,N_8049,N_8753);
nor U10864 (N_10864,N_8726,N_6921);
and U10865 (N_10865,N_7542,N_7703);
nand U10866 (N_10866,N_7431,N_8421);
and U10867 (N_10867,N_6721,N_8554);
or U10868 (N_10868,N_7469,N_6053);
or U10869 (N_10869,N_8388,N_8239);
nor U10870 (N_10870,N_8002,N_6509);
or U10871 (N_10871,N_6537,N_7511);
nor U10872 (N_10872,N_8618,N_7620);
nand U10873 (N_10873,N_6062,N_6790);
nand U10874 (N_10874,N_8516,N_7759);
and U10875 (N_10875,N_7511,N_8565);
or U10876 (N_10876,N_8954,N_6045);
nand U10877 (N_10877,N_7170,N_8778);
nand U10878 (N_10878,N_7440,N_7790);
nand U10879 (N_10879,N_8495,N_8266);
nand U10880 (N_10880,N_8339,N_8663);
and U10881 (N_10881,N_6769,N_8136);
nand U10882 (N_10882,N_6535,N_6994);
and U10883 (N_10883,N_8481,N_6778);
or U10884 (N_10884,N_7981,N_8976);
or U10885 (N_10885,N_8825,N_7797);
nor U10886 (N_10886,N_7052,N_6685);
or U10887 (N_10887,N_6984,N_7253);
or U10888 (N_10888,N_8195,N_8185);
or U10889 (N_10889,N_8687,N_7299);
nand U10890 (N_10890,N_7417,N_7087);
and U10891 (N_10891,N_6368,N_8657);
and U10892 (N_10892,N_8736,N_7901);
or U10893 (N_10893,N_7816,N_8580);
nor U10894 (N_10894,N_7409,N_6092);
nor U10895 (N_10895,N_7879,N_6270);
or U10896 (N_10896,N_8627,N_7263);
nor U10897 (N_10897,N_7967,N_7864);
nor U10898 (N_10898,N_6128,N_8129);
or U10899 (N_10899,N_6247,N_7466);
and U10900 (N_10900,N_7610,N_8570);
and U10901 (N_10901,N_8598,N_8614);
and U10902 (N_10902,N_8691,N_7917);
xnor U10903 (N_10903,N_7286,N_6078);
nand U10904 (N_10904,N_7736,N_6004);
nor U10905 (N_10905,N_7675,N_6184);
nand U10906 (N_10906,N_6941,N_6929);
nor U10907 (N_10907,N_7552,N_7213);
nor U10908 (N_10908,N_7795,N_7615);
and U10909 (N_10909,N_7158,N_6120);
and U10910 (N_10910,N_6530,N_6523);
nand U10911 (N_10911,N_8550,N_7162);
nand U10912 (N_10912,N_6306,N_7097);
and U10913 (N_10913,N_7153,N_6557);
or U10914 (N_10914,N_7748,N_7315);
or U10915 (N_10915,N_7658,N_7336);
nand U10916 (N_10916,N_6427,N_6964);
and U10917 (N_10917,N_6735,N_8277);
nor U10918 (N_10918,N_8047,N_7771);
nor U10919 (N_10919,N_6595,N_6797);
or U10920 (N_10920,N_7085,N_6589);
nor U10921 (N_10921,N_8287,N_8866);
or U10922 (N_10922,N_8671,N_7824);
and U10923 (N_10923,N_7159,N_7820);
and U10924 (N_10924,N_7221,N_8785);
and U10925 (N_10925,N_8510,N_8475);
or U10926 (N_10926,N_8739,N_7414);
nand U10927 (N_10927,N_8261,N_6349);
nor U10928 (N_10928,N_8678,N_7324);
and U10929 (N_10929,N_6570,N_6291);
nor U10930 (N_10930,N_7207,N_8284);
nor U10931 (N_10931,N_8610,N_6230);
nand U10932 (N_10932,N_6179,N_6153);
and U10933 (N_10933,N_6376,N_7618);
and U10934 (N_10934,N_6442,N_7673);
nor U10935 (N_10935,N_8964,N_7795);
nor U10936 (N_10936,N_7249,N_7875);
and U10937 (N_10937,N_6011,N_8155);
xor U10938 (N_10938,N_8061,N_7112);
and U10939 (N_10939,N_7102,N_8666);
xnor U10940 (N_10940,N_8051,N_6545);
nor U10941 (N_10941,N_6041,N_6145);
nor U10942 (N_10942,N_8472,N_6832);
or U10943 (N_10943,N_8588,N_6929);
nor U10944 (N_10944,N_6950,N_7096);
or U10945 (N_10945,N_7063,N_7006);
or U10946 (N_10946,N_7170,N_6130);
and U10947 (N_10947,N_7680,N_8269);
and U10948 (N_10948,N_7666,N_8326);
nand U10949 (N_10949,N_8777,N_8543);
or U10950 (N_10950,N_8308,N_7164);
nand U10951 (N_10951,N_8759,N_7771);
or U10952 (N_10952,N_6866,N_7592);
nand U10953 (N_10953,N_7756,N_7905);
nand U10954 (N_10954,N_7658,N_8297);
or U10955 (N_10955,N_8648,N_6483);
nand U10956 (N_10956,N_8078,N_7990);
and U10957 (N_10957,N_7302,N_7703);
and U10958 (N_10958,N_8337,N_6035);
and U10959 (N_10959,N_6313,N_8420);
nand U10960 (N_10960,N_8634,N_7430);
nand U10961 (N_10961,N_7371,N_6542);
xnor U10962 (N_10962,N_6675,N_8142);
or U10963 (N_10963,N_8277,N_7015);
nor U10964 (N_10964,N_8470,N_7792);
nand U10965 (N_10965,N_7576,N_6965);
nor U10966 (N_10966,N_7259,N_7150);
nor U10967 (N_10967,N_8821,N_6634);
nor U10968 (N_10968,N_7273,N_7161);
or U10969 (N_10969,N_7013,N_6550);
nand U10970 (N_10970,N_6327,N_8102);
nand U10971 (N_10971,N_8768,N_8436);
or U10972 (N_10972,N_6608,N_6158);
nor U10973 (N_10973,N_7700,N_6984);
or U10974 (N_10974,N_6750,N_6381);
nand U10975 (N_10975,N_8206,N_7814);
nand U10976 (N_10976,N_8898,N_6818);
and U10977 (N_10977,N_7945,N_8489);
nor U10978 (N_10978,N_6210,N_6923);
nor U10979 (N_10979,N_7642,N_8242);
nor U10980 (N_10980,N_6190,N_6330);
and U10981 (N_10981,N_6084,N_8799);
and U10982 (N_10982,N_8034,N_6956);
and U10983 (N_10983,N_7686,N_8057);
nand U10984 (N_10984,N_8425,N_7484);
nand U10985 (N_10985,N_7709,N_8194);
nand U10986 (N_10986,N_7025,N_6781);
nor U10987 (N_10987,N_7671,N_7642);
nand U10988 (N_10988,N_7065,N_7570);
nor U10989 (N_10989,N_8117,N_8697);
nor U10990 (N_10990,N_6215,N_7526);
nand U10991 (N_10991,N_8372,N_6425);
nand U10992 (N_10992,N_7156,N_6354);
nor U10993 (N_10993,N_6295,N_8569);
or U10994 (N_10994,N_6404,N_8744);
and U10995 (N_10995,N_8077,N_7251);
nand U10996 (N_10996,N_6858,N_6113);
nand U10997 (N_10997,N_7659,N_7368);
or U10998 (N_10998,N_6809,N_8120);
and U10999 (N_10999,N_7468,N_6787);
and U11000 (N_11000,N_6502,N_8114);
or U11001 (N_11001,N_6286,N_6057);
nor U11002 (N_11002,N_8099,N_7518);
nor U11003 (N_11003,N_8814,N_8110);
or U11004 (N_11004,N_8679,N_6642);
or U11005 (N_11005,N_8147,N_6458);
and U11006 (N_11006,N_8202,N_6929);
nor U11007 (N_11007,N_7233,N_6612);
nor U11008 (N_11008,N_6439,N_7831);
nor U11009 (N_11009,N_6256,N_6469);
nor U11010 (N_11010,N_7235,N_8458);
or U11011 (N_11011,N_6162,N_6881);
nor U11012 (N_11012,N_7472,N_7637);
nand U11013 (N_11013,N_8192,N_6358);
nor U11014 (N_11014,N_7165,N_8815);
nor U11015 (N_11015,N_8237,N_6911);
and U11016 (N_11016,N_6391,N_6547);
and U11017 (N_11017,N_7117,N_7319);
xnor U11018 (N_11018,N_8778,N_7146);
nand U11019 (N_11019,N_7025,N_6814);
and U11020 (N_11020,N_8329,N_8314);
nand U11021 (N_11021,N_6104,N_6506);
nand U11022 (N_11022,N_8386,N_8450);
or U11023 (N_11023,N_6679,N_8525);
nor U11024 (N_11024,N_6520,N_8183);
or U11025 (N_11025,N_6619,N_7839);
nand U11026 (N_11026,N_8682,N_6135);
and U11027 (N_11027,N_7416,N_8129);
nor U11028 (N_11028,N_6069,N_6513);
and U11029 (N_11029,N_7465,N_7892);
or U11030 (N_11030,N_7245,N_6263);
nand U11031 (N_11031,N_8929,N_6708);
nor U11032 (N_11032,N_8419,N_6600);
nand U11033 (N_11033,N_8070,N_6019);
nor U11034 (N_11034,N_6268,N_7323);
nand U11035 (N_11035,N_8200,N_7010);
nor U11036 (N_11036,N_6968,N_8521);
and U11037 (N_11037,N_7402,N_7928);
or U11038 (N_11038,N_7597,N_8375);
nand U11039 (N_11039,N_8353,N_6792);
nand U11040 (N_11040,N_7620,N_6190);
and U11041 (N_11041,N_6485,N_8783);
xnor U11042 (N_11042,N_8860,N_7469);
nor U11043 (N_11043,N_8019,N_6834);
nor U11044 (N_11044,N_6726,N_8409);
nor U11045 (N_11045,N_7845,N_8120);
nor U11046 (N_11046,N_7175,N_7495);
nand U11047 (N_11047,N_8203,N_7763);
nor U11048 (N_11048,N_8799,N_7298);
nand U11049 (N_11049,N_6201,N_7960);
or U11050 (N_11050,N_8158,N_6148);
nand U11051 (N_11051,N_7478,N_6510);
nor U11052 (N_11052,N_8130,N_6098);
nor U11053 (N_11053,N_8192,N_8958);
nor U11054 (N_11054,N_7397,N_6816);
and U11055 (N_11055,N_6538,N_8284);
and U11056 (N_11056,N_6670,N_6637);
or U11057 (N_11057,N_6999,N_6347);
and U11058 (N_11058,N_6425,N_7677);
nor U11059 (N_11059,N_7317,N_6594);
nor U11060 (N_11060,N_8745,N_7530);
nand U11061 (N_11061,N_6761,N_8988);
and U11062 (N_11062,N_6119,N_7333);
or U11063 (N_11063,N_8802,N_6014);
or U11064 (N_11064,N_7910,N_8571);
nor U11065 (N_11065,N_8411,N_6366);
and U11066 (N_11066,N_8655,N_7078);
nor U11067 (N_11067,N_7565,N_8835);
nand U11068 (N_11068,N_7191,N_7171);
nand U11069 (N_11069,N_8960,N_6131);
nor U11070 (N_11070,N_6365,N_6006);
or U11071 (N_11071,N_6128,N_6662);
or U11072 (N_11072,N_6544,N_6485);
or U11073 (N_11073,N_8771,N_6816);
nor U11074 (N_11074,N_8617,N_8370);
nand U11075 (N_11075,N_8590,N_6744);
and U11076 (N_11076,N_7357,N_6529);
nor U11077 (N_11077,N_7299,N_6836);
nor U11078 (N_11078,N_6492,N_7318);
nand U11079 (N_11079,N_8653,N_8881);
nand U11080 (N_11080,N_6681,N_8451);
and U11081 (N_11081,N_8218,N_6467);
nand U11082 (N_11082,N_6652,N_6266);
xnor U11083 (N_11083,N_7742,N_6886);
nand U11084 (N_11084,N_7020,N_7439);
and U11085 (N_11085,N_8088,N_8266);
nand U11086 (N_11086,N_6646,N_6812);
nand U11087 (N_11087,N_7551,N_8832);
and U11088 (N_11088,N_7695,N_6109);
and U11089 (N_11089,N_6408,N_7355);
and U11090 (N_11090,N_7862,N_6458);
nor U11091 (N_11091,N_6785,N_8673);
or U11092 (N_11092,N_7427,N_7373);
nor U11093 (N_11093,N_7860,N_8833);
or U11094 (N_11094,N_8179,N_7044);
nand U11095 (N_11095,N_6697,N_7300);
or U11096 (N_11096,N_8207,N_8266);
nor U11097 (N_11097,N_8778,N_8910);
and U11098 (N_11098,N_6468,N_7681);
nand U11099 (N_11099,N_8737,N_7409);
nand U11100 (N_11100,N_8948,N_6915);
nand U11101 (N_11101,N_6143,N_6246);
nor U11102 (N_11102,N_8312,N_6039);
or U11103 (N_11103,N_6514,N_7620);
or U11104 (N_11104,N_6682,N_7119);
nor U11105 (N_11105,N_7398,N_8703);
or U11106 (N_11106,N_7985,N_8815);
nand U11107 (N_11107,N_7992,N_6327);
nand U11108 (N_11108,N_6640,N_7347);
nor U11109 (N_11109,N_6745,N_6095);
nor U11110 (N_11110,N_7943,N_6993);
and U11111 (N_11111,N_8566,N_7936);
or U11112 (N_11112,N_8015,N_6783);
nand U11113 (N_11113,N_7466,N_6436);
or U11114 (N_11114,N_6803,N_6094);
or U11115 (N_11115,N_7812,N_6340);
nand U11116 (N_11116,N_8261,N_7632);
or U11117 (N_11117,N_8310,N_7576);
and U11118 (N_11118,N_8750,N_7121);
nor U11119 (N_11119,N_7237,N_6207);
and U11120 (N_11120,N_8602,N_6499);
and U11121 (N_11121,N_7359,N_6943);
and U11122 (N_11122,N_6617,N_6890);
nor U11123 (N_11123,N_6201,N_7541);
and U11124 (N_11124,N_8986,N_7111);
nand U11125 (N_11125,N_6816,N_6262);
nand U11126 (N_11126,N_6459,N_6821);
nor U11127 (N_11127,N_7845,N_6932);
nand U11128 (N_11128,N_8896,N_6770);
and U11129 (N_11129,N_8888,N_7379);
nand U11130 (N_11130,N_7818,N_6394);
and U11131 (N_11131,N_6704,N_6957);
nor U11132 (N_11132,N_7598,N_7242);
nand U11133 (N_11133,N_7198,N_7676);
nand U11134 (N_11134,N_8325,N_6116);
nand U11135 (N_11135,N_6787,N_7111);
xor U11136 (N_11136,N_7441,N_6480);
and U11137 (N_11137,N_7889,N_8704);
nand U11138 (N_11138,N_6526,N_8329);
nor U11139 (N_11139,N_6534,N_6162);
nand U11140 (N_11140,N_8914,N_8160);
nor U11141 (N_11141,N_6584,N_7442);
nand U11142 (N_11142,N_7267,N_8969);
or U11143 (N_11143,N_7834,N_8123);
nor U11144 (N_11144,N_8660,N_6539);
xnor U11145 (N_11145,N_7011,N_6206);
or U11146 (N_11146,N_6536,N_6615);
nand U11147 (N_11147,N_6945,N_7146);
nand U11148 (N_11148,N_7350,N_6500);
and U11149 (N_11149,N_7002,N_6586);
and U11150 (N_11150,N_8063,N_7820);
and U11151 (N_11151,N_6981,N_8289);
nand U11152 (N_11152,N_7674,N_8264);
and U11153 (N_11153,N_7973,N_6922);
nor U11154 (N_11154,N_8690,N_7079);
nor U11155 (N_11155,N_6399,N_8284);
nand U11156 (N_11156,N_6431,N_8405);
nor U11157 (N_11157,N_6733,N_6342);
or U11158 (N_11158,N_7643,N_7237);
and U11159 (N_11159,N_6401,N_6808);
and U11160 (N_11160,N_7804,N_6472);
or U11161 (N_11161,N_8473,N_6614);
or U11162 (N_11162,N_7283,N_7423);
nor U11163 (N_11163,N_6721,N_8232);
nor U11164 (N_11164,N_6662,N_6989);
and U11165 (N_11165,N_8035,N_6070);
nor U11166 (N_11166,N_8312,N_8393);
and U11167 (N_11167,N_6625,N_8916);
and U11168 (N_11168,N_7115,N_7586);
or U11169 (N_11169,N_6841,N_7514);
and U11170 (N_11170,N_8091,N_7773);
and U11171 (N_11171,N_7110,N_6941);
nor U11172 (N_11172,N_6516,N_6019);
or U11173 (N_11173,N_6004,N_8586);
and U11174 (N_11174,N_8323,N_8313);
and U11175 (N_11175,N_8053,N_7751);
xor U11176 (N_11176,N_7651,N_7428);
nor U11177 (N_11177,N_7356,N_6750);
or U11178 (N_11178,N_8163,N_8441);
and U11179 (N_11179,N_6998,N_6799);
or U11180 (N_11180,N_6232,N_8848);
and U11181 (N_11181,N_8306,N_7429);
nand U11182 (N_11182,N_7961,N_6284);
xnor U11183 (N_11183,N_7812,N_8507);
or U11184 (N_11184,N_6787,N_8172);
or U11185 (N_11185,N_7006,N_8814);
or U11186 (N_11186,N_7456,N_8094);
nor U11187 (N_11187,N_7354,N_8774);
or U11188 (N_11188,N_7436,N_8037);
or U11189 (N_11189,N_8372,N_8803);
and U11190 (N_11190,N_7315,N_8026);
and U11191 (N_11191,N_6594,N_7788);
nor U11192 (N_11192,N_6116,N_6754);
nand U11193 (N_11193,N_8725,N_8475);
xnor U11194 (N_11194,N_8580,N_8267);
nor U11195 (N_11195,N_8873,N_8582);
nand U11196 (N_11196,N_7638,N_6668);
and U11197 (N_11197,N_8917,N_8670);
nor U11198 (N_11198,N_6673,N_6145);
and U11199 (N_11199,N_6580,N_8197);
nor U11200 (N_11200,N_8622,N_8326);
or U11201 (N_11201,N_8692,N_7578);
and U11202 (N_11202,N_7464,N_8819);
nand U11203 (N_11203,N_6624,N_7757);
nand U11204 (N_11204,N_7361,N_7162);
and U11205 (N_11205,N_8065,N_6742);
or U11206 (N_11206,N_6359,N_8164);
nor U11207 (N_11207,N_8576,N_7882);
nor U11208 (N_11208,N_7233,N_8150);
nor U11209 (N_11209,N_8827,N_6732);
nor U11210 (N_11210,N_7123,N_8432);
and U11211 (N_11211,N_7733,N_6482);
nor U11212 (N_11212,N_6668,N_7679);
nand U11213 (N_11213,N_7433,N_8210);
nand U11214 (N_11214,N_7082,N_8151);
nand U11215 (N_11215,N_7534,N_6703);
or U11216 (N_11216,N_6222,N_6290);
nor U11217 (N_11217,N_8407,N_7714);
xnor U11218 (N_11218,N_6057,N_7179);
and U11219 (N_11219,N_8922,N_8822);
or U11220 (N_11220,N_7315,N_7510);
and U11221 (N_11221,N_6049,N_6104);
and U11222 (N_11222,N_6498,N_8157);
and U11223 (N_11223,N_7433,N_7102);
and U11224 (N_11224,N_8561,N_7969);
or U11225 (N_11225,N_8581,N_7736);
or U11226 (N_11226,N_6587,N_7222);
and U11227 (N_11227,N_6762,N_7675);
nor U11228 (N_11228,N_8573,N_7698);
nand U11229 (N_11229,N_6082,N_7901);
or U11230 (N_11230,N_6076,N_7845);
nor U11231 (N_11231,N_6743,N_7214);
nand U11232 (N_11232,N_6612,N_7339);
nor U11233 (N_11233,N_8007,N_8412);
nor U11234 (N_11234,N_7119,N_7594);
nor U11235 (N_11235,N_6085,N_6732);
nand U11236 (N_11236,N_8432,N_6233);
and U11237 (N_11237,N_7325,N_8606);
nor U11238 (N_11238,N_6805,N_8670);
nor U11239 (N_11239,N_8511,N_7717);
and U11240 (N_11240,N_7114,N_8581);
and U11241 (N_11241,N_8337,N_8931);
and U11242 (N_11242,N_8316,N_8814);
or U11243 (N_11243,N_6000,N_6592);
nor U11244 (N_11244,N_7192,N_8149);
nand U11245 (N_11245,N_7514,N_6524);
xnor U11246 (N_11246,N_8757,N_7744);
and U11247 (N_11247,N_6430,N_8697);
and U11248 (N_11248,N_7108,N_6885);
nand U11249 (N_11249,N_7947,N_7932);
and U11250 (N_11250,N_8624,N_6387);
nand U11251 (N_11251,N_6660,N_6309);
and U11252 (N_11252,N_6607,N_8859);
and U11253 (N_11253,N_7953,N_8514);
or U11254 (N_11254,N_8911,N_8821);
or U11255 (N_11255,N_6269,N_6011);
and U11256 (N_11256,N_7446,N_6417);
nor U11257 (N_11257,N_6160,N_8536);
and U11258 (N_11258,N_7363,N_8078);
or U11259 (N_11259,N_8958,N_7904);
nor U11260 (N_11260,N_6745,N_6962);
and U11261 (N_11261,N_6980,N_7937);
nand U11262 (N_11262,N_7061,N_8308);
nor U11263 (N_11263,N_7285,N_7206);
or U11264 (N_11264,N_7506,N_7785);
and U11265 (N_11265,N_7011,N_8198);
or U11266 (N_11266,N_6518,N_6153);
nand U11267 (N_11267,N_8072,N_6568);
and U11268 (N_11268,N_7367,N_8402);
nor U11269 (N_11269,N_6118,N_7230);
and U11270 (N_11270,N_6058,N_6578);
nand U11271 (N_11271,N_6274,N_7970);
nor U11272 (N_11272,N_7629,N_8995);
or U11273 (N_11273,N_8203,N_6106);
nor U11274 (N_11274,N_6214,N_7000);
nand U11275 (N_11275,N_8884,N_7642);
and U11276 (N_11276,N_8442,N_7126);
and U11277 (N_11277,N_7598,N_8530);
nand U11278 (N_11278,N_7371,N_8212);
nand U11279 (N_11279,N_8072,N_8215);
and U11280 (N_11280,N_8637,N_6399);
xnor U11281 (N_11281,N_6020,N_6018);
or U11282 (N_11282,N_7331,N_7177);
nand U11283 (N_11283,N_8342,N_7248);
nand U11284 (N_11284,N_7518,N_7779);
nor U11285 (N_11285,N_8367,N_6928);
or U11286 (N_11286,N_6403,N_6087);
nor U11287 (N_11287,N_6860,N_6613);
nand U11288 (N_11288,N_6567,N_6256);
nor U11289 (N_11289,N_7519,N_6406);
nand U11290 (N_11290,N_8913,N_8568);
or U11291 (N_11291,N_7549,N_7491);
and U11292 (N_11292,N_6317,N_6431);
or U11293 (N_11293,N_8176,N_7431);
xnor U11294 (N_11294,N_7262,N_7892);
nand U11295 (N_11295,N_6410,N_7891);
and U11296 (N_11296,N_8950,N_7043);
nand U11297 (N_11297,N_7496,N_6306);
or U11298 (N_11298,N_8182,N_8956);
or U11299 (N_11299,N_8577,N_6078);
nand U11300 (N_11300,N_8331,N_8392);
or U11301 (N_11301,N_8641,N_6966);
xnor U11302 (N_11302,N_6122,N_8660);
xnor U11303 (N_11303,N_8507,N_7787);
and U11304 (N_11304,N_8072,N_6780);
nand U11305 (N_11305,N_8448,N_6422);
or U11306 (N_11306,N_7696,N_7242);
nor U11307 (N_11307,N_8078,N_7217);
or U11308 (N_11308,N_7428,N_8451);
and U11309 (N_11309,N_8622,N_6833);
nor U11310 (N_11310,N_8625,N_7145);
nor U11311 (N_11311,N_8914,N_7042);
or U11312 (N_11312,N_7687,N_7265);
or U11313 (N_11313,N_7254,N_8061);
or U11314 (N_11314,N_7965,N_7573);
or U11315 (N_11315,N_7445,N_7930);
nor U11316 (N_11316,N_7351,N_6224);
nor U11317 (N_11317,N_7453,N_6183);
nand U11318 (N_11318,N_7072,N_7834);
and U11319 (N_11319,N_6702,N_8715);
nor U11320 (N_11320,N_7737,N_6713);
or U11321 (N_11321,N_7906,N_8786);
nor U11322 (N_11322,N_6769,N_7400);
nand U11323 (N_11323,N_7021,N_7375);
and U11324 (N_11324,N_8585,N_6612);
nor U11325 (N_11325,N_6877,N_6464);
and U11326 (N_11326,N_8103,N_6094);
nand U11327 (N_11327,N_8158,N_7619);
nor U11328 (N_11328,N_8821,N_6198);
nor U11329 (N_11329,N_8793,N_6543);
or U11330 (N_11330,N_7609,N_6027);
and U11331 (N_11331,N_6531,N_8596);
or U11332 (N_11332,N_6732,N_8052);
or U11333 (N_11333,N_8977,N_8351);
nand U11334 (N_11334,N_6060,N_6984);
nor U11335 (N_11335,N_7876,N_7706);
and U11336 (N_11336,N_8198,N_6507);
nor U11337 (N_11337,N_7862,N_6658);
nand U11338 (N_11338,N_8516,N_8775);
nand U11339 (N_11339,N_7802,N_8077);
nor U11340 (N_11340,N_6309,N_8795);
nor U11341 (N_11341,N_7960,N_8243);
or U11342 (N_11342,N_8676,N_7157);
and U11343 (N_11343,N_7978,N_6267);
nand U11344 (N_11344,N_6438,N_6625);
and U11345 (N_11345,N_8974,N_7321);
xor U11346 (N_11346,N_6704,N_8384);
and U11347 (N_11347,N_7325,N_8911);
nor U11348 (N_11348,N_8894,N_6196);
nand U11349 (N_11349,N_6520,N_8547);
nor U11350 (N_11350,N_6781,N_7614);
nor U11351 (N_11351,N_8962,N_8387);
nor U11352 (N_11352,N_8139,N_6376);
and U11353 (N_11353,N_6302,N_7116);
and U11354 (N_11354,N_7816,N_7636);
or U11355 (N_11355,N_6185,N_6441);
and U11356 (N_11356,N_7115,N_8137);
nand U11357 (N_11357,N_7517,N_7068);
nand U11358 (N_11358,N_6905,N_8403);
nor U11359 (N_11359,N_6043,N_6241);
nor U11360 (N_11360,N_8146,N_8238);
or U11361 (N_11361,N_8916,N_7673);
nor U11362 (N_11362,N_6357,N_8773);
and U11363 (N_11363,N_8334,N_7381);
nor U11364 (N_11364,N_6720,N_7414);
nor U11365 (N_11365,N_6559,N_7043);
nand U11366 (N_11366,N_6956,N_7246);
nor U11367 (N_11367,N_8533,N_8432);
or U11368 (N_11368,N_6789,N_8581);
and U11369 (N_11369,N_8016,N_7663);
nand U11370 (N_11370,N_8549,N_7058);
nand U11371 (N_11371,N_7492,N_6478);
nor U11372 (N_11372,N_8354,N_8790);
or U11373 (N_11373,N_6224,N_8652);
nand U11374 (N_11374,N_6237,N_6404);
xnor U11375 (N_11375,N_8539,N_8476);
nor U11376 (N_11376,N_6800,N_6282);
nor U11377 (N_11377,N_7231,N_6073);
nor U11378 (N_11378,N_8533,N_6997);
xnor U11379 (N_11379,N_8996,N_7730);
and U11380 (N_11380,N_8973,N_7972);
and U11381 (N_11381,N_7371,N_8270);
and U11382 (N_11382,N_8676,N_7360);
nand U11383 (N_11383,N_7329,N_8151);
and U11384 (N_11384,N_6094,N_6864);
or U11385 (N_11385,N_8567,N_8293);
and U11386 (N_11386,N_8505,N_8085);
or U11387 (N_11387,N_7933,N_7751);
nor U11388 (N_11388,N_7136,N_8534);
nand U11389 (N_11389,N_6965,N_6540);
xnor U11390 (N_11390,N_7493,N_6601);
or U11391 (N_11391,N_8266,N_7032);
xor U11392 (N_11392,N_7677,N_8565);
or U11393 (N_11393,N_8515,N_7385);
nor U11394 (N_11394,N_7428,N_6613);
nor U11395 (N_11395,N_6610,N_6758);
nor U11396 (N_11396,N_8274,N_7443);
and U11397 (N_11397,N_7649,N_8188);
or U11398 (N_11398,N_6941,N_6468);
or U11399 (N_11399,N_6069,N_8489);
nor U11400 (N_11400,N_6725,N_8983);
and U11401 (N_11401,N_7778,N_7388);
nand U11402 (N_11402,N_6688,N_8500);
nand U11403 (N_11403,N_6319,N_6522);
nor U11404 (N_11404,N_7604,N_8745);
nand U11405 (N_11405,N_8560,N_6870);
and U11406 (N_11406,N_7909,N_7389);
nor U11407 (N_11407,N_7470,N_8583);
and U11408 (N_11408,N_7574,N_7829);
nand U11409 (N_11409,N_7227,N_8680);
nand U11410 (N_11410,N_8302,N_7907);
and U11411 (N_11411,N_6802,N_6402);
nand U11412 (N_11412,N_7794,N_7061);
nand U11413 (N_11413,N_7591,N_6303);
or U11414 (N_11414,N_7292,N_8998);
nor U11415 (N_11415,N_8864,N_6519);
or U11416 (N_11416,N_7834,N_7767);
or U11417 (N_11417,N_7501,N_7362);
or U11418 (N_11418,N_7913,N_6160);
and U11419 (N_11419,N_7628,N_6637);
nand U11420 (N_11420,N_6290,N_6260);
and U11421 (N_11421,N_7924,N_8267);
and U11422 (N_11422,N_8690,N_8332);
nor U11423 (N_11423,N_8732,N_8951);
and U11424 (N_11424,N_6257,N_6602);
nand U11425 (N_11425,N_7342,N_8335);
and U11426 (N_11426,N_8105,N_7498);
or U11427 (N_11427,N_8657,N_6490);
or U11428 (N_11428,N_8953,N_8383);
nor U11429 (N_11429,N_7254,N_8327);
nand U11430 (N_11430,N_8146,N_7106);
xnor U11431 (N_11431,N_8434,N_7155);
nand U11432 (N_11432,N_8191,N_7999);
nor U11433 (N_11433,N_8710,N_6118);
nand U11434 (N_11434,N_7935,N_8137);
xnor U11435 (N_11435,N_8425,N_7462);
and U11436 (N_11436,N_6738,N_6568);
nor U11437 (N_11437,N_6546,N_8470);
or U11438 (N_11438,N_6212,N_7729);
and U11439 (N_11439,N_8479,N_7191);
and U11440 (N_11440,N_8775,N_7487);
and U11441 (N_11441,N_8527,N_7966);
and U11442 (N_11442,N_7443,N_7386);
or U11443 (N_11443,N_7467,N_6218);
nand U11444 (N_11444,N_6843,N_6539);
and U11445 (N_11445,N_6521,N_6387);
or U11446 (N_11446,N_7806,N_6991);
and U11447 (N_11447,N_6928,N_8210);
or U11448 (N_11448,N_7495,N_7284);
or U11449 (N_11449,N_8988,N_8983);
and U11450 (N_11450,N_6812,N_6008);
and U11451 (N_11451,N_7499,N_7465);
and U11452 (N_11452,N_7134,N_7239);
or U11453 (N_11453,N_8071,N_6285);
nor U11454 (N_11454,N_7538,N_6375);
nand U11455 (N_11455,N_7317,N_7228);
or U11456 (N_11456,N_7442,N_8802);
nor U11457 (N_11457,N_7013,N_7312);
nand U11458 (N_11458,N_6285,N_6521);
nor U11459 (N_11459,N_7832,N_7002);
or U11460 (N_11460,N_8849,N_7343);
and U11461 (N_11461,N_7379,N_6273);
nor U11462 (N_11462,N_6360,N_8079);
nand U11463 (N_11463,N_7539,N_7371);
nand U11464 (N_11464,N_8768,N_8793);
xnor U11465 (N_11465,N_6651,N_8556);
or U11466 (N_11466,N_7840,N_8127);
nor U11467 (N_11467,N_7074,N_6928);
and U11468 (N_11468,N_8723,N_8518);
nor U11469 (N_11469,N_6736,N_6159);
or U11470 (N_11470,N_6001,N_6133);
nand U11471 (N_11471,N_8194,N_8354);
nand U11472 (N_11472,N_8449,N_7264);
or U11473 (N_11473,N_6032,N_7501);
and U11474 (N_11474,N_8980,N_6610);
xor U11475 (N_11475,N_7258,N_7298);
nor U11476 (N_11476,N_6070,N_7368);
nand U11477 (N_11477,N_7795,N_8116);
or U11478 (N_11478,N_7956,N_7330);
or U11479 (N_11479,N_8472,N_7881);
nor U11480 (N_11480,N_8447,N_7184);
or U11481 (N_11481,N_7098,N_8444);
or U11482 (N_11482,N_6342,N_8920);
nand U11483 (N_11483,N_6568,N_8686);
nand U11484 (N_11484,N_7188,N_6517);
nand U11485 (N_11485,N_8208,N_7777);
nor U11486 (N_11486,N_8826,N_6700);
nand U11487 (N_11487,N_6466,N_7407);
and U11488 (N_11488,N_7575,N_7654);
nor U11489 (N_11489,N_8604,N_6027);
nor U11490 (N_11490,N_8206,N_6533);
nor U11491 (N_11491,N_6692,N_6305);
or U11492 (N_11492,N_6183,N_7356);
nor U11493 (N_11493,N_7623,N_8544);
or U11494 (N_11494,N_8189,N_6664);
and U11495 (N_11495,N_7216,N_8105);
nand U11496 (N_11496,N_6045,N_7023);
or U11497 (N_11497,N_8756,N_6188);
nand U11498 (N_11498,N_7200,N_6309);
nor U11499 (N_11499,N_7954,N_6278);
nand U11500 (N_11500,N_6921,N_7089);
nor U11501 (N_11501,N_7207,N_8691);
and U11502 (N_11502,N_8212,N_6741);
xor U11503 (N_11503,N_8012,N_8927);
and U11504 (N_11504,N_6690,N_6972);
or U11505 (N_11505,N_6305,N_6102);
or U11506 (N_11506,N_7400,N_6883);
or U11507 (N_11507,N_8242,N_8669);
or U11508 (N_11508,N_6166,N_6706);
or U11509 (N_11509,N_8845,N_8480);
nor U11510 (N_11510,N_7572,N_6782);
nand U11511 (N_11511,N_6089,N_7464);
nor U11512 (N_11512,N_6831,N_6414);
nor U11513 (N_11513,N_6472,N_7841);
or U11514 (N_11514,N_8344,N_6153);
and U11515 (N_11515,N_7545,N_7730);
and U11516 (N_11516,N_7163,N_6790);
nor U11517 (N_11517,N_8744,N_6252);
nand U11518 (N_11518,N_7467,N_6939);
nor U11519 (N_11519,N_7039,N_7438);
and U11520 (N_11520,N_8917,N_8843);
or U11521 (N_11521,N_6518,N_8447);
and U11522 (N_11522,N_7240,N_8931);
and U11523 (N_11523,N_8618,N_8379);
or U11524 (N_11524,N_8390,N_6618);
or U11525 (N_11525,N_6061,N_6361);
and U11526 (N_11526,N_6070,N_7749);
or U11527 (N_11527,N_7611,N_7426);
nor U11528 (N_11528,N_6869,N_8008);
or U11529 (N_11529,N_6864,N_7729);
nor U11530 (N_11530,N_7924,N_8399);
nor U11531 (N_11531,N_6092,N_6319);
nor U11532 (N_11532,N_6758,N_6010);
nor U11533 (N_11533,N_8200,N_6771);
xnor U11534 (N_11534,N_6336,N_6180);
nor U11535 (N_11535,N_6533,N_7847);
nand U11536 (N_11536,N_8243,N_8941);
nand U11537 (N_11537,N_8309,N_7853);
or U11538 (N_11538,N_8448,N_7574);
nor U11539 (N_11539,N_8325,N_7855);
or U11540 (N_11540,N_8099,N_6669);
or U11541 (N_11541,N_7458,N_6358);
or U11542 (N_11542,N_8414,N_8918);
nand U11543 (N_11543,N_7999,N_8581);
or U11544 (N_11544,N_8967,N_7887);
nand U11545 (N_11545,N_7600,N_7148);
and U11546 (N_11546,N_6951,N_7051);
and U11547 (N_11547,N_7231,N_7912);
nor U11548 (N_11548,N_8772,N_7278);
nor U11549 (N_11549,N_6339,N_6983);
nand U11550 (N_11550,N_6028,N_6125);
nor U11551 (N_11551,N_6899,N_8492);
nor U11552 (N_11552,N_7967,N_7051);
nand U11553 (N_11553,N_7671,N_7753);
nor U11554 (N_11554,N_7722,N_7616);
nor U11555 (N_11555,N_6826,N_8346);
xnor U11556 (N_11556,N_6262,N_8132);
and U11557 (N_11557,N_7915,N_8952);
or U11558 (N_11558,N_8391,N_6365);
xnor U11559 (N_11559,N_8551,N_7114);
nor U11560 (N_11560,N_6519,N_7065);
nor U11561 (N_11561,N_7062,N_7297);
nor U11562 (N_11562,N_8449,N_6477);
and U11563 (N_11563,N_6489,N_8847);
nor U11564 (N_11564,N_8033,N_6519);
nand U11565 (N_11565,N_6346,N_8284);
nor U11566 (N_11566,N_6658,N_7589);
or U11567 (N_11567,N_7428,N_6535);
or U11568 (N_11568,N_6659,N_6849);
and U11569 (N_11569,N_8991,N_6919);
nand U11570 (N_11570,N_7591,N_7466);
nor U11571 (N_11571,N_7479,N_8974);
or U11572 (N_11572,N_8005,N_7052);
nand U11573 (N_11573,N_6439,N_8748);
nand U11574 (N_11574,N_8767,N_6305);
nand U11575 (N_11575,N_6814,N_6225);
nor U11576 (N_11576,N_6051,N_6914);
nand U11577 (N_11577,N_7309,N_7610);
nand U11578 (N_11578,N_8803,N_7528);
nor U11579 (N_11579,N_7169,N_8069);
or U11580 (N_11580,N_7226,N_8196);
nand U11581 (N_11581,N_6539,N_8980);
nor U11582 (N_11582,N_7819,N_7082);
or U11583 (N_11583,N_6257,N_8375);
and U11584 (N_11584,N_7153,N_7583);
nand U11585 (N_11585,N_7946,N_7045);
or U11586 (N_11586,N_8405,N_7816);
and U11587 (N_11587,N_6819,N_7416);
and U11588 (N_11588,N_6121,N_7356);
or U11589 (N_11589,N_6110,N_8773);
nand U11590 (N_11590,N_7129,N_7316);
nand U11591 (N_11591,N_6490,N_8729);
or U11592 (N_11592,N_6704,N_7740);
and U11593 (N_11593,N_6940,N_8232);
and U11594 (N_11594,N_8601,N_6484);
nand U11595 (N_11595,N_6079,N_6909);
nor U11596 (N_11596,N_7946,N_7667);
nand U11597 (N_11597,N_7579,N_8224);
and U11598 (N_11598,N_8011,N_6945);
nor U11599 (N_11599,N_6041,N_6719);
nand U11600 (N_11600,N_7975,N_7387);
and U11601 (N_11601,N_6564,N_8410);
or U11602 (N_11602,N_6246,N_8683);
and U11603 (N_11603,N_6366,N_6811);
nor U11604 (N_11604,N_8317,N_8919);
or U11605 (N_11605,N_7147,N_7752);
xnor U11606 (N_11606,N_8123,N_7885);
and U11607 (N_11607,N_6030,N_8851);
and U11608 (N_11608,N_6397,N_7091);
or U11609 (N_11609,N_7917,N_6040);
or U11610 (N_11610,N_7957,N_6057);
nor U11611 (N_11611,N_7017,N_8886);
or U11612 (N_11612,N_7655,N_7689);
xor U11613 (N_11613,N_8721,N_6885);
nor U11614 (N_11614,N_6977,N_6354);
and U11615 (N_11615,N_6550,N_7719);
and U11616 (N_11616,N_6251,N_8897);
or U11617 (N_11617,N_8100,N_6320);
or U11618 (N_11618,N_6305,N_8788);
or U11619 (N_11619,N_8472,N_8579);
and U11620 (N_11620,N_8764,N_6594);
nand U11621 (N_11621,N_6608,N_6359);
nand U11622 (N_11622,N_6805,N_6662);
nor U11623 (N_11623,N_8413,N_6028);
or U11624 (N_11624,N_6534,N_6919);
nand U11625 (N_11625,N_8109,N_6629);
or U11626 (N_11626,N_7364,N_6931);
nand U11627 (N_11627,N_7976,N_7227);
or U11628 (N_11628,N_6865,N_7082);
nand U11629 (N_11629,N_6449,N_8755);
nand U11630 (N_11630,N_8967,N_7731);
or U11631 (N_11631,N_8232,N_6158);
nor U11632 (N_11632,N_6069,N_6509);
nor U11633 (N_11633,N_6039,N_7646);
nor U11634 (N_11634,N_7990,N_8438);
nor U11635 (N_11635,N_8958,N_8406);
nor U11636 (N_11636,N_6724,N_8248);
and U11637 (N_11637,N_6598,N_8771);
nand U11638 (N_11638,N_7807,N_8671);
or U11639 (N_11639,N_6944,N_7949);
nand U11640 (N_11640,N_8480,N_8797);
and U11641 (N_11641,N_6486,N_8573);
nor U11642 (N_11642,N_8475,N_8994);
xor U11643 (N_11643,N_6402,N_7961);
and U11644 (N_11644,N_7695,N_6588);
nand U11645 (N_11645,N_6944,N_7143);
and U11646 (N_11646,N_8150,N_6776);
and U11647 (N_11647,N_8809,N_6954);
or U11648 (N_11648,N_6595,N_6319);
and U11649 (N_11649,N_6358,N_8646);
nor U11650 (N_11650,N_7709,N_6071);
and U11651 (N_11651,N_7210,N_6551);
or U11652 (N_11652,N_8752,N_7153);
or U11653 (N_11653,N_8400,N_8573);
xor U11654 (N_11654,N_7022,N_8703);
and U11655 (N_11655,N_8363,N_8942);
or U11656 (N_11656,N_7746,N_7423);
nor U11657 (N_11657,N_7389,N_8406);
xnor U11658 (N_11658,N_6730,N_6066);
nand U11659 (N_11659,N_8954,N_7913);
xnor U11660 (N_11660,N_8092,N_7897);
xnor U11661 (N_11661,N_6369,N_6668);
nor U11662 (N_11662,N_7116,N_6248);
nand U11663 (N_11663,N_7668,N_7616);
and U11664 (N_11664,N_6972,N_8668);
nor U11665 (N_11665,N_8109,N_8260);
nor U11666 (N_11666,N_6962,N_8963);
and U11667 (N_11667,N_6056,N_6195);
nand U11668 (N_11668,N_7267,N_7069);
and U11669 (N_11669,N_7667,N_7754);
xor U11670 (N_11670,N_6878,N_8850);
and U11671 (N_11671,N_7139,N_7257);
and U11672 (N_11672,N_7619,N_6549);
or U11673 (N_11673,N_8411,N_8410);
and U11674 (N_11674,N_7369,N_7900);
and U11675 (N_11675,N_8239,N_8530);
nor U11676 (N_11676,N_8405,N_6362);
or U11677 (N_11677,N_6700,N_7235);
or U11678 (N_11678,N_6609,N_6864);
and U11679 (N_11679,N_6703,N_8945);
nand U11680 (N_11680,N_8888,N_8442);
nor U11681 (N_11681,N_8507,N_6939);
nor U11682 (N_11682,N_7559,N_7475);
or U11683 (N_11683,N_8033,N_6958);
and U11684 (N_11684,N_8735,N_6580);
nor U11685 (N_11685,N_8144,N_7837);
and U11686 (N_11686,N_7029,N_7589);
nor U11687 (N_11687,N_7167,N_7047);
and U11688 (N_11688,N_6357,N_7306);
and U11689 (N_11689,N_8857,N_6513);
nand U11690 (N_11690,N_6042,N_7051);
nand U11691 (N_11691,N_6967,N_7144);
nor U11692 (N_11692,N_8407,N_6022);
or U11693 (N_11693,N_8444,N_8627);
xor U11694 (N_11694,N_7092,N_8071);
nor U11695 (N_11695,N_8629,N_7375);
or U11696 (N_11696,N_7359,N_7670);
or U11697 (N_11697,N_7022,N_6229);
or U11698 (N_11698,N_7623,N_8057);
nand U11699 (N_11699,N_8387,N_7727);
and U11700 (N_11700,N_8696,N_7626);
and U11701 (N_11701,N_8687,N_8362);
or U11702 (N_11702,N_8486,N_8367);
nand U11703 (N_11703,N_8110,N_8936);
nor U11704 (N_11704,N_6250,N_7102);
or U11705 (N_11705,N_7724,N_6787);
nand U11706 (N_11706,N_7639,N_8427);
and U11707 (N_11707,N_8368,N_8126);
nor U11708 (N_11708,N_7472,N_7918);
nand U11709 (N_11709,N_8637,N_6809);
or U11710 (N_11710,N_8312,N_8903);
nand U11711 (N_11711,N_6097,N_6602);
or U11712 (N_11712,N_6089,N_7762);
nor U11713 (N_11713,N_7390,N_6353);
and U11714 (N_11714,N_6968,N_7250);
nand U11715 (N_11715,N_7415,N_7204);
nand U11716 (N_11716,N_8020,N_6782);
nor U11717 (N_11717,N_8845,N_7822);
or U11718 (N_11718,N_7421,N_7618);
or U11719 (N_11719,N_7560,N_6285);
and U11720 (N_11720,N_8365,N_7801);
and U11721 (N_11721,N_8345,N_7663);
nor U11722 (N_11722,N_8739,N_8523);
nor U11723 (N_11723,N_8902,N_6064);
xnor U11724 (N_11724,N_8731,N_7709);
nand U11725 (N_11725,N_7832,N_7172);
and U11726 (N_11726,N_8123,N_8852);
nand U11727 (N_11727,N_7208,N_7387);
nand U11728 (N_11728,N_6326,N_8601);
and U11729 (N_11729,N_8166,N_7818);
xnor U11730 (N_11730,N_7074,N_7427);
nor U11731 (N_11731,N_6241,N_7276);
nor U11732 (N_11732,N_8523,N_7595);
and U11733 (N_11733,N_8702,N_7440);
nand U11734 (N_11734,N_6188,N_8255);
nand U11735 (N_11735,N_8971,N_7329);
nand U11736 (N_11736,N_6609,N_6788);
nand U11737 (N_11737,N_6285,N_7536);
or U11738 (N_11738,N_6108,N_7701);
nor U11739 (N_11739,N_8317,N_8534);
nor U11740 (N_11740,N_6911,N_7374);
nand U11741 (N_11741,N_8574,N_8935);
nand U11742 (N_11742,N_7454,N_6652);
and U11743 (N_11743,N_7191,N_8858);
and U11744 (N_11744,N_8345,N_8490);
and U11745 (N_11745,N_6737,N_7990);
xor U11746 (N_11746,N_8151,N_8829);
and U11747 (N_11747,N_8864,N_7297);
or U11748 (N_11748,N_8970,N_7355);
and U11749 (N_11749,N_8360,N_6537);
nand U11750 (N_11750,N_8381,N_6417);
or U11751 (N_11751,N_7942,N_8664);
or U11752 (N_11752,N_7349,N_8478);
nor U11753 (N_11753,N_7301,N_7568);
and U11754 (N_11754,N_8876,N_7165);
nor U11755 (N_11755,N_7018,N_6791);
or U11756 (N_11756,N_6309,N_8197);
nand U11757 (N_11757,N_6788,N_7174);
nor U11758 (N_11758,N_7150,N_6145);
nor U11759 (N_11759,N_6884,N_6081);
or U11760 (N_11760,N_7741,N_6983);
or U11761 (N_11761,N_8354,N_8184);
or U11762 (N_11762,N_7614,N_6048);
nand U11763 (N_11763,N_7573,N_8085);
xnor U11764 (N_11764,N_8019,N_7837);
nor U11765 (N_11765,N_6878,N_8475);
and U11766 (N_11766,N_7781,N_6375);
nor U11767 (N_11767,N_6971,N_8028);
or U11768 (N_11768,N_6689,N_8408);
or U11769 (N_11769,N_8718,N_8638);
or U11770 (N_11770,N_6546,N_6869);
nand U11771 (N_11771,N_6393,N_7704);
nor U11772 (N_11772,N_8389,N_8328);
nor U11773 (N_11773,N_8218,N_7110);
or U11774 (N_11774,N_7692,N_8219);
nand U11775 (N_11775,N_8557,N_8696);
or U11776 (N_11776,N_8545,N_6328);
and U11777 (N_11777,N_8278,N_8575);
or U11778 (N_11778,N_8926,N_6831);
and U11779 (N_11779,N_8927,N_6033);
and U11780 (N_11780,N_8444,N_7103);
nand U11781 (N_11781,N_6520,N_8577);
nor U11782 (N_11782,N_8941,N_8208);
nand U11783 (N_11783,N_8321,N_8047);
and U11784 (N_11784,N_6825,N_6021);
or U11785 (N_11785,N_8720,N_7605);
nor U11786 (N_11786,N_7451,N_7199);
nor U11787 (N_11787,N_8253,N_8154);
or U11788 (N_11788,N_7849,N_8084);
or U11789 (N_11789,N_8244,N_8930);
nand U11790 (N_11790,N_8921,N_7629);
and U11791 (N_11791,N_6112,N_7807);
or U11792 (N_11792,N_7123,N_6984);
and U11793 (N_11793,N_6426,N_6945);
nor U11794 (N_11794,N_7815,N_8142);
nand U11795 (N_11795,N_6463,N_6926);
nor U11796 (N_11796,N_6374,N_7571);
and U11797 (N_11797,N_7041,N_8154);
and U11798 (N_11798,N_7870,N_7253);
nand U11799 (N_11799,N_7756,N_7282);
or U11800 (N_11800,N_8725,N_7542);
nand U11801 (N_11801,N_7008,N_8419);
and U11802 (N_11802,N_6012,N_7892);
and U11803 (N_11803,N_7898,N_7166);
nand U11804 (N_11804,N_6211,N_7722);
or U11805 (N_11805,N_7488,N_8929);
nor U11806 (N_11806,N_6702,N_6726);
nor U11807 (N_11807,N_8239,N_6651);
and U11808 (N_11808,N_6333,N_7096);
or U11809 (N_11809,N_8433,N_6774);
and U11810 (N_11810,N_6790,N_8869);
and U11811 (N_11811,N_7569,N_6530);
nand U11812 (N_11812,N_8319,N_7497);
nor U11813 (N_11813,N_6501,N_6887);
or U11814 (N_11814,N_8058,N_6059);
or U11815 (N_11815,N_7368,N_8782);
nor U11816 (N_11816,N_8843,N_6910);
nand U11817 (N_11817,N_7267,N_6218);
nor U11818 (N_11818,N_6530,N_8200);
or U11819 (N_11819,N_8450,N_7896);
or U11820 (N_11820,N_7170,N_6357);
nor U11821 (N_11821,N_8594,N_7893);
and U11822 (N_11822,N_7253,N_6332);
or U11823 (N_11823,N_6784,N_7015);
xor U11824 (N_11824,N_6021,N_6232);
nand U11825 (N_11825,N_6856,N_7877);
nor U11826 (N_11826,N_6410,N_7326);
and U11827 (N_11827,N_6550,N_8229);
or U11828 (N_11828,N_6919,N_8910);
or U11829 (N_11829,N_6392,N_6550);
or U11830 (N_11830,N_6307,N_8028);
nand U11831 (N_11831,N_8469,N_8275);
nor U11832 (N_11832,N_8936,N_6143);
xnor U11833 (N_11833,N_6757,N_6902);
or U11834 (N_11834,N_7940,N_8357);
nor U11835 (N_11835,N_7045,N_8841);
nor U11836 (N_11836,N_8084,N_7308);
or U11837 (N_11837,N_6881,N_8763);
nand U11838 (N_11838,N_8861,N_7527);
or U11839 (N_11839,N_7232,N_6492);
and U11840 (N_11840,N_6805,N_8428);
nor U11841 (N_11841,N_8532,N_6926);
nor U11842 (N_11842,N_6461,N_7977);
or U11843 (N_11843,N_6508,N_8335);
nand U11844 (N_11844,N_6929,N_6798);
and U11845 (N_11845,N_6433,N_6519);
nand U11846 (N_11846,N_8974,N_7485);
nand U11847 (N_11847,N_8967,N_8554);
or U11848 (N_11848,N_6402,N_6722);
nor U11849 (N_11849,N_6495,N_8002);
nand U11850 (N_11850,N_8180,N_7420);
or U11851 (N_11851,N_8850,N_8173);
nor U11852 (N_11852,N_6794,N_6549);
nand U11853 (N_11853,N_6883,N_6995);
and U11854 (N_11854,N_6755,N_6502);
nor U11855 (N_11855,N_6562,N_8643);
xnor U11856 (N_11856,N_8476,N_7165);
or U11857 (N_11857,N_8303,N_8370);
or U11858 (N_11858,N_6475,N_8352);
and U11859 (N_11859,N_7872,N_8242);
nor U11860 (N_11860,N_6943,N_8039);
nor U11861 (N_11861,N_8654,N_8859);
and U11862 (N_11862,N_6350,N_6049);
nand U11863 (N_11863,N_7579,N_7372);
or U11864 (N_11864,N_6249,N_7626);
and U11865 (N_11865,N_8109,N_6333);
nand U11866 (N_11866,N_6221,N_7074);
nor U11867 (N_11867,N_8211,N_7473);
nor U11868 (N_11868,N_7958,N_6846);
nor U11869 (N_11869,N_8151,N_6853);
nand U11870 (N_11870,N_6807,N_7397);
or U11871 (N_11871,N_7070,N_6310);
and U11872 (N_11872,N_6958,N_7914);
nor U11873 (N_11873,N_8042,N_7889);
xnor U11874 (N_11874,N_7482,N_6996);
and U11875 (N_11875,N_8039,N_6508);
and U11876 (N_11876,N_8437,N_7313);
or U11877 (N_11877,N_6032,N_8448);
or U11878 (N_11878,N_7934,N_7902);
and U11879 (N_11879,N_6977,N_7253);
and U11880 (N_11880,N_7878,N_6411);
and U11881 (N_11881,N_6234,N_7791);
nand U11882 (N_11882,N_8289,N_6508);
or U11883 (N_11883,N_7413,N_6465);
and U11884 (N_11884,N_6051,N_8694);
nand U11885 (N_11885,N_7557,N_8362);
or U11886 (N_11886,N_7170,N_8395);
and U11887 (N_11887,N_8815,N_8682);
or U11888 (N_11888,N_6412,N_6285);
or U11889 (N_11889,N_6386,N_7254);
nor U11890 (N_11890,N_7141,N_8921);
and U11891 (N_11891,N_6067,N_7848);
or U11892 (N_11892,N_6140,N_8145);
or U11893 (N_11893,N_8763,N_7161);
nor U11894 (N_11894,N_8238,N_6742);
or U11895 (N_11895,N_8726,N_8987);
nor U11896 (N_11896,N_8295,N_8312);
or U11897 (N_11897,N_6748,N_8632);
nor U11898 (N_11898,N_7595,N_7041);
and U11899 (N_11899,N_6126,N_7702);
and U11900 (N_11900,N_6194,N_8393);
and U11901 (N_11901,N_6772,N_8816);
and U11902 (N_11902,N_7428,N_6979);
and U11903 (N_11903,N_7972,N_6239);
nor U11904 (N_11904,N_7043,N_6420);
or U11905 (N_11905,N_6483,N_8629);
or U11906 (N_11906,N_7504,N_7220);
or U11907 (N_11907,N_8610,N_6941);
and U11908 (N_11908,N_8449,N_8304);
xnor U11909 (N_11909,N_7808,N_6444);
and U11910 (N_11910,N_8380,N_8675);
nor U11911 (N_11911,N_8642,N_8084);
xnor U11912 (N_11912,N_7450,N_6254);
nor U11913 (N_11913,N_8396,N_7064);
and U11914 (N_11914,N_6430,N_8096);
nand U11915 (N_11915,N_7512,N_6987);
nand U11916 (N_11916,N_7847,N_7215);
and U11917 (N_11917,N_7375,N_8538);
and U11918 (N_11918,N_7360,N_7642);
nor U11919 (N_11919,N_6997,N_8408);
and U11920 (N_11920,N_7586,N_6397);
and U11921 (N_11921,N_7844,N_8388);
nand U11922 (N_11922,N_7416,N_8975);
or U11923 (N_11923,N_8842,N_6306);
and U11924 (N_11924,N_8045,N_7044);
and U11925 (N_11925,N_6157,N_6908);
and U11926 (N_11926,N_6415,N_7157);
nor U11927 (N_11927,N_7207,N_6235);
and U11928 (N_11928,N_6768,N_6401);
nand U11929 (N_11929,N_7890,N_7147);
and U11930 (N_11930,N_6209,N_6308);
nor U11931 (N_11931,N_6798,N_7648);
nor U11932 (N_11932,N_8926,N_8076);
nand U11933 (N_11933,N_7806,N_8070);
nor U11934 (N_11934,N_8145,N_8915);
nand U11935 (N_11935,N_6335,N_6203);
nand U11936 (N_11936,N_8041,N_6178);
or U11937 (N_11937,N_7573,N_7054);
and U11938 (N_11938,N_7222,N_6044);
or U11939 (N_11939,N_8355,N_8352);
nor U11940 (N_11940,N_8798,N_6426);
and U11941 (N_11941,N_8959,N_7501);
nor U11942 (N_11942,N_7721,N_7469);
and U11943 (N_11943,N_6288,N_8062);
or U11944 (N_11944,N_7610,N_8918);
or U11945 (N_11945,N_8465,N_8128);
and U11946 (N_11946,N_6428,N_7271);
nand U11947 (N_11947,N_6647,N_7313);
nand U11948 (N_11948,N_8813,N_8314);
nor U11949 (N_11949,N_8422,N_6364);
and U11950 (N_11950,N_7909,N_7876);
nand U11951 (N_11951,N_7029,N_6332);
nor U11952 (N_11952,N_7065,N_6266);
nor U11953 (N_11953,N_8829,N_7236);
and U11954 (N_11954,N_7188,N_7530);
or U11955 (N_11955,N_6280,N_8999);
nor U11956 (N_11956,N_7127,N_6516);
nand U11957 (N_11957,N_6271,N_8765);
and U11958 (N_11958,N_8873,N_7042);
or U11959 (N_11959,N_7738,N_6286);
nor U11960 (N_11960,N_8059,N_7942);
nand U11961 (N_11961,N_6887,N_6874);
and U11962 (N_11962,N_7211,N_7516);
or U11963 (N_11963,N_7058,N_8940);
nand U11964 (N_11964,N_6839,N_7639);
nand U11965 (N_11965,N_6679,N_7733);
nor U11966 (N_11966,N_8154,N_6000);
nor U11967 (N_11967,N_8590,N_8715);
and U11968 (N_11968,N_8665,N_7920);
nand U11969 (N_11969,N_8241,N_6190);
or U11970 (N_11970,N_6260,N_8431);
nor U11971 (N_11971,N_8774,N_8980);
and U11972 (N_11972,N_7872,N_6104);
and U11973 (N_11973,N_6808,N_6219);
nor U11974 (N_11974,N_8540,N_8139);
and U11975 (N_11975,N_8176,N_6503);
nand U11976 (N_11976,N_7107,N_7593);
nor U11977 (N_11977,N_8505,N_7262);
and U11978 (N_11978,N_8248,N_6811);
nor U11979 (N_11979,N_6160,N_7449);
or U11980 (N_11980,N_8672,N_7800);
or U11981 (N_11981,N_8322,N_8978);
nand U11982 (N_11982,N_7589,N_6104);
or U11983 (N_11983,N_6712,N_6626);
and U11984 (N_11984,N_8152,N_7608);
nor U11985 (N_11985,N_8762,N_8244);
nor U11986 (N_11986,N_6365,N_8974);
or U11987 (N_11987,N_8311,N_6487);
and U11988 (N_11988,N_6951,N_6262);
or U11989 (N_11989,N_7168,N_8270);
nand U11990 (N_11990,N_8524,N_8903);
nor U11991 (N_11991,N_6276,N_8295);
nor U11992 (N_11992,N_6139,N_7961);
and U11993 (N_11993,N_6320,N_8877);
and U11994 (N_11994,N_8296,N_6230);
nor U11995 (N_11995,N_6763,N_7615);
nand U11996 (N_11996,N_7025,N_6435);
or U11997 (N_11997,N_7806,N_7375);
and U11998 (N_11998,N_8177,N_6570);
nor U11999 (N_11999,N_8271,N_8274);
nor U12000 (N_12000,N_9879,N_9687);
nand U12001 (N_12001,N_9431,N_9327);
or U12002 (N_12002,N_10321,N_10986);
or U12003 (N_12003,N_9456,N_11174);
nand U12004 (N_12004,N_10634,N_11786);
nor U12005 (N_12005,N_9516,N_11173);
nor U12006 (N_12006,N_11909,N_10237);
nor U12007 (N_12007,N_10094,N_9943);
nand U12008 (N_12008,N_11582,N_11103);
and U12009 (N_12009,N_11805,N_11009);
nor U12010 (N_12010,N_10254,N_10077);
nor U12011 (N_12011,N_9055,N_11339);
nor U12012 (N_12012,N_9486,N_10524);
and U12013 (N_12013,N_9519,N_9313);
or U12014 (N_12014,N_11350,N_11124);
nand U12015 (N_12015,N_11483,N_10633);
xor U12016 (N_12016,N_10338,N_10609);
and U12017 (N_12017,N_11808,N_10197);
or U12018 (N_12018,N_11361,N_11511);
nor U12019 (N_12019,N_9438,N_9822);
nor U12020 (N_12020,N_10411,N_11642);
or U12021 (N_12021,N_9471,N_10767);
nor U12022 (N_12022,N_10243,N_9742);
and U12023 (N_12023,N_10434,N_10643);
nor U12024 (N_12024,N_11370,N_11634);
and U12025 (N_12025,N_10562,N_10822);
or U12026 (N_12026,N_9900,N_10063);
nor U12027 (N_12027,N_10661,N_11331);
nand U12028 (N_12028,N_10070,N_11660);
and U12029 (N_12029,N_10660,N_10646);
nand U12030 (N_12030,N_10942,N_9326);
nand U12031 (N_12031,N_11600,N_10047);
or U12032 (N_12032,N_9235,N_11006);
and U12033 (N_12033,N_9083,N_9780);
or U12034 (N_12034,N_10966,N_11841);
nor U12035 (N_12035,N_10620,N_11054);
and U12036 (N_12036,N_11987,N_9772);
nor U12037 (N_12037,N_10506,N_10480);
and U12038 (N_12038,N_9854,N_10572);
nand U12039 (N_12039,N_11761,N_11056);
nor U12040 (N_12040,N_10097,N_9629);
and U12041 (N_12041,N_9549,N_11098);
nor U12042 (N_12042,N_11534,N_9881);
nand U12043 (N_12043,N_10744,N_9803);
or U12044 (N_12044,N_9414,N_11355);
and U12045 (N_12045,N_11668,N_11061);
and U12046 (N_12046,N_10726,N_10951);
and U12047 (N_12047,N_9913,N_11575);
or U12048 (N_12048,N_11209,N_9544);
xnor U12049 (N_12049,N_9116,N_11650);
nor U12050 (N_12050,N_11088,N_11547);
and U12051 (N_12051,N_11847,N_9617);
or U12052 (N_12052,N_10692,N_9616);
and U12053 (N_12053,N_9016,N_11425);
nand U12054 (N_12054,N_10812,N_10102);
nor U12055 (N_12055,N_10195,N_11110);
nor U12056 (N_12056,N_10912,N_10275);
nor U12057 (N_12057,N_11131,N_11423);
nand U12058 (N_12058,N_11401,N_10475);
and U12059 (N_12059,N_10785,N_9081);
nand U12060 (N_12060,N_11178,N_10946);
or U12061 (N_12061,N_10947,N_9265);
nand U12062 (N_12062,N_10140,N_11046);
or U12063 (N_12063,N_10561,N_10082);
nor U12064 (N_12064,N_9980,N_9305);
nor U12065 (N_12065,N_9672,N_10315);
or U12066 (N_12066,N_11719,N_10001);
and U12067 (N_12067,N_10843,N_9657);
nand U12068 (N_12068,N_11970,N_10302);
nand U12069 (N_12069,N_10326,N_11597);
nand U12070 (N_12070,N_10332,N_10239);
nand U12071 (N_12071,N_9426,N_9973);
nand U12072 (N_12072,N_9485,N_10439);
nand U12073 (N_12073,N_9407,N_10008);
nand U12074 (N_12074,N_10416,N_9206);
and U12075 (N_12075,N_9899,N_9790);
nor U12076 (N_12076,N_10152,N_11743);
and U12077 (N_12077,N_10603,N_11959);
and U12078 (N_12078,N_9513,N_9577);
or U12079 (N_12079,N_11280,N_9309);
and U12080 (N_12080,N_10975,N_9412);
or U12081 (N_12081,N_9948,N_11239);
nand U12082 (N_12082,N_11564,N_10380);
nor U12083 (N_12083,N_9766,N_10051);
or U12084 (N_12084,N_10161,N_10240);
nor U12085 (N_12085,N_9749,N_9977);
nand U12086 (N_12086,N_11321,N_10871);
or U12087 (N_12087,N_10349,N_9936);
nand U12088 (N_12088,N_11406,N_10878);
nor U12089 (N_12089,N_11151,N_11924);
nor U12090 (N_12090,N_11336,N_10473);
or U12091 (N_12091,N_11150,N_10399);
or U12092 (N_12092,N_9926,N_10917);
and U12093 (N_12093,N_11715,N_10788);
nand U12094 (N_12094,N_10700,N_10406);
nor U12095 (N_12095,N_11059,N_11857);
nand U12096 (N_12096,N_11894,N_9514);
nor U12097 (N_12097,N_10787,N_10347);
nor U12098 (N_12098,N_9022,N_9498);
nor U12099 (N_12099,N_11079,N_9808);
nor U12100 (N_12100,N_11722,N_9415);
and U12101 (N_12101,N_10096,N_10832);
nor U12102 (N_12102,N_10987,N_10731);
and U12103 (N_12103,N_10432,N_10605);
nand U12104 (N_12104,N_11739,N_9110);
or U12105 (N_12105,N_11115,N_9376);
and U12106 (N_12106,N_11246,N_10223);
or U12107 (N_12107,N_10782,N_11016);
and U12108 (N_12108,N_9205,N_10374);
and U12109 (N_12109,N_10022,N_9996);
and U12110 (N_12110,N_10383,N_9666);
or U12111 (N_12111,N_10547,N_10387);
nand U12112 (N_12112,N_11943,N_9272);
or U12113 (N_12113,N_11821,N_9994);
nor U12114 (N_12114,N_10106,N_11343);
nor U12115 (N_12115,N_10027,N_10429);
nand U12116 (N_12116,N_11696,N_11029);
and U12117 (N_12117,N_10895,N_11412);
and U12118 (N_12118,N_10104,N_10724);
nor U12119 (N_12119,N_10033,N_10886);
or U12120 (N_12120,N_9574,N_11864);
nand U12121 (N_12121,N_11887,N_10486);
nand U12122 (N_12122,N_9032,N_10068);
or U12123 (N_12123,N_11671,N_9448);
nor U12124 (N_12124,N_11153,N_10482);
nor U12125 (N_12125,N_10962,N_10307);
nand U12126 (N_12126,N_10453,N_10158);
nand U12127 (N_12127,N_10867,N_9257);
nand U12128 (N_12128,N_11207,N_10805);
nor U12129 (N_12129,N_10510,N_10126);
nand U12130 (N_12130,N_10215,N_11094);
and U12131 (N_12131,N_9964,N_10575);
xor U12132 (N_12132,N_11421,N_11745);
xor U12133 (N_12133,N_10924,N_11787);
or U12134 (N_12134,N_9774,N_10893);
nor U12135 (N_12135,N_9354,N_11905);
nand U12136 (N_12136,N_9944,N_11028);
nor U12137 (N_12137,N_9453,N_9756);
and U12138 (N_12138,N_11530,N_10284);
and U12139 (N_12139,N_9566,N_10194);
and U12140 (N_12140,N_9348,N_9674);
nor U12141 (N_12141,N_9271,N_9655);
nand U12142 (N_12142,N_9966,N_10378);
nand U12143 (N_12143,N_11895,N_11141);
or U12144 (N_12144,N_11914,N_11138);
nand U12145 (N_12145,N_10877,N_9374);
and U12146 (N_12146,N_9583,N_11477);
or U12147 (N_12147,N_9129,N_10764);
nor U12148 (N_12148,N_10268,N_9564);
nor U12149 (N_12149,N_11220,N_11972);
nor U12150 (N_12150,N_10755,N_9166);
or U12151 (N_12151,N_10998,N_11275);
or U12152 (N_12152,N_10178,N_10896);
and U12153 (N_12153,N_11169,N_10566);
nor U12154 (N_12154,N_10918,N_11128);
and U12155 (N_12155,N_11297,N_9299);
nor U12156 (N_12156,N_9955,N_9730);
xnor U12157 (N_12157,N_11121,N_9044);
nor U12158 (N_12158,N_11033,N_10624);
nor U12159 (N_12159,N_10515,N_10931);
or U12160 (N_12160,N_9723,N_9889);
nor U12161 (N_12161,N_9860,N_10250);
nor U12162 (N_12162,N_9394,N_9193);
or U12163 (N_12163,N_9492,N_11766);
and U12164 (N_12164,N_11086,N_11942);
and U12165 (N_12165,N_11049,N_11814);
or U12166 (N_12166,N_9745,N_9204);
xor U12167 (N_12167,N_10184,N_9705);
nor U12168 (N_12168,N_10181,N_10090);
nor U12169 (N_12169,N_11828,N_10211);
or U12170 (N_12170,N_9455,N_11404);
nor U12171 (N_12171,N_10465,N_10469);
or U12172 (N_12172,N_10028,N_11922);
nand U12173 (N_12173,N_9027,N_9894);
or U12174 (N_12174,N_10631,N_9863);
nor U12175 (N_12175,N_11224,N_10167);
nor U12176 (N_12176,N_11728,N_9283);
or U12177 (N_12177,N_11353,N_9421);
or U12178 (N_12178,N_11565,N_11699);
or U12179 (N_12179,N_9760,N_11946);
nor U12180 (N_12180,N_10638,N_11441);
and U12181 (N_12181,N_11409,N_11560);
nor U12182 (N_12182,N_11837,N_11559);
or U12183 (N_12183,N_10682,N_10021);
and U12184 (N_12184,N_9619,N_10351);
nand U12185 (N_12185,N_9535,N_10578);
or U12186 (N_12186,N_9097,N_10906);
or U12187 (N_12187,N_11609,N_10421);
nor U12188 (N_12188,N_9782,N_11395);
and U12189 (N_12189,N_9364,N_10990);
and U12190 (N_12190,N_10498,N_11741);
nor U12191 (N_12191,N_10288,N_11988);
nand U12192 (N_12192,N_9965,N_10289);
nand U12193 (N_12193,N_11304,N_9707);
or U12194 (N_12194,N_11114,N_11688);
nand U12195 (N_12195,N_9754,N_9626);
nand U12196 (N_12196,N_10176,N_10521);
and U12197 (N_12197,N_9391,N_11136);
and U12198 (N_12198,N_9495,N_10120);
and U12199 (N_12199,N_11817,N_10839);
and U12200 (N_12200,N_11455,N_9458);
nand U12201 (N_12201,N_11538,N_9428);
nor U12202 (N_12202,N_10736,N_11371);
nor U12203 (N_12203,N_10442,N_10031);
nand U12204 (N_12204,N_10334,N_10775);
nor U12205 (N_12205,N_10717,N_11993);
or U12206 (N_12206,N_11859,N_10807);
xnor U12207 (N_12207,N_11615,N_9114);
nand U12208 (N_12208,N_10697,N_11241);
and U12209 (N_12209,N_9999,N_9531);
or U12210 (N_12210,N_11063,N_9388);
or U12211 (N_12211,N_10776,N_11545);
nand U12212 (N_12212,N_11189,N_9623);
and U12213 (N_12213,N_11936,N_10391);
and U12214 (N_12214,N_11505,N_11288);
or U12215 (N_12215,N_9014,N_9615);
nand U12216 (N_12216,N_10777,N_10298);
and U12217 (N_12217,N_10647,N_9238);
nor U12218 (N_12218,N_9991,N_9484);
or U12219 (N_12219,N_9245,N_10907);
and U12220 (N_12220,N_9783,N_10901);
xor U12221 (N_12221,N_11374,N_10013);
and U12222 (N_12222,N_11032,N_10367);
and U12223 (N_12223,N_11208,N_11249);
or U12224 (N_12224,N_11091,N_9988);
or U12225 (N_12225,N_11733,N_9041);
nor U12226 (N_12226,N_11271,N_9671);
or U12227 (N_12227,N_10702,N_11397);
nand U12228 (N_12228,N_10122,N_11995);
and U12229 (N_12229,N_10596,N_9285);
or U12230 (N_12230,N_11272,N_10314);
nand U12231 (N_12231,N_9843,N_10039);
or U12232 (N_12232,N_10143,N_10230);
or U12233 (N_12233,N_10023,N_10329);
and U12234 (N_12234,N_11704,N_10061);
nand U12235 (N_12235,N_9154,N_11104);
nor U12236 (N_12236,N_10982,N_9897);
and U12237 (N_12237,N_9775,N_11667);
or U12238 (N_12238,N_11473,N_9013);
nand U12239 (N_12239,N_10888,N_11517);
nor U12240 (N_12240,N_11258,N_10679);
or U12241 (N_12241,N_10758,N_11148);
and U12242 (N_12242,N_10585,N_11497);
or U12243 (N_12243,N_10086,N_9602);
nor U12244 (N_12244,N_11282,N_10558);
or U12245 (N_12245,N_11955,N_9989);
nor U12246 (N_12246,N_9332,N_9054);
nor U12247 (N_12247,N_10870,N_11751);
and U12248 (N_12248,N_10535,N_10430);
nand U12249 (N_12249,N_11164,N_9761);
and U12250 (N_12250,N_10554,N_11171);
nor U12251 (N_12251,N_10500,N_9825);
nor U12252 (N_12252,N_9620,N_9532);
xnor U12253 (N_12253,N_11427,N_9281);
xnor U12254 (N_12254,N_9815,N_10376);
nand U12255 (N_12255,N_11961,N_10529);
and U12256 (N_12256,N_11315,N_10231);
nor U12257 (N_12257,N_10247,N_11450);
and U12258 (N_12258,N_11259,N_11903);
nor U12259 (N_12259,N_9470,N_10306);
xnor U12260 (N_12260,N_9115,N_9941);
nor U12261 (N_12261,N_11415,N_11599);
nor U12262 (N_12262,N_9931,N_9890);
nand U12263 (N_12263,N_9306,N_11608);
and U12264 (N_12264,N_10659,N_11165);
nor U12265 (N_12265,N_9476,N_9785);
nand U12266 (N_12266,N_10060,N_10485);
nor U12267 (N_12267,N_9318,N_10623);
or U12268 (N_12268,N_10447,N_11829);
and U12269 (N_12269,N_11064,N_10712);
nand U12270 (N_12270,N_11992,N_9106);
nor U12271 (N_12271,N_10227,N_11802);
or U12272 (N_12272,N_10502,N_11456);
nand U12273 (N_12273,N_9466,N_11812);
nor U12274 (N_12274,N_10831,N_10825);
or U12275 (N_12275,N_11702,N_11556);
and U12276 (N_12276,N_10007,N_10046);
or U12277 (N_12277,N_9356,N_11698);
and U12278 (N_12278,N_10581,N_11644);
nand U12279 (N_12279,N_10369,N_10048);
and U12280 (N_12280,N_10478,N_11732);
or U12281 (N_12281,N_10135,N_11738);
nor U12282 (N_12282,N_9869,N_10188);
nand U12283 (N_12283,N_11013,N_9915);
and U12284 (N_12284,N_11206,N_10204);
or U12285 (N_12285,N_11533,N_10327);
nand U12286 (N_12286,N_11623,N_11269);
nand U12287 (N_12287,N_10273,N_11655);
nor U12288 (N_12288,N_10412,N_9315);
nor U12289 (N_12289,N_9827,N_9888);
nand U12290 (N_12290,N_9700,N_9680);
nor U12291 (N_12291,N_10331,N_10674);
or U12292 (N_12292,N_11622,N_9568);
nand U12293 (N_12293,N_11537,N_11880);
or U12294 (N_12294,N_9224,N_9263);
and U12295 (N_12295,N_11347,N_10860);
nand U12296 (N_12296,N_9107,N_9868);
nor U12297 (N_12297,N_9248,N_11080);
nand U12298 (N_12298,N_9777,N_10846);
and U12299 (N_12299,N_11758,N_9928);
or U12300 (N_12300,N_9643,N_9231);
or U12301 (N_12301,N_9270,N_10333);
or U12302 (N_12302,N_9339,N_11492);
nor U12303 (N_12303,N_10622,N_10770);
or U12304 (N_12304,N_10248,N_9160);
nand U12305 (N_12305,N_11183,N_10256);
nor U12306 (N_12306,N_11769,N_9759);
nor U12307 (N_12307,N_10803,N_10538);
nand U12308 (N_12308,N_10219,N_9451);
or U12309 (N_12309,N_10516,N_9430);
nand U12310 (N_12310,N_9140,N_9161);
nand U12311 (N_12311,N_10342,N_11281);
and U12312 (N_12312,N_11662,N_10481);
and U12313 (N_12313,N_10232,N_11482);
or U12314 (N_12314,N_11503,N_11678);
xor U12315 (N_12315,N_9025,N_9064);
nor U12316 (N_12316,N_9738,N_9149);
or U12317 (N_12317,N_11603,N_11154);
or U12318 (N_12318,N_10363,N_9082);
nor U12319 (N_12319,N_9462,N_9904);
nand U12320 (N_12320,N_9813,N_9935);
or U12321 (N_12321,N_9523,N_11749);
nor U12322 (N_12322,N_9793,N_9891);
nand U12323 (N_12323,N_9480,N_10164);
nand U12324 (N_12324,N_11883,N_11300);
or U12325 (N_12325,N_10718,N_11057);
or U12326 (N_12326,N_10260,N_10423);
and U12327 (N_12327,N_10355,N_10295);
and U12328 (N_12328,N_11294,N_9251);
nor U12329 (N_12329,N_10956,N_11949);
or U12330 (N_12330,N_11991,N_11767);
nor U12331 (N_12331,N_10385,N_11921);
nand U12332 (N_12332,N_11167,N_11014);
nor U12333 (N_12333,N_9427,N_11161);
nor U12334 (N_12334,N_10397,N_10626);
or U12335 (N_12335,N_9938,N_9912);
nand U12336 (N_12336,N_11755,N_9320);
nand U12337 (N_12337,N_10372,N_9087);
or U12338 (N_12338,N_9651,N_9658);
nand U12339 (N_12339,N_10824,N_11038);
and U12340 (N_12340,N_11351,N_11398);
nor U12341 (N_12341,N_11686,N_10533);
or U12342 (N_12342,N_11481,N_9791);
and U12343 (N_12343,N_10542,N_10282);
nand U12344 (N_12344,N_9088,N_11390);
or U12345 (N_12345,N_10271,N_10983);
or U12346 (N_12346,N_11043,N_9393);
nand U12347 (N_12347,N_9233,N_11528);
nor U12348 (N_12348,N_11957,N_9956);
nand U12349 (N_12349,N_11192,N_10029);
and U12350 (N_12350,N_9859,N_10848);
nand U12351 (N_12351,N_9512,N_10041);
or U12352 (N_12352,N_11777,N_10503);
and U12353 (N_12353,N_11915,N_9419);
nor U12354 (N_12354,N_11015,N_11886);
and U12355 (N_12355,N_10760,N_10715);
or U12356 (N_12356,N_10226,N_9978);
nor U12357 (N_12357,N_9108,N_11865);
and U12358 (N_12358,N_9916,N_9138);
or U12359 (N_12359,N_11944,N_11568);
xor U12360 (N_12360,N_9609,N_9136);
nor U12361 (N_12361,N_9012,N_9042);
nand U12362 (N_12362,N_11718,N_10588);
and U12363 (N_12363,N_10277,N_9570);
and U12364 (N_12364,N_10491,N_11679);
nor U12365 (N_12365,N_9886,N_10970);
and U12366 (N_12366,N_9131,N_10793);
or U12367 (N_12367,N_10759,N_9555);
nand U12368 (N_12368,N_10435,N_11384);
nand U12369 (N_12369,N_11140,N_11793);
or U12370 (N_12370,N_11352,N_11203);
nor U12371 (N_12371,N_9223,N_10228);
or U12372 (N_12372,N_10939,N_11020);
or U12373 (N_12373,N_11264,N_9563);
nand U12374 (N_12374,N_11884,N_10991);
and U12375 (N_12375,N_10873,N_11897);
and U12376 (N_12376,N_10213,N_11625);
nor U12377 (N_12377,N_9538,N_11523);
and U12378 (N_12378,N_11782,N_10114);
or U12379 (N_12379,N_9024,N_11930);
and U12380 (N_12380,N_9719,N_9494);
nand U12381 (N_12381,N_9578,N_11437);
or U12382 (N_12382,N_9557,N_9591);
nand U12383 (N_12383,N_10111,N_10085);
and U12384 (N_12384,N_10173,N_11799);
nor U12385 (N_12385,N_10599,N_9817);
nor U12386 (N_12386,N_11796,N_10016);
or U12387 (N_12387,N_11024,N_10708);
or U12388 (N_12388,N_11595,N_11022);
and U12389 (N_12389,N_9870,N_10015);
nand U12390 (N_12390,N_9856,N_9954);
and U12391 (N_12391,N_9792,N_11794);
or U12392 (N_12392,N_11647,N_10706);
xnor U12393 (N_12393,N_9007,N_9947);
xnor U12394 (N_12394,N_11939,N_9392);
nor U12395 (N_12395,N_10899,N_10714);
and U12396 (N_12396,N_10501,N_11484);
or U12397 (N_12397,N_11506,N_9961);
nand U12398 (N_12398,N_9652,N_9969);
nand U12399 (N_12399,N_9622,N_9344);
nor U12400 (N_12400,N_11781,N_9840);
nor U12401 (N_12401,N_9144,N_9942);
and U12402 (N_12402,N_11596,N_11325);
nand U12403 (N_12403,N_10317,N_9001);
and U12404 (N_12404,N_10841,N_10612);
nor U12405 (N_12405,N_9066,N_11163);
nand U12406 (N_12406,N_9545,N_10748);
nand U12407 (N_12407,N_9755,N_9331);
nor U12408 (N_12408,N_9011,N_11519);
nand U12409 (N_12409,N_9992,N_10150);
nor U12410 (N_12410,N_9684,N_9352);
or U12411 (N_12411,N_11156,N_10261);
or U12412 (N_12412,N_10107,N_11290);
nand U12413 (N_12413,N_9797,N_11179);
xnor U12414 (N_12414,N_9614,N_10636);
nand U12415 (N_12415,N_10595,N_11475);
nor U12416 (N_12416,N_10433,N_10162);
nand U12417 (N_12417,N_9002,N_11866);
or U12418 (N_12418,N_9968,N_11095);
or U12419 (N_12419,N_11457,N_11377);
or U12420 (N_12420,N_10328,N_10997);
and U12421 (N_12421,N_10794,N_9148);
and U12422 (N_12422,N_9214,N_11166);
nand U12423 (N_12423,N_11674,N_11092);
nand U12424 (N_12424,N_11730,N_9252);
and U12425 (N_12425,N_9259,N_10461);
nand U12426 (N_12426,N_10032,N_10009);
nand U12427 (N_12427,N_10600,N_11432);
nand U12428 (N_12428,N_11212,N_10766);
or U12429 (N_12429,N_11573,N_10003);
nor U12430 (N_12430,N_11862,N_9565);
and U12431 (N_12431,N_11487,N_9185);
or U12432 (N_12432,N_9420,N_10673);
or U12433 (N_12433,N_9752,N_10680);
and U12434 (N_12434,N_10098,N_11932);
nand U12435 (N_12435,N_10263,N_9917);
or U12436 (N_12436,N_10088,N_10677);
nand U12437 (N_12437,N_10004,N_11222);
and U12438 (N_12438,N_9125,N_11462);
or U12439 (N_12439,N_9821,N_9794);
and U12440 (N_12440,N_11919,N_10817);
and U12441 (N_12441,N_11298,N_11843);
or U12442 (N_12442,N_11577,N_10151);
nand U12443 (N_12443,N_9333,N_10894);
xnor U12444 (N_12444,N_10402,N_11804);
nand U12445 (N_12445,N_10574,N_9158);
and U12446 (N_12446,N_9924,N_9585);
and U12447 (N_12447,N_9902,N_11792);
nand U12448 (N_12448,N_11607,N_11130);
nand U12449 (N_12449,N_11428,N_9122);
nor U12450 (N_12450,N_10444,N_9225);
nor U12451 (N_12451,N_9338,N_11904);
xor U12452 (N_12452,N_11947,N_11586);
nor U12453 (N_12453,N_10185,N_10577);
nand U12454 (N_12454,N_9475,N_10186);
and U12455 (N_12455,N_11368,N_11611);
or U12456 (N_12456,N_11504,N_11231);
nor U12457 (N_12457,N_10395,N_11724);
and U12458 (N_12458,N_11387,N_10459);
nor U12459 (N_12459,N_9950,N_11283);
or U12460 (N_12460,N_11011,N_11399);
or U12461 (N_12461,N_11574,N_10683);
or U12462 (N_12462,N_10701,N_11639);
and U12463 (N_12463,N_9449,N_10570);
nand U12464 (N_12464,N_9998,N_11005);
nand U12465 (N_12465,N_9668,N_9748);
and U12466 (N_12466,N_9173,N_11834);
nand U12467 (N_12467,N_10927,N_10310);
or U12468 (N_12468,N_10941,N_9811);
and U12469 (N_12469,N_10532,N_11122);
nand U12470 (N_12470,N_11145,N_9972);
or U12471 (N_12471,N_9734,N_11319);
or U12472 (N_12472,N_10669,N_10080);
or U12473 (N_12473,N_11149,N_9500);
nor U12474 (N_12474,N_10093,N_10555);
nand U12475 (N_12475,N_10691,N_9037);
or U12476 (N_12476,N_10354,N_10610);
and U12477 (N_12477,N_9706,N_10468);
nor U12478 (N_12478,N_9120,N_10519);
nor U12479 (N_12479,N_9653,N_10583);
nor U12480 (N_12480,N_10020,N_11007);
and U12481 (N_12481,N_10466,N_11635);
or U12482 (N_12482,N_9764,N_10458);
nand U12483 (N_12483,N_11881,N_9182);
and U12484 (N_12484,N_10280,N_10089);
nand U12485 (N_12485,N_10119,N_9239);
or U12486 (N_12486,N_10103,N_10840);
nand U12487 (N_12487,N_10483,N_9660);
or U12488 (N_12488,N_10407,N_9939);
nor U12489 (N_12489,N_11693,N_10336);
nor U12490 (N_12490,N_9312,N_10508);
or U12491 (N_12491,N_9727,N_10649);
and U12492 (N_12492,N_11845,N_11388);
or U12493 (N_12493,N_11809,N_10069);
and U12494 (N_12494,N_10722,N_9409);
nand U12495 (N_12495,N_11438,N_9307);
nand U12496 (N_12496,N_9111,N_10961);
or U12497 (N_12497,N_10055,N_11567);
and U12498 (N_12498,N_10916,N_11967);
nand U12499 (N_12499,N_10786,N_11190);
or U12500 (N_12500,N_9117,N_9515);
nand U12501 (N_12501,N_11495,N_9543);
or U12502 (N_12502,N_11176,N_9905);
or U12503 (N_12503,N_11612,N_11030);
or U12504 (N_12504,N_10976,N_11583);
nand U12505 (N_12505,N_9799,N_10553);
or U12506 (N_12506,N_11590,N_10505);
xnor U12507 (N_12507,N_9625,N_11513);
nand U12508 (N_12508,N_9946,N_11797);
or U12509 (N_12509,N_11261,N_11775);
or U12510 (N_12510,N_9028,N_9184);
nand U12511 (N_12511,N_11413,N_11302);
and U12512 (N_12512,N_9683,N_11594);
nand U12513 (N_12513,N_9167,N_9855);
nand U12514 (N_12514,N_10062,N_9696);
nand U12515 (N_12515,N_9714,N_9147);
nand U12516 (N_12516,N_11367,N_11966);
or U12517 (N_12517,N_11822,N_10614);
or U12518 (N_12518,N_9862,N_11507);
or U12519 (N_12519,N_9411,N_11587);
and U12520 (N_12520,N_9118,N_11187);
or U12521 (N_12521,N_11048,N_11172);
nand U12522 (N_12522,N_9096,N_11754);
and U12523 (N_12523,N_9035,N_9324);
nor U12524 (N_12524,N_9885,N_9406);
or U12525 (N_12525,N_11213,N_9276);
and U12526 (N_12526,N_9221,N_11296);
nand U12527 (N_12527,N_9925,N_9778);
nor U12528 (N_12528,N_9883,N_9250);
or U12529 (N_12529,N_9321,N_9624);
nor U12530 (N_12530,N_9858,N_11443);
or U12531 (N_12531,N_11251,N_11133);
xor U12532 (N_12532,N_10156,N_11381);
and U12533 (N_12533,N_11690,N_10417);
or U12534 (N_12534,N_10221,N_9378);
xor U12535 (N_12535,N_10118,N_11132);
xor U12536 (N_12536,N_10012,N_9914);
nor U12537 (N_12537,N_9715,N_11839);
nor U12538 (N_12538,N_11531,N_11096);
or U12539 (N_12539,N_11788,N_11453);
xor U12540 (N_12540,N_11899,N_11344);
nor U12541 (N_12541,N_11543,N_11958);
and U12542 (N_12542,N_10606,N_9553);
and U12543 (N_12543,N_11789,N_10765);
and U12544 (N_12544,N_10389,N_9153);
and U12545 (N_12545,N_9501,N_11807);
nand U12546 (N_12546,N_11823,N_10590);
and U12547 (N_12547,N_9253,N_9901);
or U12548 (N_12548,N_9403,N_10174);
and U12549 (N_12549,N_11476,N_9758);
nand U12550 (N_12550,N_10484,N_9310);
nor U12551 (N_12551,N_9170,N_10244);
nor U12552 (N_12552,N_10926,N_9076);
or U12553 (N_12553,N_9311,N_9690);
or U12554 (N_12554,N_10441,N_11731);
or U12555 (N_12555,N_11012,N_11451);
or U12556 (N_12556,N_9508,N_10305);
nor U12557 (N_12557,N_11465,N_11638);
or U12558 (N_12558,N_9442,N_10949);
or U12559 (N_12559,N_10863,N_10179);
or U12560 (N_12560,N_9844,N_11784);
and U12561 (N_12561,N_11860,N_10005);
nand U12562 (N_12562,N_10541,N_9552);
and U12563 (N_12563,N_11593,N_9308);
nand U12564 (N_12564,N_10981,N_10892);
or U12565 (N_12565,N_11760,N_11771);
and U12566 (N_12566,N_10160,N_10801);
nand U12567 (N_12567,N_9175,N_11137);
nor U12568 (N_12568,N_10564,N_9139);
and U12569 (N_12569,N_11727,N_11257);
or U12570 (N_12570,N_10437,N_10685);
nor U12571 (N_12571,N_10064,N_11997);
nor U12572 (N_12572,N_11950,N_10258);
nor U12573 (N_12573,N_11123,N_11037);
or U12574 (N_12574,N_9000,N_10980);
nand U12575 (N_12575,N_9983,N_9360);
nor U12576 (N_12576,N_9604,N_9478);
nand U12577 (N_12577,N_11018,N_10663);
nor U12578 (N_12578,N_10408,N_9588);
nor U12579 (N_12579,N_9744,N_11286);
and U12580 (N_12580,N_10847,N_9298);
nor U12581 (N_12581,N_10865,N_10136);
and U12582 (N_12582,N_10445,N_10903);
nor U12583 (N_12583,N_11783,N_11996);
and U12584 (N_12584,N_9551,N_9030);
nor U12585 (N_12585,N_11408,N_10364);
and U12586 (N_12586,N_9075,N_9521);
and U12587 (N_12587,N_9861,N_11309);
and U12588 (N_12588,N_10789,N_9864);
and U12589 (N_12589,N_11478,N_9260);
or U12590 (N_12590,N_11610,N_9273);
nand U12591 (N_12591,N_9729,N_10448);
nor U12592 (N_12592,N_9425,N_9788);
or U12593 (N_12593,N_11661,N_11411);
or U12594 (N_12594,N_11585,N_11083);
nand U12595 (N_12595,N_10768,N_9005);
nor U12596 (N_12596,N_11580,N_10324);
nor U12597 (N_12597,N_9046,N_11488);
nand U12598 (N_12598,N_10592,N_11791);
nor U12599 (N_12599,N_9342,N_11848);
xor U12600 (N_12600,N_9192,N_11876);
nor U12601 (N_12601,N_10798,N_11357);
nand U12602 (N_12602,N_9607,N_9819);
nor U12603 (N_12603,N_9569,N_11333);
and U12604 (N_12604,N_11287,N_10955);
nand U12605 (N_12605,N_11230,N_11237);
nor U12606 (N_12606,N_11393,N_9085);
and U12607 (N_12607,N_11736,N_10117);
nand U12608 (N_12608,N_10658,N_11752);
or U12609 (N_12609,N_9787,N_10881);
nand U12610 (N_12610,N_10550,N_10146);
nor U12611 (N_12611,N_10455,N_11579);
or U12612 (N_12612,N_9613,N_11349);
nand U12613 (N_12613,N_9921,N_9866);
and U12614 (N_12614,N_9667,N_10637);
nand U12615 (N_12615,N_9932,N_10311);
nand U12616 (N_12616,N_9801,N_11216);
nor U12617 (N_12617,N_9728,N_9317);
nand U12618 (N_12618,N_9194,N_9839);
and U12619 (N_12619,N_9853,N_9264);
nor U12620 (N_12620,N_9079,N_9586);
nand U12621 (N_12621,N_11403,N_11320);
nand U12622 (N_12622,N_9547,N_11896);
nand U12623 (N_12623,N_11326,N_11078);
or U12624 (N_12624,N_11981,N_9390);
or U12625 (N_12625,N_10169,N_10934);
nand U12626 (N_12626,N_11026,N_11877);
or U12627 (N_12627,N_9481,N_11602);
or U12628 (N_12628,N_11553,N_10889);
or U12629 (N_12629,N_10940,N_11186);
nor U12630 (N_12630,N_10656,N_10616);
nand U12631 (N_12631,N_10316,N_9196);
nand U12632 (N_12632,N_10772,N_10779);
nand U12633 (N_12633,N_9058,N_11979);
and U12634 (N_12634,N_10496,N_9807);
xor U12635 (N_12635,N_10619,N_10576);
or U12636 (N_12636,N_10175,N_11614);
or U12637 (N_12637,N_9168,N_10897);
nor U12638 (N_12638,N_11926,N_9605);
nand U12639 (N_12639,N_11641,N_10642);
or U12640 (N_12640,N_10390,N_10450);
nand U12641 (N_12641,N_11725,N_9023);
and U12642 (N_12642,N_10276,N_10115);
and U12643 (N_12643,N_9036,N_11770);
nor U12644 (N_12644,N_9191,N_9447);
and U12645 (N_12645,N_10727,N_9618);
or U12646 (N_12646,N_11912,N_11618);
and U12647 (N_12647,N_11620,N_10290);
nor U12648 (N_12648,N_10989,N_11158);
nand U12649 (N_12649,N_10121,N_11328);
nor U12650 (N_12650,N_9650,N_9268);
and U12651 (N_12651,N_11116,N_10203);
or U12652 (N_12652,N_9370,N_11496);
xnor U12653 (N_12653,N_11708,N_9489);
or U12654 (N_12654,N_9057,N_10937);
nor U12655 (N_12655,N_11363,N_10000);
and U12656 (N_12656,N_9997,N_10083);
or U12657 (N_12657,N_9896,N_10413);
and U12658 (N_12658,N_11021,N_9109);
and U12659 (N_12659,N_10038,N_10303);
nor U12660 (N_12660,N_11458,N_11819);
or U12661 (N_12661,N_10291,N_9491);
nand U12662 (N_12662,N_9382,N_11692);
and U12663 (N_12663,N_11075,N_10246);
nor U12664 (N_12664,N_11081,N_11306);
or U12665 (N_12665,N_11806,N_10965);
xor U12666 (N_12666,N_11461,N_9496);
and U12667 (N_12667,N_9849,N_11735);
nor U12668 (N_12668,N_9600,N_9599);
or U12669 (N_12669,N_10436,N_9546);
or U12670 (N_12670,N_11687,N_10866);
nand U12671 (N_12671,N_11836,N_9506);
nor U12672 (N_12672,N_10740,N_11314);
nor U12673 (N_12673,N_11196,N_9689);
and U12674 (N_12674,N_11923,N_9806);
nor U12675 (N_12675,N_9127,N_11117);
and U12676 (N_12676,N_9450,N_11968);
and U12677 (N_12677,N_11572,N_9662);
nand U12678 (N_12678,N_9210,N_10464);
nand U12679 (N_12679,N_11844,N_10493);
and U12680 (N_12680,N_9343,N_11076);
xnor U12681 (N_12681,N_9459,N_11654);
nor U12682 (N_12682,N_11027,N_9026);
or U12683 (N_12683,N_11723,N_10341);
and U12684 (N_12684,N_11778,N_9369);
nand U12685 (N_12685,N_11247,N_10147);
nand U12686 (N_12686,N_11071,N_9725);
nor U12687 (N_12687,N_11700,N_11774);
and U12688 (N_12688,N_10632,N_9798);
nand U12689 (N_12689,N_11194,N_11375);
nand U12690 (N_12690,N_9677,N_9611);
and U12691 (N_12691,N_9047,N_9113);
or U12692 (N_12692,N_10419,N_9934);
and U12693 (N_12693,N_9757,N_9830);
or U12694 (N_12694,N_9644,N_9334);
nand U12695 (N_12695,N_11311,N_9560);
nor U12696 (N_12696,N_9804,N_9654);
nor U12697 (N_12697,N_9699,N_10272);
nor U12698 (N_12698,N_9836,N_9335);
nor U12699 (N_12699,N_10954,N_10418);
nor U12700 (N_12700,N_9424,N_10137);
or U12701 (N_12701,N_11376,N_11065);
nor U12702 (N_12702,N_9610,N_11780);
or U12703 (N_12703,N_10944,N_10780);
nand U12704 (N_12704,N_11498,N_10806);
nor U12705 (N_12705,N_10675,N_9156);
and U12706 (N_12706,N_9102,N_11980);
nand U12707 (N_12707,N_9872,N_10795);
nand U12708 (N_12708,N_10887,N_9929);
nor U12709 (N_12709,N_10344,N_10325);
nor U12710 (N_12710,N_11539,N_11764);
nand U12711 (N_12711,N_11816,N_11720);
nand U12712 (N_12712,N_10218,N_10769);
and U12713 (N_12713,N_10153,N_10720);
or U12714 (N_12714,N_11566,N_11493);
nor U12715 (N_12715,N_9465,N_11680);
and U12716 (N_12716,N_11292,N_10196);
and U12717 (N_12717,N_11303,N_9630);
and U12718 (N_12718,N_9893,N_11433);
nand U12719 (N_12719,N_11868,N_11740);
nor U12720 (N_12720,N_11418,N_11204);
and U12721 (N_12721,N_11299,N_10630);
or U12722 (N_12722,N_11389,N_10409);
and U12723 (N_12723,N_9608,N_11470);
nand U12724 (N_12724,N_9119,N_9034);
and U12725 (N_12725,N_9242,N_10388);
or U12726 (N_12726,N_9355,N_10905);
and U12727 (N_12727,N_10075,N_10792);
nand U12728 (N_12728,N_11019,N_9584);
or U12729 (N_12729,N_9077,N_9303);
nand U12730 (N_12730,N_10312,N_10811);
nand U12731 (N_12731,N_9919,N_11500);
or U12732 (N_12732,N_10995,N_9637);
or U12733 (N_12733,N_11416,N_9851);
nor U12734 (N_12734,N_10902,N_10953);
and U12735 (N_12735,N_10474,N_11185);
or U12736 (N_12736,N_11323,N_9779);
or U12737 (N_12737,N_9052,N_11274);
or U12738 (N_12738,N_9053,N_9895);
or U12739 (N_12739,N_10144,N_10573);
nor U12740 (N_12740,N_9733,N_11228);
and U12741 (N_12741,N_11874,N_9207);
nor U12742 (N_12742,N_9290,N_11795);
or U12743 (N_12743,N_11305,N_11626);
nand U12744 (N_12744,N_11527,N_10133);
nor U12745 (N_12745,N_9123,N_10651);
nor U12746 (N_12746,N_9045,N_10791);
or U12747 (N_12747,N_9291,N_9445);
and U12748 (N_12748,N_11295,N_10177);
and U12749 (N_12749,N_10754,N_11756);
nor U12750 (N_12750,N_11134,N_11223);
nor U12751 (N_12751,N_10668,N_10883);
nand U12752 (N_12752,N_10264,N_9554);
nand U12753 (N_12753,N_9282,N_9739);
and U12754 (N_12754,N_11750,N_11677);
or U12755 (N_12755,N_10495,N_11546);
and U12756 (N_12756,N_10006,N_11147);
or U12757 (N_12757,N_10763,N_11360);
or U12758 (N_12758,N_11840,N_11721);
nand U12759 (N_12759,N_9048,N_11126);
and U12760 (N_12760,N_10838,N_9401);
nor U12761 (N_12761,N_11605,N_9810);
and U12762 (N_12762,N_10259,N_10019);
nor U12763 (N_12763,N_11990,N_11928);
or U12764 (N_12764,N_11265,N_11985);
or U12765 (N_12765,N_10762,N_9222);
or U12766 (N_12766,N_10978,N_10704);
or U12767 (N_12767,N_9389,N_10270);
and U12768 (N_12768,N_9151,N_11815);
nor U12769 (N_12769,N_11480,N_10932);
or U12770 (N_12770,N_9460,N_11270);
or U12771 (N_12771,N_11069,N_11501);
nand U12772 (N_12772,N_10800,N_11938);
nand U12773 (N_12773,N_9537,N_11430);
nand U12774 (N_12774,N_10224,N_9441);
nor U12775 (N_12775,N_11717,N_9824);
nor U12776 (N_12776,N_9132,N_9384);
nand U12777 (N_12777,N_11542,N_11108);
and U12778 (N_12778,N_9562,N_10569);
or U12779 (N_12779,N_10492,N_10322);
and U12780 (N_12780,N_11571,N_9632);
nand U12781 (N_12781,N_10149,N_9202);
and U12782 (N_12782,N_11113,N_11637);
nor U12783 (N_12783,N_11446,N_11440);
nand U12784 (N_12784,N_9417,N_11047);
nand U12785 (N_12785,N_9638,N_10823);
and U12786 (N_12786,N_9266,N_11978);
and U12787 (N_12787,N_10142,N_11199);
nor U12788 (N_12788,N_11025,N_9918);
nor U12789 (N_12789,N_11162,N_10362);
nor U12790 (N_12790,N_11628,N_9021);
and U12791 (N_12791,N_9820,N_11486);
or U12792 (N_12792,N_9789,N_9981);
nand U12793 (N_12793,N_10830,N_10654);
or U12794 (N_12794,N_10499,N_11676);
nor U12795 (N_12795,N_9006,N_9301);
nand U12796 (N_12796,N_10725,N_11444);
nor U12797 (N_12797,N_11691,N_9446);
nor U12798 (N_12798,N_10640,N_11541);
nand U12799 (N_12799,N_10862,N_9361);
and U12800 (N_12800,N_10814,N_10913);
nand U12801 (N_12801,N_9784,N_10035);
or U12802 (N_12802,N_11034,N_9892);
nand U12803 (N_12803,N_9678,N_10681);
nand U12804 (N_12804,N_11479,N_10065);
nor U12805 (N_12805,N_11491,N_10403);
and U12806 (N_12806,N_9726,N_9165);
and U12807 (N_12807,N_10415,N_10283);
nor U12808 (N_12808,N_11512,N_10375);
or U12809 (N_12809,N_10734,N_10353);
nor U12810 (N_12810,N_9716,N_10166);
and U12811 (N_12811,N_10220,N_11552);
nand U12812 (N_12812,N_9940,N_11729);
xnor U12813 (N_12813,N_10025,N_9256);
and U12814 (N_12814,N_9040,N_10134);
or U12815 (N_12815,N_10828,N_11826);
nor U12816 (N_12816,N_11892,N_11392);
or U12817 (N_12817,N_10826,N_10552);
and U12818 (N_12818,N_11442,N_11613);
nand U12819 (N_12819,N_9254,N_11616);
and U12820 (N_12820,N_10836,N_10462);
or U12821 (N_12821,N_11157,N_9112);
nor U12822 (N_12822,N_11332,N_9673);
or U12823 (N_12823,N_10262,N_11869);
or U12824 (N_12824,N_9509,N_11445);
nor U12825 (N_12825,N_9061,N_11256);
and U12826 (N_12826,N_11159,N_10963);
nand U12827 (N_12827,N_10292,N_11589);
nand U12828 (N_12828,N_9062,N_10930);
nor U12829 (N_12829,N_10414,N_10757);
nor U12830 (N_12830,N_10479,N_9556);
and U12831 (N_12831,N_10876,N_11245);
nor U12832 (N_12832,N_9596,N_10778);
nand U12833 (N_12833,N_9641,N_9145);
nor U12834 (N_12834,N_10379,N_10108);
and U12835 (N_12835,N_11146,N_10011);
nor U12836 (N_12836,N_10750,N_11604);
and U12837 (N_12837,N_11524,N_11318);
xnor U12838 (N_12838,N_10737,N_10530);
nor U12839 (N_12839,N_10551,N_9186);
nand U12840 (N_12840,N_9567,N_10868);
or U12841 (N_12841,N_9350,N_10582);
or U12842 (N_12842,N_11858,N_9200);
and U12843 (N_12843,N_9226,N_10512);
and U12844 (N_12844,N_10365,N_11913);
nor U12845 (N_12845,N_9358,N_9951);
nor U12846 (N_12846,N_9155,N_11901);
nor U12847 (N_12847,N_10885,N_10829);
nor U12848 (N_12848,N_10921,N_11563);
or U12849 (N_12849,N_9953,N_9261);
nor U12850 (N_12850,N_9753,N_10943);
nand U12851 (N_12851,N_10968,N_9621);
and U12852 (N_12852,N_10132,N_9633);
and U12853 (N_12853,N_9050,N_9142);
nor U12854 (N_12854,N_10320,N_10431);
nand U12855 (N_12855,N_9488,N_9212);
or U12856 (N_12856,N_9970,N_11422);
nor U12857 (N_12857,N_10579,N_11643);
nand U12858 (N_12858,N_10743,N_10170);
and U12859 (N_12859,N_11665,N_9187);
nor U12860 (N_12860,N_10155,N_9209);
nor U12861 (N_12861,N_9710,N_11229);
nand U12862 (N_12862,N_10050,N_10716);
nand U12863 (N_12863,N_9435,N_11198);
or U12864 (N_12864,N_9345,N_10190);
nor U12865 (N_12865,N_11989,N_11291);
nor U12866 (N_12866,N_10586,N_10650);
nor U12867 (N_12867,N_11983,N_9906);
and U12868 (N_12868,N_9249,N_10490);
nor U12869 (N_12869,N_11555,N_11042);
or U12870 (N_12870,N_10816,N_11976);
and U12871 (N_12871,N_9211,N_10200);
and U12872 (N_12872,N_9550,N_9300);
nor U12873 (N_12873,N_9960,N_11842);
nor U12874 (N_12874,N_11279,N_10568);
nor U12875 (N_12875,N_10255,N_11601);
nor U12876 (N_12876,N_10589,N_9418);
nor U12877 (N_12877,N_10689,N_11951);
or U12878 (N_12878,N_9400,N_9070);
nand U12879 (N_12879,N_9769,N_10818);
and U12880 (N_12880,N_10676,N_11109);
and U12881 (N_12881,N_9367,N_10460);
nor U12882 (N_12882,N_10253,N_11810);
nor U12883 (N_12883,N_9319,N_11431);
or U12884 (N_12884,N_11039,N_9682);
and U12885 (N_12885,N_10368,N_10854);
or U12886 (N_12886,N_11278,N_10183);
nor U12887 (N_12887,N_11773,N_10371);
and U12888 (N_12888,N_11459,N_9464);
and U12889 (N_12889,N_10945,N_11640);
or U12890 (N_12890,N_10517,N_10923);
nand U12891 (N_12891,N_10091,N_11139);
nor U12892 (N_12892,N_11925,N_10294);
nor U12893 (N_12893,N_10545,N_10815);
nor U12894 (N_12894,N_11310,N_11920);
nand U12895 (N_12895,N_9008,N_10182);
or U12896 (N_12896,N_11648,N_11873);
nand U12897 (N_12897,N_10130,N_10556);
or U12898 (N_12898,N_11518,N_9086);
nand U12899 (N_12899,N_10597,N_9439);
or U12900 (N_12900,N_10935,N_9540);
or U12901 (N_12901,N_10957,N_9910);
nand U12902 (N_12902,N_9247,N_11221);
or U12903 (N_12903,N_9490,N_11152);
nor U12904 (N_12904,N_10148,N_11882);
nand U12905 (N_12905,N_10773,N_11818);
nand U12906 (N_12906,N_11646,N_9126);
and U12907 (N_12907,N_11975,N_11346);
nand U12908 (N_12908,N_10381,N_11734);
or U12909 (N_12909,N_11973,N_11621);
nor U12910 (N_12910,N_10904,N_10799);
nand U12911 (N_12911,N_9104,N_10487);
nor U12912 (N_12912,N_10753,N_11945);
nor U12913 (N_12913,N_10652,N_9838);
or U12914 (N_12914,N_9218,N_10074);
and U12915 (N_12915,N_9594,N_9592);
and U12916 (N_12916,N_9199,N_9229);
and U12917 (N_12917,N_9735,N_9876);
nand U12918 (N_12918,N_10925,N_11373);
or U12919 (N_12919,N_9230,N_10452);
nor U12920 (N_12920,N_11036,N_11127);
nor U12921 (N_12921,N_9669,N_9559);
nor U12922 (N_12922,N_10404,N_11889);
nor U12923 (N_12923,N_11263,N_9635);
nand U12924 (N_12924,N_10690,N_11701);
nand U12925 (N_12925,N_9510,N_9874);
nand U12926 (N_12926,N_9482,N_9169);
nand U12927 (N_12927,N_9341,N_9704);
nor U12928 (N_12928,N_10611,N_10037);
nor U12929 (N_12929,N_9718,N_10971);
and U12930 (N_12930,N_9038,N_9911);
nand U12931 (N_12931,N_11863,N_9020);
xnor U12932 (N_12932,N_10699,N_9241);
and U12933 (N_12933,N_11998,N_10587);
and U12934 (N_12934,N_10996,N_9080);
xor U12935 (N_12935,N_11402,N_11830);
and U12936 (N_12936,N_11253,N_9100);
or U12937 (N_12937,N_9959,N_10125);
nor U12938 (N_12938,N_10977,N_10285);
or U12939 (N_12939,N_10861,N_11685);
or U12940 (N_12940,N_9487,N_11112);
and U12941 (N_12941,N_11345,N_11378);
and U12942 (N_12942,N_10522,N_11210);
nand U12943 (N_12943,N_11017,N_9511);
nor U12944 (N_12944,N_9015,N_10973);
nor U12945 (N_12945,N_11472,N_11474);
or U12946 (N_12946,N_10598,N_11910);
nor U12947 (N_12947,N_9033,N_9805);
nor U12948 (N_12948,N_11090,N_11753);
nand U12949 (N_12949,N_9809,N_11969);
and U12950 (N_12950,N_10979,N_11277);
and U12951 (N_12951,N_11673,N_11562);
xor U12952 (N_12952,N_9135,N_11188);
and U12953 (N_12953,N_10615,N_9986);
and U12954 (N_12954,N_10056,N_11898);
or U12955 (N_12955,N_11629,N_9987);
or U12956 (N_12956,N_9380,N_9737);
and U12957 (N_12957,N_10756,N_10339);
nand U12958 (N_12958,N_9743,N_10110);
nor U12959 (N_12959,N_9090,N_11856);
nor U12960 (N_12960,N_9434,N_10859);
nand U12961 (N_12961,N_9975,N_11193);
and U12962 (N_12962,N_10844,N_9497);
and U12963 (N_12963,N_10472,N_10127);
nand U12964 (N_12964,N_10154,N_10426);
nor U12965 (N_12965,N_11651,N_9072);
and U12966 (N_12966,N_10703,N_10463);
nand U12967 (N_12967,N_10053,N_11803);
nor U12968 (N_12968,N_11561,N_11243);
or U12969 (N_12969,N_10992,N_11301);
nor U12970 (N_12970,N_9386,N_9213);
or U12971 (N_12971,N_11831,N_11664);
nand U12972 (N_12972,N_9573,N_9875);
nor U12973 (N_12973,N_11205,N_9558);
and U12974 (N_12974,N_10688,N_9141);
and U12975 (N_12975,N_10410,N_9029);
and U12976 (N_12976,N_11707,N_11737);
and U12977 (N_12977,N_9217,N_11578);
and U12978 (N_12978,N_9593,N_10476);
nor U12979 (N_12979,N_10443,N_9898);
nor U12980 (N_12980,N_9984,N_10858);
and U12981 (N_12981,N_11885,N_9304);
or U12982 (N_12982,N_9065,N_10972);
nand U12983 (N_12983,N_9353,N_10201);
nand U12984 (N_12984,N_11746,N_11879);
nor U12985 (N_12985,N_9952,N_11170);
or U12986 (N_12986,N_9945,N_10042);
or U12987 (N_12987,N_11135,N_11073);
or U12988 (N_12988,N_11835,N_11948);
or U12989 (N_12989,N_9606,N_10950);
and U12990 (N_12990,N_9074,N_10489);
or U12991 (N_12991,N_10030,N_11790);
and U12992 (N_12992,N_10257,N_11581);
nand U12993 (N_12993,N_10810,N_11394);
nand U12994 (N_12994,N_9404,N_10066);
nor U12995 (N_12995,N_11584,N_11000);
or U12996 (N_12996,N_10879,N_10428);
or U12997 (N_12997,N_11324,N_9004);
and U12998 (N_12998,N_11916,N_11284);
or U12999 (N_12999,N_10054,N_9781);
nor U13000 (N_13000,N_11327,N_10300);
or U13001 (N_13001,N_10357,N_11522);
nand U13002 (N_13002,N_10225,N_11359);
or U13003 (N_13003,N_9457,N_9387);
and U13004 (N_13004,N_9373,N_10105);
and U13005 (N_13005,N_10297,N_9878);
and U13006 (N_13006,N_11362,N_10710);
and U13007 (N_13007,N_10319,N_10079);
nor U13008 (N_13008,N_10217,N_11293);
and U13009 (N_13009,N_10869,N_9314);
or U13010 (N_13010,N_10293,N_9685);
nor U13011 (N_13011,N_9831,N_9681);
or U13012 (N_13012,N_10109,N_11004);
and U13013 (N_13013,N_9698,N_11952);
nand U13014 (N_13014,N_10198,N_11931);
nor U13015 (N_13015,N_10711,N_9645);
nor U13016 (N_13016,N_9597,N_11045);
nor U13017 (N_13017,N_10959,N_9258);
nor U13018 (N_13018,N_11499,N_9220);
and U13019 (N_13019,N_10856,N_9068);
nand U13020 (N_13020,N_9473,N_9049);
or U13021 (N_13021,N_10067,N_10898);
and U13022 (N_13022,N_10567,N_9293);
nor U13023 (N_13023,N_9771,N_11619);
or U13024 (N_13024,N_9405,N_11669);
nand U13025 (N_13025,N_11762,N_9768);
or U13026 (N_13026,N_10797,N_10138);
nand U13027 (N_13027,N_9236,N_11342);
nor U13028 (N_13028,N_9410,N_11521);
or U13029 (N_13029,N_10813,N_9818);
xor U13030 (N_13030,N_10543,N_11744);
nor U13031 (N_13031,N_11954,N_11436);
and U13032 (N_13032,N_9463,N_9329);
xnor U13033 (N_13033,N_9800,N_9347);
nor U13034 (N_13034,N_9503,N_9575);
and U13035 (N_13035,N_11569,N_9847);
nor U13036 (N_13036,N_9436,N_9796);
xnor U13037 (N_13037,N_9093,N_11055);
and U13038 (N_13038,N_9958,N_9284);
nand U13039 (N_13039,N_10309,N_9648);
and U13040 (N_13040,N_9397,N_10608);
nand U13041 (N_13041,N_10629,N_11235);
nor U13042 (N_13042,N_9527,N_10208);
nor U13043 (N_13043,N_10299,N_11195);
nor U13044 (N_13044,N_11435,N_10348);
nand U13045 (N_13045,N_11001,N_10527);
nand U13046 (N_13046,N_10693,N_11893);
or U13047 (N_13047,N_9340,N_9871);
and U13048 (N_13048,N_9091,N_10279);
and U13049 (N_13049,N_9323,N_11372);
or U13050 (N_13050,N_9325,N_10168);
xnor U13051 (N_13051,N_9152,N_10187);
or U13052 (N_13052,N_11525,N_9773);
and U13053 (N_13053,N_10666,N_10471);
or U13054 (N_13054,N_9802,N_9433);
nor U13055 (N_13055,N_10116,N_10123);
nand U13056 (N_13056,N_11890,N_11653);
or U13057 (N_13057,N_9413,N_10191);
nor U13058 (N_13058,N_9534,N_10113);
or U13059 (N_13059,N_11878,N_10171);
and U13060 (N_13060,N_9089,N_11902);
nand U13061 (N_13061,N_9679,N_9437);
or U13062 (N_13062,N_9395,N_10808);
nand U13063 (N_13063,N_9071,N_11058);
or U13064 (N_13064,N_11941,N_11697);
xnor U13065 (N_13065,N_10405,N_11316);
or U13066 (N_13066,N_9228,N_9732);
or U13067 (N_13067,N_10422,N_11268);
nand U13068 (N_13068,N_10400,N_11663);
and U13069 (N_13069,N_10653,N_10286);
and U13070 (N_13070,N_9278,N_11776);
and U13071 (N_13071,N_10994,N_11380);
and U13072 (N_13072,N_10513,N_11097);
nor U13073 (N_13073,N_9279,N_11420);
and U13074 (N_13074,N_9703,N_9479);
and U13075 (N_13075,N_11536,N_9219);
nand U13076 (N_13076,N_9985,N_9069);
and U13077 (N_13077,N_10014,N_10449);
nor U13078 (N_13078,N_11820,N_9084);
or U13079 (N_13079,N_11872,N_10920);
or U13080 (N_13080,N_9659,N_11074);
nor U13081 (N_13081,N_11937,N_11077);
nand U13082 (N_13082,N_9740,N_11801);
xor U13083 (N_13083,N_9381,N_10559);
and U13084 (N_13084,N_10783,N_9177);
nand U13085 (N_13085,N_10911,N_11448);
nand U13086 (N_13086,N_9454,N_11329);
or U13087 (N_13087,N_9909,N_11354);
xnor U13088 (N_13088,N_10984,N_9443);
or U13089 (N_13089,N_11986,N_9670);
and U13090 (N_13090,N_11548,N_11386);
and U13091 (N_13091,N_11649,N_9852);
or U13092 (N_13092,N_9833,N_9665);
and U13093 (N_13093,N_10330,N_9067);
and U13094 (N_13094,N_11520,N_9372);
xor U13095 (N_13095,N_10337,N_10095);
nand U13096 (N_13096,N_9150,N_10733);
or U13097 (N_13097,N_9688,N_10591);
and U13098 (N_13098,N_9603,N_10518);
or U13099 (N_13099,N_11364,N_9143);
and U13100 (N_13100,N_11041,N_9383);
or U13101 (N_13101,N_10601,N_9159);
nor U13102 (N_13102,N_11144,N_11908);
nand U13103 (N_13103,N_11260,N_10855);
or U13104 (N_13104,N_11549,N_11215);
or U13105 (N_13105,N_10394,N_9365);
nand U13106 (N_13106,N_10141,N_10296);
nor U13107 (N_13107,N_10802,N_10594);
nor U13108 (N_13108,N_11391,N_11956);
nor U13109 (N_13109,N_9877,N_10560);
nor U13110 (N_13110,N_10157,N_11267);
or U13111 (N_13111,N_9828,N_10864);
nand U13112 (N_13112,N_10281,N_11464);
and U13113 (N_13113,N_10985,N_9043);
or U13114 (N_13114,N_11191,N_11529);
nor U13115 (N_13115,N_9472,N_10936);
xnor U13116 (N_13116,N_9098,N_11285);
nand U13117 (N_13117,N_9073,N_11825);
or U13118 (N_13118,N_11748,N_10242);
and U13119 (N_13119,N_10199,N_11852);
or U13120 (N_13120,N_11439,N_11100);
and U13121 (N_13121,N_11652,N_11008);
or U13122 (N_13122,N_10235,N_9302);
or U13123 (N_13123,N_11656,N_9366);
and U13124 (N_13124,N_9408,N_10900);
and U13125 (N_13125,N_10245,N_9349);
and U13126 (N_13126,N_11494,N_9377);
or U13127 (N_13127,N_11051,N_11485);
nand U13128 (N_13128,N_11636,N_9767);
nand U13129 (N_13129,N_9422,N_11348);
nand U13130 (N_13130,N_11526,N_11340);
and U13131 (N_13131,N_9157,N_9694);
nand U13132 (N_13132,N_9101,N_10644);
nand U13133 (N_13133,N_11953,N_9628);
nand U13134 (N_13134,N_11515,N_10967);
xor U13135 (N_13135,N_10952,N_11120);
nor U13136 (N_13136,N_9274,N_9524);
nor U13137 (N_13137,N_11846,N_11417);
xnor U13138 (N_13138,N_10988,N_11225);
nor U13139 (N_13139,N_11592,N_9507);
nor U13140 (N_13140,N_10335,N_11125);
nand U13141 (N_13141,N_10358,N_9884);
nand U13142 (N_13142,N_10964,N_9171);
or U13143 (N_13143,N_9103,N_11105);
nand U13144 (N_13144,N_10343,N_11107);
nor U13145 (N_13145,N_9533,N_10745);
or U13146 (N_13146,N_9724,N_9656);
nand U13147 (N_13147,N_9873,N_9363);
and U13148 (N_13148,N_10446,N_10323);
nand U13149 (N_13149,N_10241,N_11694);
nand U13150 (N_13150,N_11236,N_11711);
and U13151 (N_13151,N_9693,N_11250);
nand U13152 (N_13152,N_10546,N_10851);
nand U13153 (N_13153,N_9469,N_10593);
and U13154 (N_13154,N_11870,N_9018);
nor U13155 (N_13155,N_11657,N_10398);
or U13156 (N_13156,N_10267,N_10751);
nand U13157 (N_13157,N_11168,N_11960);
or U13158 (N_13158,N_11219,N_10618);
or U13159 (N_13159,N_10909,N_9502);
and U13160 (N_13160,N_11060,N_9432);
and U13161 (N_13161,N_11252,N_10129);
nor U13162 (N_13162,N_11532,N_10457);
or U13163 (N_13163,N_10738,N_9612);
nand U13164 (N_13164,N_11466,N_10210);
and U13165 (N_13165,N_10052,N_11143);
or U13166 (N_13166,N_11813,N_9832);
or U13167 (N_13167,N_10392,N_10092);
nor U13168 (N_13168,N_9640,N_11449);
xor U13169 (N_13169,N_11757,N_10124);
and U13170 (N_13170,N_10507,N_10370);
and U13171 (N_13171,N_11935,N_9094);
nand U13172 (N_13172,N_9636,N_9499);
and U13173 (N_13173,N_10278,N_11832);
or U13174 (N_13174,N_11118,N_10002);
or U13175 (N_13175,N_11489,N_10072);
nand U13176 (N_13176,N_11197,N_9776);
and U13177 (N_13177,N_9232,N_10820);
or U13178 (N_13178,N_11742,N_10948);
nor U13179 (N_13179,N_10308,N_11871);
nand U13180 (N_13180,N_9930,N_11454);
and U13181 (N_13181,N_9541,N_9051);
or U13182 (N_13182,N_9240,N_9721);
nand U13183 (N_13183,N_10837,N_11632);
nor U13184 (N_13184,N_9467,N_9188);
or U13185 (N_13185,N_11984,N_9009);
nor U13186 (N_13186,N_11160,N_10874);
or U13187 (N_13187,N_11102,N_9841);
and U13188 (N_13188,N_9702,N_9691);
and U13189 (N_13189,N_10373,N_11085);
and U13190 (N_13190,N_9017,N_11713);
nand U13191 (N_13191,N_10781,N_9751);
nor U13192 (N_13192,N_10233,N_10269);
or U13193 (N_13193,N_9137,N_11452);
nand U13194 (N_13194,N_10099,N_10884);
and U13195 (N_13195,N_9857,N_11709);
and U13196 (N_13196,N_10999,N_9539);
nor U13197 (N_13197,N_11356,N_11779);
and U13198 (N_13198,N_10627,N_11414);
nor U13199 (N_13199,N_10960,N_11933);
nand U13200 (N_13200,N_11684,N_10655);
and U13201 (N_13201,N_9572,N_11927);
or U13202 (N_13202,N_10514,N_11544);
nand U13203 (N_13203,N_10382,N_10229);
nor U13204 (N_13204,N_11226,N_11218);
nor U13205 (N_13205,N_9461,N_10670);
xnor U13206 (N_13206,N_9571,N_9227);
or U13207 (N_13207,N_11851,N_10835);
xor U13208 (N_13208,N_10018,N_10488);
nor U13209 (N_13209,N_11142,N_9267);
and U13210 (N_13210,N_11977,N_10352);
nand U13211 (N_13211,N_10548,N_9203);
nor U13212 (N_13212,N_9850,N_10087);
and U13213 (N_13213,N_9316,N_9505);
or U13214 (N_13214,N_9795,N_10922);
nor U13215 (N_13215,N_11234,N_11330);
or U13216 (N_13216,N_9741,N_9697);
and U13217 (N_13217,N_9368,N_11358);
nor U13218 (N_13218,N_10993,N_11426);
or U13219 (N_13219,N_9371,N_10207);
nand U13220 (N_13220,N_11906,N_10933);
nor U13221 (N_13221,N_10076,N_10974);
nand U13222 (N_13222,N_9396,N_9134);
nand U13223 (N_13223,N_10890,N_11369);
and U13224 (N_13224,N_11308,N_11824);
or U13225 (N_13225,N_9525,N_9190);
nand U13226 (N_13226,N_10396,N_11467);
nand U13227 (N_13227,N_10180,N_9292);
nand U13228 (N_13228,N_11365,N_9351);
or U13229 (N_13229,N_10908,N_9288);
and U13230 (N_13230,N_11867,N_9979);
nand U13231 (N_13231,N_11429,N_11338);
nand U13232 (N_13232,N_10440,N_11714);
nor U13233 (N_13233,N_11510,N_10628);
nor U13234 (N_13234,N_10425,N_10384);
nand U13235 (N_13235,N_11214,N_9598);
and U13236 (N_13236,N_9887,N_10340);
or U13237 (N_13237,N_11516,N_9949);
nor U13238 (N_13238,N_9520,N_10058);
and U13239 (N_13239,N_11312,N_11682);
or U13240 (N_13240,N_11598,N_11200);
nor U13241 (N_13241,N_9504,N_10880);
or U13242 (N_13242,N_9736,N_10915);
and U13243 (N_13243,N_10036,N_11627);
nand U13244 (N_13244,N_9908,N_9440);
nor U13245 (N_13245,N_10723,N_10318);
nor U13246 (N_13246,N_9581,N_9816);
or U13247 (N_13247,N_11624,N_11888);
nand U13248 (N_13248,N_9059,N_10266);
nor U13249 (N_13249,N_10774,N_11276);
nor U13250 (N_13250,N_9181,N_9162);
nor U13251 (N_13251,N_10845,N_11535);
and U13252 (N_13252,N_9712,N_11266);
nor U13253 (N_13253,N_9183,N_10827);
or U13254 (N_13254,N_10602,N_9483);
nor U13255 (N_13255,N_10128,N_11811);
and U13256 (N_13256,N_11383,N_9195);
and U13257 (N_13257,N_9328,N_9060);
or U13258 (N_13258,N_9105,N_10071);
or U13259 (N_13259,N_11407,N_11558);
nor U13260 (N_13260,N_9933,N_9337);
nor U13261 (N_13261,N_9092,N_11182);
nor U13262 (N_13262,N_11035,N_11747);
nand U13263 (N_13263,N_11509,N_9937);
or U13264 (N_13264,N_11551,N_11471);
nand U13265 (N_13265,N_9812,N_9234);
and U13266 (N_13266,N_9429,N_11672);
and U13267 (N_13267,N_11999,N_10705);
or U13268 (N_13268,N_9750,N_9330);
nand U13269 (N_13269,N_9770,N_11289);
and U13270 (N_13270,N_10833,N_9296);
and U13271 (N_13271,N_9542,N_9518);
nand U13272 (N_13272,N_10101,N_11658);
and U13273 (N_13273,N_9995,N_10427);
nand U13274 (N_13274,N_11469,N_11854);
nand U13275 (N_13275,N_11502,N_10928);
nor U13276 (N_13276,N_11082,N_9146);
and U13277 (N_13277,N_9375,N_10969);
or U13278 (N_13278,N_11490,N_10891);
nor U13279 (N_13279,N_9189,N_10034);
and U13280 (N_13280,N_9579,N_9846);
and U13281 (N_13281,N_9398,N_9528);
nand U13282 (N_13282,N_11337,N_11974);
nand U13283 (N_13283,N_11099,N_10857);
nand U13284 (N_13284,N_10834,N_9526);
or U13285 (N_13285,N_10205,N_10209);
nand U13286 (N_13286,N_11084,N_9920);
nor U13287 (N_13287,N_11710,N_11341);
and U13288 (N_13288,N_11833,N_11119);
nand U13289 (N_13289,N_9561,N_11010);
or U13290 (N_13290,N_11907,N_11111);
or U13291 (N_13291,N_9468,N_9837);
and U13292 (N_13292,N_9346,N_11785);
or U13293 (N_13293,N_9957,N_10057);
nand U13294 (N_13294,N_9922,N_11576);
and U13295 (N_13295,N_9180,N_9661);
nor U13296 (N_13296,N_11087,N_11716);
and U13297 (N_13297,N_10694,N_10252);
nand U13298 (N_13298,N_10451,N_9163);
nand U13299 (N_13299,N_10084,N_10687);
or U13300 (N_13300,N_10100,N_10635);
nor U13301 (N_13301,N_10531,N_10454);
or U13302 (N_13302,N_10043,N_11175);
or U13303 (N_13303,N_10707,N_9237);
nand U13304 (N_13304,N_9176,N_9208);
or U13305 (N_13305,N_10536,N_11155);
nand U13306 (N_13306,N_9589,N_9130);
nand U13307 (N_13307,N_9976,N_9845);
or U13308 (N_13308,N_11911,N_9517);
nand U13309 (N_13309,N_9197,N_11023);
or U13310 (N_13310,N_11262,N_10584);
or U13311 (N_13311,N_11964,N_11670);
or U13312 (N_13312,N_11066,N_9201);
and U13313 (N_13313,N_10523,N_10350);
nor U13314 (N_13314,N_10919,N_11468);
or U13315 (N_13315,N_11062,N_10265);
and U13316 (N_13316,N_9907,N_11689);
nand U13317 (N_13317,N_10749,N_9379);
or U13318 (N_13318,N_10719,N_10345);
and U13319 (N_13319,N_9747,N_11703);
nor U13320 (N_13320,N_11093,N_9786);
nand U13321 (N_13321,N_9982,N_10206);
or U13322 (N_13322,N_10796,N_11800);
nand U13323 (N_13323,N_9990,N_10438);
or U13324 (N_13324,N_11588,N_11307);
nor U13325 (N_13325,N_9336,N_11633);
or U13326 (N_13326,N_9003,N_9536);
nand U13327 (N_13327,N_11447,N_9720);
or U13328 (N_13328,N_11849,N_11248);
nand U13329 (N_13329,N_9695,N_10872);
and U13330 (N_13330,N_10509,N_10735);
or U13331 (N_13331,N_11002,N_10684);
nor U13332 (N_13332,N_9692,N_11463);
and U13333 (N_13333,N_10165,N_11050);
nor U13334 (N_13334,N_11962,N_9099);
and U13335 (N_13335,N_9286,N_9010);
xor U13336 (N_13336,N_11254,N_11317);
nor U13337 (N_13337,N_11630,N_10721);
and U13338 (N_13338,N_10809,N_11217);
or U13339 (N_13339,N_9423,N_10604);
or U13340 (N_13340,N_11106,N_9548);
nor U13341 (N_13341,N_10356,N_9923);
or U13342 (N_13342,N_10456,N_9880);
nor U13343 (N_13343,N_10504,N_9595);
nor U13344 (N_13344,N_11242,N_9709);
nor U13345 (N_13345,N_11554,N_10732);
nor U13346 (N_13346,N_10709,N_9746);
nand U13347 (N_13347,N_9708,N_9601);
nor U13348 (N_13348,N_11434,N_10672);
xor U13349 (N_13349,N_10112,N_11233);
or U13350 (N_13350,N_11918,N_10664);
and U13351 (N_13351,N_10761,N_10159);
or U13352 (N_13352,N_11550,N_9444);
nor U13353 (N_13353,N_10819,N_10842);
and U13354 (N_13354,N_10741,N_11366);
or U13355 (N_13355,N_9385,N_11681);
nor U13356 (N_13356,N_10366,N_10557);
nor U13357 (N_13357,N_10539,N_10665);
nand U13358 (N_13358,N_10301,N_10565);
or U13359 (N_13359,N_11712,N_10549);
or U13360 (N_13360,N_11177,N_11068);
nor U13361 (N_13361,N_9322,N_11273);
and U13362 (N_13362,N_11211,N_11695);
nand U13363 (N_13363,N_10625,N_10617);
and U13364 (N_13364,N_10359,N_10049);
nand U13365 (N_13365,N_10875,N_11683);
and U13366 (N_13366,N_9277,N_10742);
and U13367 (N_13367,N_9722,N_9246);
nor U13368 (N_13368,N_11424,N_9814);
and U13369 (N_13369,N_11855,N_10424);
or U13370 (N_13370,N_10040,N_10393);
or U13371 (N_13371,N_10494,N_10534);
nor U13372 (N_13372,N_9971,N_10852);
or U13373 (N_13373,N_10511,N_9903);
nor U13374 (N_13374,N_11875,N_9826);
and U13375 (N_13375,N_10313,N_9582);
nand U13376 (N_13376,N_10304,N_10746);
nand U13377 (N_13377,N_10238,N_9124);
or U13378 (N_13378,N_10386,N_9280);
nand U13379 (N_13379,N_10544,N_10172);
nor U13380 (N_13380,N_10024,N_9664);
or U13381 (N_13381,N_11385,N_11240);
nor U13382 (N_13382,N_11606,N_9357);
or U13383 (N_13383,N_10540,N_10131);
nand U13384 (N_13384,N_11067,N_11965);
or U13385 (N_13385,N_11982,N_9590);
nor U13386 (N_13386,N_9647,N_9198);
nor U13387 (N_13387,N_11201,N_11798);
or U13388 (N_13388,N_11940,N_11891);
and U13389 (N_13389,N_10645,N_11396);
or U13390 (N_13390,N_10163,N_10236);
and U13391 (N_13391,N_11763,N_10274);
or U13392 (N_13392,N_9178,N_11180);
or U13393 (N_13393,N_10145,N_11861);
or U13394 (N_13394,N_9717,N_9882);
nand U13395 (N_13395,N_10216,N_10214);
nor U13396 (N_13396,N_9649,N_11994);
and U13397 (N_13397,N_10739,N_10580);
or U13398 (N_13398,N_9530,N_10193);
nor U13399 (N_13399,N_9762,N_11514);
and U13400 (N_13400,N_11040,N_10078);
and U13401 (N_13401,N_10017,N_10525);
nand U13402 (N_13402,N_11772,N_10790);
nor U13403 (N_13403,N_11675,N_10696);
or U13404 (N_13404,N_10882,N_11031);
or U13405 (N_13405,N_10287,N_9867);
or U13406 (N_13406,N_11900,N_9676);
or U13407 (N_13407,N_9402,N_9842);
or U13408 (N_13408,N_10401,N_10678);
or U13409 (N_13409,N_10139,N_9993);
or U13410 (N_13410,N_10361,N_11759);
nor U13411 (N_13411,N_9289,N_10771);
or U13412 (N_13412,N_10662,N_11666);
nor U13413 (N_13413,N_11410,N_9243);
or U13414 (N_13414,N_10910,N_10849);
nand U13415 (N_13415,N_10730,N_9179);
or U13416 (N_13416,N_9576,N_9829);
or U13417 (N_13417,N_9295,N_11971);
nor U13418 (N_13418,N_10044,N_11052);
and U13419 (N_13419,N_10526,N_9056);
xor U13420 (N_13420,N_9019,N_11003);
nor U13421 (N_13421,N_10477,N_10420);
nand U13422 (N_13422,N_9848,N_9974);
and U13423 (N_13423,N_10571,N_9477);
nand U13424 (N_13424,N_10470,N_11053);
nor U13425 (N_13425,N_9493,N_11405);
or U13426 (N_13426,N_10010,N_9765);
nor U13427 (N_13427,N_10747,N_9713);
and U13428 (N_13428,N_11705,N_10377);
nor U13429 (N_13429,N_10222,N_11929);
or U13430 (N_13430,N_10641,N_10607);
nand U13431 (N_13431,N_11850,N_9663);
and U13432 (N_13432,N_10648,N_10613);
and U13433 (N_13433,N_11181,N_11419);
or U13434 (N_13434,N_11101,N_10850);
xnor U13435 (N_13435,N_9927,N_11631);
or U13436 (N_13436,N_9631,N_10657);
or U13437 (N_13437,N_10667,N_9634);
and U13438 (N_13438,N_9244,N_10914);
nand U13439 (N_13439,N_10081,N_9529);
and U13440 (N_13440,N_11400,N_11726);
nand U13441 (N_13441,N_9686,N_9095);
nor U13442 (N_13442,N_11768,N_9763);
nor U13443 (N_13443,N_10713,N_10728);
or U13444 (N_13444,N_11202,N_11334);
nand U13445 (N_13445,N_9063,N_11232);
or U13446 (N_13446,N_10752,N_9865);
or U13447 (N_13447,N_11070,N_10346);
nand U13448 (N_13448,N_10212,N_11379);
nand U13449 (N_13449,N_11853,N_11963);
nand U13450 (N_13450,N_9275,N_10563);
nor U13451 (N_13451,N_10497,N_9835);
nor U13452 (N_13452,N_9359,N_10251);
nor U13453 (N_13453,N_9646,N_9121);
or U13454 (N_13454,N_11244,N_11227);
or U13455 (N_13455,N_10520,N_11570);
and U13456 (N_13456,N_9627,N_10639);
xor U13457 (N_13457,N_9399,N_10853);
nand U13458 (N_13458,N_9963,N_10059);
nand U13459 (N_13459,N_11827,N_11072);
nor U13460 (N_13460,N_11917,N_9215);
and U13461 (N_13461,N_10695,N_9642);
nor U13462 (N_13462,N_11089,N_11382);
and U13463 (N_13463,N_10686,N_10192);
and U13464 (N_13464,N_10537,N_11255);
nand U13465 (N_13465,N_9731,N_9362);
and U13466 (N_13466,N_10729,N_11129);
nand U13467 (N_13467,N_10784,N_9031);
and U13468 (N_13468,N_11838,N_11044);
nor U13469 (N_13469,N_11591,N_11765);
nand U13470 (N_13470,N_9452,N_10821);
nand U13471 (N_13471,N_11645,N_10671);
or U13472 (N_13472,N_10234,N_11934);
nand U13473 (N_13473,N_11322,N_9834);
nor U13474 (N_13474,N_10528,N_10360);
or U13475 (N_13475,N_9967,N_9287);
nor U13476 (N_13476,N_9580,N_10929);
or U13477 (N_13477,N_11540,N_10189);
nor U13478 (N_13478,N_11617,N_11659);
nor U13479 (N_13479,N_10045,N_9255);
nor U13480 (N_13480,N_11184,N_9078);
and U13481 (N_13481,N_9039,N_9522);
and U13482 (N_13482,N_9587,N_11313);
nand U13483 (N_13483,N_9701,N_9172);
and U13484 (N_13484,N_9262,N_9164);
or U13485 (N_13485,N_9294,N_11557);
nand U13486 (N_13486,N_9216,N_9269);
and U13487 (N_13487,N_9297,N_10698);
nand U13488 (N_13488,N_9128,N_10026);
nand U13489 (N_13489,N_9474,N_11335);
and U13490 (N_13490,N_9711,N_11508);
nand U13491 (N_13491,N_11706,N_10073);
or U13492 (N_13492,N_10467,N_10804);
and U13493 (N_13493,N_9416,N_10249);
and U13494 (N_13494,N_10621,N_9133);
nor U13495 (N_13495,N_9174,N_11460);
or U13496 (N_13496,N_11238,N_10938);
nand U13497 (N_13497,N_10958,N_9823);
xnor U13498 (N_13498,N_9675,N_10202);
and U13499 (N_13499,N_9962,N_9639);
nor U13500 (N_13500,N_11279,N_11850);
and U13501 (N_13501,N_11582,N_11315);
and U13502 (N_13502,N_10492,N_10207);
nand U13503 (N_13503,N_11427,N_11918);
nor U13504 (N_13504,N_11751,N_9304);
nand U13505 (N_13505,N_10414,N_10193);
nor U13506 (N_13506,N_9071,N_9271);
and U13507 (N_13507,N_11500,N_11820);
nor U13508 (N_13508,N_9157,N_11199);
nor U13509 (N_13509,N_9772,N_10613);
and U13510 (N_13510,N_9785,N_10437);
and U13511 (N_13511,N_10826,N_9474);
and U13512 (N_13512,N_9259,N_9771);
or U13513 (N_13513,N_9806,N_11641);
or U13514 (N_13514,N_9897,N_10153);
or U13515 (N_13515,N_10993,N_9818);
and U13516 (N_13516,N_11457,N_10073);
or U13517 (N_13517,N_10206,N_11785);
nand U13518 (N_13518,N_10789,N_10092);
and U13519 (N_13519,N_9875,N_10645);
nor U13520 (N_13520,N_11903,N_11220);
or U13521 (N_13521,N_9295,N_11170);
or U13522 (N_13522,N_11876,N_9028);
nor U13523 (N_13523,N_11952,N_10199);
nand U13524 (N_13524,N_11737,N_11844);
nand U13525 (N_13525,N_10422,N_10818);
nand U13526 (N_13526,N_10184,N_10505);
nand U13527 (N_13527,N_9759,N_9733);
nand U13528 (N_13528,N_9079,N_9351);
nor U13529 (N_13529,N_9257,N_10989);
nor U13530 (N_13530,N_9415,N_11987);
nand U13531 (N_13531,N_10016,N_9534);
nand U13532 (N_13532,N_11733,N_10711);
and U13533 (N_13533,N_11163,N_10621);
nor U13534 (N_13534,N_10000,N_11444);
nand U13535 (N_13535,N_11093,N_9227);
nand U13536 (N_13536,N_9136,N_10973);
nor U13537 (N_13537,N_11325,N_10266);
or U13538 (N_13538,N_9445,N_10305);
and U13539 (N_13539,N_9257,N_10707);
nand U13540 (N_13540,N_11422,N_10360);
nand U13541 (N_13541,N_10046,N_11005);
nand U13542 (N_13542,N_11037,N_9638);
or U13543 (N_13543,N_10410,N_11419);
and U13544 (N_13544,N_11637,N_9659);
and U13545 (N_13545,N_10696,N_11284);
nor U13546 (N_13546,N_9204,N_11947);
nor U13547 (N_13547,N_9983,N_9371);
nor U13548 (N_13548,N_9680,N_9767);
nand U13549 (N_13549,N_9374,N_10474);
nand U13550 (N_13550,N_11145,N_10614);
nand U13551 (N_13551,N_9988,N_11472);
or U13552 (N_13552,N_10884,N_9411);
nor U13553 (N_13553,N_11297,N_9183);
nor U13554 (N_13554,N_9989,N_9674);
nand U13555 (N_13555,N_10066,N_10036);
nand U13556 (N_13556,N_9074,N_11681);
xnor U13557 (N_13557,N_11742,N_9393);
and U13558 (N_13558,N_10875,N_10331);
and U13559 (N_13559,N_11771,N_10786);
and U13560 (N_13560,N_10208,N_11098);
nand U13561 (N_13561,N_9439,N_10494);
nand U13562 (N_13562,N_11685,N_9777);
and U13563 (N_13563,N_11754,N_10157);
and U13564 (N_13564,N_10802,N_10523);
and U13565 (N_13565,N_9517,N_9102);
or U13566 (N_13566,N_9025,N_9809);
nand U13567 (N_13567,N_9697,N_10723);
or U13568 (N_13568,N_10380,N_10663);
nor U13569 (N_13569,N_10906,N_11488);
or U13570 (N_13570,N_9096,N_9037);
or U13571 (N_13571,N_11050,N_11564);
nand U13572 (N_13572,N_11927,N_11299);
nand U13573 (N_13573,N_11388,N_11046);
nand U13574 (N_13574,N_9605,N_11756);
xor U13575 (N_13575,N_9354,N_11971);
nand U13576 (N_13576,N_10952,N_11451);
and U13577 (N_13577,N_9073,N_10402);
and U13578 (N_13578,N_9554,N_10571);
or U13579 (N_13579,N_11327,N_10052);
nor U13580 (N_13580,N_11426,N_11849);
and U13581 (N_13581,N_9462,N_10486);
and U13582 (N_13582,N_10756,N_9511);
and U13583 (N_13583,N_10788,N_10826);
or U13584 (N_13584,N_11450,N_9054);
or U13585 (N_13585,N_11739,N_11333);
and U13586 (N_13586,N_10717,N_10240);
or U13587 (N_13587,N_9533,N_10111);
xnor U13588 (N_13588,N_10523,N_10121);
nand U13589 (N_13589,N_9423,N_9848);
or U13590 (N_13590,N_10134,N_10648);
or U13591 (N_13591,N_11316,N_11020);
or U13592 (N_13592,N_11886,N_10134);
nand U13593 (N_13593,N_10550,N_10959);
nor U13594 (N_13594,N_11217,N_9524);
nand U13595 (N_13595,N_9715,N_11858);
nand U13596 (N_13596,N_11036,N_9278);
and U13597 (N_13597,N_9421,N_9232);
nand U13598 (N_13598,N_11623,N_9768);
nand U13599 (N_13599,N_11580,N_9248);
and U13600 (N_13600,N_10794,N_10005);
and U13601 (N_13601,N_9685,N_9995);
xnor U13602 (N_13602,N_9038,N_10423);
and U13603 (N_13603,N_11252,N_11195);
or U13604 (N_13604,N_10306,N_11978);
nand U13605 (N_13605,N_11032,N_9493);
or U13606 (N_13606,N_11643,N_9889);
nand U13607 (N_13607,N_9408,N_11467);
or U13608 (N_13608,N_10268,N_11512);
nor U13609 (N_13609,N_9307,N_10163);
nor U13610 (N_13610,N_10843,N_11994);
and U13611 (N_13611,N_11907,N_9473);
or U13612 (N_13612,N_11251,N_11412);
xnor U13613 (N_13613,N_9314,N_11425);
and U13614 (N_13614,N_11695,N_10863);
nor U13615 (N_13615,N_11825,N_10081);
nand U13616 (N_13616,N_11269,N_9312);
or U13617 (N_13617,N_10574,N_9226);
nand U13618 (N_13618,N_9793,N_10279);
nor U13619 (N_13619,N_9719,N_11823);
nor U13620 (N_13620,N_9396,N_9800);
and U13621 (N_13621,N_10172,N_10845);
or U13622 (N_13622,N_10094,N_10555);
nor U13623 (N_13623,N_9613,N_11426);
nor U13624 (N_13624,N_10818,N_10329);
nor U13625 (N_13625,N_11897,N_10305);
nor U13626 (N_13626,N_11489,N_10525);
and U13627 (N_13627,N_11872,N_9863);
or U13628 (N_13628,N_11180,N_9258);
nand U13629 (N_13629,N_10837,N_11676);
nand U13630 (N_13630,N_10930,N_10097);
nor U13631 (N_13631,N_10845,N_9971);
nand U13632 (N_13632,N_10037,N_10865);
and U13633 (N_13633,N_11874,N_10928);
or U13634 (N_13634,N_9275,N_9051);
xor U13635 (N_13635,N_11149,N_10893);
or U13636 (N_13636,N_11309,N_10841);
nand U13637 (N_13637,N_11172,N_10024);
nor U13638 (N_13638,N_10777,N_10154);
nand U13639 (N_13639,N_9633,N_9775);
or U13640 (N_13640,N_10335,N_10939);
and U13641 (N_13641,N_9859,N_9563);
nand U13642 (N_13642,N_9045,N_10635);
nor U13643 (N_13643,N_9224,N_9659);
and U13644 (N_13644,N_9619,N_11157);
nand U13645 (N_13645,N_10069,N_9884);
nand U13646 (N_13646,N_10563,N_9303);
nor U13647 (N_13647,N_11960,N_9198);
and U13648 (N_13648,N_10864,N_10982);
and U13649 (N_13649,N_9175,N_10697);
or U13650 (N_13650,N_11731,N_11850);
or U13651 (N_13651,N_10203,N_11784);
nand U13652 (N_13652,N_9174,N_10475);
and U13653 (N_13653,N_10722,N_10739);
and U13654 (N_13654,N_11644,N_10881);
or U13655 (N_13655,N_9685,N_11287);
and U13656 (N_13656,N_11714,N_9610);
and U13657 (N_13657,N_10866,N_9746);
and U13658 (N_13658,N_11072,N_11338);
and U13659 (N_13659,N_10324,N_11392);
nand U13660 (N_13660,N_9662,N_11431);
nand U13661 (N_13661,N_9258,N_11253);
nor U13662 (N_13662,N_11282,N_11481);
or U13663 (N_13663,N_11414,N_9801);
or U13664 (N_13664,N_9552,N_9388);
and U13665 (N_13665,N_11328,N_9145);
and U13666 (N_13666,N_9748,N_9897);
nand U13667 (N_13667,N_10604,N_10600);
or U13668 (N_13668,N_11872,N_9521);
and U13669 (N_13669,N_10027,N_11980);
nor U13670 (N_13670,N_11406,N_9587);
nand U13671 (N_13671,N_11801,N_9077);
nor U13672 (N_13672,N_10176,N_9896);
or U13673 (N_13673,N_10843,N_9736);
or U13674 (N_13674,N_11386,N_9984);
nand U13675 (N_13675,N_9230,N_10283);
nand U13676 (N_13676,N_9702,N_9378);
nand U13677 (N_13677,N_11647,N_9336);
or U13678 (N_13678,N_10681,N_9895);
or U13679 (N_13679,N_11559,N_10355);
nand U13680 (N_13680,N_9418,N_9756);
or U13681 (N_13681,N_9757,N_11577);
nand U13682 (N_13682,N_9007,N_9404);
nor U13683 (N_13683,N_10907,N_9215);
nand U13684 (N_13684,N_10949,N_9909);
and U13685 (N_13685,N_9354,N_11322);
and U13686 (N_13686,N_11860,N_9879);
or U13687 (N_13687,N_9363,N_11023);
or U13688 (N_13688,N_11557,N_9664);
nor U13689 (N_13689,N_9737,N_11825);
and U13690 (N_13690,N_11885,N_9251);
nand U13691 (N_13691,N_9941,N_10698);
nand U13692 (N_13692,N_10643,N_11726);
or U13693 (N_13693,N_10820,N_9150);
or U13694 (N_13694,N_10478,N_11549);
nor U13695 (N_13695,N_9869,N_9542);
nand U13696 (N_13696,N_9644,N_10978);
or U13697 (N_13697,N_10266,N_10376);
nor U13698 (N_13698,N_9733,N_11790);
or U13699 (N_13699,N_11566,N_9577);
and U13700 (N_13700,N_9668,N_10744);
and U13701 (N_13701,N_10609,N_11004);
nor U13702 (N_13702,N_10410,N_10067);
nand U13703 (N_13703,N_11650,N_9368);
or U13704 (N_13704,N_9999,N_9579);
nand U13705 (N_13705,N_11378,N_10066);
nand U13706 (N_13706,N_11717,N_11966);
nor U13707 (N_13707,N_11522,N_11553);
nor U13708 (N_13708,N_9660,N_10338);
or U13709 (N_13709,N_9702,N_10285);
nand U13710 (N_13710,N_10459,N_10189);
and U13711 (N_13711,N_11764,N_11502);
nor U13712 (N_13712,N_9561,N_10756);
and U13713 (N_13713,N_11575,N_9822);
and U13714 (N_13714,N_10982,N_9929);
nor U13715 (N_13715,N_9814,N_11429);
or U13716 (N_13716,N_10676,N_10701);
nand U13717 (N_13717,N_11021,N_11416);
nand U13718 (N_13718,N_10206,N_10001);
or U13719 (N_13719,N_10525,N_10946);
and U13720 (N_13720,N_10026,N_9349);
nand U13721 (N_13721,N_11405,N_9003);
nand U13722 (N_13722,N_10708,N_10752);
nor U13723 (N_13723,N_11429,N_11009);
or U13724 (N_13724,N_10199,N_9306);
nand U13725 (N_13725,N_10924,N_10705);
nand U13726 (N_13726,N_9151,N_11150);
and U13727 (N_13727,N_9439,N_9407);
and U13728 (N_13728,N_9882,N_10897);
or U13729 (N_13729,N_11360,N_11235);
and U13730 (N_13730,N_11032,N_11894);
nand U13731 (N_13731,N_11870,N_9803);
nor U13732 (N_13732,N_11488,N_10076);
nor U13733 (N_13733,N_9169,N_9193);
and U13734 (N_13734,N_9803,N_9891);
nor U13735 (N_13735,N_11273,N_10314);
nor U13736 (N_13736,N_10840,N_11886);
or U13737 (N_13737,N_11674,N_11345);
and U13738 (N_13738,N_11642,N_11780);
and U13739 (N_13739,N_11409,N_10616);
nand U13740 (N_13740,N_11439,N_10479);
or U13741 (N_13741,N_11317,N_10307);
and U13742 (N_13742,N_10955,N_11023);
and U13743 (N_13743,N_11095,N_9588);
nand U13744 (N_13744,N_11474,N_10409);
and U13745 (N_13745,N_9216,N_9767);
or U13746 (N_13746,N_10007,N_10593);
or U13747 (N_13747,N_9745,N_9491);
and U13748 (N_13748,N_11882,N_9503);
nor U13749 (N_13749,N_10116,N_9768);
or U13750 (N_13750,N_9273,N_10665);
nand U13751 (N_13751,N_9855,N_11533);
nand U13752 (N_13752,N_9492,N_10134);
nand U13753 (N_13753,N_9431,N_10553);
or U13754 (N_13754,N_11509,N_10289);
nand U13755 (N_13755,N_9255,N_9726);
and U13756 (N_13756,N_9372,N_10385);
or U13757 (N_13757,N_11167,N_10154);
nand U13758 (N_13758,N_9434,N_9400);
nand U13759 (N_13759,N_11422,N_10945);
nor U13760 (N_13760,N_9571,N_11206);
nor U13761 (N_13761,N_10254,N_9376);
and U13762 (N_13762,N_10368,N_10223);
or U13763 (N_13763,N_9066,N_11328);
nor U13764 (N_13764,N_11346,N_10159);
and U13765 (N_13765,N_9445,N_9508);
nor U13766 (N_13766,N_11826,N_11033);
nand U13767 (N_13767,N_9019,N_9496);
or U13768 (N_13768,N_11453,N_10749);
nand U13769 (N_13769,N_10980,N_10583);
and U13770 (N_13770,N_10267,N_9301);
xor U13771 (N_13771,N_9189,N_9866);
or U13772 (N_13772,N_9949,N_9121);
nor U13773 (N_13773,N_11423,N_9336);
nand U13774 (N_13774,N_9591,N_9212);
or U13775 (N_13775,N_9466,N_9352);
nor U13776 (N_13776,N_10769,N_9624);
or U13777 (N_13777,N_9730,N_10541);
nor U13778 (N_13778,N_10251,N_11335);
or U13779 (N_13779,N_11879,N_9826);
nor U13780 (N_13780,N_11161,N_9867);
and U13781 (N_13781,N_9788,N_10473);
nand U13782 (N_13782,N_11754,N_10959);
nand U13783 (N_13783,N_11186,N_11935);
and U13784 (N_13784,N_9455,N_9055);
and U13785 (N_13785,N_9485,N_10900);
or U13786 (N_13786,N_9346,N_10658);
and U13787 (N_13787,N_11546,N_10655);
or U13788 (N_13788,N_9595,N_9963);
nor U13789 (N_13789,N_9730,N_9873);
nor U13790 (N_13790,N_10419,N_9289);
nor U13791 (N_13791,N_11243,N_10112);
nand U13792 (N_13792,N_10549,N_11237);
or U13793 (N_13793,N_11044,N_11238);
nand U13794 (N_13794,N_11122,N_11184);
and U13795 (N_13795,N_10631,N_10174);
or U13796 (N_13796,N_10954,N_9398);
nor U13797 (N_13797,N_9871,N_11963);
and U13798 (N_13798,N_10534,N_11376);
nor U13799 (N_13799,N_9818,N_9036);
and U13800 (N_13800,N_11069,N_9798);
nand U13801 (N_13801,N_9456,N_10868);
nor U13802 (N_13802,N_11900,N_10436);
nor U13803 (N_13803,N_11468,N_9335);
nand U13804 (N_13804,N_11603,N_10389);
nor U13805 (N_13805,N_10769,N_10574);
nor U13806 (N_13806,N_10125,N_9176);
and U13807 (N_13807,N_10532,N_9609);
and U13808 (N_13808,N_10693,N_10535);
or U13809 (N_13809,N_10969,N_9553);
and U13810 (N_13810,N_10172,N_11952);
nor U13811 (N_13811,N_11096,N_11136);
nor U13812 (N_13812,N_9467,N_10795);
and U13813 (N_13813,N_9823,N_9397);
nand U13814 (N_13814,N_10867,N_10795);
nand U13815 (N_13815,N_10733,N_10961);
and U13816 (N_13816,N_11861,N_11630);
xor U13817 (N_13817,N_11679,N_10348);
nand U13818 (N_13818,N_10409,N_10252);
or U13819 (N_13819,N_9968,N_9996);
nor U13820 (N_13820,N_10952,N_9129);
nand U13821 (N_13821,N_11308,N_10368);
nand U13822 (N_13822,N_10821,N_10472);
nand U13823 (N_13823,N_11745,N_10864);
nand U13824 (N_13824,N_10528,N_10463);
nor U13825 (N_13825,N_11013,N_10064);
and U13826 (N_13826,N_9335,N_10711);
or U13827 (N_13827,N_9404,N_10905);
or U13828 (N_13828,N_10003,N_10297);
nand U13829 (N_13829,N_10590,N_11642);
and U13830 (N_13830,N_11875,N_11051);
nand U13831 (N_13831,N_10858,N_9410);
nor U13832 (N_13832,N_11694,N_10328);
nor U13833 (N_13833,N_10303,N_11528);
and U13834 (N_13834,N_11555,N_11108);
nand U13835 (N_13835,N_9715,N_10678);
nand U13836 (N_13836,N_9231,N_11704);
or U13837 (N_13837,N_11508,N_10019);
or U13838 (N_13838,N_10494,N_10747);
and U13839 (N_13839,N_10534,N_10943);
nand U13840 (N_13840,N_10578,N_10490);
and U13841 (N_13841,N_10668,N_11262);
and U13842 (N_13842,N_9568,N_11382);
or U13843 (N_13843,N_9506,N_9116);
nand U13844 (N_13844,N_9919,N_10628);
nand U13845 (N_13845,N_10107,N_11471);
nand U13846 (N_13846,N_10833,N_10496);
nand U13847 (N_13847,N_10119,N_9394);
or U13848 (N_13848,N_10947,N_10870);
nor U13849 (N_13849,N_10774,N_10570);
nand U13850 (N_13850,N_11355,N_10485);
and U13851 (N_13851,N_9994,N_10402);
and U13852 (N_13852,N_11920,N_9295);
nand U13853 (N_13853,N_9868,N_10893);
nor U13854 (N_13854,N_11175,N_9350);
or U13855 (N_13855,N_10339,N_9055);
and U13856 (N_13856,N_9011,N_9359);
nor U13857 (N_13857,N_9756,N_10317);
or U13858 (N_13858,N_11688,N_11722);
nor U13859 (N_13859,N_10237,N_11236);
or U13860 (N_13860,N_9676,N_11364);
nor U13861 (N_13861,N_9327,N_9662);
or U13862 (N_13862,N_10901,N_11698);
and U13863 (N_13863,N_11941,N_11498);
nor U13864 (N_13864,N_11870,N_11695);
nor U13865 (N_13865,N_9275,N_9553);
nor U13866 (N_13866,N_11205,N_9053);
and U13867 (N_13867,N_10860,N_10475);
nand U13868 (N_13868,N_10913,N_9529);
and U13869 (N_13869,N_11509,N_9174);
and U13870 (N_13870,N_9444,N_11512);
or U13871 (N_13871,N_9602,N_11965);
nand U13872 (N_13872,N_9480,N_11520);
and U13873 (N_13873,N_11260,N_9897);
or U13874 (N_13874,N_10609,N_9667);
xor U13875 (N_13875,N_10891,N_9253);
and U13876 (N_13876,N_10047,N_10004);
or U13877 (N_13877,N_11543,N_10932);
and U13878 (N_13878,N_9891,N_9869);
nor U13879 (N_13879,N_9522,N_10390);
and U13880 (N_13880,N_11713,N_10484);
and U13881 (N_13881,N_9951,N_9335);
xnor U13882 (N_13882,N_10943,N_9980);
and U13883 (N_13883,N_9030,N_10648);
nand U13884 (N_13884,N_9691,N_11891);
or U13885 (N_13885,N_10676,N_10250);
or U13886 (N_13886,N_9126,N_11740);
nand U13887 (N_13887,N_10208,N_10603);
nand U13888 (N_13888,N_11462,N_9404);
nand U13889 (N_13889,N_9062,N_9948);
nor U13890 (N_13890,N_10470,N_11858);
nand U13891 (N_13891,N_11233,N_10483);
and U13892 (N_13892,N_11696,N_9295);
and U13893 (N_13893,N_9919,N_9465);
nor U13894 (N_13894,N_11481,N_9473);
or U13895 (N_13895,N_11060,N_10212);
xnor U13896 (N_13896,N_10865,N_9730);
nand U13897 (N_13897,N_9766,N_9746);
nor U13898 (N_13898,N_9031,N_11527);
or U13899 (N_13899,N_10235,N_9150);
nand U13900 (N_13900,N_9196,N_9697);
nand U13901 (N_13901,N_10731,N_9965);
nor U13902 (N_13902,N_10228,N_11722);
nand U13903 (N_13903,N_10601,N_10705);
nor U13904 (N_13904,N_10140,N_10342);
nand U13905 (N_13905,N_11621,N_9576);
nor U13906 (N_13906,N_9797,N_9611);
nor U13907 (N_13907,N_11479,N_9036);
and U13908 (N_13908,N_11446,N_11468);
and U13909 (N_13909,N_9772,N_10356);
and U13910 (N_13910,N_11442,N_9447);
and U13911 (N_13911,N_9767,N_9839);
and U13912 (N_13912,N_9836,N_10530);
xnor U13913 (N_13913,N_9485,N_9668);
nor U13914 (N_13914,N_10518,N_10290);
or U13915 (N_13915,N_10019,N_10268);
or U13916 (N_13916,N_9270,N_11026);
and U13917 (N_13917,N_9851,N_9239);
nand U13918 (N_13918,N_9608,N_9636);
and U13919 (N_13919,N_11573,N_10300);
or U13920 (N_13920,N_9793,N_11681);
or U13921 (N_13921,N_11212,N_9781);
nand U13922 (N_13922,N_11837,N_11842);
nor U13923 (N_13923,N_10540,N_9252);
nor U13924 (N_13924,N_10719,N_10439);
nand U13925 (N_13925,N_9979,N_11939);
and U13926 (N_13926,N_11861,N_11975);
and U13927 (N_13927,N_11737,N_10272);
and U13928 (N_13928,N_9363,N_10572);
nand U13929 (N_13929,N_11159,N_11257);
or U13930 (N_13930,N_11641,N_10778);
or U13931 (N_13931,N_10177,N_10999);
and U13932 (N_13932,N_9995,N_11084);
nand U13933 (N_13933,N_9463,N_10321);
nand U13934 (N_13934,N_10783,N_11256);
and U13935 (N_13935,N_9977,N_10149);
and U13936 (N_13936,N_11729,N_11751);
and U13937 (N_13937,N_9810,N_9831);
and U13938 (N_13938,N_9180,N_11918);
nor U13939 (N_13939,N_11160,N_11028);
nor U13940 (N_13940,N_11931,N_11939);
nand U13941 (N_13941,N_11713,N_9186);
nor U13942 (N_13942,N_10984,N_11887);
and U13943 (N_13943,N_11296,N_9507);
nand U13944 (N_13944,N_11057,N_11908);
or U13945 (N_13945,N_10276,N_11264);
nand U13946 (N_13946,N_11517,N_11805);
and U13947 (N_13947,N_10886,N_10317);
xnor U13948 (N_13948,N_9922,N_10885);
and U13949 (N_13949,N_9772,N_9458);
and U13950 (N_13950,N_11529,N_11669);
nor U13951 (N_13951,N_10520,N_11660);
or U13952 (N_13952,N_11818,N_9827);
nand U13953 (N_13953,N_11730,N_9553);
and U13954 (N_13954,N_10514,N_11591);
nor U13955 (N_13955,N_9111,N_9861);
and U13956 (N_13956,N_10540,N_9067);
nor U13957 (N_13957,N_10224,N_10423);
or U13958 (N_13958,N_9442,N_10243);
nand U13959 (N_13959,N_9979,N_10451);
and U13960 (N_13960,N_10762,N_10048);
and U13961 (N_13961,N_10821,N_11611);
nor U13962 (N_13962,N_10300,N_11777);
or U13963 (N_13963,N_9844,N_11142);
nor U13964 (N_13964,N_10127,N_11843);
and U13965 (N_13965,N_11778,N_10311);
or U13966 (N_13966,N_11583,N_9191);
or U13967 (N_13967,N_9160,N_9937);
nor U13968 (N_13968,N_9470,N_9231);
and U13969 (N_13969,N_9935,N_9082);
nand U13970 (N_13970,N_11165,N_11762);
and U13971 (N_13971,N_9475,N_11651);
xnor U13972 (N_13972,N_11334,N_11912);
and U13973 (N_13973,N_10525,N_9012);
nand U13974 (N_13974,N_9263,N_11052);
xor U13975 (N_13975,N_11335,N_11297);
nand U13976 (N_13976,N_11907,N_9139);
nor U13977 (N_13977,N_10538,N_10053);
nor U13978 (N_13978,N_10864,N_11953);
and U13979 (N_13979,N_10536,N_9186);
and U13980 (N_13980,N_11504,N_10116);
nand U13981 (N_13981,N_10654,N_9067);
nand U13982 (N_13982,N_10592,N_9357);
nor U13983 (N_13983,N_9651,N_11935);
or U13984 (N_13984,N_10234,N_9762);
and U13985 (N_13985,N_9923,N_11607);
and U13986 (N_13986,N_10573,N_10074);
nand U13987 (N_13987,N_11492,N_9337);
and U13988 (N_13988,N_10874,N_9316);
and U13989 (N_13989,N_10756,N_11456);
nand U13990 (N_13990,N_10801,N_10594);
or U13991 (N_13991,N_9126,N_11568);
or U13992 (N_13992,N_9274,N_11668);
nor U13993 (N_13993,N_9431,N_9107);
and U13994 (N_13994,N_11357,N_10750);
xor U13995 (N_13995,N_10607,N_9897);
nor U13996 (N_13996,N_9776,N_10232);
nor U13997 (N_13997,N_9610,N_9099);
nand U13998 (N_13998,N_10927,N_9393);
nor U13999 (N_13999,N_11267,N_9282);
nor U14000 (N_14000,N_9369,N_10993);
nand U14001 (N_14001,N_9115,N_10492);
and U14002 (N_14002,N_10966,N_11633);
nor U14003 (N_14003,N_11603,N_11911);
nand U14004 (N_14004,N_9833,N_10966);
nand U14005 (N_14005,N_9656,N_11455);
or U14006 (N_14006,N_10747,N_9567);
nor U14007 (N_14007,N_11033,N_11580);
nand U14008 (N_14008,N_9479,N_9501);
and U14009 (N_14009,N_10913,N_10772);
nor U14010 (N_14010,N_10957,N_11929);
nor U14011 (N_14011,N_9143,N_9318);
and U14012 (N_14012,N_9643,N_11747);
or U14013 (N_14013,N_11472,N_10423);
nor U14014 (N_14014,N_9391,N_11047);
or U14015 (N_14015,N_10630,N_11211);
nor U14016 (N_14016,N_11983,N_9511);
and U14017 (N_14017,N_11038,N_10374);
xnor U14018 (N_14018,N_9012,N_11635);
nor U14019 (N_14019,N_9934,N_9134);
and U14020 (N_14020,N_11855,N_11579);
nor U14021 (N_14021,N_10601,N_9556);
and U14022 (N_14022,N_9554,N_11655);
nor U14023 (N_14023,N_9713,N_11299);
nand U14024 (N_14024,N_9129,N_10645);
and U14025 (N_14025,N_11596,N_9562);
or U14026 (N_14026,N_11164,N_10921);
nor U14027 (N_14027,N_9872,N_10762);
and U14028 (N_14028,N_10895,N_10677);
and U14029 (N_14029,N_10449,N_10527);
or U14030 (N_14030,N_10649,N_10026);
and U14031 (N_14031,N_10880,N_10309);
nand U14032 (N_14032,N_10205,N_9504);
and U14033 (N_14033,N_9770,N_9882);
or U14034 (N_14034,N_10974,N_11084);
xor U14035 (N_14035,N_10682,N_10319);
xor U14036 (N_14036,N_11058,N_9258);
and U14037 (N_14037,N_9290,N_9166);
or U14038 (N_14038,N_11118,N_9393);
nor U14039 (N_14039,N_10556,N_9012);
nor U14040 (N_14040,N_9782,N_11434);
nand U14041 (N_14041,N_9342,N_9713);
or U14042 (N_14042,N_10447,N_10793);
or U14043 (N_14043,N_11740,N_11010);
and U14044 (N_14044,N_11780,N_11892);
and U14045 (N_14045,N_9617,N_11606);
nor U14046 (N_14046,N_10821,N_11866);
nand U14047 (N_14047,N_10443,N_10772);
or U14048 (N_14048,N_9065,N_9643);
or U14049 (N_14049,N_10817,N_11389);
and U14050 (N_14050,N_10997,N_10754);
nor U14051 (N_14051,N_9502,N_9179);
nor U14052 (N_14052,N_11908,N_10334);
nor U14053 (N_14053,N_11168,N_10760);
nor U14054 (N_14054,N_11067,N_11095);
or U14055 (N_14055,N_11015,N_10599);
or U14056 (N_14056,N_11026,N_11093);
nor U14057 (N_14057,N_10497,N_10689);
and U14058 (N_14058,N_11689,N_10788);
xor U14059 (N_14059,N_9418,N_11408);
nand U14060 (N_14060,N_9069,N_9964);
or U14061 (N_14061,N_11657,N_11858);
nor U14062 (N_14062,N_11673,N_9850);
nor U14063 (N_14063,N_11400,N_10132);
and U14064 (N_14064,N_9419,N_10278);
and U14065 (N_14065,N_11852,N_9909);
or U14066 (N_14066,N_10374,N_11963);
xnor U14067 (N_14067,N_10037,N_10661);
nor U14068 (N_14068,N_10041,N_9807);
and U14069 (N_14069,N_10135,N_9699);
or U14070 (N_14070,N_9266,N_9303);
or U14071 (N_14071,N_9204,N_11154);
nor U14072 (N_14072,N_11120,N_10330);
nand U14073 (N_14073,N_10697,N_10982);
or U14074 (N_14074,N_11319,N_11085);
nor U14075 (N_14075,N_9618,N_10717);
and U14076 (N_14076,N_10297,N_10410);
or U14077 (N_14077,N_9662,N_11177);
and U14078 (N_14078,N_11111,N_9623);
or U14079 (N_14079,N_11363,N_9812);
nor U14080 (N_14080,N_9087,N_9685);
and U14081 (N_14081,N_10028,N_10492);
or U14082 (N_14082,N_10496,N_11121);
and U14083 (N_14083,N_10878,N_9780);
nand U14084 (N_14084,N_9816,N_11781);
nor U14085 (N_14085,N_10233,N_10893);
or U14086 (N_14086,N_9192,N_11457);
and U14087 (N_14087,N_11459,N_10904);
or U14088 (N_14088,N_10233,N_10215);
and U14089 (N_14089,N_10774,N_10549);
or U14090 (N_14090,N_9940,N_9075);
nor U14091 (N_14091,N_9027,N_10994);
or U14092 (N_14092,N_9089,N_11272);
or U14093 (N_14093,N_11654,N_9166);
and U14094 (N_14094,N_11305,N_11848);
or U14095 (N_14095,N_10180,N_9660);
nor U14096 (N_14096,N_11947,N_10858);
xnor U14097 (N_14097,N_10755,N_10753);
nor U14098 (N_14098,N_9404,N_10148);
or U14099 (N_14099,N_11139,N_11865);
xor U14100 (N_14100,N_9556,N_9418);
xnor U14101 (N_14101,N_11624,N_9714);
nor U14102 (N_14102,N_10259,N_10773);
or U14103 (N_14103,N_9897,N_11748);
nand U14104 (N_14104,N_10836,N_11480);
or U14105 (N_14105,N_11359,N_10625);
and U14106 (N_14106,N_9162,N_11021);
and U14107 (N_14107,N_11652,N_11596);
nand U14108 (N_14108,N_10791,N_10510);
nand U14109 (N_14109,N_10261,N_11418);
or U14110 (N_14110,N_9334,N_10077);
and U14111 (N_14111,N_10744,N_9617);
or U14112 (N_14112,N_10621,N_9283);
and U14113 (N_14113,N_10782,N_9987);
nor U14114 (N_14114,N_9083,N_10948);
and U14115 (N_14115,N_9617,N_11889);
or U14116 (N_14116,N_11461,N_10895);
and U14117 (N_14117,N_11640,N_9049);
nor U14118 (N_14118,N_9173,N_10022);
or U14119 (N_14119,N_11126,N_10017);
nor U14120 (N_14120,N_10980,N_11763);
or U14121 (N_14121,N_10211,N_9791);
nor U14122 (N_14122,N_10555,N_11578);
and U14123 (N_14123,N_9598,N_10291);
nor U14124 (N_14124,N_11826,N_10633);
nand U14125 (N_14125,N_9345,N_9168);
nor U14126 (N_14126,N_11178,N_9501);
and U14127 (N_14127,N_10699,N_9974);
xor U14128 (N_14128,N_9671,N_9825);
and U14129 (N_14129,N_9384,N_10708);
and U14130 (N_14130,N_9230,N_9980);
nor U14131 (N_14131,N_9222,N_11765);
nor U14132 (N_14132,N_9432,N_11770);
and U14133 (N_14133,N_11844,N_10318);
or U14134 (N_14134,N_10461,N_9958);
nand U14135 (N_14135,N_10445,N_11183);
or U14136 (N_14136,N_9460,N_10492);
and U14137 (N_14137,N_9328,N_9460);
or U14138 (N_14138,N_10509,N_11572);
nor U14139 (N_14139,N_10707,N_10120);
nor U14140 (N_14140,N_11952,N_10446);
nor U14141 (N_14141,N_11041,N_9752);
nand U14142 (N_14142,N_9364,N_9284);
nand U14143 (N_14143,N_10919,N_10135);
nor U14144 (N_14144,N_9939,N_9978);
or U14145 (N_14145,N_10086,N_9225);
nor U14146 (N_14146,N_11704,N_10829);
nand U14147 (N_14147,N_10294,N_9594);
and U14148 (N_14148,N_11830,N_11463);
xor U14149 (N_14149,N_10689,N_10669);
nor U14150 (N_14150,N_10284,N_11293);
or U14151 (N_14151,N_10325,N_9433);
and U14152 (N_14152,N_11588,N_9566);
and U14153 (N_14153,N_10298,N_9659);
nand U14154 (N_14154,N_11425,N_10815);
nand U14155 (N_14155,N_10313,N_11389);
and U14156 (N_14156,N_11023,N_9423);
nand U14157 (N_14157,N_10949,N_10408);
or U14158 (N_14158,N_9610,N_9783);
nor U14159 (N_14159,N_9937,N_9216);
or U14160 (N_14160,N_11915,N_11805);
or U14161 (N_14161,N_9762,N_9032);
or U14162 (N_14162,N_10331,N_11729);
and U14163 (N_14163,N_10317,N_11065);
nor U14164 (N_14164,N_10757,N_10324);
nor U14165 (N_14165,N_9658,N_10237);
nor U14166 (N_14166,N_11328,N_11391);
nand U14167 (N_14167,N_9629,N_10047);
and U14168 (N_14168,N_11801,N_10684);
and U14169 (N_14169,N_11864,N_9989);
nor U14170 (N_14170,N_10417,N_11636);
nor U14171 (N_14171,N_11299,N_9997);
nand U14172 (N_14172,N_9236,N_11245);
and U14173 (N_14173,N_10559,N_10976);
nor U14174 (N_14174,N_11660,N_11224);
nand U14175 (N_14175,N_10296,N_9376);
nor U14176 (N_14176,N_9274,N_9284);
or U14177 (N_14177,N_11094,N_11225);
nand U14178 (N_14178,N_10690,N_11673);
nand U14179 (N_14179,N_11142,N_9222);
nor U14180 (N_14180,N_10657,N_9568);
and U14181 (N_14181,N_9723,N_11581);
nand U14182 (N_14182,N_11128,N_11809);
nor U14183 (N_14183,N_10054,N_11919);
and U14184 (N_14184,N_10051,N_10546);
nand U14185 (N_14185,N_11674,N_9471);
nor U14186 (N_14186,N_9488,N_9664);
nor U14187 (N_14187,N_11730,N_11398);
or U14188 (N_14188,N_9677,N_11373);
nand U14189 (N_14189,N_11839,N_9387);
nor U14190 (N_14190,N_9142,N_10412);
nor U14191 (N_14191,N_11914,N_10425);
nor U14192 (N_14192,N_10344,N_11879);
nor U14193 (N_14193,N_11949,N_10467);
nor U14194 (N_14194,N_10300,N_9178);
or U14195 (N_14195,N_9899,N_11363);
and U14196 (N_14196,N_10209,N_9702);
or U14197 (N_14197,N_10551,N_10586);
nor U14198 (N_14198,N_11719,N_11288);
and U14199 (N_14199,N_9271,N_11432);
or U14200 (N_14200,N_9369,N_11873);
nor U14201 (N_14201,N_9586,N_11310);
and U14202 (N_14202,N_9700,N_11241);
nand U14203 (N_14203,N_10459,N_11770);
or U14204 (N_14204,N_11164,N_10456);
nor U14205 (N_14205,N_10537,N_9062);
or U14206 (N_14206,N_11053,N_11493);
or U14207 (N_14207,N_9417,N_10154);
nand U14208 (N_14208,N_10063,N_10718);
and U14209 (N_14209,N_9876,N_10336);
or U14210 (N_14210,N_9756,N_9834);
xor U14211 (N_14211,N_11552,N_10551);
xnor U14212 (N_14212,N_10440,N_10236);
nor U14213 (N_14213,N_10101,N_9965);
xnor U14214 (N_14214,N_9820,N_9574);
and U14215 (N_14215,N_10124,N_10826);
and U14216 (N_14216,N_10410,N_10966);
or U14217 (N_14217,N_9946,N_10041);
and U14218 (N_14218,N_9363,N_11383);
nand U14219 (N_14219,N_10726,N_10989);
nor U14220 (N_14220,N_10613,N_9840);
or U14221 (N_14221,N_9371,N_11478);
and U14222 (N_14222,N_11548,N_10391);
and U14223 (N_14223,N_10682,N_9110);
or U14224 (N_14224,N_9626,N_11679);
and U14225 (N_14225,N_9836,N_11380);
or U14226 (N_14226,N_11579,N_9353);
and U14227 (N_14227,N_11437,N_9252);
nand U14228 (N_14228,N_10982,N_10548);
or U14229 (N_14229,N_9233,N_10466);
nor U14230 (N_14230,N_9227,N_9054);
or U14231 (N_14231,N_10741,N_10730);
or U14232 (N_14232,N_9013,N_10837);
nor U14233 (N_14233,N_9208,N_10544);
or U14234 (N_14234,N_9512,N_10297);
and U14235 (N_14235,N_10005,N_9717);
and U14236 (N_14236,N_9099,N_9096);
or U14237 (N_14237,N_10659,N_9956);
and U14238 (N_14238,N_11103,N_9662);
or U14239 (N_14239,N_10183,N_11066);
nor U14240 (N_14240,N_9440,N_10775);
and U14241 (N_14241,N_9046,N_11907);
and U14242 (N_14242,N_9800,N_9593);
nor U14243 (N_14243,N_11363,N_11971);
and U14244 (N_14244,N_9442,N_9505);
nand U14245 (N_14245,N_11293,N_11248);
nand U14246 (N_14246,N_10448,N_11014);
nand U14247 (N_14247,N_10955,N_9523);
or U14248 (N_14248,N_9581,N_10920);
nor U14249 (N_14249,N_9957,N_10906);
and U14250 (N_14250,N_11262,N_10725);
and U14251 (N_14251,N_11026,N_9512);
and U14252 (N_14252,N_9653,N_9323);
xor U14253 (N_14253,N_10539,N_9433);
nor U14254 (N_14254,N_10687,N_9475);
and U14255 (N_14255,N_10326,N_9502);
or U14256 (N_14256,N_10628,N_10225);
and U14257 (N_14257,N_11455,N_10138);
nor U14258 (N_14258,N_9055,N_10739);
nand U14259 (N_14259,N_10527,N_10201);
nor U14260 (N_14260,N_11419,N_11349);
nor U14261 (N_14261,N_9700,N_10516);
nor U14262 (N_14262,N_11211,N_11270);
or U14263 (N_14263,N_9421,N_10883);
nor U14264 (N_14264,N_9178,N_9981);
and U14265 (N_14265,N_10299,N_11743);
or U14266 (N_14266,N_10073,N_11944);
and U14267 (N_14267,N_11049,N_9679);
or U14268 (N_14268,N_10165,N_11468);
nor U14269 (N_14269,N_11666,N_10528);
nand U14270 (N_14270,N_11472,N_10653);
nand U14271 (N_14271,N_9160,N_10040);
and U14272 (N_14272,N_10175,N_9788);
nor U14273 (N_14273,N_10121,N_10020);
and U14274 (N_14274,N_9955,N_11451);
nand U14275 (N_14275,N_11380,N_11086);
nor U14276 (N_14276,N_11910,N_11960);
and U14277 (N_14277,N_9447,N_10282);
or U14278 (N_14278,N_9621,N_9277);
or U14279 (N_14279,N_11846,N_10373);
or U14280 (N_14280,N_9584,N_10846);
nand U14281 (N_14281,N_9218,N_10926);
nand U14282 (N_14282,N_10121,N_11818);
nor U14283 (N_14283,N_11402,N_9171);
and U14284 (N_14284,N_9421,N_9799);
nor U14285 (N_14285,N_10231,N_9904);
nand U14286 (N_14286,N_11564,N_10743);
or U14287 (N_14287,N_11430,N_10823);
nor U14288 (N_14288,N_11886,N_9557);
or U14289 (N_14289,N_11654,N_11633);
nor U14290 (N_14290,N_10412,N_10927);
or U14291 (N_14291,N_10968,N_9872);
nand U14292 (N_14292,N_11964,N_9033);
and U14293 (N_14293,N_10269,N_9397);
xnor U14294 (N_14294,N_9827,N_10080);
or U14295 (N_14295,N_11350,N_10406);
or U14296 (N_14296,N_9615,N_10613);
nand U14297 (N_14297,N_11717,N_10880);
nand U14298 (N_14298,N_10673,N_11939);
or U14299 (N_14299,N_11771,N_10338);
nor U14300 (N_14300,N_9007,N_10351);
and U14301 (N_14301,N_10052,N_9947);
nor U14302 (N_14302,N_9132,N_10008);
and U14303 (N_14303,N_10120,N_11602);
or U14304 (N_14304,N_10634,N_11772);
or U14305 (N_14305,N_10915,N_9835);
nor U14306 (N_14306,N_10419,N_10653);
or U14307 (N_14307,N_10382,N_10617);
nand U14308 (N_14308,N_11969,N_9726);
or U14309 (N_14309,N_11334,N_10684);
nand U14310 (N_14310,N_9771,N_11790);
nor U14311 (N_14311,N_9015,N_9979);
or U14312 (N_14312,N_10475,N_10067);
nor U14313 (N_14313,N_11904,N_9625);
or U14314 (N_14314,N_11907,N_9616);
and U14315 (N_14315,N_9831,N_11402);
nor U14316 (N_14316,N_9175,N_10965);
nor U14317 (N_14317,N_10877,N_10319);
nor U14318 (N_14318,N_11827,N_10670);
nor U14319 (N_14319,N_9219,N_9366);
and U14320 (N_14320,N_11551,N_11579);
nand U14321 (N_14321,N_10517,N_9350);
nor U14322 (N_14322,N_10890,N_9084);
or U14323 (N_14323,N_10119,N_9027);
nand U14324 (N_14324,N_10624,N_9858);
and U14325 (N_14325,N_11929,N_10054);
nor U14326 (N_14326,N_9418,N_9301);
and U14327 (N_14327,N_10960,N_9653);
nand U14328 (N_14328,N_10183,N_10977);
and U14329 (N_14329,N_10480,N_10168);
and U14330 (N_14330,N_9641,N_11584);
or U14331 (N_14331,N_10969,N_10195);
or U14332 (N_14332,N_10379,N_10566);
nor U14333 (N_14333,N_11705,N_10236);
or U14334 (N_14334,N_9521,N_10316);
or U14335 (N_14335,N_10378,N_11829);
nand U14336 (N_14336,N_9685,N_10774);
nand U14337 (N_14337,N_9872,N_10486);
nor U14338 (N_14338,N_11840,N_10518);
or U14339 (N_14339,N_10121,N_9628);
or U14340 (N_14340,N_10611,N_10885);
xnor U14341 (N_14341,N_9659,N_11489);
xor U14342 (N_14342,N_9167,N_10695);
nand U14343 (N_14343,N_10214,N_9575);
nor U14344 (N_14344,N_10741,N_11861);
and U14345 (N_14345,N_11823,N_10137);
and U14346 (N_14346,N_9583,N_10279);
nor U14347 (N_14347,N_10055,N_9865);
nand U14348 (N_14348,N_11003,N_10583);
nor U14349 (N_14349,N_10426,N_11877);
nor U14350 (N_14350,N_10653,N_10178);
nand U14351 (N_14351,N_9719,N_11330);
nand U14352 (N_14352,N_10271,N_9992);
and U14353 (N_14353,N_10629,N_10540);
and U14354 (N_14354,N_10979,N_10890);
nand U14355 (N_14355,N_11773,N_11379);
or U14356 (N_14356,N_9110,N_9253);
or U14357 (N_14357,N_11905,N_9077);
or U14358 (N_14358,N_9054,N_10728);
or U14359 (N_14359,N_10347,N_11260);
nand U14360 (N_14360,N_10814,N_11935);
or U14361 (N_14361,N_9164,N_9445);
nor U14362 (N_14362,N_9950,N_10548);
nand U14363 (N_14363,N_9302,N_9795);
and U14364 (N_14364,N_11840,N_10786);
nor U14365 (N_14365,N_9884,N_11160);
nand U14366 (N_14366,N_10964,N_10120);
or U14367 (N_14367,N_9572,N_11481);
or U14368 (N_14368,N_10347,N_11328);
nor U14369 (N_14369,N_9497,N_9604);
nand U14370 (N_14370,N_9966,N_10643);
and U14371 (N_14371,N_11909,N_9799);
nand U14372 (N_14372,N_9872,N_10213);
or U14373 (N_14373,N_11557,N_10342);
nor U14374 (N_14374,N_11028,N_10200);
nand U14375 (N_14375,N_10700,N_11293);
and U14376 (N_14376,N_10598,N_11402);
nor U14377 (N_14377,N_10649,N_11358);
and U14378 (N_14378,N_10083,N_9710);
or U14379 (N_14379,N_9533,N_10578);
and U14380 (N_14380,N_9570,N_10395);
nor U14381 (N_14381,N_9694,N_10171);
and U14382 (N_14382,N_10070,N_10894);
nand U14383 (N_14383,N_9735,N_11647);
and U14384 (N_14384,N_9399,N_9187);
nor U14385 (N_14385,N_11659,N_11587);
or U14386 (N_14386,N_10927,N_10330);
or U14387 (N_14387,N_9706,N_11755);
or U14388 (N_14388,N_9954,N_11343);
nor U14389 (N_14389,N_11256,N_10392);
nor U14390 (N_14390,N_11003,N_9136);
nand U14391 (N_14391,N_11499,N_9255);
nand U14392 (N_14392,N_9942,N_9743);
and U14393 (N_14393,N_11407,N_10023);
or U14394 (N_14394,N_10396,N_9823);
nor U14395 (N_14395,N_9795,N_9490);
nand U14396 (N_14396,N_10000,N_9538);
and U14397 (N_14397,N_11497,N_9150);
nand U14398 (N_14398,N_11541,N_11954);
nand U14399 (N_14399,N_11819,N_11690);
or U14400 (N_14400,N_11537,N_10799);
nor U14401 (N_14401,N_9818,N_10153);
nand U14402 (N_14402,N_11530,N_11231);
and U14403 (N_14403,N_11250,N_9110);
nand U14404 (N_14404,N_11960,N_10462);
nand U14405 (N_14405,N_9967,N_10855);
nand U14406 (N_14406,N_9144,N_10506);
nor U14407 (N_14407,N_10973,N_11993);
xor U14408 (N_14408,N_9310,N_10870);
nor U14409 (N_14409,N_11924,N_10658);
or U14410 (N_14410,N_11902,N_11652);
and U14411 (N_14411,N_10250,N_10725);
or U14412 (N_14412,N_9847,N_10511);
nand U14413 (N_14413,N_10424,N_11549);
or U14414 (N_14414,N_11644,N_11112);
nor U14415 (N_14415,N_10662,N_10793);
nand U14416 (N_14416,N_10509,N_10859);
nor U14417 (N_14417,N_9384,N_9560);
nor U14418 (N_14418,N_11772,N_10839);
xor U14419 (N_14419,N_10593,N_9605);
and U14420 (N_14420,N_9992,N_9561);
nor U14421 (N_14421,N_11380,N_11997);
or U14422 (N_14422,N_9681,N_10581);
and U14423 (N_14423,N_9892,N_10090);
nand U14424 (N_14424,N_11640,N_9219);
and U14425 (N_14425,N_10449,N_9225);
nand U14426 (N_14426,N_11427,N_9912);
nor U14427 (N_14427,N_10198,N_10827);
and U14428 (N_14428,N_10881,N_10983);
nand U14429 (N_14429,N_11501,N_9755);
nor U14430 (N_14430,N_10635,N_9780);
nand U14431 (N_14431,N_9280,N_9445);
xnor U14432 (N_14432,N_9217,N_9912);
or U14433 (N_14433,N_11135,N_9140);
or U14434 (N_14434,N_10545,N_10105);
nor U14435 (N_14435,N_11124,N_9287);
nand U14436 (N_14436,N_9790,N_9083);
or U14437 (N_14437,N_11875,N_9095);
nor U14438 (N_14438,N_9000,N_10810);
or U14439 (N_14439,N_9215,N_11041);
nor U14440 (N_14440,N_10253,N_10645);
nor U14441 (N_14441,N_10058,N_9920);
and U14442 (N_14442,N_9327,N_11007);
nor U14443 (N_14443,N_9948,N_11927);
nor U14444 (N_14444,N_10841,N_9109);
nor U14445 (N_14445,N_9904,N_9161);
nor U14446 (N_14446,N_11058,N_9680);
nand U14447 (N_14447,N_10325,N_9754);
or U14448 (N_14448,N_9869,N_9936);
nor U14449 (N_14449,N_11658,N_11560);
and U14450 (N_14450,N_9148,N_11779);
and U14451 (N_14451,N_10961,N_9624);
nand U14452 (N_14452,N_11654,N_11896);
nor U14453 (N_14453,N_9234,N_9680);
or U14454 (N_14454,N_10713,N_9746);
or U14455 (N_14455,N_9166,N_9588);
nor U14456 (N_14456,N_11411,N_11275);
and U14457 (N_14457,N_11991,N_11536);
and U14458 (N_14458,N_10574,N_11222);
nor U14459 (N_14459,N_10728,N_9666);
or U14460 (N_14460,N_10452,N_9914);
or U14461 (N_14461,N_10485,N_11486);
or U14462 (N_14462,N_11381,N_9833);
nor U14463 (N_14463,N_10304,N_10037);
or U14464 (N_14464,N_9200,N_9289);
and U14465 (N_14465,N_10077,N_11043);
or U14466 (N_14466,N_11607,N_9650);
nor U14467 (N_14467,N_9148,N_11223);
and U14468 (N_14468,N_9457,N_10770);
or U14469 (N_14469,N_11565,N_9022);
nand U14470 (N_14470,N_11594,N_10264);
nor U14471 (N_14471,N_10262,N_9810);
nand U14472 (N_14472,N_11572,N_11031);
and U14473 (N_14473,N_9351,N_9963);
and U14474 (N_14474,N_11461,N_10448);
nand U14475 (N_14475,N_9499,N_10773);
nand U14476 (N_14476,N_10256,N_11049);
nand U14477 (N_14477,N_10161,N_11090);
and U14478 (N_14478,N_9089,N_11677);
xnor U14479 (N_14479,N_11786,N_10204);
nand U14480 (N_14480,N_11865,N_10679);
and U14481 (N_14481,N_10825,N_11032);
nor U14482 (N_14482,N_11244,N_10606);
nor U14483 (N_14483,N_11408,N_11846);
nor U14484 (N_14484,N_10375,N_9642);
and U14485 (N_14485,N_9786,N_9607);
or U14486 (N_14486,N_9768,N_9677);
or U14487 (N_14487,N_9912,N_11159);
and U14488 (N_14488,N_10344,N_10272);
nand U14489 (N_14489,N_9332,N_11040);
nand U14490 (N_14490,N_9286,N_10051);
nand U14491 (N_14491,N_10084,N_11948);
nor U14492 (N_14492,N_10245,N_10798);
and U14493 (N_14493,N_11386,N_10363);
nor U14494 (N_14494,N_9688,N_11119);
or U14495 (N_14495,N_11645,N_10957);
xnor U14496 (N_14496,N_9529,N_11924);
and U14497 (N_14497,N_10273,N_11375);
nand U14498 (N_14498,N_10244,N_10446);
nand U14499 (N_14499,N_10969,N_11136);
and U14500 (N_14500,N_9630,N_10356);
nand U14501 (N_14501,N_11394,N_10541);
and U14502 (N_14502,N_9553,N_11833);
nor U14503 (N_14503,N_11117,N_10731);
xor U14504 (N_14504,N_9247,N_9731);
or U14505 (N_14505,N_11646,N_10847);
nand U14506 (N_14506,N_10099,N_9143);
or U14507 (N_14507,N_10402,N_10893);
or U14508 (N_14508,N_9409,N_10180);
nand U14509 (N_14509,N_10100,N_9955);
nor U14510 (N_14510,N_11862,N_9362);
and U14511 (N_14511,N_9770,N_10468);
nor U14512 (N_14512,N_11717,N_9780);
and U14513 (N_14513,N_10433,N_11493);
nand U14514 (N_14514,N_9740,N_11032);
or U14515 (N_14515,N_10551,N_9806);
or U14516 (N_14516,N_11199,N_10720);
and U14517 (N_14517,N_9388,N_9311);
and U14518 (N_14518,N_11170,N_10220);
nand U14519 (N_14519,N_10105,N_11955);
nor U14520 (N_14520,N_9609,N_10603);
nor U14521 (N_14521,N_10956,N_9446);
or U14522 (N_14522,N_10120,N_11798);
and U14523 (N_14523,N_9329,N_10419);
nand U14524 (N_14524,N_11981,N_11243);
or U14525 (N_14525,N_10471,N_9502);
or U14526 (N_14526,N_10515,N_9520);
and U14527 (N_14527,N_11709,N_11201);
nor U14528 (N_14528,N_10364,N_11694);
and U14529 (N_14529,N_9301,N_9415);
and U14530 (N_14530,N_11923,N_10280);
nand U14531 (N_14531,N_11854,N_11992);
nand U14532 (N_14532,N_10663,N_9571);
and U14533 (N_14533,N_10035,N_10805);
or U14534 (N_14534,N_11698,N_9696);
and U14535 (N_14535,N_10204,N_9692);
nor U14536 (N_14536,N_9228,N_10847);
and U14537 (N_14537,N_10569,N_9888);
or U14538 (N_14538,N_11809,N_11383);
nor U14539 (N_14539,N_9779,N_11590);
and U14540 (N_14540,N_11437,N_9559);
and U14541 (N_14541,N_10304,N_11319);
xor U14542 (N_14542,N_10500,N_9051);
nor U14543 (N_14543,N_11498,N_11453);
or U14544 (N_14544,N_11358,N_10163);
nor U14545 (N_14545,N_9499,N_10579);
and U14546 (N_14546,N_11957,N_11106);
nor U14547 (N_14547,N_9400,N_10550);
and U14548 (N_14548,N_9128,N_9484);
or U14549 (N_14549,N_11467,N_10352);
and U14550 (N_14550,N_9546,N_10659);
and U14551 (N_14551,N_9063,N_11743);
or U14552 (N_14552,N_10986,N_11167);
nor U14553 (N_14553,N_10759,N_11897);
nand U14554 (N_14554,N_9347,N_10141);
or U14555 (N_14555,N_10836,N_9165);
nor U14556 (N_14556,N_9603,N_9854);
nor U14557 (N_14557,N_9653,N_10363);
and U14558 (N_14558,N_11223,N_9789);
nor U14559 (N_14559,N_9787,N_9140);
nor U14560 (N_14560,N_11974,N_10856);
nor U14561 (N_14561,N_10893,N_10876);
nand U14562 (N_14562,N_11104,N_11154);
nor U14563 (N_14563,N_10586,N_9238);
nor U14564 (N_14564,N_9376,N_9477);
and U14565 (N_14565,N_9914,N_9525);
nand U14566 (N_14566,N_9470,N_10160);
nand U14567 (N_14567,N_9854,N_11184);
and U14568 (N_14568,N_11485,N_10578);
nand U14569 (N_14569,N_11362,N_10123);
nor U14570 (N_14570,N_10487,N_11272);
nor U14571 (N_14571,N_9681,N_10286);
nand U14572 (N_14572,N_11094,N_9603);
or U14573 (N_14573,N_9875,N_11491);
nand U14574 (N_14574,N_10873,N_9457);
nor U14575 (N_14575,N_10220,N_10449);
or U14576 (N_14576,N_10035,N_10853);
and U14577 (N_14577,N_10331,N_9411);
and U14578 (N_14578,N_10636,N_9525);
nand U14579 (N_14579,N_9894,N_11834);
and U14580 (N_14580,N_9584,N_10558);
nor U14581 (N_14581,N_10188,N_9550);
and U14582 (N_14582,N_10460,N_9996);
nor U14583 (N_14583,N_10989,N_10570);
and U14584 (N_14584,N_10298,N_10242);
or U14585 (N_14585,N_11167,N_10651);
nand U14586 (N_14586,N_11564,N_9789);
and U14587 (N_14587,N_11920,N_9996);
or U14588 (N_14588,N_9928,N_11649);
nor U14589 (N_14589,N_11126,N_9640);
nor U14590 (N_14590,N_9821,N_10203);
nand U14591 (N_14591,N_9663,N_9232);
nand U14592 (N_14592,N_10990,N_10054);
nor U14593 (N_14593,N_10799,N_10873);
nand U14594 (N_14594,N_10163,N_10850);
nand U14595 (N_14595,N_10357,N_11003);
nand U14596 (N_14596,N_10337,N_10375);
nor U14597 (N_14597,N_11840,N_11352);
nand U14598 (N_14598,N_11274,N_9413);
and U14599 (N_14599,N_11571,N_11738);
nor U14600 (N_14600,N_11367,N_11993);
and U14601 (N_14601,N_10951,N_11239);
or U14602 (N_14602,N_11803,N_11862);
and U14603 (N_14603,N_11362,N_10922);
and U14604 (N_14604,N_9992,N_11214);
or U14605 (N_14605,N_11113,N_9879);
nand U14606 (N_14606,N_11477,N_10307);
or U14607 (N_14607,N_9232,N_9072);
or U14608 (N_14608,N_9798,N_9445);
nor U14609 (N_14609,N_11643,N_9467);
or U14610 (N_14610,N_10002,N_11001);
nand U14611 (N_14611,N_10230,N_10768);
or U14612 (N_14612,N_9999,N_11272);
or U14613 (N_14613,N_11347,N_9592);
nor U14614 (N_14614,N_10967,N_11900);
nand U14615 (N_14615,N_9771,N_11139);
nor U14616 (N_14616,N_11451,N_10877);
or U14617 (N_14617,N_9318,N_9003);
xnor U14618 (N_14618,N_11678,N_10508);
nand U14619 (N_14619,N_10425,N_11994);
nand U14620 (N_14620,N_10940,N_9433);
nor U14621 (N_14621,N_11720,N_9172);
and U14622 (N_14622,N_10458,N_9531);
or U14623 (N_14623,N_9866,N_10318);
or U14624 (N_14624,N_10189,N_9070);
or U14625 (N_14625,N_11985,N_10068);
nand U14626 (N_14626,N_9237,N_10845);
or U14627 (N_14627,N_9345,N_10014);
or U14628 (N_14628,N_11357,N_9005);
and U14629 (N_14629,N_11850,N_11593);
nor U14630 (N_14630,N_11194,N_11838);
and U14631 (N_14631,N_11594,N_10397);
nor U14632 (N_14632,N_11730,N_11172);
or U14633 (N_14633,N_9747,N_10392);
nand U14634 (N_14634,N_11012,N_11006);
xnor U14635 (N_14635,N_10922,N_9703);
nand U14636 (N_14636,N_10839,N_9657);
nand U14637 (N_14637,N_10967,N_11517);
and U14638 (N_14638,N_11304,N_10860);
nor U14639 (N_14639,N_9046,N_10080);
or U14640 (N_14640,N_9691,N_9830);
nand U14641 (N_14641,N_9701,N_9818);
and U14642 (N_14642,N_11694,N_10332);
nand U14643 (N_14643,N_11598,N_10315);
or U14644 (N_14644,N_9698,N_11757);
nand U14645 (N_14645,N_10923,N_10605);
nor U14646 (N_14646,N_10450,N_9216);
nor U14647 (N_14647,N_10100,N_11388);
and U14648 (N_14648,N_10848,N_10758);
xnor U14649 (N_14649,N_11796,N_10326);
or U14650 (N_14650,N_11361,N_9425);
or U14651 (N_14651,N_11739,N_9939);
nand U14652 (N_14652,N_11470,N_11018);
nor U14653 (N_14653,N_11162,N_11230);
nor U14654 (N_14654,N_9948,N_11831);
nor U14655 (N_14655,N_10166,N_9916);
or U14656 (N_14656,N_9371,N_11737);
and U14657 (N_14657,N_11053,N_11761);
nor U14658 (N_14658,N_11833,N_9253);
nand U14659 (N_14659,N_11566,N_11169);
and U14660 (N_14660,N_10674,N_11918);
or U14661 (N_14661,N_11408,N_9368);
and U14662 (N_14662,N_10522,N_11919);
nor U14663 (N_14663,N_11622,N_11221);
xnor U14664 (N_14664,N_11517,N_9385);
nor U14665 (N_14665,N_9678,N_10706);
nand U14666 (N_14666,N_10736,N_10216);
nand U14667 (N_14667,N_11088,N_10078);
or U14668 (N_14668,N_11259,N_9511);
or U14669 (N_14669,N_10496,N_11475);
nand U14670 (N_14670,N_9848,N_10630);
nand U14671 (N_14671,N_10073,N_10382);
and U14672 (N_14672,N_11379,N_10421);
nand U14673 (N_14673,N_9805,N_11104);
nor U14674 (N_14674,N_9815,N_10294);
nand U14675 (N_14675,N_11257,N_9017);
nand U14676 (N_14676,N_11760,N_11904);
and U14677 (N_14677,N_10321,N_10531);
nor U14678 (N_14678,N_10291,N_9677);
nor U14679 (N_14679,N_11502,N_10285);
and U14680 (N_14680,N_10503,N_10790);
nand U14681 (N_14681,N_10039,N_9899);
or U14682 (N_14682,N_11612,N_9107);
xor U14683 (N_14683,N_10142,N_11934);
nand U14684 (N_14684,N_9429,N_10387);
nand U14685 (N_14685,N_9834,N_9605);
and U14686 (N_14686,N_10083,N_9219);
or U14687 (N_14687,N_10477,N_9708);
and U14688 (N_14688,N_10346,N_10155);
and U14689 (N_14689,N_10842,N_11671);
or U14690 (N_14690,N_11505,N_10118);
nand U14691 (N_14691,N_9039,N_9985);
or U14692 (N_14692,N_10620,N_11675);
nand U14693 (N_14693,N_9000,N_10683);
or U14694 (N_14694,N_10633,N_11781);
and U14695 (N_14695,N_10728,N_9677);
and U14696 (N_14696,N_11368,N_11281);
or U14697 (N_14697,N_11199,N_10677);
or U14698 (N_14698,N_10922,N_11878);
xor U14699 (N_14699,N_11657,N_10350);
nor U14700 (N_14700,N_11564,N_9044);
nand U14701 (N_14701,N_10824,N_10617);
nor U14702 (N_14702,N_10661,N_9585);
nand U14703 (N_14703,N_9158,N_9405);
and U14704 (N_14704,N_9795,N_9220);
nor U14705 (N_14705,N_10967,N_10655);
and U14706 (N_14706,N_9776,N_10900);
nand U14707 (N_14707,N_9237,N_9163);
nand U14708 (N_14708,N_10787,N_11026);
and U14709 (N_14709,N_9885,N_10402);
or U14710 (N_14710,N_9692,N_11458);
nor U14711 (N_14711,N_9690,N_10068);
or U14712 (N_14712,N_10952,N_11611);
or U14713 (N_14713,N_10544,N_11469);
and U14714 (N_14714,N_9721,N_10713);
nor U14715 (N_14715,N_11721,N_10499);
xnor U14716 (N_14716,N_10836,N_9952);
nor U14717 (N_14717,N_9151,N_10309);
or U14718 (N_14718,N_10631,N_10608);
nor U14719 (N_14719,N_10523,N_9483);
nor U14720 (N_14720,N_10464,N_10513);
nand U14721 (N_14721,N_9074,N_9849);
or U14722 (N_14722,N_9913,N_11709);
or U14723 (N_14723,N_10759,N_10244);
nor U14724 (N_14724,N_10571,N_10081);
or U14725 (N_14725,N_10116,N_9448);
nand U14726 (N_14726,N_11024,N_9086);
nand U14727 (N_14727,N_9372,N_9353);
nand U14728 (N_14728,N_9370,N_9540);
or U14729 (N_14729,N_9042,N_10083);
nor U14730 (N_14730,N_9980,N_10220);
xor U14731 (N_14731,N_9074,N_10128);
or U14732 (N_14732,N_10176,N_10178);
xnor U14733 (N_14733,N_9084,N_9177);
or U14734 (N_14734,N_11088,N_10907);
nor U14735 (N_14735,N_9296,N_10271);
nor U14736 (N_14736,N_10362,N_10251);
or U14737 (N_14737,N_9964,N_9384);
nor U14738 (N_14738,N_9099,N_9012);
nand U14739 (N_14739,N_9407,N_11329);
or U14740 (N_14740,N_10432,N_10497);
and U14741 (N_14741,N_10979,N_9438);
or U14742 (N_14742,N_10913,N_9523);
nor U14743 (N_14743,N_11150,N_11624);
nor U14744 (N_14744,N_9634,N_11330);
or U14745 (N_14745,N_9034,N_10324);
nand U14746 (N_14746,N_9942,N_9087);
nand U14747 (N_14747,N_10249,N_10359);
and U14748 (N_14748,N_11010,N_11585);
and U14749 (N_14749,N_10393,N_10045);
nor U14750 (N_14750,N_11386,N_11608);
nand U14751 (N_14751,N_10467,N_11869);
xor U14752 (N_14752,N_10801,N_9685);
nor U14753 (N_14753,N_9635,N_11615);
xor U14754 (N_14754,N_11448,N_11382);
nor U14755 (N_14755,N_10007,N_9552);
or U14756 (N_14756,N_10352,N_11155);
or U14757 (N_14757,N_9578,N_9829);
or U14758 (N_14758,N_10945,N_10557);
nor U14759 (N_14759,N_9995,N_11922);
nand U14760 (N_14760,N_9366,N_9623);
or U14761 (N_14761,N_10785,N_11530);
nand U14762 (N_14762,N_10160,N_9913);
or U14763 (N_14763,N_10888,N_10480);
and U14764 (N_14764,N_11751,N_11807);
and U14765 (N_14765,N_9927,N_9910);
or U14766 (N_14766,N_10763,N_11116);
nand U14767 (N_14767,N_9519,N_11111);
nand U14768 (N_14768,N_11053,N_11428);
nand U14769 (N_14769,N_10876,N_11423);
nand U14770 (N_14770,N_10380,N_9417);
or U14771 (N_14771,N_9497,N_11430);
nor U14772 (N_14772,N_9651,N_10520);
nand U14773 (N_14773,N_10680,N_9933);
nand U14774 (N_14774,N_11348,N_9384);
nand U14775 (N_14775,N_9602,N_10778);
or U14776 (N_14776,N_11930,N_10288);
nor U14777 (N_14777,N_10703,N_11092);
nand U14778 (N_14778,N_9334,N_10950);
or U14779 (N_14779,N_11952,N_9029);
nand U14780 (N_14780,N_10593,N_10744);
nor U14781 (N_14781,N_9990,N_9192);
nor U14782 (N_14782,N_9351,N_10123);
nor U14783 (N_14783,N_9956,N_11151);
nor U14784 (N_14784,N_9920,N_11991);
or U14785 (N_14785,N_9254,N_11505);
or U14786 (N_14786,N_11876,N_11242);
and U14787 (N_14787,N_11604,N_10473);
or U14788 (N_14788,N_11136,N_10357);
and U14789 (N_14789,N_9542,N_9614);
and U14790 (N_14790,N_9420,N_9058);
or U14791 (N_14791,N_10740,N_9759);
nor U14792 (N_14792,N_9951,N_10299);
nor U14793 (N_14793,N_9673,N_10388);
nor U14794 (N_14794,N_10510,N_10866);
and U14795 (N_14795,N_10765,N_10398);
nand U14796 (N_14796,N_10031,N_10585);
nand U14797 (N_14797,N_10443,N_10554);
nor U14798 (N_14798,N_9527,N_11757);
nand U14799 (N_14799,N_10113,N_9376);
nor U14800 (N_14800,N_9475,N_11969);
or U14801 (N_14801,N_10572,N_9062);
or U14802 (N_14802,N_11434,N_10251);
or U14803 (N_14803,N_10114,N_9721);
or U14804 (N_14804,N_11943,N_10916);
and U14805 (N_14805,N_11185,N_11861);
nand U14806 (N_14806,N_11927,N_10212);
nand U14807 (N_14807,N_10685,N_9499);
nand U14808 (N_14808,N_10065,N_10324);
nand U14809 (N_14809,N_9891,N_10508);
nand U14810 (N_14810,N_11452,N_10352);
nor U14811 (N_14811,N_11864,N_9804);
nor U14812 (N_14812,N_11733,N_11658);
nor U14813 (N_14813,N_9599,N_10726);
nor U14814 (N_14814,N_9311,N_9618);
nor U14815 (N_14815,N_10538,N_11079);
xnor U14816 (N_14816,N_9225,N_9555);
nand U14817 (N_14817,N_10495,N_9041);
and U14818 (N_14818,N_10317,N_9977);
or U14819 (N_14819,N_11251,N_10551);
nand U14820 (N_14820,N_11541,N_9897);
or U14821 (N_14821,N_9507,N_9305);
nand U14822 (N_14822,N_10275,N_11818);
nor U14823 (N_14823,N_9036,N_9150);
nor U14824 (N_14824,N_11490,N_9005);
or U14825 (N_14825,N_11028,N_10980);
nor U14826 (N_14826,N_9737,N_11500);
nor U14827 (N_14827,N_9835,N_11516);
or U14828 (N_14828,N_9719,N_10862);
and U14829 (N_14829,N_9388,N_9165);
nand U14830 (N_14830,N_9799,N_10108);
nor U14831 (N_14831,N_9289,N_11356);
nor U14832 (N_14832,N_9331,N_10517);
or U14833 (N_14833,N_9998,N_9789);
nand U14834 (N_14834,N_11881,N_10565);
nand U14835 (N_14835,N_11373,N_11011);
and U14836 (N_14836,N_10301,N_9729);
nand U14837 (N_14837,N_11788,N_10999);
nand U14838 (N_14838,N_11593,N_11244);
and U14839 (N_14839,N_10930,N_9708);
nand U14840 (N_14840,N_9930,N_10626);
nor U14841 (N_14841,N_10232,N_9743);
or U14842 (N_14842,N_11001,N_10652);
and U14843 (N_14843,N_10292,N_10730);
or U14844 (N_14844,N_10927,N_10115);
and U14845 (N_14845,N_11692,N_11593);
or U14846 (N_14846,N_9654,N_11171);
nand U14847 (N_14847,N_11022,N_9991);
nand U14848 (N_14848,N_9137,N_10113);
or U14849 (N_14849,N_10519,N_9057);
and U14850 (N_14850,N_11273,N_9618);
and U14851 (N_14851,N_9531,N_10248);
nand U14852 (N_14852,N_11536,N_9102);
nand U14853 (N_14853,N_11763,N_10971);
nor U14854 (N_14854,N_11995,N_10856);
or U14855 (N_14855,N_9495,N_10607);
nor U14856 (N_14856,N_9076,N_9458);
nor U14857 (N_14857,N_9572,N_11976);
nor U14858 (N_14858,N_10162,N_11798);
nor U14859 (N_14859,N_9837,N_11223);
nor U14860 (N_14860,N_9645,N_9006);
or U14861 (N_14861,N_11421,N_10482);
or U14862 (N_14862,N_9573,N_11617);
and U14863 (N_14863,N_11620,N_11546);
and U14864 (N_14864,N_10030,N_11808);
nor U14865 (N_14865,N_11592,N_11066);
xnor U14866 (N_14866,N_10938,N_11595);
or U14867 (N_14867,N_9635,N_9290);
nor U14868 (N_14868,N_11766,N_9082);
and U14869 (N_14869,N_9963,N_11609);
nor U14870 (N_14870,N_10928,N_9433);
and U14871 (N_14871,N_11445,N_11561);
nand U14872 (N_14872,N_10631,N_9327);
and U14873 (N_14873,N_10289,N_11579);
nor U14874 (N_14874,N_10836,N_9030);
nand U14875 (N_14875,N_9073,N_10392);
or U14876 (N_14876,N_9110,N_10565);
nand U14877 (N_14877,N_10810,N_9873);
nand U14878 (N_14878,N_11265,N_11580);
nand U14879 (N_14879,N_11887,N_9248);
and U14880 (N_14880,N_9931,N_11632);
xnor U14881 (N_14881,N_10684,N_10642);
nor U14882 (N_14882,N_10303,N_9244);
xnor U14883 (N_14883,N_10023,N_10728);
and U14884 (N_14884,N_11342,N_9252);
nor U14885 (N_14885,N_10894,N_11302);
or U14886 (N_14886,N_11795,N_9487);
and U14887 (N_14887,N_10962,N_10229);
or U14888 (N_14888,N_11662,N_10703);
xor U14889 (N_14889,N_11284,N_9532);
nand U14890 (N_14890,N_10660,N_11116);
nand U14891 (N_14891,N_9710,N_9837);
xor U14892 (N_14892,N_9173,N_11730);
or U14893 (N_14893,N_10744,N_11409);
nand U14894 (N_14894,N_10008,N_9239);
nor U14895 (N_14895,N_10723,N_10151);
nand U14896 (N_14896,N_11480,N_11992);
nand U14897 (N_14897,N_10627,N_11394);
or U14898 (N_14898,N_9290,N_11809);
and U14899 (N_14899,N_10262,N_9019);
nand U14900 (N_14900,N_11651,N_9677);
and U14901 (N_14901,N_11638,N_10373);
nand U14902 (N_14902,N_11337,N_10368);
nand U14903 (N_14903,N_11531,N_10840);
nand U14904 (N_14904,N_9036,N_10920);
nand U14905 (N_14905,N_10866,N_11840);
and U14906 (N_14906,N_10466,N_11974);
and U14907 (N_14907,N_10789,N_9666);
nand U14908 (N_14908,N_11490,N_10235);
or U14909 (N_14909,N_11950,N_10439);
or U14910 (N_14910,N_9085,N_9784);
nand U14911 (N_14911,N_9054,N_10426);
and U14912 (N_14912,N_11111,N_9611);
or U14913 (N_14913,N_11820,N_10893);
or U14914 (N_14914,N_11377,N_10898);
and U14915 (N_14915,N_9100,N_9660);
nand U14916 (N_14916,N_10447,N_10124);
nor U14917 (N_14917,N_11863,N_11823);
or U14918 (N_14918,N_11137,N_11740);
nand U14919 (N_14919,N_9654,N_11769);
nand U14920 (N_14920,N_10681,N_10395);
and U14921 (N_14921,N_11135,N_10171);
nor U14922 (N_14922,N_11962,N_9353);
nand U14923 (N_14923,N_10534,N_11684);
nand U14924 (N_14924,N_10620,N_11192);
nor U14925 (N_14925,N_9398,N_11898);
or U14926 (N_14926,N_9095,N_9921);
nand U14927 (N_14927,N_10343,N_9118);
or U14928 (N_14928,N_10004,N_11207);
and U14929 (N_14929,N_11714,N_9271);
or U14930 (N_14930,N_9753,N_9473);
xnor U14931 (N_14931,N_11247,N_11996);
nor U14932 (N_14932,N_10762,N_11100);
nor U14933 (N_14933,N_9472,N_9026);
or U14934 (N_14934,N_9147,N_11739);
and U14935 (N_14935,N_10982,N_10290);
and U14936 (N_14936,N_9968,N_10204);
nand U14937 (N_14937,N_10025,N_11415);
and U14938 (N_14938,N_10838,N_9817);
nor U14939 (N_14939,N_9204,N_9807);
and U14940 (N_14940,N_10200,N_9340);
nand U14941 (N_14941,N_11340,N_11192);
nor U14942 (N_14942,N_11027,N_9460);
or U14943 (N_14943,N_11105,N_11751);
or U14944 (N_14944,N_11852,N_11235);
and U14945 (N_14945,N_10348,N_11662);
or U14946 (N_14946,N_10864,N_11459);
or U14947 (N_14947,N_10666,N_11953);
nand U14948 (N_14948,N_9103,N_10298);
nor U14949 (N_14949,N_10414,N_10022);
or U14950 (N_14950,N_9081,N_10055);
nor U14951 (N_14951,N_11552,N_9894);
nor U14952 (N_14952,N_9574,N_10128);
nand U14953 (N_14953,N_9649,N_10865);
or U14954 (N_14954,N_9040,N_9341);
and U14955 (N_14955,N_10175,N_10622);
nor U14956 (N_14956,N_10132,N_9216);
nand U14957 (N_14957,N_9088,N_9332);
nand U14958 (N_14958,N_10268,N_10944);
and U14959 (N_14959,N_10537,N_10475);
nand U14960 (N_14960,N_11930,N_11371);
or U14961 (N_14961,N_11814,N_11379);
and U14962 (N_14962,N_9654,N_11035);
nor U14963 (N_14963,N_9425,N_11964);
nand U14964 (N_14964,N_10158,N_10697);
nor U14965 (N_14965,N_9085,N_11043);
and U14966 (N_14966,N_10327,N_9935);
and U14967 (N_14967,N_10457,N_10504);
nand U14968 (N_14968,N_9140,N_10711);
and U14969 (N_14969,N_9521,N_11585);
nand U14970 (N_14970,N_10045,N_10307);
or U14971 (N_14971,N_10501,N_9518);
nor U14972 (N_14972,N_10999,N_11050);
and U14973 (N_14973,N_11031,N_10637);
nand U14974 (N_14974,N_9244,N_11181);
and U14975 (N_14975,N_11288,N_10083);
or U14976 (N_14976,N_9165,N_9193);
and U14977 (N_14977,N_9586,N_9958);
nor U14978 (N_14978,N_10422,N_9951);
xor U14979 (N_14979,N_9536,N_10234);
or U14980 (N_14980,N_11362,N_9889);
or U14981 (N_14981,N_10554,N_10155);
and U14982 (N_14982,N_11406,N_9841);
or U14983 (N_14983,N_11548,N_11446);
nand U14984 (N_14984,N_9898,N_10337);
nor U14985 (N_14985,N_11862,N_11672);
nor U14986 (N_14986,N_9482,N_11105);
nor U14987 (N_14987,N_10162,N_11396);
nor U14988 (N_14988,N_9936,N_9635);
nor U14989 (N_14989,N_10672,N_10623);
or U14990 (N_14990,N_10837,N_9283);
nand U14991 (N_14991,N_9496,N_9884);
nand U14992 (N_14992,N_9058,N_11930);
or U14993 (N_14993,N_10394,N_9051);
nand U14994 (N_14994,N_9933,N_10731);
nand U14995 (N_14995,N_9661,N_11195);
nor U14996 (N_14996,N_10552,N_9266);
nor U14997 (N_14997,N_10005,N_11973);
xor U14998 (N_14998,N_11553,N_9421);
nand U14999 (N_14999,N_11587,N_10322);
nand UO_0 (O_0,N_14848,N_12741);
or UO_1 (O_1,N_13356,N_13616);
nor UO_2 (O_2,N_14014,N_13351);
nor UO_3 (O_3,N_14040,N_14179);
nor UO_4 (O_4,N_14917,N_14464);
nand UO_5 (O_5,N_13859,N_14258);
or UO_6 (O_6,N_13709,N_13358);
and UO_7 (O_7,N_12997,N_14494);
and UO_8 (O_8,N_13460,N_13874);
and UO_9 (O_9,N_13715,N_14475);
nand UO_10 (O_10,N_13169,N_13735);
or UO_11 (O_11,N_12126,N_14134);
xnor UO_12 (O_12,N_13367,N_13397);
nor UO_13 (O_13,N_13852,N_12395);
or UO_14 (O_14,N_12453,N_14244);
and UO_15 (O_15,N_13311,N_14586);
or UO_16 (O_16,N_14838,N_13039);
and UO_17 (O_17,N_14057,N_12269);
xor UO_18 (O_18,N_12617,N_12384);
or UO_19 (O_19,N_12522,N_13557);
nand UO_20 (O_20,N_13834,N_13643);
nor UO_21 (O_21,N_14532,N_13524);
xnor UO_22 (O_22,N_14441,N_14807);
nor UO_23 (O_23,N_14166,N_13334);
or UO_24 (O_24,N_14026,N_13307);
and UO_25 (O_25,N_12586,N_12454);
or UO_26 (O_26,N_14403,N_13336);
nor UO_27 (O_27,N_12035,N_14962);
nand UO_28 (O_28,N_14619,N_13604);
and UO_29 (O_29,N_13193,N_12762);
or UO_30 (O_30,N_12002,N_12468);
and UO_31 (O_31,N_14027,N_12447);
nor UO_32 (O_32,N_13914,N_13851);
and UO_33 (O_33,N_14161,N_12921);
nor UO_34 (O_34,N_13274,N_13077);
or UO_35 (O_35,N_13236,N_13017);
xor UO_36 (O_36,N_12974,N_12543);
and UO_37 (O_37,N_12017,N_12072);
nand UO_38 (O_38,N_14017,N_13197);
xnor UO_39 (O_39,N_13386,N_13092);
and UO_40 (O_40,N_12399,N_14183);
and UO_41 (O_41,N_13015,N_13510);
or UO_42 (O_42,N_14110,N_12808);
nand UO_43 (O_43,N_13498,N_13620);
nor UO_44 (O_44,N_13313,N_14467);
nand UO_45 (O_45,N_14685,N_12583);
nor UO_46 (O_46,N_13123,N_12070);
nor UO_47 (O_47,N_13088,N_12960);
and UO_48 (O_48,N_13467,N_12923);
nor UO_49 (O_49,N_12445,N_12702);
nand UO_50 (O_50,N_13479,N_13728);
nand UO_51 (O_51,N_14601,N_14985);
and UO_52 (O_52,N_13127,N_14319);
xnor UO_53 (O_53,N_13869,N_13907);
and UO_54 (O_54,N_14856,N_13565);
nand UO_55 (O_55,N_13182,N_13624);
nor UO_56 (O_56,N_13014,N_13840);
and UO_57 (O_57,N_14377,N_12486);
nand UO_58 (O_58,N_12860,N_14004);
or UO_59 (O_59,N_13156,N_12416);
or UO_60 (O_60,N_14018,N_13585);
or UO_61 (O_61,N_13960,N_14140);
and UO_62 (O_62,N_12517,N_12292);
nand UO_63 (O_63,N_12450,N_12278);
nand UO_64 (O_64,N_14331,N_12356);
nor UO_65 (O_65,N_12761,N_13913);
or UO_66 (O_66,N_13848,N_14501);
nand UO_67 (O_67,N_12625,N_12461);
and UO_68 (O_68,N_14021,N_13543);
or UO_69 (O_69,N_14311,N_13372);
nand UO_70 (O_70,N_13879,N_13833);
nor UO_71 (O_71,N_12966,N_14710);
or UO_72 (O_72,N_14712,N_13876);
xnor UO_73 (O_73,N_13562,N_13005);
and UO_74 (O_74,N_14661,N_14096);
or UO_75 (O_75,N_14681,N_12707);
and UO_76 (O_76,N_12826,N_12493);
and UO_77 (O_77,N_14785,N_12571);
nand UO_78 (O_78,N_13591,N_14776);
nand UO_79 (O_79,N_14256,N_13312);
and UO_80 (O_80,N_13207,N_13955);
nand UO_81 (O_81,N_12089,N_14976);
nor UO_82 (O_82,N_14405,N_12553);
or UO_83 (O_83,N_13481,N_14500);
nor UO_84 (O_84,N_14880,N_12955);
nand UO_85 (O_85,N_12652,N_12411);
nand UO_86 (O_86,N_14176,N_12638);
nor UO_87 (O_87,N_14059,N_13699);
nand UO_88 (O_88,N_13011,N_14382);
or UO_89 (O_89,N_12773,N_14580);
and UO_90 (O_90,N_14024,N_14704);
nor UO_91 (O_91,N_12909,N_13959);
nand UO_92 (O_92,N_12908,N_14297);
nor UO_93 (O_93,N_14592,N_14349);
nor UO_94 (O_94,N_13373,N_14939);
or UO_95 (O_95,N_14468,N_12112);
nand UO_96 (O_96,N_13910,N_12154);
and UO_97 (O_97,N_14427,N_12791);
nand UO_98 (O_98,N_13502,N_12358);
or UO_99 (O_99,N_14859,N_13981);
or UO_100 (O_100,N_13359,N_14511);
nand UO_101 (O_101,N_13215,N_14060);
nand UO_102 (O_102,N_13819,N_13789);
and UO_103 (O_103,N_13211,N_13300);
nand UO_104 (O_104,N_14127,N_12958);
nor UO_105 (O_105,N_13668,N_12579);
nand UO_106 (O_106,N_12827,N_14509);
and UO_107 (O_107,N_12385,N_14247);
nor UO_108 (O_108,N_14625,N_13820);
or UO_109 (O_109,N_13976,N_13561);
nor UO_110 (O_110,N_13506,N_12363);
and UO_111 (O_111,N_14058,N_14101);
or UO_112 (O_112,N_14341,N_14368);
and UO_113 (O_113,N_13657,N_14044);
nand UO_114 (O_114,N_13887,N_12614);
or UO_115 (O_115,N_13554,N_14234);
nand UO_116 (O_116,N_13905,N_12498);
nor UO_117 (O_117,N_13035,N_14932);
or UO_118 (O_118,N_13245,N_12813);
and UO_119 (O_119,N_14037,N_14913);
or UO_120 (O_120,N_14156,N_13755);
and UO_121 (O_121,N_14690,N_13726);
or UO_122 (O_122,N_14524,N_12423);
or UO_123 (O_123,N_14440,N_14684);
nor UO_124 (O_124,N_12562,N_13984);
or UO_125 (O_125,N_14235,N_12731);
nor UO_126 (O_126,N_13314,N_13575);
or UO_127 (O_127,N_13155,N_14131);
nor UO_128 (O_128,N_13476,N_14766);
nor UO_129 (O_129,N_12781,N_12687);
and UO_130 (O_130,N_13007,N_14790);
nor UO_131 (O_131,N_12609,N_14142);
and UO_132 (O_132,N_14143,N_12206);
and UO_133 (O_133,N_13908,N_13031);
nand UO_134 (O_134,N_14715,N_14857);
and UO_135 (O_135,N_12194,N_14695);
xor UO_136 (O_136,N_13553,N_13244);
or UO_137 (O_137,N_14056,N_12108);
and UO_138 (O_138,N_13399,N_14437);
and UO_139 (O_139,N_14254,N_14718);
and UO_140 (O_140,N_14150,N_14320);
nand UO_141 (O_141,N_14181,N_14279);
nor UO_142 (O_142,N_14429,N_14914);
and UO_143 (O_143,N_14608,N_14097);
nand UO_144 (O_144,N_14184,N_12936);
nor UO_145 (O_145,N_14599,N_13809);
nand UO_146 (O_146,N_13754,N_13600);
nor UO_147 (O_147,N_12366,N_13332);
and UO_148 (O_148,N_14365,N_12256);
nor UO_149 (O_149,N_14805,N_12326);
nand UO_150 (O_150,N_14086,N_14151);
and UO_151 (O_151,N_12729,N_14424);
nor UO_152 (O_152,N_13394,N_14271);
nor UO_153 (O_153,N_13341,N_12444);
and UO_154 (O_154,N_14222,N_14781);
nor UO_155 (O_155,N_13566,N_12127);
nor UO_156 (O_156,N_14774,N_12115);
or UO_157 (O_157,N_13659,N_12643);
and UO_158 (O_158,N_12176,N_13945);
and UO_159 (O_159,N_12215,N_14650);
or UO_160 (O_160,N_12146,N_13527);
and UO_161 (O_161,N_14470,N_12787);
and UO_162 (O_162,N_13781,N_12959);
nand UO_163 (O_163,N_14460,N_14725);
nor UO_164 (O_164,N_13004,N_14313);
or UO_165 (O_165,N_12196,N_14616);
nand UO_166 (O_166,N_12408,N_14687);
and UO_167 (O_167,N_13603,N_14105);
or UO_168 (O_168,N_14361,N_13634);
nand UO_169 (O_169,N_12873,N_13760);
nand UO_170 (O_170,N_12598,N_12841);
nor UO_171 (O_171,N_12979,N_14832);
and UO_172 (O_172,N_13222,N_13783);
nand UO_173 (O_173,N_14066,N_14287);
nor UO_174 (O_174,N_13714,N_12203);
nand UO_175 (O_175,N_13390,N_13445);
nor UO_176 (O_176,N_12412,N_14770);
nor UO_177 (O_177,N_14545,N_12043);
nand UO_178 (O_178,N_12796,N_14345);
and UO_179 (O_179,N_14121,N_13267);
and UO_180 (O_180,N_13224,N_12172);
nor UO_181 (O_181,N_12136,N_13720);
nor UO_182 (O_182,N_14485,N_14321);
nor UO_183 (O_183,N_13214,N_12480);
and UO_184 (O_184,N_14051,N_14623);
nor UO_185 (O_185,N_12164,N_12510);
nor UO_186 (O_186,N_12299,N_14339);
and UO_187 (O_187,N_13650,N_14232);
nand UO_188 (O_188,N_13271,N_12852);
nor UO_189 (O_189,N_14386,N_14617);
or UO_190 (O_190,N_12495,N_12749);
or UO_191 (O_191,N_12396,N_13348);
nand UO_192 (O_192,N_13325,N_14493);
or UO_193 (O_193,N_12027,N_12537);
nand UO_194 (O_194,N_14771,N_12378);
nor UO_195 (O_195,N_13990,N_12390);
or UO_196 (O_196,N_13582,N_12700);
or UO_197 (O_197,N_13791,N_13084);
nor UO_198 (O_198,N_12184,N_14230);
and UO_199 (O_199,N_13891,N_12050);
and UO_200 (O_200,N_14553,N_12946);
and UO_201 (O_201,N_12353,N_13592);
nor UO_202 (O_202,N_12077,N_12306);
or UO_203 (O_203,N_14828,N_12381);
nand UO_204 (O_204,N_13822,N_14558);
nor UO_205 (O_205,N_12300,N_12418);
or UO_206 (O_206,N_12682,N_13395);
and UO_207 (O_207,N_13044,N_12587);
xnor UO_208 (O_208,N_14399,N_12785);
nor UO_209 (O_209,N_12573,N_12446);
nand UO_210 (O_210,N_13861,N_13166);
nor UO_211 (O_211,N_12636,N_14251);
and UO_212 (O_212,N_14190,N_12088);
nand UO_213 (O_213,N_14536,N_14363);
and UO_214 (O_214,N_13989,N_14133);
nor UO_215 (O_215,N_14052,N_14070);
nand UO_216 (O_216,N_14912,N_14893);
nor UO_217 (O_217,N_14178,N_13256);
or UO_218 (O_218,N_14960,N_13472);
nor UO_219 (O_219,N_14074,N_14646);
nand UO_220 (O_220,N_14729,N_13048);
and UO_221 (O_221,N_12770,N_13270);
and UO_222 (O_222,N_13095,N_12844);
and UO_223 (O_223,N_12287,N_12439);
nand UO_224 (O_224,N_14043,N_12669);
nor UO_225 (O_225,N_12783,N_12951);
xnor UO_226 (O_226,N_13177,N_12521);
xor UO_227 (O_227,N_12254,N_14387);
nand UO_228 (O_228,N_14005,N_13380);
and UO_229 (O_229,N_12619,N_12057);
nand UO_230 (O_230,N_14938,N_13268);
nand UO_231 (O_231,N_14189,N_13681);
or UO_232 (O_232,N_13150,N_13019);
nor UO_233 (O_233,N_14194,N_14080);
and UO_234 (O_234,N_12015,N_14439);
and UO_235 (O_235,N_12907,N_12863);
nand UO_236 (O_236,N_13888,N_14130);
nor UO_237 (O_237,N_14242,N_12795);
nand UO_238 (O_238,N_14155,N_13132);
or UO_239 (O_239,N_13108,N_12094);
or UO_240 (O_240,N_12957,N_13694);
nor UO_241 (O_241,N_14806,N_13398);
and UO_242 (O_242,N_13052,N_14831);
nor UO_243 (O_243,N_12375,N_14731);
nand UO_244 (O_244,N_12380,N_12160);
and UO_245 (O_245,N_14624,N_14216);
nor UO_246 (O_246,N_13406,N_12168);
or UO_247 (O_247,N_14367,N_12199);
nor UO_248 (O_248,N_12058,N_13771);
nor UO_249 (O_249,N_12197,N_13381);
nor UO_250 (O_250,N_13305,N_13885);
nand UO_251 (O_251,N_12318,N_13255);
and UO_252 (O_252,N_13934,N_14449);
nand UO_253 (O_253,N_12895,N_14122);
xnor UO_254 (O_254,N_14248,N_13242);
xor UO_255 (O_255,N_14900,N_13845);
or UO_256 (O_256,N_14090,N_12110);
nor UO_257 (O_257,N_14686,N_13946);
and UO_258 (O_258,N_12584,N_12503);
or UO_259 (O_259,N_13803,N_12260);
nand UO_260 (O_260,N_13424,N_14395);
nand UO_261 (O_261,N_13648,N_12291);
or UO_262 (O_262,N_12048,N_14677);
nor UO_263 (O_263,N_14997,N_12320);
and UO_264 (O_264,N_13802,N_13702);
or UO_265 (O_265,N_14980,N_13447);
nor UO_266 (O_266,N_13601,N_13068);
nor UO_267 (O_267,N_13768,N_14490);
xnor UO_268 (O_268,N_13979,N_12743);
nand UO_269 (O_269,N_14410,N_13365);
and UO_270 (O_270,N_12793,N_14724);
nand UO_271 (O_271,N_13055,N_13873);
and UO_272 (O_272,N_13556,N_14239);
nand UO_273 (O_273,N_14591,N_14530);
nand UO_274 (O_274,N_12596,N_13435);
or UO_275 (O_275,N_14810,N_14626);
nor UO_276 (O_276,N_12520,N_13489);
nor UO_277 (O_277,N_13825,N_13992);
and UO_278 (O_278,N_12161,N_13417);
nand UO_279 (O_279,N_13409,N_14408);
nor UO_280 (O_280,N_12187,N_13228);
nor UO_281 (O_281,N_13811,N_13883);
nor UO_282 (O_282,N_12272,N_13443);
or UO_283 (O_283,N_14503,N_13520);
or UO_284 (O_284,N_12631,N_12182);
and UO_285 (O_285,N_14637,N_13546);
or UO_286 (O_286,N_13033,N_12344);
and UO_287 (O_287,N_13414,N_13954);
nor UO_288 (O_288,N_14968,N_14629);
nand UO_289 (O_289,N_14622,N_14079);
nor UO_290 (O_290,N_13844,N_12665);
nor UO_291 (O_291,N_12990,N_13862);
nand UO_292 (O_292,N_12902,N_12513);
nor UO_293 (O_293,N_13085,N_13133);
and UO_294 (O_294,N_12995,N_13724);
nand UO_295 (O_295,N_12095,N_14735);
and UO_296 (O_296,N_14041,N_12529);
or UO_297 (O_297,N_14906,N_12505);
and UO_298 (O_298,N_14691,N_14642);
nand UO_299 (O_299,N_12518,N_12142);
or UO_300 (O_300,N_13708,N_13518);
or UO_301 (O_301,N_13010,N_12107);
nor UO_302 (O_302,N_14453,N_12286);
xor UO_303 (O_303,N_14709,N_14071);
or UO_304 (O_304,N_12218,N_14539);
nand UO_305 (O_305,N_14911,N_14414);
or UO_306 (O_306,N_12588,N_12134);
nand UO_307 (O_307,N_13528,N_12970);
nand UO_308 (O_308,N_14820,N_12972);
nand UO_309 (O_309,N_12459,N_14620);
nand UO_310 (O_310,N_12345,N_14720);
nor UO_311 (O_311,N_12973,N_12975);
or UO_312 (O_312,N_12814,N_12839);
nor UO_313 (O_313,N_13751,N_13799);
nor UO_314 (O_314,N_14008,N_14948);
and UO_315 (O_315,N_13656,N_14966);
nand UO_316 (O_316,N_14604,N_14160);
and UO_317 (O_317,N_13932,N_12232);
and UO_318 (O_318,N_12823,N_14744);
nand UO_319 (O_319,N_13495,N_13471);
nor UO_320 (O_320,N_12603,N_13653);
nor UO_321 (O_321,N_12750,N_13264);
nor UO_322 (O_322,N_14109,N_12502);
nor UO_323 (O_323,N_12426,N_14396);
or UO_324 (O_324,N_12415,N_12653);
or UO_325 (O_325,N_12807,N_13260);
nand UO_326 (O_326,N_12314,N_12100);
or UO_327 (O_327,N_14890,N_12075);
nor UO_328 (O_328,N_14860,N_14739);
nand UO_329 (O_329,N_14737,N_14814);
nor UO_330 (O_330,N_13814,N_13651);
nor UO_331 (O_331,N_13164,N_14701);
and UO_332 (O_332,N_12432,N_13062);
nor UO_333 (O_333,N_14865,N_12564);
xnor UO_334 (O_334,N_14094,N_14694);
or UO_335 (O_335,N_12916,N_12305);
or UO_336 (O_336,N_14513,N_13121);
or UO_337 (O_337,N_12271,N_12786);
nor UO_338 (O_338,N_14645,N_12248);
xnor UO_339 (O_339,N_12261,N_14919);
and UO_340 (O_340,N_13266,N_12659);
and UO_341 (O_341,N_13830,N_12039);
or UO_342 (O_342,N_14708,N_12856);
nand UO_343 (O_343,N_13032,N_12087);
or UO_344 (O_344,N_13124,N_13079);
nor UO_345 (O_345,N_13776,N_14434);
and UO_346 (O_346,N_12628,N_12192);
xor UO_347 (O_347,N_14098,N_13580);
or UO_348 (O_348,N_14217,N_13344);
and UO_349 (O_349,N_14941,N_13494);
nand UO_350 (O_350,N_14447,N_13265);
nand UO_351 (O_351,N_14257,N_13596);
or UO_352 (O_352,N_14533,N_12281);
and UO_353 (O_353,N_13486,N_14585);
nand UO_354 (O_354,N_13983,N_14108);
and UO_355 (O_355,N_13737,N_13842);
or UO_356 (O_356,N_12777,N_12231);
or UO_357 (O_357,N_14680,N_12558);
or UO_358 (O_358,N_14053,N_13223);
or UO_359 (O_359,N_13966,N_12397);
nor UO_360 (O_360,N_14775,N_13078);
xnor UO_361 (O_361,N_13970,N_13466);
nand UO_362 (O_362,N_13849,N_14542);
nand UO_363 (O_363,N_14357,N_14849);
nand UO_364 (O_364,N_14202,N_12998);
or UO_365 (O_365,N_13020,N_12167);
and UO_366 (O_366,N_12884,N_13877);
nand UO_367 (O_367,N_12561,N_12273);
xnor UO_368 (O_368,N_14822,N_13162);
nand UO_369 (O_369,N_12953,N_13727);
nand UO_370 (O_370,N_14466,N_14270);
nand UO_371 (O_371,N_14001,N_13968);
and UO_372 (O_372,N_14385,N_12701);
or UO_373 (O_373,N_13323,N_12677);
nor UO_374 (O_374,N_13286,N_12313);
nor UO_375 (O_375,N_13710,N_12303);
nor UO_376 (O_376,N_12848,N_12894);
and UO_377 (O_377,N_13853,N_13287);
and UO_378 (O_378,N_13393,N_13288);
xor UO_379 (O_379,N_12671,N_13131);
nor UO_380 (O_380,N_12069,N_14438);
or UO_381 (O_381,N_14950,N_14671);
or UO_382 (O_382,N_13924,N_12162);
nand UO_383 (O_383,N_14662,N_12602);
or UO_384 (O_384,N_12066,N_12141);
and UO_385 (O_385,N_14867,N_12407);
and UO_386 (O_386,N_12912,N_14825);
and UO_387 (O_387,N_14659,N_12715);
nand UO_388 (O_388,N_14521,N_13319);
nor UO_389 (O_389,N_14336,N_14835);
or UO_390 (O_390,N_13217,N_13107);
or UO_391 (O_391,N_12179,N_13375);
nor UO_392 (O_392,N_13352,N_13626);
or UO_393 (O_393,N_12202,N_14655);
nor UO_394 (O_394,N_14378,N_13531);
nand UO_395 (O_395,N_13625,N_12428);
and UO_396 (O_396,N_13993,N_14182);
or UO_397 (O_397,N_13696,N_12725);
and UO_398 (O_398,N_12976,N_13571);
or UO_399 (O_399,N_12236,N_13280);
xor UO_400 (O_400,N_13552,N_13636);
or UO_401 (O_401,N_13067,N_14335);
nor UO_402 (O_402,N_13065,N_14442);
or UO_403 (O_403,N_13516,N_14329);
or UO_404 (O_404,N_14579,N_13559);
or UO_405 (O_405,N_12361,N_14015);
nor UO_406 (O_406,N_13804,N_14895);
nor UO_407 (O_407,N_13145,N_12433);
or UO_408 (O_408,N_13558,N_13284);
and UO_409 (O_409,N_13573,N_12947);
and UO_410 (O_410,N_12478,N_14038);
or UO_411 (O_411,N_12392,N_13744);
or UO_412 (O_412,N_12140,N_13542);
and UO_413 (O_413,N_14688,N_13655);
nor UO_414 (O_414,N_14933,N_12257);
nand UO_415 (O_415,N_13433,N_12672);
xnor UO_416 (O_416,N_12221,N_14716);
or UO_417 (O_417,N_12999,N_12714);
nand UO_418 (O_418,N_13752,N_13703);
nor UO_419 (O_419,N_13774,N_12046);
nand UO_420 (O_420,N_14995,N_13762);
nand UO_421 (O_421,N_13974,N_12800);
nand UO_422 (O_422,N_13377,N_12551);
or UO_423 (O_423,N_14212,N_13667);
nand UO_424 (O_424,N_14759,N_12533);
and UO_425 (O_425,N_12532,N_12093);
or UO_426 (O_426,N_14755,N_13196);
and UO_427 (O_427,N_13731,N_12805);
nor UO_428 (O_428,N_14484,N_13676);
and UO_429 (O_429,N_13767,N_13191);
or UO_430 (O_430,N_14237,N_13828);
and UO_431 (O_431,N_14954,N_12113);
and UO_432 (O_432,N_14366,N_14280);
nand UO_433 (O_433,N_13024,N_14355);
nor UO_434 (O_434,N_13813,N_12842);
nand UO_435 (O_435,N_13796,N_12919);
or UO_436 (O_436,N_14730,N_12983);
and UO_437 (O_437,N_14942,N_12304);
or UO_438 (O_438,N_14748,N_12920);
nand UO_439 (O_439,N_12709,N_12249);
nor UO_440 (O_440,N_12451,N_14113);
nor UO_441 (O_441,N_14561,N_14389);
and UO_442 (O_442,N_14170,N_14088);
and UO_443 (O_443,N_13790,N_13519);
nand UO_444 (O_444,N_14499,N_13545);
nor UO_445 (O_445,N_14450,N_13056);
nor UO_446 (O_446,N_12540,N_14647);
or UO_447 (O_447,N_14146,N_14083);
nand UO_448 (O_448,N_13647,N_13997);
or UO_449 (O_449,N_13644,N_13854);
nand UO_450 (O_450,N_14423,N_14419);
or UO_451 (O_451,N_13541,N_14296);
or UO_452 (O_452,N_14322,N_14411);
nor UO_453 (O_453,N_14921,N_12467);
or UO_454 (O_454,N_13185,N_14627);
nand UO_455 (O_455,N_12243,N_14243);
or UO_456 (O_456,N_12053,N_13392);
nand UO_457 (O_457,N_14702,N_13939);
and UO_458 (O_458,N_13045,N_14489);
or UO_459 (O_459,N_12803,N_14594);
nand UO_460 (O_460,N_14304,N_14293);
nand UO_461 (O_461,N_13635,N_14300);
nand UO_462 (O_462,N_14504,N_13262);
or UO_463 (O_463,N_13453,N_14836);
and UO_464 (O_464,N_12099,N_14523);
nand UO_465 (O_465,N_14751,N_14733);
nand UO_466 (O_466,N_14699,N_12012);
nor UO_467 (O_467,N_12581,N_13904);
nor UO_468 (O_468,N_12610,N_13682);
nor UO_469 (O_469,N_13687,N_14535);
or UO_470 (O_470,N_14711,N_14087);
or UO_471 (O_471,N_13415,N_12330);
or UO_472 (O_472,N_14391,N_12600);
or UO_473 (O_473,N_13446,N_14928);
nand UO_474 (O_474,N_14455,N_13547);
nand UO_475 (O_475,N_13201,N_12876);
nand UO_476 (O_476,N_14478,N_14840);
and UO_477 (O_477,N_14788,N_13619);
or UO_478 (O_478,N_12758,N_13695);
and UO_479 (O_479,N_14982,N_14075);
or UO_480 (O_480,N_14294,N_13422);
nand UO_481 (O_481,N_13778,N_14628);
nand UO_482 (O_482,N_13492,N_14589);
nand UO_483 (O_483,N_13354,N_12752);
nand UO_484 (O_484,N_13590,N_13602);
and UO_485 (O_485,N_13697,N_14153);
nor UO_486 (O_486,N_12930,N_13723);
nand UO_487 (O_487,N_12865,N_14486);
nor UO_488 (O_488,N_12080,N_13662);
and UO_489 (O_489,N_14546,N_13208);
nand UO_490 (O_490,N_14876,N_14754);
and UO_491 (O_491,N_13935,N_12157);
and UO_492 (O_492,N_14977,N_14614);
nor UO_493 (O_493,N_12952,N_13449);
and UO_494 (O_494,N_13299,N_14152);
nand UO_495 (O_495,N_12546,N_14603);
or UO_496 (O_496,N_12601,N_12476);
or UO_497 (O_497,N_13335,N_12228);
or UO_498 (O_498,N_12534,N_12574);
or UO_499 (O_499,N_13328,N_13454);
nand UO_500 (O_500,N_12590,N_13491);
nor UO_501 (O_501,N_12309,N_12728);
nor UO_502 (O_502,N_13706,N_13499);
nor UO_503 (O_503,N_14925,N_13421);
nor UO_504 (O_504,N_12794,N_12034);
or UO_505 (O_505,N_13493,N_14563);
nand UO_506 (O_506,N_13660,N_12371);
and UO_507 (O_507,N_12096,N_13452);
or UO_508 (O_508,N_13218,N_14145);
nor UO_509 (O_509,N_12689,N_13787);
nor UO_510 (O_510,N_12944,N_14303);
nand UO_511 (O_511,N_13574,N_12641);
or UO_512 (O_512,N_12190,N_14692);
or UO_513 (O_513,N_13324,N_14610);
or UO_514 (O_514,N_12116,N_13609);
or UO_515 (O_515,N_14953,N_13533);
nand UO_516 (O_516,N_13404,N_14012);
nand UO_517 (O_517,N_13841,N_14310);
and UO_518 (O_518,N_14208,N_14299);
nor UO_519 (O_519,N_12465,N_14698);
or UO_520 (O_520,N_12024,N_12866);
or UO_521 (O_521,N_13374,N_12901);
and UO_522 (O_522,N_14675,N_14889);
nor UO_523 (O_523,N_14937,N_14861);
nor UO_524 (O_524,N_13327,N_14791);
nor UO_525 (O_525,N_13899,N_12608);
nand UO_526 (O_526,N_13550,N_13961);
and UO_527 (O_527,N_12772,N_12516);
or UO_528 (O_528,N_12340,N_14007);
or UO_529 (O_529,N_13929,N_13505);
nand UO_530 (O_530,N_12489,N_14753);
nor UO_531 (O_531,N_13669,N_12222);
or UO_532 (O_532,N_14863,N_13388);
and UO_533 (O_533,N_12819,N_13940);
or UO_534 (O_534,N_13895,N_12736);
nor UO_535 (O_535,N_12797,N_12755);
xor UO_536 (O_536,N_14421,N_12023);
and UO_537 (O_537,N_14660,N_14967);
nor UO_538 (O_538,N_13522,N_12060);
or UO_539 (O_539,N_12784,N_12528);
nand UO_540 (O_540,N_13535,N_12382);
and UO_541 (O_541,N_12374,N_12373);
or UO_542 (O_542,N_14039,N_12403);
or UO_543 (O_543,N_12059,N_12545);
or UO_544 (O_544,N_14666,N_13473);
and UO_545 (O_545,N_14431,N_14118);
or UO_546 (O_546,N_12473,N_12022);
nand UO_547 (O_547,N_12217,N_14634);
or UO_548 (O_548,N_14773,N_12790);
or UO_549 (O_549,N_12992,N_12542);
and UO_550 (O_550,N_13168,N_14529);
or UO_551 (O_551,N_14502,N_14550);
and UO_552 (O_552,N_14882,N_13353);
and UO_553 (O_553,N_14342,N_13100);
and UO_554 (O_554,N_14915,N_12032);
nand UO_555 (O_555,N_14598,N_14676);
or UO_556 (O_556,N_14227,N_12560);
nor UO_557 (O_557,N_13021,N_12483);
and UO_558 (O_558,N_14444,N_13532);
nor UO_559 (O_559,N_13772,N_14615);
nor UO_560 (O_560,N_13089,N_13824);
or UO_561 (O_561,N_13362,N_13995);
nor UO_562 (O_562,N_14016,N_13029);
nor UO_563 (O_563,N_14727,N_13140);
and UO_564 (O_564,N_13151,N_14538);
and UO_565 (O_565,N_12054,N_12977);
xor UO_566 (O_566,N_12063,N_13677);
and UO_567 (O_567,N_12386,N_14549);
and UO_568 (O_568,N_12180,N_13115);
nor UO_569 (O_569,N_12047,N_14636);
nor UO_570 (O_570,N_14644,N_14940);
nand UO_571 (O_571,N_13705,N_14418);
and UO_572 (O_572,N_13649,N_12724);
nor UO_573 (O_573,N_14888,N_14957);
and UO_574 (O_574,N_12555,N_14635);
or UO_575 (O_575,N_14761,N_14246);
or UO_576 (O_576,N_13382,N_14390);
and UO_577 (O_577,N_12336,N_14456);
nor UO_578 (O_578,N_14213,N_14459);
nor UO_579 (O_579,N_13500,N_13160);
xnor UO_580 (O_580,N_13576,N_12133);
and UO_581 (O_581,N_14171,N_13186);
and UO_582 (O_582,N_12592,N_14126);
and UO_583 (O_583,N_12710,N_13322);
or UO_584 (O_584,N_13138,N_14846);
nor UO_585 (O_585,N_13239,N_14873);
and UO_586 (O_586,N_13172,N_13183);
nor UO_587 (O_587,N_12247,N_12135);
or UO_588 (O_588,N_12074,N_12723);
or UO_589 (O_589,N_12508,N_12276);
or UO_590 (O_590,N_12886,N_13765);
and UO_591 (O_591,N_13870,N_13850);
and UO_592 (O_592,N_13631,N_14316);
and UO_593 (O_593,N_13606,N_12837);
nand UO_594 (O_594,N_14104,N_14738);
nand UO_595 (O_595,N_12639,N_13865);
nand UO_596 (O_596,N_13345,N_13614);
and UO_597 (O_597,N_13878,N_13698);
nor UO_598 (O_598,N_14125,N_12933);
nand UO_599 (O_599,N_13782,N_13060);
nor UO_600 (O_600,N_12647,N_14930);
nand UO_601 (O_601,N_12836,N_13818);
nand UO_602 (O_602,N_12688,N_13564);
nand UO_603 (O_603,N_12274,N_14451);
nand UO_604 (O_604,N_12177,N_12109);
or UO_605 (O_605,N_12242,N_13901);
nand UO_606 (O_606,N_12840,N_13144);
and UO_607 (O_607,N_13061,N_12613);
or UO_608 (O_608,N_13971,N_13405);
and UO_609 (O_609,N_12499,N_14446);
and UO_610 (O_610,N_13837,N_13189);
nand UO_611 (O_611,N_13175,N_12350);
and UO_612 (O_612,N_12815,N_14764);
xor UO_613 (O_613,N_12071,N_12717);
nand UO_614 (O_614,N_14050,N_14884);
nor UO_615 (O_615,N_13700,N_14872);
and UO_616 (O_616,N_12464,N_13567);
or UO_617 (O_617,N_13387,N_14422);
nor UO_618 (O_618,N_12410,N_13973);
or UO_619 (O_619,N_14777,N_14205);
and UO_620 (O_620,N_13611,N_12897);
and UO_621 (O_621,N_12233,N_12768);
and UO_622 (O_622,N_14430,N_13722);
and UO_623 (O_623,N_13936,N_14689);
nor UO_624 (O_624,N_13957,N_14282);
or UO_625 (O_625,N_13922,N_14165);
nand UO_626 (O_626,N_12213,N_14225);
or UO_627 (O_627,N_12241,N_12942);
nand UO_628 (O_628,N_12387,N_14261);
and UO_629 (O_629,N_12016,N_13586);
nor UO_630 (O_630,N_14106,N_14481);
and UO_631 (O_631,N_12754,N_13972);
or UO_632 (O_632,N_12185,N_12918);
and UO_633 (O_633,N_13712,N_12929);
nor UO_634 (O_634,N_14630,N_14406);
nor UO_635 (O_635,N_14085,N_13836);
nand UO_636 (O_636,N_12801,N_12905);
and UO_637 (O_637,N_12475,N_12870);
nor UO_638 (O_638,N_13301,N_14575);
or UO_639 (O_639,N_13594,N_12861);
and UO_640 (O_640,N_14657,N_13054);
nand UO_641 (O_641,N_12675,N_14344);
nand UO_642 (O_642,N_12346,N_14621);
or UO_643 (O_643,N_13827,N_14670);
nand UO_644 (O_644,N_12899,N_14990);
and UO_645 (O_645,N_14034,N_12938);
nand UO_646 (O_646,N_13640,N_14826);
and UO_647 (O_647,N_13234,N_12441);
nor UO_648 (O_648,N_14866,N_14308);
or UO_649 (O_649,N_13254,N_14307);
or UO_650 (O_650,N_13763,N_12519);
and UO_651 (O_651,N_14705,N_13190);
or UO_652 (O_652,N_14376,N_12994);
and UO_653 (O_653,N_13610,N_12940);
and UO_654 (O_654,N_14844,N_12234);
or UO_655 (O_655,N_14023,N_13378);
nand UO_656 (O_656,N_14428,N_12949);
and UO_657 (O_657,N_12525,N_12151);
xnor UO_658 (O_658,N_12854,N_14054);
or UO_659 (O_659,N_14746,N_12252);
nand UO_660 (O_660,N_14192,N_12120);
or UO_661 (O_661,N_14618,N_14259);
and UO_662 (O_662,N_13279,N_12114);
nand UO_663 (O_663,N_14180,N_14762);
nand UO_664 (O_664,N_12851,N_12575);
and UO_665 (O_665,N_12541,N_12991);
nor UO_666 (O_666,N_12130,N_12436);
and UO_667 (O_667,N_13738,N_13137);
nand UO_668 (O_668,N_13231,N_12487);
or UO_669 (O_669,N_14816,N_13087);
or UO_670 (O_670,N_13599,N_13037);
nand UO_671 (O_671,N_14465,N_14173);
and UO_672 (O_672,N_14672,N_12118);
nand UO_673 (O_673,N_13074,N_13198);
nand UO_674 (O_674,N_13663,N_13187);
and UO_675 (O_675,N_12697,N_13202);
and UO_676 (O_676,N_14934,N_14115);
nand UO_677 (O_677,N_13831,N_13418);
nor UO_678 (O_678,N_12020,N_12398);
nand UO_679 (O_679,N_12890,N_12316);
nand UO_680 (O_680,N_14283,N_14528);
and UO_681 (O_681,N_12853,N_12835);
nor UO_682 (O_682,N_13537,N_12948);
nor UO_683 (O_683,N_12219,N_12357);
and UO_684 (O_684,N_12722,N_12457);
nor UO_685 (O_685,N_12985,N_14559);
or UO_686 (O_686,N_12106,N_14883);
or UO_687 (O_687,N_12402,N_14042);
nand UO_688 (O_688,N_13379,N_13766);
or UO_689 (O_689,N_12137,N_14274);
nor UO_690 (O_690,N_12552,N_14218);
or UO_691 (O_691,N_14061,N_14330);
and UO_692 (O_692,N_12055,N_12364);
or UO_693 (O_693,N_12500,N_12068);
or UO_694 (O_694,N_13097,N_14245);
or UO_695 (O_695,N_13838,N_14784);
xor UO_696 (O_696,N_12898,N_12474);
and UO_697 (O_697,N_13867,N_14332);
and UO_698 (O_698,N_13953,N_14112);
nor UO_699 (O_699,N_12210,N_14369);
nand UO_700 (O_700,N_12253,N_14590);
and UO_701 (O_701,N_12523,N_12810);
and UO_702 (O_702,N_14829,N_12081);
nand UO_703 (O_703,N_12746,N_13366);
nand UO_704 (O_704,N_13812,N_13428);
nor UO_705 (O_705,N_14947,N_12621);
and UO_706 (O_706,N_14819,N_13745);
nand UO_707 (O_707,N_13258,N_12900);
nand UO_708 (O_708,N_12341,N_13568);
nor UO_709 (O_709,N_14808,N_12181);
nand UO_710 (O_710,N_14476,N_13617);
and UO_711 (O_711,N_14157,N_13321);
or UO_712 (O_712,N_14062,N_12227);
and UO_713 (O_713,N_12315,N_12981);
xor UO_714 (O_714,N_13081,N_14507);
or UO_715 (O_715,N_12526,N_12595);
and UO_716 (O_716,N_12765,N_13013);
nor UO_717 (O_717,N_12565,N_13049);
or UO_718 (O_718,N_14743,N_12466);
and UO_719 (O_719,N_12824,N_13192);
nor UO_720 (O_720,N_12582,N_12913);
or UO_721 (O_721,N_13718,N_12240);
nand UO_722 (O_722,N_12424,N_12143);
nor UO_723 (O_723,N_13444,N_13882);
and UO_724 (O_724,N_14996,N_13680);
nor UO_725 (O_725,N_13350,N_13785);
xnor UO_726 (O_726,N_13176,N_14845);
and UO_727 (O_727,N_12443,N_13605);
and UO_728 (O_728,N_14392,N_13978);
nand UO_729 (O_729,N_12650,N_12915);
and UO_730 (O_730,N_13034,N_14552);
and UO_731 (O_731,N_14760,N_14817);
nor UO_732 (O_732,N_13607,N_12351);
and UO_733 (O_733,N_13503,N_13272);
and UO_734 (O_734,N_13943,N_12634);
nor UO_735 (O_735,N_14172,N_13478);
and UO_736 (O_736,N_13009,N_13534);
and UO_737 (O_737,N_13497,N_12442);
or UO_738 (O_738,N_14868,N_14284);
nor UO_739 (O_739,N_14309,N_13282);
and UO_740 (O_740,N_14898,N_14963);
nor UO_741 (O_741,N_12329,N_13240);
nor UO_742 (O_742,N_12557,N_13117);
and UO_743 (O_743,N_14482,N_12391);
nand UO_744 (O_744,N_13504,N_13487);
or UO_745 (O_745,N_12036,N_12084);
and UO_746 (O_746,N_13360,N_13174);
and UO_747 (O_747,N_12667,N_14656);
nor UO_748 (O_748,N_13143,N_12389);
and UO_749 (O_749,N_14164,N_12616);
nor UO_750 (O_750,N_14314,N_13181);
xor UO_751 (O_751,N_12492,N_12406);
nor UO_752 (O_752,N_14994,N_13965);
nor UO_753 (O_753,N_12515,N_13050);
nand UO_754 (O_754,N_14479,N_14457);
nor UO_755 (O_755,N_13578,N_13469);
nand UO_756 (O_756,N_14658,N_12904);
and UO_757 (O_757,N_14541,N_13514);
or UO_758 (O_758,N_14811,N_13237);
or UO_759 (O_759,N_14292,N_13209);
xnor UO_760 (O_760,N_12238,N_14973);
nand UO_761 (O_761,N_12097,N_13956);
nand UO_762 (O_762,N_13101,N_13194);
nand UO_763 (O_763,N_12119,N_13304);
xor UO_764 (O_764,N_12308,N_13800);
nor UO_765 (O_765,N_13329,N_14103);
or UO_766 (O_766,N_12527,N_13507);
and UO_767 (O_767,N_12906,N_13688);
nand UO_768 (O_768,N_14100,N_13484);
and UO_769 (O_769,N_13886,N_14983);
nor UO_770 (O_770,N_14077,N_12400);
or UO_771 (O_771,N_12775,N_13898);
nor UO_772 (O_772,N_12307,N_14198);
and UO_773 (O_773,N_12988,N_14250);
nand UO_774 (O_774,N_12296,N_12360);
nand UO_775 (O_775,N_12914,N_12355);
xnor UO_776 (O_776,N_12969,N_13438);
and UO_777 (O_777,N_12352,N_14853);
or UO_778 (O_778,N_14483,N_12323);
or UO_779 (O_779,N_13432,N_14841);
and UO_780 (O_780,N_14517,N_14169);
or UO_781 (O_781,N_12372,N_14272);
nor UO_782 (O_782,N_13252,N_14548);
nor UO_783 (O_783,N_12239,N_14668);
nor UO_784 (O_784,N_14852,N_12627);
or UO_785 (O_785,N_13047,N_14818);
nand UO_786 (O_786,N_12117,N_14388);
or UO_787 (O_787,N_12481,N_13863);
nand UO_788 (O_788,N_12747,N_12766);
or UO_789 (O_789,N_14804,N_13950);
or UO_790 (O_790,N_14886,N_13843);
nor UO_791 (O_791,N_12668,N_13333);
nand UO_792 (O_792,N_14286,N_13579);
nand UO_793 (O_793,N_14570,N_13391);
nand UO_794 (O_794,N_13900,N_14512);
nand UO_795 (O_795,N_12311,N_13051);
nor UO_796 (O_796,N_14581,N_12855);
nand UO_797 (O_797,N_12462,N_12295);
or UO_798 (O_798,N_12939,N_14400);
nor UO_799 (O_799,N_14031,N_14273);
or UO_800 (O_800,N_14350,N_13216);
xor UO_801 (O_801,N_12347,N_14420);
nor UO_802 (O_802,N_13918,N_14000);
nor UO_803 (O_803,N_13769,N_14537);
and UO_804 (O_804,N_13801,N_13999);
nand UO_805 (O_805,N_13159,N_12818);
or UO_806 (O_806,N_14752,N_13788);
or UO_807 (O_807,N_14837,N_13458);
and UO_808 (O_808,N_13521,N_14800);
nor UO_809 (O_809,N_13630,N_12365);
nor UO_810 (O_810,N_13793,N_13385);
or UO_811 (O_811,N_14167,N_12440);
or UO_812 (O_812,N_13633,N_14742);
and UO_813 (O_813,N_13310,N_14128);
or UO_814 (O_814,N_12756,N_13919);
or UO_815 (O_815,N_12414,N_12605);
or UO_816 (O_816,N_12954,N_14824);
or UO_817 (O_817,N_14830,N_12152);
and UO_818 (O_818,N_14301,N_12597);
nor UO_819 (O_819,N_12599,N_14547);
or UO_820 (O_820,N_12536,N_13338);
or UO_821 (O_821,N_14206,N_12158);
nand UO_822 (O_822,N_12251,N_14064);
or UO_823 (O_823,N_12744,N_14252);
and UO_824 (O_824,N_12809,N_13431);
or UO_825 (O_825,N_12778,N_13548);
nor UO_826 (O_826,N_12270,N_13118);
nor UO_827 (O_827,N_12690,N_14196);
nor UO_828 (O_828,N_13470,N_12868);
or UO_829 (O_829,N_14340,N_13523);
or UO_830 (O_830,N_12028,N_14177);
nor UO_831 (O_831,N_13410,N_14556);
and UO_832 (O_832,N_13815,N_12511);
or UO_833 (O_833,N_13423,N_14203);
nor UO_834 (O_834,N_14055,N_12706);
and UO_835 (O_835,N_13808,N_14958);
nor UO_836 (O_836,N_13184,N_13784);
or UO_837 (O_837,N_13581,N_12891);
and UO_838 (O_838,N_12550,N_14417);
nor UO_839 (O_839,N_14238,N_13026);
or UO_840 (O_840,N_13179,N_14780);
or UO_841 (O_841,N_13149,N_14162);
nand UO_842 (O_842,N_14663,N_14432);
and UO_843 (O_843,N_12166,N_12338);
nor UO_844 (O_844,N_13756,N_14679);
and UO_845 (O_845,N_13639,N_13170);
nand UO_846 (O_846,N_14035,N_12965);
nor UO_847 (O_847,N_13915,N_12448);
or UO_848 (O_848,N_13082,N_14989);
and UO_849 (O_849,N_12052,N_13587);
and UO_850 (O_850,N_14516,N_12896);
or UO_851 (O_851,N_14929,N_12417);
nor UO_852 (O_852,N_13583,N_12789);
and UO_853 (O_853,N_12339,N_14955);
nand UO_854 (O_854,N_14260,N_13730);
nand UO_855 (O_855,N_13560,N_14003);
nand UO_856 (O_856,N_12121,N_12820);
and UO_857 (O_857,N_13871,N_14899);
nor UO_858 (O_858,N_12479,N_12009);
nor UO_859 (O_859,N_12211,N_13315);
nand UO_860 (O_860,N_12277,N_14892);
nand UO_861 (O_861,N_14030,N_14916);
and UO_862 (O_862,N_12774,N_12193);
and UO_863 (O_863,N_12716,N_14573);
nor UO_864 (O_864,N_12859,N_12284);
and UO_865 (O_865,N_12324,N_13401);
and UO_866 (O_866,N_13920,N_12751);
xor UO_867 (O_867,N_13227,N_12691);
and UO_868 (O_868,N_12494,N_14343);
and UO_869 (O_869,N_14554,N_14137);
nand UO_870 (O_870,N_12229,N_14974);
and UO_871 (O_871,N_13530,N_12704);
or UO_872 (O_872,N_12937,N_14117);
nand UO_873 (O_873,N_13749,N_12945);
nor UO_874 (O_874,N_13090,N_12681);
nand UO_875 (O_875,N_13894,N_13403);
and UO_876 (O_876,N_12175,N_14187);
xor UO_877 (O_877,N_12924,N_13511);
nor UO_878 (O_878,N_12220,N_14135);
or UO_879 (O_879,N_13364,N_13621);
nor UO_880 (O_880,N_14943,N_12530);
nand UO_881 (O_881,N_14374,N_12148);
nand UO_882 (O_882,N_12547,N_13347);
and UO_883 (O_883,N_14120,N_13099);
nor UO_884 (O_884,N_13269,N_13949);
nand UO_885 (O_885,N_14649,N_13980);
nand UO_886 (O_886,N_13283,N_13468);
nand UO_887 (O_887,N_12833,N_12258);
nor UO_888 (O_888,N_12178,N_13002);
and UO_889 (O_889,N_13128,N_13986);
nor UO_890 (O_890,N_12713,N_12005);
or UO_891 (O_891,N_13721,N_14908);
xnor UO_892 (O_892,N_13941,N_12968);
nor UO_893 (O_893,N_12204,N_12153);
or UO_894 (O_894,N_14163,N_12779);
nand UO_895 (O_895,N_13316,N_13719);
nand UO_896 (O_896,N_12570,N_13474);
or UO_897 (O_897,N_14063,N_12684);
nor UO_898 (O_898,N_14643,N_14089);
nor UO_899 (O_899,N_14065,N_12001);
nand UO_900 (O_900,N_13584,N_13407);
or UO_901 (O_901,N_12950,N_13238);
nand UO_902 (O_902,N_14924,N_13858);
and UO_903 (O_903,N_14723,N_12266);
nand UO_904 (O_904,N_14652,N_13806);
nor UO_905 (O_905,N_12963,N_13916);
or UO_906 (O_906,N_13249,N_14641);
or UO_907 (O_907,N_14611,N_12369);
nand UO_908 (O_908,N_13674,N_14792);
nand UO_909 (O_909,N_12090,N_13797);
and UO_910 (O_910,N_14904,N_12275);
and UO_911 (O_911,N_12802,N_14722);
nand UO_912 (O_912,N_14697,N_13437);
nand UO_913 (O_913,N_13028,N_12348);
nand UO_914 (O_914,N_14095,N_13147);
nand UO_915 (O_915,N_14956,N_13308);
nand UO_916 (O_916,N_14175,N_13829);
and UO_917 (O_917,N_14338,N_12593);
nor UO_918 (O_918,N_13664,N_12556);
and UO_919 (O_919,N_12332,N_13230);
or UO_920 (O_920,N_14263,N_13346);
nand UO_921 (O_921,N_14596,N_14813);
nand UO_922 (O_922,N_14362,N_13921);
or UO_923 (O_923,N_12987,N_14076);
nor UO_924 (O_924,N_14576,N_14285);
or UO_925 (O_925,N_14946,N_14448);
nor UO_926 (O_926,N_12828,N_13058);
and UO_927 (O_927,N_13952,N_12812);
or UO_928 (O_928,N_13538,N_14901);
and UO_929 (O_929,N_12246,N_12935);
and UO_930 (O_930,N_14025,N_12214);
nor UO_931 (O_931,N_12051,N_13597);
and UO_932 (O_932,N_13761,N_12554);
or UO_933 (O_933,N_14567,N_13294);
or UO_934 (O_934,N_12244,N_12325);
xnor UO_935 (O_935,N_12040,N_12869);
and UO_936 (O_936,N_12298,N_13349);
xor UO_937 (O_937,N_12205,N_12883);
or UO_938 (O_938,N_12504,N_14673);
and UO_939 (O_939,N_13967,N_12437);
xor UO_940 (O_940,N_12811,N_14381);
nor UO_941 (O_941,N_13396,N_13001);
or UO_942 (O_942,N_12695,N_13509);
or UO_943 (O_943,N_12056,N_13442);
nand UO_944 (O_944,N_13823,N_12576);
nand UO_945 (O_945,N_12734,N_14226);
nor UO_946 (O_946,N_13490,N_14199);
or UO_947 (O_947,N_13302,N_13259);
nor UO_948 (O_948,N_13786,N_12629);
xor UO_949 (O_949,N_14964,N_12816);
nor UO_950 (O_950,N_14487,N_13129);
nand UO_951 (O_951,N_14969,N_14373);
and UO_952 (O_952,N_12250,N_13152);
nand UO_953 (O_953,N_13890,N_14756);
nor UO_954 (O_954,N_13041,N_12917);
nor UO_955 (O_955,N_12769,N_14462);
nor UO_956 (O_956,N_13595,N_14520);
or UO_957 (O_957,N_12128,N_12656);
nand UO_958 (O_958,N_13477,N_12589);
or UO_959 (O_959,N_12882,N_14812);
and UO_960 (O_960,N_13627,N_13969);
nand UO_961 (O_961,N_14740,N_12376);
or UO_962 (O_962,N_12674,N_12922);
or UO_963 (O_963,N_13764,N_13928);
or UO_964 (O_964,N_13463,N_13296);
nand UO_965 (O_965,N_12753,N_14905);
nand UO_966 (O_966,N_12010,N_13003);
and UO_967 (O_967,N_14569,N_14732);
nand UO_968 (O_968,N_13293,N_12484);
nand UO_969 (O_969,N_13753,N_13770);
nand UO_970 (O_970,N_13593,N_14975);
or UO_971 (O_971,N_12062,N_12881);
nor UO_972 (O_972,N_13642,N_13629);
nand UO_973 (O_973,N_14255,N_12216);
or UO_974 (O_974,N_14291,N_13450);
or UO_975 (O_975,N_13572,N_14091);
or UO_976 (O_976,N_14714,N_14278);
xor UO_977 (O_977,N_12189,N_13742);
nor UO_978 (O_978,N_13339,N_13281);
nor UO_979 (O_979,N_13794,N_14713);
or UO_980 (O_980,N_14305,N_14002);
nor UO_981 (O_981,N_14082,N_13440);
or UO_982 (O_982,N_13944,N_13171);
and UO_983 (O_983,N_14333,N_12230);
or UO_984 (O_984,N_13725,N_13342);
and UO_985 (O_985,N_14220,N_12721);
nand UO_986 (O_986,N_12578,N_12262);
and UO_987 (O_987,N_13539,N_14168);
or UO_988 (O_988,N_13235,N_13134);
nand UO_989 (O_989,N_14734,N_14445);
and UO_990 (O_990,N_13008,N_14046);
nand UO_991 (O_991,N_14458,N_13158);
and UO_992 (O_992,N_14211,N_13866);
nor UO_993 (O_993,N_13337,N_14275);
nor UO_994 (O_994,N_13439,N_12718);
and UO_995 (O_995,N_12104,N_14269);
xnor UO_996 (O_996,N_13340,N_14665);
nand UO_997 (O_997,N_12200,N_12927);
or UO_998 (O_998,N_12843,N_13091);
and UO_999 (O_999,N_12477,N_14703);
nor UO_1000 (O_1000,N_12019,N_14186);
and UO_1001 (O_1001,N_14011,N_13707);
or UO_1002 (O_1002,N_13195,N_14609);
nand UO_1003 (O_1003,N_14749,N_12661);
and UO_1004 (O_1004,N_12740,N_12705);
nand UO_1005 (O_1005,N_14249,N_12003);
and UO_1006 (O_1006,N_14638,N_13991);
nand UO_1007 (O_1007,N_13136,N_12712);
nand UO_1008 (O_1008,N_12237,N_14551);
or UO_1009 (O_1009,N_13792,N_14639);
and UO_1010 (O_1010,N_12648,N_13563);
and UO_1011 (O_1011,N_13114,N_13613);
nor UO_1012 (O_1012,N_14185,N_14877);
nor UO_1013 (O_1013,N_12362,N_12925);
or UO_1014 (O_1014,N_13740,N_13104);
nand UO_1015 (O_1015,N_14081,N_13330);
or UO_1016 (O_1016,N_12150,N_13670);
nor UO_1017 (O_1017,N_12585,N_13246);
nand UO_1018 (O_1018,N_14936,N_14869);
nand UO_1019 (O_1019,N_14452,N_13750);
nor UO_1020 (O_1020,N_14067,N_12065);
nor UO_1021 (O_1021,N_12044,N_14325);
or UO_1022 (O_1022,N_12078,N_14028);
xnor UO_1023 (O_1023,N_13434,N_13297);
and UO_1024 (O_1024,N_13075,N_14068);
and UO_1025 (O_1025,N_14772,N_14597);
nand UO_1026 (O_1026,N_13427,N_12732);
and UO_1027 (O_1027,N_14009,N_12188);
or UO_1028 (O_1028,N_12698,N_14909);
and UO_1029 (O_1029,N_14803,N_13652);
nand UO_1030 (O_1030,N_14488,N_13426);
nor UO_1031 (O_1031,N_14221,N_14842);
or UO_1032 (O_1032,N_13063,N_12265);
nor UO_1033 (O_1033,N_13775,N_12821);
nand UO_1034 (O_1034,N_12401,N_12149);
nand UO_1035 (O_1035,N_13893,N_13646);
and UO_1036 (O_1036,N_14918,N_13213);
nor UO_1037 (O_1037,N_13113,N_13717);
nor UO_1038 (O_1038,N_12615,N_13678);
nor UO_1039 (O_1039,N_14998,N_12225);
or UO_1040 (O_1040,N_13743,N_12235);
xor UO_1041 (O_1041,N_13086,N_14891);
nand UO_1042 (O_1042,N_13030,N_14745);
nor UO_1043 (O_1043,N_14945,N_13331);
and UO_1044 (O_1044,N_13816,N_12031);
nor UO_1045 (O_1045,N_14839,N_12926);
and UO_1046 (O_1046,N_13693,N_14506);
or UO_1047 (O_1047,N_14833,N_13622);
xnor UO_1048 (O_1048,N_14669,N_13309);
and UO_1049 (O_1049,N_13975,N_14923);
xnor UO_1050 (O_1050,N_12567,N_12858);
or UO_1051 (O_1051,N_14870,N_14847);
and UO_1052 (O_1052,N_12507,N_14436);
nand UO_1053 (O_1053,N_14298,N_12267);
xor UO_1054 (O_1054,N_13038,N_14477);
or UO_1055 (O_1055,N_14522,N_12463);
or UO_1056 (O_1056,N_14757,N_14116);
or UO_1057 (O_1057,N_14834,N_14871);
nand UO_1058 (O_1058,N_12834,N_14324);
and UO_1059 (O_1059,N_12155,N_12125);
nand UO_1060 (O_1060,N_12144,N_13475);
nand UO_1061 (O_1061,N_12941,N_12383);
and UO_1062 (O_1062,N_14949,N_12033);
nor UO_1063 (O_1063,N_12147,N_14970);
nor UO_1064 (O_1064,N_13411,N_14147);
or UO_1065 (O_1065,N_14048,N_13998);
nor UO_1066 (O_1066,N_13985,N_13540);
and UO_1067 (O_1067,N_14571,N_13512);
nand UO_1068 (O_1068,N_14209,N_13204);
xnor UO_1069 (O_1069,N_13306,N_14463);
or UO_1070 (O_1070,N_14469,N_14364);
nand UO_1071 (O_1071,N_12739,N_13902);
and UO_1072 (O_1072,N_12719,N_14266);
xnor UO_1073 (O_1073,N_13263,N_13103);
or UO_1074 (O_1074,N_14191,N_14069);
or UO_1075 (O_1075,N_12379,N_13931);
nor UO_1076 (O_1076,N_14952,N_14566);
nand UO_1077 (O_1077,N_13420,N_12085);
or UO_1078 (O_1078,N_14606,N_13923);
nor UO_1079 (O_1079,N_12014,N_12285);
and UO_1080 (O_1080,N_13416,N_14613);
nor UO_1081 (O_1081,N_14534,N_12129);
or UO_1082 (O_1082,N_12838,N_13889);
xnor UO_1083 (O_1083,N_13247,N_13291);
or UO_1084 (O_1084,N_12405,N_13076);
or UO_1085 (O_1085,N_14508,N_14758);
nand UO_1086 (O_1086,N_12509,N_14809);
and UO_1087 (O_1087,N_14763,N_12301);
or UO_1088 (O_1088,N_13389,N_14875);
or UO_1089 (O_1089,N_12660,N_12889);
nor UO_1090 (O_1090,N_13042,N_14993);
or UO_1091 (O_1091,N_12996,N_13221);
or UO_1092 (O_1092,N_13673,N_12822);
or UO_1093 (O_1093,N_13225,N_12849);
nor UO_1094 (O_1094,N_14584,N_12632);
and UO_1095 (O_1095,N_13779,N_12798);
or UO_1096 (O_1096,N_12524,N_12377);
nor UO_1097 (O_1097,N_14631,N_13933);
or UO_1098 (O_1098,N_14593,N_13684);
or UO_1099 (O_1099,N_12328,N_14768);
nor UO_1100 (O_1100,N_13135,N_12212);
and UO_1101 (O_1101,N_14394,N_13232);
nand UO_1102 (O_1102,N_12434,N_12943);
or UO_1103 (O_1103,N_14987,N_12934);
and UO_1104 (O_1104,N_14514,N_12961);
or UO_1105 (O_1105,N_14233,N_13692);
and UO_1106 (O_1106,N_14371,N_13897);
or UO_1107 (O_1107,N_12435,N_13958);
or UO_1108 (O_1108,N_13826,N_13690);
or UO_1109 (O_1109,N_12419,N_14317);
nor UO_1110 (O_1110,N_14887,N_12782);
or UO_1111 (O_1111,N_12760,N_13073);
nor UO_1112 (O_1112,N_13112,N_12984);
and UO_1113 (O_1113,N_12030,N_12449);
and UO_1114 (O_1114,N_14999,N_12651);
or UO_1115 (O_1115,N_13361,N_14544);
or UO_1116 (O_1116,N_14959,N_13686);
nand UO_1117 (O_1117,N_12566,N_12207);
nor UO_1118 (O_1118,N_13043,N_14653);
nor UO_1119 (O_1119,N_13821,N_14241);
or UO_1120 (O_1120,N_12642,N_13963);
and UO_1121 (O_1121,N_12759,N_14927);
nor UO_1122 (O_1122,N_13508,N_13355);
or UO_1123 (O_1123,N_13122,N_14526);
and UO_1124 (O_1124,N_12335,N_13459);
nand UO_1125 (O_1125,N_13608,N_14736);
or UO_1126 (O_1126,N_13675,N_13053);
or UO_1127 (O_1127,N_14204,N_14302);
nor UO_1128 (O_1128,N_13102,N_12086);
and UO_1129 (O_1129,N_13628,N_13810);
and UO_1130 (O_1130,N_14965,N_14497);
nor UO_1131 (O_1131,N_14854,N_13116);
nand UO_1132 (O_1132,N_13292,N_13106);
and UO_1133 (O_1133,N_12845,N_13679);
or UO_1134 (O_1134,N_12911,N_12623);
and UO_1135 (O_1135,N_14565,N_12037);
or UO_1136 (O_1136,N_14049,N_12730);
nand UO_1137 (O_1137,N_12531,N_12874);
nand UO_1138 (O_1138,N_13072,N_12425);
and UO_1139 (O_1139,N_12429,N_14093);
nor UO_1140 (O_1140,N_14612,N_14767);
nand UO_1141 (O_1141,N_12622,N_14583);
nand UO_1142 (O_1142,N_12767,N_14159);
or UO_1143 (O_1143,N_14352,N_12191);
and UO_1144 (O_1144,N_13180,N_14557);
or UO_1145 (O_1145,N_12482,N_14188);
nand UO_1146 (O_1146,N_12679,N_14750);
nand UO_1147 (O_1147,N_12893,N_13369);
nand UO_1148 (O_1148,N_13278,N_14560);
nand UO_1149 (O_1149,N_14896,N_12655);
and UO_1150 (O_1150,N_14407,N_12283);
or UO_1151 (O_1151,N_12804,N_14779);
nand UO_1152 (O_1152,N_12067,N_13098);
and UO_1153 (O_1153,N_12496,N_14380);
or UO_1154 (O_1154,N_14201,N_12038);
nor UO_1155 (O_1155,N_13875,N_14119);
or UO_1156 (O_1156,N_13513,N_12611);
or UO_1157 (O_1157,N_12021,N_13817);
nand UO_1158 (O_1158,N_14413,N_13947);
nand UO_1159 (O_1159,N_14099,N_14010);
and UO_1160 (O_1160,N_13716,N_14174);
nand UO_1161 (O_1161,N_14029,N_13250);
nor UO_1162 (O_1162,N_13370,N_12577);
nand UO_1163 (O_1163,N_13964,N_12159);
and UO_1164 (O_1164,N_13059,N_14801);
or UO_1165 (O_1165,N_13517,N_12198);
nand UO_1166 (O_1166,N_14991,N_12594);
nand UO_1167 (O_1167,N_13501,N_12456);
nor UO_1168 (O_1168,N_13632,N_14802);
nand UO_1169 (O_1169,N_14683,N_12430);
and UO_1170 (O_1170,N_12692,N_12259);
nor UO_1171 (O_1171,N_13739,N_14019);
nor UO_1172 (O_1172,N_12393,N_12658);
and UO_1173 (O_1173,N_13982,N_12726);
and UO_1174 (O_1174,N_14402,N_13732);
nand UO_1175 (O_1175,N_13996,N_14926);
nand UO_1176 (O_1176,N_13371,N_14633);
nor UO_1177 (O_1177,N_14798,N_12864);
or UO_1178 (O_1178,N_14602,N_13212);
nor UO_1179 (O_1179,N_12131,N_12871);
and UO_1180 (O_1180,N_13071,N_12288);
or UO_1181 (O_1181,N_14102,N_12978);
or UO_1182 (O_1182,N_13057,N_13412);
nor UO_1183 (O_1183,N_13430,N_13303);
nor UO_1184 (O_1184,N_14111,N_13515);
and UO_1185 (O_1185,N_14518,N_12105);
and UO_1186 (O_1186,N_12438,N_14543);
or UO_1187 (O_1187,N_12422,N_13130);
and UO_1188 (O_1188,N_12607,N_14496);
nor UO_1189 (O_1189,N_14318,N_13153);
nand UO_1190 (O_1190,N_14706,N_13402);
nand UO_1191 (O_1191,N_14334,N_12354);
or UO_1192 (O_1192,N_13615,N_12703);
nand UO_1193 (O_1193,N_13988,N_12964);
xor UO_1194 (O_1194,N_13253,N_12367);
or UO_1195 (O_1195,N_13529,N_14214);
xor UO_1196 (O_1196,N_14073,N_12862);
and UO_1197 (O_1197,N_12013,N_13220);
and UO_1198 (O_1198,N_12245,N_12004);
or UO_1199 (O_1199,N_14276,N_14498);
nor UO_1200 (O_1200,N_12264,N_12654);
or UO_1201 (O_1201,N_13671,N_12549);
xnor UO_1202 (O_1202,N_12806,N_14519);
and UO_1203 (O_1203,N_14264,N_13461);
and UO_1204 (O_1204,N_13154,N_13846);
and UO_1205 (O_1205,N_13526,N_13142);
nor UO_1206 (O_1206,N_14897,N_14231);
and UO_1207 (O_1207,N_14200,N_14971);
nor UO_1208 (O_1208,N_14323,N_12359);
nor UO_1209 (O_1209,N_12170,N_13109);
nand UO_1210 (O_1210,N_12903,N_12337);
nor UO_1211 (O_1211,N_13173,N_13080);
nor UO_1212 (O_1212,N_12388,N_13163);
xnor UO_1213 (O_1213,N_14789,N_14114);
and UO_1214 (O_1214,N_12342,N_13120);
and UO_1215 (O_1215,N_12708,N_14219);
and UO_1216 (O_1216,N_12006,N_14326);
and UO_1217 (O_1217,N_13691,N_13638);
and UO_1218 (O_1218,N_13413,N_14290);
nor UO_1219 (O_1219,N_13069,N_12169);
nor UO_1220 (O_1220,N_12678,N_13200);
or UO_1221 (O_1221,N_14401,N_14425);
nand UO_1222 (O_1222,N_12472,N_13096);
nand UO_1223 (O_1223,N_14984,N_14492);
nand UO_1224 (O_1224,N_12061,N_14572);
nor UO_1225 (O_1225,N_12606,N_13588);
or UO_1226 (O_1226,N_14907,N_14013);
nor UO_1227 (O_1227,N_12640,N_13805);
and UO_1228 (O_1228,N_13464,N_13525);
or UO_1229 (O_1229,N_13661,N_14799);
and UO_1230 (O_1230,N_12470,N_14433);
nand UO_1231 (O_1231,N_14281,N_13938);
nor UO_1232 (O_1232,N_12327,N_13551);
or UO_1233 (O_1233,N_12413,N_14787);
nand UO_1234 (O_1234,N_12711,N_12201);
and UO_1235 (O_1235,N_13868,N_13683);
or UO_1236 (O_1236,N_12720,N_12645);
and UO_1237 (O_1237,N_14881,N_13612);
and UO_1238 (O_1238,N_12857,N_14765);
nand UO_1239 (O_1239,N_12649,N_13906);
nor UO_1240 (O_1240,N_12563,N_14384);
nand UO_1241 (O_1241,N_12742,N_14793);
and UO_1242 (O_1242,N_13139,N_12535);
nand UO_1243 (O_1243,N_12007,N_14510);
nand UO_1244 (O_1244,N_14393,N_13835);
nand UO_1245 (O_1245,N_12263,N_14288);
nand UO_1246 (O_1246,N_14337,N_12626);
nor UO_1247 (O_1247,N_14531,N_14769);
or UO_1248 (O_1248,N_12737,N_13962);
or UO_1249 (O_1249,N_12064,N_12512);
or UO_1250 (O_1250,N_14505,N_12174);
or UO_1251 (O_1251,N_13141,N_12982);
and UO_1252 (O_1252,N_13012,N_12310);
nand UO_1253 (O_1253,N_12612,N_14992);
nand UO_1254 (O_1254,N_13927,N_12624);
or UO_1255 (O_1255,N_12092,N_12676);
and UO_1256 (O_1256,N_13773,N_12165);
or UO_1257 (O_1257,N_12370,N_14903);
and UO_1258 (O_1258,N_14555,N_13780);
nor UO_1259 (O_1259,N_14092,N_13383);
nor UO_1260 (O_1260,N_14375,N_14821);
nor UO_1261 (O_1261,N_14696,N_12000);
nand UO_1262 (O_1262,N_14006,N_14577);
nor UO_1263 (O_1263,N_14295,N_14358);
nor UO_1264 (O_1264,N_14796,N_12618);
and UO_1265 (O_1265,N_14397,N_12967);
or UO_1266 (O_1266,N_13857,N_12831);
nor UO_1267 (O_1267,N_12872,N_14783);
nor UO_1268 (O_1268,N_14461,N_14347);
nand UO_1269 (O_1269,N_13777,N_13289);
nand UO_1270 (O_1270,N_12497,N_14527);
or UO_1271 (O_1271,N_12317,N_14398);
or UO_1272 (O_1272,N_12042,N_13036);
nor UO_1273 (O_1273,N_12488,N_12455);
xnor UO_1274 (O_1274,N_14693,N_12322);
and UO_1275 (O_1275,N_12637,N_14578);
nand UO_1276 (O_1276,N_13892,N_14047);
nor UO_1277 (O_1277,N_12145,N_14210);
or UO_1278 (O_1278,N_12223,N_12471);
and UO_1279 (O_1279,N_13376,N_14726);
nor UO_1280 (O_1280,N_12073,N_13860);
and UO_1281 (O_1281,N_12123,N_14651);
or UO_1282 (O_1282,N_14144,N_14648);
or UO_1283 (O_1283,N_13734,N_13665);
or UO_1284 (O_1284,N_12183,N_12103);
nand UO_1285 (O_1285,N_12173,N_12091);
nand UO_1286 (O_1286,N_12138,N_14253);
nand UO_1287 (O_1287,N_12333,N_13994);
nand UO_1288 (O_1288,N_13896,N_14370);
or UO_1289 (O_1289,N_14360,N_13110);
nand UO_1290 (O_1290,N_12680,N_12792);
nor UO_1291 (O_1291,N_14747,N_12748);
nand UO_1292 (O_1292,N_13758,N_14404);
nand UO_1293 (O_1293,N_14587,N_14786);
nand UO_1294 (O_1294,N_12879,N_13126);
nor UO_1295 (O_1295,N_13343,N_14474);
and UO_1296 (O_1296,N_14078,N_12686);
and UO_1297 (O_1297,N_14045,N_12139);
nor UO_1298 (O_1298,N_12098,N_13881);
xnor UO_1299 (O_1299,N_13937,N_13022);
or UO_1300 (O_1300,N_14879,N_12124);
nor UO_1301 (O_1301,N_12409,N_13326);
nor UO_1302 (O_1302,N_13589,N_13419);
nand UO_1303 (O_1303,N_14795,N_13741);
nand UO_1304 (O_1304,N_14678,N_12633);
or UO_1305 (O_1305,N_13884,N_13093);
nor UO_1306 (O_1306,N_14471,N_13569);
nand UO_1307 (O_1307,N_12620,N_14682);
nand UO_1308 (O_1308,N_14961,N_13119);
xnor UO_1309 (O_1309,N_13480,N_14564);
nor UO_1310 (O_1310,N_14262,N_12289);
xnor UO_1311 (O_1311,N_13188,N_12163);
and UO_1312 (O_1312,N_13598,N_14032);
or UO_1313 (O_1313,N_13226,N_13025);
or UO_1314 (O_1314,N_13926,N_14864);
nor UO_1315 (O_1315,N_14267,N_14348);
nand UO_1316 (O_1316,N_13248,N_12506);
nor UO_1317 (O_1317,N_12971,N_12224);
nand UO_1318 (O_1318,N_13623,N_14902);
or UO_1319 (O_1319,N_13951,N_14020);
and UO_1320 (O_1320,N_12572,N_14717);
nor UO_1321 (O_1321,N_14922,N_14158);
nor UO_1322 (O_1322,N_14136,N_13448);
nand UO_1323 (O_1323,N_14574,N_14728);
or UO_1324 (O_1324,N_14741,N_13666);
nor UO_1325 (O_1325,N_14353,N_13298);
or UO_1326 (O_1326,N_12171,N_14778);
and UO_1327 (O_1327,N_12548,N_12727);
and UO_1328 (O_1328,N_14495,N_12693);
or UO_1329 (O_1329,N_13275,N_14582);
nor UO_1330 (O_1330,N_14084,N_12368);
nand UO_1331 (O_1331,N_12018,N_13046);
xor UO_1332 (O_1332,N_12580,N_13798);
nor UO_1333 (O_1333,N_13465,N_13165);
nor UO_1334 (O_1334,N_14480,N_13257);
nand UO_1335 (O_1335,N_12186,N_13429);
nand UO_1336 (O_1336,N_14129,N_12630);
or UO_1337 (O_1337,N_12757,N_13488);
and UO_1338 (O_1338,N_13847,N_12887);
and UO_1339 (O_1339,N_12302,N_12568);
nand UO_1340 (O_1340,N_13701,N_14981);
nor UO_1341 (O_1341,N_12460,N_12764);
and UO_1342 (O_1342,N_13408,N_14372);
nand UO_1343 (O_1343,N_14138,N_14328);
or UO_1344 (O_1344,N_13105,N_13205);
nor UO_1345 (O_1345,N_12101,N_12293);
nand UO_1346 (O_1346,N_13148,N_14139);
nor UO_1347 (O_1347,N_13977,N_12928);
nor UO_1348 (O_1348,N_13482,N_14525);
and UO_1349 (O_1349,N_14379,N_14265);
and UO_1350 (O_1350,N_12735,N_14409);
and UO_1351 (O_1351,N_14383,N_14972);
nand UO_1352 (O_1352,N_12544,N_12888);
nand UO_1353 (O_1353,N_13203,N_12799);
nand UO_1354 (O_1354,N_12825,N_12738);
or UO_1355 (O_1355,N_13384,N_13167);
nand UO_1356 (O_1356,N_12111,N_14207);
and UO_1357 (O_1357,N_14141,N_14851);
nor UO_1358 (O_1358,N_12559,N_12268);
or UO_1359 (O_1359,N_13276,N_13400);
xor UO_1360 (O_1360,N_13451,N_14910);
or UO_1361 (O_1361,N_14312,N_12156);
or UO_1362 (O_1362,N_13855,N_14588);
nor UO_1363 (O_1363,N_13637,N_14986);
nor UO_1364 (O_1364,N_12282,N_12780);
and UO_1365 (O_1365,N_14036,N_12501);
or UO_1366 (O_1366,N_13243,N_12343);
and UO_1367 (O_1367,N_12733,N_14033);
nor UO_1368 (O_1368,N_12280,N_12045);
nor UO_1369 (O_1369,N_12102,N_14197);
or UO_1370 (O_1370,N_12491,N_12817);
nor UO_1371 (O_1371,N_14491,N_12662);
nor UO_1372 (O_1372,N_14354,N_12083);
nand UO_1373 (O_1373,N_12331,N_12082);
nor UO_1374 (O_1374,N_13094,N_13711);
nor UO_1375 (O_1375,N_12312,N_12421);
nor UO_1376 (O_1376,N_12132,N_13206);
and UO_1377 (O_1377,N_12657,N_12699);
xor UO_1378 (O_1378,N_14223,N_14815);
and UO_1379 (O_1379,N_14920,N_13747);
or UO_1380 (O_1380,N_12079,N_14632);
nor UO_1381 (O_1381,N_12604,N_14664);
or UO_1382 (O_1382,N_13425,N_12666);
nand UO_1383 (O_1383,N_14878,N_13832);
nand UO_1384 (O_1384,N_12663,N_13290);
nor UO_1385 (O_1385,N_12029,N_14107);
xnor UO_1386 (O_1386,N_13146,N_13462);
nand UO_1387 (O_1387,N_12931,N_13318);
nand UO_1388 (O_1388,N_12694,N_14515);
nand UO_1389 (O_1389,N_14894,N_14605);
and UO_1390 (O_1390,N_13456,N_12763);
nand UO_1391 (O_1391,N_13157,N_14193);
and UO_1392 (O_1392,N_12685,N_13909);
nor UO_1393 (O_1393,N_14667,N_12635);
nor UO_1394 (O_1394,N_13807,N_12646);
or UO_1395 (O_1395,N_14359,N_12956);
nand UO_1396 (O_1396,N_13555,N_14931);
and UO_1397 (O_1397,N_12846,N_13689);
nor UO_1398 (O_1398,N_14472,N_14850);
nor UO_1399 (O_1399,N_12334,N_12829);
and UO_1400 (O_1400,N_13736,N_12490);
or UO_1401 (O_1401,N_14443,N_14224);
and UO_1402 (O_1402,N_13357,N_12011);
nor UO_1403 (O_1403,N_14148,N_13618);
nor UO_1404 (O_1404,N_13930,N_12993);
nand UO_1405 (O_1405,N_13178,N_13948);
nand UO_1406 (O_1406,N_14951,N_13544);
or UO_1407 (O_1407,N_13023,N_13759);
nor UO_1408 (O_1408,N_13219,N_14229);
and UO_1409 (O_1409,N_12591,N_13748);
nand UO_1410 (O_1410,N_14858,N_13645);
nand UO_1411 (O_1411,N_14416,N_12771);
nand UO_1412 (O_1412,N_13713,N_13903);
or UO_1413 (O_1413,N_13457,N_14123);
nand UO_1414 (O_1414,N_12255,N_14595);
and UO_1415 (O_1415,N_14435,N_13864);
and UO_1416 (O_1416,N_12427,N_14412);
and UO_1417 (O_1417,N_14640,N_12877);
xor UO_1418 (O_1418,N_13251,N_12932);
nand UO_1419 (O_1419,N_13016,N_13485);
nand UO_1420 (O_1420,N_12962,N_12485);
nand UO_1421 (O_1421,N_12989,N_12847);
nand UO_1422 (O_1422,N_13911,N_13006);
or UO_1423 (O_1423,N_14072,N_12788);
xor UO_1424 (O_1424,N_13317,N_12420);
nor UO_1425 (O_1425,N_13856,N_13161);
and UO_1426 (O_1426,N_14327,N_14568);
nor UO_1427 (O_1427,N_14979,N_12832);
nor UO_1428 (O_1428,N_13261,N_13441);
nor UO_1429 (O_1429,N_12297,N_13368);
and UO_1430 (O_1430,N_13654,N_13641);
nand UO_1431 (O_1431,N_12321,N_12664);
or UO_1432 (O_1432,N_14236,N_14874);
nand UO_1433 (O_1433,N_13040,N_14797);
nor UO_1434 (O_1434,N_12431,N_14855);
nor UO_1435 (O_1435,N_12850,N_14346);
nor UO_1436 (O_1436,N_13549,N_14149);
and UO_1437 (O_1437,N_13757,N_13577);
or UO_1438 (O_1438,N_13363,N_14988);
and UO_1439 (O_1439,N_14654,N_14540);
and UO_1440 (O_1440,N_12910,N_13199);
nand UO_1441 (O_1441,N_14268,N_14719);
or UO_1442 (O_1442,N_14823,N_12538);
nor UO_1443 (O_1443,N_13233,N_12867);
nand UO_1444 (O_1444,N_13746,N_14124);
nand UO_1445 (O_1445,N_13570,N_12830);
or UO_1446 (O_1446,N_14022,N_12880);
or UO_1447 (O_1447,N_14277,N_12049);
and UO_1448 (O_1448,N_14827,N_12673);
nand UO_1449 (O_1449,N_14978,N_12026);
and UO_1450 (O_1450,N_12745,N_13285);
nand UO_1451 (O_1451,N_12569,N_13729);
or UO_1452 (O_1452,N_13733,N_13064);
nor UO_1453 (O_1453,N_13925,N_12670);
nand UO_1454 (O_1454,N_12875,N_13083);
and UO_1455 (O_1455,N_12290,N_14154);
nand UO_1456 (O_1456,N_14315,N_12885);
or UO_1457 (O_1457,N_12892,N_14885);
nor UO_1458 (O_1458,N_12644,N_13066);
nand UO_1459 (O_1459,N_13111,N_14862);
nor UO_1460 (O_1460,N_12294,N_13872);
nand UO_1461 (O_1461,N_13241,N_13320);
nor UO_1462 (O_1462,N_13942,N_12458);
nor UO_1463 (O_1463,N_14415,N_12683);
xnor UO_1464 (O_1464,N_12404,N_14306);
nor UO_1465 (O_1465,N_12209,N_12452);
or UO_1466 (O_1466,N_14794,N_13125);
and UO_1467 (O_1467,N_12195,N_12469);
xor UO_1468 (O_1468,N_14707,N_12226);
and UO_1469 (O_1469,N_14454,N_14356);
nor UO_1470 (O_1470,N_13839,N_14782);
nor UO_1471 (O_1471,N_12514,N_13210);
or UO_1472 (O_1472,N_12208,N_13436);
nor UO_1473 (O_1473,N_12394,N_13027);
and UO_1474 (O_1474,N_14721,N_13277);
or UO_1475 (O_1475,N_14473,N_12980);
nor UO_1476 (O_1476,N_12878,N_13000);
or UO_1477 (O_1477,N_13704,N_12279);
or UO_1478 (O_1478,N_13685,N_13229);
nor UO_1479 (O_1479,N_12041,N_13496);
nor UO_1480 (O_1480,N_14674,N_14944);
and UO_1481 (O_1481,N_13987,N_14607);
xnor UO_1482 (O_1482,N_12122,N_12696);
and UO_1483 (O_1483,N_13880,N_13455);
nor UO_1484 (O_1484,N_13070,N_13295);
nand UO_1485 (O_1485,N_14700,N_14351);
nand UO_1486 (O_1486,N_13917,N_14562);
or UO_1487 (O_1487,N_13483,N_12025);
or UO_1488 (O_1488,N_12986,N_14215);
nor UO_1489 (O_1489,N_13658,N_12539);
or UO_1490 (O_1490,N_14600,N_12076);
xnor UO_1491 (O_1491,N_14426,N_13273);
or UO_1492 (O_1492,N_13536,N_14132);
nand UO_1493 (O_1493,N_12008,N_14289);
nand UO_1494 (O_1494,N_13672,N_14195);
nand UO_1495 (O_1495,N_13912,N_14228);
or UO_1496 (O_1496,N_12319,N_12776);
nor UO_1497 (O_1497,N_12349,N_14935);
nand UO_1498 (O_1498,N_14843,N_13795);
or UO_1499 (O_1499,N_13018,N_14240);
xor UO_1500 (O_1500,N_13066,N_12117);
and UO_1501 (O_1501,N_13675,N_12657);
nor UO_1502 (O_1502,N_13196,N_13066);
and UO_1503 (O_1503,N_12524,N_14757);
or UO_1504 (O_1504,N_12774,N_14580);
nor UO_1505 (O_1505,N_14727,N_14100);
and UO_1506 (O_1506,N_13843,N_12136);
nand UO_1507 (O_1507,N_13832,N_12245);
and UO_1508 (O_1508,N_13204,N_14846);
nand UO_1509 (O_1509,N_12331,N_14827);
nor UO_1510 (O_1510,N_14016,N_12532);
or UO_1511 (O_1511,N_12946,N_14121);
and UO_1512 (O_1512,N_12874,N_12592);
xor UO_1513 (O_1513,N_13091,N_12079);
or UO_1514 (O_1514,N_12770,N_14653);
and UO_1515 (O_1515,N_14256,N_12799);
nor UO_1516 (O_1516,N_14414,N_13191);
or UO_1517 (O_1517,N_12736,N_14047);
nor UO_1518 (O_1518,N_13679,N_14314);
or UO_1519 (O_1519,N_13640,N_14346);
nor UO_1520 (O_1520,N_14162,N_14590);
or UO_1521 (O_1521,N_13871,N_12731);
nand UO_1522 (O_1522,N_14617,N_14721);
or UO_1523 (O_1523,N_13372,N_14443);
nor UO_1524 (O_1524,N_13578,N_14928);
or UO_1525 (O_1525,N_12391,N_12576);
and UO_1526 (O_1526,N_12937,N_14595);
nand UO_1527 (O_1527,N_14917,N_13532);
nor UO_1528 (O_1528,N_12120,N_14324);
or UO_1529 (O_1529,N_13741,N_12639);
or UO_1530 (O_1530,N_12993,N_12947);
xnor UO_1531 (O_1531,N_14238,N_12308);
nand UO_1532 (O_1532,N_14402,N_13886);
nor UO_1533 (O_1533,N_13497,N_14041);
nor UO_1534 (O_1534,N_12673,N_14006);
nor UO_1535 (O_1535,N_13661,N_13200);
nand UO_1536 (O_1536,N_14958,N_12435);
nor UO_1537 (O_1537,N_13013,N_12453);
or UO_1538 (O_1538,N_12275,N_12712);
xnor UO_1539 (O_1539,N_12807,N_14100);
or UO_1540 (O_1540,N_14517,N_14791);
nand UO_1541 (O_1541,N_13181,N_12725);
nor UO_1542 (O_1542,N_13380,N_13941);
nand UO_1543 (O_1543,N_13221,N_14927);
nand UO_1544 (O_1544,N_12047,N_14233);
or UO_1545 (O_1545,N_12744,N_14314);
or UO_1546 (O_1546,N_13330,N_13364);
or UO_1547 (O_1547,N_12855,N_13396);
or UO_1548 (O_1548,N_14670,N_13254);
or UO_1549 (O_1549,N_14405,N_14506);
or UO_1550 (O_1550,N_12546,N_14859);
nor UO_1551 (O_1551,N_12222,N_14056);
nand UO_1552 (O_1552,N_12531,N_14920);
or UO_1553 (O_1553,N_12005,N_13986);
nand UO_1554 (O_1554,N_12124,N_13739);
or UO_1555 (O_1555,N_12388,N_13384);
nor UO_1556 (O_1556,N_12216,N_13525);
or UO_1557 (O_1557,N_12337,N_14009);
nor UO_1558 (O_1558,N_13189,N_12237);
nor UO_1559 (O_1559,N_14461,N_12053);
nor UO_1560 (O_1560,N_12705,N_13668);
and UO_1561 (O_1561,N_12883,N_14068);
nand UO_1562 (O_1562,N_12065,N_14866);
and UO_1563 (O_1563,N_13300,N_14889);
xor UO_1564 (O_1564,N_14421,N_14435);
nor UO_1565 (O_1565,N_13107,N_14551);
or UO_1566 (O_1566,N_13245,N_14856);
nand UO_1567 (O_1567,N_14519,N_13006);
nand UO_1568 (O_1568,N_13768,N_14898);
and UO_1569 (O_1569,N_14536,N_13519);
xnor UO_1570 (O_1570,N_13598,N_14264);
nand UO_1571 (O_1571,N_12608,N_13805);
or UO_1572 (O_1572,N_12574,N_12739);
or UO_1573 (O_1573,N_12136,N_12466);
and UO_1574 (O_1574,N_12714,N_12421);
or UO_1575 (O_1575,N_13993,N_12726);
or UO_1576 (O_1576,N_14763,N_13482);
nand UO_1577 (O_1577,N_12986,N_13698);
nand UO_1578 (O_1578,N_14417,N_13330);
nand UO_1579 (O_1579,N_14444,N_14228);
or UO_1580 (O_1580,N_13229,N_14357);
nand UO_1581 (O_1581,N_14179,N_12187);
nand UO_1582 (O_1582,N_12625,N_14675);
and UO_1583 (O_1583,N_12207,N_14764);
nor UO_1584 (O_1584,N_14594,N_14235);
nor UO_1585 (O_1585,N_13060,N_13531);
and UO_1586 (O_1586,N_14200,N_13914);
nand UO_1587 (O_1587,N_13514,N_13752);
or UO_1588 (O_1588,N_13021,N_12033);
nand UO_1589 (O_1589,N_13233,N_14278);
nor UO_1590 (O_1590,N_13862,N_12528);
and UO_1591 (O_1591,N_12094,N_14590);
nor UO_1592 (O_1592,N_14070,N_14794);
nand UO_1593 (O_1593,N_13168,N_14980);
or UO_1594 (O_1594,N_13160,N_13446);
nand UO_1595 (O_1595,N_13244,N_12794);
and UO_1596 (O_1596,N_12548,N_14058);
nor UO_1597 (O_1597,N_12163,N_12446);
or UO_1598 (O_1598,N_12426,N_14713);
or UO_1599 (O_1599,N_12510,N_14150);
nand UO_1600 (O_1600,N_12799,N_13419);
nand UO_1601 (O_1601,N_13720,N_14195);
nand UO_1602 (O_1602,N_12603,N_14925);
or UO_1603 (O_1603,N_14094,N_13111);
nand UO_1604 (O_1604,N_12056,N_14672);
or UO_1605 (O_1605,N_12700,N_14166);
xnor UO_1606 (O_1606,N_12760,N_12142);
and UO_1607 (O_1607,N_14183,N_14525);
nand UO_1608 (O_1608,N_14016,N_12604);
nand UO_1609 (O_1609,N_13447,N_12756);
or UO_1610 (O_1610,N_13940,N_14962);
and UO_1611 (O_1611,N_13973,N_14936);
xor UO_1612 (O_1612,N_14910,N_12278);
nand UO_1613 (O_1613,N_14774,N_14285);
nor UO_1614 (O_1614,N_12922,N_12755);
or UO_1615 (O_1615,N_13817,N_14865);
or UO_1616 (O_1616,N_13562,N_12225);
or UO_1617 (O_1617,N_14976,N_13053);
nor UO_1618 (O_1618,N_13158,N_13363);
nand UO_1619 (O_1619,N_13327,N_13197);
and UO_1620 (O_1620,N_12378,N_12617);
nor UO_1621 (O_1621,N_14499,N_14871);
nor UO_1622 (O_1622,N_14905,N_14294);
and UO_1623 (O_1623,N_12331,N_14758);
nor UO_1624 (O_1624,N_14074,N_13733);
or UO_1625 (O_1625,N_12128,N_12721);
or UO_1626 (O_1626,N_14694,N_13844);
or UO_1627 (O_1627,N_12424,N_14544);
and UO_1628 (O_1628,N_14356,N_12294);
nor UO_1629 (O_1629,N_14243,N_13940);
and UO_1630 (O_1630,N_13543,N_13033);
and UO_1631 (O_1631,N_13766,N_14599);
nor UO_1632 (O_1632,N_13447,N_14279);
and UO_1633 (O_1633,N_14051,N_14567);
nand UO_1634 (O_1634,N_14241,N_14071);
and UO_1635 (O_1635,N_13104,N_14128);
nand UO_1636 (O_1636,N_14769,N_14912);
nor UO_1637 (O_1637,N_12443,N_13752);
and UO_1638 (O_1638,N_14824,N_14914);
nor UO_1639 (O_1639,N_12228,N_13531);
or UO_1640 (O_1640,N_14778,N_12393);
and UO_1641 (O_1641,N_12406,N_12489);
nor UO_1642 (O_1642,N_14378,N_14951);
nor UO_1643 (O_1643,N_12363,N_12236);
xnor UO_1644 (O_1644,N_13216,N_14094);
nor UO_1645 (O_1645,N_12357,N_13455);
or UO_1646 (O_1646,N_13139,N_12672);
nor UO_1647 (O_1647,N_14282,N_12915);
and UO_1648 (O_1648,N_14468,N_13579);
and UO_1649 (O_1649,N_12206,N_13041);
nand UO_1650 (O_1650,N_12433,N_13197);
xnor UO_1651 (O_1651,N_14540,N_14579);
and UO_1652 (O_1652,N_13327,N_13932);
nand UO_1653 (O_1653,N_13139,N_13257);
nor UO_1654 (O_1654,N_13302,N_13529);
nand UO_1655 (O_1655,N_13237,N_13167);
and UO_1656 (O_1656,N_13468,N_14890);
and UO_1657 (O_1657,N_13178,N_12417);
nor UO_1658 (O_1658,N_12901,N_13058);
nor UO_1659 (O_1659,N_12326,N_12136);
nand UO_1660 (O_1660,N_14153,N_12669);
and UO_1661 (O_1661,N_13089,N_13560);
and UO_1662 (O_1662,N_12498,N_12233);
or UO_1663 (O_1663,N_13472,N_12906);
and UO_1664 (O_1664,N_12832,N_13267);
or UO_1665 (O_1665,N_13606,N_13214);
nand UO_1666 (O_1666,N_13083,N_13380);
nand UO_1667 (O_1667,N_14646,N_13345);
or UO_1668 (O_1668,N_14440,N_13274);
and UO_1669 (O_1669,N_14786,N_14152);
or UO_1670 (O_1670,N_13402,N_12396);
and UO_1671 (O_1671,N_14175,N_12685);
nand UO_1672 (O_1672,N_13927,N_13505);
or UO_1673 (O_1673,N_13359,N_12606);
nand UO_1674 (O_1674,N_12293,N_12863);
nand UO_1675 (O_1675,N_14485,N_14386);
xnor UO_1676 (O_1676,N_13664,N_13433);
or UO_1677 (O_1677,N_13419,N_12443);
nor UO_1678 (O_1678,N_13890,N_13299);
and UO_1679 (O_1679,N_13073,N_14407);
or UO_1680 (O_1680,N_13213,N_13482);
nor UO_1681 (O_1681,N_14206,N_14494);
or UO_1682 (O_1682,N_12215,N_13724);
and UO_1683 (O_1683,N_13613,N_12025);
nor UO_1684 (O_1684,N_14882,N_13476);
nand UO_1685 (O_1685,N_14780,N_14144);
nor UO_1686 (O_1686,N_12585,N_13094);
nand UO_1687 (O_1687,N_13366,N_14147);
nor UO_1688 (O_1688,N_12790,N_12422);
and UO_1689 (O_1689,N_14909,N_13629);
nor UO_1690 (O_1690,N_13874,N_14990);
nor UO_1691 (O_1691,N_13080,N_13853);
or UO_1692 (O_1692,N_12571,N_12229);
nor UO_1693 (O_1693,N_12392,N_12676);
and UO_1694 (O_1694,N_14931,N_12518);
nand UO_1695 (O_1695,N_14314,N_13871);
or UO_1696 (O_1696,N_13327,N_14353);
nand UO_1697 (O_1697,N_12073,N_12139);
and UO_1698 (O_1698,N_12271,N_14949);
and UO_1699 (O_1699,N_14277,N_14252);
and UO_1700 (O_1700,N_12971,N_13598);
nor UO_1701 (O_1701,N_13024,N_12182);
and UO_1702 (O_1702,N_12161,N_14239);
xor UO_1703 (O_1703,N_12057,N_12170);
and UO_1704 (O_1704,N_12058,N_12749);
xor UO_1705 (O_1705,N_12333,N_12752);
or UO_1706 (O_1706,N_13381,N_12892);
or UO_1707 (O_1707,N_12540,N_14682);
and UO_1708 (O_1708,N_13715,N_12593);
nand UO_1709 (O_1709,N_12552,N_12736);
nand UO_1710 (O_1710,N_13265,N_12941);
or UO_1711 (O_1711,N_12151,N_12028);
and UO_1712 (O_1712,N_14635,N_13108);
and UO_1713 (O_1713,N_14280,N_12408);
nor UO_1714 (O_1714,N_13207,N_13433);
nor UO_1715 (O_1715,N_13673,N_13645);
nor UO_1716 (O_1716,N_14372,N_13807);
xor UO_1717 (O_1717,N_14573,N_12615);
and UO_1718 (O_1718,N_13968,N_12950);
nand UO_1719 (O_1719,N_12538,N_12891);
or UO_1720 (O_1720,N_13477,N_13317);
nor UO_1721 (O_1721,N_12923,N_12314);
nand UO_1722 (O_1722,N_14314,N_13162);
and UO_1723 (O_1723,N_13254,N_13262);
and UO_1724 (O_1724,N_12774,N_12054);
nor UO_1725 (O_1725,N_12544,N_12975);
or UO_1726 (O_1726,N_14487,N_12932);
or UO_1727 (O_1727,N_12325,N_14152);
nor UO_1728 (O_1728,N_14738,N_13676);
nor UO_1729 (O_1729,N_13472,N_13287);
nor UO_1730 (O_1730,N_13949,N_13320);
nor UO_1731 (O_1731,N_13347,N_14538);
nor UO_1732 (O_1732,N_12048,N_12291);
and UO_1733 (O_1733,N_14355,N_12854);
nor UO_1734 (O_1734,N_14918,N_14945);
or UO_1735 (O_1735,N_12933,N_13646);
nand UO_1736 (O_1736,N_13213,N_12915);
nor UO_1737 (O_1737,N_12752,N_12841);
nand UO_1738 (O_1738,N_14773,N_14307);
nand UO_1739 (O_1739,N_12260,N_13775);
nand UO_1740 (O_1740,N_13394,N_13912);
nor UO_1741 (O_1741,N_13650,N_12402);
nand UO_1742 (O_1742,N_13427,N_12094);
or UO_1743 (O_1743,N_12246,N_14311);
nor UO_1744 (O_1744,N_12383,N_13146);
nor UO_1745 (O_1745,N_13721,N_12921);
nand UO_1746 (O_1746,N_12012,N_12401);
and UO_1747 (O_1747,N_13568,N_14971);
or UO_1748 (O_1748,N_13154,N_12210);
or UO_1749 (O_1749,N_12671,N_12262);
nor UO_1750 (O_1750,N_12271,N_13085);
and UO_1751 (O_1751,N_12857,N_14897);
nor UO_1752 (O_1752,N_14302,N_13939);
or UO_1753 (O_1753,N_14553,N_14829);
nor UO_1754 (O_1754,N_12078,N_14070);
and UO_1755 (O_1755,N_13670,N_14428);
nand UO_1756 (O_1756,N_14824,N_14223);
nor UO_1757 (O_1757,N_12830,N_13531);
or UO_1758 (O_1758,N_14847,N_12803);
nand UO_1759 (O_1759,N_13651,N_14846);
nor UO_1760 (O_1760,N_12567,N_12739);
and UO_1761 (O_1761,N_14140,N_13414);
nand UO_1762 (O_1762,N_13089,N_14452);
or UO_1763 (O_1763,N_14024,N_12295);
and UO_1764 (O_1764,N_13844,N_13490);
nand UO_1765 (O_1765,N_12181,N_12062);
nor UO_1766 (O_1766,N_12874,N_13228);
nand UO_1767 (O_1767,N_13923,N_14977);
xnor UO_1768 (O_1768,N_14370,N_13479);
nand UO_1769 (O_1769,N_12479,N_14083);
xor UO_1770 (O_1770,N_14290,N_13136);
or UO_1771 (O_1771,N_14264,N_13940);
nand UO_1772 (O_1772,N_14330,N_12912);
and UO_1773 (O_1773,N_14994,N_12471);
nor UO_1774 (O_1774,N_13207,N_13654);
and UO_1775 (O_1775,N_12535,N_12906);
nand UO_1776 (O_1776,N_13804,N_12164);
nand UO_1777 (O_1777,N_13706,N_14394);
and UO_1778 (O_1778,N_12111,N_13559);
and UO_1779 (O_1779,N_13504,N_14943);
nor UO_1780 (O_1780,N_13118,N_14863);
nor UO_1781 (O_1781,N_13186,N_13533);
nor UO_1782 (O_1782,N_14333,N_13405);
nand UO_1783 (O_1783,N_14305,N_13729);
and UO_1784 (O_1784,N_13229,N_12190);
and UO_1785 (O_1785,N_14672,N_12928);
nor UO_1786 (O_1786,N_13306,N_13038);
and UO_1787 (O_1787,N_13301,N_13711);
xor UO_1788 (O_1788,N_12635,N_12072);
or UO_1789 (O_1789,N_13206,N_13958);
nor UO_1790 (O_1790,N_13352,N_12680);
and UO_1791 (O_1791,N_12608,N_13129);
and UO_1792 (O_1792,N_12168,N_12104);
or UO_1793 (O_1793,N_12464,N_12880);
nand UO_1794 (O_1794,N_13584,N_13286);
or UO_1795 (O_1795,N_12130,N_12808);
or UO_1796 (O_1796,N_13756,N_14159);
nor UO_1797 (O_1797,N_13282,N_13946);
and UO_1798 (O_1798,N_13877,N_14973);
or UO_1799 (O_1799,N_14903,N_12669);
or UO_1800 (O_1800,N_12074,N_12434);
and UO_1801 (O_1801,N_14142,N_13489);
nand UO_1802 (O_1802,N_12980,N_13351);
nor UO_1803 (O_1803,N_12504,N_14185);
nand UO_1804 (O_1804,N_12989,N_13061);
nor UO_1805 (O_1805,N_12654,N_13815);
or UO_1806 (O_1806,N_12087,N_14300);
and UO_1807 (O_1807,N_13546,N_13400);
nor UO_1808 (O_1808,N_13137,N_14685);
or UO_1809 (O_1809,N_12901,N_12746);
or UO_1810 (O_1810,N_14940,N_14130);
nand UO_1811 (O_1811,N_12658,N_12349);
nor UO_1812 (O_1812,N_12212,N_12226);
or UO_1813 (O_1813,N_12725,N_12560);
or UO_1814 (O_1814,N_13104,N_14176);
nor UO_1815 (O_1815,N_14860,N_13177);
or UO_1816 (O_1816,N_12017,N_14793);
and UO_1817 (O_1817,N_13951,N_13448);
and UO_1818 (O_1818,N_12675,N_14700);
nand UO_1819 (O_1819,N_13667,N_14946);
or UO_1820 (O_1820,N_12575,N_14496);
nand UO_1821 (O_1821,N_12368,N_14190);
or UO_1822 (O_1822,N_14055,N_12310);
nor UO_1823 (O_1823,N_13144,N_12889);
nand UO_1824 (O_1824,N_14692,N_14103);
or UO_1825 (O_1825,N_14747,N_14082);
or UO_1826 (O_1826,N_12038,N_12863);
nor UO_1827 (O_1827,N_12559,N_12691);
nor UO_1828 (O_1828,N_13946,N_13462);
nor UO_1829 (O_1829,N_13533,N_14011);
nor UO_1830 (O_1830,N_14846,N_12439);
and UO_1831 (O_1831,N_13722,N_13199);
nor UO_1832 (O_1832,N_14771,N_12581);
nand UO_1833 (O_1833,N_13607,N_13927);
and UO_1834 (O_1834,N_12404,N_13484);
or UO_1835 (O_1835,N_14187,N_14702);
and UO_1836 (O_1836,N_13664,N_14535);
nand UO_1837 (O_1837,N_14100,N_13231);
and UO_1838 (O_1838,N_13701,N_14061);
and UO_1839 (O_1839,N_14257,N_13395);
nand UO_1840 (O_1840,N_12566,N_13165);
nor UO_1841 (O_1841,N_13923,N_13965);
nor UO_1842 (O_1842,N_12344,N_13036);
nand UO_1843 (O_1843,N_12923,N_12674);
or UO_1844 (O_1844,N_13635,N_13094);
or UO_1845 (O_1845,N_14812,N_12485);
nor UO_1846 (O_1846,N_13425,N_14534);
nand UO_1847 (O_1847,N_13681,N_12822);
nand UO_1848 (O_1848,N_14963,N_12627);
or UO_1849 (O_1849,N_13377,N_13200);
nor UO_1850 (O_1850,N_12359,N_12858);
nor UO_1851 (O_1851,N_13053,N_14376);
nand UO_1852 (O_1852,N_12990,N_12336);
nand UO_1853 (O_1853,N_13509,N_14871);
nor UO_1854 (O_1854,N_13982,N_14865);
and UO_1855 (O_1855,N_12700,N_13093);
or UO_1856 (O_1856,N_12476,N_13136);
nor UO_1857 (O_1857,N_12941,N_13384);
or UO_1858 (O_1858,N_12119,N_14010);
nand UO_1859 (O_1859,N_14045,N_13208);
and UO_1860 (O_1860,N_14092,N_12044);
nor UO_1861 (O_1861,N_13818,N_12779);
nand UO_1862 (O_1862,N_14771,N_12021);
nor UO_1863 (O_1863,N_13305,N_13569);
nor UO_1864 (O_1864,N_14530,N_13935);
xor UO_1865 (O_1865,N_14063,N_12616);
xor UO_1866 (O_1866,N_12037,N_13250);
or UO_1867 (O_1867,N_12099,N_12159);
and UO_1868 (O_1868,N_14854,N_12776);
or UO_1869 (O_1869,N_13795,N_12797);
and UO_1870 (O_1870,N_12442,N_12740);
or UO_1871 (O_1871,N_13302,N_12540);
nand UO_1872 (O_1872,N_14017,N_12593);
or UO_1873 (O_1873,N_14566,N_13834);
nor UO_1874 (O_1874,N_13116,N_13481);
nand UO_1875 (O_1875,N_12174,N_12987);
and UO_1876 (O_1876,N_12227,N_12572);
and UO_1877 (O_1877,N_12961,N_12470);
or UO_1878 (O_1878,N_14517,N_14440);
nand UO_1879 (O_1879,N_14810,N_14819);
or UO_1880 (O_1880,N_12146,N_12482);
nand UO_1881 (O_1881,N_13394,N_14850);
nand UO_1882 (O_1882,N_12758,N_12230);
or UO_1883 (O_1883,N_13250,N_14703);
nor UO_1884 (O_1884,N_14512,N_12283);
and UO_1885 (O_1885,N_12737,N_13570);
nor UO_1886 (O_1886,N_12660,N_14569);
nand UO_1887 (O_1887,N_14586,N_13680);
and UO_1888 (O_1888,N_13097,N_13769);
and UO_1889 (O_1889,N_13834,N_13282);
or UO_1890 (O_1890,N_14890,N_13843);
nand UO_1891 (O_1891,N_13456,N_13221);
nor UO_1892 (O_1892,N_12903,N_12052);
nand UO_1893 (O_1893,N_12829,N_12495);
nor UO_1894 (O_1894,N_14803,N_14487);
and UO_1895 (O_1895,N_13392,N_14755);
nor UO_1896 (O_1896,N_14599,N_14026);
and UO_1897 (O_1897,N_13491,N_14729);
and UO_1898 (O_1898,N_14631,N_13401);
or UO_1899 (O_1899,N_14418,N_13556);
and UO_1900 (O_1900,N_12792,N_13709);
nor UO_1901 (O_1901,N_14942,N_13679);
nor UO_1902 (O_1902,N_12626,N_13720);
and UO_1903 (O_1903,N_12119,N_13344);
nor UO_1904 (O_1904,N_14274,N_12858);
or UO_1905 (O_1905,N_12361,N_13843);
nor UO_1906 (O_1906,N_14024,N_14666);
nor UO_1907 (O_1907,N_12465,N_14202);
nor UO_1908 (O_1908,N_13695,N_14408);
or UO_1909 (O_1909,N_14585,N_12615);
xnor UO_1910 (O_1910,N_14858,N_12055);
or UO_1911 (O_1911,N_12110,N_14813);
and UO_1912 (O_1912,N_12685,N_14448);
and UO_1913 (O_1913,N_12892,N_14761);
or UO_1914 (O_1914,N_13765,N_13115);
nor UO_1915 (O_1915,N_13032,N_13782);
nor UO_1916 (O_1916,N_12525,N_12067);
nor UO_1917 (O_1917,N_12847,N_13262);
and UO_1918 (O_1918,N_14721,N_13832);
or UO_1919 (O_1919,N_14385,N_13400);
nand UO_1920 (O_1920,N_13400,N_13802);
and UO_1921 (O_1921,N_14910,N_14959);
nand UO_1922 (O_1922,N_14399,N_14022);
or UO_1923 (O_1923,N_14298,N_13651);
and UO_1924 (O_1924,N_14816,N_13483);
or UO_1925 (O_1925,N_14044,N_14036);
nand UO_1926 (O_1926,N_12679,N_13578);
or UO_1927 (O_1927,N_14831,N_13674);
nand UO_1928 (O_1928,N_14920,N_13600);
and UO_1929 (O_1929,N_12370,N_14260);
nor UO_1930 (O_1930,N_14492,N_14726);
or UO_1931 (O_1931,N_14141,N_13471);
nor UO_1932 (O_1932,N_14377,N_13959);
or UO_1933 (O_1933,N_13713,N_12915);
xnor UO_1934 (O_1934,N_14158,N_14336);
and UO_1935 (O_1935,N_13496,N_13734);
or UO_1936 (O_1936,N_14166,N_14436);
nor UO_1937 (O_1937,N_14427,N_12038);
nor UO_1938 (O_1938,N_12237,N_14687);
or UO_1939 (O_1939,N_14296,N_12735);
nand UO_1940 (O_1940,N_12770,N_13981);
nand UO_1941 (O_1941,N_14284,N_13460);
or UO_1942 (O_1942,N_14309,N_14863);
nor UO_1943 (O_1943,N_14619,N_13450);
and UO_1944 (O_1944,N_12313,N_14931);
and UO_1945 (O_1945,N_12668,N_14628);
or UO_1946 (O_1946,N_14344,N_13388);
nor UO_1947 (O_1947,N_14300,N_14472);
nor UO_1948 (O_1948,N_14264,N_12790);
and UO_1949 (O_1949,N_13835,N_12260);
nor UO_1950 (O_1950,N_12105,N_13420);
nor UO_1951 (O_1951,N_13594,N_13074);
nand UO_1952 (O_1952,N_13094,N_12415);
nor UO_1953 (O_1953,N_14765,N_12940);
and UO_1954 (O_1954,N_13639,N_12013);
nand UO_1955 (O_1955,N_12734,N_12840);
nand UO_1956 (O_1956,N_12267,N_13526);
nor UO_1957 (O_1957,N_12762,N_13937);
and UO_1958 (O_1958,N_12777,N_13580);
or UO_1959 (O_1959,N_14532,N_13726);
and UO_1960 (O_1960,N_14268,N_12287);
nor UO_1961 (O_1961,N_13054,N_14750);
and UO_1962 (O_1962,N_14559,N_14039);
nand UO_1963 (O_1963,N_12429,N_12484);
nand UO_1964 (O_1964,N_13201,N_12598);
nand UO_1965 (O_1965,N_14900,N_14871);
or UO_1966 (O_1966,N_13191,N_14651);
nor UO_1967 (O_1967,N_14112,N_14395);
nand UO_1968 (O_1968,N_14726,N_12945);
nor UO_1969 (O_1969,N_13464,N_13705);
and UO_1970 (O_1970,N_14194,N_14638);
or UO_1971 (O_1971,N_13392,N_14121);
nand UO_1972 (O_1972,N_14586,N_13578);
or UO_1973 (O_1973,N_13172,N_14155);
nand UO_1974 (O_1974,N_12100,N_12602);
nor UO_1975 (O_1975,N_14590,N_12973);
nand UO_1976 (O_1976,N_13564,N_13903);
nand UO_1977 (O_1977,N_13247,N_13115);
nor UO_1978 (O_1978,N_13621,N_12406);
or UO_1979 (O_1979,N_14520,N_13712);
nand UO_1980 (O_1980,N_12360,N_14434);
nand UO_1981 (O_1981,N_14838,N_14082);
or UO_1982 (O_1982,N_13463,N_14560);
and UO_1983 (O_1983,N_13249,N_14623);
nor UO_1984 (O_1984,N_14754,N_12811);
or UO_1985 (O_1985,N_13751,N_12973);
and UO_1986 (O_1986,N_13064,N_14031);
nor UO_1987 (O_1987,N_13162,N_12977);
xnor UO_1988 (O_1988,N_12534,N_12567);
nor UO_1989 (O_1989,N_13153,N_13458);
and UO_1990 (O_1990,N_14809,N_14621);
nor UO_1991 (O_1991,N_12386,N_13804);
nor UO_1992 (O_1992,N_13127,N_14363);
or UO_1993 (O_1993,N_12345,N_13776);
nand UO_1994 (O_1994,N_13467,N_14128);
nor UO_1995 (O_1995,N_13983,N_12447);
nand UO_1996 (O_1996,N_13711,N_14606);
or UO_1997 (O_1997,N_13367,N_12853);
nor UO_1998 (O_1998,N_14680,N_12098);
nor UO_1999 (O_1999,N_13452,N_13240);
endmodule