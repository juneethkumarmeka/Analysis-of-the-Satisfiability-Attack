module basic_1500_15000_2000_20_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_739,In_439);
nor U1 (N_1,In_1241,In_1455);
nand U2 (N_2,In_7,In_394);
and U3 (N_3,In_370,In_1458);
nand U4 (N_4,In_565,In_538);
or U5 (N_5,In_485,In_1035);
and U6 (N_6,In_218,In_558);
nand U7 (N_7,In_285,In_411);
xnor U8 (N_8,In_268,In_1341);
and U9 (N_9,In_647,In_964);
nand U10 (N_10,In_543,In_1115);
nand U11 (N_11,In_881,In_573);
xnor U12 (N_12,In_862,In_621);
and U13 (N_13,In_2,In_1183);
xor U14 (N_14,In_101,In_1057);
nand U15 (N_15,In_900,In_474);
and U16 (N_16,In_1348,In_1365);
nor U17 (N_17,In_884,In_904);
or U18 (N_18,In_89,In_1310);
or U19 (N_19,In_898,In_812);
nor U20 (N_20,In_859,In_1405);
or U21 (N_21,In_288,In_144);
nand U22 (N_22,In_1077,In_530);
and U23 (N_23,In_194,In_691);
nand U24 (N_24,In_374,In_779);
nor U25 (N_25,In_954,In_238);
xor U26 (N_26,In_1097,In_567);
nor U27 (N_27,In_1076,In_1343);
nand U28 (N_28,In_293,In_1132);
nand U29 (N_29,In_979,In_86);
nand U30 (N_30,In_639,In_1443);
and U31 (N_31,In_1095,In_211);
nor U32 (N_32,In_1001,In_1224);
nor U33 (N_33,In_416,In_1431);
nand U34 (N_34,In_1047,In_927);
nand U35 (N_35,In_747,In_1049);
nand U36 (N_36,In_432,In_174);
xor U37 (N_37,In_891,In_1473);
nor U38 (N_38,In_600,In_939);
nand U39 (N_39,In_789,In_1381);
nor U40 (N_40,In_1475,In_1158);
nor U41 (N_41,In_1075,In_1402);
nand U42 (N_42,In_1234,In_1248);
xor U43 (N_43,In_69,In_913);
or U44 (N_44,In_460,In_990);
or U45 (N_45,In_188,In_1321);
nor U46 (N_46,In_157,In_1331);
and U47 (N_47,In_824,In_88);
xnor U48 (N_48,In_587,In_1229);
or U49 (N_49,In_822,In_741);
nor U50 (N_50,In_933,In_1033);
nor U51 (N_51,In_1476,In_865);
nor U52 (N_52,In_793,In_477);
or U53 (N_53,In_184,In_1399);
and U54 (N_54,In_58,In_1107);
or U55 (N_55,In_611,In_751);
nand U56 (N_56,In_29,In_577);
xnor U57 (N_57,In_199,In_1154);
nand U58 (N_58,In_914,In_1459);
or U59 (N_59,In_1019,In_254);
nand U60 (N_60,In_905,In_450);
nor U61 (N_61,In_415,In_584);
or U62 (N_62,In_269,In_81);
xor U63 (N_63,In_483,In_546);
or U64 (N_64,In_1171,In_452);
nand U65 (N_65,In_1370,In_471);
xnor U66 (N_66,In_1438,In_781);
xnor U67 (N_67,In_361,In_1194);
and U68 (N_68,In_1336,In_1188);
and U69 (N_69,In_1034,In_770);
xor U70 (N_70,In_16,In_245);
and U71 (N_71,In_892,In_1000);
xnor U72 (N_72,In_632,In_1065);
and U73 (N_73,In_1299,In_518);
nor U74 (N_74,In_1307,In_65);
nor U75 (N_75,In_525,In_1335);
nor U76 (N_76,In_1182,In_1123);
nor U77 (N_77,In_1017,In_1113);
xnor U78 (N_78,In_523,In_240);
nor U79 (N_79,In_602,In_138);
nand U80 (N_80,In_903,In_1337);
and U81 (N_81,In_668,In_1340);
or U82 (N_82,In_740,In_942);
nand U83 (N_83,In_513,In_412);
and U84 (N_84,In_986,In_1009);
xnor U85 (N_85,In_1302,In_329);
and U86 (N_86,In_1084,In_236);
and U87 (N_87,In_10,In_1108);
nor U88 (N_88,In_266,In_360);
and U89 (N_89,In_938,In_868);
xor U90 (N_90,In_1435,In_826);
and U91 (N_91,In_794,In_335);
nand U92 (N_92,In_461,In_953);
or U93 (N_93,In_1347,In_612);
nand U94 (N_94,In_1413,In_975);
or U95 (N_95,In_1338,In_931);
xor U96 (N_96,In_1414,In_478);
and U97 (N_97,In_589,In_1135);
or U98 (N_98,In_1373,In_897);
xor U99 (N_99,In_50,In_212);
or U100 (N_100,In_948,In_465);
and U101 (N_101,In_1282,In_1324);
nand U102 (N_102,In_1422,In_665);
nor U103 (N_103,In_1040,In_800);
or U104 (N_104,In_338,In_99);
nor U105 (N_105,In_76,In_133);
nand U106 (N_106,In_1272,In_278);
or U107 (N_107,In_634,In_977);
or U108 (N_108,In_108,In_12);
nand U109 (N_109,In_104,In_1225);
and U110 (N_110,In_1051,In_1385);
and U111 (N_111,In_425,In_858);
xnor U112 (N_112,In_150,In_1472);
xnor U113 (N_113,In_1279,In_141);
xnor U114 (N_114,In_1327,In_701);
and U115 (N_115,In_856,In_274);
or U116 (N_116,In_493,In_875);
xor U117 (N_117,In_1,In_1316);
nand U118 (N_118,In_1461,In_1334);
nor U119 (N_119,In_857,In_289);
and U120 (N_120,In_429,In_186);
nor U121 (N_121,In_1361,In_291);
or U122 (N_122,In_733,In_275);
and U123 (N_123,In_1203,In_735);
or U124 (N_124,In_1469,In_1128);
and U125 (N_125,In_135,In_974);
nor U126 (N_126,In_785,In_1221);
and U127 (N_127,In_1322,In_1101);
and U128 (N_128,In_656,In_41);
xnor U129 (N_129,In_315,In_702);
and U130 (N_130,In_1199,In_165);
nor U131 (N_131,In_198,In_396);
xor U132 (N_132,In_1064,In_1265);
nor U133 (N_133,In_1329,In_154);
xnor U134 (N_134,In_455,In_514);
and U135 (N_135,In_623,In_916);
nor U136 (N_136,In_225,In_286);
xor U137 (N_137,In_220,In_1180);
nand U138 (N_138,In_1445,In_519);
nand U139 (N_139,In_322,In_1215);
nor U140 (N_140,In_579,In_1191);
or U141 (N_141,In_1434,In_1169);
xnor U142 (N_142,In_512,In_496);
or U143 (N_143,In_257,In_1484);
or U144 (N_144,In_724,In_805);
or U145 (N_145,In_1058,In_1143);
nor U146 (N_146,In_1492,In_379);
xor U147 (N_147,In_316,In_422);
nor U148 (N_148,In_1367,In_673);
nor U149 (N_149,In_405,In_1167);
nand U150 (N_150,In_552,In_105);
nand U151 (N_151,In_231,In_480);
nor U152 (N_152,In_1228,In_183);
xnor U153 (N_153,In_944,In_427);
or U154 (N_154,In_170,In_1004);
or U155 (N_155,In_797,In_290);
xor U156 (N_156,In_1111,In_633);
and U157 (N_157,In_676,In_593);
or U158 (N_158,In_835,In_766);
nand U159 (N_159,In_731,In_36);
and U160 (N_160,In_1073,In_949);
and U161 (N_161,In_339,In_851);
or U162 (N_162,In_517,In_428);
or U163 (N_163,In_650,In_524);
or U164 (N_164,In_988,In_1467);
xor U165 (N_165,In_119,In_486);
or U166 (N_166,In_1270,In_712);
nor U167 (N_167,In_147,In_1003);
xor U168 (N_168,In_1189,In_221);
nor U169 (N_169,In_31,In_1100);
or U170 (N_170,In_348,In_487);
and U171 (N_171,In_327,In_928);
xor U172 (N_172,In_1320,In_498);
nand U173 (N_173,In_1396,In_981);
nand U174 (N_174,In_784,In_210);
xor U175 (N_175,In_39,In_768);
and U176 (N_176,In_969,In_44);
and U177 (N_177,In_1330,In_372);
nand U178 (N_178,In_1397,In_957);
and U179 (N_179,In_753,In_57);
and U180 (N_180,In_1144,In_576);
or U181 (N_181,In_947,In_383);
or U182 (N_182,In_17,In_85);
nand U183 (N_183,In_1391,In_1301);
nand U184 (N_184,In_1355,In_355);
xnor U185 (N_185,In_500,In_1437);
xor U186 (N_186,In_1488,In_758);
xor U187 (N_187,In_563,In_532);
and U188 (N_188,In_259,In_759);
or U189 (N_189,In_306,In_201);
or U190 (N_190,In_582,In_746);
or U191 (N_191,In_219,In_677);
nand U192 (N_192,In_443,In_890);
or U193 (N_193,In_43,In_1202);
nor U194 (N_194,In_1483,In_776);
nor U195 (N_195,In_228,In_1345);
or U196 (N_196,In_1464,In_1263);
nor U197 (N_197,In_213,In_671);
nor U198 (N_198,In_510,In_205);
xnor U199 (N_199,In_653,In_1067);
nand U200 (N_200,In_490,In_566);
nand U201 (N_201,In_341,In_1403);
xor U202 (N_202,In_166,In_1031);
xor U203 (N_203,In_848,In_690);
and U204 (N_204,In_882,In_730);
nor U205 (N_205,In_49,In_1291);
or U206 (N_206,In_1247,In_1463);
and U207 (N_207,In_132,In_1448);
or U208 (N_208,In_1059,In_469);
xnor U209 (N_209,In_997,In_426);
or U210 (N_210,In_1447,In_375);
or U211 (N_211,In_1099,In_1262);
xnor U212 (N_212,In_5,In_630);
and U213 (N_213,In_1465,In_64);
xor U214 (N_214,In_1319,In_839);
nand U215 (N_215,In_25,In_273);
or U216 (N_216,In_63,In_707);
and U217 (N_217,In_1168,In_922);
nand U218 (N_218,In_161,In_276);
nor U219 (N_219,In_3,In_911);
or U220 (N_220,In_497,In_590);
and U221 (N_221,In_1214,In_755);
nand U222 (N_222,In_390,In_1245);
or U223 (N_223,In_686,In_1315);
and U224 (N_224,In_887,In_359);
nand U225 (N_225,In_271,In_1278);
xor U226 (N_226,In_818,In_795);
or U227 (N_227,In_651,In_1201);
xnor U228 (N_228,In_540,In_82);
or U229 (N_229,In_1333,In_1460);
and U230 (N_230,In_1165,In_125);
nor U231 (N_231,In_912,In_693);
nor U232 (N_232,In_1462,In_966);
and U233 (N_233,In_983,In_642);
and U234 (N_234,In_134,In_83);
and U235 (N_235,In_1032,In_610);
xor U236 (N_236,In_644,In_1478);
and U237 (N_237,In_246,In_1081);
or U238 (N_238,In_472,In_1028);
or U239 (N_239,In_1217,In_727);
nor U240 (N_240,In_773,In_250);
nand U241 (N_241,In_588,In_585);
or U242 (N_242,In_935,In_509);
or U243 (N_243,In_227,In_908);
xnor U244 (N_244,In_100,In_209);
xor U245 (N_245,In_629,In_1125);
nand U246 (N_246,In_403,In_237);
xor U247 (N_247,In_13,In_637);
nor U248 (N_248,In_1487,In_732);
nand U249 (N_249,In_1176,In_685);
xnor U250 (N_250,In_140,In_402);
or U251 (N_251,In_961,In_129);
xnor U252 (N_252,In_744,In_1060);
nor U253 (N_253,In_120,In_417);
nor U254 (N_254,In_1253,In_937);
nand U255 (N_255,In_247,In_958);
or U256 (N_256,In_813,In_1052);
nand U257 (N_257,In_1013,In_1016);
nor U258 (N_258,In_683,In_442);
or U259 (N_259,In_436,In_667);
nor U260 (N_260,In_1106,In_37);
or U261 (N_261,In_1486,In_24);
nor U262 (N_262,In_1219,In_548);
and U263 (N_263,In_204,In_745);
nand U264 (N_264,In_516,In_1220);
and U265 (N_265,In_466,In_243);
or U266 (N_266,In_1433,In_1091);
and U267 (N_267,In_754,In_1269);
xnor U268 (N_268,In_876,In_841);
nand U269 (N_269,In_762,In_896);
nand U270 (N_270,In_1145,In_367);
and U271 (N_271,In_815,In_1498);
or U272 (N_272,In_21,In_1493);
and U273 (N_273,In_458,In_777);
or U274 (N_274,In_94,In_714);
nor U275 (N_275,In_553,In_1120);
or U276 (N_276,In_222,In_1196);
and U277 (N_277,In_1292,In_114);
and U278 (N_278,In_1374,In_718);
or U279 (N_279,In_906,In_936);
and U280 (N_280,In_300,In_295);
nand U281 (N_281,In_309,In_711);
xnor U282 (N_282,In_1023,In_678);
xnor U283 (N_283,In_1068,In_1200);
or U284 (N_284,In_1139,In_1173);
nand U285 (N_285,In_200,In_1137);
nand U286 (N_286,In_1018,In_307);
nor U287 (N_287,In_583,In_993);
xnor U288 (N_288,In_454,In_726);
nand U289 (N_289,In_1179,In_1415);
and U290 (N_290,In_350,In_662);
nor U291 (N_291,In_998,In_457);
nor U292 (N_292,In_1131,In_1339);
xnor U293 (N_293,In_1261,In_1133);
nand U294 (N_294,In_84,In_654);
nand U295 (N_295,In_1376,In_1046);
or U296 (N_296,In_305,In_1289);
xnor U297 (N_297,In_1452,In_1477);
nor U298 (N_298,In_279,In_1369);
nand U299 (N_299,In_527,In_595);
nor U300 (N_300,In_1074,In_502);
xor U301 (N_301,In_929,In_470);
or U302 (N_302,In_1240,In_146);
xnor U303 (N_303,In_4,In_494);
nor U304 (N_304,In_111,In_1312);
nor U305 (N_305,In_399,In_169);
nand U306 (N_306,In_1386,In_202);
xnor U307 (N_307,In_1495,In_1233);
xor U308 (N_308,In_666,In_627);
or U309 (N_309,In_889,In_340);
nand U310 (N_310,In_575,In_1162);
nor U311 (N_311,In_1086,In_287);
nand U312 (N_312,In_301,In_1193);
xor U313 (N_313,In_1406,In_251);
nand U314 (N_314,In_1457,In_1147);
or U315 (N_315,In_915,In_734);
nand U316 (N_316,In_1436,In_1249);
and U317 (N_317,In_765,In_831);
nand U318 (N_318,In_1298,In_35);
nor U319 (N_319,In_1276,In_1407);
nor U320 (N_320,In_468,In_729);
nor U321 (N_321,In_1449,In_333);
xnor U322 (N_322,In_1371,In_1377);
and U323 (N_323,In_167,In_1104);
nand U324 (N_324,In_1260,In_413);
xnor U325 (N_325,In_453,In_349);
xnor U326 (N_326,In_825,In_449);
nor U327 (N_327,In_1366,In_385);
nand U328 (N_328,In_529,In_956);
xnor U329 (N_329,In_750,In_1379);
nor U330 (N_330,In_1204,In_657);
and U331 (N_331,In_456,In_1007);
or U332 (N_332,In_177,In_1134);
or U333 (N_333,In_572,In_1267);
or U334 (N_334,In_1352,In_1083);
xnor U335 (N_335,In_1071,In_294);
and U336 (N_336,In_79,In_946);
and U337 (N_337,In_122,In_680);
nor U338 (N_338,In_118,In_1286);
xor U339 (N_339,In_1208,In_767);
or U340 (N_340,In_814,In_1206);
nor U341 (N_341,In_811,In_854);
xor U342 (N_342,In_864,In_1395);
and U343 (N_343,In_550,In_708);
xnor U344 (N_344,In_1170,In_431);
or U345 (N_345,In_995,In_1116);
and U346 (N_346,In_1417,In_280);
and U347 (N_347,In_581,In_533);
nand U348 (N_348,In_55,In_207);
nor U349 (N_349,In_378,In_934);
nand U350 (N_350,In_192,In_670);
nand U351 (N_351,In_725,In_1491);
xnor U352 (N_352,In_796,In_253);
xnor U353 (N_353,In_447,In_596);
or U354 (N_354,In_1243,In_778);
and U355 (N_355,In_531,In_311);
or U356 (N_356,In_679,In_1103);
xnor U357 (N_357,In_604,In_156);
nand U358 (N_358,In_1470,In_1372);
xor U359 (N_359,In_51,In_809);
or U360 (N_360,In_418,In_646);
nand U361 (N_361,In_1236,In_717);
xnor U362 (N_362,In_392,In_1063);
or U363 (N_363,In_1011,In_462);
and U364 (N_364,In_1380,In_1494);
xor U365 (N_365,In_866,In_823);
nand U366 (N_366,In_842,In_1479);
or U367 (N_367,In_1184,In_391);
xor U368 (N_368,In_1141,In_1306);
and U369 (N_369,In_1080,In_860);
nand U370 (N_370,In_1257,In_941);
or U371 (N_371,In_555,In_1497);
nand U372 (N_372,In_1044,In_902);
and U373 (N_373,In_420,In_560);
nor U374 (N_374,In_1042,In_663);
or U375 (N_375,In_499,In_1266);
nand U376 (N_376,In_505,In_96);
xor U377 (N_377,In_960,In_1002);
xnor U378 (N_378,In_1237,In_249);
or U379 (N_379,In_609,In_1079);
nand U380 (N_380,In_395,In_989);
xnor U381 (N_381,In_364,In_1358);
or U382 (N_382,In_414,In_47);
xor U383 (N_383,In_1037,In_551);
and U384 (N_384,In_1264,In_1281);
nand U385 (N_385,In_1382,In_782);
or U386 (N_386,In_1238,In_682);
nand U387 (N_387,In_557,In_388);
or U388 (N_388,In_821,In_780);
xor U389 (N_389,In_987,In_649);
and U390 (N_390,In_1275,In_318);
nor U391 (N_391,In_930,In_1378);
xnor U392 (N_392,In_74,In_615);
and U393 (N_393,In_1295,In_1025);
and U394 (N_394,In_334,In_508);
or U395 (N_395,In_1305,In_699);
nand U396 (N_396,In_863,In_636);
nand U397 (N_397,In_326,In_1129);
or U398 (N_398,In_27,In_121);
and U399 (N_399,In_586,In_1014);
xnor U400 (N_400,In_1485,In_262);
nor U401 (N_401,In_1441,In_526);
and U402 (N_402,In_893,In_1303);
nor U403 (N_403,In_445,In_397);
or U404 (N_404,In_536,In_234);
xor U405 (N_405,In_323,In_845);
and U406 (N_406,In_97,In_321);
nor U407 (N_407,In_1185,In_830);
xor U408 (N_408,In_808,In_1362);
nor U409 (N_409,In_115,In_1072);
nand U410 (N_410,In_272,In_1050);
nand U411 (N_411,In_534,In_8);
nand U412 (N_412,In_1251,In_233);
and U413 (N_413,In_599,In_45);
and U414 (N_414,In_410,In_68);
nand U415 (N_415,In_310,In_371);
nand U416 (N_416,In_1400,In_1450);
and U417 (N_417,In_232,In_1172);
xnor U418 (N_418,In_267,In_325);
nor U419 (N_419,In_87,In_1043);
or U420 (N_420,In_675,In_1187);
or U421 (N_421,In_330,In_1294);
nand U422 (N_422,In_1412,In_1232);
xor U423 (N_423,In_819,In_1440);
nor U424 (N_424,In_1235,In_1216);
xnor U425 (N_425,In_1122,In_1280);
nand U426 (N_426,In_520,In_515);
and U427 (N_427,In_190,In_1388);
or U428 (N_428,In_1259,In_806);
nand U429 (N_429,In_1323,In_1268);
nand U430 (N_430,In_886,In_568);
xnor U431 (N_431,In_265,In_1480);
or U432 (N_432,In_1140,In_384);
nand U433 (N_433,In_924,In_26);
nor U434 (N_434,In_569,In_803);
xnor U435 (N_435,In_158,In_365);
and U436 (N_436,In_996,In_18);
nand U437 (N_437,In_737,In_570);
nor U438 (N_438,In_1242,In_620);
or U439 (N_439,In_1098,In_304);
and U440 (N_440,In_380,In_720);
or U441 (N_441,In_578,In_230);
xnor U442 (N_442,In_423,In_719);
nor U443 (N_443,In_95,In_828);
xnor U444 (N_444,In_1346,In_542);
xor U445 (N_445,In_674,In_1390);
and U446 (N_446,In_377,In_102);
and U447 (N_447,In_638,In_1102);
xor U448 (N_448,In_1421,In_1481);
or U449 (N_449,In_1246,In_624);
or U450 (N_450,In_888,In_482);
nand U451 (N_451,In_319,In_217);
xnor U452 (N_452,In_698,In_116);
or U453 (N_453,In_1420,In_1054);
nand U454 (N_454,In_1094,In_363);
xnor U455 (N_455,In_1062,In_464);
or U456 (N_456,In_618,In_879);
or U457 (N_457,In_343,In_208);
nor U458 (N_458,In_162,In_722);
nor U459 (N_459,In_761,In_258);
nand U460 (N_460,In_1112,In_645);
or U461 (N_461,In_625,In_1359);
or U462 (N_462,In_1138,In_1114);
and U463 (N_463,In_123,In_728);
nand U464 (N_464,In_910,In_742);
nand U465 (N_465,In_846,In_1451);
or U466 (N_466,In_78,In_107);
xnor U467 (N_467,In_992,In_738);
xnor U468 (N_468,In_1496,In_827);
nand U469 (N_469,In_131,In_715);
xnor U470 (N_470,In_556,In_664);
xnor U471 (N_471,In_605,In_149);
nor U472 (N_472,In_1087,In_829);
nor U473 (N_473,In_950,In_109);
xor U474 (N_474,In_1029,In_6);
xor U475 (N_475,In_537,In_1368);
nor U476 (N_476,In_571,In_619);
nand U477 (N_477,In_435,In_28);
nand U478 (N_478,In_895,In_919);
xnor U479 (N_479,In_283,In_959);
nor U480 (N_480,In_196,In_72);
nand U481 (N_481,In_172,In_1157);
or U482 (N_482,In_117,In_1078);
xnor U483 (N_483,In_346,In_985);
xnor U484 (N_484,In_491,In_978);
and U485 (N_485,In_1300,In_1210);
nor U486 (N_486,In_1211,In_23);
and U487 (N_487,In_313,In_790);
xnor U488 (N_488,In_106,In_607);
nand U489 (N_489,In_299,In_869);
nor U490 (N_490,In_1041,In_475);
xnor U491 (N_491,In_616,In_635);
nand U492 (N_492,In_1363,In_688);
or U493 (N_493,In_126,In_195);
nand U494 (N_494,In_434,In_1213);
nor U495 (N_495,In_332,In_277);
nor U496 (N_496,In_1296,In_270);
or U497 (N_497,In_788,In_539);
and U498 (N_498,In_226,In_59);
and U499 (N_499,In_446,In_393);
nand U500 (N_500,In_92,In_139);
and U501 (N_501,In_1012,In_1222);
or U502 (N_502,In_541,In_982);
nor U503 (N_503,In_1198,In_401);
xnor U504 (N_504,In_1432,In_1231);
or U505 (N_505,In_695,In_1288);
nor U506 (N_506,In_603,In_19);
nor U507 (N_507,In_1425,In_1411);
xor U508 (N_508,In_1332,In_1121);
xor U509 (N_509,In_1293,In_1124);
xnor U510 (N_510,In_574,In_820);
nand U511 (N_511,In_705,In_783);
nor U512 (N_512,In_1195,In_775);
nor U513 (N_513,In_1313,In_369);
nor U514 (N_514,In_554,In_504);
xnor U515 (N_515,In_1155,In_352);
and U516 (N_516,In_424,In_894);
xor U517 (N_517,In_984,In_1244);
or U518 (N_518,In_356,In_951);
nand U519 (N_519,In_203,In_1283);
nor U520 (N_520,In_873,In_1127);
nor U521 (N_521,In_362,In_93);
or U522 (N_522,In_20,In_175);
and U523 (N_523,In_713,In_489);
xnor U524 (N_524,In_689,In_1088);
xnor U525 (N_525,In_836,In_907);
nor U526 (N_526,In_1166,In_155);
nor U527 (N_527,In_791,In_849);
or U528 (N_528,In_1163,In_1252);
or U529 (N_529,In_1393,In_160);
and U530 (N_530,In_235,In_1178);
or U531 (N_531,In_1105,In_206);
nand U532 (N_532,In_66,In_774);
nor U533 (N_533,In_1285,In_1159);
and U534 (N_534,In_1349,In_127);
or U535 (N_535,In_952,In_967);
xnor U536 (N_536,In_1325,In_844);
xor U537 (N_537,In_77,In_1350);
nand U538 (N_538,In_792,In_448);
and U539 (N_539,In_264,In_580);
xnor U540 (N_540,In_1148,In_1021);
xnor U541 (N_541,In_53,In_798);
or U542 (N_542,In_302,In_787);
and U543 (N_543,In_973,In_853);
nand U544 (N_544,In_1468,In_9);
and U545 (N_545,In_430,In_103);
nor U546 (N_546,In_1297,In_1416);
nor U547 (N_547,In_142,In_917);
nor U548 (N_548,In_1230,In_56);
or U549 (N_549,In_1174,In_1039);
xnor U550 (N_550,In_1177,In_617);
xor U551 (N_551,In_1284,In_506);
nand U552 (N_552,In_354,In_521);
nand U553 (N_553,In_655,In_337);
nor U554 (N_554,In_451,In_764);
or U555 (N_555,In_921,In_1093);
nor U556 (N_556,In_1326,In_613);
or U557 (N_557,In_381,In_1151);
xnor U558 (N_558,In_252,In_622);
nand U559 (N_559,In_312,In_1056);
nand U560 (N_560,In_296,In_769);
xnor U561 (N_561,In_871,In_1375);
nor U562 (N_562,In_706,In_672);
or U563 (N_563,In_970,In_1212);
and U564 (N_564,In_1454,In_1142);
nor U565 (N_565,In_816,In_11);
nor U566 (N_566,In_1256,In_837);
nand U567 (N_567,In_1197,In_54);
or U568 (N_568,In_877,In_626);
and U569 (N_569,In_1149,In_723);
nand U570 (N_570,In_999,In_382);
nor U571 (N_571,In_152,In_760);
nand U572 (N_572,In_1038,In_476);
nor U573 (N_573,In_182,In_168);
nand U574 (N_574,In_861,In_1356);
xor U575 (N_575,In_197,In_433);
xor U576 (N_576,In_492,In_178);
or U577 (N_577,In_899,In_242);
or U578 (N_578,In_669,In_965);
and U579 (N_579,In_73,In_1427);
nand U580 (N_580,In_511,In_32);
nor U581 (N_581,In_328,In_15);
nor U582 (N_582,In_223,In_1273);
and U583 (N_583,In_255,In_1353);
or U584 (N_584,In_153,In_1090);
nor U585 (N_585,In_692,In_389);
or U586 (N_586,In_1022,In_1453);
or U587 (N_587,In_34,In_641);
nand U588 (N_588,In_547,In_1401);
and U589 (N_589,In_1027,In_1156);
nor U590 (N_590,In_1255,In_185);
xnor U591 (N_591,In_991,In_62);
xor U592 (N_592,In_878,In_1398);
or U593 (N_593,In_628,In_1499);
nor U594 (N_594,In_592,In_1070);
and U595 (N_595,In_799,In_810);
and U596 (N_596,In_1389,In_1239);
nand U597 (N_597,In_923,In_801);
nand U598 (N_598,In_1392,In_358);
nand U599 (N_599,In_159,In_920);
nand U600 (N_600,In_357,In_976);
or U601 (N_601,In_1092,In_1429);
or U602 (N_602,In_1066,In_696);
xnor U603 (N_603,In_1344,In_1471);
nand U604 (N_604,In_1419,In_1410);
or U605 (N_605,In_867,In_1020);
or U606 (N_606,In_1360,In_400);
nand U607 (N_607,In_1126,In_260);
or U608 (N_608,In_1005,In_256);
xnor U609 (N_609,In_239,In_75);
or U610 (N_610,In_1418,In_344);
nand U611 (N_611,In_1164,In_1036);
and U612 (N_612,In_1010,In_1277);
nor U613 (N_613,In_709,In_98);
and U614 (N_614,In_33,In_1474);
xnor U615 (N_615,In_1423,In_872);
nand U616 (N_616,In_901,In_870);
and U617 (N_617,In_1110,In_855);
and U618 (N_618,In_1342,In_1318);
and U619 (N_619,In_112,In_61);
xnor U620 (N_620,In_67,In_1152);
nor U621 (N_621,In_704,In_187);
xnor U622 (N_622,In_1308,In_535);
nand U623 (N_623,In_1311,In_70);
and U624 (N_624,In_661,In_314);
xor U625 (N_625,In_601,In_324);
xnor U626 (N_626,In_1439,In_136);
and U627 (N_627,In_694,In_681);
xnor U628 (N_628,In_945,In_488);
nand U629 (N_629,In_1205,In_22);
and U630 (N_630,In_833,In_110);
nand U631 (N_631,In_1136,In_282);
nor U632 (N_632,In_748,In_561);
and U633 (N_633,In_351,In_1045);
nand U634 (N_634,In_926,In_1055);
and U635 (N_635,In_652,In_366);
nand U636 (N_636,In_1192,In_1085);
or U637 (N_637,In_1430,In_215);
or U638 (N_638,In_331,In_1364);
and U639 (N_639,In_137,In_438);
and U640 (N_640,In_697,In_522);
xnor U641 (N_641,In_163,In_216);
or U642 (N_642,In_376,In_549);
xor U643 (N_643,In_971,In_387);
xor U644 (N_644,In_749,In_1384);
nor U645 (N_645,In_559,In_467);
nand U646 (N_646,In_786,In_1008);
nor U647 (N_647,In_716,In_598);
and U648 (N_648,In_643,In_1109);
nand U649 (N_649,In_721,In_407);
nor U650 (N_650,In_1271,In_148);
and U651 (N_651,In_48,In_736);
xor U652 (N_652,In_398,In_320);
nand U653 (N_653,In_1409,In_38);
nand U654 (N_654,In_440,In_71);
and U655 (N_655,In_345,In_193);
nand U656 (N_656,In_308,In_1024);
nor U657 (N_657,In_180,In_1490);
and U658 (N_658,In_838,In_0);
or U659 (N_659,In_91,In_963);
xnor U660 (N_660,In_191,In_281);
or U661 (N_661,In_176,In_703);
and U662 (N_662,In_42,In_317);
xor U663 (N_663,In_80,In_687);
nor U664 (N_664,In_40,In_437);
xnor U665 (N_665,In_463,In_1404);
xor U666 (N_666,In_248,In_292);
xnor U667 (N_667,In_128,In_757);
and U668 (N_668,In_1328,In_1048);
nand U669 (N_669,In_1181,In_503);
nand U670 (N_670,In_444,In_1190);
nand U671 (N_671,In_684,In_479);
nand U672 (N_672,In_885,In_1226);
and U673 (N_673,In_495,In_484);
nand U674 (N_674,In_124,In_189);
nand U675 (N_675,In_342,In_1274);
nor U676 (N_676,In_880,In_752);
and U677 (N_677,In_90,In_261);
nor U678 (N_678,In_113,In_459);
xor U679 (N_679,In_631,In_883);
xor U680 (N_680,In_284,In_597);
and U681 (N_681,In_807,In_771);
nor U682 (N_682,In_473,In_1254);
or U683 (N_683,In_481,In_60);
xor U684 (N_684,In_772,In_421);
and U685 (N_685,In_817,In_528);
nor U686 (N_686,In_336,In_1482);
or U687 (N_687,In_710,In_1150);
nand U688 (N_688,In_244,In_659);
nand U689 (N_689,In_46,In_130);
or U690 (N_690,In_1146,In_297);
nand U691 (N_691,In_419,In_1309);
and U692 (N_692,In_1314,In_1444);
xor U693 (N_693,In_1096,In_368);
nor U694 (N_694,In_606,In_1466);
nor U695 (N_695,In_145,In_840);
and U696 (N_696,In_501,In_1026);
and U697 (N_697,In_1258,In_962);
nor U698 (N_698,In_648,In_1118);
and U699 (N_699,In_850,In_1387);
or U700 (N_700,In_1354,In_1304);
nand U701 (N_701,In_658,In_1119);
nand U702 (N_702,In_834,In_179);
nand U703 (N_703,In_241,In_1061);
nor U704 (N_704,In_1117,In_1351);
nor U705 (N_705,In_1456,In_1069);
nand U706 (N_706,In_544,In_224);
and U707 (N_707,In_1082,In_1489);
nand U708 (N_708,In_171,In_1428);
or U709 (N_709,In_386,In_562);
or U710 (N_710,In_994,In_743);
or U711 (N_711,In_263,In_1227);
xnor U712 (N_712,In_1290,In_1357);
nand U713 (N_713,In_52,In_1130);
xor U714 (N_714,In_1250,In_1160);
or U715 (N_715,In_1030,In_1153);
nand U716 (N_716,In_832,In_164);
or U717 (N_717,In_406,In_847);
nand U718 (N_718,In_1207,In_972);
xnor U719 (N_719,In_980,In_564);
or U720 (N_720,In_441,In_1317);
nor U721 (N_721,In_614,In_143);
nor U722 (N_722,In_918,In_1394);
or U723 (N_723,In_909,In_173);
and U724 (N_724,In_660,In_874);
and U725 (N_725,In_852,In_408);
and U726 (N_726,In_932,In_404);
xor U727 (N_727,In_1218,In_802);
xor U728 (N_728,In_1383,In_1424);
xnor U729 (N_729,In_700,In_14);
or U730 (N_730,In_373,In_214);
or U731 (N_731,In_1015,In_1186);
or U732 (N_732,In_940,In_943);
nand U733 (N_733,In_763,In_1287);
nor U734 (N_734,In_968,In_1209);
and U735 (N_735,In_1006,In_181);
xor U736 (N_736,In_229,In_608);
and U737 (N_737,In_1446,In_594);
xnor U738 (N_738,In_804,In_545);
and U739 (N_739,In_298,In_409);
nand U740 (N_740,In_1442,In_591);
and U741 (N_741,In_1426,In_353);
and U742 (N_742,In_955,In_925);
nand U743 (N_743,In_1223,In_843);
and U744 (N_744,In_1408,In_30);
nand U745 (N_745,In_507,In_1053);
or U746 (N_746,In_347,In_151);
xnor U747 (N_747,In_640,In_1089);
nor U748 (N_748,In_1175,In_303);
nor U749 (N_749,In_756,In_1161);
nor U750 (N_750,N_146,N_587);
nand U751 (N_751,N_433,N_705);
nor U752 (N_752,N_684,N_621);
or U753 (N_753,N_330,N_21);
or U754 (N_754,N_106,N_565);
or U755 (N_755,N_525,N_137);
xor U756 (N_756,N_456,N_409);
or U757 (N_757,N_553,N_595);
and U758 (N_758,N_218,N_288);
or U759 (N_759,N_650,N_102);
and U760 (N_760,N_643,N_632);
xnor U761 (N_761,N_669,N_350);
nand U762 (N_762,N_136,N_356);
and U763 (N_763,N_361,N_37);
xor U764 (N_764,N_489,N_642);
and U765 (N_765,N_312,N_362);
nand U766 (N_766,N_408,N_316);
or U767 (N_767,N_130,N_385);
xnor U768 (N_768,N_484,N_696);
and U769 (N_769,N_543,N_220);
nand U770 (N_770,N_373,N_222);
xnor U771 (N_771,N_683,N_729);
nand U772 (N_772,N_129,N_503);
and U773 (N_773,N_331,N_521);
and U774 (N_774,N_282,N_675);
xnor U775 (N_775,N_631,N_386);
and U776 (N_776,N_510,N_244);
xnor U777 (N_777,N_44,N_536);
or U778 (N_778,N_89,N_736);
and U779 (N_779,N_267,N_325);
nor U780 (N_780,N_113,N_480);
nand U781 (N_781,N_114,N_431);
or U782 (N_782,N_402,N_201);
or U783 (N_783,N_447,N_699);
nor U784 (N_784,N_566,N_237);
xnor U785 (N_785,N_158,N_176);
xnor U786 (N_786,N_671,N_370);
nor U787 (N_787,N_294,N_628);
and U788 (N_788,N_550,N_27);
nand U789 (N_789,N_459,N_173);
xor U790 (N_790,N_403,N_635);
nand U791 (N_791,N_496,N_191);
or U792 (N_792,N_592,N_269);
or U793 (N_793,N_725,N_538);
xor U794 (N_794,N_345,N_138);
nand U795 (N_795,N_713,N_260);
and U796 (N_796,N_13,N_700);
nor U797 (N_797,N_453,N_31);
nand U798 (N_798,N_718,N_383);
xnor U799 (N_799,N_209,N_673);
xor U800 (N_800,N_71,N_256);
and U801 (N_801,N_1,N_227);
or U802 (N_802,N_142,N_380);
nor U803 (N_803,N_552,N_51);
xor U804 (N_804,N_285,N_300);
and U805 (N_805,N_240,N_667);
xnor U806 (N_806,N_69,N_309);
xnor U807 (N_807,N_108,N_66);
nand U808 (N_808,N_514,N_691);
xor U809 (N_809,N_204,N_81);
xnor U810 (N_810,N_737,N_645);
nor U811 (N_811,N_265,N_359);
nor U812 (N_812,N_687,N_225);
nand U813 (N_813,N_707,N_622);
and U814 (N_814,N_368,N_262);
or U815 (N_815,N_446,N_195);
and U816 (N_816,N_589,N_588);
xor U817 (N_817,N_630,N_103);
or U818 (N_818,N_732,N_636);
xnor U819 (N_819,N_374,N_463);
and U820 (N_820,N_223,N_170);
xnor U821 (N_821,N_164,N_407);
nor U822 (N_822,N_413,N_15);
nand U823 (N_823,N_96,N_284);
or U824 (N_824,N_17,N_697);
and U825 (N_825,N_417,N_556);
and U826 (N_826,N_723,N_199);
xnor U827 (N_827,N_353,N_275);
nand U828 (N_828,N_304,N_692);
nor U829 (N_829,N_662,N_612);
nand U830 (N_830,N_93,N_562);
or U831 (N_831,N_423,N_593);
xor U832 (N_832,N_286,N_245);
nand U833 (N_833,N_43,N_340);
and U834 (N_834,N_393,N_211);
or U835 (N_835,N_625,N_375);
xor U836 (N_836,N_726,N_418);
and U837 (N_837,N_255,N_336);
nand U838 (N_838,N_166,N_465);
xnor U839 (N_839,N_156,N_477);
nand U840 (N_840,N_695,N_348);
nor U841 (N_841,N_440,N_685);
nand U842 (N_842,N_523,N_122);
or U843 (N_843,N_689,N_185);
xor U844 (N_844,N_45,N_620);
or U845 (N_845,N_187,N_739);
nor U846 (N_846,N_357,N_711);
xnor U847 (N_847,N_399,N_243);
nor U848 (N_848,N_633,N_358);
xor U849 (N_849,N_470,N_153);
xor U850 (N_850,N_246,N_132);
xnor U851 (N_851,N_659,N_266);
xnor U852 (N_852,N_609,N_498);
xor U853 (N_853,N_35,N_747);
or U854 (N_854,N_61,N_268);
xnor U855 (N_855,N_213,N_212);
xor U856 (N_856,N_10,N_554);
nand U857 (N_857,N_60,N_454);
nand U858 (N_858,N_273,N_111);
xnor U859 (N_859,N_354,N_8);
nor U860 (N_860,N_257,N_512);
nor U861 (N_861,N_528,N_499);
and U862 (N_862,N_559,N_427);
xor U863 (N_863,N_253,N_539);
nand U864 (N_864,N_421,N_558);
nor U865 (N_865,N_75,N_67);
xnor U866 (N_866,N_197,N_139);
nor U867 (N_867,N_624,N_112);
and U868 (N_868,N_679,N_73);
nand U869 (N_869,N_120,N_363);
or U870 (N_870,N_604,N_742);
xor U871 (N_871,N_181,N_372);
nor U872 (N_872,N_657,N_546);
nor U873 (N_873,N_524,N_186);
or U874 (N_874,N_228,N_563);
and U875 (N_875,N_258,N_724);
nand U876 (N_876,N_339,N_264);
or U877 (N_877,N_730,N_200);
nand U878 (N_878,N_494,N_337);
xnor U879 (N_879,N_627,N_693);
or U880 (N_880,N_39,N_281);
and U881 (N_881,N_640,N_151);
nor U882 (N_882,N_59,N_414);
xor U883 (N_883,N_719,N_76);
xor U884 (N_884,N_492,N_217);
xnor U885 (N_885,N_46,N_415);
xnor U886 (N_886,N_475,N_276);
nand U887 (N_887,N_485,N_352);
or U888 (N_888,N_236,N_476);
nand U889 (N_889,N_332,N_449);
xor U890 (N_890,N_149,N_405);
or U891 (N_891,N_295,N_572);
nand U892 (N_892,N_99,N_749);
xor U893 (N_893,N_493,N_469);
nand U894 (N_894,N_569,N_517);
or U895 (N_895,N_157,N_148);
nor U896 (N_896,N_9,N_289);
nor U897 (N_897,N_184,N_744);
nand U898 (N_898,N_233,N_333);
and U899 (N_899,N_135,N_232);
nand U900 (N_900,N_655,N_457);
or U901 (N_901,N_500,N_63);
and U902 (N_902,N_670,N_717);
nor U903 (N_903,N_90,N_12);
and U904 (N_904,N_545,N_254);
and U905 (N_905,N_381,N_661);
xor U906 (N_906,N_682,N_419);
or U907 (N_907,N_637,N_490);
nand U908 (N_908,N_0,N_605);
nand U909 (N_909,N_516,N_586);
xnor U910 (N_910,N_634,N_389);
or U911 (N_911,N_28,N_377);
nand U912 (N_912,N_371,N_607);
or U913 (N_913,N_411,N_505);
xnor U914 (N_914,N_177,N_251);
nand U915 (N_915,N_443,N_664);
nand U916 (N_916,N_196,N_80);
or U917 (N_917,N_647,N_656);
nor U918 (N_918,N_74,N_585);
or U919 (N_919,N_384,N_648);
xnor U920 (N_920,N_738,N_573);
nand U921 (N_921,N_548,N_107);
xnor U922 (N_922,N_702,N_152);
xnor U923 (N_923,N_313,N_105);
nand U924 (N_924,N_714,N_745);
nand U925 (N_925,N_24,N_171);
or U926 (N_926,N_497,N_250);
or U927 (N_927,N_161,N_147);
nor U928 (N_928,N_83,N_663);
xor U929 (N_929,N_189,N_519);
nand U930 (N_930,N_29,N_610);
and U931 (N_931,N_623,N_50);
or U932 (N_932,N_396,N_513);
xor U933 (N_933,N_676,N_248);
or U934 (N_934,N_743,N_210);
nor U935 (N_935,N_561,N_296);
nor U936 (N_936,N_603,N_461);
nand U937 (N_937,N_509,N_401);
nand U938 (N_938,N_568,N_19);
xor U939 (N_939,N_133,N_551);
xor U940 (N_940,N_127,N_613);
xnor U941 (N_941,N_224,N_531);
xor U942 (N_942,N_507,N_712);
nand U943 (N_943,N_144,N_315);
and U944 (N_944,N_444,N_436);
xor U945 (N_945,N_704,N_741);
xnor U946 (N_946,N_291,N_540);
xor U947 (N_947,N_672,N_326);
nor U948 (N_948,N_280,N_347);
xnor U949 (N_949,N_279,N_706);
nor U950 (N_950,N_342,N_272);
nand U951 (N_951,N_644,N_159);
nor U952 (N_952,N_141,N_478);
and U953 (N_953,N_155,N_638);
nor U954 (N_954,N_52,N_508);
nor U955 (N_955,N_482,N_651);
and U956 (N_956,N_328,N_448);
or U957 (N_957,N_410,N_721);
xnor U958 (N_958,N_34,N_3);
and U959 (N_959,N_6,N_422);
xor U960 (N_960,N_307,N_179);
xnor U961 (N_961,N_183,N_581);
xnor U962 (N_962,N_247,N_343);
nand U963 (N_963,N_597,N_677);
nor U964 (N_964,N_302,N_178);
xor U965 (N_965,N_234,N_305);
or U966 (N_966,N_11,N_4);
xnor U967 (N_967,N_252,N_334);
nand U968 (N_968,N_594,N_488);
nand U969 (N_969,N_394,N_277);
or U970 (N_970,N_38,N_118);
nand U971 (N_971,N_733,N_101);
nand U972 (N_972,N_471,N_674);
nor U973 (N_973,N_95,N_53);
nand U974 (N_974,N_42,N_16);
or U975 (N_975,N_32,N_22);
or U976 (N_976,N_82,N_150);
nor U977 (N_977,N_208,N_533);
or U978 (N_978,N_263,N_278);
xor U979 (N_979,N_169,N_502);
or U980 (N_980,N_530,N_686);
nand U981 (N_981,N_270,N_117);
and U982 (N_982,N_207,N_165);
or U983 (N_983,N_694,N_221);
or U984 (N_984,N_335,N_583);
xor U985 (N_985,N_346,N_329);
nor U986 (N_986,N_420,N_626);
and U987 (N_987,N_481,N_703);
xnor U988 (N_988,N_571,N_229);
nand U989 (N_989,N_542,N_468);
and U990 (N_990,N_495,N_460);
nand U991 (N_991,N_33,N_549);
or U992 (N_992,N_190,N_48);
nor U993 (N_993,N_49,N_580);
nand U994 (N_994,N_297,N_445);
xnor U995 (N_995,N_7,N_64);
and U996 (N_996,N_491,N_666);
nand U997 (N_997,N_720,N_501);
xor U998 (N_998,N_526,N_698);
or U999 (N_999,N_483,N_474);
nor U1000 (N_1000,N_611,N_600);
and U1001 (N_1001,N_274,N_678);
and U1002 (N_1002,N_424,N_615);
nor U1003 (N_1003,N_646,N_175);
or U1004 (N_1004,N_716,N_654);
nor U1005 (N_1005,N_560,N_168);
nand U1006 (N_1006,N_437,N_355);
nor U1007 (N_1007,N_54,N_5);
or U1008 (N_1008,N_579,N_577);
nor U1009 (N_1009,N_570,N_665);
xor U1010 (N_1010,N_344,N_601);
xnor U1011 (N_1011,N_639,N_77);
and U1012 (N_1012,N_109,N_728);
nand U1013 (N_1013,N_504,N_55);
nor U1014 (N_1014,N_205,N_194);
nor U1015 (N_1015,N_486,N_219);
and U1016 (N_1016,N_544,N_430);
and U1017 (N_1017,N_608,N_230);
nor U1018 (N_1018,N_668,N_616);
nand U1019 (N_1019,N_464,N_40);
nand U1020 (N_1020,N_439,N_727);
nor U1021 (N_1021,N_557,N_391);
xnor U1022 (N_1022,N_319,N_310);
xnor U1023 (N_1023,N_215,N_462);
and U1024 (N_1024,N_203,N_72);
nor U1025 (N_1025,N_324,N_390);
nor U1026 (N_1026,N_681,N_429);
and U1027 (N_1027,N_351,N_534);
or U1028 (N_1028,N_473,N_41);
nand U1029 (N_1029,N_649,N_690);
or U1030 (N_1030,N_575,N_323);
nor U1031 (N_1031,N_116,N_366);
or U1032 (N_1032,N_110,N_365);
nor U1033 (N_1033,N_522,N_259);
nand U1034 (N_1034,N_172,N_98);
and U1035 (N_1035,N_94,N_740);
xnor U1036 (N_1036,N_126,N_541);
or U1037 (N_1037,N_722,N_92);
nor U1038 (N_1038,N_367,N_198);
nand U1039 (N_1039,N_748,N_14);
and U1040 (N_1040,N_458,N_70);
xnor U1041 (N_1041,N_596,N_584);
and U1042 (N_1042,N_65,N_62);
and U1043 (N_1043,N_360,N_341);
or U1044 (N_1044,N_241,N_452);
or U1045 (N_1045,N_283,N_406);
or U1046 (N_1046,N_78,N_298);
nor U1047 (N_1047,N_369,N_701);
xnor U1048 (N_1048,N_658,N_308);
nor U1049 (N_1049,N_314,N_617);
xor U1050 (N_1050,N_322,N_397);
xor U1051 (N_1051,N_97,N_472);
nand U1052 (N_1052,N_599,N_416);
nand U1053 (N_1053,N_555,N_709);
or U1054 (N_1054,N_85,N_487);
xor U1055 (N_1055,N_376,N_18);
nand U1056 (N_1056,N_746,N_455);
xor U1057 (N_1057,N_467,N_708);
nand U1058 (N_1058,N_364,N_321);
xnor U1059 (N_1059,N_518,N_123);
nand U1060 (N_1060,N_653,N_606);
nand U1061 (N_1061,N_84,N_134);
and U1062 (N_1062,N_602,N_162);
nor U1063 (N_1063,N_582,N_338);
nand U1064 (N_1064,N_388,N_527);
nand U1065 (N_1065,N_180,N_428);
and U1066 (N_1066,N_25,N_547);
xnor U1067 (N_1067,N_574,N_688);
nand U1068 (N_1068,N_680,N_404);
or U1069 (N_1069,N_154,N_578);
xnor U1070 (N_1070,N_271,N_400);
or U1071 (N_1071,N_318,N_249);
nor U1072 (N_1072,N_618,N_438);
nor U1073 (N_1073,N_327,N_140);
nor U1074 (N_1074,N_30,N_435);
nand U1075 (N_1075,N_731,N_2);
nand U1076 (N_1076,N_293,N_511);
nand U1077 (N_1077,N_299,N_590);
xnor U1078 (N_1078,N_192,N_231);
nor U1079 (N_1079,N_128,N_214);
or U1080 (N_1080,N_537,N_412);
or U1081 (N_1081,N_23,N_193);
nand U1082 (N_1082,N_124,N_104);
or U1083 (N_1083,N_660,N_182);
xnor U1084 (N_1084,N_317,N_652);
or U1085 (N_1085,N_379,N_292);
nand U1086 (N_1086,N_614,N_57);
xnor U1087 (N_1087,N_91,N_441);
xor U1088 (N_1088,N_68,N_506);
nor U1089 (N_1089,N_26,N_576);
xor U1090 (N_1090,N_529,N_515);
nand U1091 (N_1091,N_206,N_290);
or U1092 (N_1092,N_131,N_160);
nand U1093 (N_1093,N_301,N_567);
and U1094 (N_1094,N_392,N_479);
xnor U1095 (N_1095,N_320,N_303);
or U1096 (N_1096,N_202,N_629);
and U1097 (N_1097,N_242,N_710);
and U1098 (N_1098,N_86,N_36);
xnor U1099 (N_1099,N_735,N_216);
nor U1100 (N_1100,N_466,N_425);
nand U1101 (N_1101,N_306,N_115);
xor U1102 (N_1102,N_287,N_226);
nand U1103 (N_1103,N_87,N_100);
xor U1104 (N_1104,N_20,N_451);
nand U1105 (N_1105,N_235,N_398);
or U1106 (N_1106,N_167,N_520);
nand U1107 (N_1107,N_56,N_535);
nor U1108 (N_1108,N_311,N_734);
nor U1109 (N_1109,N_715,N_125);
nand U1110 (N_1110,N_532,N_619);
nor U1111 (N_1111,N_58,N_119);
xnor U1112 (N_1112,N_88,N_442);
or U1113 (N_1113,N_163,N_450);
or U1114 (N_1114,N_79,N_378);
xor U1115 (N_1115,N_434,N_143);
and U1116 (N_1116,N_598,N_174);
and U1117 (N_1117,N_395,N_261);
or U1118 (N_1118,N_382,N_239);
or U1119 (N_1119,N_47,N_641);
xnor U1120 (N_1120,N_432,N_426);
xor U1121 (N_1121,N_121,N_387);
xor U1122 (N_1122,N_591,N_238);
or U1123 (N_1123,N_564,N_145);
xor U1124 (N_1124,N_188,N_349);
nor U1125 (N_1125,N_9,N_182);
nor U1126 (N_1126,N_732,N_327);
or U1127 (N_1127,N_197,N_646);
xor U1128 (N_1128,N_620,N_344);
nor U1129 (N_1129,N_231,N_94);
xor U1130 (N_1130,N_723,N_129);
or U1131 (N_1131,N_365,N_654);
or U1132 (N_1132,N_713,N_39);
or U1133 (N_1133,N_469,N_608);
or U1134 (N_1134,N_663,N_521);
nand U1135 (N_1135,N_374,N_559);
and U1136 (N_1136,N_622,N_500);
and U1137 (N_1137,N_93,N_302);
nor U1138 (N_1138,N_137,N_328);
or U1139 (N_1139,N_541,N_630);
and U1140 (N_1140,N_695,N_195);
xnor U1141 (N_1141,N_193,N_174);
or U1142 (N_1142,N_534,N_43);
and U1143 (N_1143,N_24,N_368);
nor U1144 (N_1144,N_476,N_697);
nor U1145 (N_1145,N_196,N_172);
nand U1146 (N_1146,N_225,N_445);
nand U1147 (N_1147,N_133,N_276);
nand U1148 (N_1148,N_45,N_242);
nor U1149 (N_1149,N_515,N_255);
or U1150 (N_1150,N_426,N_428);
xor U1151 (N_1151,N_465,N_446);
xnor U1152 (N_1152,N_579,N_249);
nand U1153 (N_1153,N_549,N_621);
xnor U1154 (N_1154,N_625,N_671);
nand U1155 (N_1155,N_115,N_152);
nand U1156 (N_1156,N_692,N_22);
or U1157 (N_1157,N_580,N_571);
and U1158 (N_1158,N_259,N_691);
and U1159 (N_1159,N_656,N_26);
nand U1160 (N_1160,N_321,N_642);
nor U1161 (N_1161,N_324,N_648);
and U1162 (N_1162,N_570,N_118);
and U1163 (N_1163,N_224,N_494);
and U1164 (N_1164,N_436,N_52);
nor U1165 (N_1165,N_198,N_726);
xnor U1166 (N_1166,N_629,N_648);
and U1167 (N_1167,N_363,N_723);
xor U1168 (N_1168,N_410,N_589);
nand U1169 (N_1169,N_600,N_30);
nand U1170 (N_1170,N_296,N_15);
or U1171 (N_1171,N_723,N_30);
xnor U1172 (N_1172,N_462,N_560);
and U1173 (N_1173,N_320,N_389);
xnor U1174 (N_1174,N_235,N_681);
nor U1175 (N_1175,N_401,N_623);
nand U1176 (N_1176,N_585,N_691);
xor U1177 (N_1177,N_505,N_497);
or U1178 (N_1178,N_710,N_613);
and U1179 (N_1179,N_573,N_78);
nor U1180 (N_1180,N_707,N_356);
or U1181 (N_1181,N_442,N_226);
xnor U1182 (N_1182,N_273,N_6);
nor U1183 (N_1183,N_199,N_182);
xor U1184 (N_1184,N_694,N_129);
and U1185 (N_1185,N_396,N_297);
nor U1186 (N_1186,N_150,N_5);
and U1187 (N_1187,N_518,N_105);
nand U1188 (N_1188,N_396,N_261);
xor U1189 (N_1189,N_12,N_396);
or U1190 (N_1190,N_340,N_331);
or U1191 (N_1191,N_299,N_523);
or U1192 (N_1192,N_737,N_142);
or U1193 (N_1193,N_196,N_658);
nor U1194 (N_1194,N_664,N_687);
nand U1195 (N_1195,N_279,N_465);
and U1196 (N_1196,N_62,N_726);
and U1197 (N_1197,N_163,N_13);
nand U1198 (N_1198,N_242,N_108);
or U1199 (N_1199,N_215,N_540);
xnor U1200 (N_1200,N_168,N_305);
nand U1201 (N_1201,N_256,N_357);
nand U1202 (N_1202,N_174,N_370);
or U1203 (N_1203,N_719,N_603);
or U1204 (N_1204,N_152,N_153);
and U1205 (N_1205,N_23,N_710);
xor U1206 (N_1206,N_160,N_549);
xnor U1207 (N_1207,N_166,N_55);
and U1208 (N_1208,N_567,N_238);
nor U1209 (N_1209,N_718,N_153);
and U1210 (N_1210,N_370,N_47);
or U1211 (N_1211,N_4,N_142);
nand U1212 (N_1212,N_606,N_642);
or U1213 (N_1213,N_636,N_716);
nand U1214 (N_1214,N_141,N_105);
xnor U1215 (N_1215,N_532,N_324);
xor U1216 (N_1216,N_599,N_529);
nor U1217 (N_1217,N_313,N_257);
or U1218 (N_1218,N_218,N_567);
nand U1219 (N_1219,N_392,N_734);
or U1220 (N_1220,N_274,N_370);
xnor U1221 (N_1221,N_218,N_22);
nand U1222 (N_1222,N_264,N_515);
xor U1223 (N_1223,N_65,N_276);
nor U1224 (N_1224,N_92,N_422);
nand U1225 (N_1225,N_436,N_181);
xor U1226 (N_1226,N_449,N_723);
nor U1227 (N_1227,N_504,N_30);
or U1228 (N_1228,N_5,N_646);
nand U1229 (N_1229,N_631,N_358);
or U1230 (N_1230,N_283,N_193);
nand U1231 (N_1231,N_159,N_594);
or U1232 (N_1232,N_521,N_618);
and U1233 (N_1233,N_334,N_269);
or U1234 (N_1234,N_305,N_518);
xnor U1235 (N_1235,N_243,N_383);
nor U1236 (N_1236,N_634,N_663);
nand U1237 (N_1237,N_566,N_522);
nor U1238 (N_1238,N_225,N_418);
or U1239 (N_1239,N_190,N_79);
and U1240 (N_1240,N_539,N_84);
nor U1241 (N_1241,N_700,N_77);
xor U1242 (N_1242,N_488,N_315);
nand U1243 (N_1243,N_572,N_213);
and U1244 (N_1244,N_67,N_204);
or U1245 (N_1245,N_554,N_71);
or U1246 (N_1246,N_520,N_86);
nor U1247 (N_1247,N_633,N_99);
xor U1248 (N_1248,N_90,N_273);
xnor U1249 (N_1249,N_612,N_319);
and U1250 (N_1250,N_65,N_478);
or U1251 (N_1251,N_125,N_438);
nand U1252 (N_1252,N_339,N_588);
nor U1253 (N_1253,N_343,N_479);
or U1254 (N_1254,N_370,N_291);
or U1255 (N_1255,N_55,N_547);
or U1256 (N_1256,N_265,N_594);
nand U1257 (N_1257,N_524,N_405);
or U1258 (N_1258,N_220,N_670);
nand U1259 (N_1259,N_238,N_462);
xor U1260 (N_1260,N_722,N_213);
nand U1261 (N_1261,N_11,N_542);
and U1262 (N_1262,N_22,N_341);
or U1263 (N_1263,N_76,N_524);
or U1264 (N_1264,N_392,N_443);
nand U1265 (N_1265,N_466,N_697);
nor U1266 (N_1266,N_487,N_35);
or U1267 (N_1267,N_102,N_210);
nand U1268 (N_1268,N_680,N_324);
or U1269 (N_1269,N_118,N_462);
nor U1270 (N_1270,N_648,N_421);
nor U1271 (N_1271,N_169,N_44);
xnor U1272 (N_1272,N_254,N_37);
and U1273 (N_1273,N_142,N_179);
nand U1274 (N_1274,N_133,N_697);
and U1275 (N_1275,N_247,N_706);
and U1276 (N_1276,N_350,N_82);
xor U1277 (N_1277,N_144,N_731);
nand U1278 (N_1278,N_303,N_606);
nor U1279 (N_1279,N_88,N_167);
nand U1280 (N_1280,N_53,N_45);
nor U1281 (N_1281,N_186,N_391);
xnor U1282 (N_1282,N_383,N_634);
and U1283 (N_1283,N_533,N_106);
and U1284 (N_1284,N_61,N_309);
or U1285 (N_1285,N_31,N_505);
nor U1286 (N_1286,N_187,N_726);
nor U1287 (N_1287,N_186,N_419);
nor U1288 (N_1288,N_539,N_643);
xor U1289 (N_1289,N_245,N_642);
xor U1290 (N_1290,N_288,N_355);
nand U1291 (N_1291,N_202,N_90);
xnor U1292 (N_1292,N_520,N_113);
nand U1293 (N_1293,N_103,N_447);
nand U1294 (N_1294,N_456,N_598);
nor U1295 (N_1295,N_147,N_85);
nor U1296 (N_1296,N_122,N_191);
nand U1297 (N_1297,N_34,N_19);
nor U1298 (N_1298,N_223,N_96);
or U1299 (N_1299,N_600,N_569);
nand U1300 (N_1300,N_537,N_156);
nor U1301 (N_1301,N_459,N_655);
or U1302 (N_1302,N_445,N_438);
nor U1303 (N_1303,N_295,N_90);
nor U1304 (N_1304,N_659,N_116);
nand U1305 (N_1305,N_339,N_255);
and U1306 (N_1306,N_3,N_488);
and U1307 (N_1307,N_335,N_681);
or U1308 (N_1308,N_554,N_436);
xnor U1309 (N_1309,N_373,N_62);
nand U1310 (N_1310,N_182,N_488);
nor U1311 (N_1311,N_732,N_562);
or U1312 (N_1312,N_608,N_37);
nor U1313 (N_1313,N_415,N_98);
and U1314 (N_1314,N_339,N_169);
or U1315 (N_1315,N_322,N_239);
xor U1316 (N_1316,N_606,N_567);
and U1317 (N_1317,N_500,N_300);
or U1318 (N_1318,N_330,N_396);
or U1319 (N_1319,N_310,N_468);
or U1320 (N_1320,N_44,N_205);
nor U1321 (N_1321,N_162,N_374);
and U1322 (N_1322,N_462,N_211);
and U1323 (N_1323,N_118,N_101);
xnor U1324 (N_1324,N_689,N_710);
nor U1325 (N_1325,N_24,N_592);
nand U1326 (N_1326,N_512,N_663);
and U1327 (N_1327,N_638,N_605);
xor U1328 (N_1328,N_173,N_62);
nand U1329 (N_1329,N_698,N_79);
nand U1330 (N_1330,N_599,N_494);
nand U1331 (N_1331,N_237,N_253);
xnor U1332 (N_1332,N_116,N_257);
and U1333 (N_1333,N_436,N_561);
xor U1334 (N_1334,N_342,N_266);
or U1335 (N_1335,N_337,N_432);
xnor U1336 (N_1336,N_517,N_239);
and U1337 (N_1337,N_694,N_704);
nor U1338 (N_1338,N_638,N_199);
xnor U1339 (N_1339,N_585,N_480);
xnor U1340 (N_1340,N_622,N_135);
and U1341 (N_1341,N_377,N_176);
and U1342 (N_1342,N_654,N_81);
and U1343 (N_1343,N_364,N_215);
nand U1344 (N_1344,N_46,N_325);
nand U1345 (N_1345,N_302,N_288);
or U1346 (N_1346,N_99,N_314);
or U1347 (N_1347,N_436,N_665);
or U1348 (N_1348,N_174,N_707);
xor U1349 (N_1349,N_85,N_678);
xor U1350 (N_1350,N_488,N_578);
xor U1351 (N_1351,N_396,N_721);
nand U1352 (N_1352,N_37,N_538);
nand U1353 (N_1353,N_223,N_357);
xor U1354 (N_1354,N_233,N_427);
and U1355 (N_1355,N_421,N_30);
or U1356 (N_1356,N_585,N_571);
xor U1357 (N_1357,N_192,N_30);
nand U1358 (N_1358,N_120,N_46);
or U1359 (N_1359,N_55,N_560);
and U1360 (N_1360,N_82,N_44);
or U1361 (N_1361,N_46,N_265);
and U1362 (N_1362,N_463,N_125);
and U1363 (N_1363,N_361,N_467);
xnor U1364 (N_1364,N_307,N_740);
nand U1365 (N_1365,N_28,N_487);
nand U1366 (N_1366,N_672,N_230);
xnor U1367 (N_1367,N_509,N_309);
nand U1368 (N_1368,N_460,N_21);
nand U1369 (N_1369,N_447,N_492);
nor U1370 (N_1370,N_563,N_334);
or U1371 (N_1371,N_555,N_643);
nor U1372 (N_1372,N_280,N_207);
nand U1373 (N_1373,N_455,N_437);
xnor U1374 (N_1374,N_560,N_209);
xnor U1375 (N_1375,N_117,N_525);
nand U1376 (N_1376,N_135,N_337);
nand U1377 (N_1377,N_625,N_253);
nor U1378 (N_1378,N_411,N_603);
xnor U1379 (N_1379,N_674,N_232);
xor U1380 (N_1380,N_746,N_370);
nand U1381 (N_1381,N_313,N_298);
nand U1382 (N_1382,N_456,N_68);
or U1383 (N_1383,N_113,N_363);
and U1384 (N_1384,N_592,N_529);
nand U1385 (N_1385,N_42,N_701);
or U1386 (N_1386,N_416,N_748);
or U1387 (N_1387,N_425,N_666);
nand U1388 (N_1388,N_175,N_65);
nor U1389 (N_1389,N_465,N_623);
nor U1390 (N_1390,N_325,N_464);
or U1391 (N_1391,N_530,N_543);
nor U1392 (N_1392,N_152,N_701);
xnor U1393 (N_1393,N_126,N_363);
and U1394 (N_1394,N_7,N_46);
or U1395 (N_1395,N_411,N_129);
nor U1396 (N_1396,N_735,N_237);
nor U1397 (N_1397,N_33,N_294);
and U1398 (N_1398,N_183,N_546);
nand U1399 (N_1399,N_505,N_709);
and U1400 (N_1400,N_664,N_477);
xnor U1401 (N_1401,N_153,N_117);
and U1402 (N_1402,N_726,N_686);
and U1403 (N_1403,N_27,N_470);
nor U1404 (N_1404,N_309,N_301);
and U1405 (N_1405,N_498,N_359);
or U1406 (N_1406,N_429,N_315);
nand U1407 (N_1407,N_99,N_26);
and U1408 (N_1408,N_140,N_116);
xnor U1409 (N_1409,N_560,N_428);
nand U1410 (N_1410,N_162,N_534);
nand U1411 (N_1411,N_579,N_122);
and U1412 (N_1412,N_709,N_335);
or U1413 (N_1413,N_360,N_354);
or U1414 (N_1414,N_87,N_487);
and U1415 (N_1415,N_434,N_432);
and U1416 (N_1416,N_74,N_212);
nor U1417 (N_1417,N_88,N_264);
xor U1418 (N_1418,N_488,N_613);
nand U1419 (N_1419,N_64,N_148);
xor U1420 (N_1420,N_517,N_654);
nand U1421 (N_1421,N_309,N_262);
nand U1422 (N_1422,N_51,N_318);
nor U1423 (N_1423,N_344,N_375);
or U1424 (N_1424,N_330,N_653);
nor U1425 (N_1425,N_159,N_620);
or U1426 (N_1426,N_48,N_571);
nand U1427 (N_1427,N_706,N_132);
nand U1428 (N_1428,N_730,N_697);
nand U1429 (N_1429,N_391,N_81);
xor U1430 (N_1430,N_457,N_104);
and U1431 (N_1431,N_301,N_683);
nand U1432 (N_1432,N_173,N_189);
or U1433 (N_1433,N_331,N_694);
nand U1434 (N_1434,N_602,N_559);
xnor U1435 (N_1435,N_332,N_136);
xor U1436 (N_1436,N_586,N_448);
and U1437 (N_1437,N_690,N_702);
xor U1438 (N_1438,N_304,N_126);
or U1439 (N_1439,N_344,N_404);
or U1440 (N_1440,N_646,N_485);
nor U1441 (N_1441,N_674,N_505);
nand U1442 (N_1442,N_477,N_186);
xor U1443 (N_1443,N_320,N_319);
and U1444 (N_1444,N_408,N_345);
xnor U1445 (N_1445,N_321,N_648);
nand U1446 (N_1446,N_361,N_117);
nor U1447 (N_1447,N_202,N_745);
and U1448 (N_1448,N_661,N_196);
nor U1449 (N_1449,N_522,N_691);
nor U1450 (N_1450,N_533,N_118);
and U1451 (N_1451,N_260,N_708);
xor U1452 (N_1452,N_149,N_460);
and U1453 (N_1453,N_717,N_410);
nor U1454 (N_1454,N_460,N_737);
nor U1455 (N_1455,N_141,N_738);
and U1456 (N_1456,N_532,N_442);
and U1457 (N_1457,N_670,N_678);
xnor U1458 (N_1458,N_88,N_62);
or U1459 (N_1459,N_456,N_207);
nor U1460 (N_1460,N_325,N_288);
nand U1461 (N_1461,N_24,N_643);
nand U1462 (N_1462,N_266,N_264);
nor U1463 (N_1463,N_336,N_160);
nor U1464 (N_1464,N_108,N_475);
nor U1465 (N_1465,N_9,N_0);
xnor U1466 (N_1466,N_507,N_82);
nand U1467 (N_1467,N_562,N_156);
nor U1468 (N_1468,N_88,N_202);
or U1469 (N_1469,N_222,N_278);
or U1470 (N_1470,N_417,N_319);
nor U1471 (N_1471,N_546,N_685);
or U1472 (N_1472,N_589,N_556);
nand U1473 (N_1473,N_718,N_407);
and U1474 (N_1474,N_364,N_139);
nor U1475 (N_1475,N_360,N_398);
or U1476 (N_1476,N_309,N_599);
nand U1477 (N_1477,N_99,N_572);
and U1478 (N_1478,N_95,N_147);
nand U1479 (N_1479,N_401,N_302);
and U1480 (N_1480,N_309,N_464);
and U1481 (N_1481,N_564,N_456);
or U1482 (N_1482,N_399,N_678);
and U1483 (N_1483,N_44,N_203);
nand U1484 (N_1484,N_222,N_257);
and U1485 (N_1485,N_510,N_627);
or U1486 (N_1486,N_443,N_222);
or U1487 (N_1487,N_130,N_419);
xor U1488 (N_1488,N_721,N_361);
nor U1489 (N_1489,N_372,N_496);
nor U1490 (N_1490,N_259,N_126);
and U1491 (N_1491,N_203,N_63);
and U1492 (N_1492,N_656,N_709);
nand U1493 (N_1493,N_545,N_739);
or U1494 (N_1494,N_233,N_660);
nand U1495 (N_1495,N_577,N_32);
and U1496 (N_1496,N_595,N_207);
nor U1497 (N_1497,N_258,N_119);
and U1498 (N_1498,N_489,N_178);
or U1499 (N_1499,N_123,N_621);
xnor U1500 (N_1500,N_973,N_1058);
and U1501 (N_1501,N_1015,N_978);
and U1502 (N_1502,N_1399,N_1413);
or U1503 (N_1503,N_1451,N_1461);
xnor U1504 (N_1504,N_1245,N_870);
or U1505 (N_1505,N_1377,N_1119);
and U1506 (N_1506,N_876,N_1427);
and U1507 (N_1507,N_948,N_1246);
or U1508 (N_1508,N_1044,N_1491);
or U1509 (N_1509,N_842,N_752);
nand U1510 (N_1510,N_1325,N_1169);
or U1511 (N_1511,N_883,N_1237);
nor U1512 (N_1512,N_985,N_1443);
or U1513 (N_1513,N_1390,N_925);
and U1514 (N_1514,N_972,N_1046);
nor U1515 (N_1515,N_1032,N_1197);
nand U1516 (N_1516,N_951,N_926);
nand U1517 (N_1517,N_1388,N_924);
nand U1518 (N_1518,N_846,N_1161);
nand U1519 (N_1519,N_817,N_778);
or U1520 (N_1520,N_1230,N_788);
xor U1521 (N_1521,N_1269,N_920);
and U1522 (N_1522,N_1051,N_1167);
nand U1523 (N_1523,N_1407,N_1344);
or U1524 (N_1524,N_851,N_881);
nand U1525 (N_1525,N_1057,N_1188);
xor U1526 (N_1526,N_879,N_783);
nand U1527 (N_1527,N_1153,N_1128);
xnor U1528 (N_1528,N_1067,N_1482);
xor U1529 (N_1529,N_1373,N_790);
and U1530 (N_1530,N_1265,N_1484);
and U1531 (N_1531,N_910,N_998);
xor U1532 (N_1532,N_884,N_963);
nand U1533 (N_1533,N_1165,N_1178);
xor U1534 (N_1534,N_761,N_1066);
xor U1535 (N_1535,N_1437,N_889);
nand U1536 (N_1536,N_1329,N_933);
and U1537 (N_1537,N_869,N_1412);
nor U1538 (N_1538,N_1406,N_1037);
and U1539 (N_1539,N_1025,N_1072);
nand U1540 (N_1540,N_1334,N_1022);
nand U1541 (N_1541,N_1054,N_1131);
xor U1542 (N_1542,N_1438,N_1419);
xnor U1543 (N_1543,N_1376,N_912);
nand U1544 (N_1544,N_1220,N_862);
xor U1545 (N_1545,N_1240,N_1367);
and U1546 (N_1546,N_750,N_832);
or U1547 (N_1547,N_1450,N_1366);
or U1548 (N_1548,N_1073,N_1341);
nor U1549 (N_1549,N_1086,N_1403);
nor U1550 (N_1550,N_1241,N_999);
nor U1551 (N_1551,N_1053,N_809);
or U1552 (N_1552,N_882,N_766);
nand U1553 (N_1553,N_988,N_1079);
and U1554 (N_1554,N_1127,N_1000);
nand U1555 (N_1555,N_1260,N_1418);
or U1556 (N_1556,N_1088,N_1476);
nor U1557 (N_1557,N_1436,N_1183);
nor U1558 (N_1558,N_1486,N_930);
and U1559 (N_1559,N_1300,N_1034);
or U1560 (N_1560,N_1007,N_1288);
xor U1561 (N_1561,N_1179,N_1322);
and U1562 (N_1562,N_1468,N_1039);
and U1563 (N_1563,N_798,N_772);
and U1564 (N_1564,N_855,N_854);
xor U1565 (N_1565,N_949,N_1487);
nor U1566 (N_1566,N_980,N_1004);
or U1567 (N_1567,N_1055,N_1361);
xor U1568 (N_1568,N_825,N_1247);
nor U1569 (N_1569,N_1157,N_1394);
nand U1570 (N_1570,N_865,N_1492);
nor U1571 (N_1571,N_1281,N_1229);
or U1572 (N_1572,N_1035,N_867);
nand U1573 (N_1573,N_1218,N_990);
nor U1574 (N_1574,N_1173,N_1184);
nor U1575 (N_1575,N_1099,N_1424);
or U1576 (N_1576,N_1094,N_1404);
xnor U1577 (N_1577,N_1308,N_943);
and U1578 (N_1578,N_1107,N_1452);
nand U1579 (N_1579,N_757,N_1429);
nor U1580 (N_1580,N_1190,N_1315);
or U1581 (N_1581,N_782,N_1417);
xor U1582 (N_1582,N_1239,N_1499);
and U1583 (N_1583,N_1462,N_1122);
xor U1584 (N_1584,N_1309,N_962);
xnor U1585 (N_1585,N_1393,N_1435);
xnor U1586 (N_1586,N_952,N_1112);
or U1587 (N_1587,N_903,N_1392);
xor U1588 (N_1588,N_1222,N_1148);
xor U1589 (N_1589,N_1110,N_1162);
nand U1590 (N_1590,N_1209,N_1456);
and U1591 (N_1591,N_987,N_1180);
and U1592 (N_1592,N_1370,N_983);
or U1593 (N_1593,N_848,N_1048);
xnor U1594 (N_1594,N_1142,N_921);
or U1595 (N_1595,N_1196,N_1194);
nor U1596 (N_1596,N_1001,N_1335);
and U1597 (N_1597,N_800,N_845);
nor U1598 (N_1598,N_833,N_1149);
xor U1599 (N_1599,N_1002,N_1172);
nor U1600 (N_1600,N_1278,N_1011);
xor U1601 (N_1601,N_1279,N_1242);
and U1602 (N_1602,N_1307,N_1075);
nor U1603 (N_1603,N_822,N_1310);
xnor U1604 (N_1604,N_1356,N_1323);
and U1605 (N_1605,N_1158,N_1005);
nand U1606 (N_1606,N_816,N_1089);
and U1607 (N_1607,N_939,N_1474);
nor U1608 (N_1608,N_1297,N_1291);
and U1609 (N_1609,N_1358,N_756);
xor U1610 (N_1610,N_1012,N_878);
nor U1611 (N_1611,N_1017,N_1340);
and U1612 (N_1612,N_944,N_902);
or U1613 (N_1613,N_1111,N_784);
nand U1614 (N_1614,N_1466,N_866);
xnor U1615 (N_1615,N_1430,N_1449);
or U1616 (N_1616,N_1401,N_986);
or U1617 (N_1617,N_1217,N_1263);
nand U1618 (N_1618,N_1347,N_781);
or U1619 (N_1619,N_1043,N_1441);
and U1620 (N_1620,N_1348,N_754);
nand U1621 (N_1621,N_1493,N_1159);
and U1622 (N_1622,N_1185,N_852);
nand U1623 (N_1623,N_994,N_1250);
and U1624 (N_1624,N_1285,N_828);
nor U1625 (N_1625,N_1116,N_1052);
nand U1626 (N_1626,N_931,N_1305);
xor U1627 (N_1627,N_1331,N_1191);
xnor U1628 (N_1628,N_1258,N_1163);
xor U1629 (N_1629,N_1410,N_1069);
nor U1630 (N_1630,N_1349,N_1207);
and U1631 (N_1631,N_896,N_1372);
nand U1632 (N_1632,N_830,N_858);
xor U1633 (N_1633,N_915,N_810);
and U1634 (N_1634,N_1092,N_1343);
nor U1635 (N_1635,N_1455,N_1087);
xor U1636 (N_1636,N_1354,N_1375);
and U1637 (N_1637,N_806,N_975);
nand U1638 (N_1638,N_1405,N_1342);
or U1639 (N_1639,N_981,N_1221);
nand U1640 (N_1640,N_1262,N_914);
or U1641 (N_1641,N_820,N_839);
xnor U1642 (N_1642,N_906,N_1383);
nor U1643 (N_1643,N_1074,N_787);
nand U1644 (N_1644,N_1371,N_803);
xnor U1645 (N_1645,N_1319,N_1332);
xnor U1646 (N_1646,N_1336,N_1444);
nor U1647 (N_1647,N_1447,N_1226);
nand U1648 (N_1648,N_843,N_1176);
and U1649 (N_1649,N_1299,N_769);
nor U1650 (N_1650,N_1369,N_1238);
nor U1651 (N_1651,N_946,N_970);
and U1652 (N_1652,N_1359,N_1078);
nand U1653 (N_1653,N_1432,N_829);
xnor U1654 (N_1654,N_1013,N_1495);
or U1655 (N_1655,N_1140,N_1350);
or U1656 (N_1656,N_1214,N_909);
xor U1657 (N_1657,N_1024,N_1268);
and U1658 (N_1658,N_950,N_1193);
nand U1659 (N_1659,N_908,N_1030);
nor U1660 (N_1660,N_1266,N_1314);
nand U1661 (N_1661,N_877,N_916);
nor U1662 (N_1662,N_1120,N_1085);
nor U1663 (N_1663,N_1275,N_857);
nor U1664 (N_1664,N_1264,N_1204);
nand U1665 (N_1665,N_1113,N_823);
xnor U1666 (N_1666,N_1151,N_936);
nor U1667 (N_1667,N_890,N_947);
nand U1668 (N_1668,N_1497,N_997);
or U1669 (N_1669,N_1227,N_1216);
nor U1670 (N_1670,N_1494,N_838);
xnor U1671 (N_1671,N_1253,N_1132);
and U1672 (N_1672,N_753,N_791);
or U1673 (N_1673,N_1312,N_1199);
or U1674 (N_1674,N_1133,N_1306);
nor U1675 (N_1675,N_1473,N_1063);
nor U1676 (N_1676,N_1355,N_1465);
xnor U1677 (N_1677,N_1421,N_1286);
nor U1678 (N_1678,N_841,N_1463);
xnor U1679 (N_1679,N_969,N_901);
or U1680 (N_1680,N_1397,N_875);
or U1681 (N_1681,N_1177,N_1283);
nand U1682 (N_1682,N_1289,N_1065);
and U1683 (N_1683,N_1431,N_955);
nor U1684 (N_1684,N_1198,N_868);
and U1685 (N_1685,N_1382,N_1234);
nor U1686 (N_1686,N_1061,N_1248);
nor U1687 (N_1687,N_1125,N_1206);
and U1688 (N_1688,N_1175,N_1105);
and U1689 (N_1689,N_898,N_1321);
and U1690 (N_1690,N_1235,N_1021);
and U1691 (N_1691,N_1498,N_953);
nor U1692 (N_1692,N_923,N_904);
and U1693 (N_1693,N_1143,N_850);
or U1694 (N_1694,N_1439,N_1181);
xor U1695 (N_1695,N_1064,N_1302);
and U1696 (N_1696,N_1118,N_1475);
and U1697 (N_1697,N_1244,N_1422);
xor U1698 (N_1698,N_780,N_1490);
nand U1699 (N_1699,N_815,N_1280);
xor U1700 (N_1700,N_957,N_913);
nor U1701 (N_1701,N_1135,N_1201);
nand U1702 (N_1702,N_1047,N_938);
nand U1703 (N_1703,N_805,N_1464);
or U1704 (N_1704,N_1313,N_1212);
xor U1705 (N_1705,N_1378,N_1324);
and U1706 (N_1706,N_1357,N_1290);
or U1707 (N_1707,N_1036,N_1311);
and U1708 (N_1708,N_1130,N_1480);
xor U1709 (N_1709,N_1211,N_1284);
or U1710 (N_1710,N_1006,N_1136);
nor U1711 (N_1711,N_1028,N_1428);
nand U1712 (N_1712,N_812,N_860);
and U1713 (N_1713,N_1170,N_1445);
or U1714 (N_1714,N_1433,N_1470);
nor U1715 (N_1715,N_827,N_1203);
and U1716 (N_1716,N_807,N_1338);
or U1717 (N_1717,N_1081,N_945);
and U1718 (N_1718,N_977,N_1472);
and U1719 (N_1719,N_1020,N_1328);
or U1720 (N_1720,N_1317,N_1381);
or U1721 (N_1721,N_1337,N_993);
xor U1722 (N_1722,N_966,N_1147);
or U1723 (N_1723,N_834,N_961);
and U1724 (N_1724,N_1009,N_1156);
or U1725 (N_1725,N_1489,N_861);
or U1726 (N_1726,N_1384,N_1330);
or U1727 (N_1727,N_1144,N_1385);
nand U1728 (N_1728,N_1353,N_1208);
and U1729 (N_1729,N_777,N_1224);
nand U1730 (N_1730,N_864,N_1272);
nor U1731 (N_1731,N_1071,N_1182);
nand U1732 (N_1732,N_849,N_1060);
xor U1733 (N_1733,N_774,N_992);
nor U1734 (N_1734,N_1287,N_1326);
xnor U1735 (N_1735,N_1213,N_1010);
or U1736 (N_1736,N_1123,N_1346);
nand U1737 (N_1737,N_1440,N_1045);
nand U1738 (N_1738,N_1134,N_1301);
nor U1739 (N_1739,N_856,N_1068);
nor U1740 (N_1740,N_1483,N_871);
nand U1741 (N_1741,N_818,N_1114);
nor U1742 (N_1742,N_1379,N_1104);
or U1743 (N_1743,N_794,N_785);
nor U1744 (N_1744,N_1189,N_954);
and U1745 (N_1745,N_1256,N_1496);
xor U1746 (N_1746,N_928,N_853);
nand U1747 (N_1747,N_1254,N_991);
or U1748 (N_1748,N_1391,N_888);
or U1749 (N_1749,N_1205,N_895);
and U1750 (N_1750,N_797,N_960);
nand U1751 (N_1751,N_1100,N_1408);
xnor U1752 (N_1752,N_897,N_932);
nor U1753 (N_1753,N_899,N_1202);
nand U1754 (N_1754,N_976,N_1049);
nor U1755 (N_1755,N_762,N_1457);
xnor U1756 (N_1756,N_1479,N_1080);
and U1757 (N_1757,N_1031,N_979);
or U1758 (N_1758,N_1270,N_1387);
xor U1759 (N_1759,N_1296,N_1426);
xnor U1760 (N_1760,N_984,N_894);
nand U1761 (N_1761,N_887,N_821);
and U1762 (N_1762,N_1327,N_1228);
or U1763 (N_1763,N_1467,N_1187);
xnor U1764 (N_1764,N_824,N_1292);
nand U1765 (N_1765,N_802,N_1316);
or U1766 (N_1766,N_1477,N_1362);
nand U1767 (N_1767,N_1026,N_911);
or U1768 (N_1768,N_1333,N_789);
nor U1769 (N_1769,N_768,N_1084);
xnor U1770 (N_1770,N_1014,N_1223);
nand U1771 (N_1771,N_974,N_1124);
nor U1772 (N_1772,N_919,N_1374);
and U1773 (N_1773,N_1033,N_837);
or U1774 (N_1774,N_1303,N_826);
and U1775 (N_1775,N_1298,N_760);
xor U1776 (N_1776,N_1339,N_840);
or U1777 (N_1777,N_917,N_886);
xnor U1778 (N_1778,N_942,N_1027);
nand U1779 (N_1779,N_1137,N_1093);
or U1780 (N_1780,N_965,N_1231);
nor U1781 (N_1781,N_1411,N_1236);
nor U1782 (N_1782,N_1360,N_1101);
or U1783 (N_1783,N_1138,N_795);
nor U1784 (N_1784,N_1402,N_1282);
or U1785 (N_1785,N_1059,N_1488);
and U1786 (N_1786,N_1090,N_775);
or U1787 (N_1787,N_922,N_940);
xor U1788 (N_1788,N_1146,N_1117);
or U1789 (N_1789,N_937,N_1155);
or U1790 (N_1790,N_1019,N_1050);
nor U1791 (N_1791,N_773,N_1023);
nand U1792 (N_1792,N_1109,N_801);
xor U1793 (N_1793,N_1446,N_771);
nor U1794 (N_1794,N_1160,N_1215);
and U1795 (N_1795,N_1448,N_1164);
nor U1796 (N_1796,N_1380,N_880);
or U1797 (N_1797,N_1274,N_907);
or U1798 (N_1798,N_799,N_764);
nand U1799 (N_1799,N_893,N_964);
and U1800 (N_1800,N_1108,N_836);
nand U1801 (N_1801,N_819,N_765);
nor U1802 (N_1802,N_763,N_941);
nor U1803 (N_1803,N_1442,N_1293);
nor U1804 (N_1804,N_905,N_996);
xnor U1805 (N_1805,N_1168,N_835);
and U1806 (N_1806,N_967,N_1386);
and U1807 (N_1807,N_1096,N_1273);
nand U1808 (N_1808,N_1232,N_1416);
and U1809 (N_1809,N_935,N_1166);
and U1810 (N_1810,N_751,N_968);
and U1811 (N_1811,N_1318,N_1038);
nand U1812 (N_1812,N_1460,N_755);
and U1813 (N_1813,N_1018,N_1016);
and U1814 (N_1814,N_1454,N_1368);
or U1815 (N_1815,N_1083,N_1364);
nor U1816 (N_1816,N_786,N_1106);
and U1817 (N_1817,N_1103,N_1481);
nand U1818 (N_1818,N_1252,N_776);
or U1819 (N_1819,N_1095,N_767);
nand U1820 (N_1820,N_959,N_982);
or U1821 (N_1821,N_1415,N_1192);
and U1822 (N_1822,N_1070,N_1139);
and U1823 (N_1823,N_1056,N_995);
xor U1824 (N_1824,N_793,N_779);
or U1825 (N_1825,N_1225,N_1423);
nand U1826 (N_1826,N_1459,N_844);
nor U1827 (N_1827,N_1171,N_1097);
nor U1828 (N_1828,N_1150,N_1008);
or U1829 (N_1829,N_1102,N_900);
nand U1830 (N_1830,N_918,N_831);
and U1831 (N_1831,N_1082,N_1098);
nand U1832 (N_1832,N_1062,N_873);
or U1833 (N_1833,N_1294,N_1469);
nor U1834 (N_1834,N_1115,N_1261);
nand U1835 (N_1835,N_1414,N_1257);
nor U1836 (N_1836,N_804,N_1091);
nor U1837 (N_1837,N_1271,N_1409);
nand U1838 (N_1838,N_1210,N_758);
nor U1839 (N_1839,N_929,N_1365);
nand U1840 (N_1840,N_1154,N_1458);
nor U1841 (N_1841,N_927,N_1145);
xor U1842 (N_1842,N_1453,N_1295);
xnor U1843 (N_1843,N_770,N_1152);
nand U1844 (N_1844,N_1277,N_1121);
or U1845 (N_1845,N_1320,N_1041);
or U1846 (N_1846,N_874,N_971);
xor U1847 (N_1847,N_1255,N_1396);
xnor U1848 (N_1848,N_891,N_1485);
xor U1849 (N_1849,N_792,N_1077);
or U1850 (N_1850,N_1400,N_1126);
or U1851 (N_1851,N_814,N_1040);
or U1852 (N_1852,N_1141,N_863);
nand U1853 (N_1853,N_1389,N_847);
xor U1854 (N_1854,N_1425,N_1200);
or U1855 (N_1855,N_1304,N_1249);
or U1856 (N_1856,N_892,N_1233);
and U1857 (N_1857,N_1129,N_859);
xor U1858 (N_1858,N_811,N_1395);
xor U1859 (N_1859,N_813,N_759);
nor U1860 (N_1860,N_1478,N_1076);
nand U1861 (N_1861,N_872,N_1351);
and U1862 (N_1862,N_796,N_1251);
nand U1863 (N_1863,N_1259,N_1029);
xnor U1864 (N_1864,N_956,N_1042);
xnor U1865 (N_1865,N_1471,N_808);
and U1866 (N_1866,N_1003,N_1276);
and U1867 (N_1867,N_1267,N_1243);
or U1868 (N_1868,N_885,N_989);
nand U1869 (N_1869,N_1174,N_1195);
xnor U1870 (N_1870,N_934,N_1345);
and U1871 (N_1871,N_1352,N_1420);
and U1872 (N_1872,N_1434,N_1219);
nand U1873 (N_1873,N_1363,N_1398);
or U1874 (N_1874,N_958,N_1186);
nor U1875 (N_1875,N_1349,N_783);
nand U1876 (N_1876,N_844,N_943);
or U1877 (N_1877,N_1103,N_1345);
or U1878 (N_1878,N_1416,N_844);
or U1879 (N_1879,N_1188,N_1123);
and U1880 (N_1880,N_786,N_1148);
nand U1881 (N_1881,N_759,N_786);
xnor U1882 (N_1882,N_1369,N_911);
nor U1883 (N_1883,N_1431,N_1488);
nor U1884 (N_1884,N_1213,N_1269);
nand U1885 (N_1885,N_1417,N_922);
and U1886 (N_1886,N_1355,N_1289);
xor U1887 (N_1887,N_855,N_760);
xor U1888 (N_1888,N_1420,N_1229);
xnor U1889 (N_1889,N_949,N_1239);
nand U1890 (N_1890,N_757,N_907);
and U1891 (N_1891,N_1056,N_906);
nor U1892 (N_1892,N_829,N_950);
nor U1893 (N_1893,N_1032,N_1352);
nand U1894 (N_1894,N_1155,N_1144);
xor U1895 (N_1895,N_1496,N_1143);
nand U1896 (N_1896,N_1324,N_811);
xnor U1897 (N_1897,N_928,N_1366);
and U1898 (N_1898,N_1190,N_1499);
nand U1899 (N_1899,N_799,N_1068);
and U1900 (N_1900,N_832,N_1394);
nor U1901 (N_1901,N_829,N_1062);
nor U1902 (N_1902,N_1218,N_1216);
xor U1903 (N_1903,N_1263,N_1151);
or U1904 (N_1904,N_1303,N_1476);
xor U1905 (N_1905,N_895,N_1101);
xor U1906 (N_1906,N_1083,N_1395);
or U1907 (N_1907,N_1160,N_802);
xor U1908 (N_1908,N_1201,N_1436);
and U1909 (N_1909,N_1435,N_1427);
nor U1910 (N_1910,N_895,N_1290);
or U1911 (N_1911,N_777,N_1434);
xor U1912 (N_1912,N_1008,N_1436);
and U1913 (N_1913,N_1088,N_1104);
or U1914 (N_1914,N_1486,N_1002);
and U1915 (N_1915,N_1407,N_789);
xor U1916 (N_1916,N_1465,N_797);
xnor U1917 (N_1917,N_934,N_1298);
nor U1918 (N_1918,N_890,N_1370);
nor U1919 (N_1919,N_1114,N_954);
xor U1920 (N_1920,N_1035,N_783);
and U1921 (N_1921,N_819,N_1457);
and U1922 (N_1922,N_1203,N_1392);
nor U1923 (N_1923,N_915,N_1056);
nor U1924 (N_1924,N_1332,N_1103);
nand U1925 (N_1925,N_762,N_969);
nand U1926 (N_1926,N_1445,N_1173);
and U1927 (N_1927,N_962,N_1316);
nor U1928 (N_1928,N_1079,N_1427);
xnor U1929 (N_1929,N_1290,N_1242);
nor U1930 (N_1930,N_1267,N_1381);
and U1931 (N_1931,N_1004,N_1045);
and U1932 (N_1932,N_1335,N_1445);
nand U1933 (N_1933,N_1076,N_757);
and U1934 (N_1934,N_1146,N_1211);
and U1935 (N_1935,N_1153,N_1060);
and U1936 (N_1936,N_1293,N_1341);
nand U1937 (N_1937,N_1463,N_1112);
nand U1938 (N_1938,N_917,N_1263);
nor U1939 (N_1939,N_794,N_900);
xnor U1940 (N_1940,N_1333,N_1228);
and U1941 (N_1941,N_878,N_853);
or U1942 (N_1942,N_1491,N_878);
and U1943 (N_1943,N_1471,N_885);
and U1944 (N_1944,N_1258,N_793);
nand U1945 (N_1945,N_857,N_924);
nor U1946 (N_1946,N_1107,N_922);
nor U1947 (N_1947,N_824,N_1416);
nor U1948 (N_1948,N_984,N_878);
xnor U1949 (N_1949,N_1175,N_1417);
nand U1950 (N_1950,N_1014,N_1361);
xor U1951 (N_1951,N_882,N_860);
and U1952 (N_1952,N_1057,N_1458);
nor U1953 (N_1953,N_1115,N_1220);
and U1954 (N_1954,N_961,N_1161);
nor U1955 (N_1955,N_1117,N_1256);
xnor U1956 (N_1956,N_1131,N_1342);
nand U1957 (N_1957,N_1000,N_1095);
xnor U1958 (N_1958,N_1019,N_1188);
or U1959 (N_1959,N_1039,N_1322);
xnor U1960 (N_1960,N_1299,N_1201);
and U1961 (N_1961,N_1373,N_850);
nor U1962 (N_1962,N_821,N_1363);
or U1963 (N_1963,N_1250,N_1344);
and U1964 (N_1964,N_1474,N_1401);
nand U1965 (N_1965,N_1351,N_1488);
or U1966 (N_1966,N_1391,N_864);
nor U1967 (N_1967,N_1137,N_940);
or U1968 (N_1968,N_1203,N_1369);
or U1969 (N_1969,N_1332,N_758);
nand U1970 (N_1970,N_908,N_772);
xnor U1971 (N_1971,N_936,N_1325);
and U1972 (N_1972,N_756,N_830);
xor U1973 (N_1973,N_1200,N_1482);
and U1974 (N_1974,N_1332,N_1169);
or U1975 (N_1975,N_1343,N_898);
xnor U1976 (N_1976,N_1420,N_1468);
nand U1977 (N_1977,N_1082,N_761);
nand U1978 (N_1978,N_809,N_1158);
and U1979 (N_1979,N_767,N_1499);
nor U1980 (N_1980,N_1371,N_1228);
and U1981 (N_1981,N_885,N_1050);
nand U1982 (N_1982,N_836,N_1206);
nand U1983 (N_1983,N_1494,N_1381);
nand U1984 (N_1984,N_1331,N_970);
xnor U1985 (N_1985,N_936,N_1197);
nor U1986 (N_1986,N_1457,N_975);
and U1987 (N_1987,N_1110,N_834);
nand U1988 (N_1988,N_1444,N_1174);
nand U1989 (N_1989,N_1192,N_771);
or U1990 (N_1990,N_1377,N_957);
and U1991 (N_1991,N_916,N_1115);
nand U1992 (N_1992,N_936,N_1490);
xor U1993 (N_1993,N_1440,N_1488);
xnor U1994 (N_1994,N_1012,N_767);
nor U1995 (N_1995,N_1112,N_1314);
nand U1996 (N_1996,N_1019,N_1220);
and U1997 (N_1997,N_1042,N_1448);
xor U1998 (N_1998,N_1324,N_1485);
nand U1999 (N_1999,N_815,N_845);
nand U2000 (N_2000,N_1196,N_1148);
nand U2001 (N_2001,N_1187,N_1350);
or U2002 (N_2002,N_1481,N_1230);
nand U2003 (N_2003,N_1015,N_869);
nor U2004 (N_2004,N_1081,N_1131);
or U2005 (N_2005,N_1123,N_890);
or U2006 (N_2006,N_1131,N_885);
or U2007 (N_2007,N_849,N_1130);
nand U2008 (N_2008,N_1258,N_1370);
nor U2009 (N_2009,N_874,N_1060);
nor U2010 (N_2010,N_878,N_775);
or U2011 (N_2011,N_1403,N_1388);
and U2012 (N_2012,N_872,N_1169);
or U2013 (N_2013,N_1306,N_1430);
xnor U2014 (N_2014,N_1017,N_987);
or U2015 (N_2015,N_951,N_811);
xnor U2016 (N_2016,N_1112,N_949);
nand U2017 (N_2017,N_1167,N_1436);
or U2018 (N_2018,N_1188,N_1141);
nor U2019 (N_2019,N_1494,N_793);
or U2020 (N_2020,N_1039,N_1304);
or U2021 (N_2021,N_1157,N_1149);
and U2022 (N_2022,N_1035,N_1013);
and U2023 (N_2023,N_1433,N_1008);
and U2024 (N_2024,N_1237,N_1375);
nand U2025 (N_2025,N_1115,N_827);
nor U2026 (N_2026,N_931,N_814);
and U2027 (N_2027,N_1172,N_1481);
nand U2028 (N_2028,N_1308,N_1146);
nand U2029 (N_2029,N_1192,N_824);
nand U2030 (N_2030,N_1451,N_864);
and U2031 (N_2031,N_1012,N_959);
nand U2032 (N_2032,N_782,N_1469);
xnor U2033 (N_2033,N_1274,N_1049);
or U2034 (N_2034,N_753,N_1295);
or U2035 (N_2035,N_1473,N_935);
xor U2036 (N_2036,N_1046,N_1481);
and U2037 (N_2037,N_912,N_938);
nand U2038 (N_2038,N_988,N_1212);
nor U2039 (N_2039,N_995,N_965);
nor U2040 (N_2040,N_1069,N_1341);
xor U2041 (N_2041,N_1010,N_1050);
or U2042 (N_2042,N_1364,N_1168);
and U2043 (N_2043,N_1180,N_1357);
nand U2044 (N_2044,N_1005,N_894);
xnor U2045 (N_2045,N_1439,N_1399);
nand U2046 (N_2046,N_1196,N_1269);
and U2047 (N_2047,N_1143,N_907);
and U2048 (N_2048,N_802,N_1034);
and U2049 (N_2049,N_1076,N_840);
and U2050 (N_2050,N_1483,N_837);
or U2051 (N_2051,N_850,N_754);
nand U2052 (N_2052,N_1421,N_751);
or U2053 (N_2053,N_884,N_1464);
and U2054 (N_2054,N_1331,N_1312);
xor U2055 (N_2055,N_997,N_1040);
nand U2056 (N_2056,N_1301,N_831);
nand U2057 (N_2057,N_903,N_823);
nor U2058 (N_2058,N_969,N_804);
xor U2059 (N_2059,N_1208,N_850);
and U2060 (N_2060,N_1124,N_982);
and U2061 (N_2061,N_1456,N_1034);
nand U2062 (N_2062,N_999,N_1385);
nand U2063 (N_2063,N_1395,N_1153);
nand U2064 (N_2064,N_1188,N_751);
nor U2065 (N_2065,N_1127,N_863);
nor U2066 (N_2066,N_811,N_1022);
and U2067 (N_2067,N_1245,N_769);
and U2068 (N_2068,N_1235,N_1264);
nand U2069 (N_2069,N_1064,N_1230);
xnor U2070 (N_2070,N_1178,N_1466);
and U2071 (N_2071,N_1259,N_1217);
xnor U2072 (N_2072,N_1102,N_1140);
or U2073 (N_2073,N_808,N_1236);
nor U2074 (N_2074,N_1072,N_1094);
nand U2075 (N_2075,N_1046,N_905);
or U2076 (N_2076,N_1081,N_1041);
and U2077 (N_2077,N_839,N_1374);
nand U2078 (N_2078,N_1490,N_938);
and U2079 (N_2079,N_1019,N_1189);
and U2080 (N_2080,N_1277,N_821);
and U2081 (N_2081,N_1453,N_1090);
xor U2082 (N_2082,N_1328,N_1330);
nand U2083 (N_2083,N_856,N_1114);
and U2084 (N_2084,N_799,N_1048);
and U2085 (N_2085,N_1442,N_796);
or U2086 (N_2086,N_1177,N_1227);
and U2087 (N_2087,N_1173,N_1345);
or U2088 (N_2088,N_805,N_1229);
nor U2089 (N_2089,N_1460,N_1364);
and U2090 (N_2090,N_847,N_1469);
nor U2091 (N_2091,N_1130,N_1443);
and U2092 (N_2092,N_1304,N_900);
xnor U2093 (N_2093,N_953,N_832);
and U2094 (N_2094,N_1294,N_1086);
or U2095 (N_2095,N_1300,N_888);
nand U2096 (N_2096,N_1343,N_972);
xnor U2097 (N_2097,N_1201,N_1466);
and U2098 (N_2098,N_1143,N_1345);
xnor U2099 (N_2099,N_1405,N_1073);
xnor U2100 (N_2100,N_1100,N_1006);
nor U2101 (N_2101,N_1005,N_1400);
nor U2102 (N_2102,N_1425,N_896);
and U2103 (N_2103,N_805,N_1481);
and U2104 (N_2104,N_1014,N_901);
nand U2105 (N_2105,N_1244,N_819);
or U2106 (N_2106,N_1216,N_790);
nor U2107 (N_2107,N_1290,N_990);
and U2108 (N_2108,N_762,N_1137);
or U2109 (N_2109,N_863,N_1134);
nand U2110 (N_2110,N_1201,N_1048);
xnor U2111 (N_2111,N_1487,N_960);
and U2112 (N_2112,N_805,N_786);
nand U2113 (N_2113,N_840,N_1190);
and U2114 (N_2114,N_793,N_803);
and U2115 (N_2115,N_1393,N_757);
or U2116 (N_2116,N_1133,N_991);
and U2117 (N_2117,N_851,N_803);
xor U2118 (N_2118,N_828,N_1290);
nor U2119 (N_2119,N_982,N_812);
nand U2120 (N_2120,N_1478,N_1452);
xor U2121 (N_2121,N_1215,N_1201);
or U2122 (N_2122,N_1461,N_1285);
or U2123 (N_2123,N_951,N_857);
xor U2124 (N_2124,N_1038,N_765);
nand U2125 (N_2125,N_1077,N_909);
nor U2126 (N_2126,N_1195,N_1053);
xor U2127 (N_2127,N_1123,N_947);
nor U2128 (N_2128,N_975,N_1373);
xnor U2129 (N_2129,N_795,N_1404);
and U2130 (N_2130,N_1109,N_1173);
or U2131 (N_2131,N_1212,N_1420);
and U2132 (N_2132,N_1357,N_1080);
and U2133 (N_2133,N_1365,N_866);
nand U2134 (N_2134,N_851,N_1087);
nand U2135 (N_2135,N_1055,N_890);
and U2136 (N_2136,N_982,N_1061);
or U2137 (N_2137,N_1459,N_930);
and U2138 (N_2138,N_1426,N_930);
xnor U2139 (N_2139,N_1047,N_1439);
nand U2140 (N_2140,N_1089,N_1060);
or U2141 (N_2141,N_1300,N_1007);
or U2142 (N_2142,N_1237,N_878);
xnor U2143 (N_2143,N_1220,N_1067);
and U2144 (N_2144,N_1440,N_1448);
or U2145 (N_2145,N_952,N_1149);
nor U2146 (N_2146,N_997,N_1358);
nand U2147 (N_2147,N_1464,N_1183);
nand U2148 (N_2148,N_1109,N_1111);
nand U2149 (N_2149,N_1185,N_1480);
and U2150 (N_2150,N_1326,N_1100);
xnor U2151 (N_2151,N_1314,N_759);
nand U2152 (N_2152,N_1116,N_1477);
or U2153 (N_2153,N_1498,N_1097);
or U2154 (N_2154,N_1009,N_753);
nor U2155 (N_2155,N_969,N_916);
and U2156 (N_2156,N_1125,N_1023);
or U2157 (N_2157,N_1184,N_840);
nor U2158 (N_2158,N_1095,N_957);
nand U2159 (N_2159,N_1280,N_1090);
xnor U2160 (N_2160,N_1074,N_763);
or U2161 (N_2161,N_1148,N_751);
nor U2162 (N_2162,N_1256,N_1481);
xnor U2163 (N_2163,N_1338,N_765);
and U2164 (N_2164,N_1463,N_1184);
xor U2165 (N_2165,N_1040,N_1373);
xnor U2166 (N_2166,N_1362,N_1158);
and U2167 (N_2167,N_1051,N_941);
xnor U2168 (N_2168,N_1152,N_1153);
nor U2169 (N_2169,N_1468,N_1058);
and U2170 (N_2170,N_1478,N_980);
nor U2171 (N_2171,N_1129,N_1395);
nor U2172 (N_2172,N_976,N_1275);
nand U2173 (N_2173,N_1475,N_1352);
or U2174 (N_2174,N_782,N_1116);
nand U2175 (N_2175,N_1227,N_1300);
or U2176 (N_2176,N_1270,N_1326);
and U2177 (N_2177,N_800,N_1322);
nor U2178 (N_2178,N_845,N_1433);
or U2179 (N_2179,N_1166,N_784);
or U2180 (N_2180,N_1387,N_758);
nor U2181 (N_2181,N_1080,N_1325);
and U2182 (N_2182,N_858,N_817);
nor U2183 (N_2183,N_774,N_777);
or U2184 (N_2184,N_1092,N_1151);
nand U2185 (N_2185,N_853,N_1397);
or U2186 (N_2186,N_1286,N_887);
or U2187 (N_2187,N_1168,N_1128);
and U2188 (N_2188,N_785,N_841);
nand U2189 (N_2189,N_1477,N_837);
nor U2190 (N_2190,N_1086,N_1226);
nand U2191 (N_2191,N_1099,N_1496);
nor U2192 (N_2192,N_1160,N_1139);
xor U2193 (N_2193,N_1302,N_1369);
nor U2194 (N_2194,N_1135,N_889);
nor U2195 (N_2195,N_1366,N_1180);
xor U2196 (N_2196,N_1016,N_1112);
or U2197 (N_2197,N_1304,N_1470);
nand U2198 (N_2198,N_1299,N_1369);
and U2199 (N_2199,N_974,N_1437);
or U2200 (N_2200,N_1015,N_895);
nand U2201 (N_2201,N_939,N_1453);
nor U2202 (N_2202,N_1037,N_1431);
or U2203 (N_2203,N_1381,N_834);
nor U2204 (N_2204,N_1219,N_1107);
nand U2205 (N_2205,N_1329,N_1372);
nand U2206 (N_2206,N_1273,N_1348);
xor U2207 (N_2207,N_1173,N_1459);
xor U2208 (N_2208,N_1372,N_1187);
nor U2209 (N_2209,N_856,N_1281);
and U2210 (N_2210,N_1465,N_785);
nor U2211 (N_2211,N_1325,N_771);
xnor U2212 (N_2212,N_758,N_1020);
xor U2213 (N_2213,N_1170,N_1325);
xnor U2214 (N_2214,N_1264,N_1093);
and U2215 (N_2215,N_1318,N_1284);
or U2216 (N_2216,N_829,N_1331);
nor U2217 (N_2217,N_1494,N_1362);
xor U2218 (N_2218,N_1473,N_1472);
or U2219 (N_2219,N_952,N_1143);
nand U2220 (N_2220,N_1485,N_1076);
nand U2221 (N_2221,N_969,N_822);
nor U2222 (N_2222,N_1195,N_1299);
and U2223 (N_2223,N_1181,N_1370);
or U2224 (N_2224,N_1135,N_1073);
xor U2225 (N_2225,N_913,N_1314);
xor U2226 (N_2226,N_846,N_881);
or U2227 (N_2227,N_1257,N_1129);
nand U2228 (N_2228,N_1275,N_1030);
nand U2229 (N_2229,N_1293,N_1170);
and U2230 (N_2230,N_764,N_1267);
or U2231 (N_2231,N_839,N_1426);
or U2232 (N_2232,N_872,N_926);
or U2233 (N_2233,N_1194,N_971);
xnor U2234 (N_2234,N_935,N_1410);
or U2235 (N_2235,N_1144,N_1020);
nand U2236 (N_2236,N_1498,N_849);
or U2237 (N_2237,N_1243,N_973);
xor U2238 (N_2238,N_1264,N_1160);
nand U2239 (N_2239,N_1316,N_972);
or U2240 (N_2240,N_1263,N_792);
and U2241 (N_2241,N_1049,N_1098);
nand U2242 (N_2242,N_1299,N_980);
and U2243 (N_2243,N_1091,N_1165);
or U2244 (N_2244,N_1258,N_907);
and U2245 (N_2245,N_1422,N_974);
nand U2246 (N_2246,N_1006,N_947);
xnor U2247 (N_2247,N_1377,N_968);
nor U2248 (N_2248,N_1233,N_1114);
xor U2249 (N_2249,N_1312,N_756);
and U2250 (N_2250,N_1588,N_2035);
xor U2251 (N_2251,N_1921,N_1638);
nand U2252 (N_2252,N_1955,N_1594);
nor U2253 (N_2253,N_2042,N_2131);
and U2254 (N_2254,N_1583,N_2130);
nor U2255 (N_2255,N_1937,N_1502);
or U2256 (N_2256,N_1501,N_1766);
or U2257 (N_2257,N_1891,N_1818);
or U2258 (N_2258,N_1535,N_1702);
xnor U2259 (N_2259,N_1500,N_1799);
xor U2260 (N_2260,N_1716,N_2145);
and U2261 (N_2261,N_1731,N_2040);
xnor U2262 (N_2262,N_1811,N_2037);
or U2263 (N_2263,N_1862,N_2069);
and U2264 (N_2264,N_2210,N_2054);
nor U2265 (N_2265,N_1659,N_2128);
nand U2266 (N_2266,N_2193,N_1604);
and U2267 (N_2267,N_1873,N_2142);
nand U2268 (N_2268,N_1795,N_1900);
xnor U2269 (N_2269,N_1568,N_1925);
nand U2270 (N_2270,N_1929,N_2133);
xnor U2271 (N_2271,N_2020,N_2228);
nor U2272 (N_2272,N_1561,N_1732);
or U2273 (N_2273,N_2244,N_2125);
nand U2274 (N_2274,N_1758,N_1781);
and U2275 (N_2275,N_2078,N_1817);
or U2276 (N_2276,N_2219,N_2099);
and U2277 (N_2277,N_1895,N_1786);
xor U2278 (N_2278,N_1866,N_1823);
nor U2279 (N_2279,N_2033,N_1717);
nor U2280 (N_2280,N_1868,N_1595);
and U2281 (N_2281,N_2190,N_1938);
xor U2282 (N_2282,N_1787,N_2029);
and U2283 (N_2283,N_1510,N_1765);
nand U2284 (N_2284,N_1850,N_1618);
nor U2285 (N_2285,N_1832,N_1773);
nor U2286 (N_2286,N_1730,N_1532);
and U2287 (N_2287,N_1951,N_2081);
nor U2288 (N_2288,N_2160,N_2138);
nor U2289 (N_2289,N_1623,N_2249);
nor U2290 (N_2290,N_1724,N_1720);
and U2291 (N_2291,N_1715,N_1693);
xor U2292 (N_2292,N_2047,N_1905);
xnor U2293 (N_2293,N_1919,N_2007);
or U2294 (N_2294,N_1512,N_1779);
or U2295 (N_2295,N_1549,N_1942);
nor U2296 (N_2296,N_2098,N_1993);
or U2297 (N_2297,N_1975,N_1592);
nor U2298 (N_2298,N_1711,N_1918);
nor U2299 (N_2299,N_1685,N_1644);
nand U2300 (N_2300,N_1987,N_1982);
nand U2301 (N_2301,N_1827,N_2001);
nor U2302 (N_2302,N_1761,N_2004);
or U2303 (N_2303,N_1852,N_1701);
or U2304 (N_2304,N_1760,N_1869);
or U2305 (N_2305,N_2218,N_1762);
nand U2306 (N_2306,N_1603,N_2167);
nand U2307 (N_2307,N_1554,N_2231);
nor U2308 (N_2308,N_2154,N_2019);
and U2309 (N_2309,N_1718,N_1859);
or U2310 (N_2310,N_1733,N_2215);
and U2311 (N_2311,N_1804,N_1681);
and U2312 (N_2312,N_1943,N_1930);
nor U2313 (N_2313,N_2191,N_2075);
nand U2314 (N_2314,N_2089,N_1609);
nand U2315 (N_2315,N_1646,N_2000);
or U2316 (N_2316,N_1573,N_1547);
and U2317 (N_2317,N_1524,N_1962);
and U2318 (N_2318,N_1727,N_2065);
or U2319 (N_2319,N_2158,N_2101);
or U2320 (N_2320,N_2073,N_1700);
nor U2321 (N_2321,N_1843,N_1589);
xor U2322 (N_2322,N_1878,N_2083);
or U2323 (N_2323,N_1548,N_2201);
nor U2324 (N_2324,N_1751,N_1519);
xnor U2325 (N_2325,N_1771,N_1793);
xor U2326 (N_2326,N_1876,N_1617);
xor U2327 (N_2327,N_1903,N_2064);
xor U2328 (N_2328,N_2150,N_1995);
nand U2329 (N_2329,N_1841,N_1978);
nor U2330 (N_2330,N_2076,N_2161);
or U2331 (N_2331,N_1775,N_2146);
and U2332 (N_2332,N_1965,N_1916);
or U2333 (N_2333,N_1650,N_1739);
nor U2334 (N_2334,N_1531,N_1879);
nand U2335 (N_2335,N_1522,N_1507);
nand U2336 (N_2336,N_2237,N_1714);
nand U2337 (N_2337,N_2038,N_1536);
nor U2338 (N_2338,N_1577,N_1661);
nand U2339 (N_2339,N_1515,N_2196);
xnor U2340 (N_2340,N_1503,N_2238);
and U2341 (N_2341,N_2002,N_1858);
or U2342 (N_2342,N_1648,N_1846);
and U2343 (N_2343,N_1587,N_2243);
and U2344 (N_2344,N_1822,N_1719);
and U2345 (N_2345,N_1615,N_2032);
or U2346 (N_2346,N_1584,N_1655);
or U2347 (N_2347,N_2119,N_1602);
and U2348 (N_2348,N_1516,N_2204);
nand U2349 (N_2349,N_1687,N_1541);
and U2350 (N_2350,N_1863,N_1520);
or U2351 (N_2351,N_1745,N_1525);
nor U2352 (N_2352,N_1576,N_2009);
or U2353 (N_2353,N_2071,N_2092);
nand U2354 (N_2354,N_1906,N_1941);
and U2355 (N_2355,N_1569,N_2124);
nand U2356 (N_2356,N_1729,N_2107);
xnor U2357 (N_2357,N_1979,N_1922);
xor U2358 (N_2358,N_2012,N_2052);
nor U2359 (N_2359,N_1657,N_1959);
nand U2360 (N_2360,N_1805,N_1580);
or U2361 (N_2361,N_1593,N_1776);
nor U2362 (N_2362,N_1754,N_2147);
nand U2363 (N_2363,N_1808,N_1660);
xor U2364 (N_2364,N_1677,N_1509);
xnor U2365 (N_2365,N_2227,N_1894);
nand U2366 (N_2366,N_1986,N_1964);
xor U2367 (N_2367,N_1789,N_1728);
nor U2368 (N_2368,N_2139,N_1833);
nor U2369 (N_2369,N_2159,N_1777);
and U2370 (N_2370,N_2212,N_1981);
or U2371 (N_2371,N_1713,N_1667);
nor U2372 (N_2372,N_1997,N_2103);
or U2373 (N_2373,N_1600,N_2061);
nand U2374 (N_2374,N_2121,N_1813);
or U2375 (N_2375,N_2077,N_1632);
or U2376 (N_2376,N_1668,N_1526);
nor U2377 (N_2377,N_1924,N_1555);
nand U2378 (N_2378,N_1613,N_1690);
xnor U2379 (N_2379,N_1725,N_1686);
xor U2380 (N_2380,N_1505,N_1723);
nand U2381 (N_2381,N_1735,N_1898);
or U2382 (N_2382,N_1683,N_1630);
nor U2383 (N_2383,N_1865,N_1666);
xnor U2384 (N_2384,N_2053,N_1738);
nor U2385 (N_2385,N_1904,N_1742);
nor U2386 (N_2386,N_1928,N_2187);
or U2387 (N_2387,N_2015,N_1886);
nor U2388 (N_2388,N_1802,N_1971);
or U2389 (N_2389,N_1914,N_1896);
xor U2390 (N_2390,N_2156,N_1881);
nor U2391 (N_2391,N_1992,N_1910);
or U2392 (N_2392,N_1639,N_2174);
xnor U2393 (N_2393,N_2030,N_2140);
nor U2394 (N_2394,N_1734,N_2018);
xnor U2395 (N_2395,N_1698,N_2118);
nor U2396 (N_2396,N_1557,N_1750);
xor U2397 (N_2397,N_2178,N_2005);
or U2398 (N_2398,N_2200,N_2134);
and U2399 (N_2399,N_2149,N_2170);
nor U2400 (N_2400,N_1736,N_1915);
or U2401 (N_2401,N_2136,N_1572);
and U2402 (N_2402,N_1926,N_1917);
xor U2403 (N_2403,N_1949,N_1848);
nor U2404 (N_2404,N_2006,N_1860);
nand U2405 (N_2405,N_1958,N_1670);
nand U2406 (N_2406,N_1744,N_1654);
nor U2407 (N_2407,N_1882,N_1829);
xnor U2408 (N_2408,N_2180,N_1712);
nand U2409 (N_2409,N_1820,N_1796);
nand U2410 (N_2410,N_1642,N_1633);
nand U2411 (N_2411,N_1870,N_1601);
or U2412 (N_2412,N_1697,N_1912);
nand U2413 (N_2413,N_1945,N_2176);
nor U2414 (N_2414,N_1977,N_2059);
and U2415 (N_2415,N_2116,N_2230);
or U2416 (N_2416,N_1983,N_1556);
nand U2417 (N_2417,N_1991,N_2063);
or U2418 (N_2418,N_1647,N_1880);
or U2419 (N_2419,N_2179,N_1980);
or U2420 (N_2420,N_1746,N_2185);
and U2421 (N_2421,N_2085,N_1560);
nand U2422 (N_2422,N_1902,N_1952);
nor U2423 (N_2423,N_1994,N_1907);
or U2424 (N_2424,N_1830,N_1884);
xnor U2425 (N_2425,N_2031,N_2127);
and U2426 (N_2426,N_2143,N_2206);
nor U2427 (N_2427,N_1612,N_1790);
or U2428 (N_2428,N_1857,N_1757);
nor U2429 (N_2429,N_2199,N_1565);
nor U2430 (N_2430,N_1671,N_1707);
xor U2431 (N_2431,N_1631,N_1996);
nor U2432 (N_2432,N_1944,N_2025);
nor U2433 (N_2433,N_2056,N_2144);
nand U2434 (N_2434,N_1564,N_1774);
and U2435 (N_2435,N_1756,N_1570);
or U2436 (N_2436,N_1845,N_1598);
or U2437 (N_2437,N_2216,N_2241);
xor U2438 (N_2438,N_2057,N_1544);
nor U2439 (N_2439,N_1798,N_1956);
and U2440 (N_2440,N_1933,N_1967);
xnor U2441 (N_2441,N_2095,N_1622);
and U2442 (N_2442,N_1763,N_2058);
and U2443 (N_2443,N_1923,N_2188);
nand U2444 (N_2444,N_1663,N_1546);
xnor U2445 (N_2445,N_1567,N_1909);
and U2446 (N_2446,N_1726,N_1741);
and U2447 (N_2447,N_2202,N_2235);
or U2448 (N_2448,N_1606,N_2164);
nor U2449 (N_2449,N_2186,N_1966);
and U2450 (N_2450,N_1753,N_1940);
or U2451 (N_2451,N_1534,N_1699);
xnor U2452 (N_2452,N_1759,N_1785);
or U2453 (N_2453,N_2106,N_1538);
xor U2454 (N_2454,N_1575,N_2192);
or U2455 (N_2455,N_1597,N_1984);
nor U2456 (N_2456,N_1563,N_1792);
nor U2457 (N_2457,N_1935,N_2181);
and U2458 (N_2458,N_1769,N_1694);
or U2459 (N_2459,N_2036,N_2114);
or U2460 (N_2460,N_1607,N_1772);
xor U2461 (N_2461,N_2189,N_1897);
xnor U2462 (N_2462,N_1559,N_2248);
xor U2463 (N_2463,N_1801,N_1871);
nand U2464 (N_2464,N_2122,N_1619);
nand U2465 (N_2465,N_1558,N_2014);
xnor U2466 (N_2466,N_1540,N_1616);
xnor U2467 (N_2467,N_1867,N_2112);
nand U2468 (N_2468,N_2003,N_2080);
xor U2469 (N_2469,N_2104,N_1627);
xnor U2470 (N_2470,N_1851,N_1810);
xor U2471 (N_2471,N_1842,N_2207);
nor U2472 (N_2472,N_1674,N_2166);
nand U2473 (N_2473,N_1614,N_1824);
and U2474 (N_2474,N_1656,N_1834);
nand U2475 (N_2475,N_1840,N_1770);
xor U2476 (N_2476,N_1913,N_1853);
nor U2477 (N_2477,N_2108,N_1875);
and U2478 (N_2478,N_1936,N_2022);
and U2479 (N_2479,N_1528,N_2197);
xor U2480 (N_2480,N_2094,N_2070);
nand U2481 (N_2481,N_1791,N_1826);
or U2482 (N_2482,N_1571,N_1856);
or U2483 (N_2483,N_2162,N_2229);
or U2484 (N_2484,N_2152,N_1696);
or U2485 (N_2485,N_2110,N_1839);
xor U2486 (N_2486,N_2087,N_1539);
and U2487 (N_2487,N_2232,N_1678);
and U2488 (N_2488,N_1920,N_1947);
nor U2489 (N_2489,N_2100,N_2097);
xnor U2490 (N_2490,N_1518,N_1585);
nor U2491 (N_2491,N_1797,N_2026);
xor U2492 (N_2492,N_2074,N_2226);
xnor U2493 (N_2493,N_1970,N_1605);
xnor U2494 (N_2494,N_1838,N_2214);
or U2495 (N_2495,N_2165,N_2048);
or U2496 (N_2496,N_2023,N_2046);
and U2497 (N_2497,N_2172,N_1809);
nor U2498 (N_2498,N_1523,N_2184);
nand U2499 (N_2499,N_1888,N_1596);
xor U2500 (N_2500,N_1625,N_2039);
nand U2501 (N_2501,N_1533,N_2017);
and U2502 (N_2502,N_1511,N_1844);
and U2503 (N_2503,N_1504,N_1855);
nor U2504 (N_2504,N_1662,N_1957);
and U2505 (N_2505,N_2011,N_1768);
nor U2506 (N_2506,N_2247,N_1645);
or U2507 (N_2507,N_1961,N_1643);
nand U2508 (N_2508,N_2240,N_2008);
nand U2509 (N_2509,N_1553,N_2067);
nand U2510 (N_2510,N_1931,N_1691);
xor U2511 (N_2511,N_2105,N_1954);
xnor U2512 (N_2512,N_2091,N_1972);
nor U2513 (N_2513,N_1989,N_1828);
or U2514 (N_2514,N_1579,N_2126);
nor U2515 (N_2515,N_2177,N_2198);
and U2516 (N_2516,N_2169,N_1883);
and U2517 (N_2517,N_2123,N_1819);
and U2518 (N_2518,N_2088,N_2168);
or U2519 (N_2519,N_1665,N_1621);
nand U2520 (N_2520,N_2148,N_1710);
or U2521 (N_2521,N_1749,N_1658);
xnor U2522 (N_2522,N_2044,N_1814);
nor U2523 (N_2523,N_2171,N_2084);
or U2524 (N_2524,N_1529,N_1624);
or U2525 (N_2525,N_2027,N_2221);
and U2526 (N_2526,N_1651,N_2217);
xnor U2527 (N_2527,N_2157,N_1586);
nor U2528 (N_2528,N_1740,N_1752);
nor U2529 (N_2529,N_2109,N_1543);
or U2530 (N_2530,N_1517,N_2016);
and U2531 (N_2531,N_1976,N_1927);
xor U2532 (N_2532,N_1675,N_2111);
and U2533 (N_2533,N_1590,N_2024);
nand U2534 (N_2534,N_1889,N_1950);
nor U2535 (N_2535,N_1704,N_1932);
or U2536 (N_2536,N_1599,N_2141);
nor U2537 (N_2537,N_2233,N_1640);
xor U2538 (N_2538,N_1649,N_1849);
xnor U2539 (N_2539,N_1591,N_1999);
xor U2540 (N_2540,N_1684,N_1626);
and U2541 (N_2541,N_1953,N_1706);
nand U2542 (N_2542,N_1708,N_1688);
xnor U2543 (N_2543,N_1821,N_1969);
nor U2544 (N_2544,N_1815,N_1676);
or U2545 (N_2545,N_2153,N_2209);
and U2546 (N_2546,N_1506,N_1783);
nand U2547 (N_2547,N_2182,N_2137);
and U2548 (N_2548,N_1721,N_1990);
xor U2549 (N_2549,N_2183,N_1737);
nor U2550 (N_2550,N_1514,N_2203);
or U2551 (N_2551,N_1610,N_1861);
and U2552 (N_2552,N_1872,N_1825);
nand U2553 (N_2553,N_2055,N_2050);
xnor U2554 (N_2554,N_2090,N_2086);
and U2555 (N_2555,N_1934,N_1703);
and U2556 (N_2556,N_1582,N_2068);
or U2557 (N_2557,N_2102,N_2021);
or U2558 (N_2558,N_2060,N_1963);
nand U2559 (N_2559,N_1530,N_1574);
nor U2560 (N_2560,N_1545,N_1669);
nand U2561 (N_2561,N_1782,N_1513);
xnor U2562 (N_2562,N_2010,N_1911);
nor U2563 (N_2563,N_1835,N_2028);
and U2564 (N_2564,N_1709,N_2041);
nor U2565 (N_2565,N_2173,N_1901);
nor U2566 (N_2566,N_2245,N_1641);
or U2567 (N_2567,N_1946,N_2223);
or U2568 (N_2568,N_1695,N_1508);
and U2569 (N_2569,N_2096,N_2163);
xnor U2570 (N_2570,N_2205,N_2155);
nor U2571 (N_2571,N_2062,N_2082);
nand U2572 (N_2572,N_2093,N_2213);
nand U2573 (N_2573,N_2222,N_1784);
nand U2574 (N_2574,N_1974,N_2120);
nor U2575 (N_2575,N_2113,N_2234);
nand U2576 (N_2576,N_1988,N_1664);
or U2577 (N_2577,N_1652,N_1800);
nand U2578 (N_2578,N_1635,N_1854);
nand U2579 (N_2579,N_1973,N_1885);
nor U2580 (N_2580,N_1620,N_1679);
xnor U2581 (N_2581,N_1899,N_1550);
and U2582 (N_2582,N_2220,N_2049);
xnor U2583 (N_2583,N_1836,N_2208);
xor U2584 (N_2584,N_1890,N_1521);
nor U2585 (N_2585,N_1755,N_1788);
nand U2586 (N_2586,N_1968,N_1780);
and U2587 (N_2587,N_2225,N_1552);
and U2588 (N_2588,N_1743,N_1812);
or U2589 (N_2589,N_1893,N_2045);
and U2590 (N_2590,N_1998,N_1634);
nor U2591 (N_2591,N_1939,N_1537);
nand U2592 (N_2592,N_1837,N_1673);
or U2593 (N_2593,N_1611,N_1689);
nor U2594 (N_2594,N_1892,N_2115);
nor U2595 (N_2595,N_1747,N_1985);
nand U2596 (N_2596,N_1692,N_2211);
or U2597 (N_2597,N_2239,N_1562);
and U2598 (N_2598,N_2034,N_1672);
or U2599 (N_2599,N_1764,N_2194);
xnor U2600 (N_2600,N_2224,N_2236);
xor U2601 (N_2601,N_1566,N_1551);
nor U2602 (N_2602,N_2079,N_1803);
or U2603 (N_2603,N_1581,N_1960);
and U2604 (N_2604,N_2195,N_2151);
or U2605 (N_2605,N_2242,N_1908);
nand U2606 (N_2606,N_1847,N_1637);
nand U2607 (N_2607,N_1608,N_1794);
nand U2608 (N_2608,N_1887,N_1874);
and U2609 (N_2609,N_1767,N_1722);
nand U2610 (N_2610,N_1542,N_1877);
and U2611 (N_2611,N_1527,N_2043);
nand U2612 (N_2612,N_2246,N_2117);
nor U2613 (N_2613,N_2013,N_1831);
and U2614 (N_2614,N_1682,N_2072);
and U2615 (N_2615,N_1748,N_2175);
nand U2616 (N_2616,N_1806,N_1816);
or U2617 (N_2617,N_1807,N_1948);
nand U2618 (N_2618,N_1705,N_1628);
nor U2619 (N_2619,N_1629,N_1864);
nand U2620 (N_2620,N_2129,N_1778);
nand U2621 (N_2621,N_2051,N_2132);
or U2622 (N_2622,N_1636,N_1680);
or U2623 (N_2623,N_2066,N_1578);
xor U2624 (N_2624,N_1653,N_2135);
nand U2625 (N_2625,N_1755,N_1656);
xnor U2626 (N_2626,N_2119,N_1552);
nand U2627 (N_2627,N_1600,N_1604);
nand U2628 (N_2628,N_1569,N_1620);
and U2629 (N_2629,N_1712,N_1980);
nor U2630 (N_2630,N_2025,N_2045);
nand U2631 (N_2631,N_1626,N_1771);
and U2632 (N_2632,N_1667,N_1619);
xnor U2633 (N_2633,N_1981,N_1920);
or U2634 (N_2634,N_1860,N_1714);
xor U2635 (N_2635,N_2012,N_2233);
xor U2636 (N_2636,N_1617,N_2073);
nor U2637 (N_2637,N_1523,N_1605);
xor U2638 (N_2638,N_2232,N_2197);
and U2639 (N_2639,N_1963,N_1802);
nor U2640 (N_2640,N_2175,N_2172);
or U2641 (N_2641,N_1564,N_1830);
xor U2642 (N_2642,N_1778,N_1915);
nand U2643 (N_2643,N_1782,N_1970);
or U2644 (N_2644,N_1987,N_1542);
xnor U2645 (N_2645,N_2198,N_2027);
nand U2646 (N_2646,N_1957,N_1709);
nand U2647 (N_2647,N_1891,N_1905);
nor U2648 (N_2648,N_2055,N_1771);
nor U2649 (N_2649,N_1808,N_2198);
and U2650 (N_2650,N_1620,N_2157);
nor U2651 (N_2651,N_2047,N_1925);
nor U2652 (N_2652,N_1999,N_1985);
and U2653 (N_2653,N_1875,N_1591);
nand U2654 (N_2654,N_2175,N_1959);
nand U2655 (N_2655,N_1774,N_2033);
and U2656 (N_2656,N_2153,N_1526);
nand U2657 (N_2657,N_2010,N_2211);
and U2658 (N_2658,N_1866,N_2052);
xnor U2659 (N_2659,N_1791,N_2048);
and U2660 (N_2660,N_2018,N_1755);
nand U2661 (N_2661,N_1802,N_1705);
nand U2662 (N_2662,N_1978,N_1635);
xor U2663 (N_2663,N_2132,N_1573);
or U2664 (N_2664,N_2202,N_1729);
or U2665 (N_2665,N_1678,N_1947);
and U2666 (N_2666,N_1584,N_1896);
or U2667 (N_2667,N_2189,N_1658);
nor U2668 (N_2668,N_2242,N_1864);
xnor U2669 (N_2669,N_2152,N_2189);
xnor U2670 (N_2670,N_1544,N_1968);
or U2671 (N_2671,N_2220,N_1969);
xnor U2672 (N_2672,N_2038,N_1783);
xnor U2673 (N_2673,N_1652,N_1859);
nand U2674 (N_2674,N_1938,N_1846);
nand U2675 (N_2675,N_1756,N_1852);
nor U2676 (N_2676,N_2039,N_1801);
xor U2677 (N_2677,N_1831,N_2067);
xor U2678 (N_2678,N_1873,N_1815);
nand U2679 (N_2679,N_1837,N_2236);
nor U2680 (N_2680,N_2039,N_2244);
xnor U2681 (N_2681,N_1867,N_1754);
nand U2682 (N_2682,N_2018,N_1600);
and U2683 (N_2683,N_2158,N_2047);
nand U2684 (N_2684,N_1883,N_2152);
nand U2685 (N_2685,N_1553,N_1944);
nor U2686 (N_2686,N_1991,N_2171);
or U2687 (N_2687,N_1958,N_1983);
and U2688 (N_2688,N_1750,N_2095);
xnor U2689 (N_2689,N_1775,N_1705);
xor U2690 (N_2690,N_1720,N_2054);
nand U2691 (N_2691,N_1845,N_2124);
and U2692 (N_2692,N_2149,N_2013);
and U2693 (N_2693,N_1821,N_1763);
nor U2694 (N_2694,N_1931,N_1683);
nor U2695 (N_2695,N_1700,N_1681);
or U2696 (N_2696,N_1765,N_2073);
xor U2697 (N_2697,N_1740,N_1660);
nand U2698 (N_2698,N_1725,N_2057);
nor U2699 (N_2699,N_2123,N_1736);
or U2700 (N_2700,N_1765,N_1687);
or U2701 (N_2701,N_1530,N_2056);
xor U2702 (N_2702,N_1576,N_1949);
nor U2703 (N_2703,N_1591,N_1771);
or U2704 (N_2704,N_2000,N_1909);
and U2705 (N_2705,N_2126,N_2090);
nand U2706 (N_2706,N_2186,N_1654);
nand U2707 (N_2707,N_2021,N_2027);
nand U2708 (N_2708,N_1529,N_2242);
nor U2709 (N_2709,N_1877,N_1507);
nor U2710 (N_2710,N_2101,N_2078);
nor U2711 (N_2711,N_1798,N_2059);
and U2712 (N_2712,N_2013,N_2109);
or U2713 (N_2713,N_2098,N_1956);
xor U2714 (N_2714,N_1866,N_1796);
and U2715 (N_2715,N_1573,N_2211);
and U2716 (N_2716,N_1560,N_2133);
nor U2717 (N_2717,N_1846,N_2034);
xor U2718 (N_2718,N_1739,N_2094);
xnor U2719 (N_2719,N_1982,N_1737);
or U2720 (N_2720,N_1691,N_1755);
and U2721 (N_2721,N_1549,N_2190);
nor U2722 (N_2722,N_2153,N_1623);
nor U2723 (N_2723,N_1657,N_1786);
xor U2724 (N_2724,N_2171,N_1701);
and U2725 (N_2725,N_2218,N_2123);
nand U2726 (N_2726,N_1670,N_2139);
or U2727 (N_2727,N_2223,N_1953);
or U2728 (N_2728,N_2054,N_1567);
nand U2729 (N_2729,N_2063,N_2057);
nor U2730 (N_2730,N_2003,N_1756);
or U2731 (N_2731,N_2035,N_2108);
or U2732 (N_2732,N_1830,N_1559);
nand U2733 (N_2733,N_1759,N_1522);
and U2734 (N_2734,N_1999,N_2145);
xnor U2735 (N_2735,N_2160,N_1829);
nand U2736 (N_2736,N_2208,N_1703);
nand U2737 (N_2737,N_1654,N_1709);
nor U2738 (N_2738,N_2063,N_1849);
nand U2739 (N_2739,N_2221,N_1606);
and U2740 (N_2740,N_1695,N_1767);
or U2741 (N_2741,N_2242,N_1632);
nor U2742 (N_2742,N_1837,N_2024);
nor U2743 (N_2743,N_2063,N_1759);
nand U2744 (N_2744,N_2131,N_2150);
nor U2745 (N_2745,N_1881,N_1725);
and U2746 (N_2746,N_1980,N_1937);
xor U2747 (N_2747,N_1986,N_2059);
xnor U2748 (N_2748,N_1718,N_1768);
and U2749 (N_2749,N_1881,N_1708);
xor U2750 (N_2750,N_1656,N_1717);
or U2751 (N_2751,N_2100,N_2028);
xor U2752 (N_2752,N_1599,N_1654);
xor U2753 (N_2753,N_1572,N_1605);
and U2754 (N_2754,N_2145,N_2115);
nand U2755 (N_2755,N_2117,N_1569);
or U2756 (N_2756,N_1788,N_2197);
and U2757 (N_2757,N_1895,N_1957);
and U2758 (N_2758,N_1890,N_1765);
nor U2759 (N_2759,N_2200,N_1736);
xor U2760 (N_2760,N_1894,N_1845);
nand U2761 (N_2761,N_1783,N_2138);
or U2762 (N_2762,N_1544,N_1890);
or U2763 (N_2763,N_1946,N_2219);
nor U2764 (N_2764,N_1904,N_1738);
nor U2765 (N_2765,N_2027,N_1616);
xor U2766 (N_2766,N_2024,N_1692);
xor U2767 (N_2767,N_1885,N_1575);
xor U2768 (N_2768,N_1634,N_2189);
or U2769 (N_2769,N_2019,N_1724);
and U2770 (N_2770,N_1955,N_1588);
or U2771 (N_2771,N_2151,N_2223);
nor U2772 (N_2772,N_1862,N_2126);
nor U2773 (N_2773,N_1755,N_1649);
nand U2774 (N_2774,N_1853,N_1606);
nand U2775 (N_2775,N_1748,N_1815);
xnor U2776 (N_2776,N_2025,N_1639);
nor U2777 (N_2777,N_1921,N_2044);
nand U2778 (N_2778,N_1808,N_1864);
or U2779 (N_2779,N_1964,N_2180);
or U2780 (N_2780,N_2050,N_1665);
nand U2781 (N_2781,N_1576,N_1880);
xor U2782 (N_2782,N_2201,N_1842);
nor U2783 (N_2783,N_2035,N_1621);
or U2784 (N_2784,N_1603,N_1774);
and U2785 (N_2785,N_2022,N_2005);
nor U2786 (N_2786,N_1835,N_1608);
nand U2787 (N_2787,N_1915,N_1840);
nand U2788 (N_2788,N_2125,N_1689);
nand U2789 (N_2789,N_2072,N_2080);
or U2790 (N_2790,N_2167,N_1659);
xnor U2791 (N_2791,N_1628,N_1901);
nand U2792 (N_2792,N_1769,N_1876);
nor U2793 (N_2793,N_1888,N_1546);
nor U2794 (N_2794,N_1685,N_1869);
nor U2795 (N_2795,N_1986,N_1769);
and U2796 (N_2796,N_1688,N_2153);
or U2797 (N_2797,N_1869,N_1705);
nand U2798 (N_2798,N_1505,N_2102);
and U2799 (N_2799,N_1562,N_2109);
xnor U2800 (N_2800,N_1528,N_2245);
and U2801 (N_2801,N_2111,N_1797);
nor U2802 (N_2802,N_1604,N_2048);
or U2803 (N_2803,N_1603,N_1706);
or U2804 (N_2804,N_2039,N_2238);
or U2805 (N_2805,N_1661,N_1923);
nor U2806 (N_2806,N_1872,N_1575);
and U2807 (N_2807,N_1954,N_1642);
nor U2808 (N_2808,N_1981,N_1568);
xor U2809 (N_2809,N_2164,N_1805);
nand U2810 (N_2810,N_2237,N_1713);
xor U2811 (N_2811,N_2130,N_1982);
and U2812 (N_2812,N_1983,N_2075);
or U2813 (N_2813,N_1671,N_1929);
nand U2814 (N_2814,N_1906,N_1705);
nand U2815 (N_2815,N_1715,N_1646);
xor U2816 (N_2816,N_1934,N_1919);
or U2817 (N_2817,N_1980,N_1758);
or U2818 (N_2818,N_1626,N_2153);
and U2819 (N_2819,N_2102,N_1594);
or U2820 (N_2820,N_1700,N_2070);
xnor U2821 (N_2821,N_1717,N_2105);
nor U2822 (N_2822,N_2022,N_1998);
nor U2823 (N_2823,N_1971,N_1817);
nor U2824 (N_2824,N_1671,N_2236);
nand U2825 (N_2825,N_2197,N_2043);
nand U2826 (N_2826,N_2119,N_1524);
nand U2827 (N_2827,N_1893,N_2109);
or U2828 (N_2828,N_1761,N_2201);
nand U2829 (N_2829,N_2015,N_1817);
and U2830 (N_2830,N_2129,N_1767);
nor U2831 (N_2831,N_1902,N_1671);
nand U2832 (N_2832,N_1731,N_1712);
nor U2833 (N_2833,N_1780,N_1857);
nand U2834 (N_2834,N_1736,N_1868);
or U2835 (N_2835,N_1923,N_1626);
nor U2836 (N_2836,N_1677,N_1806);
nor U2837 (N_2837,N_2208,N_1970);
and U2838 (N_2838,N_2079,N_2176);
xor U2839 (N_2839,N_1561,N_1955);
xor U2840 (N_2840,N_1802,N_1901);
nor U2841 (N_2841,N_1949,N_1943);
and U2842 (N_2842,N_1923,N_2213);
and U2843 (N_2843,N_2043,N_1683);
nand U2844 (N_2844,N_2237,N_2157);
xnor U2845 (N_2845,N_2106,N_1573);
nor U2846 (N_2846,N_1991,N_2196);
and U2847 (N_2847,N_2236,N_1976);
and U2848 (N_2848,N_1993,N_1560);
nor U2849 (N_2849,N_1914,N_1535);
xor U2850 (N_2850,N_2174,N_2239);
nor U2851 (N_2851,N_1899,N_1837);
and U2852 (N_2852,N_1871,N_1739);
or U2853 (N_2853,N_1747,N_1905);
xnor U2854 (N_2854,N_1658,N_1672);
nand U2855 (N_2855,N_2247,N_1736);
nor U2856 (N_2856,N_1950,N_2159);
nor U2857 (N_2857,N_2240,N_1818);
xnor U2858 (N_2858,N_1856,N_1854);
xor U2859 (N_2859,N_1526,N_2110);
nor U2860 (N_2860,N_2176,N_2039);
xor U2861 (N_2861,N_2085,N_2222);
nor U2862 (N_2862,N_2120,N_2100);
xnor U2863 (N_2863,N_1580,N_2071);
xnor U2864 (N_2864,N_2118,N_1682);
nand U2865 (N_2865,N_1503,N_1726);
and U2866 (N_2866,N_2228,N_1785);
nor U2867 (N_2867,N_1890,N_1944);
xnor U2868 (N_2868,N_2038,N_1507);
or U2869 (N_2869,N_1937,N_2165);
xor U2870 (N_2870,N_2189,N_1841);
nor U2871 (N_2871,N_2149,N_1623);
or U2872 (N_2872,N_1932,N_2171);
or U2873 (N_2873,N_1708,N_1607);
and U2874 (N_2874,N_2109,N_1530);
nor U2875 (N_2875,N_1564,N_2124);
xor U2876 (N_2876,N_2059,N_1837);
nand U2877 (N_2877,N_2074,N_1693);
and U2878 (N_2878,N_1921,N_2057);
xnor U2879 (N_2879,N_1823,N_1888);
nand U2880 (N_2880,N_2089,N_2026);
xor U2881 (N_2881,N_1850,N_2143);
or U2882 (N_2882,N_1662,N_1791);
xnor U2883 (N_2883,N_1671,N_1863);
and U2884 (N_2884,N_2196,N_1665);
and U2885 (N_2885,N_1785,N_1566);
nor U2886 (N_2886,N_2183,N_2155);
xor U2887 (N_2887,N_1980,N_1511);
nor U2888 (N_2888,N_1908,N_1501);
xor U2889 (N_2889,N_1807,N_2065);
xnor U2890 (N_2890,N_2150,N_1965);
nor U2891 (N_2891,N_1580,N_2176);
nor U2892 (N_2892,N_1889,N_1554);
nor U2893 (N_2893,N_2004,N_1802);
or U2894 (N_2894,N_1691,N_1525);
xor U2895 (N_2895,N_1886,N_1723);
and U2896 (N_2896,N_2044,N_1931);
nor U2897 (N_2897,N_1515,N_2173);
nor U2898 (N_2898,N_2083,N_1799);
xor U2899 (N_2899,N_1926,N_1836);
or U2900 (N_2900,N_2218,N_2065);
nand U2901 (N_2901,N_1978,N_1988);
and U2902 (N_2902,N_2015,N_2245);
xor U2903 (N_2903,N_2152,N_2083);
xor U2904 (N_2904,N_2190,N_1718);
nor U2905 (N_2905,N_1706,N_1545);
nor U2906 (N_2906,N_2169,N_1517);
and U2907 (N_2907,N_2025,N_1910);
xor U2908 (N_2908,N_1574,N_1816);
nor U2909 (N_2909,N_2078,N_1724);
nor U2910 (N_2910,N_2062,N_1704);
or U2911 (N_2911,N_1884,N_1725);
xnor U2912 (N_2912,N_1979,N_1604);
xor U2913 (N_2913,N_1742,N_2093);
nand U2914 (N_2914,N_1706,N_1613);
nand U2915 (N_2915,N_1569,N_2062);
or U2916 (N_2916,N_2068,N_2054);
or U2917 (N_2917,N_2096,N_1579);
or U2918 (N_2918,N_1942,N_1936);
or U2919 (N_2919,N_1993,N_2246);
nor U2920 (N_2920,N_1760,N_2032);
xnor U2921 (N_2921,N_1599,N_1850);
or U2922 (N_2922,N_1723,N_1688);
or U2923 (N_2923,N_2226,N_1537);
or U2924 (N_2924,N_1777,N_1982);
xnor U2925 (N_2925,N_2166,N_1572);
nand U2926 (N_2926,N_1896,N_1726);
nand U2927 (N_2927,N_2045,N_1944);
nor U2928 (N_2928,N_1890,N_1595);
nor U2929 (N_2929,N_1859,N_2120);
or U2930 (N_2930,N_1672,N_1856);
nor U2931 (N_2931,N_2174,N_1710);
and U2932 (N_2932,N_1890,N_1533);
or U2933 (N_2933,N_1975,N_1520);
nand U2934 (N_2934,N_2193,N_2056);
nor U2935 (N_2935,N_2013,N_1617);
nand U2936 (N_2936,N_1745,N_2185);
nor U2937 (N_2937,N_1781,N_2119);
nor U2938 (N_2938,N_1825,N_2170);
nor U2939 (N_2939,N_2195,N_2159);
xnor U2940 (N_2940,N_1921,N_1929);
nand U2941 (N_2941,N_1523,N_2180);
and U2942 (N_2942,N_2007,N_1895);
nor U2943 (N_2943,N_1967,N_1617);
nor U2944 (N_2944,N_1623,N_1822);
nand U2945 (N_2945,N_1574,N_1626);
and U2946 (N_2946,N_1638,N_1510);
xnor U2947 (N_2947,N_2094,N_2041);
nor U2948 (N_2948,N_1879,N_2001);
xor U2949 (N_2949,N_1755,N_1598);
or U2950 (N_2950,N_1825,N_1796);
nor U2951 (N_2951,N_2165,N_1932);
xnor U2952 (N_2952,N_1868,N_2001);
xnor U2953 (N_2953,N_1655,N_1795);
or U2954 (N_2954,N_1754,N_1595);
nor U2955 (N_2955,N_1892,N_1681);
or U2956 (N_2956,N_2059,N_2105);
xor U2957 (N_2957,N_2161,N_1683);
nand U2958 (N_2958,N_1614,N_2015);
xor U2959 (N_2959,N_1993,N_2004);
or U2960 (N_2960,N_1591,N_1945);
or U2961 (N_2961,N_1838,N_1951);
nor U2962 (N_2962,N_1536,N_1630);
nor U2963 (N_2963,N_2077,N_2074);
or U2964 (N_2964,N_1920,N_2182);
nand U2965 (N_2965,N_2141,N_1884);
xnor U2966 (N_2966,N_1641,N_2079);
nand U2967 (N_2967,N_1964,N_1536);
nand U2968 (N_2968,N_2109,N_1896);
nor U2969 (N_2969,N_1858,N_1699);
nand U2970 (N_2970,N_1783,N_2097);
and U2971 (N_2971,N_1744,N_1626);
nor U2972 (N_2972,N_2198,N_1917);
xor U2973 (N_2973,N_2007,N_1739);
xnor U2974 (N_2974,N_1963,N_2086);
nand U2975 (N_2975,N_2196,N_1777);
nor U2976 (N_2976,N_2080,N_1923);
xor U2977 (N_2977,N_1536,N_1530);
nand U2978 (N_2978,N_1706,N_1814);
xnor U2979 (N_2979,N_2215,N_1647);
xnor U2980 (N_2980,N_2168,N_1721);
or U2981 (N_2981,N_1846,N_2210);
or U2982 (N_2982,N_1691,N_1989);
nand U2983 (N_2983,N_1716,N_1867);
and U2984 (N_2984,N_1572,N_1597);
nand U2985 (N_2985,N_1527,N_1610);
nor U2986 (N_2986,N_1928,N_1673);
nand U2987 (N_2987,N_2144,N_1709);
xor U2988 (N_2988,N_2172,N_1689);
and U2989 (N_2989,N_1669,N_1557);
xor U2990 (N_2990,N_1686,N_2044);
or U2991 (N_2991,N_1755,N_2008);
nand U2992 (N_2992,N_2147,N_2120);
and U2993 (N_2993,N_2206,N_1681);
nand U2994 (N_2994,N_2149,N_1720);
and U2995 (N_2995,N_2003,N_2127);
and U2996 (N_2996,N_1702,N_1943);
or U2997 (N_2997,N_2048,N_1696);
nor U2998 (N_2998,N_1538,N_2088);
and U2999 (N_2999,N_1510,N_1609);
xnor U3000 (N_3000,N_2853,N_2495);
or U3001 (N_3001,N_2475,N_2644);
nand U3002 (N_3002,N_2604,N_2898);
nor U3003 (N_3003,N_2537,N_2378);
xor U3004 (N_3004,N_2479,N_2956);
nor U3005 (N_3005,N_2919,N_2271);
xor U3006 (N_3006,N_2549,N_2630);
nand U3007 (N_3007,N_2651,N_2995);
nor U3008 (N_3008,N_2424,N_2946);
or U3009 (N_3009,N_2838,N_2429);
and U3010 (N_3010,N_2509,N_2610);
and U3011 (N_3011,N_2771,N_2832);
xnor U3012 (N_3012,N_2453,N_2886);
and U3013 (N_3013,N_2804,N_2550);
or U3014 (N_3014,N_2326,N_2599);
nor U3015 (N_3015,N_2953,N_2904);
or U3016 (N_3016,N_2951,N_2837);
xnor U3017 (N_3017,N_2350,N_2680);
and U3018 (N_3018,N_2567,N_2615);
xnor U3019 (N_3019,N_2897,N_2278);
or U3020 (N_3020,N_2258,N_2583);
or U3021 (N_3021,N_2913,N_2260);
nand U3022 (N_3022,N_2961,N_2374);
or U3023 (N_3023,N_2557,N_2908);
nor U3024 (N_3024,N_2574,N_2686);
nor U3025 (N_3025,N_2456,N_2394);
nor U3026 (N_3026,N_2398,N_2872);
nand U3027 (N_3027,N_2367,N_2526);
and U3028 (N_3028,N_2609,N_2745);
nor U3029 (N_3029,N_2722,N_2347);
or U3030 (N_3030,N_2331,N_2314);
nor U3031 (N_3031,N_2750,N_2847);
or U3032 (N_3032,N_2380,N_2654);
nand U3033 (N_3033,N_2887,N_2994);
xor U3034 (N_3034,N_2282,N_2264);
or U3035 (N_3035,N_2540,N_2254);
or U3036 (N_3036,N_2877,N_2344);
nor U3037 (N_3037,N_2287,N_2524);
nor U3038 (N_3038,N_2998,N_2516);
nand U3039 (N_3039,N_2706,N_2581);
xor U3040 (N_3040,N_2856,N_2588);
xor U3041 (N_3041,N_2770,N_2551);
nand U3042 (N_3042,N_2738,N_2385);
or U3043 (N_3043,N_2922,N_2437);
nand U3044 (N_3044,N_2726,N_2859);
or U3045 (N_3045,N_2262,N_2703);
or U3046 (N_3046,N_2836,N_2596);
and U3047 (N_3047,N_2778,N_2642);
xor U3048 (N_3048,N_2755,N_2895);
xnor U3049 (N_3049,N_2957,N_2503);
xor U3050 (N_3050,N_2816,N_2619);
xor U3051 (N_3051,N_2341,N_2938);
nor U3052 (N_3052,N_2829,N_2334);
and U3053 (N_3053,N_2364,N_2692);
or U3054 (N_3054,N_2346,N_2512);
or U3055 (N_3055,N_2421,N_2677);
nand U3056 (N_3056,N_2869,N_2477);
xor U3057 (N_3057,N_2487,N_2308);
and U3058 (N_3058,N_2841,N_2404);
xnor U3059 (N_3059,N_2839,N_2284);
or U3060 (N_3060,N_2541,N_2565);
xnor U3061 (N_3061,N_2426,N_2389);
nor U3062 (N_3062,N_2656,N_2734);
nor U3063 (N_3063,N_2451,N_2452);
nor U3064 (N_3064,N_2330,N_2785);
xor U3065 (N_3065,N_2999,N_2440);
nor U3066 (N_3066,N_2365,N_2890);
nor U3067 (N_3067,N_2305,N_2562);
and U3068 (N_3068,N_2807,N_2593);
and U3069 (N_3069,N_2783,N_2940);
xnor U3070 (N_3070,N_2851,N_2301);
or U3071 (N_3071,N_2513,N_2587);
and U3072 (N_3072,N_2544,N_2405);
nand U3073 (N_3073,N_2658,N_2375);
xnor U3074 (N_3074,N_2752,N_2875);
and U3075 (N_3075,N_2844,N_2884);
nor U3076 (N_3076,N_2371,N_2276);
xor U3077 (N_3077,N_2339,N_2721);
nand U3078 (N_3078,N_2407,N_2580);
or U3079 (N_3079,N_2812,N_2473);
or U3080 (N_3080,N_2273,N_2775);
nor U3081 (N_3081,N_2834,N_2751);
or U3082 (N_3082,N_2962,N_2379);
nor U3083 (N_3083,N_2931,N_2607);
xor U3084 (N_3084,N_2799,N_2633);
nand U3085 (N_3085,N_2865,N_2942);
or U3086 (N_3086,N_2765,N_2848);
nor U3087 (N_3087,N_2514,N_2556);
nor U3088 (N_3088,N_2277,N_2930);
xor U3089 (N_3089,N_2650,N_2910);
nor U3090 (N_3090,N_2740,N_2422);
and U3091 (N_3091,N_2572,N_2489);
or U3092 (N_3092,N_2622,N_2434);
and U3093 (N_3093,N_2532,N_2854);
nand U3094 (N_3094,N_2470,N_2432);
nand U3095 (N_3095,N_2861,N_2723);
nor U3096 (N_3096,N_2693,N_2767);
nor U3097 (N_3097,N_2697,N_2779);
or U3098 (N_3098,N_2535,N_2830);
or U3099 (N_3099,N_2490,N_2678);
nand U3100 (N_3100,N_2733,N_2893);
and U3101 (N_3101,N_2529,N_2410);
and U3102 (N_3102,N_2705,N_2792);
or U3103 (N_3103,N_2253,N_2665);
nor U3104 (N_3104,N_2416,N_2757);
and U3105 (N_3105,N_2608,N_2283);
xnor U3106 (N_3106,N_2388,N_2794);
or U3107 (N_3107,N_2871,N_2618);
nor U3108 (N_3108,N_2261,N_2821);
xor U3109 (N_3109,N_2486,N_2924);
or U3110 (N_3110,N_2802,N_2760);
nor U3111 (N_3111,N_2846,N_2967);
nor U3112 (N_3112,N_2519,N_2787);
nand U3113 (N_3113,N_2579,N_2880);
and U3114 (N_3114,N_2554,N_2614);
nand U3115 (N_3115,N_2545,N_2517);
nor U3116 (N_3116,N_2510,N_2932);
xor U3117 (N_3117,N_2318,N_2840);
xnor U3118 (N_3118,N_2762,N_2307);
or U3119 (N_3119,N_2466,N_2891);
nand U3120 (N_3120,N_2270,N_2612);
nand U3121 (N_3121,N_2358,N_2862);
nand U3122 (N_3122,N_2643,N_2945);
nand U3123 (N_3123,N_2906,N_2742);
nor U3124 (N_3124,N_2605,N_2467);
and U3125 (N_3125,N_2590,N_2362);
nor U3126 (N_3126,N_2573,N_2555);
nor U3127 (N_3127,N_2559,N_2806);
nor U3128 (N_3128,N_2303,N_2496);
nor U3129 (N_3129,N_2764,N_2885);
or U3130 (N_3130,N_2417,N_2291);
nor U3131 (N_3131,N_2881,N_2427);
nand U3132 (N_3132,N_2298,N_2739);
nor U3133 (N_3133,N_2805,N_2329);
or U3134 (N_3134,N_2668,N_2639);
and U3135 (N_3135,N_2458,N_2664);
nor U3136 (N_3136,N_2297,N_2386);
nand U3137 (N_3137,N_2383,N_2809);
nor U3138 (N_3138,N_2800,N_2506);
nor U3139 (N_3139,N_2631,N_2731);
and U3140 (N_3140,N_2689,N_2585);
or U3141 (N_3141,N_2624,N_2568);
or U3142 (N_3142,N_2413,N_2718);
nor U3143 (N_3143,N_2813,N_2667);
or U3144 (N_3144,N_2707,N_2483);
and U3145 (N_3145,N_2373,N_2730);
nor U3146 (N_3146,N_2746,N_2634);
xor U3147 (N_3147,N_2719,N_2449);
or U3148 (N_3148,N_2657,N_2370);
or U3149 (N_3149,N_2876,N_2903);
nand U3150 (N_3150,N_2281,N_2533);
nand U3151 (N_3151,N_2300,N_2652);
and U3152 (N_3152,N_2336,N_2695);
xnor U3153 (N_3153,N_2469,N_2597);
and U3154 (N_3154,N_2814,N_2611);
xnor U3155 (N_3155,N_2754,N_2598);
nand U3156 (N_3156,N_2316,N_2811);
nor U3157 (N_3157,N_2338,N_2257);
or U3158 (N_3158,N_2737,N_2251);
xnor U3159 (N_3159,N_2729,N_2274);
nand U3160 (N_3160,N_2408,N_2553);
and U3161 (N_3161,N_2711,N_2396);
or U3162 (N_3162,N_2663,N_2543);
nor U3163 (N_3163,N_2603,N_2646);
xor U3164 (N_3164,N_2431,N_2672);
and U3165 (N_3165,N_2842,N_2858);
and U3166 (N_3166,N_2915,N_2454);
nand U3167 (N_3167,N_2947,N_2828);
nand U3168 (N_3168,N_2978,N_2632);
and U3169 (N_3169,N_2969,N_2402);
nand U3170 (N_3170,N_2337,N_2445);
nand U3171 (N_3171,N_2691,N_2638);
or U3172 (N_3172,N_2822,N_2296);
nand U3173 (N_3173,N_2295,N_2774);
nand U3174 (N_3174,N_2340,N_2860);
or U3175 (N_3175,N_2870,N_2833);
nor U3176 (N_3176,N_2332,N_2592);
nand U3177 (N_3177,N_2810,N_2661);
and U3178 (N_3178,N_2987,N_2328);
or U3179 (N_3179,N_2460,N_2481);
xor U3180 (N_3180,N_2763,N_2293);
or U3181 (N_3181,N_2977,N_2671);
xnor U3182 (N_3182,N_2419,N_2753);
xnor U3183 (N_3183,N_2289,N_2360);
xnor U3184 (N_3184,N_2527,N_2530);
and U3185 (N_3185,N_2361,N_2868);
or U3186 (N_3186,N_2323,N_2497);
xnor U3187 (N_3187,N_2867,N_2280);
and U3188 (N_3188,N_2436,N_2866);
and U3189 (N_3189,N_2443,N_2472);
and U3190 (N_3190,N_2521,N_2626);
nand U3191 (N_3191,N_2403,N_2925);
nand U3192 (N_3192,N_2768,N_2983);
or U3193 (N_3193,N_2928,N_2687);
or U3194 (N_3194,N_2500,N_2625);
nor U3195 (N_3195,N_2899,N_2259);
or U3196 (N_3196,N_2727,N_2879);
nand U3197 (N_3197,N_2666,N_2411);
or U3198 (N_3198,N_2493,N_2415);
nand U3199 (N_3199,N_2414,N_2351);
and U3200 (N_3200,N_2941,N_2345);
or U3201 (N_3201,N_2484,N_2462);
or U3202 (N_3202,N_2523,N_2476);
xnor U3203 (N_3203,N_2699,N_2474);
nor U3204 (N_3204,N_2704,N_2939);
and U3205 (N_3205,N_2918,N_2905);
and U3206 (N_3206,N_2439,N_2773);
nor U3207 (N_3207,N_2594,N_2744);
xor U3208 (N_3208,N_2935,N_2309);
nand U3209 (N_3209,N_2943,N_2808);
and U3210 (N_3210,N_2463,N_2892);
or U3211 (N_3211,N_2269,N_2628);
nand U3212 (N_3212,N_2465,N_2790);
nor U3213 (N_3213,N_2515,N_2522);
and U3214 (N_3214,N_2929,N_2902);
or U3215 (N_3215,N_2491,N_2640);
and U3216 (N_3216,N_2569,N_2675);
xnor U3217 (N_3217,N_2996,N_2570);
nor U3218 (N_3218,N_2252,N_2395);
or U3219 (N_3219,N_2412,N_2348);
nand U3220 (N_3220,N_2366,N_2578);
or U3221 (N_3221,N_2817,N_2818);
nor U3222 (N_3222,N_2505,N_2647);
nand U3223 (N_3223,N_2613,N_2717);
and U3224 (N_3224,N_2450,N_2965);
nor U3225 (N_3225,N_2724,N_2321);
and U3226 (N_3226,N_2747,N_2911);
xor U3227 (N_3227,N_2518,N_2782);
xor U3228 (N_3228,N_2715,N_2709);
xor U3229 (N_3229,N_2976,N_2606);
nand U3230 (N_3230,N_2425,N_2447);
and U3231 (N_3231,N_2835,N_2285);
nand U3232 (N_3232,N_2758,N_2485);
xor U3233 (N_3233,N_2420,N_2390);
xor U3234 (N_3234,N_2649,N_2448);
nor U3235 (N_3235,N_2888,N_2827);
or U3236 (N_3236,N_2315,N_2874);
nor U3237 (N_3237,N_2756,N_2279);
xor U3238 (N_3238,N_2688,N_2552);
or U3239 (N_3239,N_2438,N_2302);
nand U3240 (N_3240,N_2914,N_2982);
xnor U3241 (N_3241,N_2531,N_2972);
xor U3242 (N_3242,N_2777,N_2442);
nand U3243 (N_3243,N_2849,N_2561);
xor U3244 (N_3244,N_2542,N_2327);
or U3245 (N_3245,N_2979,N_2716);
or U3246 (N_3246,N_2966,N_2560);
or U3247 (N_3247,N_2852,N_2363);
and U3248 (N_3248,N_2660,N_2992);
nor U3249 (N_3249,N_2268,N_2850);
nor U3250 (N_3250,N_2873,N_2907);
xnor U3251 (N_3251,N_2710,N_2823);
or U3252 (N_3252,N_2648,N_2418);
nor U3253 (N_3253,N_2662,N_2728);
nor U3254 (N_3254,N_2937,N_2256);
xnor U3255 (N_3255,N_2312,N_2824);
xnor U3256 (N_3256,N_2894,N_2798);
nand U3257 (N_3257,N_2698,N_2968);
or U3258 (N_3258,N_2571,N_2319);
xnor U3259 (N_3259,N_2306,N_2653);
nand U3260 (N_3260,N_2714,N_2955);
nand U3261 (N_3261,N_2589,N_2320);
or U3262 (N_3262,N_2669,N_2355);
xnor U3263 (N_3263,N_2696,N_2989);
or U3264 (N_3264,N_2720,N_2934);
and U3265 (N_3265,N_2399,N_2973);
or U3266 (N_3266,N_2255,N_2288);
nor U3267 (N_3267,N_2324,N_2793);
nor U3268 (N_3268,N_2499,N_2801);
nor U3269 (N_3269,N_2674,N_2952);
nand U3270 (N_3270,N_2304,N_2936);
xnor U3271 (N_3271,N_2901,N_2963);
and U3272 (N_3272,N_2455,N_2636);
and U3273 (N_3273,N_2681,N_2325);
and U3274 (N_3274,N_2769,N_2641);
xnor U3275 (N_3275,N_2595,N_2993);
and U3276 (N_3276,N_2926,N_2343);
xor U3277 (N_3277,N_2392,N_2815);
nand U3278 (N_3278,N_2921,N_2525);
nor U3279 (N_3279,N_2786,N_2317);
xor U3280 (N_3280,N_2444,N_2310);
nor U3281 (N_3281,N_2601,N_2423);
and U3282 (N_3282,N_2701,N_2984);
nor U3283 (N_3283,N_2685,N_2912);
nor U3284 (N_3284,N_2397,N_2735);
nand U3285 (N_3285,N_2428,N_2508);
nor U3286 (N_3286,N_2393,N_2292);
xor U3287 (N_3287,N_2974,N_2272);
nand U3288 (N_3288,N_2534,N_2960);
and U3289 (N_3289,N_2250,N_2520);
and U3290 (N_3290,N_2311,N_2547);
nor U3291 (N_3291,N_2882,N_2795);
nor U3292 (N_3292,N_2819,N_2864);
and U3293 (N_3293,N_2975,N_2863);
and U3294 (N_3294,N_2369,N_2825);
nand U3295 (N_3295,N_2637,N_2602);
and U3296 (N_3296,N_2743,N_2382);
or U3297 (N_3297,N_2948,N_2673);
or U3298 (N_3298,N_2927,N_2684);
and U3299 (N_3299,N_2826,N_2629);
nand U3300 (N_3300,N_2539,N_2725);
and U3301 (N_3301,N_2528,N_2435);
nor U3302 (N_3302,N_2889,N_2676);
xnor U3303 (N_3303,N_2635,N_2997);
nor U3304 (N_3304,N_2409,N_2920);
or U3305 (N_3305,N_2909,N_2796);
nand U3306 (N_3306,N_2488,N_2381);
nor U3307 (N_3307,N_2275,N_2538);
and U3308 (N_3308,N_2845,N_2857);
nand U3309 (N_3309,N_2883,N_2576);
or U3310 (N_3310,N_2313,N_2694);
and U3311 (N_3311,N_2878,N_2659);
xnor U3312 (N_3312,N_2356,N_2492);
or U3313 (N_3313,N_2406,N_2501);
xor U3314 (N_3314,N_2563,N_2267);
and U3315 (N_3315,N_2788,N_2981);
nor U3316 (N_3316,N_2843,N_2349);
xor U3317 (N_3317,N_2917,N_2988);
and U3318 (N_3318,N_2781,N_2504);
or U3319 (N_3319,N_2372,N_2482);
nor U3320 (N_3320,N_2708,N_2645);
or U3321 (N_3321,N_2780,N_2461);
and U3322 (N_3322,N_2376,N_2964);
xnor U3323 (N_3323,N_2991,N_2971);
xor U3324 (N_3324,N_2582,N_2958);
nand U3325 (N_3325,N_2368,N_2584);
xor U3326 (N_3326,N_2335,N_2294);
and U3327 (N_3327,N_2591,N_2950);
and U3328 (N_3328,N_2690,N_2949);
nor U3329 (N_3329,N_2655,N_2400);
or U3330 (N_3330,N_2498,N_2749);
or U3331 (N_3331,N_2357,N_2621);
or U3332 (N_3332,N_2970,N_2766);
and U3333 (N_3333,N_2401,N_2468);
nand U3334 (N_3334,N_2457,N_2617);
nor U3335 (N_3335,N_2577,N_2430);
xor U3336 (N_3336,N_2713,N_2916);
xor U3337 (N_3337,N_2441,N_2679);
nor U3338 (N_3338,N_2494,N_2536);
nand U3339 (N_3339,N_2748,N_2923);
or U3340 (N_3340,N_2265,N_2712);
or U3341 (N_3341,N_2896,N_2627);
xnor U3342 (N_3342,N_2616,N_2575);
xor U3343 (N_3343,N_2286,N_2464);
xnor U3344 (N_3344,N_2831,N_2959);
or U3345 (N_3345,N_2342,N_2359);
nand U3346 (N_3346,N_2741,N_2290);
and U3347 (N_3347,N_2263,N_2511);
and U3348 (N_3348,N_2784,N_2702);
xnor U3349 (N_3349,N_2558,N_2759);
or U3350 (N_3350,N_2507,N_2564);
and U3351 (N_3351,N_2322,N_2546);
or U3352 (N_3352,N_2954,N_2985);
xor U3353 (N_3353,N_2944,N_2682);
nand U3354 (N_3354,N_2480,N_2586);
nor U3355 (N_3355,N_2736,N_2820);
nor U3356 (N_3356,N_2670,N_2266);
nand U3357 (N_3357,N_2446,N_2761);
nor U3358 (N_3358,N_2700,N_2789);
or U3359 (N_3359,N_2377,N_2352);
nand U3360 (N_3360,N_2986,N_2548);
nor U3361 (N_3361,N_2459,N_2354);
and U3362 (N_3362,N_2391,N_2803);
xor U3363 (N_3363,N_2502,N_2933);
and U3364 (N_3364,N_2478,N_2471);
nor U3365 (N_3365,N_2732,N_2353);
nor U3366 (N_3366,N_2566,N_2776);
nand U3367 (N_3367,N_2791,N_2387);
nand U3368 (N_3368,N_2384,N_2990);
xnor U3369 (N_3369,N_2980,N_2433);
or U3370 (N_3370,N_2855,N_2683);
xnor U3371 (N_3371,N_2900,N_2600);
and U3372 (N_3372,N_2797,N_2299);
xor U3373 (N_3373,N_2620,N_2772);
and U3374 (N_3374,N_2333,N_2623);
nor U3375 (N_3375,N_2657,N_2251);
and U3376 (N_3376,N_2446,N_2570);
nand U3377 (N_3377,N_2701,N_2932);
or U3378 (N_3378,N_2906,N_2292);
or U3379 (N_3379,N_2882,N_2525);
or U3380 (N_3380,N_2625,N_2277);
xor U3381 (N_3381,N_2941,N_2253);
nor U3382 (N_3382,N_2327,N_2800);
and U3383 (N_3383,N_2667,N_2798);
xnor U3384 (N_3384,N_2801,N_2570);
or U3385 (N_3385,N_2939,N_2741);
nor U3386 (N_3386,N_2380,N_2872);
nand U3387 (N_3387,N_2881,N_2819);
xnor U3388 (N_3388,N_2263,N_2483);
or U3389 (N_3389,N_2716,N_2727);
xor U3390 (N_3390,N_2353,N_2461);
nor U3391 (N_3391,N_2739,N_2262);
and U3392 (N_3392,N_2722,N_2827);
nand U3393 (N_3393,N_2845,N_2746);
and U3394 (N_3394,N_2608,N_2595);
nor U3395 (N_3395,N_2814,N_2276);
xor U3396 (N_3396,N_2410,N_2706);
xor U3397 (N_3397,N_2572,N_2422);
nor U3398 (N_3398,N_2503,N_2852);
or U3399 (N_3399,N_2727,N_2351);
and U3400 (N_3400,N_2968,N_2655);
or U3401 (N_3401,N_2253,N_2287);
nor U3402 (N_3402,N_2920,N_2848);
nand U3403 (N_3403,N_2397,N_2652);
nand U3404 (N_3404,N_2775,N_2655);
xor U3405 (N_3405,N_2435,N_2694);
and U3406 (N_3406,N_2445,N_2622);
xnor U3407 (N_3407,N_2788,N_2488);
nor U3408 (N_3408,N_2326,N_2888);
xor U3409 (N_3409,N_2443,N_2889);
nand U3410 (N_3410,N_2934,N_2388);
and U3411 (N_3411,N_2489,N_2415);
xnor U3412 (N_3412,N_2654,N_2334);
xnor U3413 (N_3413,N_2473,N_2956);
nor U3414 (N_3414,N_2760,N_2996);
nand U3415 (N_3415,N_2714,N_2849);
xnor U3416 (N_3416,N_2343,N_2381);
nand U3417 (N_3417,N_2833,N_2606);
xor U3418 (N_3418,N_2690,N_2744);
nand U3419 (N_3419,N_2378,N_2352);
and U3420 (N_3420,N_2467,N_2640);
nor U3421 (N_3421,N_2605,N_2849);
and U3422 (N_3422,N_2673,N_2343);
or U3423 (N_3423,N_2669,N_2828);
xnor U3424 (N_3424,N_2639,N_2767);
nand U3425 (N_3425,N_2253,N_2970);
and U3426 (N_3426,N_2667,N_2514);
and U3427 (N_3427,N_2269,N_2524);
xnor U3428 (N_3428,N_2256,N_2729);
nand U3429 (N_3429,N_2992,N_2937);
nand U3430 (N_3430,N_2742,N_2881);
nand U3431 (N_3431,N_2809,N_2569);
nor U3432 (N_3432,N_2531,N_2314);
and U3433 (N_3433,N_2930,N_2967);
nor U3434 (N_3434,N_2335,N_2782);
nand U3435 (N_3435,N_2781,N_2818);
nor U3436 (N_3436,N_2981,N_2834);
xor U3437 (N_3437,N_2807,N_2655);
nand U3438 (N_3438,N_2563,N_2658);
nand U3439 (N_3439,N_2279,N_2694);
and U3440 (N_3440,N_2811,N_2601);
nand U3441 (N_3441,N_2483,N_2350);
nand U3442 (N_3442,N_2474,N_2299);
xor U3443 (N_3443,N_2321,N_2684);
nor U3444 (N_3444,N_2699,N_2941);
or U3445 (N_3445,N_2820,N_2726);
and U3446 (N_3446,N_2481,N_2803);
xnor U3447 (N_3447,N_2595,N_2362);
and U3448 (N_3448,N_2738,N_2892);
and U3449 (N_3449,N_2714,N_2646);
and U3450 (N_3450,N_2342,N_2770);
nand U3451 (N_3451,N_2780,N_2837);
nand U3452 (N_3452,N_2283,N_2649);
or U3453 (N_3453,N_2443,N_2662);
or U3454 (N_3454,N_2696,N_2451);
nor U3455 (N_3455,N_2559,N_2713);
nor U3456 (N_3456,N_2579,N_2273);
xor U3457 (N_3457,N_2983,N_2907);
and U3458 (N_3458,N_2860,N_2563);
or U3459 (N_3459,N_2442,N_2540);
and U3460 (N_3460,N_2360,N_2730);
xor U3461 (N_3461,N_2504,N_2985);
xor U3462 (N_3462,N_2631,N_2341);
or U3463 (N_3463,N_2577,N_2429);
or U3464 (N_3464,N_2342,N_2698);
or U3465 (N_3465,N_2303,N_2534);
nand U3466 (N_3466,N_2412,N_2855);
nor U3467 (N_3467,N_2827,N_2594);
nor U3468 (N_3468,N_2534,N_2633);
and U3469 (N_3469,N_2486,N_2645);
nor U3470 (N_3470,N_2499,N_2427);
nor U3471 (N_3471,N_2977,N_2287);
xor U3472 (N_3472,N_2478,N_2580);
xor U3473 (N_3473,N_2578,N_2736);
nor U3474 (N_3474,N_2304,N_2536);
nor U3475 (N_3475,N_2552,N_2828);
nand U3476 (N_3476,N_2723,N_2762);
nand U3477 (N_3477,N_2506,N_2988);
nor U3478 (N_3478,N_2999,N_2821);
and U3479 (N_3479,N_2297,N_2705);
nand U3480 (N_3480,N_2293,N_2430);
nor U3481 (N_3481,N_2627,N_2682);
xnor U3482 (N_3482,N_2273,N_2705);
or U3483 (N_3483,N_2608,N_2313);
xnor U3484 (N_3484,N_2574,N_2423);
xor U3485 (N_3485,N_2588,N_2547);
xor U3486 (N_3486,N_2585,N_2358);
and U3487 (N_3487,N_2638,N_2813);
or U3488 (N_3488,N_2482,N_2874);
or U3489 (N_3489,N_2376,N_2390);
and U3490 (N_3490,N_2260,N_2948);
nand U3491 (N_3491,N_2816,N_2738);
nor U3492 (N_3492,N_2520,N_2883);
xor U3493 (N_3493,N_2299,N_2575);
nand U3494 (N_3494,N_2583,N_2959);
nand U3495 (N_3495,N_2918,N_2641);
nand U3496 (N_3496,N_2433,N_2810);
and U3497 (N_3497,N_2553,N_2630);
and U3498 (N_3498,N_2758,N_2373);
nor U3499 (N_3499,N_2665,N_2639);
or U3500 (N_3500,N_2441,N_2937);
nor U3501 (N_3501,N_2932,N_2680);
or U3502 (N_3502,N_2363,N_2787);
or U3503 (N_3503,N_2723,N_2523);
xnor U3504 (N_3504,N_2731,N_2467);
and U3505 (N_3505,N_2282,N_2275);
or U3506 (N_3506,N_2807,N_2561);
and U3507 (N_3507,N_2602,N_2472);
nand U3508 (N_3508,N_2495,N_2428);
xnor U3509 (N_3509,N_2849,N_2595);
or U3510 (N_3510,N_2340,N_2575);
xor U3511 (N_3511,N_2666,N_2970);
and U3512 (N_3512,N_2273,N_2823);
xor U3513 (N_3513,N_2313,N_2427);
nand U3514 (N_3514,N_2930,N_2831);
and U3515 (N_3515,N_2981,N_2877);
nand U3516 (N_3516,N_2712,N_2795);
or U3517 (N_3517,N_2889,N_2380);
xor U3518 (N_3518,N_2933,N_2803);
nor U3519 (N_3519,N_2350,N_2711);
or U3520 (N_3520,N_2359,N_2893);
nand U3521 (N_3521,N_2803,N_2395);
or U3522 (N_3522,N_2754,N_2971);
and U3523 (N_3523,N_2775,N_2286);
xor U3524 (N_3524,N_2987,N_2618);
or U3525 (N_3525,N_2688,N_2968);
nor U3526 (N_3526,N_2416,N_2627);
and U3527 (N_3527,N_2889,N_2973);
nor U3528 (N_3528,N_2902,N_2685);
and U3529 (N_3529,N_2638,N_2467);
nor U3530 (N_3530,N_2805,N_2464);
nor U3531 (N_3531,N_2830,N_2593);
or U3532 (N_3532,N_2753,N_2381);
and U3533 (N_3533,N_2465,N_2580);
xor U3534 (N_3534,N_2322,N_2353);
nand U3535 (N_3535,N_2807,N_2632);
xnor U3536 (N_3536,N_2443,N_2968);
xnor U3537 (N_3537,N_2735,N_2260);
and U3538 (N_3538,N_2260,N_2413);
nand U3539 (N_3539,N_2360,N_2857);
nand U3540 (N_3540,N_2287,N_2486);
or U3541 (N_3541,N_2403,N_2735);
xor U3542 (N_3542,N_2894,N_2694);
xor U3543 (N_3543,N_2868,N_2982);
and U3544 (N_3544,N_2580,N_2571);
nor U3545 (N_3545,N_2470,N_2626);
xnor U3546 (N_3546,N_2404,N_2304);
nand U3547 (N_3547,N_2560,N_2561);
and U3548 (N_3548,N_2271,N_2800);
or U3549 (N_3549,N_2540,N_2884);
nor U3550 (N_3550,N_2805,N_2553);
nand U3551 (N_3551,N_2765,N_2907);
nand U3552 (N_3552,N_2640,N_2295);
nor U3553 (N_3553,N_2760,N_2797);
xnor U3554 (N_3554,N_2555,N_2982);
and U3555 (N_3555,N_2516,N_2977);
xor U3556 (N_3556,N_2373,N_2993);
nand U3557 (N_3557,N_2341,N_2399);
and U3558 (N_3558,N_2698,N_2597);
and U3559 (N_3559,N_2560,N_2786);
nor U3560 (N_3560,N_2690,N_2420);
and U3561 (N_3561,N_2465,N_2344);
xor U3562 (N_3562,N_2590,N_2545);
nor U3563 (N_3563,N_2786,N_2513);
xnor U3564 (N_3564,N_2721,N_2894);
nand U3565 (N_3565,N_2698,N_2387);
nor U3566 (N_3566,N_2922,N_2790);
or U3567 (N_3567,N_2834,N_2918);
xnor U3568 (N_3568,N_2703,N_2278);
nor U3569 (N_3569,N_2268,N_2689);
nand U3570 (N_3570,N_2690,N_2349);
nand U3571 (N_3571,N_2531,N_2832);
nor U3572 (N_3572,N_2713,N_2781);
or U3573 (N_3573,N_2882,N_2655);
nor U3574 (N_3574,N_2941,N_2899);
and U3575 (N_3575,N_2892,N_2413);
or U3576 (N_3576,N_2836,N_2445);
nor U3577 (N_3577,N_2630,N_2530);
nand U3578 (N_3578,N_2838,N_2378);
nand U3579 (N_3579,N_2504,N_2452);
or U3580 (N_3580,N_2497,N_2256);
xor U3581 (N_3581,N_2514,N_2916);
xnor U3582 (N_3582,N_2927,N_2468);
xnor U3583 (N_3583,N_2737,N_2770);
and U3584 (N_3584,N_2659,N_2413);
nor U3585 (N_3585,N_2813,N_2437);
or U3586 (N_3586,N_2653,N_2470);
nor U3587 (N_3587,N_2659,N_2956);
and U3588 (N_3588,N_2735,N_2875);
or U3589 (N_3589,N_2252,N_2942);
nor U3590 (N_3590,N_2467,N_2808);
xnor U3591 (N_3591,N_2845,N_2749);
and U3592 (N_3592,N_2510,N_2252);
nor U3593 (N_3593,N_2562,N_2822);
nand U3594 (N_3594,N_2500,N_2541);
nand U3595 (N_3595,N_2792,N_2462);
xnor U3596 (N_3596,N_2438,N_2990);
nor U3597 (N_3597,N_2506,N_2709);
nor U3598 (N_3598,N_2485,N_2916);
or U3599 (N_3599,N_2505,N_2332);
nand U3600 (N_3600,N_2507,N_2786);
and U3601 (N_3601,N_2308,N_2656);
and U3602 (N_3602,N_2936,N_2986);
nand U3603 (N_3603,N_2550,N_2988);
nor U3604 (N_3604,N_2343,N_2994);
nor U3605 (N_3605,N_2410,N_2948);
and U3606 (N_3606,N_2793,N_2548);
nand U3607 (N_3607,N_2652,N_2518);
or U3608 (N_3608,N_2781,N_2588);
nor U3609 (N_3609,N_2497,N_2945);
nand U3610 (N_3610,N_2740,N_2535);
nor U3611 (N_3611,N_2751,N_2892);
nor U3612 (N_3612,N_2517,N_2729);
and U3613 (N_3613,N_2529,N_2284);
and U3614 (N_3614,N_2896,N_2897);
or U3615 (N_3615,N_2870,N_2963);
xor U3616 (N_3616,N_2950,N_2593);
and U3617 (N_3617,N_2439,N_2285);
nand U3618 (N_3618,N_2668,N_2715);
nand U3619 (N_3619,N_2400,N_2577);
and U3620 (N_3620,N_2999,N_2601);
nor U3621 (N_3621,N_2552,N_2859);
nand U3622 (N_3622,N_2614,N_2992);
or U3623 (N_3623,N_2475,N_2499);
xor U3624 (N_3624,N_2969,N_2545);
nand U3625 (N_3625,N_2771,N_2363);
nand U3626 (N_3626,N_2632,N_2890);
and U3627 (N_3627,N_2324,N_2963);
and U3628 (N_3628,N_2389,N_2404);
or U3629 (N_3629,N_2511,N_2726);
or U3630 (N_3630,N_2910,N_2667);
nor U3631 (N_3631,N_2893,N_2501);
nand U3632 (N_3632,N_2310,N_2656);
and U3633 (N_3633,N_2329,N_2981);
xnor U3634 (N_3634,N_2715,N_2411);
and U3635 (N_3635,N_2856,N_2725);
nor U3636 (N_3636,N_2798,N_2636);
xor U3637 (N_3637,N_2745,N_2856);
nand U3638 (N_3638,N_2561,N_2673);
nor U3639 (N_3639,N_2436,N_2293);
xnor U3640 (N_3640,N_2652,N_2594);
nand U3641 (N_3641,N_2373,N_2434);
nor U3642 (N_3642,N_2812,N_2499);
nor U3643 (N_3643,N_2666,N_2551);
or U3644 (N_3644,N_2739,N_2445);
nand U3645 (N_3645,N_2824,N_2537);
xor U3646 (N_3646,N_2289,N_2651);
nor U3647 (N_3647,N_2865,N_2846);
or U3648 (N_3648,N_2563,N_2318);
and U3649 (N_3649,N_2470,N_2790);
or U3650 (N_3650,N_2419,N_2644);
or U3651 (N_3651,N_2370,N_2550);
and U3652 (N_3652,N_2851,N_2591);
and U3653 (N_3653,N_2920,N_2288);
nor U3654 (N_3654,N_2732,N_2518);
and U3655 (N_3655,N_2536,N_2275);
xor U3656 (N_3656,N_2273,N_2599);
or U3657 (N_3657,N_2920,N_2660);
nand U3658 (N_3658,N_2738,N_2608);
nor U3659 (N_3659,N_2910,N_2737);
and U3660 (N_3660,N_2542,N_2836);
and U3661 (N_3661,N_2901,N_2915);
xnor U3662 (N_3662,N_2918,N_2890);
nand U3663 (N_3663,N_2294,N_2325);
and U3664 (N_3664,N_2877,N_2566);
xnor U3665 (N_3665,N_2832,N_2352);
nor U3666 (N_3666,N_2459,N_2616);
nand U3667 (N_3667,N_2580,N_2777);
or U3668 (N_3668,N_2846,N_2363);
nor U3669 (N_3669,N_2915,N_2823);
and U3670 (N_3670,N_2391,N_2410);
nand U3671 (N_3671,N_2676,N_2368);
and U3672 (N_3672,N_2282,N_2656);
or U3673 (N_3673,N_2896,N_2725);
or U3674 (N_3674,N_2736,N_2922);
nor U3675 (N_3675,N_2950,N_2841);
and U3676 (N_3676,N_2663,N_2844);
nor U3677 (N_3677,N_2663,N_2546);
xor U3678 (N_3678,N_2493,N_2982);
nor U3679 (N_3679,N_2936,N_2739);
nand U3680 (N_3680,N_2516,N_2957);
nor U3681 (N_3681,N_2287,N_2912);
and U3682 (N_3682,N_2299,N_2899);
or U3683 (N_3683,N_2527,N_2572);
and U3684 (N_3684,N_2632,N_2863);
xnor U3685 (N_3685,N_2835,N_2341);
nor U3686 (N_3686,N_2987,N_2294);
or U3687 (N_3687,N_2879,N_2699);
xor U3688 (N_3688,N_2548,N_2691);
xnor U3689 (N_3689,N_2262,N_2841);
xnor U3690 (N_3690,N_2885,N_2401);
xnor U3691 (N_3691,N_2297,N_2463);
and U3692 (N_3692,N_2482,N_2673);
nor U3693 (N_3693,N_2685,N_2532);
or U3694 (N_3694,N_2332,N_2637);
nor U3695 (N_3695,N_2837,N_2330);
xnor U3696 (N_3696,N_2654,N_2779);
or U3697 (N_3697,N_2543,N_2273);
or U3698 (N_3698,N_2436,N_2940);
nand U3699 (N_3699,N_2372,N_2264);
nor U3700 (N_3700,N_2803,N_2593);
nand U3701 (N_3701,N_2822,N_2718);
nor U3702 (N_3702,N_2292,N_2901);
or U3703 (N_3703,N_2779,N_2509);
nand U3704 (N_3704,N_2918,N_2973);
and U3705 (N_3705,N_2488,N_2609);
and U3706 (N_3706,N_2764,N_2449);
nor U3707 (N_3707,N_2360,N_2287);
and U3708 (N_3708,N_2806,N_2777);
or U3709 (N_3709,N_2398,N_2607);
and U3710 (N_3710,N_2975,N_2410);
nand U3711 (N_3711,N_2317,N_2572);
xor U3712 (N_3712,N_2457,N_2382);
or U3713 (N_3713,N_2894,N_2572);
nor U3714 (N_3714,N_2931,N_2724);
xor U3715 (N_3715,N_2347,N_2732);
nand U3716 (N_3716,N_2831,N_2419);
or U3717 (N_3717,N_2347,N_2604);
xnor U3718 (N_3718,N_2690,N_2724);
nor U3719 (N_3719,N_2970,N_2954);
nand U3720 (N_3720,N_2292,N_2423);
or U3721 (N_3721,N_2309,N_2445);
and U3722 (N_3722,N_2456,N_2694);
or U3723 (N_3723,N_2745,N_2664);
nand U3724 (N_3724,N_2597,N_2830);
nand U3725 (N_3725,N_2801,N_2296);
xnor U3726 (N_3726,N_2252,N_2310);
nor U3727 (N_3727,N_2300,N_2691);
nand U3728 (N_3728,N_2541,N_2580);
xor U3729 (N_3729,N_2339,N_2839);
xnor U3730 (N_3730,N_2691,N_2433);
or U3731 (N_3731,N_2487,N_2323);
nand U3732 (N_3732,N_2298,N_2398);
nand U3733 (N_3733,N_2495,N_2728);
or U3734 (N_3734,N_2367,N_2779);
or U3735 (N_3735,N_2683,N_2767);
and U3736 (N_3736,N_2360,N_2791);
nor U3737 (N_3737,N_2822,N_2543);
and U3738 (N_3738,N_2856,N_2558);
and U3739 (N_3739,N_2273,N_2651);
nor U3740 (N_3740,N_2421,N_2564);
and U3741 (N_3741,N_2733,N_2807);
or U3742 (N_3742,N_2664,N_2536);
and U3743 (N_3743,N_2501,N_2688);
nand U3744 (N_3744,N_2605,N_2859);
nor U3745 (N_3745,N_2327,N_2622);
and U3746 (N_3746,N_2435,N_2646);
nor U3747 (N_3747,N_2971,N_2250);
xor U3748 (N_3748,N_2627,N_2688);
and U3749 (N_3749,N_2729,N_2526);
nor U3750 (N_3750,N_3689,N_3311);
nand U3751 (N_3751,N_3151,N_3411);
nand U3752 (N_3752,N_3699,N_3389);
and U3753 (N_3753,N_3108,N_3303);
and U3754 (N_3754,N_3336,N_3348);
xor U3755 (N_3755,N_3481,N_3164);
xnor U3756 (N_3756,N_3667,N_3593);
xnor U3757 (N_3757,N_3557,N_3673);
xnor U3758 (N_3758,N_3437,N_3296);
nand U3759 (N_3759,N_3020,N_3726);
nand U3760 (N_3760,N_3721,N_3188);
xnor U3761 (N_3761,N_3310,N_3200);
and U3762 (N_3762,N_3217,N_3220);
or U3763 (N_3763,N_3376,N_3226);
xor U3764 (N_3764,N_3280,N_3459);
nor U3765 (N_3765,N_3306,N_3498);
nand U3766 (N_3766,N_3416,N_3566);
or U3767 (N_3767,N_3021,N_3698);
nor U3768 (N_3768,N_3506,N_3493);
nand U3769 (N_3769,N_3354,N_3187);
nor U3770 (N_3770,N_3583,N_3071);
xor U3771 (N_3771,N_3167,N_3214);
nor U3772 (N_3772,N_3251,N_3610);
or U3773 (N_3773,N_3120,N_3049);
xor U3774 (N_3774,N_3160,N_3588);
or U3775 (N_3775,N_3561,N_3028);
nor U3776 (N_3776,N_3736,N_3706);
and U3777 (N_3777,N_3563,N_3009);
nand U3778 (N_3778,N_3692,N_3714);
xor U3779 (N_3779,N_3138,N_3513);
nor U3780 (N_3780,N_3109,N_3095);
or U3781 (N_3781,N_3398,N_3162);
and U3782 (N_3782,N_3539,N_3479);
xnor U3783 (N_3783,N_3036,N_3233);
or U3784 (N_3784,N_3700,N_3456);
nor U3785 (N_3785,N_3397,N_3207);
and U3786 (N_3786,N_3253,N_3205);
xnor U3787 (N_3787,N_3068,N_3367);
and U3788 (N_3788,N_3345,N_3744);
and U3789 (N_3789,N_3091,N_3551);
nand U3790 (N_3790,N_3150,N_3523);
nand U3791 (N_3791,N_3299,N_3648);
nand U3792 (N_3792,N_3055,N_3461);
nor U3793 (N_3793,N_3022,N_3199);
xor U3794 (N_3794,N_3618,N_3453);
nor U3795 (N_3795,N_3635,N_3050);
and U3796 (N_3796,N_3438,N_3460);
and U3797 (N_3797,N_3037,N_3595);
and U3798 (N_3798,N_3391,N_3381);
xor U3799 (N_3799,N_3195,N_3190);
and U3800 (N_3800,N_3653,N_3155);
or U3801 (N_3801,N_3284,N_3517);
nand U3802 (N_3802,N_3556,N_3218);
xnor U3803 (N_3803,N_3526,N_3173);
xnor U3804 (N_3804,N_3156,N_3603);
nor U3805 (N_3805,N_3185,N_3463);
nor U3806 (N_3806,N_3694,N_3685);
or U3807 (N_3807,N_3027,N_3549);
or U3808 (N_3808,N_3419,N_3269);
and U3809 (N_3809,N_3198,N_3257);
or U3810 (N_3810,N_3490,N_3112);
xor U3811 (N_3811,N_3208,N_3383);
xnor U3812 (N_3812,N_3740,N_3168);
and U3813 (N_3813,N_3728,N_3647);
nor U3814 (N_3814,N_3633,N_3450);
nor U3815 (N_3815,N_3682,N_3090);
and U3816 (N_3816,N_3626,N_3040);
nor U3817 (N_3817,N_3165,N_3189);
or U3818 (N_3818,N_3123,N_3402);
nor U3819 (N_3819,N_3237,N_3042);
nand U3820 (N_3820,N_3489,N_3430);
nand U3821 (N_3821,N_3136,N_3514);
or U3822 (N_3822,N_3007,N_3606);
and U3823 (N_3823,N_3175,N_3325);
nor U3824 (N_3824,N_3641,N_3079);
xor U3825 (N_3825,N_3148,N_3576);
or U3826 (N_3826,N_3536,N_3425);
nand U3827 (N_3827,N_3743,N_3435);
xnor U3828 (N_3828,N_3439,N_3312);
and U3829 (N_3829,N_3403,N_3033);
or U3830 (N_3830,N_3255,N_3114);
nor U3831 (N_3831,N_3562,N_3624);
xnor U3832 (N_3832,N_3720,N_3180);
and U3833 (N_3833,N_3605,N_3627);
nand U3834 (N_3834,N_3695,N_3361);
or U3835 (N_3835,N_3067,N_3103);
nand U3836 (N_3836,N_3451,N_3204);
or U3837 (N_3837,N_3745,N_3322);
and U3838 (N_3838,N_3072,N_3659);
nor U3839 (N_3839,N_3499,N_3182);
or U3840 (N_3840,N_3572,N_3666);
nand U3841 (N_3841,N_3056,N_3192);
nor U3842 (N_3842,N_3544,N_3238);
and U3843 (N_3843,N_3739,N_3340);
nor U3844 (N_3844,N_3053,N_3116);
and U3845 (N_3845,N_3107,N_3362);
xnor U3846 (N_3846,N_3410,N_3476);
and U3847 (N_3847,N_3283,N_3552);
nor U3848 (N_3848,N_3297,N_3289);
and U3849 (N_3849,N_3330,N_3343);
xnor U3850 (N_3850,N_3074,N_3111);
nand U3851 (N_3851,N_3276,N_3528);
or U3852 (N_3852,N_3708,N_3623);
nor U3853 (N_3853,N_3683,N_3326);
nand U3854 (N_3854,N_3084,N_3329);
and U3855 (N_3855,N_3351,N_3130);
or U3856 (N_3856,N_3527,N_3712);
nand U3857 (N_3857,N_3599,N_3270);
nor U3858 (N_3858,N_3719,N_3742);
and U3859 (N_3859,N_3632,N_3678);
xnor U3860 (N_3860,N_3124,N_3664);
or U3861 (N_3861,N_3424,N_3364);
nand U3862 (N_3862,N_3365,N_3069);
or U3863 (N_3863,N_3333,N_3203);
nor U3864 (N_3864,N_3738,N_3570);
nand U3865 (N_3865,N_3642,N_3224);
and U3866 (N_3866,N_3015,N_3387);
or U3867 (N_3867,N_3581,N_3426);
and U3868 (N_3868,N_3264,N_3480);
or U3869 (N_3869,N_3206,N_3619);
nand U3870 (N_3870,N_3656,N_3702);
or U3871 (N_3871,N_3250,N_3645);
xor U3872 (N_3872,N_3468,N_3375);
or U3873 (N_3873,N_3675,N_3510);
nor U3874 (N_3874,N_3186,N_3637);
nand U3875 (N_3875,N_3129,N_3670);
xnor U3876 (N_3876,N_3302,N_3414);
nand U3877 (N_3877,N_3152,N_3620);
nor U3878 (N_3878,N_3134,N_3242);
xor U3879 (N_3879,N_3234,N_3500);
xor U3880 (N_3880,N_3611,N_3677);
xor U3881 (N_3881,N_3540,N_3693);
nor U3882 (N_3882,N_3569,N_3530);
nor U3883 (N_3883,N_3607,N_3229);
nor U3884 (N_3884,N_3358,N_3535);
nand U3885 (N_3885,N_3550,N_3448);
nor U3886 (N_3886,N_3723,N_3013);
nor U3887 (N_3887,N_3121,N_3184);
xnor U3888 (N_3888,N_3105,N_3406);
and U3889 (N_3889,N_3650,N_3469);
nand U3890 (N_3890,N_3082,N_3057);
xnor U3891 (N_3891,N_3147,N_3665);
nor U3892 (N_3892,N_3118,N_3360);
or U3893 (N_3893,N_3286,N_3249);
nand U3894 (N_3894,N_3625,N_3290);
xor U3895 (N_3895,N_3711,N_3565);
or U3896 (N_3896,N_3405,N_3212);
xnor U3897 (N_3897,N_3163,N_3559);
nand U3898 (N_3898,N_3592,N_3341);
or U3899 (N_3899,N_3386,N_3433);
nand U3900 (N_3900,N_3707,N_3064);
nor U3901 (N_3901,N_3231,N_3445);
nand U3902 (N_3902,N_3132,N_3002);
xnor U3903 (N_3903,N_3545,N_3616);
xnor U3904 (N_3904,N_3273,N_3140);
xor U3905 (N_3905,N_3649,N_3268);
or U3906 (N_3906,N_3235,N_3066);
xor U3907 (N_3907,N_3194,N_3221);
or U3908 (N_3908,N_3636,N_3478);
xor U3909 (N_3909,N_3244,N_3359);
xnor U3910 (N_3910,N_3317,N_3591);
or U3911 (N_3911,N_3101,N_3172);
xnor U3912 (N_3912,N_3690,N_3413);
xnor U3913 (N_3913,N_3658,N_3327);
nand U3914 (N_3914,N_3574,N_3024);
or U3915 (N_3915,N_3373,N_3347);
nor U3916 (N_3916,N_3328,N_3612);
or U3917 (N_3917,N_3573,N_3525);
or U3918 (N_3918,N_3051,N_3575);
nand U3919 (N_3919,N_3177,N_3582);
nor U3920 (N_3920,N_3701,N_3104);
nor U3921 (N_3921,N_3586,N_3447);
xnor U3922 (N_3922,N_3225,N_3272);
and U3923 (N_3923,N_3628,N_3202);
nand U3924 (N_3924,N_3298,N_3578);
or U3925 (N_3925,N_3457,N_3041);
xor U3926 (N_3926,N_3031,N_3254);
or U3927 (N_3927,N_3128,N_3331);
and U3928 (N_3928,N_3567,N_3725);
nand U3929 (N_3929,N_3314,N_3388);
xnor U3930 (N_3930,N_3560,N_3355);
xor U3931 (N_3931,N_3594,N_3503);
and U3932 (N_3932,N_3639,N_3651);
or U3933 (N_3933,N_3474,N_3732);
nand U3934 (N_3934,N_3598,N_3183);
nor U3935 (N_3935,N_3613,N_3704);
nand U3936 (N_3936,N_3577,N_3571);
xnor U3937 (N_3937,N_3589,N_3553);
nand U3938 (N_3938,N_3038,N_3219);
nand U3939 (N_3939,N_3223,N_3356);
xor U3940 (N_3940,N_3243,N_3094);
nor U3941 (N_3941,N_3232,N_3729);
xnor U3942 (N_3942,N_3004,N_3688);
nand U3943 (N_3943,N_3193,N_3409);
xor U3944 (N_3944,N_3029,N_3497);
or U3945 (N_3945,N_3087,N_3222);
or U3946 (N_3946,N_3423,N_3488);
xnor U3947 (N_3947,N_3098,N_3014);
nand U3948 (N_3948,N_3263,N_3546);
nand U3949 (N_3949,N_3088,N_3191);
xnor U3950 (N_3950,N_3371,N_3174);
and U3951 (N_3951,N_3722,N_3246);
and U3952 (N_3952,N_3696,N_3541);
nor U3953 (N_3953,N_3176,N_3379);
and U3954 (N_3954,N_3660,N_3640);
or U3955 (N_3955,N_3608,N_3534);
xor U3956 (N_3956,N_3097,N_3334);
xor U3957 (N_3957,N_3643,N_3078);
or U3958 (N_3958,N_3075,N_3139);
nor U3959 (N_3959,N_3215,N_3077);
and U3960 (N_3960,N_3412,N_3003);
nor U3961 (N_3961,N_3522,N_3106);
or U3962 (N_3962,N_3652,N_3294);
nand U3963 (N_3963,N_3023,N_3505);
or U3964 (N_3964,N_3495,N_3579);
nor U3965 (N_3965,N_3400,N_3515);
or U3966 (N_3966,N_3399,N_3520);
nand U3967 (N_3967,N_3321,N_3662);
and U3968 (N_3968,N_3256,N_3377);
or U3969 (N_3969,N_3127,N_3178);
nor U3970 (N_3970,N_3032,N_3166);
nand U3971 (N_3971,N_3507,N_3717);
nor U3972 (N_3972,N_3275,N_3063);
nor U3973 (N_3973,N_3604,N_3631);
or U3974 (N_3974,N_3271,N_3143);
xnor U3975 (N_3975,N_3313,N_3279);
nand U3976 (N_3976,N_3646,N_3467);
nand U3977 (N_3977,N_3282,N_3596);
xor U3978 (N_3978,N_3715,N_3407);
nand U3979 (N_3979,N_3025,N_3547);
nand U3980 (N_3980,N_3352,N_3730);
or U3981 (N_3981,N_3543,N_3252);
nor U3982 (N_3982,N_3141,N_3393);
nand U3983 (N_3983,N_3230,N_3564);
and U3984 (N_3984,N_3501,N_3216);
nor U3985 (N_3985,N_3157,N_3171);
and U3986 (N_3986,N_3008,N_3724);
nor U3987 (N_3987,N_3644,N_3201);
nor U3988 (N_3988,N_3170,N_3076);
nor U3989 (N_3989,N_3486,N_3471);
nand U3990 (N_3990,N_3372,N_3320);
and U3991 (N_3991,N_3718,N_3668);
xor U3992 (N_3992,N_3687,N_3260);
xor U3993 (N_3993,N_3676,N_3019);
nand U3994 (N_3994,N_3496,N_3309);
xor U3995 (N_3995,N_3709,N_3006);
xnor U3996 (N_3996,N_3342,N_3558);
or U3997 (N_3997,N_3259,N_3454);
nor U3998 (N_3998,N_3737,N_3401);
nor U3999 (N_3999,N_3086,N_3159);
and U4000 (N_4000,N_3061,N_3408);
nor U4001 (N_4001,N_3304,N_3052);
and U4002 (N_4002,N_3300,N_3179);
or U4003 (N_4003,N_3046,N_3703);
or U4004 (N_4004,N_3096,N_3432);
and U4005 (N_4005,N_3368,N_3630);
or U4006 (N_4006,N_3621,N_3366);
nor U4007 (N_4007,N_3385,N_3126);
nand U4008 (N_4008,N_3516,N_3236);
or U4009 (N_4009,N_3420,N_3600);
nor U4010 (N_4010,N_3679,N_3404);
nor U4011 (N_4011,N_3262,N_3070);
xnor U4012 (N_4012,N_3502,N_3370);
nand U4013 (N_4013,N_3227,N_3092);
xor U4014 (N_4014,N_3415,N_3374);
nand U4015 (N_4015,N_3710,N_3292);
or U4016 (N_4016,N_3661,N_3153);
or U4017 (N_4017,N_3197,N_3012);
or U4018 (N_4018,N_3281,N_3083);
xor U4019 (N_4019,N_3532,N_3080);
nand U4020 (N_4020,N_3035,N_3663);
nor U4021 (N_4021,N_3261,N_3017);
nor U4022 (N_4022,N_3034,N_3350);
and U4023 (N_4023,N_3054,N_3440);
nand U4024 (N_4024,N_3016,N_3568);
nand U4025 (N_4025,N_3245,N_3161);
or U4026 (N_4026,N_3135,N_3145);
nor U4027 (N_4027,N_3154,N_3258);
nand U4028 (N_4028,N_3301,N_3427);
nor U4029 (N_4029,N_3395,N_3248);
or U4030 (N_4030,N_3073,N_3308);
and U4031 (N_4031,N_3746,N_3554);
nor U4032 (N_4032,N_3697,N_3018);
or U4033 (N_4033,N_3392,N_3210);
nor U4034 (N_4034,N_3531,N_3512);
xor U4035 (N_4035,N_3537,N_3655);
nand U4036 (N_4036,N_3492,N_3615);
nor U4037 (N_4037,N_3339,N_3735);
or U4038 (N_4038,N_3524,N_3684);
nor U4039 (N_4039,N_3181,N_3102);
xnor U4040 (N_4040,N_3060,N_3511);
xnor U4041 (N_4041,N_3209,N_3099);
nor U4042 (N_4042,N_3734,N_3601);
xor U4043 (N_4043,N_3324,N_3382);
nand U4044 (N_4044,N_3265,N_3000);
and U4045 (N_4045,N_3727,N_3518);
or U4046 (N_4046,N_3473,N_3691);
xor U4047 (N_4047,N_3485,N_3716);
or U4048 (N_4048,N_3713,N_3119);
nand U4049 (N_4049,N_3026,N_3357);
and U4050 (N_4050,N_3671,N_3005);
or U4051 (N_4051,N_3529,N_3266);
or U4052 (N_4052,N_3455,N_3274);
nor U4053 (N_4053,N_3384,N_3295);
or U4054 (N_4054,N_3291,N_3521);
nor U4055 (N_4055,N_3418,N_3674);
or U4056 (N_4056,N_3115,N_3487);
nand U4057 (N_4057,N_3509,N_3555);
or U4058 (N_4058,N_3749,N_3100);
nor U4059 (N_4059,N_3464,N_3081);
nor U4060 (N_4060,N_3417,N_3443);
and U4061 (N_4061,N_3142,N_3748);
xor U4062 (N_4062,N_3133,N_3125);
nand U4063 (N_4063,N_3587,N_3278);
nand U4064 (N_4064,N_3538,N_3349);
or U4065 (N_4065,N_3444,N_3484);
xor U4066 (N_4066,N_3030,N_3584);
nor U4067 (N_4067,N_3634,N_3504);
and U4068 (N_4068,N_3346,N_3307);
or U4069 (N_4069,N_3483,N_3731);
xnor U4070 (N_4070,N_3267,N_3470);
nand U4071 (N_4071,N_3747,N_3369);
and U4072 (N_4072,N_3614,N_3240);
nor U4073 (N_4073,N_3318,N_3542);
nor U4074 (N_4074,N_3247,N_3196);
xnor U4075 (N_4075,N_3044,N_3434);
or U4076 (N_4076,N_3043,N_3344);
xnor U4077 (N_4077,N_3001,N_3323);
and U4078 (N_4078,N_3548,N_3602);
and U4079 (N_4079,N_3277,N_3158);
xor U4080 (N_4080,N_3137,N_3363);
nand U4081 (N_4081,N_3638,N_3213);
nor U4082 (N_4082,N_3533,N_3039);
nor U4083 (N_4083,N_3093,N_3431);
nand U4084 (N_4084,N_3241,N_3353);
nand U4085 (N_4085,N_3396,N_3122);
or U4086 (N_4086,N_3285,N_3228);
and U4087 (N_4087,N_3169,N_3065);
nand U4088 (N_4088,N_3390,N_3211);
and U4089 (N_4089,N_3590,N_3477);
nor U4090 (N_4090,N_3332,N_3422);
xor U4091 (N_4091,N_3669,N_3048);
xor U4092 (N_4092,N_3672,N_3394);
xor U4093 (N_4093,N_3421,N_3047);
nand U4094 (N_4094,N_3617,N_3622);
or U4095 (N_4095,N_3491,N_3472);
nand U4096 (N_4096,N_3058,N_3085);
or U4097 (N_4097,N_3335,N_3686);
nand U4098 (N_4098,N_3597,N_3337);
xnor U4099 (N_4099,N_3465,N_3315);
and U4100 (N_4100,N_3741,N_3305);
or U4101 (N_4101,N_3629,N_3288);
and U4102 (N_4102,N_3287,N_3089);
or U4103 (N_4103,N_3657,N_3059);
nor U4104 (N_4104,N_3475,N_3446);
nor U4105 (N_4105,N_3378,N_3585);
nand U4106 (N_4106,N_3117,N_3580);
nor U4107 (N_4107,N_3519,N_3458);
and U4108 (N_4108,N_3429,N_3449);
xnor U4109 (N_4109,N_3494,N_3482);
nor U4110 (N_4110,N_3441,N_3144);
nor U4111 (N_4111,N_3113,N_3705);
nor U4112 (N_4112,N_3380,N_3010);
and U4113 (N_4113,N_3131,N_3316);
nor U4114 (N_4114,N_3462,N_3110);
nand U4115 (N_4115,N_3338,N_3654);
nand U4116 (N_4116,N_3452,N_3239);
nand U4117 (N_4117,N_3149,N_3442);
or U4118 (N_4118,N_3680,N_3733);
nand U4119 (N_4119,N_3681,N_3436);
nor U4120 (N_4120,N_3045,N_3466);
xnor U4121 (N_4121,N_3508,N_3011);
xor U4122 (N_4122,N_3428,N_3609);
and U4123 (N_4123,N_3293,N_3146);
xor U4124 (N_4124,N_3062,N_3319);
xor U4125 (N_4125,N_3740,N_3702);
nor U4126 (N_4126,N_3568,N_3288);
or U4127 (N_4127,N_3465,N_3368);
or U4128 (N_4128,N_3042,N_3156);
nor U4129 (N_4129,N_3266,N_3081);
nand U4130 (N_4130,N_3304,N_3044);
or U4131 (N_4131,N_3285,N_3726);
nor U4132 (N_4132,N_3350,N_3110);
xor U4133 (N_4133,N_3552,N_3024);
xnor U4134 (N_4134,N_3216,N_3044);
nor U4135 (N_4135,N_3010,N_3016);
nand U4136 (N_4136,N_3524,N_3212);
and U4137 (N_4137,N_3050,N_3301);
and U4138 (N_4138,N_3486,N_3052);
and U4139 (N_4139,N_3025,N_3218);
and U4140 (N_4140,N_3602,N_3579);
or U4141 (N_4141,N_3225,N_3614);
or U4142 (N_4142,N_3477,N_3357);
xnor U4143 (N_4143,N_3543,N_3315);
xor U4144 (N_4144,N_3178,N_3122);
xor U4145 (N_4145,N_3524,N_3461);
xnor U4146 (N_4146,N_3722,N_3083);
nor U4147 (N_4147,N_3437,N_3177);
xnor U4148 (N_4148,N_3397,N_3169);
and U4149 (N_4149,N_3534,N_3148);
nor U4150 (N_4150,N_3436,N_3733);
xor U4151 (N_4151,N_3001,N_3288);
and U4152 (N_4152,N_3717,N_3040);
nor U4153 (N_4153,N_3590,N_3347);
xor U4154 (N_4154,N_3039,N_3558);
xor U4155 (N_4155,N_3115,N_3320);
and U4156 (N_4156,N_3291,N_3107);
or U4157 (N_4157,N_3507,N_3473);
or U4158 (N_4158,N_3224,N_3581);
xnor U4159 (N_4159,N_3014,N_3603);
or U4160 (N_4160,N_3403,N_3031);
xnor U4161 (N_4161,N_3745,N_3051);
nor U4162 (N_4162,N_3338,N_3677);
or U4163 (N_4163,N_3485,N_3612);
xor U4164 (N_4164,N_3405,N_3392);
or U4165 (N_4165,N_3196,N_3058);
nor U4166 (N_4166,N_3205,N_3515);
nand U4167 (N_4167,N_3695,N_3230);
or U4168 (N_4168,N_3069,N_3514);
or U4169 (N_4169,N_3746,N_3613);
nor U4170 (N_4170,N_3496,N_3502);
xor U4171 (N_4171,N_3592,N_3267);
and U4172 (N_4172,N_3183,N_3403);
and U4173 (N_4173,N_3736,N_3077);
or U4174 (N_4174,N_3638,N_3304);
or U4175 (N_4175,N_3424,N_3133);
nand U4176 (N_4176,N_3054,N_3411);
nor U4177 (N_4177,N_3299,N_3294);
xnor U4178 (N_4178,N_3091,N_3193);
and U4179 (N_4179,N_3211,N_3678);
nor U4180 (N_4180,N_3579,N_3076);
nand U4181 (N_4181,N_3566,N_3059);
nor U4182 (N_4182,N_3518,N_3591);
nand U4183 (N_4183,N_3152,N_3411);
nand U4184 (N_4184,N_3357,N_3674);
nand U4185 (N_4185,N_3250,N_3604);
and U4186 (N_4186,N_3384,N_3277);
nor U4187 (N_4187,N_3291,N_3424);
or U4188 (N_4188,N_3172,N_3429);
or U4189 (N_4189,N_3683,N_3045);
xor U4190 (N_4190,N_3222,N_3280);
or U4191 (N_4191,N_3693,N_3593);
xor U4192 (N_4192,N_3342,N_3094);
xor U4193 (N_4193,N_3524,N_3497);
and U4194 (N_4194,N_3052,N_3273);
nand U4195 (N_4195,N_3683,N_3462);
nor U4196 (N_4196,N_3052,N_3600);
or U4197 (N_4197,N_3377,N_3542);
xnor U4198 (N_4198,N_3384,N_3240);
nor U4199 (N_4199,N_3710,N_3655);
or U4200 (N_4200,N_3343,N_3543);
nor U4201 (N_4201,N_3142,N_3718);
or U4202 (N_4202,N_3219,N_3729);
and U4203 (N_4203,N_3672,N_3587);
nand U4204 (N_4204,N_3322,N_3675);
nand U4205 (N_4205,N_3503,N_3591);
and U4206 (N_4206,N_3707,N_3630);
nand U4207 (N_4207,N_3559,N_3661);
and U4208 (N_4208,N_3343,N_3473);
nor U4209 (N_4209,N_3326,N_3522);
or U4210 (N_4210,N_3091,N_3326);
or U4211 (N_4211,N_3293,N_3068);
or U4212 (N_4212,N_3496,N_3246);
xnor U4213 (N_4213,N_3499,N_3530);
or U4214 (N_4214,N_3061,N_3522);
or U4215 (N_4215,N_3507,N_3546);
xnor U4216 (N_4216,N_3625,N_3101);
xnor U4217 (N_4217,N_3434,N_3014);
nand U4218 (N_4218,N_3717,N_3012);
and U4219 (N_4219,N_3347,N_3073);
xnor U4220 (N_4220,N_3521,N_3585);
nand U4221 (N_4221,N_3276,N_3716);
nand U4222 (N_4222,N_3471,N_3358);
nand U4223 (N_4223,N_3275,N_3330);
nand U4224 (N_4224,N_3398,N_3179);
or U4225 (N_4225,N_3431,N_3718);
xnor U4226 (N_4226,N_3379,N_3077);
xor U4227 (N_4227,N_3380,N_3467);
nand U4228 (N_4228,N_3057,N_3504);
nor U4229 (N_4229,N_3026,N_3656);
nand U4230 (N_4230,N_3279,N_3713);
nor U4231 (N_4231,N_3267,N_3460);
or U4232 (N_4232,N_3009,N_3484);
xnor U4233 (N_4233,N_3350,N_3548);
nor U4234 (N_4234,N_3514,N_3188);
and U4235 (N_4235,N_3678,N_3656);
nor U4236 (N_4236,N_3747,N_3468);
and U4237 (N_4237,N_3184,N_3288);
nor U4238 (N_4238,N_3225,N_3130);
and U4239 (N_4239,N_3209,N_3635);
nor U4240 (N_4240,N_3675,N_3615);
nor U4241 (N_4241,N_3126,N_3059);
and U4242 (N_4242,N_3035,N_3351);
or U4243 (N_4243,N_3418,N_3648);
nor U4244 (N_4244,N_3384,N_3132);
xnor U4245 (N_4245,N_3246,N_3230);
nand U4246 (N_4246,N_3662,N_3246);
or U4247 (N_4247,N_3437,N_3353);
xor U4248 (N_4248,N_3241,N_3159);
nand U4249 (N_4249,N_3188,N_3655);
xnor U4250 (N_4250,N_3652,N_3321);
or U4251 (N_4251,N_3100,N_3514);
nand U4252 (N_4252,N_3204,N_3310);
nor U4253 (N_4253,N_3239,N_3428);
xor U4254 (N_4254,N_3697,N_3100);
or U4255 (N_4255,N_3366,N_3700);
and U4256 (N_4256,N_3573,N_3148);
nand U4257 (N_4257,N_3326,N_3314);
nor U4258 (N_4258,N_3397,N_3010);
nor U4259 (N_4259,N_3091,N_3357);
nand U4260 (N_4260,N_3135,N_3448);
and U4261 (N_4261,N_3381,N_3388);
nand U4262 (N_4262,N_3331,N_3137);
xnor U4263 (N_4263,N_3027,N_3706);
nor U4264 (N_4264,N_3212,N_3055);
nand U4265 (N_4265,N_3062,N_3265);
nor U4266 (N_4266,N_3661,N_3111);
or U4267 (N_4267,N_3531,N_3431);
or U4268 (N_4268,N_3163,N_3218);
and U4269 (N_4269,N_3447,N_3540);
nand U4270 (N_4270,N_3334,N_3401);
nor U4271 (N_4271,N_3476,N_3103);
xor U4272 (N_4272,N_3476,N_3554);
nor U4273 (N_4273,N_3677,N_3109);
and U4274 (N_4274,N_3092,N_3343);
xor U4275 (N_4275,N_3104,N_3262);
nand U4276 (N_4276,N_3101,N_3122);
nor U4277 (N_4277,N_3229,N_3485);
or U4278 (N_4278,N_3002,N_3242);
nand U4279 (N_4279,N_3595,N_3675);
nor U4280 (N_4280,N_3250,N_3523);
nand U4281 (N_4281,N_3665,N_3039);
nand U4282 (N_4282,N_3732,N_3356);
xor U4283 (N_4283,N_3128,N_3339);
or U4284 (N_4284,N_3095,N_3573);
or U4285 (N_4285,N_3646,N_3540);
or U4286 (N_4286,N_3587,N_3060);
nor U4287 (N_4287,N_3244,N_3514);
or U4288 (N_4288,N_3696,N_3671);
xnor U4289 (N_4289,N_3651,N_3749);
and U4290 (N_4290,N_3636,N_3517);
nor U4291 (N_4291,N_3605,N_3728);
nor U4292 (N_4292,N_3524,N_3334);
nor U4293 (N_4293,N_3097,N_3383);
nor U4294 (N_4294,N_3408,N_3570);
xnor U4295 (N_4295,N_3534,N_3384);
and U4296 (N_4296,N_3287,N_3054);
and U4297 (N_4297,N_3601,N_3686);
nor U4298 (N_4298,N_3699,N_3617);
and U4299 (N_4299,N_3706,N_3689);
or U4300 (N_4300,N_3622,N_3020);
xor U4301 (N_4301,N_3364,N_3656);
or U4302 (N_4302,N_3530,N_3071);
nand U4303 (N_4303,N_3062,N_3448);
nor U4304 (N_4304,N_3562,N_3589);
or U4305 (N_4305,N_3618,N_3524);
nand U4306 (N_4306,N_3306,N_3315);
nor U4307 (N_4307,N_3585,N_3457);
nand U4308 (N_4308,N_3518,N_3714);
nor U4309 (N_4309,N_3359,N_3224);
and U4310 (N_4310,N_3126,N_3642);
xor U4311 (N_4311,N_3703,N_3202);
nor U4312 (N_4312,N_3024,N_3629);
nand U4313 (N_4313,N_3633,N_3220);
or U4314 (N_4314,N_3508,N_3355);
nand U4315 (N_4315,N_3104,N_3748);
or U4316 (N_4316,N_3415,N_3346);
or U4317 (N_4317,N_3395,N_3591);
nor U4318 (N_4318,N_3267,N_3588);
xor U4319 (N_4319,N_3685,N_3567);
and U4320 (N_4320,N_3525,N_3545);
nor U4321 (N_4321,N_3276,N_3532);
xnor U4322 (N_4322,N_3690,N_3653);
nor U4323 (N_4323,N_3745,N_3010);
and U4324 (N_4324,N_3278,N_3306);
or U4325 (N_4325,N_3520,N_3724);
or U4326 (N_4326,N_3233,N_3707);
xnor U4327 (N_4327,N_3691,N_3010);
nand U4328 (N_4328,N_3125,N_3535);
xor U4329 (N_4329,N_3143,N_3077);
nand U4330 (N_4330,N_3734,N_3249);
nand U4331 (N_4331,N_3618,N_3295);
nor U4332 (N_4332,N_3579,N_3747);
and U4333 (N_4333,N_3460,N_3513);
xnor U4334 (N_4334,N_3025,N_3011);
or U4335 (N_4335,N_3684,N_3653);
and U4336 (N_4336,N_3340,N_3585);
and U4337 (N_4337,N_3277,N_3200);
or U4338 (N_4338,N_3604,N_3320);
and U4339 (N_4339,N_3096,N_3424);
xnor U4340 (N_4340,N_3249,N_3280);
nor U4341 (N_4341,N_3404,N_3011);
nand U4342 (N_4342,N_3694,N_3084);
xnor U4343 (N_4343,N_3001,N_3636);
nor U4344 (N_4344,N_3660,N_3421);
nand U4345 (N_4345,N_3401,N_3297);
or U4346 (N_4346,N_3563,N_3490);
xnor U4347 (N_4347,N_3477,N_3560);
or U4348 (N_4348,N_3381,N_3412);
nand U4349 (N_4349,N_3273,N_3325);
xor U4350 (N_4350,N_3731,N_3345);
and U4351 (N_4351,N_3556,N_3605);
nand U4352 (N_4352,N_3546,N_3254);
and U4353 (N_4353,N_3004,N_3727);
or U4354 (N_4354,N_3299,N_3551);
and U4355 (N_4355,N_3070,N_3486);
or U4356 (N_4356,N_3688,N_3048);
and U4357 (N_4357,N_3390,N_3624);
xor U4358 (N_4358,N_3724,N_3302);
xor U4359 (N_4359,N_3308,N_3403);
nand U4360 (N_4360,N_3674,N_3564);
nor U4361 (N_4361,N_3242,N_3701);
nand U4362 (N_4362,N_3344,N_3695);
or U4363 (N_4363,N_3251,N_3092);
and U4364 (N_4364,N_3325,N_3246);
xor U4365 (N_4365,N_3078,N_3109);
nand U4366 (N_4366,N_3544,N_3637);
nor U4367 (N_4367,N_3700,N_3668);
or U4368 (N_4368,N_3205,N_3018);
nor U4369 (N_4369,N_3613,N_3453);
and U4370 (N_4370,N_3174,N_3332);
or U4371 (N_4371,N_3129,N_3372);
nor U4372 (N_4372,N_3688,N_3388);
xor U4373 (N_4373,N_3328,N_3182);
nor U4374 (N_4374,N_3288,N_3084);
nand U4375 (N_4375,N_3062,N_3638);
or U4376 (N_4376,N_3071,N_3117);
xor U4377 (N_4377,N_3287,N_3154);
and U4378 (N_4378,N_3133,N_3377);
or U4379 (N_4379,N_3305,N_3037);
nor U4380 (N_4380,N_3351,N_3207);
xnor U4381 (N_4381,N_3039,N_3630);
xor U4382 (N_4382,N_3582,N_3450);
or U4383 (N_4383,N_3406,N_3461);
and U4384 (N_4384,N_3630,N_3680);
nor U4385 (N_4385,N_3653,N_3159);
and U4386 (N_4386,N_3384,N_3129);
and U4387 (N_4387,N_3334,N_3602);
xnor U4388 (N_4388,N_3145,N_3194);
or U4389 (N_4389,N_3349,N_3680);
nor U4390 (N_4390,N_3266,N_3667);
xor U4391 (N_4391,N_3263,N_3358);
and U4392 (N_4392,N_3239,N_3158);
nor U4393 (N_4393,N_3132,N_3038);
and U4394 (N_4394,N_3532,N_3180);
xnor U4395 (N_4395,N_3263,N_3146);
xor U4396 (N_4396,N_3427,N_3106);
and U4397 (N_4397,N_3177,N_3369);
and U4398 (N_4398,N_3094,N_3216);
and U4399 (N_4399,N_3102,N_3425);
nand U4400 (N_4400,N_3286,N_3312);
and U4401 (N_4401,N_3618,N_3334);
and U4402 (N_4402,N_3746,N_3581);
and U4403 (N_4403,N_3599,N_3488);
or U4404 (N_4404,N_3494,N_3689);
xor U4405 (N_4405,N_3569,N_3200);
nor U4406 (N_4406,N_3136,N_3122);
xnor U4407 (N_4407,N_3555,N_3110);
and U4408 (N_4408,N_3396,N_3067);
nor U4409 (N_4409,N_3551,N_3548);
nor U4410 (N_4410,N_3742,N_3589);
and U4411 (N_4411,N_3464,N_3225);
and U4412 (N_4412,N_3168,N_3450);
nand U4413 (N_4413,N_3121,N_3381);
nor U4414 (N_4414,N_3161,N_3521);
and U4415 (N_4415,N_3323,N_3279);
nor U4416 (N_4416,N_3532,N_3558);
nor U4417 (N_4417,N_3147,N_3532);
or U4418 (N_4418,N_3537,N_3344);
nor U4419 (N_4419,N_3231,N_3154);
xnor U4420 (N_4420,N_3516,N_3687);
nand U4421 (N_4421,N_3392,N_3458);
or U4422 (N_4422,N_3646,N_3199);
nand U4423 (N_4423,N_3033,N_3562);
xnor U4424 (N_4424,N_3731,N_3370);
nor U4425 (N_4425,N_3330,N_3655);
xor U4426 (N_4426,N_3590,N_3132);
nor U4427 (N_4427,N_3060,N_3201);
nor U4428 (N_4428,N_3219,N_3221);
and U4429 (N_4429,N_3000,N_3477);
nand U4430 (N_4430,N_3314,N_3301);
xnor U4431 (N_4431,N_3469,N_3461);
nand U4432 (N_4432,N_3339,N_3258);
and U4433 (N_4433,N_3407,N_3435);
or U4434 (N_4434,N_3438,N_3001);
and U4435 (N_4435,N_3597,N_3328);
xor U4436 (N_4436,N_3223,N_3163);
nor U4437 (N_4437,N_3136,N_3269);
or U4438 (N_4438,N_3415,N_3225);
or U4439 (N_4439,N_3077,N_3321);
nor U4440 (N_4440,N_3025,N_3174);
xor U4441 (N_4441,N_3726,N_3149);
nand U4442 (N_4442,N_3701,N_3515);
xnor U4443 (N_4443,N_3261,N_3520);
or U4444 (N_4444,N_3499,N_3656);
or U4445 (N_4445,N_3059,N_3188);
or U4446 (N_4446,N_3713,N_3475);
xnor U4447 (N_4447,N_3016,N_3011);
nand U4448 (N_4448,N_3331,N_3482);
or U4449 (N_4449,N_3058,N_3545);
nor U4450 (N_4450,N_3080,N_3403);
or U4451 (N_4451,N_3371,N_3082);
and U4452 (N_4452,N_3468,N_3084);
xnor U4453 (N_4453,N_3163,N_3092);
xnor U4454 (N_4454,N_3144,N_3022);
nor U4455 (N_4455,N_3279,N_3235);
xnor U4456 (N_4456,N_3432,N_3039);
xor U4457 (N_4457,N_3258,N_3306);
or U4458 (N_4458,N_3625,N_3292);
xnor U4459 (N_4459,N_3272,N_3148);
nor U4460 (N_4460,N_3585,N_3681);
or U4461 (N_4461,N_3569,N_3070);
or U4462 (N_4462,N_3385,N_3655);
or U4463 (N_4463,N_3124,N_3604);
nor U4464 (N_4464,N_3235,N_3172);
and U4465 (N_4465,N_3487,N_3106);
or U4466 (N_4466,N_3710,N_3484);
or U4467 (N_4467,N_3501,N_3612);
xor U4468 (N_4468,N_3353,N_3511);
nor U4469 (N_4469,N_3045,N_3140);
nor U4470 (N_4470,N_3376,N_3363);
or U4471 (N_4471,N_3614,N_3290);
nor U4472 (N_4472,N_3542,N_3378);
nor U4473 (N_4473,N_3555,N_3386);
and U4474 (N_4474,N_3264,N_3523);
nor U4475 (N_4475,N_3483,N_3354);
xor U4476 (N_4476,N_3525,N_3669);
nand U4477 (N_4477,N_3293,N_3353);
and U4478 (N_4478,N_3575,N_3272);
nor U4479 (N_4479,N_3361,N_3628);
nor U4480 (N_4480,N_3433,N_3466);
xnor U4481 (N_4481,N_3538,N_3625);
nor U4482 (N_4482,N_3542,N_3383);
nor U4483 (N_4483,N_3683,N_3100);
nor U4484 (N_4484,N_3535,N_3626);
and U4485 (N_4485,N_3659,N_3341);
and U4486 (N_4486,N_3488,N_3140);
or U4487 (N_4487,N_3428,N_3263);
or U4488 (N_4488,N_3121,N_3108);
or U4489 (N_4489,N_3227,N_3294);
and U4490 (N_4490,N_3136,N_3314);
nand U4491 (N_4491,N_3293,N_3252);
nor U4492 (N_4492,N_3398,N_3203);
or U4493 (N_4493,N_3674,N_3306);
nor U4494 (N_4494,N_3406,N_3675);
xor U4495 (N_4495,N_3453,N_3540);
or U4496 (N_4496,N_3349,N_3365);
nor U4497 (N_4497,N_3097,N_3004);
nand U4498 (N_4498,N_3518,N_3003);
nand U4499 (N_4499,N_3551,N_3080);
nor U4500 (N_4500,N_4430,N_4049);
nor U4501 (N_4501,N_4034,N_4067);
and U4502 (N_4502,N_4189,N_4433);
xor U4503 (N_4503,N_3905,N_4284);
or U4504 (N_4504,N_4353,N_4064);
nand U4505 (N_4505,N_4416,N_3880);
nor U4506 (N_4506,N_4315,N_4331);
nand U4507 (N_4507,N_4458,N_4287);
or U4508 (N_4508,N_4440,N_3857);
nor U4509 (N_4509,N_4383,N_4467);
or U4510 (N_4510,N_4148,N_4031);
or U4511 (N_4511,N_4276,N_3862);
xnor U4512 (N_4512,N_4496,N_4329);
nor U4513 (N_4513,N_4468,N_3988);
or U4514 (N_4514,N_3996,N_4402);
nand U4515 (N_4515,N_4495,N_3801);
or U4516 (N_4516,N_4098,N_3950);
or U4517 (N_4517,N_4474,N_4165);
nand U4518 (N_4518,N_4424,N_3838);
or U4519 (N_4519,N_3972,N_3964);
nor U4520 (N_4520,N_4001,N_4293);
nand U4521 (N_4521,N_4312,N_3762);
nor U4522 (N_4522,N_4217,N_4183);
and U4523 (N_4523,N_3915,N_4026);
xor U4524 (N_4524,N_4393,N_4214);
nor U4525 (N_4525,N_4074,N_4066);
nor U4526 (N_4526,N_4203,N_3881);
nand U4527 (N_4527,N_3751,N_4309);
and U4528 (N_4528,N_3969,N_4053);
nor U4529 (N_4529,N_4477,N_4472);
nand U4530 (N_4530,N_4490,N_4033);
nor U4531 (N_4531,N_3882,N_4149);
or U4532 (N_4532,N_4313,N_4350);
nand U4533 (N_4533,N_3923,N_4004);
nor U4534 (N_4534,N_4438,N_4168);
or U4535 (N_4535,N_4377,N_4073);
nand U4536 (N_4536,N_3924,N_4447);
nand U4537 (N_4537,N_3804,N_4325);
nor U4538 (N_4538,N_3831,N_4157);
nand U4539 (N_4539,N_3901,N_4288);
nand U4540 (N_4540,N_4125,N_3788);
nor U4541 (N_4541,N_4206,N_4258);
or U4542 (N_4542,N_4057,N_4326);
nand U4543 (N_4543,N_4365,N_4340);
nor U4544 (N_4544,N_3778,N_4009);
or U4545 (N_4545,N_4105,N_4109);
xor U4546 (N_4546,N_4221,N_3820);
nand U4547 (N_4547,N_4442,N_4230);
nor U4548 (N_4548,N_4235,N_4186);
xor U4549 (N_4549,N_4298,N_4341);
and U4550 (N_4550,N_4114,N_4352);
nand U4551 (N_4551,N_4172,N_3761);
nand U4552 (N_4552,N_4311,N_4076);
xnor U4553 (N_4553,N_3998,N_3891);
nand U4554 (N_4554,N_4346,N_4348);
nand U4555 (N_4555,N_4054,N_4334);
xor U4556 (N_4556,N_3949,N_3987);
nand U4557 (N_4557,N_4027,N_4407);
or U4558 (N_4558,N_3877,N_3848);
and U4559 (N_4559,N_4238,N_3911);
and U4560 (N_4560,N_4279,N_4497);
nand U4561 (N_4561,N_4386,N_3819);
nor U4562 (N_4562,N_4421,N_3758);
nor U4563 (N_4563,N_4249,N_4261);
or U4564 (N_4564,N_3780,N_4469);
or U4565 (N_4565,N_4108,N_4146);
or U4566 (N_4566,N_3883,N_4161);
or U4567 (N_4567,N_4318,N_4178);
nand U4568 (N_4568,N_4151,N_3928);
nand U4569 (N_4569,N_3767,N_4166);
or U4570 (N_4570,N_3948,N_4111);
or U4571 (N_4571,N_3990,N_4107);
xnor U4572 (N_4572,N_4250,N_4256);
and U4573 (N_4573,N_4461,N_4139);
nor U4574 (N_4574,N_4251,N_4374);
nor U4575 (N_4575,N_4022,N_4381);
nor U4576 (N_4576,N_4450,N_3887);
nor U4577 (N_4577,N_3763,N_3843);
or U4578 (N_4578,N_3782,N_3930);
nand U4579 (N_4579,N_4291,N_4234);
xor U4580 (N_4580,N_4084,N_4127);
nor U4581 (N_4581,N_4017,N_4434);
and U4582 (N_4582,N_3892,N_4006);
and U4583 (N_4583,N_4343,N_4223);
nor U4584 (N_4584,N_3976,N_3863);
nand U4585 (N_4585,N_3884,N_4356);
and U4586 (N_4586,N_4129,N_4038);
nor U4587 (N_4587,N_4457,N_3844);
xor U4588 (N_4588,N_3773,N_4220);
xnor U4589 (N_4589,N_4039,N_3897);
or U4590 (N_4590,N_3939,N_4498);
and U4591 (N_4591,N_4056,N_4379);
nor U4592 (N_4592,N_4021,N_3834);
nor U4593 (N_4593,N_4182,N_4015);
nor U4594 (N_4594,N_3845,N_3798);
and U4595 (N_4595,N_4385,N_4248);
nor U4596 (N_4596,N_4337,N_3833);
and U4597 (N_4597,N_4414,N_4306);
and U4598 (N_4598,N_4427,N_3753);
or U4599 (N_4599,N_3854,N_3941);
nor U4600 (N_4600,N_4032,N_4283);
nor U4601 (N_4601,N_4308,N_3997);
nor U4602 (N_4602,N_4491,N_4000);
nand U4603 (N_4603,N_3992,N_4211);
nor U4604 (N_4604,N_4304,N_4411);
xnor U4605 (N_4605,N_4141,N_4364);
nor U4606 (N_4606,N_4366,N_4226);
nor U4607 (N_4607,N_4269,N_3955);
or U4608 (N_4608,N_4199,N_4347);
nor U4609 (N_4609,N_3828,N_4289);
xor U4610 (N_4610,N_4042,N_3817);
or U4611 (N_4611,N_4236,N_3959);
or U4612 (N_4612,N_4167,N_3971);
nand U4613 (N_4613,N_4476,N_4462);
xor U4614 (N_4614,N_4130,N_4398);
or U4615 (N_4615,N_4263,N_3846);
nand U4616 (N_4616,N_4224,N_4436);
and U4617 (N_4617,N_3864,N_3812);
nor U4618 (N_4618,N_4390,N_4209);
or U4619 (N_4619,N_4323,N_4344);
nor U4620 (N_4620,N_4321,N_4371);
xor U4621 (N_4621,N_3945,N_4210);
nand U4622 (N_4622,N_4378,N_3919);
nor U4623 (N_4623,N_4155,N_3821);
and U4624 (N_4624,N_4181,N_4142);
xnor U4625 (N_4625,N_4216,N_4271);
or U4626 (N_4626,N_4092,N_3755);
nor U4627 (N_4627,N_3847,N_3985);
nand U4628 (N_4628,N_4445,N_4062);
and U4629 (N_4629,N_3837,N_3965);
nand U4630 (N_4630,N_4011,N_4116);
or U4631 (N_4631,N_4426,N_4302);
and U4632 (N_4632,N_4046,N_4449);
xnor U4633 (N_4633,N_4078,N_3994);
xor U4634 (N_4634,N_3807,N_4484);
nand U4635 (N_4635,N_4425,N_4035);
or U4636 (N_4636,N_4012,N_3760);
nand U4637 (N_4637,N_4025,N_4136);
xnor U4638 (N_4638,N_3876,N_4100);
nor U4639 (N_4639,N_4405,N_4095);
nand U4640 (N_4640,N_4252,N_4133);
or U4641 (N_4641,N_4071,N_4154);
and U4642 (N_4642,N_3787,N_4264);
nor U4643 (N_4643,N_4205,N_3800);
and U4644 (N_4644,N_4389,N_4265);
xor U4645 (N_4645,N_4094,N_3826);
and U4646 (N_4646,N_4396,N_4110);
nand U4647 (N_4647,N_4330,N_4124);
xor U4648 (N_4648,N_4406,N_3858);
nor U4649 (N_4649,N_3774,N_4020);
xor U4650 (N_4650,N_4227,N_3866);
and U4651 (N_4651,N_4455,N_4336);
or U4652 (N_4652,N_4065,N_3810);
nand U4653 (N_4653,N_4409,N_4314);
nor U4654 (N_4654,N_3789,N_3870);
nand U4655 (N_4655,N_4176,N_4218);
nand U4656 (N_4656,N_3806,N_3783);
or U4657 (N_4657,N_3960,N_3829);
or U4658 (N_4658,N_3979,N_4204);
or U4659 (N_4659,N_3865,N_3791);
nand U4660 (N_4660,N_3898,N_4091);
nand U4661 (N_4661,N_4104,N_3794);
and U4662 (N_4662,N_4088,N_4096);
and U4663 (N_4663,N_3759,N_4454);
or U4664 (N_4664,N_4499,N_3793);
nand U4665 (N_4665,N_4040,N_3776);
and U4666 (N_4666,N_4122,N_3902);
nor U4667 (N_4667,N_4101,N_4202);
or U4668 (N_4668,N_4037,N_4192);
nand U4669 (N_4669,N_4069,N_3951);
or U4670 (N_4670,N_4175,N_4429);
or U4671 (N_4671,N_3920,N_3896);
or U4672 (N_4672,N_3961,N_4355);
or U4673 (N_4673,N_4362,N_3932);
or U4674 (N_4674,N_4145,N_4401);
xnor U4675 (N_4675,N_4131,N_3940);
nor U4676 (N_4676,N_3904,N_4241);
nor U4677 (N_4677,N_4085,N_4392);
nor U4678 (N_4678,N_4010,N_4063);
nand U4679 (N_4679,N_4187,N_4090);
or U4680 (N_4680,N_4296,N_3859);
or U4681 (N_4681,N_4008,N_3918);
nor U4682 (N_4682,N_4123,N_4068);
and U4683 (N_4683,N_4059,N_4135);
xnor U4684 (N_4684,N_3910,N_4003);
and U4685 (N_4685,N_4316,N_4338);
nand U4686 (N_4686,N_4297,N_4232);
nand U4687 (N_4687,N_4201,N_3768);
and U4688 (N_4688,N_4043,N_3893);
or U4689 (N_4689,N_4270,N_3764);
nor U4690 (N_4690,N_3995,N_3832);
nor U4691 (N_4691,N_4388,N_4475);
and U4692 (N_4692,N_3840,N_4075);
or U4693 (N_4693,N_3873,N_4333);
nand U4694 (N_4694,N_4119,N_4262);
and U4695 (N_4695,N_3936,N_3909);
or U4696 (N_4696,N_4048,N_3977);
or U4697 (N_4697,N_4115,N_4013);
or U4698 (N_4698,N_3824,N_4327);
nand U4699 (N_4699,N_4273,N_4354);
nor U4700 (N_4700,N_3903,N_4277);
nor U4701 (N_4701,N_4050,N_4415);
nor U4702 (N_4702,N_3795,N_4492);
xor U4703 (N_4703,N_4198,N_4132);
xnor U4704 (N_4704,N_3850,N_4358);
xnor U4705 (N_4705,N_4185,N_3856);
nand U4706 (N_4706,N_3906,N_3975);
xor U4707 (N_4707,N_3852,N_4267);
nor U4708 (N_4708,N_4222,N_3802);
nand U4709 (N_4709,N_4300,N_3953);
and U4710 (N_4710,N_4134,N_4180);
or U4711 (N_4711,N_3855,N_3929);
xnor U4712 (N_4712,N_4349,N_4400);
and U4713 (N_4713,N_4128,N_4086);
nand U4714 (N_4714,N_4439,N_3869);
nor U4715 (N_4715,N_3899,N_3885);
nand U4716 (N_4716,N_3931,N_3769);
or U4717 (N_4717,N_3750,N_3808);
nor U4718 (N_4718,N_4423,N_4137);
xor U4719 (N_4719,N_4479,N_3942);
nand U4720 (N_4720,N_3890,N_4058);
xor U4721 (N_4721,N_3839,N_4410);
or U4722 (N_4722,N_4370,N_4272);
or U4723 (N_4723,N_3927,N_4305);
or U4724 (N_4724,N_4482,N_3818);
nand U4725 (N_4725,N_4106,N_3967);
nand U4726 (N_4726,N_4233,N_4412);
xnor U4727 (N_4727,N_3874,N_4029);
and U4728 (N_4728,N_3842,N_4244);
or U4729 (N_4729,N_4219,N_4229);
and U4730 (N_4730,N_4237,N_3779);
xor U4731 (N_4731,N_4169,N_3963);
xnor U4732 (N_4732,N_3888,N_4159);
and U4733 (N_4733,N_4282,N_4324);
or U4734 (N_4734,N_3922,N_4303);
nor U4735 (N_4735,N_4367,N_3803);
or U4736 (N_4736,N_3886,N_4170);
xnor U4737 (N_4737,N_3926,N_3786);
xor U4738 (N_4738,N_4481,N_4120);
xnor U4739 (N_4739,N_4144,N_4443);
nor U4740 (N_4740,N_3777,N_4399);
xnor U4741 (N_4741,N_4420,N_4463);
xor U4742 (N_4742,N_4488,N_4342);
or U4743 (N_4743,N_4072,N_4275);
xnor U4744 (N_4744,N_4382,N_4268);
and U4745 (N_4745,N_4018,N_4422);
nand U4746 (N_4746,N_3784,N_4404);
or U4747 (N_4747,N_4152,N_4190);
nand U4748 (N_4748,N_4239,N_4322);
or U4749 (N_4749,N_4471,N_4257);
or U4750 (N_4750,N_3815,N_4156);
xnor U4751 (N_4751,N_4451,N_3813);
and U4752 (N_4752,N_4281,N_3772);
xnor U4753 (N_4753,N_4278,N_4081);
nor U4754 (N_4754,N_3861,N_4369);
or U4755 (N_4755,N_4162,N_4207);
xor U4756 (N_4756,N_4197,N_4339);
xnor U4757 (N_4757,N_4184,N_4486);
and U4758 (N_4758,N_4179,N_3796);
and U4759 (N_4759,N_4014,N_4002);
nand U4760 (N_4760,N_4375,N_4243);
or U4761 (N_4761,N_3809,N_4225);
or U4762 (N_4762,N_3993,N_3836);
nor U4763 (N_4763,N_4351,N_4024);
nor U4764 (N_4764,N_4387,N_4143);
and U4765 (N_4765,N_4394,N_3871);
or U4766 (N_4766,N_4016,N_3894);
or U4767 (N_4767,N_4335,N_4260);
nor U4768 (N_4768,N_4373,N_4254);
xnor U4769 (N_4769,N_3830,N_4290);
or U4770 (N_4770,N_4193,N_3968);
and U4771 (N_4771,N_4286,N_4310);
nand U4772 (N_4772,N_4147,N_3766);
nand U4773 (N_4773,N_4483,N_4140);
xor U4774 (N_4774,N_4307,N_3925);
or U4775 (N_4775,N_4470,N_4087);
xnor U4776 (N_4776,N_4395,N_4099);
nand U4777 (N_4777,N_4453,N_3878);
or U4778 (N_4778,N_3935,N_4007);
and U4779 (N_4779,N_4478,N_4295);
xnor U4780 (N_4780,N_3756,N_3805);
nor U4781 (N_4781,N_4195,N_4174);
and U4782 (N_4782,N_4391,N_4177);
nor U4783 (N_4783,N_3966,N_4208);
nor U4784 (N_4784,N_4055,N_3981);
xnor U4785 (N_4785,N_4245,N_4444);
and U4786 (N_4786,N_4158,N_4052);
and U4787 (N_4787,N_3860,N_4357);
and U4788 (N_4788,N_3872,N_4036);
or U4789 (N_4789,N_4372,N_4464);
xnor U4790 (N_4790,N_4044,N_4419);
nor U4791 (N_4791,N_4060,N_3868);
or U4792 (N_4792,N_4240,N_4089);
nor U4793 (N_4793,N_3814,N_3849);
xor U4794 (N_4794,N_4319,N_3991);
xor U4795 (N_4795,N_3785,N_4465);
nand U4796 (N_4796,N_4045,N_4380);
nor U4797 (N_4797,N_3917,N_3816);
nand U4798 (N_4798,N_4097,N_4079);
and U4799 (N_4799,N_4196,N_4126);
or U4800 (N_4800,N_4118,N_4191);
nor U4801 (N_4801,N_4408,N_4160);
nor U4802 (N_4802,N_3914,N_4317);
xnor U4803 (N_4803,N_4431,N_4494);
or U4804 (N_4804,N_3853,N_3811);
or U4805 (N_4805,N_4292,N_4173);
nand U4806 (N_4806,N_3956,N_4121);
xor U4807 (N_4807,N_4274,N_4441);
and U4808 (N_4808,N_4452,N_4361);
nand U4809 (N_4809,N_3933,N_4345);
xnor U4810 (N_4810,N_3989,N_4320);
xor U4811 (N_4811,N_4456,N_3916);
or U4812 (N_4812,N_3775,N_4487);
nand U4813 (N_4813,N_4359,N_3970);
or U4814 (N_4814,N_3825,N_4299);
and U4815 (N_4815,N_3912,N_3974);
xor U4816 (N_4816,N_4432,N_4077);
and U4817 (N_4817,N_3752,N_3841);
nand U4818 (N_4818,N_4150,N_4047);
nand U4819 (N_4819,N_4363,N_4360);
nor U4820 (N_4820,N_4448,N_4188);
xnor U4821 (N_4821,N_4212,N_3757);
xor U4822 (N_4822,N_4376,N_4294);
and U4823 (N_4823,N_4466,N_3900);
and U4824 (N_4824,N_4051,N_3962);
xnor U4825 (N_4825,N_3822,N_4083);
and U4826 (N_4826,N_4397,N_3952);
or U4827 (N_4827,N_4242,N_3827);
nor U4828 (N_4828,N_4493,N_4213);
and U4829 (N_4829,N_4164,N_3867);
or U4830 (N_4830,N_4019,N_3984);
xnor U4831 (N_4831,N_3851,N_4112);
xnor U4832 (N_4832,N_4061,N_3879);
or U4833 (N_4833,N_4023,N_4460);
nor U4834 (N_4834,N_4417,N_3986);
nor U4835 (N_4835,N_4080,N_4041);
nand U4836 (N_4836,N_3973,N_3908);
xor U4837 (N_4837,N_4247,N_3770);
and U4838 (N_4838,N_3797,N_4103);
or U4839 (N_4839,N_4485,N_3790);
and U4840 (N_4840,N_4093,N_3875);
nor U4841 (N_4841,N_4117,N_4030);
and U4842 (N_4842,N_4194,N_3958);
nor U4843 (N_4843,N_4200,N_3921);
nor U4844 (N_4844,N_4070,N_4437);
and U4845 (N_4845,N_3980,N_3982);
and U4846 (N_4846,N_3954,N_3907);
and U4847 (N_4847,N_3937,N_4231);
nor U4848 (N_4848,N_4259,N_4418);
xnor U4849 (N_4849,N_4028,N_3938);
nor U4850 (N_4850,N_4413,N_3913);
nand U4851 (N_4851,N_4082,N_4332);
nor U4852 (N_4852,N_3792,N_4280);
nand U4853 (N_4853,N_4138,N_3934);
nand U4854 (N_4854,N_4228,N_3754);
xor U4855 (N_4855,N_4253,N_4246);
nand U4856 (N_4856,N_4301,N_4171);
and U4857 (N_4857,N_4459,N_3781);
or U4858 (N_4858,N_3946,N_4005);
or U4859 (N_4859,N_4285,N_4368);
xnor U4860 (N_4860,N_3944,N_4266);
xor U4861 (N_4861,N_4328,N_3835);
nor U4862 (N_4862,N_4102,N_4163);
and U4863 (N_4863,N_4215,N_4384);
xnor U4864 (N_4864,N_4489,N_3978);
xnor U4865 (N_4865,N_4255,N_3895);
nand U4866 (N_4866,N_4446,N_3983);
nor U4867 (N_4867,N_3799,N_4473);
xnor U4868 (N_4868,N_4403,N_3957);
nor U4869 (N_4869,N_3771,N_3947);
and U4870 (N_4870,N_4428,N_3823);
nand U4871 (N_4871,N_3943,N_4113);
nor U4872 (N_4872,N_3889,N_3765);
and U4873 (N_4873,N_4480,N_4435);
xor U4874 (N_4874,N_4153,N_3999);
nor U4875 (N_4875,N_4022,N_4049);
xnor U4876 (N_4876,N_3986,N_4457);
or U4877 (N_4877,N_4249,N_4279);
nand U4878 (N_4878,N_3858,N_3987);
xor U4879 (N_4879,N_3855,N_4467);
nor U4880 (N_4880,N_4015,N_4006);
nand U4881 (N_4881,N_3890,N_3897);
nor U4882 (N_4882,N_4256,N_4355);
nor U4883 (N_4883,N_3974,N_4171);
or U4884 (N_4884,N_4211,N_3905);
xnor U4885 (N_4885,N_4148,N_3760);
xor U4886 (N_4886,N_3849,N_3815);
or U4887 (N_4887,N_4267,N_3857);
or U4888 (N_4888,N_4441,N_4128);
xnor U4889 (N_4889,N_4049,N_4272);
xor U4890 (N_4890,N_4101,N_4337);
xor U4891 (N_4891,N_3951,N_4185);
nor U4892 (N_4892,N_3971,N_4374);
xor U4893 (N_4893,N_4127,N_4097);
nand U4894 (N_4894,N_3991,N_4119);
or U4895 (N_4895,N_4326,N_4141);
xnor U4896 (N_4896,N_3766,N_4478);
and U4897 (N_4897,N_3980,N_4431);
and U4898 (N_4898,N_3988,N_4352);
xor U4899 (N_4899,N_3910,N_3862);
xor U4900 (N_4900,N_4408,N_3810);
nand U4901 (N_4901,N_4470,N_3845);
nand U4902 (N_4902,N_4453,N_4358);
xnor U4903 (N_4903,N_3948,N_3944);
xor U4904 (N_4904,N_4496,N_4219);
nor U4905 (N_4905,N_4058,N_4457);
xor U4906 (N_4906,N_4410,N_4487);
and U4907 (N_4907,N_3794,N_3821);
nand U4908 (N_4908,N_4063,N_4174);
or U4909 (N_4909,N_3881,N_4345);
xor U4910 (N_4910,N_4491,N_4070);
or U4911 (N_4911,N_3983,N_3932);
and U4912 (N_4912,N_4245,N_4250);
nor U4913 (N_4913,N_4026,N_4284);
or U4914 (N_4914,N_4465,N_4338);
nand U4915 (N_4915,N_4191,N_3950);
nand U4916 (N_4916,N_4489,N_4205);
or U4917 (N_4917,N_4275,N_3862);
or U4918 (N_4918,N_4016,N_4248);
nand U4919 (N_4919,N_4349,N_4286);
nor U4920 (N_4920,N_4342,N_4184);
nand U4921 (N_4921,N_3803,N_4081);
nor U4922 (N_4922,N_4273,N_4488);
nor U4923 (N_4923,N_4037,N_4176);
xnor U4924 (N_4924,N_4486,N_4134);
or U4925 (N_4925,N_4272,N_3831);
xor U4926 (N_4926,N_4375,N_4202);
or U4927 (N_4927,N_3975,N_4406);
nor U4928 (N_4928,N_4191,N_4474);
xnor U4929 (N_4929,N_3839,N_4441);
and U4930 (N_4930,N_4090,N_3852);
xnor U4931 (N_4931,N_3754,N_4380);
nor U4932 (N_4932,N_3875,N_4484);
xor U4933 (N_4933,N_4326,N_3971);
and U4934 (N_4934,N_4395,N_4344);
and U4935 (N_4935,N_4226,N_4124);
and U4936 (N_4936,N_4217,N_4052);
xnor U4937 (N_4937,N_4450,N_4153);
nor U4938 (N_4938,N_4474,N_3774);
nor U4939 (N_4939,N_3877,N_3846);
or U4940 (N_4940,N_4199,N_4059);
nand U4941 (N_4941,N_4264,N_3797);
nor U4942 (N_4942,N_4072,N_4193);
nand U4943 (N_4943,N_3793,N_4231);
nand U4944 (N_4944,N_4084,N_4110);
or U4945 (N_4945,N_3762,N_4362);
nor U4946 (N_4946,N_3949,N_4279);
and U4947 (N_4947,N_4276,N_3760);
nand U4948 (N_4948,N_3916,N_4366);
and U4949 (N_4949,N_4062,N_3966);
and U4950 (N_4950,N_3807,N_4070);
and U4951 (N_4951,N_4498,N_4349);
xnor U4952 (N_4952,N_4275,N_3827);
and U4953 (N_4953,N_4145,N_4200);
nand U4954 (N_4954,N_4037,N_4286);
or U4955 (N_4955,N_4490,N_4351);
or U4956 (N_4956,N_4335,N_4445);
nand U4957 (N_4957,N_3869,N_4325);
xnor U4958 (N_4958,N_4163,N_4189);
nand U4959 (N_4959,N_3834,N_4449);
nor U4960 (N_4960,N_3987,N_4381);
xor U4961 (N_4961,N_4407,N_4498);
or U4962 (N_4962,N_4050,N_4402);
or U4963 (N_4963,N_3885,N_3769);
or U4964 (N_4964,N_4111,N_3985);
nand U4965 (N_4965,N_3942,N_4451);
xnor U4966 (N_4966,N_4313,N_3888);
or U4967 (N_4967,N_3788,N_4387);
and U4968 (N_4968,N_4101,N_3794);
nor U4969 (N_4969,N_3974,N_4118);
nand U4970 (N_4970,N_4135,N_4309);
nand U4971 (N_4971,N_4401,N_4362);
nor U4972 (N_4972,N_4182,N_4009);
and U4973 (N_4973,N_3758,N_4304);
or U4974 (N_4974,N_4473,N_4341);
and U4975 (N_4975,N_4316,N_4378);
xnor U4976 (N_4976,N_4406,N_4417);
and U4977 (N_4977,N_4210,N_4413);
xor U4978 (N_4978,N_4279,N_3803);
xnor U4979 (N_4979,N_4348,N_3757);
and U4980 (N_4980,N_4368,N_4033);
nand U4981 (N_4981,N_4337,N_4332);
nand U4982 (N_4982,N_4423,N_4313);
and U4983 (N_4983,N_3936,N_4289);
and U4984 (N_4984,N_3848,N_3934);
nand U4985 (N_4985,N_3977,N_4372);
xnor U4986 (N_4986,N_3805,N_4231);
or U4987 (N_4987,N_3846,N_4301);
xor U4988 (N_4988,N_3817,N_3997);
xor U4989 (N_4989,N_4371,N_4415);
xor U4990 (N_4990,N_3924,N_4270);
nand U4991 (N_4991,N_4245,N_4120);
and U4992 (N_4992,N_4483,N_4101);
xor U4993 (N_4993,N_4313,N_4065);
nor U4994 (N_4994,N_3947,N_4256);
nor U4995 (N_4995,N_3883,N_4234);
nor U4996 (N_4996,N_4239,N_3937);
xor U4997 (N_4997,N_4273,N_3770);
nand U4998 (N_4998,N_3780,N_4338);
nor U4999 (N_4999,N_4485,N_4272);
and U5000 (N_5000,N_4097,N_3752);
and U5001 (N_5001,N_4106,N_4326);
nor U5002 (N_5002,N_4421,N_3913);
or U5003 (N_5003,N_4388,N_4447);
xnor U5004 (N_5004,N_4187,N_4291);
nand U5005 (N_5005,N_3931,N_4005);
xnor U5006 (N_5006,N_3792,N_3807);
xor U5007 (N_5007,N_3881,N_4412);
and U5008 (N_5008,N_4170,N_4320);
and U5009 (N_5009,N_3864,N_4338);
nand U5010 (N_5010,N_4187,N_3989);
nor U5011 (N_5011,N_4335,N_4447);
xnor U5012 (N_5012,N_3782,N_3898);
or U5013 (N_5013,N_3873,N_4216);
nor U5014 (N_5014,N_4037,N_4214);
or U5015 (N_5015,N_3786,N_3812);
xor U5016 (N_5016,N_3914,N_3926);
nand U5017 (N_5017,N_4022,N_4058);
nor U5018 (N_5018,N_3835,N_4285);
nor U5019 (N_5019,N_3809,N_4482);
xnor U5020 (N_5020,N_3784,N_4497);
and U5021 (N_5021,N_4063,N_4460);
or U5022 (N_5022,N_4395,N_4168);
nand U5023 (N_5023,N_3977,N_4335);
xor U5024 (N_5024,N_4258,N_4490);
and U5025 (N_5025,N_4277,N_4259);
and U5026 (N_5026,N_3881,N_3896);
nor U5027 (N_5027,N_3965,N_4300);
nand U5028 (N_5028,N_4270,N_3856);
nor U5029 (N_5029,N_3800,N_4233);
and U5030 (N_5030,N_4465,N_4479);
nor U5031 (N_5031,N_3916,N_4063);
nor U5032 (N_5032,N_3983,N_3828);
nor U5033 (N_5033,N_4160,N_4100);
or U5034 (N_5034,N_4258,N_4096);
xor U5035 (N_5035,N_4217,N_3920);
nand U5036 (N_5036,N_4113,N_4335);
xor U5037 (N_5037,N_4246,N_4426);
nand U5038 (N_5038,N_3769,N_4455);
nor U5039 (N_5039,N_4488,N_4306);
or U5040 (N_5040,N_3766,N_4052);
nand U5041 (N_5041,N_3799,N_3996);
xor U5042 (N_5042,N_4298,N_3904);
and U5043 (N_5043,N_4495,N_4197);
xnor U5044 (N_5044,N_4288,N_4052);
xor U5045 (N_5045,N_4267,N_4395);
or U5046 (N_5046,N_3836,N_4084);
nand U5047 (N_5047,N_3935,N_3864);
xor U5048 (N_5048,N_4470,N_4372);
nand U5049 (N_5049,N_3755,N_3989);
nand U5050 (N_5050,N_4015,N_4232);
and U5051 (N_5051,N_4026,N_4438);
xnor U5052 (N_5052,N_4246,N_4140);
nand U5053 (N_5053,N_3838,N_4436);
and U5054 (N_5054,N_3810,N_3945);
or U5055 (N_5055,N_3937,N_4335);
or U5056 (N_5056,N_4320,N_4104);
nand U5057 (N_5057,N_4396,N_4219);
or U5058 (N_5058,N_3868,N_3862);
nor U5059 (N_5059,N_4149,N_4249);
and U5060 (N_5060,N_4383,N_4412);
or U5061 (N_5061,N_4323,N_4049);
nand U5062 (N_5062,N_4445,N_4115);
or U5063 (N_5063,N_4254,N_3771);
xor U5064 (N_5064,N_3918,N_3751);
and U5065 (N_5065,N_4460,N_4310);
nor U5066 (N_5066,N_3751,N_4068);
xnor U5067 (N_5067,N_4197,N_4026);
xor U5068 (N_5068,N_3998,N_4009);
and U5069 (N_5069,N_4132,N_4121);
or U5070 (N_5070,N_3786,N_4161);
xnor U5071 (N_5071,N_4214,N_4177);
nand U5072 (N_5072,N_4340,N_3840);
or U5073 (N_5073,N_3833,N_3978);
nor U5074 (N_5074,N_4130,N_4122);
nand U5075 (N_5075,N_4149,N_4457);
nand U5076 (N_5076,N_4463,N_4154);
and U5077 (N_5077,N_4005,N_4393);
nand U5078 (N_5078,N_3936,N_4136);
xor U5079 (N_5079,N_3918,N_4437);
and U5080 (N_5080,N_4196,N_3871);
xnor U5081 (N_5081,N_4331,N_4373);
or U5082 (N_5082,N_4265,N_3992);
xnor U5083 (N_5083,N_3828,N_4431);
nand U5084 (N_5084,N_4439,N_4098);
nor U5085 (N_5085,N_3810,N_4355);
and U5086 (N_5086,N_4057,N_3825);
or U5087 (N_5087,N_4095,N_4215);
and U5088 (N_5088,N_3878,N_3959);
nor U5089 (N_5089,N_4078,N_3908);
or U5090 (N_5090,N_4218,N_4220);
or U5091 (N_5091,N_4278,N_4040);
nor U5092 (N_5092,N_4132,N_4197);
or U5093 (N_5093,N_4428,N_4152);
xnor U5094 (N_5094,N_3910,N_4450);
and U5095 (N_5095,N_3942,N_3826);
xor U5096 (N_5096,N_3959,N_4040);
nand U5097 (N_5097,N_4060,N_3812);
nand U5098 (N_5098,N_4423,N_4328);
xor U5099 (N_5099,N_3858,N_3760);
and U5100 (N_5100,N_4271,N_3924);
xor U5101 (N_5101,N_4499,N_4383);
xor U5102 (N_5102,N_3804,N_3889);
nor U5103 (N_5103,N_4370,N_3811);
nor U5104 (N_5104,N_4458,N_4472);
and U5105 (N_5105,N_4358,N_4307);
nor U5106 (N_5106,N_4145,N_4284);
nor U5107 (N_5107,N_4421,N_4444);
nor U5108 (N_5108,N_4256,N_4217);
and U5109 (N_5109,N_4066,N_4023);
or U5110 (N_5110,N_4051,N_4256);
nand U5111 (N_5111,N_4091,N_4033);
nor U5112 (N_5112,N_3771,N_4441);
nand U5113 (N_5113,N_4044,N_3780);
and U5114 (N_5114,N_4121,N_4464);
or U5115 (N_5115,N_3934,N_3854);
nor U5116 (N_5116,N_3779,N_4230);
or U5117 (N_5117,N_3795,N_4229);
xnor U5118 (N_5118,N_4353,N_3974);
xnor U5119 (N_5119,N_4176,N_4366);
xnor U5120 (N_5120,N_4215,N_4254);
and U5121 (N_5121,N_4000,N_4321);
or U5122 (N_5122,N_4377,N_3957);
and U5123 (N_5123,N_4187,N_3949);
and U5124 (N_5124,N_3755,N_3962);
nand U5125 (N_5125,N_3831,N_4161);
nor U5126 (N_5126,N_4357,N_3960);
or U5127 (N_5127,N_3793,N_4298);
and U5128 (N_5128,N_4383,N_4361);
xnor U5129 (N_5129,N_3843,N_3974);
xnor U5130 (N_5130,N_3871,N_4386);
or U5131 (N_5131,N_4312,N_4352);
nand U5132 (N_5132,N_4350,N_4046);
nand U5133 (N_5133,N_4372,N_4277);
or U5134 (N_5134,N_4107,N_4329);
nor U5135 (N_5135,N_3856,N_4032);
xor U5136 (N_5136,N_4093,N_4472);
nand U5137 (N_5137,N_4053,N_4469);
and U5138 (N_5138,N_4403,N_4352);
or U5139 (N_5139,N_4112,N_4000);
nor U5140 (N_5140,N_4048,N_4377);
and U5141 (N_5141,N_4351,N_3851);
or U5142 (N_5142,N_4380,N_4155);
nand U5143 (N_5143,N_4393,N_4003);
nand U5144 (N_5144,N_4015,N_4390);
xor U5145 (N_5145,N_4422,N_4150);
or U5146 (N_5146,N_4465,N_3761);
xnor U5147 (N_5147,N_4110,N_4059);
xor U5148 (N_5148,N_4441,N_4345);
nand U5149 (N_5149,N_4117,N_4116);
or U5150 (N_5150,N_4163,N_3788);
and U5151 (N_5151,N_4336,N_4089);
or U5152 (N_5152,N_4082,N_3888);
or U5153 (N_5153,N_4295,N_3912);
nor U5154 (N_5154,N_4326,N_3869);
nor U5155 (N_5155,N_4323,N_4317);
or U5156 (N_5156,N_3805,N_4014);
and U5157 (N_5157,N_4344,N_4441);
and U5158 (N_5158,N_4464,N_3880);
or U5159 (N_5159,N_3822,N_4243);
and U5160 (N_5160,N_4327,N_4347);
xnor U5161 (N_5161,N_4297,N_3884);
nor U5162 (N_5162,N_4187,N_3947);
nand U5163 (N_5163,N_3805,N_4184);
nand U5164 (N_5164,N_4297,N_4256);
xor U5165 (N_5165,N_3806,N_4109);
or U5166 (N_5166,N_4404,N_4036);
nor U5167 (N_5167,N_3885,N_3900);
nor U5168 (N_5168,N_4047,N_4423);
or U5169 (N_5169,N_3820,N_4472);
nand U5170 (N_5170,N_4153,N_4454);
xor U5171 (N_5171,N_3854,N_4237);
xor U5172 (N_5172,N_3887,N_3964);
and U5173 (N_5173,N_3806,N_4309);
xnor U5174 (N_5174,N_4412,N_3901);
xor U5175 (N_5175,N_3996,N_4367);
or U5176 (N_5176,N_3901,N_4104);
or U5177 (N_5177,N_3835,N_3859);
and U5178 (N_5178,N_4089,N_3763);
nor U5179 (N_5179,N_3983,N_4152);
nor U5180 (N_5180,N_4226,N_4193);
nand U5181 (N_5181,N_3904,N_3804);
nand U5182 (N_5182,N_4004,N_4401);
or U5183 (N_5183,N_3873,N_4455);
xnor U5184 (N_5184,N_4137,N_4038);
or U5185 (N_5185,N_3753,N_4433);
nand U5186 (N_5186,N_3918,N_4055);
nand U5187 (N_5187,N_4255,N_3766);
nor U5188 (N_5188,N_3758,N_4277);
xnor U5189 (N_5189,N_3836,N_4347);
nand U5190 (N_5190,N_3842,N_4307);
and U5191 (N_5191,N_4054,N_4322);
or U5192 (N_5192,N_4457,N_4276);
or U5193 (N_5193,N_4286,N_3901);
nand U5194 (N_5194,N_3777,N_4042);
and U5195 (N_5195,N_3892,N_4466);
and U5196 (N_5196,N_3800,N_3883);
or U5197 (N_5197,N_4169,N_4251);
nand U5198 (N_5198,N_4357,N_4156);
nand U5199 (N_5199,N_3905,N_3951);
or U5200 (N_5200,N_3880,N_4233);
and U5201 (N_5201,N_4105,N_3789);
nor U5202 (N_5202,N_3986,N_4002);
nand U5203 (N_5203,N_3905,N_4157);
and U5204 (N_5204,N_4032,N_3774);
nand U5205 (N_5205,N_3871,N_4165);
nand U5206 (N_5206,N_4380,N_4023);
nand U5207 (N_5207,N_4088,N_4074);
xor U5208 (N_5208,N_3934,N_3793);
or U5209 (N_5209,N_4473,N_4201);
xnor U5210 (N_5210,N_4383,N_4199);
nor U5211 (N_5211,N_4105,N_4417);
or U5212 (N_5212,N_4463,N_4321);
or U5213 (N_5213,N_4029,N_3785);
nand U5214 (N_5214,N_4221,N_4177);
and U5215 (N_5215,N_3817,N_4001);
and U5216 (N_5216,N_4132,N_3838);
or U5217 (N_5217,N_4332,N_4011);
or U5218 (N_5218,N_4203,N_4371);
and U5219 (N_5219,N_4413,N_3823);
xor U5220 (N_5220,N_3866,N_4156);
nand U5221 (N_5221,N_3923,N_3989);
or U5222 (N_5222,N_4140,N_4235);
nor U5223 (N_5223,N_4110,N_4497);
nand U5224 (N_5224,N_3854,N_4119);
nand U5225 (N_5225,N_3834,N_3816);
nor U5226 (N_5226,N_4369,N_4094);
or U5227 (N_5227,N_4308,N_4347);
nor U5228 (N_5228,N_4053,N_4299);
and U5229 (N_5229,N_4101,N_3866);
and U5230 (N_5230,N_4047,N_4086);
nor U5231 (N_5231,N_4228,N_4153);
nor U5232 (N_5232,N_3915,N_4002);
or U5233 (N_5233,N_4004,N_4234);
or U5234 (N_5234,N_3785,N_4007);
and U5235 (N_5235,N_4181,N_3901);
xnor U5236 (N_5236,N_4110,N_4281);
nand U5237 (N_5237,N_4085,N_4159);
or U5238 (N_5238,N_4129,N_4025);
xnor U5239 (N_5239,N_3982,N_3803);
or U5240 (N_5240,N_4182,N_4493);
xor U5241 (N_5241,N_3860,N_3760);
and U5242 (N_5242,N_4234,N_3832);
nand U5243 (N_5243,N_4445,N_4419);
and U5244 (N_5244,N_3978,N_4150);
nand U5245 (N_5245,N_4099,N_3757);
nand U5246 (N_5246,N_4363,N_4428);
and U5247 (N_5247,N_3859,N_4065);
or U5248 (N_5248,N_4442,N_3830);
nand U5249 (N_5249,N_4016,N_3861);
or U5250 (N_5250,N_5057,N_4855);
nand U5251 (N_5251,N_5234,N_4861);
xor U5252 (N_5252,N_4710,N_5032);
nand U5253 (N_5253,N_5218,N_5094);
xor U5254 (N_5254,N_4675,N_4956);
and U5255 (N_5255,N_5046,N_5073);
nor U5256 (N_5256,N_5037,N_4909);
nor U5257 (N_5257,N_4862,N_4978);
and U5258 (N_5258,N_4959,N_5161);
nor U5259 (N_5259,N_5059,N_5210);
nand U5260 (N_5260,N_5103,N_4774);
and U5261 (N_5261,N_5199,N_4766);
nand U5262 (N_5262,N_4526,N_4795);
and U5263 (N_5263,N_4874,N_4512);
xor U5264 (N_5264,N_4760,N_4998);
nand U5265 (N_5265,N_5206,N_5130);
or U5266 (N_5266,N_4528,N_5166);
nor U5267 (N_5267,N_4812,N_4727);
and U5268 (N_5268,N_4858,N_5208);
xor U5269 (N_5269,N_4669,N_5101);
nand U5270 (N_5270,N_4676,N_4977);
and U5271 (N_5271,N_4860,N_4896);
xnor U5272 (N_5272,N_5223,N_4993);
nor U5273 (N_5273,N_5027,N_4831);
nor U5274 (N_5274,N_4797,N_4634);
or U5275 (N_5275,N_4563,N_4782);
nor U5276 (N_5276,N_4626,N_4725);
and U5277 (N_5277,N_5061,N_4814);
nand U5278 (N_5278,N_5247,N_4913);
nor U5279 (N_5279,N_5115,N_4648);
xnor U5280 (N_5280,N_4990,N_4531);
and U5281 (N_5281,N_4992,N_5140);
nor U5282 (N_5282,N_5200,N_4728);
xnor U5283 (N_5283,N_5096,N_4985);
and U5284 (N_5284,N_4940,N_5152);
and U5285 (N_5285,N_4566,N_5156);
or U5286 (N_5286,N_5080,N_4951);
and U5287 (N_5287,N_4519,N_4817);
or U5288 (N_5288,N_4661,N_4621);
xor U5289 (N_5289,N_4527,N_5054);
xor U5290 (N_5290,N_5085,N_4771);
xor U5291 (N_5291,N_5207,N_4687);
or U5292 (N_5292,N_5226,N_4640);
and U5293 (N_5293,N_5087,N_5240);
nand U5294 (N_5294,N_4964,N_4847);
xor U5295 (N_5295,N_5246,N_4917);
and U5296 (N_5296,N_4843,N_4561);
nor U5297 (N_5297,N_4942,N_4735);
nor U5298 (N_5298,N_4919,N_5084);
nor U5299 (N_5299,N_4718,N_4800);
and U5300 (N_5300,N_5248,N_4853);
or U5301 (N_5301,N_4813,N_5179);
xor U5302 (N_5302,N_4620,N_4671);
xnor U5303 (N_5303,N_4601,N_4715);
nor U5304 (N_5304,N_5109,N_5201);
xnor U5305 (N_5305,N_5168,N_4918);
nor U5306 (N_5306,N_5058,N_4971);
or U5307 (N_5307,N_4697,N_5172);
nand U5308 (N_5308,N_4598,N_4827);
xor U5309 (N_5309,N_5099,N_5193);
nand U5310 (N_5310,N_5186,N_4741);
nor U5311 (N_5311,N_5146,N_4607);
and U5312 (N_5312,N_4974,N_5159);
xor U5313 (N_5313,N_5078,N_4933);
and U5314 (N_5314,N_4970,N_5178);
xor U5315 (N_5315,N_5129,N_4679);
and U5316 (N_5316,N_4529,N_4820);
or U5317 (N_5317,N_5117,N_5167);
xnor U5318 (N_5318,N_4571,N_5076);
or U5319 (N_5319,N_5092,N_4881);
nor U5320 (N_5320,N_4958,N_4726);
xnor U5321 (N_5321,N_4761,N_4890);
xnor U5322 (N_5322,N_4508,N_5025);
or U5323 (N_5323,N_5197,N_5068);
and U5324 (N_5324,N_4724,N_4844);
nor U5325 (N_5325,N_4744,N_4645);
and U5326 (N_5326,N_4945,N_5072);
nor U5327 (N_5327,N_5018,N_4522);
and U5328 (N_5328,N_5041,N_5143);
and U5329 (N_5329,N_5036,N_4551);
nor U5330 (N_5330,N_4886,N_5162);
nand U5331 (N_5331,N_4574,N_5075);
and U5332 (N_5332,N_5153,N_4712);
or U5333 (N_5333,N_4908,N_4898);
xnor U5334 (N_5334,N_5222,N_5015);
or U5335 (N_5335,N_4547,N_5102);
nor U5336 (N_5336,N_5225,N_4716);
xor U5337 (N_5337,N_4879,N_4805);
and U5338 (N_5338,N_4558,N_4680);
and U5339 (N_5339,N_5031,N_4854);
nor U5340 (N_5340,N_5194,N_4905);
xor U5341 (N_5341,N_4932,N_5147);
nand U5342 (N_5342,N_4511,N_5139);
nor U5343 (N_5343,N_5209,N_5042);
and U5344 (N_5344,N_5128,N_4931);
and U5345 (N_5345,N_4674,N_4962);
nor U5346 (N_5346,N_5136,N_4734);
nor U5347 (N_5347,N_4589,N_4807);
or U5348 (N_5348,N_5034,N_5134);
nand U5349 (N_5349,N_5188,N_5028);
nand U5350 (N_5350,N_5195,N_4901);
and U5351 (N_5351,N_4754,N_5055);
xor U5352 (N_5352,N_4973,N_4891);
xor U5353 (N_5353,N_4723,N_5244);
or U5354 (N_5354,N_4623,N_4586);
nor U5355 (N_5355,N_4729,N_5003);
nor U5356 (N_5356,N_5187,N_5013);
and U5357 (N_5357,N_4757,N_4832);
nand U5358 (N_5358,N_4987,N_4668);
nor U5359 (N_5359,N_4981,N_4767);
and U5360 (N_5360,N_5113,N_4641);
nand U5361 (N_5361,N_4678,N_4644);
xor U5362 (N_5362,N_4949,N_4610);
or U5363 (N_5363,N_5175,N_4880);
and U5364 (N_5364,N_5030,N_4897);
xnor U5365 (N_5365,N_5024,N_5126);
nand U5366 (N_5366,N_4849,N_4836);
and U5367 (N_5367,N_5150,N_4846);
or U5368 (N_5368,N_5064,N_4991);
xor U5369 (N_5369,N_5231,N_4708);
or U5370 (N_5370,N_5163,N_4520);
nand U5371 (N_5371,N_4944,N_5241);
or U5372 (N_5372,N_4632,N_5086);
nor U5373 (N_5373,N_4848,N_5125);
xor U5374 (N_5374,N_4811,N_4694);
nor U5375 (N_5375,N_4752,N_4720);
and U5376 (N_5376,N_5014,N_5141);
and U5377 (N_5377,N_4747,N_4777);
nor U5378 (N_5378,N_4967,N_4906);
nor U5379 (N_5379,N_4762,N_5090);
and U5380 (N_5380,N_4877,N_5051);
xnor U5381 (N_5381,N_4695,N_4525);
or U5382 (N_5382,N_4655,N_4955);
and U5383 (N_5383,N_4732,N_4542);
or U5384 (N_5384,N_4979,N_4592);
and U5385 (N_5385,N_4614,N_4646);
xor U5386 (N_5386,N_4983,N_4530);
nand U5387 (N_5387,N_5007,N_4600);
nor U5388 (N_5388,N_4654,N_4660);
or U5389 (N_5389,N_4873,N_5165);
or U5390 (N_5390,N_4534,N_4662);
nand U5391 (N_5391,N_5052,N_5249);
and U5392 (N_5392,N_4790,N_4915);
nand U5393 (N_5393,N_4587,N_4749);
nand U5394 (N_5394,N_4875,N_4609);
xnor U5395 (N_5395,N_5211,N_4773);
nand U5396 (N_5396,N_4809,N_4535);
nand U5397 (N_5397,N_5144,N_4857);
and U5398 (N_5398,N_5157,N_4840);
nor U5399 (N_5399,N_4622,N_4670);
xor U5400 (N_5400,N_5079,N_4755);
nand U5401 (N_5401,N_4605,N_5082);
or U5402 (N_5402,N_4633,N_5227);
nor U5403 (N_5403,N_4612,N_4930);
nand U5404 (N_5404,N_4546,N_4500);
xnor U5405 (N_5405,N_5012,N_5169);
or U5406 (N_5406,N_5142,N_4579);
and U5407 (N_5407,N_4540,N_4653);
and U5408 (N_5408,N_4871,N_4663);
and U5409 (N_5409,N_4872,N_4794);
and U5410 (N_5410,N_4664,N_5216);
or U5411 (N_5411,N_4988,N_4736);
nor U5412 (N_5412,N_4748,N_5035);
and U5413 (N_5413,N_4883,N_4521);
and U5414 (N_5414,N_4625,N_4939);
nand U5415 (N_5415,N_5050,N_4900);
nor U5416 (N_5416,N_4953,N_5237);
nor U5417 (N_5417,N_4556,N_5033);
xnor U5418 (N_5418,N_4829,N_5121);
nand U5419 (N_5419,N_5077,N_4989);
nor U5420 (N_5420,N_4785,N_5158);
nand U5421 (N_5421,N_4510,N_4709);
xnor U5422 (N_5422,N_4696,N_4681);
nor U5423 (N_5423,N_5095,N_4649);
xnor U5424 (N_5424,N_4851,N_5198);
xnor U5425 (N_5425,N_4544,N_4565);
or U5426 (N_5426,N_5236,N_5056);
nor U5427 (N_5427,N_4801,N_4513);
nand U5428 (N_5428,N_4618,N_5243);
and U5429 (N_5429,N_5174,N_4700);
xor U5430 (N_5430,N_4869,N_4691);
nand U5431 (N_5431,N_5173,N_4714);
and U5432 (N_5432,N_5232,N_4783);
and U5433 (N_5433,N_5016,N_4798);
nor U5434 (N_5434,N_4532,N_4686);
nor U5435 (N_5435,N_4759,N_4580);
and U5436 (N_5436,N_5189,N_4683);
nor U5437 (N_5437,N_4870,N_4509);
xnor U5438 (N_5438,N_5045,N_4786);
and U5439 (N_5439,N_4722,N_4927);
or U5440 (N_5440,N_4845,N_5149);
and U5441 (N_5441,N_5148,N_4789);
and U5442 (N_5442,N_4784,N_5235);
and U5443 (N_5443,N_4799,N_4758);
nand U5444 (N_5444,N_4514,N_4776);
or U5445 (N_5445,N_4611,N_4994);
and U5446 (N_5446,N_4504,N_5040);
nand U5447 (N_5447,N_4667,N_4731);
nand U5448 (N_5448,N_4823,N_4926);
nand U5449 (N_5449,N_4745,N_5132);
or U5450 (N_5450,N_5022,N_4863);
or U5451 (N_5451,N_5047,N_5185);
and U5452 (N_5452,N_4878,N_4980);
xor U5453 (N_5453,N_4515,N_4682);
or U5454 (N_5454,N_4868,N_4608);
and U5455 (N_5455,N_4503,N_4910);
nand U5456 (N_5456,N_5214,N_4772);
and U5457 (N_5457,N_4938,N_4567);
nand U5458 (N_5458,N_4740,N_4637);
nor U5459 (N_5459,N_4575,N_4864);
and U5460 (N_5460,N_5192,N_4577);
nand U5461 (N_5461,N_4775,N_4781);
and U5462 (N_5462,N_5233,N_4582);
nand U5463 (N_5463,N_4924,N_4833);
nor U5464 (N_5464,N_5049,N_4584);
or U5465 (N_5465,N_4912,N_5154);
nand U5466 (N_5466,N_4523,N_4613);
xor U5467 (N_5467,N_4658,N_4719);
and U5468 (N_5468,N_4842,N_4516);
nor U5469 (N_5469,N_4765,N_5212);
nor U5470 (N_5470,N_4717,N_4976);
nand U5471 (N_5471,N_4787,N_4882);
or U5472 (N_5472,N_5017,N_4506);
and U5473 (N_5473,N_4911,N_5088);
nor U5474 (N_5474,N_5093,N_4636);
xnor U5475 (N_5475,N_4538,N_5089);
nand U5476 (N_5476,N_5124,N_4764);
nand U5477 (N_5477,N_4922,N_5038);
nand U5478 (N_5478,N_5123,N_4793);
and U5479 (N_5479,N_4892,N_4585);
nand U5480 (N_5480,N_4803,N_5119);
and U5481 (N_5481,N_4541,N_4756);
nand U5482 (N_5482,N_4884,N_4539);
and U5483 (N_5483,N_5008,N_4835);
nor U5484 (N_5484,N_4562,N_4837);
or U5485 (N_5485,N_5137,N_4665);
xor U5486 (N_5486,N_4689,N_4972);
and U5487 (N_5487,N_4948,N_5006);
nor U5488 (N_5488,N_4867,N_5023);
or U5489 (N_5489,N_4738,N_4619);
or U5490 (N_5490,N_5204,N_5122);
nor U5491 (N_5491,N_4721,N_4965);
nor U5492 (N_5492,N_5005,N_4688);
or U5493 (N_5493,N_4818,N_4631);
and U5494 (N_5494,N_4690,N_4925);
and U5495 (N_5495,N_4583,N_4672);
nand U5496 (N_5496,N_4730,N_4704);
and U5497 (N_5497,N_4802,N_4995);
nand U5498 (N_5498,N_4502,N_5002);
and U5499 (N_5499,N_4916,N_4770);
and U5500 (N_5500,N_4548,N_5021);
nor U5501 (N_5501,N_5228,N_5203);
or U5502 (N_5502,N_4627,N_4692);
xnor U5503 (N_5503,N_4753,N_5107);
or U5504 (N_5504,N_5091,N_5155);
xnor U5505 (N_5505,N_4713,N_5138);
nor U5506 (N_5506,N_4946,N_4570);
nand U5507 (N_5507,N_5081,N_5245);
xnor U5508 (N_5508,N_4824,N_4711);
nor U5509 (N_5509,N_4769,N_5060);
nor U5510 (N_5510,N_5114,N_4739);
xnor U5511 (N_5511,N_5238,N_4652);
or U5512 (N_5512,N_5104,N_5063);
nand U5513 (N_5513,N_5011,N_4921);
or U5514 (N_5514,N_5181,N_5111);
nor U5515 (N_5515,N_4685,N_5120);
nand U5516 (N_5516,N_5066,N_4830);
or U5517 (N_5517,N_4923,N_4865);
nor U5518 (N_5518,N_4635,N_4590);
nand U5519 (N_5519,N_4703,N_4560);
or U5520 (N_5520,N_5108,N_4804);
or U5521 (N_5521,N_5048,N_4596);
or U5522 (N_5522,N_4693,N_4578);
nand U5523 (N_5523,N_5230,N_4763);
xnor U5524 (N_5524,N_5026,N_4996);
or U5525 (N_5525,N_4742,N_4552);
xor U5526 (N_5526,N_4796,N_5171);
or U5527 (N_5527,N_5202,N_4602);
xnor U5528 (N_5528,N_4543,N_4569);
nor U5529 (N_5529,N_5010,N_4572);
nor U5530 (N_5530,N_4969,N_4903);
nand U5531 (N_5531,N_4606,N_5242);
or U5532 (N_5532,N_4705,N_4594);
xor U5533 (N_5533,N_5219,N_4647);
or U5534 (N_5534,N_4555,N_5215);
or U5535 (N_5535,N_4876,N_4986);
or U5536 (N_5536,N_4524,N_4554);
nor U5537 (N_5537,N_4517,N_4894);
nor U5538 (N_5538,N_4624,N_5160);
and U5539 (N_5539,N_4701,N_5029);
xor U5540 (N_5540,N_4656,N_5170);
xor U5541 (N_5541,N_4779,N_5224);
xnor U5542 (N_5542,N_4581,N_4750);
nor U5543 (N_5543,N_4999,N_4549);
nor U5544 (N_5544,N_4642,N_4778);
xor U5545 (N_5545,N_4659,N_5229);
xnor U5546 (N_5546,N_4595,N_5098);
and U5547 (N_5547,N_5133,N_5070);
nor U5548 (N_5548,N_4568,N_4792);
or U5549 (N_5549,N_4960,N_4839);
xnor U5550 (N_5550,N_4591,N_4615);
or U5551 (N_5551,N_5217,N_4698);
nand U5552 (N_5552,N_5164,N_4791);
nor U5553 (N_5553,N_5205,N_4826);
nor U5554 (N_5554,N_4935,N_5004);
or U5555 (N_5555,N_4603,N_4657);
or U5556 (N_5556,N_4997,N_4838);
and U5557 (N_5557,N_4968,N_4628);
and U5558 (N_5558,N_4651,N_4505);
and U5559 (N_5559,N_4780,N_4819);
and U5560 (N_5560,N_4597,N_5135);
or U5561 (N_5561,N_5131,N_5184);
or U5562 (N_5562,N_4961,N_4743);
and U5563 (N_5563,N_5180,N_5177);
and U5564 (N_5564,N_5112,N_5065);
nand U5565 (N_5565,N_4904,N_4617);
nand U5566 (N_5566,N_4950,N_4533);
and U5567 (N_5567,N_4815,N_4593);
xor U5568 (N_5568,N_5220,N_4852);
or U5569 (N_5569,N_4825,N_5190);
and U5570 (N_5570,N_4934,N_5116);
xnor U5571 (N_5571,N_4677,N_5000);
and U5572 (N_5572,N_5069,N_4929);
xor U5573 (N_5573,N_5097,N_4733);
nand U5574 (N_5574,N_4707,N_4936);
nand U5575 (N_5575,N_5221,N_5182);
xor U5576 (N_5576,N_4553,N_4537);
nand U5577 (N_5577,N_4914,N_4599);
or U5578 (N_5578,N_4684,N_4902);
and U5579 (N_5579,N_5009,N_4501);
or U5580 (N_5580,N_4629,N_5118);
nor U5581 (N_5581,N_5196,N_4816);
xor U5582 (N_5582,N_4856,N_4893);
nor U5583 (N_5583,N_5151,N_4937);
nor U5584 (N_5584,N_4887,N_5001);
xnor U5585 (N_5585,N_4810,N_5110);
nand U5586 (N_5586,N_5067,N_5183);
and U5587 (N_5587,N_4536,N_4889);
nand U5588 (N_5588,N_5053,N_4963);
or U5589 (N_5589,N_4841,N_4975);
or U5590 (N_5590,N_4828,N_4643);
nand U5591 (N_5591,N_4639,N_4941);
nor U5592 (N_5592,N_4518,N_4788);
and U5593 (N_5593,N_4545,N_4920);
and U5594 (N_5594,N_5100,N_5039);
and U5595 (N_5595,N_4638,N_4966);
xor U5596 (N_5596,N_4834,N_5106);
and U5597 (N_5597,N_4673,N_4947);
and U5598 (N_5598,N_4822,N_4984);
nand U5599 (N_5599,N_4559,N_4666);
nand U5600 (N_5600,N_5213,N_4630);
and U5601 (N_5601,N_5145,N_5239);
xor U5602 (N_5602,N_4768,N_4573);
or U5603 (N_5603,N_5019,N_4957);
nand U5604 (N_5604,N_5191,N_5074);
nand U5605 (N_5605,N_4588,N_4888);
and U5606 (N_5606,N_4806,N_4859);
xor U5607 (N_5607,N_4885,N_4952);
and U5608 (N_5608,N_4616,N_4507);
nand U5609 (N_5609,N_4907,N_4895);
and U5610 (N_5610,N_5071,N_4850);
nor U5611 (N_5611,N_4866,N_5020);
or U5612 (N_5612,N_4943,N_4982);
nand U5613 (N_5613,N_4576,N_4821);
and U5614 (N_5614,N_5105,N_4564);
or U5615 (N_5615,N_4557,N_4737);
nand U5616 (N_5616,N_5083,N_4746);
nor U5617 (N_5617,N_5062,N_5043);
xor U5618 (N_5618,N_4751,N_4706);
nor U5619 (N_5619,N_4604,N_4808);
xor U5620 (N_5620,N_4550,N_5044);
nand U5621 (N_5621,N_4650,N_4702);
or U5622 (N_5622,N_4928,N_5127);
nand U5623 (N_5623,N_5176,N_4699);
or U5624 (N_5624,N_4899,N_4954);
and U5625 (N_5625,N_4598,N_4704);
nor U5626 (N_5626,N_4789,N_5234);
nand U5627 (N_5627,N_5172,N_5159);
nor U5628 (N_5628,N_4925,N_4871);
and U5629 (N_5629,N_4972,N_4657);
nand U5630 (N_5630,N_5195,N_4945);
nor U5631 (N_5631,N_4909,N_4544);
and U5632 (N_5632,N_4768,N_4566);
nor U5633 (N_5633,N_4902,N_5007);
or U5634 (N_5634,N_5018,N_5144);
and U5635 (N_5635,N_4530,N_5141);
or U5636 (N_5636,N_4615,N_4912);
nand U5637 (N_5637,N_4888,N_5034);
nor U5638 (N_5638,N_4540,N_5144);
nand U5639 (N_5639,N_4536,N_5080);
and U5640 (N_5640,N_5074,N_4834);
nand U5641 (N_5641,N_5079,N_4698);
nand U5642 (N_5642,N_4512,N_4537);
nand U5643 (N_5643,N_4990,N_5120);
and U5644 (N_5644,N_4791,N_4799);
nand U5645 (N_5645,N_4862,N_4523);
and U5646 (N_5646,N_5155,N_4927);
or U5647 (N_5647,N_4969,N_4776);
or U5648 (N_5648,N_4862,N_4764);
or U5649 (N_5649,N_4876,N_4642);
nor U5650 (N_5650,N_5076,N_4995);
or U5651 (N_5651,N_4727,N_4908);
and U5652 (N_5652,N_4579,N_5145);
and U5653 (N_5653,N_4706,N_4692);
and U5654 (N_5654,N_4636,N_5111);
nor U5655 (N_5655,N_4573,N_5010);
or U5656 (N_5656,N_4938,N_5038);
nor U5657 (N_5657,N_4997,N_4594);
xor U5658 (N_5658,N_4953,N_4509);
and U5659 (N_5659,N_4761,N_5205);
and U5660 (N_5660,N_5107,N_4883);
or U5661 (N_5661,N_4563,N_4735);
nand U5662 (N_5662,N_4929,N_4577);
or U5663 (N_5663,N_4938,N_5199);
nand U5664 (N_5664,N_5228,N_4858);
nor U5665 (N_5665,N_4895,N_5094);
nor U5666 (N_5666,N_4971,N_5242);
or U5667 (N_5667,N_4989,N_5037);
and U5668 (N_5668,N_5088,N_5086);
nor U5669 (N_5669,N_4673,N_4964);
and U5670 (N_5670,N_5185,N_4931);
nor U5671 (N_5671,N_5114,N_4680);
or U5672 (N_5672,N_5164,N_5093);
nor U5673 (N_5673,N_4758,N_5214);
nor U5674 (N_5674,N_5227,N_5183);
xor U5675 (N_5675,N_4817,N_4752);
and U5676 (N_5676,N_5206,N_5177);
and U5677 (N_5677,N_4881,N_4777);
xor U5678 (N_5678,N_4971,N_4878);
xor U5679 (N_5679,N_4566,N_5205);
and U5680 (N_5680,N_4644,N_4760);
nand U5681 (N_5681,N_4914,N_4902);
or U5682 (N_5682,N_4856,N_4777);
and U5683 (N_5683,N_5220,N_5164);
or U5684 (N_5684,N_5010,N_4854);
nand U5685 (N_5685,N_4544,N_5075);
nand U5686 (N_5686,N_5067,N_4705);
xor U5687 (N_5687,N_4943,N_4664);
xnor U5688 (N_5688,N_4766,N_4701);
xor U5689 (N_5689,N_5089,N_4648);
nand U5690 (N_5690,N_4783,N_4709);
nand U5691 (N_5691,N_4525,N_5142);
nand U5692 (N_5692,N_4574,N_5168);
or U5693 (N_5693,N_5050,N_4953);
nand U5694 (N_5694,N_4805,N_4756);
or U5695 (N_5695,N_4877,N_4636);
or U5696 (N_5696,N_4681,N_4979);
or U5697 (N_5697,N_4649,N_4989);
xnor U5698 (N_5698,N_5163,N_4589);
and U5699 (N_5699,N_5096,N_4515);
xor U5700 (N_5700,N_4842,N_4748);
and U5701 (N_5701,N_4726,N_4661);
or U5702 (N_5702,N_4706,N_4756);
and U5703 (N_5703,N_4794,N_4739);
nand U5704 (N_5704,N_5063,N_5163);
or U5705 (N_5705,N_5028,N_4545);
or U5706 (N_5706,N_4786,N_5097);
nor U5707 (N_5707,N_4909,N_5023);
nand U5708 (N_5708,N_5019,N_4554);
nor U5709 (N_5709,N_4734,N_4993);
nand U5710 (N_5710,N_4977,N_5211);
and U5711 (N_5711,N_4601,N_4654);
xor U5712 (N_5712,N_4590,N_4532);
or U5713 (N_5713,N_5155,N_5013);
xor U5714 (N_5714,N_4913,N_4756);
nor U5715 (N_5715,N_5172,N_5125);
and U5716 (N_5716,N_5008,N_5175);
nand U5717 (N_5717,N_4765,N_4757);
and U5718 (N_5718,N_4724,N_4822);
nand U5719 (N_5719,N_5103,N_4574);
xnor U5720 (N_5720,N_5201,N_4950);
and U5721 (N_5721,N_4626,N_5191);
and U5722 (N_5722,N_4976,N_5194);
nor U5723 (N_5723,N_5112,N_4685);
xnor U5724 (N_5724,N_4992,N_5010);
xnor U5725 (N_5725,N_5202,N_5163);
xnor U5726 (N_5726,N_5000,N_5074);
or U5727 (N_5727,N_4636,N_5009);
nand U5728 (N_5728,N_4749,N_4644);
nand U5729 (N_5729,N_4696,N_5037);
nor U5730 (N_5730,N_4632,N_4577);
and U5731 (N_5731,N_5221,N_4968);
nand U5732 (N_5732,N_5083,N_4913);
nand U5733 (N_5733,N_4595,N_4822);
nor U5734 (N_5734,N_4753,N_4659);
or U5735 (N_5735,N_4568,N_4576);
nand U5736 (N_5736,N_5169,N_5052);
nor U5737 (N_5737,N_5058,N_4515);
or U5738 (N_5738,N_5146,N_5116);
and U5739 (N_5739,N_5209,N_4671);
or U5740 (N_5740,N_4530,N_4780);
nor U5741 (N_5741,N_5014,N_5176);
nor U5742 (N_5742,N_5145,N_5085);
xor U5743 (N_5743,N_4782,N_4628);
xor U5744 (N_5744,N_4887,N_5190);
or U5745 (N_5745,N_4646,N_5204);
nor U5746 (N_5746,N_4862,N_5231);
xor U5747 (N_5747,N_4672,N_5212);
xnor U5748 (N_5748,N_4909,N_5124);
and U5749 (N_5749,N_4608,N_4504);
and U5750 (N_5750,N_5013,N_4639);
and U5751 (N_5751,N_4774,N_5208);
and U5752 (N_5752,N_4828,N_4978);
or U5753 (N_5753,N_4542,N_4847);
or U5754 (N_5754,N_4596,N_5229);
nor U5755 (N_5755,N_5161,N_4942);
xnor U5756 (N_5756,N_5102,N_4606);
nor U5757 (N_5757,N_4630,N_4566);
and U5758 (N_5758,N_4659,N_5200);
nand U5759 (N_5759,N_5234,N_4743);
xnor U5760 (N_5760,N_4979,N_4674);
or U5761 (N_5761,N_4935,N_4543);
xor U5762 (N_5762,N_4525,N_5195);
xor U5763 (N_5763,N_5194,N_4773);
and U5764 (N_5764,N_4977,N_4882);
and U5765 (N_5765,N_4828,N_4881);
xor U5766 (N_5766,N_5222,N_4511);
or U5767 (N_5767,N_4919,N_4672);
and U5768 (N_5768,N_4579,N_5247);
nand U5769 (N_5769,N_4871,N_5001);
or U5770 (N_5770,N_4790,N_4914);
or U5771 (N_5771,N_4665,N_5197);
nand U5772 (N_5772,N_5109,N_5112);
and U5773 (N_5773,N_5212,N_4930);
xnor U5774 (N_5774,N_4945,N_5012);
nand U5775 (N_5775,N_4719,N_5186);
nor U5776 (N_5776,N_4976,N_5052);
xor U5777 (N_5777,N_5026,N_4922);
or U5778 (N_5778,N_4924,N_5014);
nand U5779 (N_5779,N_4832,N_4894);
xnor U5780 (N_5780,N_4585,N_4804);
and U5781 (N_5781,N_4748,N_4872);
and U5782 (N_5782,N_4876,N_5111);
nand U5783 (N_5783,N_4898,N_4606);
nor U5784 (N_5784,N_4939,N_4941);
or U5785 (N_5785,N_5208,N_4568);
or U5786 (N_5786,N_4839,N_4668);
and U5787 (N_5787,N_5031,N_4728);
or U5788 (N_5788,N_4868,N_4631);
xnor U5789 (N_5789,N_4646,N_5155);
xor U5790 (N_5790,N_5125,N_4925);
nor U5791 (N_5791,N_4526,N_4675);
nor U5792 (N_5792,N_5103,N_4941);
nor U5793 (N_5793,N_4866,N_4780);
and U5794 (N_5794,N_4681,N_5080);
xor U5795 (N_5795,N_4510,N_5079);
or U5796 (N_5796,N_4502,N_4518);
and U5797 (N_5797,N_4734,N_5118);
xor U5798 (N_5798,N_5056,N_5201);
and U5799 (N_5799,N_4982,N_4717);
and U5800 (N_5800,N_4869,N_4723);
nor U5801 (N_5801,N_4785,N_4524);
nand U5802 (N_5802,N_4665,N_5059);
and U5803 (N_5803,N_5053,N_5047);
nor U5804 (N_5804,N_4870,N_4524);
xnor U5805 (N_5805,N_4843,N_5232);
or U5806 (N_5806,N_4831,N_4955);
nand U5807 (N_5807,N_4785,N_5157);
nand U5808 (N_5808,N_4976,N_5050);
and U5809 (N_5809,N_5208,N_5203);
xnor U5810 (N_5810,N_4740,N_4768);
nor U5811 (N_5811,N_4690,N_4994);
nand U5812 (N_5812,N_4842,N_5068);
or U5813 (N_5813,N_4974,N_5063);
nand U5814 (N_5814,N_4745,N_4995);
or U5815 (N_5815,N_4732,N_5008);
nand U5816 (N_5816,N_4926,N_4903);
nand U5817 (N_5817,N_4803,N_4903);
nor U5818 (N_5818,N_4804,N_5018);
and U5819 (N_5819,N_4762,N_4617);
xnor U5820 (N_5820,N_5177,N_4603);
or U5821 (N_5821,N_4926,N_5095);
nor U5822 (N_5822,N_5097,N_4613);
nand U5823 (N_5823,N_5083,N_4737);
xnor U5824 (N_5824,N_4915,N_4507);
and U5825 (N_5825,N_4625,N_4611);
and U5826 (N_5826,N_4662,N_4558);
or U5827 (N_5827,N_5164,N_4819);
nor U5828 (N_5828,N_4990,N_4882);
or U5829 (N_5829,N_4974,N_4725);
xnor U5830 (N_5830,N_4826,N_4503);
or U5831 (N_5831,N_4735,N_4637);
nor U5832 (N_5832,N_5240,N_4688);
and U5833 (N_5833,N_4914,N_5070);
or U5834 (N_5834,N_4951,N_4953);
nand U5835 (N_5835,N_4560,N_4702);
and U5836 (N_5836,N_4990,N_4808);
or U5837 (N_5837,N_4854,N_5038);
and U5838 (N_5838,N_5194,N_4808);
nand U5839 (N_5839,N_4812,N_4777);
xor U5840 (N_5840,N_4717,N_4770);
or U5841 (N_5841,N_4596,N_5034);
nor U5842 (N_5842,N_5182,N_4606);
or U5843 (N_5843,N_5180,N_5055);
nand U5844 (N_5844,N_4667,N_5203);
nor U5845 (N_5845,N_4721,N_5125);
xor U5846 (N_5846,N_5015,N_4869);
and U5847 (N_5847,N_4765,N_4501);
and U5848 (N_5848,N_5011,N_5157);
nor U5849 (N_5849,N_4727,N_4871);
or U5850 (N_5850,N_5117,N_4553);
or U5851 (N_5851,N_4906,N_5188);
nor U5852 (N_5852,N_5202,N_4671);
or U5853 (N_5853,N_5227,N_4857);
or U5854 (N_5854,N_4620,N_5190);
xnor U5855 (N_5855,N_4742,N_4821);
or U5856 (N_5856,N_4729,N_4770);
xnor U5857 (N_5857,N_4927,N_5126);
xnor U5858 (N_5858,N_4940,N_4544);
xnor U5859 (N_5859,N_4908,N_5148);
nor U5860 (N_5860,N_5146,N_5153);
xor U5861 (N_5861,N_4996,N_5199);
nand U5862 (N_5862,N_5018,N_5086);
nand U5863 (N_5863,N_4943,N_5106);
nor U5864 (N_5864,N_5034,N_4677);
or U5865 (N_5865,N_5087,N_4830);
xnor U5866 (N_5866,N_4614,N_4839);
nand U5867 (N_5867,N_5096,N_5133);
nor U5868 (N_5868,N_4931,N_4620);
nor U5869 (N_5869,N_4984,N_5110);
nand U5870 (N_5870,N_4885,N_5246);
nand U5871 (N_5871,N_5154,N_5190);
nand U5872 (N_5872,N_4676,N_4647);
or U5873 (N_5873,N_4948,N_4852);
and U5874 (N_5874,N_4989,N_4694);
xnor U5875 (N_5875,N_4675,N_5107);
xor U5876 (N_5876,N_4670,N_4960);
xor U5877 (N_5877,N_4643,N_5024);
nand U5878 (N_5878,N_4655,N_4700);
or U5879 (N_5879,N_5085,N_4632);
and U5880 (N_5880,N_4762,N_4880);
nand U5881 (N_5881,N_5033,N_4543);
and U5882 (N_5882,N_4923,N_5112);
nand U5883 (N_5883,N_4647,N_4535);
and U5884 (N_5884,N_5235,N_4660);
nand U5885 (N_5885,N_5062,N_4944);
or U5886 (N_5886,N_5216,N_4637);
or U5887 (N_5887,N_4746,N_5155);
nor U5888 (N_5888,N_5139,N_5093);
or U5889 (N_5889,N_5097,N_5046);
xor U5890 (N_5890,N_4782,N_4827);
and U5891 (N_5891,N_5016,N_4520);
or U5892 (N_5892,N_4760,N_4797);
nand U5893 (N_5893,N_4827,N_4770);
nor U5894 (N_5894,N_5219,N_4833);
and U5895 (N_5895,N_4981,N_5132);
xnor U5896 (N_5896,N_4512,N_5067);
xnor U5897 (N_5897,N_4929,N_5060);
xor U5898 (N_5898,N_5154,N_4782);
or U5899 (N_5899,N_4604,N_4860);
xnor U5900 (N_5900,N_4582,N_5065);
nor U5901 (N_5901,N_4866,N_4822);
xor U5902 (N_5902,N_4856,N_5121);
and U5903 (N_5903,N_4744,N_4907);
nor U5904 (N_5904,N_4953,N_4934);
and U5905 (N_5905,N_4830,N_4811);
nor U5906 (N_5906,N_4604,N_5130);
xnor U5907 (N_5907,N_4807,N_4861);
nand U5908 (N_5908,N_5195,N_5176);
or U5909 (N_5909,N_4752,N_5124);
xor U5910 (N_5910,N_4536,N_4615);
or U5911 (N_5911,N_4911,N_4503);
or U5912 (N_5912,N_4733,N_4821);
or U5913 (N_5913,N_4961,N_5237);
xnor U5914 (N_5914,N_4710,N_4690);
or U5915 (N_5915,N_4883,N_4610);
xor U5916 (N_5916,N_4585,N_4902);
or U5917 (N_5917,N_4964,N_4586);
and U5918 (N_5918,N_4949,N_4772);
and U5919 (N_5919,N_4679,N_4808);
nand U5920 (N_5920,N_5043,N_4825);
or U5921 (N_5921,N_4956,N_4554);
and U5922 (N_5922,N_4717,N_4860);
or U5923 (N_5923,N_5028,N_4923);
xor U5924 (N_5924,N_4748,N_4533);
or U5925 (N_5925,N_4533,N_4849);
xnor U5926 (N_5926,N_4905,N_5037);
nand U5927 (N_5927,N_4630,N_4536);
nor U5928 (N_5928,N_4649,N_4744);
or U5929 (N_5929,N_4968,N_4825);
nand U5930 (N_5930,N_4821,N_5008);
xor U5931 (N_5931,N_5187,N_4745);
and U5932 (N_5932,N_4700,N_4503);
and U5933 (N_5933,N_4856,N_4911);
xor U5934 (N_5934,N_4943,N_5010);
or U5935 (N_5935,N_4889,N_5210);
nand U5936 (N_5936,N_4755,N_4655);
or U5937 (N_5937,N_4649,N_4844);
and U5938 (N_5938,N_5002,N_4929);
nand U5939 (N_5939,N_5008,N_5184);
or U5940 (N_5940,N_4582,N_4736);
nor U5941 (N_5941,N_4829,N_5050);
or U5942 (N_5942,N_4617,N_4767);
or U5943 (N_5943,N_5008,N_4631);
nor U5944 (N_5944,N_5185,N_5021);
nor U5945 (N_5945,N_4711,N_4545);
nor U5946 (N_5946,N_4877,N_5179);
and U5947 (N_5947,N_4744,N_4677);
nor U5948 (N_5948,N_4898,N_5058);
and U5949 (N_5949,N_4865,N_5048);
nand U5950 (N_5950,N_4841,N_4505);
xor U5951 (N_5951,N_4576,N_4659);
or U5952 (N_5952,N_4712,N_5077);
nor U5953 (N_5953,N_4549,N_4700);
and U5954 (N_5954,N_4550,N_4800);
or U5955 (N_5955,N_4831,N_4933);
and U5956 (N_5956,N_4991,N_4573);
nand U5957 (N_5957,N_4569,N_4741);
or U5958 (N_5958,N_5083,N_4776);
nand U5959 (N_5959,N_5168,N_5053);
and U5960 (N_5960,N_4624,N_5152);
nand U5961 (N_5961,N_5143,N_4969);
and U5962 (N_5962,N_5239,N_4854);
and U5963 (N_5963,N_4881,N_5144);
nand U5964 (N_5964,N_4973,N_4967);
xnor U5965 (N_5965,N_4587,N_4692);
nor U5966 (N_5966,N_5073,N_4554);
and U5967 (N_5967,N_4885,N_4817);
or U5968 (N_5968,N_5194,N_4943);
xor U5969 (N_5969,N_4758,N_4722);
xnor U5970 (N_5970,N_4584,N_4540);
or U5971 (N_5971,N_4946,N_5041);
nor U5972 (N_5972,N_4832,N_4623);
nand U5973 (N_5973,N_5035,N_5013);
or U5974 (N_5974,N_5044,N_4592);
xor U5975 (N_5975,N_5172,N_5232);
xnor U5976 (N_5976,N_4923,N_4930);
xnor U5977 (N_5977,N_5211,N_4602);
or U5978 (N_5978,N_4777,N_5020);
or U5979 (N_5979,N_4708,N_5238);
nand U5980 (N_5980,N_4562,N_4647);
and U5981 (N_5981,N_5198,N_4896);
nor U5982 (N_5982,N_5051,N_4573);
and U5983 (N_5983,N_4666,N_4542);
nand U5984 (N_5984,N_4608,N_4731);
and U5985 (N_5985,N_5143,N_5031);
xor U5986 (N_5986,N_5237,N_4712);
nor U5987 (N_5987,N_4803,N_5060);
nand U5988 (N_5988,N_4562,N_4890);
nand U5989 (N_5989,N_4621,N_5110);
or U5990 (N_5990,N_4790,N_4852);
xnor U5991 (N_5991,N_4658,N_4608);
or U5992 (N_5992,N_4686,N_4582);
xor U5993 (N_5993,N_4955,N_4667);
nand U5994 (N_5994,N_5013,N_4734);
xnor U5995 (N_5995,N_5141,N_5149);
xnor U5996 (N_5996,N_5145,N_4768);
nand U5997 (N_5997,N_4855,N_4646);
xor U5998 (N_5998,N_4840,N_4833);
nor U5999 (N_5999,N_4801,N_4602);
nand U6000 (N_6000,N_5468,N_5529);
xor U6001 (N_6001,N_5258,N_5405);
nand U6002 (N_6002,N_5677,N_5358);
nand U6003 (N_6003,N_5997,N_5985);
and U6004 (N_6004,N_5304,N_5667);
or U6005 (N_6005,N_5681,N_5607);
nand U6006 (N_6006,N_5673,N_5441);
and U6007 (N_6007,N_5579,N_5920);
xor U6008 (N_6008,N_5551,N_5763);
nor U6009 (N_6009,N_5801,N_5438);
and U6010 (N_6010,N_5538,N_5302);
and U6011 (N_6011,N_5996,N_5932);
nor U6012 (N_6012,N_5444,N_5622);
or U6013 (N_6013,N_5783,N_5536);
nor U6014 (N_6014,N_5955,N_5994);
nand U6015 (N_6015,N_5824,N_5850);
nand U6016 (N_6016,N_5612,N_5715);
and U6017 (N_6017,N_5528,N_5696);
nor U6018 (N_6018,N_5625,N_5534);
or U6019 (N_6019,N_5657,N_5694);
nand U6020 (N_6020,N_5706,N_5780);
xor U6021 (N_6021,N_5383,N_5844);
nand U6022 (N_6022,N_5627,N_5557);
nor U6023 (N_6023,N_5718,N_5922);
or U6024 (N_6024,N_5340,N_5788);
xor U6025 (N_6025,N_5930,N_5290);
or U6026 (N_6026,N_5637,N_5511);
nand U6027 (N_6027,N_5581,N_5375);
or U6028 (N_6028,N_5870,N_5835);
nand U6029 (N_6029,N_5826,N_5466);
or U6030 (N_6030,N_5273,N_5446);
and U6031 (N_6031,N_5613,N_5286);
xor U6032 (N_6032,N_5815,N_5717);
nand U6033 (N_6033,N_5900,N_5882);
nor U6034 (N_6034,N_5682,N_5250);
xor U6035 (N_6035,N_5925,N_5705);
or U6036 (N_6036,N_5561,N_5614);
nand U6037 (N_6037,N_5431,N_5299);
nor U6038 (N_6038,N_5811,N_5867);
or U6039 (N_6039,N_5336,N_5838);
nand U6040 (N_6040,N_5411,N_5828);
xor U6041 (N_6041,N_5585,N_5822);
nand U6042 (N_6042,N_5461,N_5751);
and U6043 (N_6043,N_5573,N_5460);
xnor U6044 (N_6044,N_5889,N_5720);
xnor U6045 (N_6045,N_5301,N_5496);
and U6046 (N_6046,N_5753,N_5542);
xnor U6047 (N_6047,N_5470,N_5965);
nor U6048 (N_6048,N_5387,N_5707);
and U6049 (N_6049,N_5523,N_5531);
nor U6050 (N_6050,N_5426,N_5962);
and U6051 (N_6051,N_5728,N_5462);
nor U6052 (N_6052,N_5685,N_5265);
nor U6053 (N_6053,N_5809,N_5799);
and U6054 (N_6054,N_5797,N_5660);
or U6055 (N_6055,N_5597,N_5908);
xnor U6056 (N_6056,N_5964,N_5782);
nand U6057 (N_6057,N_5634,N_5623);
nor U6058 (N_6058,N_5862,N_5888);
nor U6059 (N_6059,N_5818,N_5716);
and U6060 (N_6060,N_5476,N_5594);
nor U6061 (N_6061,N_5562,N_5356);
and U6062 (N_6062,N_5950,N_5598);
and U6063 (N_6063,N_5544,N_5732);
and U6064 (N_6064,N_5848,N_5734);
or U6065 (N_6065,N_5432,N_5812);
nand U6066 (N_6066,N_5568,N_5400);
nand U6067 (N_6067,N_5659,N_5784);
xnor U6068 (N_6068,N_5467,N_5686);
and U6069 (N_6069,N_5790,N_5399);
nand U6070 (N_6070,N_5272,N_5830);
nor U6071 (N_6071,N_5499,N_5892);
and U6072 (N_6072,N_5669,N_5516);
and U6073 (N_6073,N_5970,N_5498);
or U6074 (N_6074,N_5390,N_5695);
xnor U6075 (N_6075,N_5591,N_5719);
nand U6076 (N_6076,N_5646,N_5367);
nor U6077 (N_6077,N_5891,N_5588);
nor U6078 (N_6078,N_5342,N_5972);
and U6079 (N_6079,N_5554,N_5624);
and U6080 (N_6080,N_5368,N_5877);
nand U6081 (N_6081,N_5550,N_5449);
xnor U6082 (N_6082,N_5934,N_5580);
nand U6083 (N_6083,N_5522,N_5979);
nor U6084 (N_6084,N_5350,N_5424);
xnor U6085 (N_6085,N_5495,N_5626);
xnor U6086 (N_6086,N_5911,N_5963);
or U6087 (N_6087,N_5489,N_5312);
nand U6088 (N_6088,N_5451,N_5689);
nand U6089 (N_6089,N_5491,N_5372);
and U6090 (N_6090,N_5916,N_5337);
or U6091 (N_6091,N_5297,N_5709);
nand U6092 (N_6092,N_5683,N_5508);
nand U6093 (N_6093,N_5457,N_5282);
xnor U6094 (N_6094,N_5430,N_5989);
or U6095 (N_6095,N_5703,N_5280);
nor U6096 (N_6096,N_5354,N_5629);
or U6097 (N_6097,N_5725,N_5558);
nor U6098 (N_6098,N_5913,N_5519);
and U6099 (N_6099,N_5264,N_5803);
or U6100 (N_6100,N_5982,N_5262);
or U6101 (N_6101,N_5688,N_5611);
xnor U6102 (N_6102,N_5313,N_5795);
xnor U6103 (N_6103,N_5714,N_5915);
nand U6104 (N_6104,N_5408,N_5565);
nand U6105 (N_6105,N_5310,N_5764);
or U6106 (N_6106,N_5663,N_5933);
or U6107 (N_6107,N_5546,N_5407);
or U6108 (N_6108,N_5630,N_5724);
nor U6109 (N_6109,N_5307,N_5700);
nand U6110 (N_6110,N_5593,N_5995);
or U6111 (N_6111,N_5761,N_5991);
and U6112 (N_6112,N_5391,N_5287);
xor U6113 (N_6113,N_5279,N_5873);
xor U6114 (N_6114,N_5566,N_5890);
nand U6115 (N_6115,N_5649,N_5886);
or U6116 (N_6116,N_5404,N_5481);
nand U6117 (N_6117,N_5482,N_5604);
nand U6118 (N_6118,N_5841,N_5907);
xor U6119 (N_6119,N_5652,N_5434);
and U6120 (N_6120,N_5447,N_5608);
and U6121 (N_6121,N_5276,N_5417);
nor U6122 (N_6122,N_5433,N_5651);
xnor U6123 (N_6123,N_5628,N_5768);
and U6124 (N_6124,N_5693,N_5535);
xnor U6125 (N_6125,N_5993,N_5545);
xnor U6126 (N_6126,N_5373,N_5345);
nand U6127 (N_6127,N_5807,N_5800);
or U6128 (N_6128,N_5261,N_5733);
or U6129 (N_6129,N_5300,N_5760);
nor U6130 (N_6130,N_5474,N_5515);
and U6131 (N_6131,N_5389,N_5757);
nand U6132 (N_6132,N_5382,N_5395);
and U6133 (N_6133,N_5638,N_5854);
nand U6134 (N_6134,N_5817,N_5746);
xnor U6135 (N_6135,N_5394,N_5569);
or U6136 (N_6136,N_5269,N_5931);
or U6137 (N_6137,N_5619,N_5602);
or U6138 (N_6138,N_5610,N_5284);
nand U6139 (N_6139,N_5392,N_5819);
xor U6140 (N_6140,N_5855,N_5315);
and U6141 (N_6141,N_5324,N_5338);
nor U6142 (N_6142,N_5712,N_5567);
nand U6143 (N_6143,N_5874,N_5277);
nand U6144 (N_6144,N_5289,N_5947);
or U6145 (N_6145,N_5547,N_5865);
or U6146 (N_6146,N_5737,N_5906);
nand U6147 (N_6147,N_5633,N_5251);
nand U6148 (N_6148,N_5736,N_5977);
and U6149 (N_6149,N_5897,N_5512);
xor U6150 (N_6150,N_5999,N_5674);
or U6151 (N_6151,N_5770,N_5420);
nor U6152 (N_6152,N_5257,N_5750);
xor U6153 (N_6153,N_5314,N_5576);
and U6154 (N_6154,N_5926,N_5339);
xnor U6155 (N_6155,N_5923,N_5465);
nor U6156 (N_6156,N_5921,N_5679);
nand U6157 (N_6157,N_5487,N_5548);
nand U6158 (N_6158,N_5332,N_5747);
xor U6159 (N_6159,N_5680,N_5283);
xor U6160 (N_6160,N_5857,N_5653);
xor U6161 (N_6161,N_5692,N_5904);
nand U6162 (N_6162,N_5861,N_5268);
xor U6163 (N_6163,N_5978,N_5412);
xnor U6164 (N_6164,N_5928,N_5988);
nand U6165 (N_6165,N_5912,N_5735);
and U6166 (N_6166,N_5590,N_5829);
nor U6167 (N_6167,N_5666,N_5423);
nand U6168 (N_6168,N_5506,N_5293);
and U6169 (N_6169,N_5296,N_5847);
nand U6170 (N_6170,N_5401,N_5518);
xor U6171 (N_6171,N_5909,N_5924);
nor U6172 (N_6172,N_5259,N_5537);
or U6173 (N_6173,N_5274,N_5364);
nand U6174 (N_6174,N_5946,N_5502);
nand U6175 (N_6175,N_5976,N_5710);
nor U6176 (N_6176,N_5871,N_5632);
or U6177 (N_6177,N_5295,N_5642);
xnor U6178 (N_6178,N_5899,N_5843);
or U6179 (N_6179,N_5959,N_5486);
nand U6180 (N_6180,N_5351,N_5984);
nor U6181 (N_6181,N_5986,N_5530);
nand U6182 (N_6182,N_5472,N_5675);
or U6183 (N_6183,N_5406,N_5344);
nor U6184 (N_6184,N_5553,N_5776);
nand U6185 (N_6185,N_5347,N_5388);
and U6186 (N_6186,N_5883,N_5773);
xnor U6187 (N_6187,N_5559,N_5766);
and U6188 (N_6188,N_5587,N_5731);
xor U6189 (N_6189,N_5664,N_5458);
nor U6190 (N_6190,N_5656,N_5325);
xor U6191 (N_6191,N_5943,N_5371);
or U6192 (N_6192,N_5644,N_5711);
xor U6193 (N_6193,N_5549,N_5343);
nand U6194 (N_6194,N_5464,N_5599);
or U6195 (N_6195,N_5798,N_5601);
nor U6196 (N_6196,N_5285,N_5836);
and U6197 (N_6197,N_5771,N_5298);
xor U6198 (N_6198,N_5386,N_5839);
xor U6199 (N_6199,N_5759,N_5729);
or U6200 (N_6200,N_5856,N_5514);
and U6201 (N_6201,N_5501,N_5456);
or U6202 (N_6202,N_5742,N_5333);
nor U6203 (N_6203,N_5526,N_5589);
or U6204 (N_6204,N_5256,N_5267);
nor U6205 (N_6205,N_5863,N_5439);
and U6206 (N_6206,N_5524,N_5306);
nor U6207 (N_6207,N_5834,N_5485);
or U6208 (N_6208,N_5321,N_5577);
xnor U6209 (N_6209,N_5951,N_5416);
nand U6210 (N_6210,N_5945,N_5254);
xor U6211 (N_6211,N_5748,N_5318);
and U6212 (N_6212,N_5713,N_5403);
or U6213 (N_6213,N_5749,N_5702);
and U6214 (N_6214,N_5918,N_5635);
and U6215 (N_6215,N_5820,N_5381);
nor U6216 (N_6216,N_5308,N_5992);
nand U6217 (N_6217,N_5410,N_5435);
xor U6218 (N_6218,N_5596,N_5840);
nor U6219 (N_6219,N_5492,N_5726);
and U6220 (N_6220,N_5473,N_5291);
or U6221 (N_6221,N_5641,N_5661);
nand U6222 (N_6222,N_5505,N_5582);
xnor U6223 (N_6223,N_5958,N_5691);
xor U6224 (N_6224,N_5743,N_5378);
xnor U6225 (N_6225,N_5754,N_5459);
nand U6226 (N_6226,N_5796,N_5429);
nor U6227 (N_6227,N_5758,N_5781);
and U6228 (N_6228,N_5357,N_5805);
xnor U6229 (N_6229,N_5353,N_5821);
nor U6230 (N_6230,N_5440,N_5377);
xor U6231 (N_6231,N_5436,N_5366);
xor U6232 (N_6232,N_5937,N_5939);
nor U6233 (N_6233,N_5876,N_5775);
nand U6234 (N_6234,N_5833,N_5935);
or U6235 (N_6235,N_5842,N_5393);
nor U6236 (N_6236,N_5359,N_5563);
nor U6237 (N_6237,N_5330,N_5636);
xor U6238 (N_6238,N_5755,N_5520);
and U6239 (N_6239,N_5278,N_5902);
nand U6240 (N_6240,N_5827,N_5360);
xor U6241 (N_6241,N_5510,N_5645);
or U6242 (N_6242,N_5415,N_5252);
and U6243 (N_6243,N_5648,N_5885);
nor U6244 (N_6244,N_5592,N_5525);
and U6245 (N_6245,N_5665,N_5319);
or U6246 (N_6246,N_5793,N_5288);
xnor U6247 (N_6247,N_5570,N_5938);
xor U6248 (N_6248,N_5864,N_5334);
nand U6249 (N_6249,N_5521,N_5872);
nand U6250 (N_6250,N_5650,N_5739);
and U6251 (N_6251,N_5445,N_5898);
or U6252 (N_6252,N_5969,N_5341);
xor U6253 (N_6253,N_5957,N_5352);
nand U6254 (N_6254,N_5309,N_5671);
xnor U6255 (N_6255,N_5832,N_5294);
nor U6256 (N_6256,N_5777,N_5363);
nor U6257 (N_6257,N_5572,N_5361);
xor U6258 (N_6258,N_5980,N_5896);
nor U6259 (N_6259,N_5794,N_5500);
xnor U6260 (N_6260,N_5413,N_5533);
nand U6261 (N_6261,N_5949,N_5328);
xnor U6262 (N_6262,N_5831,N_5575);
xor U6263 (N_6263,N_5253,N_5745);
and U6264 (N_6264,N_5956,N_5397);
and U6265 (N_6265,N_5609,N_5376);
nand U6266 (N_6266,N_5884,N_5584);
or U6267 (N_6267,N_5981,N_5792);
and U6268 (N_6268,N_5621,N_5418);
nand U6269 (N_6269,N_5655,N_5849);
nor U6270 (N_6270,N_5292,N_5605);
nand U6271 (N_6271,N_5603,N_5973);
nor U6272 (N_6272,N_5813,N_5668);
xnor U6273 (N_6273,N_5443,N_5654);
xnor U6274 (N_6274,N_5756,N_5425);
xnor U6275 (N_6275,N_5823,N_5769);
nand U6276 (N_6276,N_5852,N_5452);
xnor U6277 (N_6277,N_5708,N_5851);
xor U6278 (N_6278,N_5987,N_5966);
xor U6279 (N_6279,N_5539,N_5741);
and U6280 (N_6280,N_5600,N_5369);
nand U6281 (N_6281,N_5914,N_5868);
xor U6282 (N_6282,N_5929,N_5260);
nor U6283 (N_6283,N_5952,N_5471);
and U6284 (N_6284,N_5428,N_5878);
and U6285 (N_6285,N_5860,N_5422);
xor U6286 (N_6286,N_5774,N_5846);
xor U6287 (N_6287,N_5374,N_5323);
nor U6288 (N_6288,N_5779,N_5697);
or U6289 (N_6289,N_5327,N_5905);
and U6290 (N_6290,N_5331,N_5453);
nor U6291 (N_6291,N_5606,N_5786);
xor U6292 (N_6292,N_5701,N_5647);
nor U6293 (N_6293,N_5617,N_5527);
and U6294 (N_6294,N_5483,N_5990);
nor U6295 (N_6295,N_5772,N_5919);
xnor U6296 (N_6296,N_5640,N_5463);
nand U6297 (N_6297,N_5311,N_5355);
or U6298 (N_6298,N_5478,N_5998);
nor U6299 (N_6299,N_5414,N_5560);
or U6300 (N_6300,N_5936,N_5541);
nand U6301 (N_6301,N_5326,N_5266);
or U6302 (N_6302,N_5532,N_5643);
nand U6303 (N_6303,N_5722,N_5879);
nand U6304 (N_6304,N_5574,N_5903);
and U6305 (N_6305,N_5479,N_5493);
nand U6306 (N_6306,N_5927,N_5362);
or U6307 (N_6307,N_5942,N_5762);
xor U6308 (N_6308,N_5837,N_5730);
xor U6309 (N_6309,N_5670,N_5480);
xor U6310 (N_6310,N_5421,N_5765);
and U6311 (N_6311,N_5586,N_5419);
and U6312 (N_6312,N_5954,N_5804);
or U6313 (N_6313,N_5975,N_5895);
nor U6314 (N_6314,N_5490,N_5370);
or U6315 (N_6315,N_5869,N_5917);
and U6316 (N_6316,N_5396,N_5808);
and U6317 (N_6317,N_5791,N_5752);
nor U6318 (N_6318,N_5556,N_5853);
xor U6319 (N_6319,N_5983,N_5303);
or U6320 (N_6320,N_5620,N_5583);
or U6321 (N_6321,N_5785,N_5901);
nor U6322 (N_6322,N_5316,N_5402);
nand U6323 (N_6323,N_5721,N_5740);
nand U6324 (N_6324,N_5484,N_5723);
nor U6325 (N_6325,N_5814,N_5427);
xnor U6326 (N_6326,N_5940,N_5968);
and U6327 (N_6327,N_5503,N_5944);
or U6328 (N_6328,N_5941,N_5379);
nor U6329 (N_6329,N_5442,N_5744);
nor U6330 (N_6330,N_5875,N_5616);
or U6331 (N_6331,N_5380,N_5455);
and U6332 (N_6332,N_5974,N_5346);
and U6333 (N_6333,N_5910,N_5893);
and U6334 (N_6334,N_5450,N_5454);
nor U6335 (N_6335,N_5806,N_5517);
xor U6336 (N_6336,N_5384,N_5858);
xor U6337 (N_6337,N_5477,N_5787);
nor U6338 (N_6338,N_5409,N_5631);
xor U6339 (N_6339,N_5317,N_5349);
nor U6340 (N_6340,N_5595,N_5967);
nand U6341 (N_6341,N_5564,N_5880);
or U6342 (N_6342,N_5639,N_5271);
nor U6343 (N_6343,N_5555,N_5507);
or U6344 (N_6344,N_5690,N_5270);
xor U6345 (N_6345,N_5509,N_5320);
nand U6346 (N_6346,N_5698,N_5727);
and U6347 (N_6347,N_5329,N_5365);
xor U6348 (N_6348,N_5866,N_5859);
or U6349 (N_6349,N_5504,N_5335);
nor U6350 (N_6350,N_5845,N_5322);
xor U6351 (N_6351,N_5348,N_5618);
nand U6352 (N_6352,N_5816,N_5494);
or U6353 (N_6353,N_5810,N_5540);
xor U6354 (N_6354,N_5658,N_5513);
nand U6355 (N_6355,N_5543,N_5385);
nor U6356 (N_6356,N_5398,N_5255);
xnor U6357 (N_6357,N_5825,N_5953);
nor U6358 (N_6358,N_5894,N_5475);
or U6359 (N_6359,N_5662,N_5469);
and U6360 (N_6360,N_5802,N_5437);
nand U6361 (N_6361,N_5960,N_5615);
or U6362 (N_6362,N_5497,N_5687);
nor U6363 (N_6363,N_5448,N_5971);
nand U6364 (N_6364,N_5488,N_5778);
or U6365 (N_6365,N_5789,N_5263);
and U6366 (N_6366,N_5948,N_5767);
and U6367 (N_6367,N_5738,N_5676);
or U6368 (N_6368,N_5578,N_5281);
xor U6369 (N_6369,N_5305,N_5704);
and U6370 (N_6370,N_5672,N_5571);
or U6371 (N_6371,N_5678,N_5552);
nand U6372 (N_6372,N_5881,N_5699);
xnor U6373 (N_6373,N_5275,N_5961);
or U6374 (N_6374,N_5684,N_5887);
or U6375 (N_6375,N_5830,N_5358);
and U6376 (N_6376,N_5260,N_5483);
nor U6377 (N_6377,N_5474,N_5972);
nand U6378 (N_6378,N_5615,N_5604);
nand U6379 (N_6379,N_5532,N_5821);
and U6380 (N_6380,N_5912,N_5638);
and U6381 (N_6381,N_5330,N_5361);
or U6382 (N_6382,N_5889,N_5746);
nor U6383 (N_6383,N_5578,N_5841);
or U6384 (N_6384,N_5649,N_5647);
xor U6385 (N_6385,N_5392,N_5769);
nand U6386 (N_6386,N_5808,N_5335);
and U6387 (N_6387,N_5801,N_5282);
xor U6388 (N_6388,N_5980,N_5267);
xor U6389 (N_6389,N_5911,N_5277);
nand U6390 (N_6390,N_5635,N_5259);
or U6391 (N_6391,N_5746,N_5809);
nand U6392 (N_6392,N_5567,N_5855);
nor U6393 (N_6393,N_5755,N_5762);
or U6394 (N_6394,N_5947,N_5374);
xnor U6395 (N_6395,N_5391,N_5268);
or U6396 (N_6396,N_5928,N_5544);
nor U6397 (N_6397,N_5901,N_5755);
or U6398 (N_6398,N_5251,N_5564);
xor U6399 (N_6399,N_5655,N_5526);
xor U6400 (N_6400,N_5521,N_5309);
xnor U6401 (N_6401,N_5387,N_5886);
or U6402 (N_6402,N_5907,N_5514);
or U6403 (N_6403,N_5860,N_5263);
nand U6404 (N_6404,N_5592,N_5449);
xor U6405 (N_6405,N_5919,N_5620);
xor U6406 (N_6406,N_5701,N_5492);
and U6407 (N_6407,N_5769,N_5836);
or U6408 (N_6408,N_5469,N_5997);
xnor U6409 (N_6409,N_5829,N_5311);
xor U6410 (N_6410,N_5588,N_5344);
nand U6411 (N_6411,N_5636,N_5582);
and U6412 (N_6412,N_5263,N_5480);
or U6413 (N_6413,N_5573,N_5671);
nor U6414 (N_6414,N_5384,N_5665);
or U6415 (N_6415,N_5663,N_5865);
and U6416 (N_6416,N_5851,N_5751);
nor U6417 (N_6417,N_5305,N_5373);
nand U6418 (N_6418,N_5860,N_5507);
and U6419 (N_6419,N_5849,N_5709);
nand U6420 (N_6420,N_5552,N_5342);
and U6421 (N_6421,N_5782,N_5553);
nor U6422 (N_6422,N_5669,N_5567);
xor U6423 (N_6423,N_5788,N_5488);
nand U6424 (N_6424,N_5964,N_5555);
xnor U6425 (N_6425,N_5877,N_5921);
and U6426 (N_6426,N_5903,N_5619);
nand U6427 (N_6427,N_5887,N_5503);
nand U6428 (N_6428,N_5994,N_5636);
and U6429 (N_6429,N_5421,N_5558);
nor U6430 (N_6430,N_5520,N_5760);
nand U6431 (N_6431,N_5252,N_5736);
nor U6432 (N_6432,N_5255,N_5890);
xnor U6433 (N_6433,N_5540,N_5870);
nand U6434 (N_6434,N_5988,N_5647);
xor U6435 (N_6435,N_5421,N_5805);
xor U6436 (N_6436,N_5774,N_5839);
nor U6437 (N_6437,N_5356,N_5601);
xor U6438 (N_6438,N_5827,N_5370);
nand U6439 (N_6439,N_5987,N_5944);
nand U6440 (N_6440,N_5825,N_5366);
nor U6441 (N_6441,N_5747,N_5608);
nor U6442 (N_6442,N_5314,N_5859);
xor U6443 (N_6443,N_5709,N_5854);
nand U6444 (N_6444,N_5731,N_5610);
xnor U6445 (N_6445,N_5524,N_5657);
nand U6446 (N_6446,N_5637,N_5570);
nand U6447 (N_6447,N_5881,N_5884);
xnor U6448 (N_6448,N_5630,N_5938);
xor U6449 (N_6449,N_5332,N_5558);
and U6450 (N_6450,N_5912,N_5731);
or U6451 (N_6451,N_5953,N_5354);
nand U6452 (N_6452,N_5799,N_5721);
and U6453 (N_6453,N_5464,N_5800);
nor U6454 (N_6454,N_5702,N_5723);
nand U6455 (N_6455,N_5769,N_5390);
or U6456 (N_6456,N_5481,N_5401);
and U6457 (N_6457,N_5484,N_5681);
nor U6458 (N_6458,N_5422,N_5732);
nand U6459 (N_6459,N_5825,N_5971);
nand U6460 (N_6460,N_5602,N_5813);
or U6461 (N_6461,N_5539,N_5707);
and U6462 (N_6462,N_5545,N_5564);
nor U6463 (N_6463,N_5458,N_5401);
xnor U6464 (N_6464,N_5415,N_5922);
xor U6465 (N_6465,N_5899,N_5504);
and U6466 (N_6466,N_5850,N_5525);
xnor U6467 (N_6467,N_5896,N_5489);
nor U6468 (N_6468,N_5277,N_5614);
nor U6469 (N_6469,N_5642,N_5778);
and U6470 (N_6470,N_5539,N_5949);
xnor U6471 (N_6471,N_5518,N_5865);
or U6472 (N_6472,N_5991,N_5737);
and U6473 (N_6473,N_5412,N_5929);
xor U6474 (N_6474,N_5261,N_5831);
xor U6475 (N_6475,N_5520,N_5854);
nand U6476 (N_6476,N_5946,N_5285);
and U6477 (N_6477,N_5839,N_5775);
or U6478 (N_6478,N_5312,N_5844);
nor U6479 (N_6479,N_5706,N_5920);
and U6480 (N_6480,N_5842,N_5413);
xnor U6481 (N_6481,N_5684,N_5865);
or U6482 (N_6482,N_5648,N_5658);
nor U6483 (N_6483,N_5338,N_5304);
nor U6484 (N_6484,N_5551,N_5692);
and U6485 (N_6485,N_5616,N_5424);
or U6486 (N_6486,N_5511,N_5602);
nor U6487 (N_6487,N_5715,N_5286);
and U6488 (N_6488,N_5829,N_5287);
and U6489 (N_6489,N_5986,N_5648);
xnor U6490 (N_6490,N_5943,N_5945);
nor U6491 (N_6491,N_5541,N_5999);
nand U6492 (N_6492,N_5749,N_5812);
nand U6493 (N_6493,N_5918,N_5373);
and U6494 (N_6494,N_5856,N_5775);
or U6495 (N_6495,N_5405,N_5973);
and U6496 (N_6496,N_5484,N_5845);
xor U6497 (N_6497,N_5678,N_5474);
nand U6498 (N_6498,N_5602,N_5336);
and U6499 (N_6499,N_5557,N_5289);
nor U6500 (N_6500,N_5253,N_5824);
xor U6501 (N_6501,N_5825,N_5292);
xnor U6502 (N_6502,N_5315,N_5545);
xor U6503 (N_6503,N_5460,N_5764);
nand U6504 (N_6504,N_5784,N_5908);
and U6505 (N_6505,N_5401,N_5689);
and U6506 (N_6506,N_5738,N_5955);
and U6507 (N_6507,N_5701,N_5260);
and U6508 (N_6508,N_5427,N_5623);
nand U6509 (N_6509,N_5263,N_5433);
nor U6510 (N_6510,N_5308,N_5311);
nor U6511 (N_6511,N_5285,N_5254);
xor U6512 (N_6512,N_5606,N_5932);
xor U6513 (N_6513,N_5973,N_5557);
nor U6514 (N_6514,N_5477,N_5612);
xor U6515 (N_6515,N_5406,N_5906);
nor U6516 (N_6516,N_5478,N_5933);
nand U6517 (N_6517,N_5532,N_5665);
and U6518 (N_6518,N_5322,N_5650);
or U6519 (N_6519,N_5554,N_5296);
nor U6520 (N_6520,N_5576,N_5301);
or U6521 (N_6521,N_5669,N_5900);
nor U6522 (N_6522,N_5510,N_5871);
and U6523 (N_6523,N_5553,N_5777);
nand U6524 (N_6524,N_5594,N_5874);
or U6525 (N_6525,N_5320,N_5944);
nand U6526 (N_6526,N_5324,N_5640);
and U6527 (N_6527,N_5749,N_5654);
and U6528 (N_6528,N_5309,N_5380);
and U6529 (N_6529,N_5328,N_5310);
nand U6530 (N_6530,N_5602,N_5355);
xor U6531 (N_6531,N_5852,N_5463);
nand U6532 (N_6532,N_5946,N_5279);
nor U6533 (N_6533,N_5682,N_5886);
nor U6534 (N_6534,N_5506,N_5944);
xor U6535 (N_6535,N_5345,N_5504);
nand U6536 (N_6536,N_5895,N_5649);
nor U6537 (N_6537,N_5675,N_5667);
nor U6538 (N_6538,N_5664,N_5614);
xor U6539 (N_6539,N_5499,N_5867);
and U6540 (N_6540,N_5395,N_5912);
and U6541 (N_6541,N_5410,N_5905);
or U6542 (N_6542,N_5620,N_5505);
xor U6543 (N_6543,N_5960,N_5563);
nand U6544 (N_6544,N_5664,N_5702);
nand U6545 (N_6545,N_5546,N_5921);
or U6546 (N_6546,N_5661,N_5649);
nor U6547 (N_6547,N_5827,N_5259);
nor U6548 (N_6548,N_5758,N_5931);
or U6549 (N_6549,N_5542,N_5413);
xor U6550 (N_6550,N_5704,N_5416);
or U6551 (N_6551,N_5730,N_5854);
nor U6552 (N_6552,N_5897,N_5532);
xor U6553 (N_6553,N_5597,N_5316);
or U6554 (N_6554,N_5705,N_5587);
xor U6555 (N_6555,N_5750,N_5579);
and U6556 (N_6556,N_5405,N_5492);
xor U6557 (N_6557,N_5657,N_5910);
or U6558 (N_6558,N_5716,N_5347);
xnor U6559 (N_6559,N_5979,N_5746);
xnor U6560 (N_6560,N_5700,N_5297);
or U6561 (N_6561,N_5689,N_5590);
nor U6562 (N_6562,N_5314,N_5329);
nand U6563 (N_6563,N_5694,N_5466);
nor U6564 (N_6564,N_5304,N_5356);
or U6565 (N_6565,N_5769,N_5465);
nor U6566 (N_6566,N_5926,N_5699);
or U6567 (N_6567,N_5880,N_5408);
xor U6568 (N_6568,N_5861,N_5383);
nor U6569 (N_6569,N_5794,N_5545);
or U6570 (N_6570,N_5889,N_5658);
nor U6571 (N_6571,N_5901,N_5560);
or U6572 (N_6572,N_5533,N_5987);
nor U6573 (N_6573,N_5530,N_5310);
and U6574 (N_6574,N_5924,N_5283);
nand U6575 (N_6575,N_5363,N_5251);
or U6576 (N_6576,N_5795,N_5318);
and U6577 (N_6577,N_5282,N_5633);
xnor U6578 (N_6578,N_5756,N_5621);
nand U6579 (N_6579,N_5774,N_5979);
and U6580 (N_6580,N_5567,N_5560);
and U6581 (N_6581,N_5726,N_5524);
xnor U6582 (N_6582,N_5928,N_5664);
and U6583 (N_6583,N_5572,N_5704);
or U6584 (N_6584,N_5899,N_5524);
xor U6585 (N_6585,N_5422,N_5807);
nand U6586 (N_6586,N_5824,N_5810);
nor U6587 (N_6587,N_5716,N_5790);
nor U6588 (N_6588,N_5940,N_5782);
and U6589 (N_6589,N_5781,N_5367);
nor U6590 (N_6590,N_5366,N_5377);
xor U6591 (N_6591,N_5422,N_5453);
nand U6592 (N_6592,N_5699,N_5995);
nor U6593 (N_6593,N_5863,N_5605);
nor U6594 (N_6594,N_5322,N_5378);
nor U6595 (N_6595,N_5557,N_5567);
nand U6596 (N_6596,N_5499,N_5441);
or U6597 (N_6597,N_5629,N_5399);
or U6598 (N_6598,N_5960,N_5298);
nor U6599 (N_6599,N_5348,N_5519);
nand U6600 (N_6600,N_5256,N_5305);
and U6601 (N_6601,N_5942,N_5860);
and U6602 (N_6602,N_5901,N_5275);
nand U6603 (N_6603,N_5824,N_5311);
and U6604 (N_6604,N_5850,N_5402);
or U6605 (N_6605,N_5927,N_5630);
or U6606 (N_6606,N_5944,N_5272);
and U6607 (N_6607,N_5387,N_5682);
and U6608 (N_6608,N_5931,N_5797);
or U6609 (N_6609,N_5805,N_5425);
and U6610 (N_6610,N_5728,N_5855);
nor U6611 (N_6611,N_5334,N_5894);
nand U6612 (N_6612,N_5370,N_5843);
nand U6613 (N_6613,N_5605,N_5977);
xor U6614 (N_6614,N_5476,N_5649);
xor U6615 (N_6615,N_5301,N_5700);
xor U6616 (N_6616,N_5576,N_5715);
nor U6617 (N_6617,N_5414,N_5472);
nand U6618 (N_6618,N_5364,N_5783);
nand U6619 (N_6619,N_5312,N_5602);
or U6620 (N_6620,N_5982,N_5701);
and U6621 (N_6621,N_5819,N_5815);
nand U6622 (N_6622,N_5845,N_5946);
and U6623 (N_6623,N_5735,N_5522);
nand U6624 (N_6624,N_5465,N_5921);
and U6625 (N_6625,N_5714,N_5542);
and U6626 (N_6626,N_5513,N_5376);
nand U6627 (N_6627,N_5685,N_5324);
or U6628 (N_6628,N_5766,N_5668);
or U6629 (N_6629,N_5737,N_5488);
or U6630 (N_6630,N_5679,N_5576);
nand U6631 (N_6631,N_5983,N_5835);
nor U6632 (N_6632,N_5669,N_5868);
nand U6633 (N_6633,N_5346,N_5640);
nand U6634 (N_6634,N_5871,N_5990);
and U6635 (N_6635,N_5810,N_5500);
or U6636 (N_6636,N_5880,N_5270);
xor U6637 (N_6637,N_5344,N_5538);
nand U6638 (N_6638,N_5984,N_5964);
and U6639 (N_6639,N_5709,N_5787);
and U6640 (N_6640,N_5337,N_5592);
xnor U6641 (N_6641,N_5325,N_5745);
and U6642 (N_6642,N_5661,N_5656);
or U6643 (N_6643,N_5362,N_5576);
and U6644 (N_6644,N_5974,N_5698);
and U6645 (N_6645,N_5583,N_5830);
xnor U6646 (N_6646,N_5449,N_5364);
nand U6647 (N_6647,N_5322,N_5554);
or U6648 (N_6648,N_5344,N_5722);
or U6649 (N_6649,N_5908,N_5565);
xnor U6650 (N_6650,N_5549,N_5985);
xnor U6651 (N_6651,N_5480,N_5699);
nor U6652 (N_6652,N_5622,N_5536);
nor U6653 (N_6653,N_5544,N_5504);
xor U6654 (N_6654,N_5388,N_5524);
nor U6655 (N_6655,N_5922,N_5417);
and U6656 (N_6656,N_5481,N_5398);
xor U6657 (N_6657,N_5338,N_5377);
xnor U6658 (N_6658,N_5891,N_5739);
nor U6659 (N_6659,N_5912,N_5405);
nor U6660 (N_6660,N_5702,N_5886);
nand U6661 (N_6661,N_5253,N_5737);
nor U6662 (N_6662,N_5762,N_5880);
nand U6663 (N_6663,N_5538,N_5952);
and U6664 (N_6664,N_5607,N_5355);
nand U6665 (N_6665,N_5576,N_5677);
nor U6666 (N_6666,N_5887,N_5625);
nand U6667 (N_6667,N_5642,N_5494);
and U6668 (N_6668,N_5444,N_5857);
nand U6669 (N_6669,N_5260,N_5740);
xnor U6670 (N_6670,N_5325,N_5879);
nand U6671 (N_6671,N_5863,N_5961);
nand U6672 (N_6672,N_5807,N_5613);
or U6673 (N_6673,N_5844,N_5492);
or U6674 (N_6674,N_5517,N_5412);
nand U6675 (N_6675,N_5547,N_5686);
xnor U6676 (N_6676,N_5936,N_5655);
and U6677 (N_6677,N_5927,N_5890);
xor U6678 (N_6678,N_5320,N_5758);
and U6679 (N_6679,N_5618,N_5265);
xnor U6680 (N_6680,N_5279,N_5370);
or U6681 (N_6681,N_5920,N_5871);
or U6682 (N_6682,N_5506,N_5791);
xor U6683 (N_6683,N_5308,N_5965);
nand U6684 (N_6684,N_5354,N_5739);
xnor U6685 (N_6685,N_5887,N_5616);
nor U6686 (N_6686,N_5255,N_5674);
and U6687 (N_6687,N_5505,N_5358);
xnor U6688 (N_6688,N_5807,N_5510);
or U6689 (N_6689,N_5749,N_5370);
or U6690 (N_6690,N_5597,N_5886);
and U6691 (N_6691,N_5685,N_5396);
or U6692 (N_6692,N_5654,N_5526);
or U6693 (N_6693,N_5942,N_5599);
xor U6694 (N_6694,N_5663,N_5840);
or U6695 (N_6695,N_5692,N_5286);
nor U6696 (N_6696,N_5418,N_5623);
xnor U6697 (N_6697,N_5634,N_5691);
or U6698 (N_6698,N_5461,N_5767);
nand U6699 (N_6699,N_5326,N_5652);
and U6700 (N_6700,N_5488,N_5557);
xor U6701 (N_6701,N_5746,N_5996);
xor U6702 (N_6702,N_5801,N_5502);
xor U6703 (N_6703,N_5914,N_5849);
xor U6704 (N_6704,N_5282,N_5446);
nor U6705 (N_6705,N_5886,N_5911);
xnor U6706 (N_6706,N_5449,N_5403);
and U6707 (N_6707,N_5880,N_5658);
or U6708 (N_6708,N_5839,N_5413);
nand U6709 (N_6709,N_5783,N_5652);
nand U6710 (N_6710,N_5937,N_5883);
nand U6711 (N_6711,N_5320,N_5542);
nand U6712 (N_6712,N_5961,N_5447);
nor U6713 (N_6713,N_5688,N_5358);
nor U6714 (N_6714,N_5717,N_5656);
nand U6715 (N_6715,N_5491,N_5565);
and U6716 (N_6716,N_5989,N_5559);
or U6717 (N_6717,N_5651,N_5500);
nor U6718 (N_6718,N_5700,N_5726);
xor U6719 (N_6719,N_5562,N_5310);
and U6720 (N_6720,N_5369,N_5739);
nand U6721 (N_6721,N_5599,N_5613);
or U6722 (N_6722,N_5525,N_5292);
and U6723 (N_6723,N_5940,N_5801);
and U6724 (N_6724,N_5999,N_5354);
nand U6725 (N_6725,N_5988,N_5392);
xor U6726 (N_6726,N_5418,N_5942);
and U6727 (N_6727,N_5514,N_5799);
or U6728 (N_6728,N_5687,N_5918);
and U6729 (N_6729,N_5344,N_5584);
or U6730 (N_6730,N_5382,N_5443);
nand U6731 (N_6731,N_5450,N_5483);
and U6732 (N_6732,N_5467,N_5983);
or U6733 (N_6733,N_5380,N_5654);
nor U6734 (N_6734,N_5326,N_5553);
xnor U6735 (N_6735,N_5903,N_5776);
xor U6736 (N_6736,N_5465,N_5314);
nor U6737 (N_6737,N_5686,N_5485);
nand U6738 (N_6738,N_5475,N_5533);
and U6739 (N_6739,N_5707,N_5709);
and U6740 (N_6740,N_5608,N_5750);
and U6741 (N_6741,N_5963,N_5285);
xnor U6742 (N_6742,N_5770,N_5899);
and U6743 (N_6743,N_5565,N_5396);
and U6744 (N_6744,N_5636,N_5991);
or U6745 (N_6745,N_5415,N_5779);
nand U6746 (N_6746,N_5561,N_5515);
and U6747 (N_6747,N_5338,N_5535);
and U6748 (N_6748,N_5272,N_5744);
and U6749 (N_6749,N_5350,N_5634);
nand U6750 (N_6750,N_6399,N_6257);
nor U6751 (N_6751,N_6183,N_6255);
or U6752 (N_6752,N_6552,N_6386);
xor U6753 (N_6753,N_6131,N_6001);
nand U6754 (N_6754,N_6007,N_6330);
nand U6755 (N_6755,N_6317,N_6042);
xor U6756 (N_6756,N_6199,N_6073);
nor U6757 (N_6757,N_6032,N_6563);
or U6758 (N_6758,N_6024,N_6151);
nand U6759 (N_6759,N_6018,N_6260);
xnor U6760 (N_6760,N_6282,N_6542);
xor U6761 (N_6761,N_6556,N_6631);
and U6762 (N_6762,N_6075,N_6414);
or U6763 (N_6763,N_6017,N_6342);
and U6764 (N_6764,N_6059,N_6186);
and U6765 (N_6765,N_6663,N_6671);
and U6766 (N_6766,N_6160,N_6510);
and U6767 (N_6767,N_6606,N_6412);
or U6768 (N_6768,N_6102,N_6016);
nor U6769 (N_6769,N_6006,N_6576);
nand U6770 (N_6770,N_6082,N_6624);
xor U6771 (N_6771,N_6424,N_6713);
nand U6772 (N_6772,N_6425,N_6190);
xnor U6773 (N_6773,N_6246,N_6258);
and U6774 (N_6774,N_6309,N_6578);
nand U6775 (N_6775,N_6251,N_6459);
nor U6776 (N_6776,N_6277,N_6435);
or U6777 (N_6777,N_6140,N_6261);
or U6778 (N_6778,N_6478,N_6376);
and U6779 (N_6779,N_6534,N_6544);
nand U6780 (N_6780,N_6736,N_6543);
nand U6781 (N_6781,N_6422,N_6152);
and U6782 (N_6782,N_6270,N_6148);
xnor U6783 (N_6783,N_6276,N_6492);
nand U6784 (N_6784,N_6746,N_6494);
xor U6785 (N_6785,N_6182,N_6648);
and U6786 (N_6786,N_6033,N_6395);
xnor U6787 (N_6787,N_6592,N_6045);
xor U6788 (N_6788,N_6333,N_6515);
nand U6789 (N_6789,N_6288,N_6083);
xnor U6790 (N_6790,N_6575,N_6044);
nor U6791 (N_6791,N_6585,N_6672);
and U6792 (N_6792,N_6105,N_6472);
nand U6793 (N_6793,N_6539,N_6476);
and U6794 (N_6794,N_6571,N_6323);
nand U6795 (N_6795,N_6615,N_6526);
nor U6796 (N_6796,N_6292,N_6189);
nand U6797 (N_6797,N_6030,N_6621);
xor U6798 (N_6798,N_6020,N_6013);
or U6799 (N_6799,N_6058,N_6240);
and U6800 (N_6800,N_6065,N_6532);
nand U6801 (N_6801,N_6324,N_6206);
and U6802 (N_6802,N_6410,N_6647);
nand U6803 (N_6803,N_6328,N_6245);
nand U6804 (N_6804,N_6745,N_6369);
xor U6805 (N_6805,N_6721,N_6703);
xnor U6806 (N_6806,N_6594,N_6620);
and U6807 (N_6807,N_6726,N_6359);
xor U6808 (N_6808,N_6164,N_6372);
nand U6809 (N_6809,N_6008,N_6715);
xnor U6810 (N_6810,N_6043,N_6431);
xnor U6811 (N_6811,N_6389,N_6450);
and U6812 (N_6812,N_6128,N_6373);
or U6813 (N_6813,N_6747,N_6439);
nand U6814 (N_6814,N_6092,N_6391);
nand U6815 (N_6815,N_6191,N_6172);
xnor U6816 (N_6816,N_6656,N_6582);
xor U6817 (N_6817,N_6619,N_6505);
and U6818 (N_6818,N_6235,N_6290);
and U6819 (N_6819,N_6451,N_6602);
xnor U6820 (N_6820,N_6162,N_6285);
and U6821 (N_6821,N_6327,N_6400);
xnor U6822 (N_6822,N_6433,N_6081);
nor U6823 (N_6823,N_6562,N_6355);
xnor U6824 (N_6824,N_6237,N_6627);
nor U6825 (N_6825,N_6192,N_6470);
xor U6826 (N_6826,N_6286,N_6012);
and U6827 (N_6827,N_6229,N_6232);
xnor U6828 (N_6828,N_6074,N_6497);
nand U6829 (N_6829,N_6717,N_6474);
and U6830 (N_6830,N_6460,N_6679);
nor U6831 (N_6831,N_6638,N_6112);
or U6832 (N_6832,N_6301,N_6654);
xor U6833 (N_6833,N_6611,N_6367);
or U6834 (N_6834,N_6274,N_6479);
nor U6835 (N_6835,N_6567,N_6210);
or U6836 (N_6836,N_6166,N_6674);
or U6837 (N_6837,N_6499,N_6040);
nor U6838 (N_6838,N_6196,N_6436);
nor U6839 (N_6839,N_6377,N_6614);
xor U6840 (N_6840,N_6749,N_6710);
nor U6841 (N_6841,N_6720,N_6050);
nand U6842 (N_6842,N_6402,N_6593);
nor U6843 (N_6843,N_6605,N_6429);
and U6844 (N_6844,N_6089,N_6573);
nand U6845 (N_6845,N_6444,N_6486);
and U6846 (N_6846,N_6052,N_6417);
nand U6847 (N_6847,N_6533,N_6256);
and U6848 (N_6848,N_6354,N_6714);
nand U6849 (N_6849,N_6347,N_6063);
xor U6850 (N_6850,N_6003,N_6150);
nor U6851 (N_6851,N_6336,N_6156);
or U6852 (N_6852,N_6019,N_6313);
xor U6853 (N_6853,N_6490,N_6649);
and U6854 (N_6854,N_6031,N_6618);
or U6855 (N_6855,N_6712,N_6241);
nand U6856 (N_6856,N_6467,N_6180);
or U6857 (N_6857,N_6111,N_6218);
or U6858 (N_6858,N_6316,N_6302);
and U6859 (N_6859,N_6034,N_6334);
or U6860 (N_6860,N_6743,N_6310);
nor U6861 (N_6861,N_6087,N_6315);
xor U6862 (N_6862,N_6384,N_6697);
nor U6863 (N_6863,N_6167,N_6742);
nand U6864 (N_6864,N_6363,N_6155);
nor U6865 (N_6865,N_6652,N_6070);
xnor U6866 (N_6866,N_6265,N_6493);
nor U6867 (N_6867,N_6056,N_6587);
or U6868 (N_6868,N_6072,N_6094);
nand U6869 (N_6869,N_6568,N_6064);
or U6870 (N_6870,N_6360,N_6341);
and U6871 (N_6871,N_6047,N_6343);
xor U6872 (N_6872,N_6053,N_6512);
and U6873 (N_6873,N_6076,N_6465);
or U6874 (N_6874,N_6250,N_6491);
and U6875 (N_6875,N_6642,N_6570);
xnor U6876 (N_6876,N_6254,N_6035);
nand U6877 (N_6877,N_6550,N_6427);
or U6878 (N_6878,N_6187,N_6731);
and U6879 (N_6879,N_6695,N_6121);
nor U6880 (N_6880,N_6730,N_6722);
xor U6881 (N_6881,N_6516,N_6116);
and U6882 (N_6882,N_6421,N_6095);
nand U6883 (N_6883,N_6634,N_6509);
nor U6884 (N_6884,N_6234,N_6666);
or U6885 (N_6885,N_6120,N_6272);
or U6886 (N_6886,N_6049,N_6464);
nand U6887 (N_6887,N_6704,N_6590);
and U6888 (N_6888,N_6549,N_6134);
nand U6889 (N_6889,N_6737,N_6716);
xnor U6890 (N_6890,N_6597,N_6688);
nand U6891 (N_6891,N_6370,N_6572);
nand U6892 (N_6892,N_6247,N_6209);
nor U6893 (N_6893,N_6548,N_6078);
nand U6894 (N_6894,N_6280,N_6732);
and U6895 (N_6895,N_6705,N_6362);
nor U6896 (N_6896,N_6036,N_6657);
xnor U6897 (N_6897,N_6293,N_6104);
xor U6898 (N_6898,N_6356,N_6238);
and U6899 (N_6899,N_6170,N_6506);
xor U6900 (N_6900,N_6419,N_6067);
nand U6901 (N_6901,N_6588,N_6253);
nor U6902 (N_6902,N_6616,N_6368);
and U6903 (N_6903,N_6346,N_6482);
nand U6904 (N_6904,N_6338,N_6441);
nand U6905 (N_6905,N_6311,N_6096);
or U6906 (N_6906,N_6744,N_6066);
nand U6907 (N_6907,N_6584,N_6623);
or U6908 (N_6908,N_6469,N_6735);
and U6909 (N_6909,N_6650,N_6084);
or U6910 (N_6910,N_6527,N_6204);
nor U6911 (N_6911,N_6653,N_6138);
or U6912 (N_6912,N_6269,N_6103);
nor U6913 (N_6913,N_6561,N_6268);
or U6914 (N_6914,N_6109,N_6503);
nand U6915 (N_6915,N_6243,N_6188);
nor U6916 (N_6916,N_6039,N_6521);
and U6917 (N_6917,N_6348,N_6706);
and U6918 (N_6918,N_6297,N_6291);
xnor U6919 (N_6919,N_6669,N_6118);
xnor U6920 (N_6920,N_6130,N_6723);
nor U6921 (N_6921,N_6227,N_6122);
and U6922 (N_6922,N_6353,N_6644);
nor U6923 (N_6923,N_6021,N_6530);
nor U6924 (N_6924,N_6380,N_6404);
nor U6925 (N_6925,N_6004,N_6212);
nor U6926 (N_6926,N_6147,N_6379);
xor U6927 (N_6927,N_6179,N_6077);
and U6928 (N_6928,N_6434,N_6242);
and U6929 (N_6929,N_6686,N_6358);
or U6930 (N_6930,N_6289,N_6536);
and U6931 (N_6931,N_6197,N_6423);
nor U6932 (N_6932,N_6633,N_6683);
or U6933 (N_6933,N_6696,N_6603);
and U6934 (N_6934,N_6655,N_6388);
or U6935 (N_6935,N_6393,N_6524);
xnor U6936 (N_6936,N_6387,N_6739);
nand U6937 (N_6937,N_6418,N_6217);
nand U6938 (N_6938,N_6296,N_6681);
nor U6939 (N_6939,N_6060,N_6629);
nor U6940 (N_6940,N_6127,N_6287);
nand U6941 (N_6941,N_6248,N_6511);
or U6942 (N_6942,N_6124,N_6284);
or U6943 (N_6943,N_6264,N_6734);
and U6944 (N_6944,N_6177,N_6661);
or U6945 (N_6945,N_6225,N_6143);
and U6946 (N_6946,N_6537,N_6061);
xnor U6947 (N_6947,N_6529,N_6086);
and U6948 (N_6948,N_6098,N_6591);
and U6949 (N_6949,N_6660,N_6080);
nor U6950 (N_6950,N_6553,N_6741);
and U6951 (N_6951,N_6322,N_6205);
and U6952 (N_6952,N_6097,N_6538);
xor U6953 (N_6953,N_6673,N_6230);
nand U6954 (N_6954,N_6306,N_6129);
xnor U6955 (N_6955,N_6701,N_6279);
xnor U6956 (N_6956,N_6038,N_6107);
or U6957 (N_6957,N_6161,N_6055);
and U6958 (N_6958,N_6228,N_6202);
or U6959 (N_6959,N_6498,N_6068);
and U6960 (N_6960,N_6637,N_6557);
or U6961 (N_6961,N_6294,N_6522);
xnor U6962 (N_6962,N_6687,N_6407);
or U6963 (N_6963,N_6325,N_6119);
and U6964 (N_6964,N_6171,N_6565);
or U6965 (N_6965,N_6437,N_6223);
or U6966 (N_6966,N_6484,N_6636);
xor U6967 (N_6967,N_6321,N_6026);
or U6968 (N_6968,N_6513,N_6520);
and U6969 (N_6969,N_6331,N_6233);
nor U6970 (N_6970,N_6579,N_6022);
nand U6971 (N_6971,N_6707,N_6612);
xor U6972 (N_6972,N_6574,N_6165);
and U6973 (N_6973,N_6169,N_6304);
nor U6974 (N_6974,N_6485,N_6011);
xnor U6975 (N_6975,N_6483,N_6403);
nor U6976 (N_6976,N_6298,N_6193);
and U6977 (N_6977,N_6662,N_6528);
or U6978 (N_6978,N_6569,N_6443);
and U6979 (N_6979,N_6224,N_6184);
nand U6980 (N_6980,N_6014,N_6617);
xor U6981 (N_6981,N_6699,N_6468);
or U6982 (N_6982,N_6028,N_6259);
nand U6983 (N_6983,N_6420,N_6106);
and U6984 (N_6984,N_6231,N_6303);
xnor U6985 (N_6985,N_6453,N_6025);
nor U6986 (N_6986,N_6378,N_6397);
nand U6987 (N_6987,N_6555,N_6609);
nand U6988 (N_6988,N_6554,N_6300);
or U6989 (N_6989,N_6689,N_6738);
xnor U6990 (N_6990,N_6239,N_6314);
xor U6991 (N_6991,N_6023,N_6275);
nor U6992 (N_6992,N_6525,N_6219);
or U6993 (N_6993,N_6589,N_6339);
nor U6994 (N_6994,N_6471,N_6222);
xnor U6995 (N_6995,N_6457,N_6708);
xnor U6996 (N_6996,N_6366,N_6487);
xnor U6997 (N_6997,N_6266,N_6110);
nand U6998 (N_6998,N_6643,N_6062);
xnor U6999 (N_6999,N_6684,N_6508);
or U7000 (N_7000,N_6027,N_6607);
and U7001 (N_7001,N_6691,N_6091);
and U7002 (N_7002,N_6159,N_6142);
or U7003 (N_7003,N_6117,N_6108);
and U7004 (N_7004,N_6394,N_6215);
nor U7005 (N_7005,N_6740,N_6307);
or U7006 (N_7006,N_6599,N_6085);
and U7007 (N_7007,N_6176,N_6583);
and U7008 (N_7008,N_6178,N_6639);
xor U7009 (N_7009,N_6320,N_6630);
nor U7010 (N_7010,N_6145,N_6153);
xor U7011 (N_7011,N_6480,N_6271);
nor U7012 (N_7012,N_6724,N_6440);
or U7013 (N_7013,N_6398,N_6430);
nand U7014 (N_7014,N_6625,N_6519);
or U7015 (N_7015,N_6560,N_6201);
or U7016 (N_7016,N_6473,N_6329);
xor U7017 (N_7017,N_6299,N_6729);
or U7018 (N_7018,N_6318,N_6452);
nor U7019 (N_7019,N_6651,N_6203);
nor U7020 (N_7020,N_6405,N_6670);
nand U7021 (N_7021,N_6481,N_6458);
and U7022 (N_7022,N_6711,N_6694);
nor U7023 (N_7023,N_6319,N_6531);
xnor U7024 (N_7024,N_6048,N_6496);
and U7025 (N_7025,N_6401,N_6613);
or U7026 (N_7026,N_6278,N_6728);
nand U7027 (N_7027,N_6415,N_6438);
and U7028 (N_7028,N_6344,N_6181);
and U7029 (N_7029,N_6502,N_6194);
nor U7030 (N_7030,N_6396,N_6216);
or U7031 (N_7031,N_6665,N_6658);
and U7032 (N_7032,N_6002,N_6682);
nand U7033 (N_7033,N_6685,N_6409);
and U7034 (N_7034,N_6079,N_6680);
nand U7035 (N_7035,N_6364,N_6208);
xnor U7036 (N_7036,N_6340,N_6071);
nand U7037 (N_7037,N_6295,N_6586);
nor U7038 (N_7038,N_6069,N_6518);
and U7039 (N_7039,N_6226,N_6361);
or U7040 (N_7040,N_6454,N_6381);
xor U7041 (N_7041,N_6382,N_6600);
xnor U7042 (N_7042,N_6220,N_6645);
nor U7043 (N_7043,N_6173,N_6113);
and U7044 (N_7044,N_6558,N_6351);
xnor U7045 (N_7045,N_6447,N_6385);
xor U7046 (N_7046,N_6632,N_6137);
nor U7047 (N_7047,N_6676,N_6046);
or U7048 (N_7048,N_6523,N_6664);
nand U7049 (N_7049,N_6088,N_6326);
xnor U7050 (N_7050,N_6628,N_6267);
and U7051 (N_7051,N_6305,N_6535);
nand U7052 (N_7052,N_6365,N_6559);
and U7053 (N_7053,N_6345,N_6604);
or U7054 (N_7054,N_6211,N_6371);
and U7055 (N_7055,N_6236,N_6037);
or U7056 (N_7056,N_6010,N_6174);
nor U7057 (N_7057,N_6154,N_6641);
xnor U7058 (N_7058,N_6659,N_6350);
or U7059 (N_7059,N_6580,N_6335);
nand U7060 (N_7060,N_6308,N_6709);
xor U7061 (N_7061,N_6125,N_6375);
nor U7062 (N_7062,N_6009,N_6207);
nor U7063 (N_7063,N_6114,N_6426);
nor U7064 (N_7064,N_6698,N_6262);
and U7065 (N_7065,N_6352,N_6123);
or U7066 (N_7066,N_6115,N_6136);
and U7067 (N_7067,N_6135,N_6195);
nor U7068 (N_7068,N_6332,N_6337);
nor U7069 (N_7069,N_6626,N_6719);
nor U7070 (N_7070,N_6545,N_6392);
nor U7071 (N_7071,N_6727,N_6132);
xor U7072 (N_7072,N_6540,N_6428);
and U7073 (N_7073,N_6564,N_6501);
and U7074 (N_7074,N_6445,N_6667);
or U7075 (N_7075,N_6514,N_6610);
nand U7076 (N_7076,N_6668,N_6581);
and U7077 (N_7077,N_6463,N_6718);
nor U7078 (N_7078,N_6133,N_6507);
and U7079 (N_7079,N_6495,N_6595);
xnor U7080 (N_7080,N_6432,N_6244);
nor U7081 (N_7081,N_6489,N_6000);
nand U7082 (N_7082,N_6390,N_6475);
xnor U7083 (N_7083,N_6541,N_6601);
xnor U7084 (N_7084,N_6283,N_6677);
nand U7085 (N_7085,N_6690,N_6263);
nor U7086 (N_7086,N_6051,N_6598);
and U7087 (N_7087,N_6101,N_6157);
or U7088 (N_7088,N_6700,N_6163);
and U7089 (N_7089,N_6646,N_6733);
or U7090 (N_7090,N_6139,N_6141);
xor U7091 (N_7091,N_6596,N_6200);
and U7092 (N_7092,N_6213,N_6146);
or U7093 (N_7093,N_6057,N_6408);
xnor U7094 (N_7094,N_6547,N_6273);
xnor U7095 (N_7095,N_6488,N_6281);
nand U7096 (N_7096,N_6640,N_6214);
nor U7097 (N_7097,N_6357,N_6041);
or U7098 (N_7098,N_6455,N_6546);
or U7099 (N_7099,N_6456,N_6413);
or U7100 (N_7100,N_6252,N_6517);
or U7101 (N_7101,N_6374,N_6149);
or U7102 (N_7102,N_6168,N_6312);
or U7103 (N_7103,N_6005,N_6100);
nand U7104 (N_7104,N_6678,N_6349);
nor U7105 (N_7105,N_6477,N_6093);
xor U7106 (N_7106,N_6198,N_6144);
and U7107 (N_7107,N_6462,N_6692);
and U7108 (N_7108,N_6551,N_6702);
nor U7109 (N_7109,N_6577,N_6221);
nor U7110 (N_7110,N_6029,N_6175);
xor U7111 (N_7111,N_6383,N_6126);
nand U7112 (N_7112,N_6504,N_6442);
xnor U7113 (N_7113,N_6675,N_6461);
and U7114 (N_7114,N_6406,N_6448);
nor U7115 (N_7115,N_6449,N_6249);
nor U7116 (N_7116,N_6054,N_6416);
or U7117 (N_7117,N_6446,N_6158);
nor U7118 (N_7118,N_6748,N_6099);
xnor U7119 (N_7119,N_6693,N_6635);
or U7120 (N_7120,N_6500,N_6566);
and U7121 (N_7121,N_6608,N_6015);
xnor U7122 (N_7122,N_6090,N_6466);
xor U7123 (N_7123,N_6622,N_6725);
nand U7124 (N_7124,N_6411,N_6185);
nand U7125 (N_7125,N_6084,N_6565);
or U7126 (N_7126,N_6632,N_6175);
nand U7127 (N_7127,N_6632,N_6431);
and U7128 (N_7128,N_6738,N_6422);
xor U7129 (N_7129,N_6639,N_6217);
nor U7130 (N_7130,N_6530,N_6419);
nand U7131 (N_7131,N_6248,N_6482);
nand U7132 (N_7132,N_6081,N_6129);
and U7133 (N_7133,N_6713,N_6098);
nor U7134 (N_7134,N_6149,N_6253);
and U7135 (N_7135,N_6280,N_6201);
nor U7136 (N_7136,N_6334,N_6563);
and U7137 (N_7137,N_6250,N_6256);
and U7138 (N_7138,N_6126,N_6031);
and U7139 (N_7139,N_6046,N_6334);
or U7140 (N_7140,N_6313,N_6302);
or U7141 (N_7141,N_6332,N_6489);
nand U7142 (N_7142,N_6139,N_6612);
nor U7143 (N_7143,N_6650,N_6581);
nor U7144 (N_7144,N_6338,N_6109);
or U7145 (N_7145,N_6548,N_6070);
nand U7146 (N_7146,N_6429,N_6568);
or U7147 (N_7147,N_6700,N_6353);
and U7148 (N_7148,N_6234,N_6689);
xor U7149 (N_7149,N_6131,N_6355);
and U7150 (N_7150,N_6285,N_6083);
or U7151 (N_7151,N_6356,N_6640);
nand U7152 (N_7152,N_6587,N_6654);
nor U7153 (N_7153,N_6399,N_6647);
and U7154 (N_7154,N_6691,N_6415);
xor U7155 (N_7155,N_6439,N_6561);
xor U7156 (N_7156,N_6142,N_6153);
or U7157 (N_7157,N_6230,N_6431);
or U7158 (N_7158,N_6606,N_6683);
nand U7159 (N_7159,N_6258,N_6537);
nor U7160 (N_7160,N_6748,N_6741);
or U7161 (N_7161,N_6440,N_6304);
xnor U7162 (N_7162,N_6479,N_6458);
nor U7163 (N_7163,N_6250,N_6009);
nor U7164 (N_7164,N_6146,N_6616);
xor U7165 (N_7165,N_6124,N_6312);
and U7166 (N_7166,N_6274,N_6259);
xnor U7167 (N_7167,N_6129,N_6605);
nand U7168 (N_7168,N_6685,N_6369);
xnor U7169 (N_7169,N_6244,N_6095);
nor U7170 (N_7170,N_6697,N_6310);
and U7171 (N_7171,N_6424,N_6541);
nand U7172 (N_7172,N_6345,N_6254);
nor U7173 (N_7173,N_6176,N_6489);
nor U7174 (N_7174,N_6390,N_6079);
nand U7175 (N_7175,N_6029,N_6394);
or U7176 (N_7176,N_6680,N_6646);
nor U7177 (N_7177,N_6499,N_6377);
or U7178 (N_7178,N_6600,N_6173);
xnor U7179 (N_7179,N_6489,N_6369);
xnor U7180 (N_7180,N_6124,N_6678);
nor U7181 (N_7181,N_6411,N_6676);
and U7182 (N_7182,N_6180,N_6017);
nand U7183 (N_7183,N_6108,N_6458);
xor U7184 (N_7184,N_6260,N_6600);
and U7185 (N_7185,N_6306,N_6034);
and U7186 (N_7186,N_6127,N_6467);
xor U7187 (N_7187,N_6717,N_6473);
or U7188 (N_7188,N_6037,N_6596);
nand U7189 (N_7189,N_6545,N_6133);
xor U7190 (N_7190,N_6396,N_6279);
nor U7191 (N_7191,N_6535,N_6068);
nor U7192 (N_7192,N_6549,N_6234);
xnor U7193 (N_7193,N_6008,N_6619);
xnor U7194 (N_7194,N_6705,N_6119);
nand U7195 (N_7195,N_6518,N_6178);
nor U7196 (N_7196,N_6151,N_6726);
xor U7197 (N_7197,N_6354,N_6027);
nand U7198 (N_7198,N_6052,N_6704);
nand U7199 (N_7199,N_6119,N_6027);
nor U7200 (N_7200,N_6602,N_6408);
or U7201 (N_7201,N_6023,N_6472);
and U7202 (N_7202,N_6094,N_6279);
nor U7203 (N_7203,N_6203,N_6247);
xnor U7204 (N_7204,N_6697,N_6417);
xnor U7205 (N_7205,N_6708,N_6505);
nor U7206 (N_7206,N_6369,N_6283);
nor U7207 (N_7207,N_6611,N_6453);
and U7208 (N_7208,N_6492,N_6358);
nand U7209 (N_7209,N_6154,N_6106);
or U7210 (N_7210,N_6230,N_6607);
nor U7211 (N_7211,N_6108,N_6611);
nor U7212 (N_7212,N_6724,N_6431);
and U7213 (N_7213,N_6605,N_6688);
and U7214 (N_7214,N_6495,N_6519);
nor U7215 (N_7215,N_6075,N_6605);
nor U7216 (N_7216,N_6558,N_6644);
nor U7217 (N_7217,N_6237,N_6015);
and U7218 (N_7218,N_6081,N_6365);
nor U7219 (N_7219,N_6360,N_6187);
or U7220 (N_7220,N_6711,N_6609);
nand U7221 (N_7221,N_6008,N_6675);
and U7222 (N_7222,N_6173,N_6716);
xor U7223 (N_7223,N_6215,N_6560);
or U7224 (N_7224,N_6549,N_6334);
or U7225 (N_7225,N_6624,N_6109);
nand U7226 (N_7226,N_6701,N_6255);
nand U7227 (N_7227,N_6161,N_6099);
nor U7228 (N_7228,N_6114,N_6130);
xnor U7229 (N_7229,N_6390,N_6600);
xor U7230 (N_7230,N_6103,N_6492);
and U7231 (N_7231,N_6708,N_6399);
or U7232 (N_7232,N_6271,N_6710);
nor U7233 (N_7233,N_6598,N_6551);
or U7234 (N_7234,N_6444,N_6321);
nand U7235 (N_7235,N_6480,N_6032);
xnor U7236 (N_7236,N_6020,N_6123);
nor U7237 (N_7237,N_6466,N_6143);
nand U7238 (N_7238,N_6426,N_6079);
nand U7239 (N_7239,N_6276,N_6471);
or U7240 (N_7240,N_6331,N_6440);
nor U7241 (N_7241,N_6021,N_6382);
nand U7242 (N_7242,N_6347,N_6210);
nand U7243 (N_7243,N_6233,N_6066);
nand U7244 (N_7244,N_6387,N_6036);
nand U7245 (N_7245,N_6153,N_6319);
or U7246 (N_7246,N_6187,N_6123);
nand U7247 (N_7247,N_6395,N_6339);
xnor U7248 (N_7248,N_6261,N_6100);
nand U7249 (N_7249,N_6332,N_6564);
nor U7250 (N_7250,N_6720,N_6100);
nand U7251 (N_7251,N_6152,N_6467);
nor U7252 (N_7252,N_6198,N_6051);
xor U7253 (N_7253,N_6114,N_6028);
nand U7254 (N_7254,N_6694,N_6674);
or U7255 (N_7255,N_6186,N_6398);
or U7256 (N_7256,N_6407,N_6371);
and U7257 (N_7257,N_6216,N_6229);
nand U7258 (N_7258,N_6610,N_6587);
or U7259 (N_7259,N_6414,N_6370);
or U7260 (N_7260,N_6595,N_6467);
nand U7261 (N_7261,N_6665,N_6175);
nand U7262 (N_7262,N_6280,N_6557);
nand U7263 (N_7263,N_6277,N_6677);
and U7264 (N_7264,N_6333,N_6581);
xnor U7265 (N_7265,N_6691,N_6719);
and U7266 (N_7266,N_6072,N_6543);
or U7267 (N_7267,N_6137,N_6534);
nand U7268 (N_7268,N_6471,N_6185);
nand U7269 (N_7269,N_6731,N_6647);
nand U7270 (N_7270,N_6316,N_6550);
or U7271 (N_7271,N_6374,N_6332);
xor U7272 (N_7272,N_6416,N_6642);
xor U7273 (N_7273,N_6449,N_6681);
xnor U7274 (N_7274,N_6373,N_6039);
nor U7275 (N_7275,N_6433,N_6354);
nor U7276 (N_7276,N_6378,N_6121);
xnor U7277 (N_7277,N_6272,N_6537);
or U7278 (N_7278,N_6325,N_6613);
nand U7279 (N_7279,N_6104,N_6374);
nand U7280 (N_7280,N_6058,N_6572);
xnor U7281 (N_7281,N_6273,N_6714);
or U7282 (N_7282,N_6591,N_6038);
nor U7283 (N_7283,N_6509,N_6013);
or U7284 (N_7284,N_6297,N_6503);
or U7285 (N_7285,N_6487,N_6389);
or U7286 (N_7286,N_6217,N_6156);
xnor U7287 (N_7287,N_6629,N_6599);
nand U7288 (N_7288,N_6658,N_6033);
or U7289 (N_7289,N_6265,N_6597);
or U7290 (N_7290,N_6018,N_6701);
and U7291 (N_7291,N_6277,N_6193);
and U7292 (N_7292,N_6564,N_6402);
nand U7293 (N_7293,N_6626,N_6487);
or U7294 (N_7294,N_6430,N_6095);
nand U7295 (N_7295,N_6405,N_6501);
or U7296 (N_7296,N_6673,N_6578);
and U7297 (N_7297,N_6343,N_6347);
and U7298 (N_7298,N_6034,N_6405);
and U7299 (N_7299,N_6665,N_6590);
and U7300 (N_7300,N_6627,N_6517);
nand U7301 (N_7301,N_6635,N_6622);
nand U7302 (N_7302,N_6469,N_6284);
xor U7303 (N_7303,N_6527,N_6309);
or U7304 (N_7304,N_6633,N_6533);
or U7305 (N_7305,N_6040,N_6178);
and U7306 (N_7306,N_6221,N_6085);
and U7307 (N_7307,N_6496,N_6022);
xor U7308 (N_7308,N_6675,N_6501);
or U7309 (N_7309,N_6123,N_6218);
and U7310 (N_7310,N_6596,N_6593);
nor U7311 (N_7311,N_6711,N_6587);
and U7312 (N_7312,N_6383,N_6525);
xnor U7313 (N_7313,N_6025,N_6662);
xnor U7314 (N_7314,N_6024,N_6406);
nor U7315 (N_7315,N_6564,N_6000);
xnor U7316 (N_7316,N_6226,N_6538);
xor U7317 (N_7317,N_6445,N_6041);
and U7318 (N_7318,N_6001,N_6343);
and U7319 (N_7319,N_6116,N_6604);
and U7320 (N_7320,N_6716,N_6506);
nor U7321 (N_7321,N_6393,N_6548);
nor U7322 (N_7322,N_6542,N_6007);
or U7323 (N_7323,N_6446,N_6003);
xnor U7324 (N_7324,N_6349,N_6015);
nand U7325 (N_7325,N_6725,N_6277);
xor U7326 (N_7326,N_6131,N_6023);
xor U7327 (N_7327,N_6025,N_6364);
nor U7328 (N_7328,N_6292,N_6630);
and U7329 (N_7329,N_6619,N_6612);
or U7330 (N_7330,N_6113,N_6118);
or U7331 (N_7331,N_6693,N_6433);
or U7332 (N_7332,N_6667,N_6670);
nor U7333 (N_7333,N_6413,N_6636);
and U7334 (N_7334,N_6081,N_6027);
xnor U7335 (N_7335,N_6440,N_6618);
nor U7336 (N_7336,N_6611,N_6606);
xor U7337 (N_7337,N_6004,N_6592);
nand U7338 (N_7338,N_6741,N_6353);
or U7339 (N_7339,N_6351,N_6288);
or U7340 (N_7340,N_6129,N_6402);
and U7341 (N_7341,N_6286,N_6455);
nand U7342 (N_7342,N_6119,N_6186);
xor U7343 (N_7343,N_6516,N_6466);
nand U7344 (N_7344,N_6576,N_6353);
xor U7345 (N_7345,N_6718,N_6731);
or U7346 (N_7346,N_6585,N_6560);
or U7347 (N_7347,N_6022,N_6187);
and U7348 (N_7348,N_6711,N_6333);
and U7349 (N_7349,N_6326,N_6469);
nand U7350 (N_7350,N_6135,N_6086);
nand U7351 (N_7351,N_6540,N_6743);
or U7352 (N_7352,N_6382,N_6441);
nor U7353 (N_7353,N_6195,N_6496);
or U7354 (N_7354,N_6541,N_6232);
xor U7355 (N_7355,N_6211,N_6007);
nor U7356 (N_7356,N_6042,N_6435);
xnor U7357 (N_7357,N_6188,N_6512);
nor U7358 (N_7358,N_6021,N_6043);
and U7359 (N_7359,N_6636,N_6664);
nand U7360 (N_7360,N_6451,N_6093);
and U7361 (N_7361,N_6465,N_6114);
nor U7362 (N_7362,N_6091,N_6259);
nor U7363 (N_7363,N_6059,N_6383);
nor U7364 (N_7364,N_6749,N_6743);
or U7365 (N_7365,N_6611,N_6382);
or U7366 (N_7366,N_6567,N_6045);
and U7367 (N_7367,N_6675,N_6650);
nor U7368 (N_7368,N_6264,N_6008);
nand U7369 (N_7369,N_6323,N_6375);
nor U7370 (N_7370,N_6433,N_6150);
xor U7371 (N_7371,N_6378,N_6179);
nand U7372 (N_7372,N_6164,N_6668);
and U7373 (N_7373,N_6499,N_6467);
nand U7374 (N_7374,N_6350,N_6487);
and U7375 (N_7375,N_6155,N_6679);
xnor U7376 (N_7376,N_6714,N_6442);
nor U7377 (N_7377,N_6576,N_6735);
or U7378 (N_7378,N_6496,N_6394);
nand U7379 (N_7379,N_6679,N_6184);
nor U7380 (N_7380,N_6223,N_6120);
and U7381 (N_7381,N_6327,N_6517);
or U7382 (N_7382,N_6628,N_6169);
and U7383 (N_7383,N_6593,N_6297);
and U7384 (N_7384,N_6031,N_6691);
nor U7385 (N_7385,N_6332,N_6329);
xnor U7386 (N_7386,N_6534,N_6071);
or U7387 (N_7387,N_6007,N_6589);
or U7388 (N_7388,N_6287,N_6720);
nor U7389 (N_7389,N_6113,N_6484);
or U7390 (N_7390,N_6722,N_6020);
nand U7391 (N_7391,N_6263,N_6643);
or U7392 (N_7392,N_6330,N_6327);
and U7393 (N_7393,N_6359,N_6241);
xor U7394 (N_7394,N_6428,N_6700);
nor U7395 (N_7395,N_6583,N_6392);
xnor U7396 (N_7396,N_6400,N_6094);
and U7397 (N_7397,N_6371,N_6037);
nand U7398 (N_7398,N_6744,N_6653);
nand U7399 (N_7399,N_6602,N_6175);
nor U7400 (N_7400,N_6537,N_6626);
nor U7401 (N_7401,N_6664,N_6142);
or U7402 (N_7402,N_6647,N_6738);
or U7403 (N_7403,N_6169,N_6231);
or U7404 (N_7404,N_6589,N_6545);
nor U7405 (N_7405,N_6503,N_6079);
or U7406 (N_7406,N_6499,N_6011);
nand U7407 (N_7407,N_6045,N_6067);
xor U7408 (N_7408,N_6726,N_6450);
or U7409 (N_7409,N_6205,N_6668);
nand U7410 (N_7410,N_6546,N_6723);
xnor U7411 (N_7411,N_6393,N_6649);
nand U7412 (N_7412,N_6264,N_6514);
and U7413 (N_7413,N_6638,N_6660);
or U7414 (N_7414,N_6427,N_6322);
xnor U7415 (N_7415,N_6446,N_6553);
or U7416 (N_7416,N_6549,N_6734);
xnor U7417 (N_7417,N_6243,N_6510);
xnor U7418 (N_7418,N_6051,N_6444);
nor U7419 (N_7419,N_6313,N_6176);
nor U7420 (N_7420,N_6489,N_6042);
xor U7421 (N_7421,N_6095,N_6263);
and U7422 (N_7422,N_6311,N_6529);
xor U7423 (N_7423,N_6616,N_6013);
xor U7424 (N_7424,N_6229,N_6697);
and U7425 (N_7425,N_6090,N_6344);
or U7426 (N_7426,N_6553,N_6585);
and U7427 (N_7427,N_6033,N_6037);
nor U7428 (N_7428,N_6509,N_6103);
or U7429 (N_7429,N_6182,N_6076);
xnor U7430 (N_7430,N_6015,N_6325);
nor U7431 (N_7431,N_6470,N_6031);
xnor U7432 (N_7432,N_6285,N_6127);
nand U7433 (N_7433,N_6619,N_6184);
or U7434 (N_7434,N_6123,N_6497);
nor U7435 (N_7435,N_6319,N_6029);
and U7436 (N_7436,N_6083,N_6722);
xor U7437 (N_7437,N_6361,N_6674);
xnor U7438 (N_7438,N_6198,N_6050);
or U7439 (N_7439,N_6141,N_6227);
and U7440 (N_7440,N_6237,N_6466);
xnor U7441 (N_7441,N_6025,N_6353);
nor U7442 (N_7442,N_6106,N_6060);
nor U7443 (N_7443,N_6383,N_6214);
and U7444 (N_7444,N_6005,N_6033);
or U7445 (N_7445,N_6711,N_6448);
xor U7446 (N_7446,N_6675,N_6715);
nor U7447 (N_7447,N_6300,N_6534);
or U7448 (N_7448,N_6320,N_6357);
nand U7449 (N_7449,N_6149,N_6282);
nor U7450 (N_7450,N_6630,N_6730);
nor U7451 (N_7451,N_6381,N_6070);
or U7452 (N_7452,N_6188,N_6598);
xor U7453 (N_7453,N_6497,N_6136);
nor U7454 (N_7454,N_6556,N_6627);
and U7455 (N_7455,N_6672,N_6076);
or U7456 (N_7456,N_6524,N_6162);
or U7457 (N_7457,N_6712,N_6047);
and U7458 (N_7458,N_6722,N_6220);
nor U7459 (N_7459,N_6340,N_6538);
nor U7460 (N_7460,N_6173,N_6743);
nand U7461 (N_7461,N_6709,N_6494);
and U7462 (N_7462,N_6173,N_6669);
xor U7463 (N_7463,N_6409,N_6544);
nor U7464 (N_7464,N_6619,N_6703);
and U7465 (N_7465,N_6355,N_6628);
nor U7466 (N_7466,N_6070,N_6605);
nand U7467 (N_7467,N_6617,N_6625);
and U7468 (N_7468,N_6413,N_6564);
nor U7469 (N_7469,N_6341,N_6026);
and U7470 (N_7470,N_6067,N_6372);
or U7471 (N_7471,N_6281,N_6429);
xor U7472 (N_7472,N_6512,N_6316);
nand U7473 (N_7473,N_6327,N_6545);
or U7474 (N_7474,N_6534,N_6030);
or U7475 (N_7475,N_6147,N_6199);
or U7476 (N_7476,N_6430,N_6107);
xnor U7477 (N_7477,N_6075,N_6602);
nor U7478 (N_7478,N_6594,N_6250);
nor U7479 (N_7479,N_6127,N_6212);
or U7480 (N_7480,N_6437,N_6719);
xor U7481 (N_7481,N_6117,N_6050);
nand U7482 (N_7482,N_6609,N_6303);
nor U7483 (N_7483,N_6704,N_6144);
xnor U7484 (N_7484,N_6435,N_6406);
nand U7485 (N_7485,N_6636,N_6558);
nor U7486 (N_7486,N_6656,N_6730);
nor U7487 (N_7487,N_6561,N_6569);
or U7488 (N_7488,N_6667,N_6207);
nor U7489 (N_7489,N_6313,N_6620);
and U7490 (N_7490,N_6545,N_6179);
or U7491 (N_7491,N_6437,N_6362);
nand U7492 (N_7492,N_6598,N_6438);
nand U7493 (N_7493,N_6205,N_6593);
nand U7494 (N_7494,N_6378,N_6692);
nand U7495 (N_7495,N_6598,N_6420);
nor U7496 (N_7496,N_6230,N_6331);
nand U7497 (N_7497,N_6237,N_6329);
nor U7498 (N_7498,N_6389,N_6293);
xor U7499 (N_7499,N_6638,N_6429);
nand U7500 (N_7500,N_7219,N_6765);
xor U7501 (N_7501,N_6970,N_7190);
nand U7502 (N_7502,N_7448,N_6793);
and U7503 (N_7503,N_7263,N_6859);
xnor U7504 (N_7504,N_7353,N_6821);
or U7505 (N_7505,N_7460,N_7212);
xnor U7506 (N_7506,N_7282,N_7450);
and U7507 (N_7507,N_7485,N_6911);
xnor U7508 (N_7508,N_7453,N_6833);
or U7509 (N_7509,N_6852,N_6902);
or U7510 (N_7510,N_7250,N_7126);
xor U7511 (N_7511,N_7171,N_6758);
xor U7512 (N_7512,N_6941,N_7444);
and U7513 (N_7513,N_7103,N_7370);
or U7514 (N_7514,N_7314,N_6888);
or U7515 (N_7515,N_6994,N_7050);
nand U7516 (N_7516,N_6950,N_7145);
xnor U7517 (N_7517,N_7328,N_7043);
or U7518 (N_7518,N_7333,N_6928);
or U7519 (N_7519,N_6820,N_7120);
or U7520 (N_7520,N_6894,N_7433);
nor U7521 (N_7521,N_6929,N_7170);
and U7522 (N_7522,N_6880,N_7028);
nor U7523 (N_7523,N_7494,N_7239);
nand U7524 (N_7524,N_6862,N_7240);
xnor U7525 (N_7525,N_7369,N_6787);
nand U7526 (N_7526,N_7044,N_7217);
xnor U7527 (N_7527,N_7130,N_7462);
nor U7528 (N_7528,N_7270,N_7306);
or U7529 (N_7529,N_7286,N_7459);
xor U7530 (N_7530,N_6913,N_7027);
xnor U7531 (N_7531,N_7200,N_7291);
xor U7532 (N_7532,N_7260,N_7072);
nand U7533 (N_7533,N_6799,N_7497);
or U7534 (N_7534,N_6891,N_7268);
xnor U7535 (N_7535,N_6858,N_6757);
nand U7536 (N_7536,N_7408,N_7352);
nor U7537 (N_7537,N_7019,N_7151);
nand U7538 (N_7538,N_6770,N_7054);
nor U7539 (N_7539,N_6829,N_7199);
nand U7540 (N_7540,N_6752,N_7457);
xnor U7541 (N_7541,N_6936,N_6992);
and U7542 (N_7542,N_7318,N_7451);
xnor U7543 (N_7543,N_7482,N_7074);
xor U7544 (N_7544,N_6877,N_6952);
nor U7545 (N_7545,N_7376,N_7039);
nand U7546 (N_7546,N_6791,N_6882);
xnor U7547 (N_7547,N_7499,N_6892);
nand U7548 (N_7548,N_7165,N_7473);
nor U7549 (N_7549,N_7022,N_7327);
nor U7550 (N_7550,N_7234,N_7104);
nor U7551 (N_7551,N_7128,N_7017);
nand U7552 (N_7552,N_7413,N_7067);
nand U7553 (N_7553,N_7096,N_7026);
xor U7554 (N_7554,N_6767,N_7066);
and U7555 (N_7555,N_7311,N_6938);
nand U7556 (N_7556,N_6860,N_6873);
or U7557 (N_7557,N_6934,N_6867);
and U7558 (N_7558,N_7317,N_7257);
and U7559 (N_7559,N_6993,N_7015);
nand U7560 (N_7560,N_7107,N_6750);
and U7561 (N_7561,N_6930,N_6908);
and U7562 (N_7562,N_7059,N_6948);
nand U7563 (N_7563,N_6960,N_7225);
or U7564 (N_7564,N_7078,N_7228);
nand U7565 (N_7565,N_7038,N_7283);
nand U7566 (N_7566,N_7351,N_7011);
or U7567 (N_7567,N_7407,N_7127);
nand U7568 (N_7568,N_7492,N_7479);
and U7569 (N_7569,N_7045,N_7255);
nand U7570 (N_7570,N_6887,N_6837);
and U7571 (N_7571,N_7013,N_6853);
nand U7572 (N_7572,N_7428,N_7266);
and U7573 (N_7573,N_7300,N_7297);
nand U7574 (N_7574,N_7086,N_7055);
xor U7575 (N_7575,N_7491,N_7105);
nor U7576 (N_7576,N_7033,N_6855);
xnor U7577 (N_7577,N_7488,N_7337);
nand U7578 (N_7578,N_6847,N_7301);
xnor U7579 (N_7579,N_7242,N_6806);
nand U7580 (N_7580,N_6940,N_7336);
nand U7581 (N_7581,N_7204,N_7342);
or U7582 (N_7582,N_7247,N_7281);
or U7583 (N_7583,N_7160,N_6762);
nor U7584 (N_7584,N_6983,N_7395);
xnor U7585 (N_7585,N_6916,N_7032);
and U7586 (N_7586,N_6876,N_7269);
nand U7587 (N_7587,N_6985,N_7070);
nand U7588 (N_7588,N_7287,N_6818);
xnor U7589 (N_7589,N_7476,N_7495);
and U7590 (N_7590,N_6907,N_7076);
or U7591 (N_7591,N_6986,N_7243);
nand U7592 (N_7592,N_7422,N_6984);
or U7593 (N_7593,N_6857,N_6832);
nor U7594 (N_7594,N_6807,N_6999);
or U7595 (N_7595,N_7463,N_6898);
and U7596 (N_7596,N_6954,N_7423);
xor U7597 (N_7597,N_7124,N_7275);
and U7598 (N_7598,N_7177,N_6964);
and U7599 (N_7599,N_6966,N_7335);
nor U7600 (N_7600,N_6760,N_7053);
or U7601 (N_7601,N_6864,N_7440);
and U7602 (N_7602,N_7374,N_7155);
xnor U7603 (N_7603,N_6845,N_7009);
xor U7604 (N_7604,N_7321,N_6878);
nand U7605 (N_7605,N_7248,N_6872);
nor U7606 (N_7606,N_7475,N_7345);
nand U7607 (N_7607,N_6794,N_6951);
or U7608 (N_7608,N_7144,N_7489);
xnor U7609 (N_7609,N_6819,N_7481);
and U7610 (N_7610,N_7496,N_6896);
xor U7611 (N_7611,N_7343,N_7386);
xor U7612 (N_7612,N_7304,N_6836);
nor U7613 (N_7613,N_7418,N_7088);
or U7614 (N_7614,N_7073,N_6967);
or U7615 (N_7615,N_6927,N_6924);
nor U7616 (N_7616,N_7172,N_6763);
or U7617 (N_7617,N_7349,N_7195);
or U7618 (N_7618,N_6841,N_7010);
xor U7619 (N_7619,N_7480,N_7285);
nand U7620 (N_7620,N_6849,N_7427);
nor U7621 (N_7621,N_7307,N_6904);
or U7622 (N_7622,N_7157,N_6842);
or U7623 (N_7623,N_6766,N_7261);
and U7624 (N_7624,N_7143,N_7443);
xor U7625 (N_7625,N_7030,N_7042);
xnor U7626 (N_7626,N_6775,N_6825);
nor U7627 (N_7627,N_6823,N_6844);
nor U7628 (N_7628,N_7372,N_7135);
and U7629 (N_7629,N_6759,N_6835);
or U7630 (N_7630,N_7452,N_7003);
nand U7631 (N_7631,N_7310,N_7487);
or U7632 (N_7632,N_6895,N_7246);
nor U7633 (N_7633,N_7071,N_7419);
or U7634 (N_7634,N_7005,N_6786);
xnor U7635 (N_7635,N_6871,N_7409);
nand U7636 (N_7636,N_7431,N_7467);
xnor U7637 (N_7637,N_7305,N_7137);
or U7638 (N_7638,N_7278,N_7233);
or U7639 (N_7639,N_7062,N_7154);
xor U7640 (N_7640,N_6785,N_6885);
or U7641 (N_7641,N_6834,N_7194);
xnor U7642 (N_7642,N_7102,N_6809);
nor U7643 (N_7643,N_7312,N_7432);
nor U7644 (N_7644,N_7118,N_7169);
or U7645 (N_7645,N_7037,N_7414);
nor U7646 (N_7646,N_7403,N_7398);
nor U7647 (N_7647,N_7141,N_7220);
or U7648 (N_7648,N_6863,N_7394);
or U7649 (N_7649,N_6840,N_7158);
or U7650 (N_7650,N_7437,N_7230);
nand U7651 (N_7651,N_7175,N_6771);
and U7652 (N_7652,N_7081,N_7012);
and U7653 (N_7653,N_7184,N_6980);
xor U7654 (N_7654,N_6805,N_6991);
xnor U7655 (N_7655,N_6764,N_6774);
xor U7656 (N_7656,N_7400,N_6797);
nand U7657 (N_7657,N_7093,N_7371);
nand U7658 (N_7658,N_6843,N_7138);
xnor U7659 (N_7659,N_6811,N_7430);
xnor U7660 (N_7660,N_7173,N_7415);
nand U7661 (N_7661,N_6953,N_7231);
and U7662 (N_7662,N_7139,N_7302);
or U7663 (N_7663,N_6995,N_6889);
nand U7664 (N_7664,N_7410,N_7441);
and U7665 (N_7665,N_6933,N_6879);
nand U7666 (N_7666,N_7202,N_6976);
xnor U7667 (N_7667,N_7241,N_6925);
or U7668 (N_7668,N_7316,N_7092);
nor U7669 (N_7669,N_6893,N_6920);
nor U7670 (N_7670,N_7186,N_7446);
nand U7671 (N_7671,N_6881,N_7229);
xor U7672 (N_7672,N_7163,N_7429);
or U7673 (N_7673,N_7363,N_6866);
nand U7674 (N_7674,N_7252,N_6814);
nand U7675 (N_7675,N_7256,N_6909);
nand U7676 (N_7676,N_7134,N_7399);
nand U7677 (N_7677,N_7277,N_7346);
xnor U7678 (N_7678,N_7004,N_7434);
nor U7679 (N_7679,N_7035,N_7136);
nor U7680 (N_7680,N_7332,N_6949);
or U7681 (N_7681,N_6804,N_7490);
or U7682 (N_7682,N_7174,N_7162);
xor U7683 (N_7683,N_6973,N_6861);
and U7684 (N_7684,N_6946,N_7357);
xor U7685 (N_7685,N_7356,N_7320);
nor U7686 (N_7686,N_7344,N_7461);
or U7687 (N_7687,N_7361,N_7358);
nor U7688 (N_7688,N_6795,N_7486);
or U7689 (N_7689,N_6828,N_6754);
or U7690 (N_7690,N_6851,N_6988);
and U7691 (N_7691,N_6977,N_7117);
nand U7692 (N_7692,N_6957,N_7132);
and U7693 (N_7693,N_7040,N_7365);
nand U7694 (N_7694,N_7087,N_6974);
xor U7695 (N_7695,N_6796,N_7329);
and U7696 (N_7696,N_6782,N_7056);
xor U7697 (N_7697,N_6962,N_6827);
and U7698 (N_7698,N_7036,N_7292);
xor U7699 (N_7699,N_6943,N_6884);
or U7700 (N_7700,N_7483,N_7471);
nand U7701 (N_7701,N_7382,N_7390);
nor U7702 (N_7702,N_7142,N_7447);
nor U7703 (N_7703,N_7227,N_7469);
or U7704 (N_7704,N_7235,N_7161);
nand U7705 (N_7705,N_7341,N_7378);
nand U7706 (N_7706,N_7290,N_7082);
and U7707 (N_7707,N_7330,N_7384);
nand U7708 (N_7708,N_7181,N_6839);
or U7709 (N_7709,N_7455,N_6917);
xor U7710 (N_7710,N_6987,N_7191);
and U7711 (N_7711,N_7421,N_7426);
xnor U7712 (N_7712,N_7084,N_6926);
and U7713 (N_7713,N_6846,N_6815);
nor U7714 (N_7714,N_7046,N_6975);
nor U7715 (N_7715,N_7065,N_7198);
or U7716 (N_7716,N_7299,N_7416);
nand U7717 (N_7717,N_7014,N_6777);
xor U7718 (N_7718,N_7484,N_6778);
nor U7719 (N_7719,N_7354,N_7392);
xnor U7720 (N_7720,N_7339,N_7322);
nand U7721 (N_7721,N_7366,N_6810);
xor U7722 (N_7722,N_7420,N_7276);
and U7723 (N_7723,N_7034,N_7208);
xor U7724 (N_7724,N_7064,N_7449);
or U7725 (N_7725,N_7406,N_7466);
xor U7726 (N_7726,N_7188,N_6856);
xnor U7727 (N_7727,N_7213,N_7383);
nand U7728 (N_7728,N_7123,N_7401);
xnor U7729 (N_7729,N_6923,N_7244);
or U7730 (N_7730,N_7493,N_7280);
xor U7731 (N_7731,N_6921,N_7267);
nor U7732 (N_7732,N_7016,N_7001);
and U7733 (N_7733,N_7180,N_6808);
xor U7734 (N_7734,N_7131,N_6822);
or U7735 (N_7735,N_6761,N_7355);
nor U7736 (N_7736,N_7264,N_7458);
nor U7737 (N_7737,N_6997,N_7176);
or U7738 (N_7738,N_7211,N_6769);
nor U7739 (N_7739,N_7079,N_7101);
nor U7740 (N_7740,N_6935,N_7417);
xnor U7741 (N_7741,N_7115,N_7197);
and U7742 (N_7742,N_7007,N_6803);
xnor U7743 (N_7743,N_7253,N_6961);
nor U7744 (N_7744,N_7122,N_6798);
or U7745 (N_7745,N_7379,N_7439);
or U7746 (N_7746,N_7309,N_7298);
or U7747 (N_7747,N_6801,N_6830);
or U7748 (N_7748,N_7214,N_7498);
nor U7749 (N_7749,N_7405,N_7391);
and U7750 (N_7750,N_7058,N_7098);
nor U7751 (N_7751,N_7156,N_7245);
and U7752 (N_7752,N_6918,N_7221);
and U7753 (N_7753,N_7119,N_7116);
nand U7754 (N_7754,N_7296,N_7259);
nand U7755 (N_7755,N_6919,N_6932);
xor U7756 (N_7756,N_7129,N_6812);
nand U7757 (N_7757,N_7152,N_7097);
nand U7758 (N_7758,N_7274,N_7293);
nor U7759 (N_7759,N_7367,N_7273);
xnor U7760 (N_7760,N_6989,N_6912);
nand U7761 (N_7761,N_7080,N_7089);
xor U7762 (N_7762,N_7167,N_7251);
nor U7763 (N_7763,N_6897,N_7090);
xnor U7764 (N_7764,N_6968,N_7023);
nor U7765 (N_7765,N_7049,N_7404);
xnor U7766 (N_7766,N_7334,N_7477);
and U7767 (N_7767,N_7393,N_7438);
and U7768 (N_7768,N_7468,N_7381);
and U7769 (N_7769,N_7373,N_7362);
nand U7770 (N_7770,N_7435,N_6751);
or U7771 (N_7771,N_7020,N_6824);
nand U7772 (N_7772,N_7470,N_7295);
xor U7773 (N_7773,N_7402,N_6788);
nand U7774 (N_7774,N_7085,N_7187);
xor U7775 (N_7775,N_6959,N_7031);
nand U7776 (N_7776,N_7340,N_7024);
and U7777 (N_7777,N_6756,N_6958);
xnor U7778 (N_7778,N_7068,N_7052);
xnor U7779 (N_7779,N_6813,N_6792);
nor U7780 (N_7780,N_6955,N_6773);
nand U7781 (N_7781,N_7121,N_7232);
and U7782 (N_7782,N_6890,N_7226);
xnor U7783 (N_7783,N_6915,N_7478);
and U7784 (N_7784,N_7193,N_7325);
or U7785 (N_7785,N_7380,N_7289);
and U7786 (N_7786,N_6875,N_7223);
xor U7787 (N_7787,N_7436,N_7347);
xnor U7788 (N_7788,N_7094,N_7178);
xnor U7789 (N_7789,N_7008,N_7218);
and U7790 (N_7790,N_7140,N_7359);
or U7791 (N_7791,N_6865,N_7047);
nand U7792 (N_7792,N_6945,N_7150);
nor U7793 (N_7793,N_7196,N_7396);
nor U7794 (N_7794,N_7029,N_7166);
xor U7795 (N_7795,N_6906,N_7474);
and U7796 (N_7796,N_7083,N_6874);
or U7797 (N_7797,N_6768,N_6789);
nor U7798 (N_7798,N_7313,N_7271);
nand U7799 (N_7799,N_7111,N_7108);
nor U7800 (N_7800,N_7018,N_6998);
xnor U7801 (N_7801,N_7206,N_6922);
nor U7802 (N_7802,N_7210,N_7075);
nand U7803 (N_7803,N_7060,N_6790);
and U7804 (N_7804,N_6850,N_6854);
nor U7805 (N_7805,N_7249,N_7388);
nand U7806 (N_7806,N_6753,N_6883);
xnor U7807 (N_7807,N_6870,N_7360);
or U7808 (N_7808,N_6905,N_6779);
nand U7809 (N_7809,N_7308,N_7303);
and U7810 (N_7810,N_6965,N_6971);
nor U7811 (N_7811,N_6931,N_7222);
nand U7812 (N_7812,N_7215,N_7051);
or U7813 (N_7813,N_6848,N_7099);
and U7814 (N_7814,N_7442,N_7364);
or U7815 (N_7815,N_6972,N_6910);
xor U7816 (N_7816,N_7201,N_7182);
nor U7817 (N_7817,N_7472,N_7025);
nand U7818 (N_7818,N_7385,N_6990);
nor U7819 (N_7819,N_6963,N_7041);
nand U7820 (N_7820,N_7254,N_6755);
nor U7821 (N_7821,N_7057,N_7265);
and U7822 (N_7822,N_7323,N_7324);
or U7823 (N_7823,N_6800,N_7209);
nand U7824 (N_7824,N_7189,N_7284);
xor U7825 (N_7825,N_7109,N_7113);
or U7826 (N_7826,N_7133,N_7465);
and U7827 (N_7827,N_7192,N_7179);
or U7828 (N_7828,N_6996,N_6868);
nor U7829 (N_7829,N_6900,N_7000);
and U7830 (N_7830,N_7100,N_6939);
nor U7831 (N_7831,N_6979,N_6982);
nor U7832 (N_7832,N_7464,N_6816);
or U7833 (N_7833,N_6886,N_7368);
or U7834 (N_7834,N_7203,N_7456);
and U7835 (N_7835,N_7091,N_7061);
nor U7836 (N_7836,N_7411,N_6869);
and U7837 (N_7837,N_7153,N_6981);
xnor U7838 (N_7838,N_7216,N_7224);
or U7839 (N_7839,N_7006,N_7205);
nor U7840 (N_7840,N_7389,N_7021);
nor U7841 (N_7841,N_7319,N_7294);
nor U7842 (N_7842,N_7112,N_6817);
or U7843 (N_7843,N_6784,N_7149);
and U7844 (N_7844,N_7164,N_6781);
or U7845 (N_7845,N_6826,N_7454);
and U7846 (N_7846,N_6776,N_7350);
nand U7847 (N_7847,N_7183,N_7114);
xor U7848 (N_7848,N_7425,N_7146);
nor U7849 (N_7849,N_7207,N_7168);
or U7850 (N_7850,N_6903,N_7326);
or U7851 (N_7851,N_6831,N_6838);
xor U7852 (N_7852,N_6901,N_7110);
nor U7853 (N_7853,N_7397,N_6802);
or U7854 (N_7854,N_7445,N_7185);
or U7855 (N_7855,N_7063,N_6944);
xor U7856 (N_7856,N_7315,N_7095);
nand U7857 (N_7857,N_7338,N_7377);
and U7858 (N_7858,N_6780,N_7375);
xor U7859 (N_7859,N_7002,N_7148);
or U7860 (N_7860,N_6772,N_7069);
nand U7861 (N_7861,N_7279,N_6937);
nor U7862 (N_7862,N_7348,N_7262);
and U7863 (N_7863,N_6914,N_7258);
and U7864 (N_7864,N_7331,N_6969);
xnor U7865 (N_7865,N_7288,N_6942);
or U7866 (N_7866,N_7387,N_7238);
nor U7867 (N_7867,N_7412,N_6978);
nor U7868 (N_7868,N_7077,N_7272);
nor U7869 (N_7869,N_7147,N_6956);
nor U7870 (N_7870,N_7424,N_7237);
and U7871 (N_7871,N_6899,N_6947);
xnor U7872 (N_7872,N_7125,N_6783);
nand U7873 (N_7873,N_7236,N_7159);
xnor U7874 (N_7874,N_7048,N_7106);
and U7875 (N_7875,N_7268,N_6869);
and U7876 (N_7876,N_6814,N_7064);
nand U7877 (N_7877,N_7495,N_7468);
nor U7878 (N_7878,N_7496,N_7179);
xnor U7879 (N_7879,N_7246,N_7347);
or U7880 (N_7880,N_6814,N_6954);
xor U7881 (N_7881,N_7479,N_7083);
and U7882 (N_7882,N_7126,N_7319);
nand U7883 (N_7883,N_7109,N_6947);
nor U7884 (N_7884,N_7177,N_7142);
xor U7885 (N_7885,N_6969,N_6872);
xnor U7886 (N_7886,N_7018,N_7314);
nor U7887 (N_7887,N_7190,N_6838);
xnor U7888 (N_7888,N_6995,N_6964);
and U7889 (N_7889,N_6855,N_7146);
nor U7890 (N_7890,N_6918,N_7310);
nor U7891 (N_7891,N_7011,N_7362);
nand U7892 (N_7892,N_7169,N_7341);
nor U7893 (N_7893,N_6915,N_7172);
xor U7894 (N_7894,N_7411,N_7087);
xor U7895 (N_7895,N_7034,N_7190);
and U7896 (N_7896,N_7100,N_7031);
xor U7897 (N_7897,N_6996,N_7024);
nor U7898 (N_7898,N_7399,N_7275);
xor U7899 (N_7899,N_7468,N_6954);
nand U7900 (N_7900,N_6996,N_7004);
and U7901 (N_7901,N_7026,N_6783);
nor U7902 (N_7902,N_7158,N_6943);
xor U7903 (N_7903,N_7345,N_7220);
and U7904 (N_7904,N_7442,N_7321);
xor U7905 (N_7905,N_7480,N_7365);
nor U7906 (N_7906,N_7237,N_6799);
and U7907 (N_7907,N_7146,N_7406);
xnor U7908 (N_7908,N_7348,N_6770);
xnor U7909 (N_7909,N_7163,N_6778);
xor U7910 (N_7910,N_7389,N_6751);
and U7911 (N_7911,N_7186,N_7481);
nor U7912 (N_7912,N_6974,N_7109);
and U7913 (N_7913,N_7055,N_7433);
nand U7914 (N_7914,N_7389,N_7356);
nor U7915 (N_7915,N_7135,N_7282);
nor U7916 (N_7916,N_6876,N_7165);
xor U7917 (N_7917,N_6777,N_6774);
nor U7918 (N_7918,N_6863,N_6761);
and U7919 (N_7919,N_7393,N_7432);
or U7920 (N_7920,N_6911,N_6882);
nand U7921 (N_7921,N_6759,N_6862);
and U7922 (N_7922,N_7139,N_7046);
or U7923 (N_7923,N_7074,N_7396);
and U7924 (N_7924,N_6866,N_6821);
nor U7925 (N_7925,N_6910,N_6946);
xnor U7926 (N_7926,N_7315,N_6924);
xor U7927 (N_7927,N_7024,N_6951);
and U7928 (N_7928,N_6903,N_7186);
nand U7929 (N_7929,N_7061,N_7294);
and U7930 (N_7930,N_6814,N_7051);
nand U7931 (N_7931,N_7230,N_7245);
nand U7932 (N_7932,N_7490,N_6824);
or U7933 (N_7933,N_7101,N_7472);
xnor U7934 (N_7934,N_6809,N_6849);
xnor U7935 (N_7935,N_7173,N_7300);
nand U7936 (N_7936,N_7401,N_6764);
nor U7937 (N_7937,N_7046,N_6887);
or U7938 (N_7938,N_7390,N_7386);
and U7939 (N_7939,N_7208,N_7399);
nor U7940 (N_7940,N_7182,N_7046);
nand U7941 (N_7941,N_7397,N_7174);
nor U7942 (N_7942,N_7345,N_7105);
or U7943 (N_7943,N_6998,N_6926);
and U7944 (N_7944,N_7276,N_7442);
nor U7945 (N_7945,N_6809,N_7301);
xor U7946 (N_7946,N_7429,N_6993);
xor U7947 (N_7947,N_7444,N_6901);
nor U7948 (N_7948,N_7118,N_6949);
nand U7949 (N_7949,N_7272,N_7273);
or U7950 (N_7950,N_7121,N_7362);
nand U7951 (N_7951,N_7326,N_7163);
or U7952 (N_7952,N_7326,N_6934);
xnor U7953 (N_7953,N_6859,N_7417);
nand U7954 (N_7954,N_7120,N_7004);
and U7955 (N_7955,N_6896,N_6772);
nand U7956 (N_7956,N_7381,N_7136);
xor U7957 (N_7957,N_7064,N_7409);
and U7958 (N_7958,N_6956,N_7213);
or U7959 (N_7959,N_6979,N_7227);
or U7960 (N_7960,N_7093,N_7462);
or U7961 (N_7961,N_7104,N_7319);
and U7962 (N_7962,N_7471,N_7050);
or U7963 (N_7963,N_7247,N_7354);
or U7964 (N_7964,N_7113,N_7341);
nor U7965 (N_7965,N_7365,N_7252);
or U7966 (N_7966,N_6869,N_7049);
nor U7967 (N_7967,N_7076,N_7459);
nor U7968 (N_7968,N_6868,N_7073);
or U7969 (N_7969,N_7452,N_7405);
nor U7970 (N_7970,N_7274,N_6950);
or U7971 (N_7971,N_6919,N_6894);
nand U7972 (N_7972,N_6972,N_7181);
and U7973 (N_7973,N_6761,N_7065);
and U7974 (N_7974,N_6932,N_7158);
nor U7975 (N_7975,N_7469,N_7433);
nor U7976 (N_7976,N_7396,N_7486);
xor U7977 (N_7977,N_7441,N_7452);
and U7978 (N_7978,N_6828,N_7391);
nor U7979 (N_7979,N_7053,N_7161);
and U7980 (N_7980,N_7200,N_6924);
nor U7981 (N_7981,N_7217,N_7490);
nor U7982 (N_7982,N_7424,N_7358);
or U7983 (N_7983,N_6908,N_7161);
xor U7984 (N_7984,N_6999,N_7242);
nand U7985 (N_7985,N_6796,N_6867);
and U7986 (N_7986,N_7344,N_6961);
nor U7987 (N_7987,N_6873,N_6974);
nand U7988 (N_7988,N_7481,N_7373);
xor U7989 (N_7989,N_6967,N_7161);
xnor U7990 (N_7990,N_7234,N_6978);
xnor U7991 (N_7991,N_7112,N_7116);
and U7992 (N_7992,N_7071,N_7099);
nor U7993 (N_7993,N_7113,N_7269);
nand U7994 (N_7994,N_7225,N_7409);
xor U7995 (N_7995,N_7199,N_6789);
or U7996 (N_7996,N_7126,N_6957);
nand U7997 (N_7997,N_6863,N_7225);
and U7998 (N_7998,N_7292,N_6960);
xor U7999 (N_7999,N_7099,N_7295);
or U8000 (N_8000,N_6878,N_6814);
nor U8001 (N_8001,N_6754,N_6885);
or U8002 (N_8002,N_7001,N_7175);
or U8003 (N_8003,N_7058,N_7067);
nand U8004 (N_8004,N_7163,N_7021);
or U8005 (N_8005,N_7494,N_7194);
nand U8006 (N_8006,N_7483,N_7129);
nor U8007 (N_8007,N_7274,N_7158);
nand U8008 (N_8008,N_7049,N_7454);
xnor U8009 (N_8009,N_7255,N_6770);
or U8010 (N_8010,N_7014,N_6812);
nor U8011 (N_8011,N_6787,N_7203);
or U8012 (N_8012,N_7054,N_7227);
or U8013 (N_8013,N_7052,N_7312);
or U8014 (N_8014,N_6932,N_7116);
xnor U8015 (N_8015,N_7022,N_7352);
or U8016 (N_8016,N_7225,N_6888);
xor U8017 (N_8017,N_7322,N_7052);
xor U8018 (N_8018,N_7178,N_7097);
nor U8019 (N_8019,N_7008,N_6851);
xor U8020 (N_8020,N_7372,N_7086);
xor U8021 (N_8021,N_6834,N_7425);
nor U8022 (N_8022,N_7068,N_7272);
nand U8023 (N_8023,N_7353,N_6880);
or U8024 (N_8024,N_6783,N_6819);
nor U8025 (N_8025,N_6803,N_7240);
xnor U8026 (N_8026,N_7037,N_6750);
or U8027 (N_8027,N_7181,N_7490);
and U8028 (N_8028,N_6855,N_7405);
nand U8029 (N_8029,N_6841,N_7179);
nand U8030 (N_8030,N_6775,N_7194);
xnor U8031 (N_8031,N_6867,N_7317);
or U8032 (N_8032,N_7113,N_7238);
and U8033 (N_8033,N_7299,N_6820);
or U8034 (N_8034,N_6914,N_7379);
or U8035 (N_8035,N_7344,N_6894);
and U8036 (N_8036,N_6848,N_6928);
or U8037 (N_8037,N_7450,N_7171);
and U8038 (N_8038,N_7005,N_7068);
nor U8039 (N_8039,N_6794,N_6787);
nand U8040 (N_8040,N_7068,N_7140);
xor U8041 (N_8041,N_6913,N_6873);
nor U8042 (N_8042,N_6896,N_6949);
nor U8043 (N_8043,N_6908,N_7224);
and U8044 (N_8044,N_7240,N_7015);
xor U8045 (N_8045,N_7166,N_6768);
or U8046 (N_8046,N_6796,N_7247);
nor U8047 (N_8047,N_7404,N_7388);
nand U8048 (N_8048,N_7143,N_7319);
and U8049 (N_8049,N_7171,N_7131);
or U8050 (N_8050,N_7338,N_7339);
nand U8051 (N_8051,N_6777,N_6974);
and U8052 (N_8052,N_6945,N_7240);
or U8053 (N_8053,N_7393,N_6803);
or U8054 (N_8054,N_7217,N_6946);
nand U8055 (N_8055,N_7066,N_7426);
or U8056 (N_8056,N_7156,N_7301);
xnor U8057 (N_8057,N_6961,N_7093);
nor U8058 (N_8058,N_7079,N_7414);
and U8059 (N_8059,N_7061,N_7436);
nor U8060 (N_8060,N_6987,N_7246);
or U8061 (N_8061,N_6836,N_6763);
nor U8062 (N_8062,N_7383,N_7499);
and U8063 (N_8063,N_6940,N_6834);
nor U8064 (N_8064,N_7247,N_7149);
xnor U8065 (N_8065,N_7421,N_7055);
nor U8066 (N_8066,N_7275,N_7184);
nor U8067 (N_8067,N_7089,N_7474);
xor U8068 (N_8068,N_6836,N_7162);
xnor U8069 (N_8069,N_7313,N_7261);
nand U8070 (N_8070,N_6802,N_7104);
nand U8071 (N_8071,N_6789,N_7081);
nand U8072 (N_8072,N_6765,N_7181);
nor U8073 (N_8073,N_6835,N_6824);
nor U8074 (N_8074,N_7202,N_7445);
nor U8075 (N_8075,N_7408,N_7151);
nor U8076 (N_8076,N_7092,N_7299);
nor U8077 (N_8077,N_6858,N_7280);
nor U8078 (N_8078,N_7087,N_7259);
nand U8079 (N_8079,N_7301,N_7115);
nor U8080 (N_8080,N_7400,N_7112);
or U8081 (N_8081,N_7092,N_6986);
nand U8082 (N_8082,N_7390,N_7357);
nor U8083 (N_8083,N_7455,N_6776);
xor U8084 (N_8084,N_7131,N_7496);
nand U8085 (N_8085,N_7334,N_7402);
nor U8086 (N_8086,N_6874,N_7037);
or U8087 (N_8087,N_6874,N_7029);
or U8088 (N_8088,N_6974,N_7475);
or U8089 (N_8089,N_7470,N_7230);
nor U8090 (N_8090,N_7180,N_7281);
nor U8091 (N_8091,N_7455,N_6794);
nand U8092 (N_8092,N_7138,N_7259);
or U8093 (N_8093,N_7031,N_6944);
nand U8094 (N_8094,N_6898,N_6952);
nor U8095 (N_8095,N_6795,N_7188);
and U8096 (N_8096,N_6967,N_7194);
nor U8097 (N_8097,N_6989,N_7447);
xnor U8098 (N_8098,N_6954,N_7003);
nor U8099 (N_8099,N_7328,N_6883);
nand U8100 (N_8100,N_7195,N_6854);
or U8101 (N_8101,N_6939,N_7337);
or U8102 (N_8102,N_7442,N_7100);
nor U8103 (N_8103,N_7440,N_7414);
nor U8104 (N_8104,N_7447,N_6826);
nand U8105 (N_8105,N_7451,N_6891);
or U8106 (N_8106,N_7029,N_6940);
nand U8107 (N_8107,N_7352,N_6973);
or U8108 (N_8108,N_6928,N_7422);
xor U8109 (N_8109,N_6890,N_7411);
xor U8110 (N_8110,N_7064,N_7456);
nand U8111 (N_8111,N_7483,N_6810);
nand U8112 (N_8112,N_6855,N_6878);
xor U8113 (N_8113,N_7379,N_7478);
nand U8114 (N_8114,N_6799,N_7202);
nand U8115 (N_8115,N_7005,N_7468);
or U8116 (N_8116,N_6877,N_6895);
nor U8117 (N_8117,N_6839,N_7493);
and U8118 (N_8118,N_7073,N_7445);
nor U8119 (N_8119,N_7246,N_7482);
or U8120 (N_8120,N_7161,N_7374);
nand U8121 (N_8121,N_6898,N_7362);
nand U8122 (N_8122,N_7247,N_6896);
nand U8123 (N_8123,N_7242,N_7389);
nand U8124 (N_8124,N_6966,N_6822);
or U8125 (N_8125,N_7491,N_7247);
nand U8126 (N_8126,N_7231,N_7200);
and U8127 (N_8127,N_7435,N_7063);
nor U8128 (N_8128,N_6961,N_6764);
or U8129 (N_8129,N_7322,N_7145);
nand U8130 (N_8130,N_7084,N_6770);
and U8131 (N_8131,N_6768,N_7175);
xnor U8132 (N_8132,N_7453,N_6946);
nor U8133 (N_8133,N_7299,N_7297);
nand U8134 (N_8134,N_6774,N_6763);
and U8135 (N_8135,N_7389,N_6902);
xor U8136 (N_8136,N_7362,N_7440);
and U8137 (N_8137,N_7445,N_7285);
or U8138 (N_8138,N_7161,N_7372);
or U8139 (N_8139,N_7106,N_7259);
or U8140 (N_8140,N_6772,N_6852);
xnor U8141 (N_8141,N_7493,N_7162);
or U8142 (N_8142,N_7218,N_6805);
and U8143 (N_8143,N_7207,N_7059);
nor U8144 (N_8144,N_7339,N_7275);
or U8145 (N_8145,N_7432,N_7364);
xnor U8146 (N_8146,N_7102,N_7375);
or U8147 (N_8147,N_7156,N_7476);
xor U8148 (N_8148,N_7178,N_7199);
or U8149 (N_8149,N_6843,N_7012);
nor U8150 (N_8150,N_7023,N_7220);
or U8151 (N_8151,N_7332,N_6823);
and U8152 (N_8152,N_6970,N_7185);
nor U8153 (N_8153,N_7237,N_7389);
nor U8154 (N_8154,N_7493,N_7498);
or U8155 (N_8155,N_7321,N_6876);
or U8156 (N_8156,N_7164,N_7215);
xnor U8157 (N_8157,N_7235,N_7084);
or U8158 (N_8158,N_7150,N_6810);
nor U8159 (N_8159,N_7090,N_6774);
and U8160 (N_8160,N_7382,N_7237);
or U8161 (N_8161,N_7230,N_7339);
nor U8162 (N_8162,N_6795,N_6988);
or U8163 (N_8163,N_7095,N_7442);
nor U8164 (N_8164,N_7290,N_7378);
nand U8165 (N_8165,N_7396,N_7490);
nor U8166 (N_8166,N_7300,N_7252);
nand U8167 (N_8167,N_7399,N_7170);
or U8168 (N_8168,N_7200,N_7215);
xor U8169 (N_8169,N_7170,N_6828);
and U8170 (N_8170,N_6917,N_6891);
xnor U8171 (N_8171,N_6887,N_6750);
and U8172 (N_8172,N_6879,N_6850);
xnor U8173 (N_8173,N_7483,N_7180);
and U8174 (N_8174,N_7208,N_7035);
and U8175 (N_8175,N_7022,N_6780);
nand U8176 (N_8176,N_6831,N_7146);
xor U8177 (N_8177,N_7474,N_6875);
nor U8178 (N_8178,N_7286,N_7310);
or U8179 (N_8179,N_6893,N_6817);
and U8180 (N_8180,N_7462,N_6942);
nand U8181 (N_8181,N_6875,N_7469);
and U8182 (N_8182,N_7085,N_6932);
nor U8183 (N_8183,N_6808,N_6847);
nor U8184 (N_8184,N_7138,N_6971);
and U8185 (N_8185,N_7076,N_6835);
and U8186 (N_8186,N_7175,N_7093);
or U8187 (N_8187,N_6916,N_7197);
xnor U8188 (N_8188,N_7180,N_7160);
and U8189 (N_8189,N_7244,N_7136);
or U8190 (N_8190,N_6938,N_7285);
xnor U8191 (N_8191,N_7185,N_7416);
nor U8192 (N_8192,N_7200,N_7468);
and U8193 (N_8193,N_7442,N_6953);
nor U8194 (N_8194,N_6763,N_6855);
and U8195 (N_8195,N_7440,N_6881);
xor U8196 (N_8196,N_7016,N_6915);
and U8197 (N_8197,N_7433,N_6789);
and U8198 (N_8198,N_6904,N_7481);
nand U8199 (N_8199,N_7440,N_7147);
nand U8200 (N_8200,N_7448,N_7142);
or U8201 (N_8201,N_6895,N_7383);
or U8202 (N_8202,N_7132,N_6952);
nand U8203 (N_8203,N_7498,N_6974);
nand U8204 (N_8204,N_7155,N_7326);
or U8205 (N_8205,N_6806,N_7351);
nor U8206 (N_8206,N_7318,N_7375);
and U8207 (N_8207,N_6896,N_7270);
nand U8208 (N_8208,N_7300,N_6814);
or U8209 (N_8209,N_7452,N_7344);
nand U8210 (N_8210,N_7370,N_7336);
and U8211 (N_8211,N_7397,N_7352);
xnor U8212 (N_8212,N_7139,N_6779);
xnor U8213 (N_8213,N_7066,N_6797);
xnor U8214 (N_8214,N_7305,N_7421);
and U8215 (N_8215,N_6928,N_7451);
xor U8216 (N_8216,N_7355,N_7095);
and U8217 (N_8217,N_7427,N_7249);
nor U8218 (N_8218,N_6873,N_7421);
nor U8219 (N_8219,N_6931,N_7004);
and U8220 (N_8220,N_7265,N_7152);
nand U8221 (N_8221,N_6755,N_7300);
and U8222 (N_8222,N_7066,N_7089);
xor U8223 (N_8223,N_7135,N_6814);
nand U8224 (N_8224,N_7029,N_7140);
nor U8225 (N_8225,N_6988,N_7194);
nand U8226 (N_8226,N_7215,N_6816);
xnor U8227 (N_8227,N_7081,N_6962);
and U8228 (N_8228,N_7416,N_6941);
nand U8229 (N_8229,N_7006,N_7222);
or U8230 (N_8230,N_7260,N_6975);
nor U8231 (N_8231,N_6853,N_7261);
and U8232 (N_8232,N_6791,N_6990);
or U8233 (N_8233,N_7374,N_6757);
nand U8234 (N_8234,N_6941,N_7403);
nand U8235 (N_8235,N_7353,N_7086);
and U8236 (N_8236,N_6785,N_6887);
or U8237 (N_8237,N_7138,N_7371);
nor U8238 (N_8238,N_6867,N_7214);
nand U8239 (N_8239,N_6902,N_7190);
xor U8240 (N_8240,N_7290,N_6781);
nor U8241 (N_8241,N_6826,N_6968);
and U8242 (N_8242,N_7326,N_6881);
or U8243 (N_8243,N_7303,N_7390);
nor U8244 (N_8244,N_7249,N_7033);
and U8245 (N_8245,N_7254,N_7216);
nand U8246 (N_8246,N_7222,N_6882);
and U8247 (N_8247,N_6878,N_7431);
or U8248 (N_8248,N_7195,N_7083);
and U8249 (N_8249,N_7285,N_6914);
nand U8250 (N_8250,N_7704,N_7567);
or U8251 (N_8251,N_8087,N_7714);
or U8252 (N_8252,N_7951,N_7796);
xor U8253 (N_8253,N_7591,N_8018);
nand U8254 (N_8254,N_7914,N_7845);
nor U8255 (N_8255,N_7729,N_7604);
nor U8256 (N_8256,N_8076,N_8025);
nand U8257 (N_8257,N_7755,N_7840);
and U8258 (N_8258,N_7507,N_8145);
and U8259 (N_8259,N_7803,N_8219);
nand U8260 (N_8260,N_7780,N_8075);
or U8261 (N_8261,N_8071,N_8080);
and U8262 (N_8262,N_7614,N_8051);
nor U8263 (N_8263,N_7898,N_8154);
xnor U8264 (N_8264,N_7957,N_7732);
and U8265 (N_8265,N_7717,N_8216);
xor U8266 (N_8266,N_7745,N_8188);
and U8267 (N_8267,N_8237,N_8163);
xnor U8268 (N_8268,N_7968,N_7777);
and U8269 (N_8269,N_8200,N_7514);
and U8270 (N_8270,N_7910,N_7743);
and U8271 (N_8271,N_7931,N_7685);
or U8272 (N_8272,N_7920,N_7683);
or U8273 (N_8273,N_7628,N_7657);
nand U8274 (N_8274,N_7859,N_7692);
and U8275 (N_8275,N_7577,N_8113);
or U8276 (N_8276,N_8125,N_7650);
nand U8277 (N_8277,N_7618,N_7593);
or U8278 (N_8278,N_7706,N_8088);
and U8279 (N_8279,N_7695,N_8225);
or U8280 (N_8280,N_7633,N_8244);
or U8281 (N_8281,N_7802,N_7876);
xnor U8282 (N_8282,N_8063,N_8126);
and U8283 (N_8283,N_7874,N_8109);
nand U8284 (N_8284,N_8082,N_8010);
nand U8285 (N_8285,N_8226,N_7986);
nand U8286 (N_8286,N_8050,N_7613);
or U8287 (N_8287,N_7915,N_8045);
xnor U8288 (N_8288,N_7554,N_7902);
and U8289 (N_8289,N_7697,N_7655);
nor U8290 (N_8290,N_8083,N_8224);
xor U8291 (N_8291,N_7636,N_8085);
or U8292 (N_8292,N_7763,N_8236);
xor U8293 (N_8293,N_7982,N_7983);
nand U8294 (N_8294,N_8141,N_7820);
nand U8295 (N_8295,N_7927,N_7976);
nor U8296 (N_8296,N_8049,N_7620);
or U8297 (N_8297,N_7853,N_7959);
nor U8298 (N_8298,N_7929,N_7900);
xor U8299 (N_8299,N_7998,N_8160);
nor U8300 (N_8300,N_7839,N_8165);
nand U8301 (N_8301,N_7922,N_8061);
xor U8302 (N_8302,N_7879,N_7975);
nor U8303 (N_8303,N_7793,N_8030);
nand U8304 (N_8304,N_7981,N_8022);
and U8305 (N_8305,N_8129,N_7863);
and U8306 (N_8306,N_7662,N_7587);
and U8307 (N_8307,N_7851,N_7737);
nand U8308 (N_8308,N_7778,N_8029);
xnor U8309 (N_8309,N_7792,N_7724);
or U8310 (N_8310,N_8211,N_7974);
nand U8311 (N_8311,N_8077,N_7795);
nand U8312 (N_8312,N_7945,N_7538);
and U8313 (N_8313,N_7557,N_7949);
nor U8314 (N_8314,N_8215,N_7622);
nand U8315 (N_8315,N_7516,N_7580);
and U8316 (N_8316,N_7666,N_7877);
nor U8317 (N_8317,N_7581,N_7635);
or U8318 (N_8318,N_7601,N_7800);
or U8319 (N_8319,N_7680,N_7590);
or U8320 (N_8320,N_7781,N_7540);
nor U8321 (N_8321,N_8228,N_8150);
xor U8322 (N_8322,N_8020,N_7947);
or U8323 (N_8323,N_8016,N_7543);
nor U8324 (N_8324,N_7659,N_7679);
nor U8325 (N_8325,N_7574,N_7824);
or U8326 (N_8326,N_8127,N_7977);
nor U8327 (N_8327,N_7999,N_8038);
xor U8328 (N_8328,N_7596,N_7742);
nor U8329 (N_8329,N_7885,N_7728);
nor U8330 (N_8330,N_7558,N_7735);
xor U8331 (N_8331,N_7653,N_8013);
and U8332 (N_8332,N_7531,N_7640);
and U8333 (N_8333,N_8248,N_7843);
nor U8334 (N_8334,N_8190,N_7855);
xnor U8335 (N_8335,N_8206,N_8173);
nor U8336 (N_8336,N_8197,N_7753);
and U8337 (N_8337,N_7571,N_7568);
xor U8338 (N_8338,N_8186,N_8170);
nand U8339 (N_8339,N_7869,N_8212);
nor U8340 (N_8340,N_7708,N_7705);
and U8341 (N_8341,N_7850,N_7806);
nand U8342 (N_8342,N_7858,N_7592);
nor U8343 (N_8343,N_8138,N_7736);
and U8344 (N_8344,N_7608,N_8181);
nand U8345 (N_8345,N_7688,N_8232);
xor U8346 (N_8346,N_7602,N_7825);
nor U8347 (N_8347,N_8246,N_7672);
nor U8348 (N_8348,N_8155,N_7619);
xor U8349 (N_8349,N_7721,N_8166);
nand U8350 (N_8350,N_7738,N_7921);
nand U8351 (N_8351,N_8169,N_7519);
or U8352 (N_8352,N_8217,N_8218);
xor U8353 (N_8353,N_7751,N_8073);
nor U8354 (N_8354,N_7617,N_7637);
and U8355 (N_8355,N_7675,N_7582);
nand U8356 (N_8356,N_7799,N_8157);
nand U8357 (N_8357,N_8052,N_7651);
nor U8358 (N_8358,N_7701,N_7849);
nor U8359 (N_8359,N_7993,N_8176);
and U8360 (N_8360,N_8098,N_8072);
and U8361 (N_8361,N_7754,N_7541);
nand U8362 (N_8362,N_8070,N_7854);
and U8363 (N_8363,N_8179,N_7757);
nor U8364 (N_8364,N_7684,N_7994);
or U8365 (N_8365,N_8012,N_7926);
and U8366 (N_8366,N_7860,N_8091);
and U8367 (N_8367,N_7572,N_7693);
and U8368 (N_8368,N_8021,N_7956);
or U8369 (N_8369,N_7527,N_7819);
and U8370 (N_8370,N_7932,N_7727);
or U8371 (N_8371,N_7969,N_8147);
xnor U8372 (N_8372,N_8005,N_7864);
or U8373 (N_8373,N_8123,N_8078);
or U8374 (N_8374,N_7747,N_8131);
or U8375 (N_8375,N_7689,N_7676);
xnor U8376 (N_8376,N_8065,N_7595);
nor U8377 (N_8377,N_7534,N_7775);
nor U8378 (N_8378,N_7783,N_7913);
nor U8379 (N_8379,N_7546,N_8238);
xor U8380 (N_8380,N_8067,N_8231);
or U8381 (N_8381,N_7875,N_8137);
nand U8382 (N_8382,N_7579,N_7548);
and U8383 (N_8383,N_8144,N_8112);
nor U8384 (N_8384,N_8039,N_8048);
nor U8385 (N_8385,N_8011,N_8132);
nor U8386 (N_8386,N_7646,N_8019);
or U8387 (N_8387,N_7690,N_7872);
nand U8388 (N_8388,N_8032,N_7607);
and U8389 (N_8389,N_7862,N_8036);
xnor U8390 (N_8390,N_7537,N_8079);
nand U8391 (N_8391,N_8159,N_7606);
xnor U8392 (N_8392,N_8153,N_8222);
xnor U8393 (N_8393,N_7817,N_8040);
xor U8394 (N_8394,N_7542,N_7699);
nor U8395 (N_8395,N_7642,N_7648);
or U8396 (N_8396,N_7517,N_8074);
or U8397 (N_8397,N_7535,N_7924);
or U8398 (N_8398,N_7609,N_7985);
xnor U8399 (N_8399,N_8142,N_7656);
nand U8400 (N_8400,N_7928,N_7630);
xor U8401 (N_8401,N_7887,N_7502);
nor U8402 (N_8402,N_8214,N_8046);
or U8403 (N_8403,N_7884,N_8026);
nand U8404 (N_8404,N_7955,N_7629);
nor U8405 (N_8405,N_7739,N_8041);
xor U8406 (N_8406,N_8174,N_8024);
or U8407 (N_8407,N_8033,N_8148);
or U8408 (N_8408,N_7812,N_7918);
and U8409 (N_8409,N_7823,N_8223);
and U8410 (N_8410,N_7847,N_7575);
or U8411 (N_8411,N_7828,N_8001);
nor U8412 (N_8412,N_7631,N_7809);
xor U8413 (N_8413,N_7661,N_7550);
nand U8414 (N_8414,N_7681,N_7936);
nand U8415 (N_8415,N_7668,N_8108);
or U8416 (N_8416,N_8162,N_7696);
nor U8417 (N_8417,N_8156,N_7573);
nor U8418 (N_8418,N_7944,N_7711);
nand U8419 (N_8419,N_8002,N_7776);
or U8420 (N_8420,N_7551,N_7643);
nor U8421 (N_8421,N_7505,N_7518);
nor U8422 (N_8422,N_7678,N_7821);
or U8423 (N_8423,N_8117,N_7564);
and U8424 (N_8424,N_7907,N_8086);
nand U8425 (N_8425,N_7987,N_7605);
or U8426 (N_8426,N_8007,N_7774);
nand U8427 (N_8427,N_7830,N_7810);
nor U8428 (N_8428,N_8208,N_7808);
or U8429 (N_8429,N_8135,N_8089);
or U8430 (N_8430,N_7912,N_7988);
nand U8431 (N_8431,N_7756,N_7698);
or U8432 (N_8432,N_7649,N_7647);
xnor U8433 (N_8433,N_7815,N_8053);
or U8434 (N_8434,N_7677,N_7515);
nand U8435 (N_8435,N_7664,N_7669);
nor U8436 (N_8436,N_7513,N_7552);
xnor U8437 (N_8437,N_8161,N_7788);
or U8438 (N_8438,N_7621,N_7765);
nand U8439 (N_8439,N_7952,N_7663);
and U8440 (N_8440,N_8171,N_8202);
and U8441 (N_8441,N_7733,N_8207);
nand U8442 (N_8442,N_7967,N_8104);
nand U8443 (N_8443,N_7510,N_7991);
nand U8444 (N_8444,N_8192,N_7521);
nand U8445 (N_8445,N_7566,N_8092);
xor U8446 (N_8446,N_7589,N_7771);
and U8447 (N_8447,N_7709,N_7893);
or U8448 (N_8448,N_7827,N_7962);
xor U8449 (N_8449,N_7719,N_8118);
or U8450 (N_8450,N_7897,N_7826);
nor U8451 (N_8451,N_7761,N_7702);
xnor U8452 (N_8452,N_7807,N_8189);
xnor U8453 (N_8453,N_7835,N_8119);
or U8454 (N_8454,N_8247,N_7509);
xor U8455 (N_8455,N_8064,N_8096);
nor U8456 (N_8456,N_8178,N_8114);
and U8457 (N_8457,N_8003,N_7950);
xor U8458 (N_8458,N_7730,N_7559);
xnor U8459 (N_8459,N_7805,N_8240);
xor U8460 (N_8460,N_8062,N_7822);
and U8461 (N_8461,N_8249,N_8035);
nor U8462 (N_8462,N_7954,N_8069);
and U8463 (N_8463,N_7856,N_7801);
xor U8464 (N_8464,N_7644,N_7645);
nand U8465 (N_8465,N_7995,N_7748);
and U8466 (N_8466,N_7996,N_7989);
nand U8467 (N_8467,N_7682,N_8205);
nor U8468 (N_8468,N_8037,N_7789);
nand U8469 (N_8469,N_7916,N_7848);
nand U8470 (N_8470,N_7966,N_7923);
nor U8471 (N_8471,N_8198,N_8124);
nor U8472 (N_8472,N_7578,N_7707);
and U8473 (N_8473,N_7686,N_7533);
nand U8474 (N_8474,N_7787,N_7597);
xor U8475 (N_8475,N_7726,N_7943);
xnor U8476 (N_8476,N_7615,N_7600);
nor U8477 (N_8477,N_7791,N_7846);
nor U8478 (N_8478,N_7536,N_8168);
or U8479 (N_8479,N_7710,N_8149);
or U8480 (N_8480,N_7794,N_7836);
xnor U8481 (N_8481,N_7798,N_8056);
nand U8482 (N_8482,N_7603,N_8044);
nand U8483 (N_8483,N_8047,N_7948);
nand U8484 (N_8484,N_8110,N_7674);
xor U8485 (N_8485,N_7837,N_8146);
or U8486 (N_8486,N_7569,N_7671);
nand U8487 (N_8487,N_7960,N_8060);
and U8488 (N_8488,N_7694,N_8006);
and U8489 (N_8489,N_8136,N_7971);
and U8490 (N_8490,N_8101,N_7841);
or U8491 (N_8491,N_8213,N_8008);
xnor U8492 (N_8492,N_7888,N_7861);
xor U8493 (N_8493,N_7834,N_8116);
or U8494 (N_8494,N_7886,N_7524);
nand U8495 (N_8495,N_7731,N_8175);
and U8496 (N_8496,N_8164,N_8133);
nor U8497 (N_8497,N_7520,N_7526);
nor U8498 (N_8498,N_8042,N_7811);
and U8499 (N_8499,N_8245,N_8107);
nand U8500 (N_8500,N_7766,N_7925);
xor U8501 (N_8501,N_7634,N_8199);
and U8502 (N_8502,N_7865,N_7549);
or U8503 (N_8503,N_7503,N_7984);
nand U8504 (N_8504,N_8182,N_7866);
nor U8505 (N_8505,N_8054,N_7561);
nor U8506 (N_8506,N_7940,N_8177);
and U8507 (N_8507,N_7570,N_7911);
nand U8508 (N_8508,N_8028,N_7703);
xor U8509 (N_8509,N_7530,N_7720);
nand U8510 (N_8510,N_7556,N_7616);
nor U8511 (N_8511,N_7673,N_7746);
and U8512 (N_8512,N_7980,N_7909);
nand U8513 (N_8513,N_7715,N_7942);
or U8514 (N_8514,N_7725,N_7588);
nand U8515 (N_8515,N_8220,N_7665);
and U8516 (N_8516,N_7716,N_8004);
nand U8517 (N_8517,N_8187,N_7818);
and U8518 (N_8518,N_7598,N_7785);
and U8519 (N_8519,N_8058,N_8140);
xnor U8520 (N_8520,N_8196,N_8242);
nand U8521 (N_8521,N_8128,N_7930);
xnor U8522 (N_8522,N_7599,N_8233);
and U8523 (N_8523,N_7937,N_8201);
xor U8524 (N_8524,N_7842,N_7623);
or U8525 (N_8525,N_7660,N_8120);
xor U8526 (N_8526,N_7508,N_7584);
xor U8527 (N_8527,N_7889,N_7953);
or U8528 (N_8528,N_7903,N_7905);
and U8529 (N_8529,N_7868,N_8094);
xnor U8530 (N_8530,N_7700,N_8130);
or U8531 (N_8531,N_7528,N_7760);
or U8532 (N_8532,N_7831,N_8000);
nand U8533 (N_8533,N_8167,N_8183);
and U8534 (N_8534,N_7563,N_8017);
nor U8535 (N_8535,N_8221,N_7654);
nor U8536 (N_8536,N_7857,N_7938);
nor U8537 (N_8537,N_7908,N_8015);
or U8538 (N_8538,N_8121,N_8227);
nor U8539 (N_8539,N_8234,N_8239);
and U8540 (N_8540,N_7667,N_7752);
xnor U8541 (N_8541,N_7741,N_7946);
or U8542 (N_8542,N_8151,N_7764);
and U8543 (N_8543,N_7973,N_7612);
nand U8544 (N_8544,N_8180,N_7941);
nor U8545 (N_8545,N_7734,N_7624);
nand U8546 (N_8546,N_7813,N_8152);
nor U8547 (N_8547,N_8134,N_7670);
nor U8548 (N_8548,N_7768,N_7500);
nor U8549 (N_8549,N_7544,N_8111);
or U8550 (N_8550,N_8185,N_7758);
or U8551 (N_8551,N_7687,N_8093);
or U8552 (N_8552,N_7770,N_8191);
nand U8553 (N_8553,N_8057,N_7625);
xnor U8554 (N_8554,N_7652,N_7904);
or U8555 (N_8555,N_8204,N_8209);
xnor U8556 (N_8556,N_7829,N_7786);
or U8557 (N_8557,N_8243,N_7529);
nand U8558 (N_8558,N_8158,N_7782);
or U8559 (N_8559,N_7565,N_7832);
nor U8560 (N_8560,N_7804,N_7779);
xnor U8561 (N_8561,N_7773,N_8014);
xor U8562 (N_8562,N_7626,N_8068);
or U8563 (N_8563,N_7744,N_7632);
nor U8564 (N_8564,N_7740,N_8027);
and U8565 (N_8565,N_8115,N_7772);
xnor U8566 (N_8566,N_8103,N_7992);
xnor U8567 (N_8567,N_7749,N_7833);
xnor U8568 (N_8568,N_7658,N_7852);
nor U8569 (N_8569,N_8172,N_8241);
xor U8570 (N_8570,N_8023,N_7990);
and U8571 (N_8571,N_8139,N_7867);
nand U8572 (N_8572,N_7769,N_7878);
xnor U8573 (N_8573,N_7545,N_7958);
xor U8574 (N_8574,N_8102,N_7501);
nand U8575 (N_8575,N_7762,N_7512);
or U8576 (N_8576,N_7504,N_7562);
xor U8577 (N_8577,N_7611,N_7891);
or U8578 (N_8578,N_8143,N_7641);
xnor U8579 (N_8579,N_8081,N_7934);
nor U8580 (N_8580,N_7979,N_7576);
nor U8581 (N_8581,N_7871,N_7759);
nand U8582 (N_8582,N_7881,N_8066);
or U8583 (N_8583,N_7713,N_7594);
xor U8584 (N_8584,N_8084,N_7712);
nand U8585 (N_8585,N_7880,N_7978);
nor U8586 (N_8586,N_8203,N_7718);
nor U8587 (N_8587,N_7522,N_7883);
nor U8588 (N_8588,N_7511,N_7899);
or U8589 (N_8589,N_7585,N_7906);
xnor U8590 (N_8590,N_7767,N_7939);
or U8591 (N_8591,N_8229,N_8195);
xor U8592 (N_8592,N_8100,N_7691);
and U8593 (N_8593,N_7814,N_7539);
and U8594 (N_8594,N_7532,N_7919);
and U8595 (N_8595,N_7997,N_8090);
nand U8596 (N_8596,N_7547,N_8194);
or U8597 (N_8597,N_7882,N_7722);
nor U8598 (N_8598,N_7555,N_7816);
nand U8599 (N_8599,N_7894,N_7586);
or U8600 (N_8600,N_8031,N_8099);
or U8601 (N_8601,N_7525,N_8193);
and U8602 (N_8602,N_8095,N_7784);
nor U8603 (N_8603,N_7964,N_7972);
nand U8604 (N_8604,N_7895,N_7935);
nor U8605 (N_8605,N_7750,N_7970);
nor U8606 (N_8606,N_8009,N_7965);
xnor U8607 (N_8607,N_8210,N_7892);
and U8608 (N_8608,N_7933,N_7553);
xnor U8609 (N_8609,N_8043,N_8230);
nand U8610 (N_8610,N_7506,N_7844);
or U8611 (N_8611,N_7838,N_7917);
nand U8612 (N_8612,N_7560,N_7639);
and U8613 (N_8613,N_8055,N_7901);
and U8614 (N_8614,N_8106,N_8122);
and U8615 (N_8615,N_8059,N_7963);
and U8616 (N_8616,N_7890,N_7790);
nor U8617 (N_8617,N_7896,N_7873);
nand U8618 (N_8618,N_7797,N_7961);
nand U8619 (N_8619,N_8034,N_7638);
xor U8620 (N_8620,N_7870,N_7583);
or U8621 (N_8621,N_8105,N_7523);
xor U8622 (N_8622,N_7610,N_8235);
nor U8623 (N_8623,N_8184,N_8097);
and U8624 (N_8624,N_7723,N_7627);
nand U8625 (N_8625,N_8237,N_7639);
xor U8626 (N_8626,N_7954,N_7698);
nand U8627 (N_8627,N_7894,N_7852);
nor U8628 (N_8628,N_8094,N_7867);
nor U8629 (N_8629,N_7504,N_8016);
nand U8630 (N_8630,N_8241,N_7792);
nor U8631 (N_8631,N_7542,N_7648);
and U8632 (N_8632,N_7870,N_7910);
or U8633 (N_8633,N_7998,N_8046);
nand U8634 (N_8634,N_7952,N_7584);
nor U8635 (N_8635,N_8229,N_8029);
xor U8636 (N_8636,N_7846,N_7873);
and U8637 (N_8637,N_8039,N_8224);
or U8638 (N_8638,N_7679,N_7921);
xnor U8639 (N_8639,N_7730,N_7770);
or U8640 (N_8640,N_8003,N_8155);
or U8641 (N_8641,N_7618,N_7608);
xor U8642 (N_8642,N_8022,N_7687);
xnor U8643 (N_8643,N_8095,N_7504);
nor U8644 (N_8644,N_8053,N_7716);
or U8645 (N_8645,N_7985,N_7613);
and U8646 (N_8646,N_7970,N_7942);
nand U8647 (N_8647,N_8226,N_7751);
nor U8648 (N_8648,N_7586,N_8032);
or U8649 (N_8649,N_7508,N_7520);
xnor U8650 (N_8650,N_8242,N_7503);
or U8651 (N_8651,N_7692,N_7759);
and U8652 (N_8652,N_8001,N_8167);
nor U8653 (N_8653,N_7949,N_7729);
nor U8654 (N_8654,N_7839,N_7656);
nor U8655 (N_8655,N_7547,N_8085);
or U8656 (N_8656,N_8017,N_8045);
nand U8657 (N_8657,N_8137,N_7955);
and U8658 (N_8658,N_7511,N_7702);
nor U8659 (N_8659,N_7720,N_8143);
or U8660 (N_8660,N_7717,N_8106);
and U8661 (N_8661,N_8159,N_8043);
nand U8662 (N_8662,N_8177,N_7738);
and U8663 (N_8663,N_8206,N_8119);
nand U8664 (N_8664,N_7557,N_8171);
or U8665 (N_8665,N_7878,N_7784);
or U8666 (N_8666,N_7740,N_7845);
nor U8667 (N_8667,N_7943,N_7938);
nand U8668 (N_8668,N_7700,N_8100);
nand U8669 (N_8669,N_7997,N_7966);
nand U8670 (N_8670,N_7848,N_8246);
nor U8671 (N_8671,N_8073,N_7879);
and U8672 (N_8672,N_7557,N_7980);
xor U8673 (N_8673,N_7901,N_7926);
and U8674 (N_8674,N_7953,N_7564);
xnor U8675 (N_8675,N_8247,N_7677);
and U8676 (N_8676,N_7744,N_8156);
nor U8677 (N_8677,N_8070,N_8171);
nand U8678 (N_8678,N_8100,N_8024);
or U8679 (N_8679,N_7724,N_7715);
or U8680 (N_8680,N_8239,N_8018);
and U8681 (N_8681,N_8126,N_8101);
nor U8682 (N_8682,N_8083,N_8112);
nor U8683 (N_8683,N_8169,N_7528);
nor U8684 (N_8684,N_7512,N_7952);
nor U8685 (N_8685,N_7862,N_7822);
xnor U8686 (N_8686,N_8015,N_7891);
and U8687 (N_8687,N_7740,N_7671);
nand U8688 (N_8688,N_7575,N_7688);
nand U8689 (N_8689,N_7759,N_8091);
or U8690 (N_8690,N_8189,N_7612);
xor U8691 (N_8691,N_8133,N_8192);
nor U8692 (N_8692,N_7855,N_7575);
xnor U8693 (N_8693,N_8080,N_7930);
nor U8694 (N_8694,N_7546,N_7554);
nand U8695 (N_8695,N_7571,N_7537);
nor U8696 (N_8696,N_7566,N_8200);
xnor U8697 (N_8697,N_7966,N_7850);
nor U8698 (N_8698,N_7640,N_7748);
nand U8699 (N_8699,N_7757,N_7962);
and U8700 (N_8700,N_7696,N_7573);
nand U8701 (N_8701,N_7891,N_7857);
or U8702 (N_8702,N_7611,N_8006);
and U8703 (N_8703,N_7726,N_8052);
and U8704 (N_8704,N_7737,N_7776);
and U8705 (N_8705,N_7765,N_7655);
and U8706 (N_8706,N_8006,N_8030);
or U8707 (N_8707,N_7560,N_7932);
nor U8708 (N_8708,N_8184,N_7783);
and U8709 (N_8709,N_7695,N_7909);
and U8710 (N_8710,N_7578,N_7949);
xor U8711 (N_8711,N_7942,N_7847);
nand U8712 (N_8712,N_7883,N_7776);
xnor U8713 (N_8713,N_7546,N_8000);
or U8714 (N_8714,N_8216,N_7750);
and U8715 (N_8715,N_7918,N_7919);
nor U8716 (N_8716,N_7657,N_7613);
nor U8717 (N_8717,N_7896,N_7544);
nor U8718 (N_8718,N_7802,N_7871);
nand U8719 (N_8719,N_7662,N_7996);
nor U8720 (N_8720,N_7910,N_7895);
xor U8721 (N_8721,N_8061,N_7510);
and U8722 (N_8722,N_7576,N_7713);
xnor U8723 (N_8723,N_7799,N_8086);
nand U8724 (N_8724,N_8114,N_7869);
nand U8725 (N_8725,N_8192,N_8037);
xnor U8726 (N_8726,N_7746,N_7569);
nand U8727 (N_8727,N_8012,N_7603);
and U8728 (N_8728,N_7963,N_7522);
or U8729 (N_8729,N_8157,N_7877);
nor U8730 (N_8730,N_7930,N_8163);
and U8731 (N_8731,N_7725,N_7916);
or U8732 (N_8732,N_7876,N_8187);
nand U8733 (N_8733,N_7902,N_8229);
nand U8734 (N_8734,N_7503,N_7916);
xor U8735 (N_8735,N_7642,N_7633);
xnor U8736 (N_8736,N_8248,N_7951);
nor U8737 (N_8737,N_7903,N_7998);
xor U8738 (N_8738,N_8214,N_7805);
nand U8739 (N_8739,N_7500,N_7846);
xnor U8740 (N_8740,N_7753,N_7876);
and U8741 (N_8741,N_8148,N_7622);
xor U8742 (N_8742,N_8079,N_8103);
xor U8743 (N_8743,N_8117,N_7857);
or U8744 (N_8744,N_7950,N_8028);
nor U8745 (N_8745,N_7693,N_8165);
xor U8746 (N_8746,N_7635,N_7906);
nand U8747 (N_8747,N_7596,N_7781);
nor U8748 (N_8748,N_7810,N_7550);
and U8749 (N_8749,N_7629,N_8114);
nand U8750 (N_8750,N_8106,N_8166);
nor U8751 (N_8751,N_7978,N_7549);
nand U8752 (N_8752,N_7989,N_7562);
nand U8753 (N_8753,N_7508,N_7749);
and U8754 (N_8754,N_8123,N_8042);
nor U8755 (N_8755,N_7983,N_7665);
and U8756 (N_8756,N_8100,N_7605);
xnor U8757 (N_8757,N_7887,N_7787);
or U8758 (N_8758,N_7998,N_7906);
nand U8759 (N_8759,N_8000,N_7955);
nand U8760 (N_8760,N_7972,N_8227);
nor U8761 (N_8761,N_7963,N_7773);
nand U8762 (N_8762,N_7772,N_8090);
nor U8763 (N_8763,N_8159,N_7855);
or U8764 (N_8764,N_7529,N_7511);
nand U8765 (N_8765,N_7768,N_7633);
and U8766 (N_8766,N_7971,N_7934);
or U8767 (N_8767,N_7919,N_8091);
nor U8768 (N_8768,N_8124,N_8150);
nor U8769 (N_8769,N_8018,N_7887);
nand U8770 (N_8770,N_8008,N_7853);
xnor U8771 (N_8771,N_7852,N_7646);
or U8772 (N_8772,N_7597,N_8162);
nand U8773 (N_8773,N_7750,N_7668);
and U8774 (N_8774,N_7524,N_7617);
or U8775 (N_8775,N_7959,N_7556);
xor U8776 (N_8776,N_7807,N_7593);
nand U8777 (N_8777,N_7738,N_7672);
xnor U8778 (N_8778,N_7888,N_7614);
and U8779 (N_8779,N_8111,N_8148);
xnor U8780 (N_8780,N_8099,N_7508);
and U8781 (N_8781,N_7805,N_7969);
or U8782 (N_8782,N_7808,N_7894);
xnor U8783 (N_8783,N_7927,N_7999);
and U8784 (N_8784,N_7829,N_8007);
nand U8785 (N_8785,N_7786,N_8071);
nand U8786 (N_8786,N_7986,N_7588);
or U8787 (N_8787,N_7952,N_8188);
and U8788 (N_8788,N_7517,N_8007);
nor U8789 (N_8789,N_7926,N_7516);
nand U8790 (N_8790,N_7848,N_8191);
or U8791 (N_8791,N_7799,N_7907);
and U8792 (N_8792,N_7989,N_8101);
nand U8793 (N_8793,N_7690,N_8032);
or U8794 (N_8794,N_7894,N_7953);
xor U8795 (N_8795,N_8151,N_8216);
and U8796 (N_8796,N_7508,N_7629);
or U8797 (N_8797,N_8170,N_7792);
xor U8798 (N_8798,N_7807,N_8111);
and U8799 (N_8799,N_7546,N_7869);
nor U8800 (N_8800,N_7515,N_7620);
nor U8801 (N_8801,N_7604,N_7759);
nand U8802 (N_8802,N_7760,N_7693);
nand U8803 (N_8803,N_7766,N_8246);
nand U8804 (N_8804,N_7809,N_7586);
or U8805 (N_8805,N_7659,N_8057);
or U8806 (N_8806,N_8098,N_8212);
nand U8807 (N_8807,N_8011,N_8110);
xnor U8808 (N_8808,N_7991,N_7695);
nand U8809 (N_8809,N_7755,N_7681);
and U8810 (N_8810,N_8193,N_7890);
nor U8811 (N_8811,N_7894,N_7960);
xnor U8812 (N_8812,N_8051,N_7671);
nand U8813 (N_8813,N_8051,N_7531);
xnor U8814 (N_8814,N_8070,N_7957);
xnor U8815 (N_8815,N_7632,N_8157);
or U8816 (N_8816,N_7683,N_7881);
nor U8817 (N_8817,N_7902,N_7518);
or U8818 (N_8818,N_7698,N_7782);
and U8819 (N_8819,N_7573,N_7946);
nand U8820 (N_8820,N_7614,N_7952);
nor U8821 (N_8821,N_7892,N_8038);
and U8822 (N_8822,N_7522,N_7692);
and U8823 (N_8823,N_8075,N_7513);
nand U8824 (N_8824,N_7899,N_7500);
nand U8825 (N_8825,N_8060,N_8208);
xor U8826 (N_8826,N_8028,N_8008);
xnor U8827 (N_8827,N_7922,N_7605);
or U8828 (N_8828,N_7540,N_8159);
nor U8829 (N_8829,N_7969,N_7800);
and U8830 (N_8830,N_7960,N_7758);
or U8831 (N_8831,N_7961,N_8104);
or U8832 (N_8832,N_8045,N_7756);
nand U8833 (N_8833,N_8103,N_7939);
or U8834 (N_8834,N_7521,N_7702);
and U8835 (N_8835,N_7845,N_8137);
xor U8836 (N_8836,N_7928,N_8103);
and U8837 (N_8837,N_7528,N_8231);
nand U8838 (N_8838,N_7884,N_7656);
and U8839 (N_8839,N_7686,N_7783);
or U8840 (N_8840,N_7658,N_7866);
nor U8841 (N_8841,N_8119,N_7940);
nand U8842 (N_8842,N_7933,N_7711);
nand U8843 (N_8843,N_7942,N_7976);
and U8844 (N_8844,N_8218,N_7555);
nor U8845 (N_8845,N_7608,N_7535);
xnor U8846 (N_8846,N_8086,N_8109);
nor U8847 (N_8847,N_7542,N_8018);
xnor U8848 (N_8848,N_8093,N_8073);
nor U8849 (N_8849,N_7976,N_7645);
nand U8850 (N_8850,N_8236,N_7955);
nor U8851 (N_8851,N_7904,N_7733);
nand U8852 (N_8852,N_7876,N_7941);
xnor U8853 (N_8853,N_7740,N_7820);
xor U8854 (N_8854,N_7693,N_8157);
nand U8855 (N_8855,N_8238,N_7558);
nor U8856 (N_8856,N_7673,N_7901);
and U8857 (N_8857,N_7719,N_7687);
and U8858 (N_8858,N_8060,N_8143);
nand U8859 (N_8859,N_8146,N_8238);
nor U8860 (N_8860,N_7630,N_8204);
xnor U8861 (N_8861,N_8027,N_7987);
or U8862 (N_8862,N_7872,N_8203);
nor U8863 (N_8863,N_7934,N_8018);
and U8864 (N_8864,N_8227,N_7980);
or U8865 (N_8865,N_7637,N_7836);
or U8866 (N_8866,N_8009,N_8087);
or U8867 (N_8867,N_7804,N_8177);
or U8868 (N_8868,N_7673,N_7818);
nor U8869 (N_8869,N_7874,N_7744);
and U8870 (N_8870,N_7886,N_7989);
or U8871 (N_8871,N_7680,N_7809);
nand U8872 (N_8872,N_7868,N_7568);
or U8873 (N_8873,N_8038,N_7857);
xnor U8874 (N_8874,N_7779,N_8106);
and U8875 (N_8875,N_8201,N_7718);
or U8876 (N_8876,N_7997,N_7818);
nor U8877 (N_8877,N_7686,N_7827);
nor U8878 (N_8878,N_7782,N_7692);
nand U8879 (N_8879,N_8034,N_7814);
and U8880 (N_8880,N_7950,N_7835);
nor U8881 (N_8881,N_8149,N_8229);
nand U8882 (N_8882,N_7684,N_8196);
or U8883 (N_8883,N_7963,N_8198);
nand U8884 (N_8884,N_8099,N_8119);
or U8885 (N_8885,N_7584,N_7941);
and U8886 (N_8886,N_8132,N_8128);
or U8887 (N_8887,N_7592,N_8097);
xor U8888 (N_8888,N_7910,N_7542);
or U8889 (N_8889,N_7565,N_7908);
and U8890 (N_8890,N_8028,N_8153);
xnor U8891 (N_8891,N_8155,N_7584);
or U8892 (N_8892,N_7665,N_7688);
nand U8893 (N_8893,N_7530,N_8183);
xor U8894 (N_8894,N_7850,N_7843);
nand U8895 (N_8895,N_7771,N_7720);
xnor U8896 (N_8896,N_7985,N_8035);
or U8897 (N_8897,N_8130,N_8043);
and U8898 (N_8898,N_8116,N_7819);
or U8899 (N_8899,N_8085,N_7891);
xnor U8900 (N_8900,N_7768,N_7588);
and U8901 (N_8901,N_8190,N_7589);
nand U8902 (N_8902,N_7961,N_7742);
and U8903 (N_8903,N_7644,N_7923);
or U8904 (N_8904,N_7573,N_7897);
xor U8905 (N_8905,N_8102,N_8210);
and U8906 (N_8906,N_8120,N_7994);
or U8907 (N_8907,N_7822,N_7652);
nor U8908 (N_8908,N_8021,N_8068);
nand U8909 (N_8909,N_8035,N_7969);
and U8910 (N_8910,N_7869,N_7760);
nand U8911 (N_8911,N_7903,N_7964);
nor U8912 (N_8912,N_7784,N_7504);
xnor U8913 (N_8913,N_7943,N_8064);
and U8914 (N_8914,N_8175,N_7715);
nor U8915 (N_8915,N_8149,N_7773);
xnor U8916 (N_8916,N_8216,N_7850);
or U8917 (N_8917,N_7917,N_8027);
and U8918 (N_8918,N_7528,N_7794);
xnor U8919 (N_8919,N_7811,N_7690);
and U8920 (N_8920,N_7737,N_8208);
nand U8921 (N_8921,N_8212,N_7780);
xor U8922 (N_8922,N_7710,N_8192);
and U8923 (N_8923,N_7687,N_7663);
nor U8924 (N_8924,N_7571,N_7513);
nand U8925 (N_8925,N_7860,N_7683);
nand U8926 (N_8926,N_8178,N_8011);
nor U8927 (N_8927,N_7750,N_8215);
and U8928 (N_8928,N_7616,N_8016);
nand U8929 (N_8929,N_8228,N_8005);
nor U8930 (N_8930,N_7929,N_7976);
and U8931 (N_8931,N_8210,N_7742);
nor U8932 (N_8932,N_7890,N_7784);
nor U8933 (N_8933,N_7927,N_8208);
or U8934 (N_8934,N_8068,N_7674);
nand U8935 (N_8935,N_8038,N_7602);
xor U8936 (N_8936,N_7804,N_8010);
nor U8937 (N_8937,N_7531,N_7858);
xnor U8938 (N_8938,N_7898,N_7615);
xnor U8939 (N_8939,N_8138,N_7866);
nand U8940 (N_8940,N_8115,N_7805);
xnor U8941 (N_8941,N_7833,N_8117);
and U8942 (N_8942,N_7600,N_7667);
and U8943 (N_8943,N_7758,N_8065);
nand U8944 (N_8944,N_7543,N_7709);
xnor U8945 (N_8945,N_8229,N_8147);
xnor U8946 (N_8946,N_7561,N_7858);
or U8947 (N_8947,N_7984,N_8243);
xnor U8948 (N_8948,N_7577,N_7583);
and U8949 (N_8949,N_7852,N_7781);
or U8950 (N_8950,N_7989,N_7619);
nand U8951 (N_8951,N_7527,N_8026);
or U8952 (N_8952,N_7656,N_7525);
or U8953 (N_8953,N_8070,N_7921);
or U8954 (N_8954,N_7848,N_7607);
nor U8955 (N_8955,N_7720,N_8097);
xor U8956 (N_8956,N_8026,N_7875);
xor U8957 (N_8957,N_8189,N_7913);
nor U8958 (N_8958,N_8091,N_7933);
nor U8959 (N_8959,N_7612,N_8231);
or U8960 (N_8960,N_8063,N_7576);
nand U8961 (N_8961,N_8190,N_7510);
nor U8962 (N_8962,N_7746,N_7531);
nand U8963 (N_8963,N_7878,N_7892);
and U8964 (N_8964,N_7976,N_8093);
xor U8965 (N_8965,N_7943,N_7680);
nand U8966 (N_8966,N_8242,N_7562);
nand U8967 (N_8967,N_8236,N_8168);
nand U8968 (N_8968,N_8137,N_8153);
and U8969 (N_8969,N_8184,N_7634);
and U8970 (N_8970,N_7608,N_7773);
or U8971 (N_8971,N_7930,N_7970);
xor U8972 (N_8972,N_8094,N_7511);
or U8973 (N_8973,N_7542,N_7797);
xnor U8974 (N_8974,N_7884,N_7981);
nor U8975 (N_8975,N_7847,N_8010);
nor U8976 (N_8976,N_7844,N_8095);
xor U8977 (N_8977,N_8073,N_7766);
nand U8978 (N_8978,N_7890,N_8247);
xnor U8979 (N_8979,N_7556,N_7835);
or U8980 (N_8980,N_7670,N_7688);
and U8981 (N_8981,N_7947,N_7710);
nand U8982 (N_8982,N_8077,N_7845);
and U8983 (N_8983,N_8177,N_7883);
xor U8984 (N_8984,N_7945,N_8058);
nand U8985 (N_8985,N_8179,N_7574);
xnor U8986 (N_8986,N_7920,N_7971);
nand U8987 (N_8987,N_8241,N_7892);
nor U8988 (N_8988,N_7638,N_8182);
nor U8989 (N_8989,N_7611,N_7772);
xor U8990 (N_8990,N_7934,N_7883);
or U8991 (N_8991,N_7510,N_7664);
nand U8992 (N_8992,N_7728,N_7947);
and U8993 (N_8993,N_8190,N_7963);
xnor U8994 (N_8994,N_7724,N_8112);
and U8995 (N_8995,N_7662,N_8095);
nand U8996 (N_8996,N_7809,N_8219);
nor U8997 (N_8997,N_7731,N_7781);
xnor U8998 (N_8998,N_8103,N_8205);
nand U8999 (N_8999,N_8131,N_7554);
nor U9000 (N_9000,N_8468,N_8741);
nand U9001 (N_9001,N_8650,N_8317);
and U9002 (N_9002,N_8471,N_8911);
or U9003 (N_9003,N_8441,N_8601);
or U9004 (N_9004,N_8591,N_8937);
and U9005 (N_9005,N_8993,N_8967);
nand U9006 (N_9006,N_8836,N_8657);
nand U9007 (N_9007,N_8602,N_8496);
nand U9008 (N_9008,N_8369,N_8400);
and U9009 (N_9009,N_8992,N_8768);
and U9010 (N_9010,N_8887,N_8856);
or U9011 (N_9011,N_8345,N_8855);
nor U9012 (N_9012,N_8448,N_8430);
or U9013 (N_9013,N_8339,N_8793);
or U9014 (N_9014,N_8579,N_8853);
and U9015 (N_9015,N_8407,N_8551);
nor U9016 (N_9016,N_8279,N_8909);
and U9017 (N_9017,N_8882,N_8832);
or U9018 (N_9018,N_8978,N_8559);
nand U9019 (N_9019,N_8338,N_8402);
nand U9020 (N_9020,N_8800,N_8418);
nand U9021 (N_9021,N_8844,N_8865);
or U9022 (N_9022,N_8944,N_8336);
nor U9023 (N_9023,N_8974,N_8361);
nand U9024 (N_9024,N_8305,N_8782);
xnor U9025 (N_9025,N_8296,N_8850);
nor U9026 (N_9026,N_8566,N_8811);
nor U9027 (N_9027,N_8473,N_8946);
xor U9028 (N_9028,N_8633,N_8900);
xor U9029 (N_9029,N_8731,N_8714);
and U9030 (N_9030,N_8669,N_8392);
nand U9031 (N_9031,N_8763,N_8991);
nand U9032 (N_9032,N_8627,N_8895);
xnor U9033 (N_9033,N_8482,N_8457);
and U9034 (N_9034,N_8507,N_8340);
and U9035 (N_9035,N_8437,N_8569);
nand U9036 (N_9036,N_8480,N_8863);
or U9037 (N_9037,N_8784,N_8474);
and U9038 (N_9038,N_8764,N_8631);
nor U9039 (N_9039,N_8302,N_8290);
and U9040 (N_9040,N_8554,N_8977);
nand U9041 (N_9041,N_8729,N_8349);
nand U9042 (N_9042,N_8427,N_8259);
or U9043 (N_9043,N_8924,N_8861);
nor U9044 (N_9044,N_8699,N_8723);
xnor U9045 (N_9045,N_8454,N_8726);
or U9046 (N_9046,N_8623,N_8772);
or U9047 (N_9047,N_8287,N_8923);
or U9048 (N_9048,N_8616,N_8310);
or U9049 (N_9049,N_8817,N_8385);
xor U9050 (N_9050,N_8269,N_8506);
nor U9051 (N_9051,N_8486,N_8769);
and U9052 (N_9052,N_8845,N_8456);
xnor U9053 (N_9053,N_8278,N_8268);
nand U9054 (N_9054,N_8393,N_8495);
and U9055 (N_9055,N_8678,N_8801);
nor U9056 (N_9056,N_8711,N_8710);
xnor U9057 (N_9057,N_8491,N_8894);
xor U9058 (N_9058,N_8692,N_8460);
nor U9059 (N_9059,N_8819,N_8914);
or U9060 (N_9060,N_8280,N_8462);
and U9061 (N_9061,N_8775,N_8813);
nor U9062 (N_9062,N_8690,N_8922);
and U9063 (N_9063,N_8368,N_8553);
and U9064 (N_9064,N_8286,N_8440);
xor U9065 (N_9065,N_8847,N_8805);
nor U9066 (N_9066,N_8425,N_8382);
and U9067 (N_9067,N_8572,N_8334);
xor U9068 (N_9068,N_8527,N_8637);
and U9069 (N_9069,N_8646,N_8372);
nand U9070 (N_9070,N_8258,N_8335);
xor U9071 (N_9071,N_8304,N_8717);
or U9072 (N_9072,N_8774,N_8919);
nor U9073 (N_9073,N_8276,N_8724);
and U9074 (N_9074,N_8698,N_8595);
and U9075 (N_9075,N_8549,N_8423);
nand U9076 (N_9076,N_8376,N_8373);
nand U9077 (N_9077,N_8634,N_8940);
or U9078 (N_9078,N_8799,N_8896);
xnor U9079 (N_9079,N_8500,N_8614);
and U9080 (N_9080,N_8628,N_8556);
xnor U9081 (N_9081,N_8792,N_8300);
xor U9082 (N_9082,N_8464,N_8785);
nand U9083 (N_9083,N_8539,N_8434);
and U9084 (N_9084,N_8273,N_8484);
or U9085 (N_9085,N_8607,N_8687);
xnor U9086 (N_9086,N_8585,N_8688);
xor U9087 (N_9087,N_8933,N_8830);
nor U9088 (N_9088,N_8884,N_8860);
xor U9089 (N_9089,N_8673,N_8907);
nand U9090 (N_9090,N_8390,N_8550);
xnor U9091 (N_9091,N_8446,N_8790);
nor U9092 (N_9092,N_8416,N_8583);
nor U9093 (N_9093,N_8435,N_8684);
nand U9094 (N_9094,N_8875,N_8449);
xnor U9095 (N_9095,N_8864,N_8939);
xor U9096 (N_9096,N_8765,N_8750);
nor U9097 (N_9097,N_8325,N_8695);
nor U9098 (N_9098,N_8727,N_8777);
or U9099 (N_9099,N_8709,N_8834);
nand U9100 (N_9100,N_8309,N_8512);
nor U9101 (N_9101,N_8315,N_8851);
and U9102 (N_9102,N_8251,N_8472);
nand U9103 (N_9103,N_8580,N_8959);
or U9104 (N_9104,N_8685,N_8270);
or U9105 (N_9105,N_8635,N_8739);
xor U9106 (N_9106,N_8523,N_8327);
nor U9107 (N_9107,N_8271,N_8351);
and U9108 (N_9108,N_8973,N_8526);
nor U9109 (N_9109,N_8771,N_8916);
nand U9110 (N_9110,N_8942,N_8363);
nand U9111 (N_9111,N_8749,N_8455);
or U9112 (N_9112,N_8333,N_8878);
nand U9113 (N_9113,N_8778,N_8316);
nor U9114 (N_9114,N_8516,N_8356);
or U9115 (N_9115,N_8615,N_8510);
xor U9116 (N_9116,N_8406,N_8371);
nor U9117 (N_9117,N_8467,N_8842);
nand U9118 (N_9118,N_8822,N_8901);
or U9119 (N_9119,N_8643,N_8653);
nand U9120 (N_9120,N_8783,N_8951);
and U9121 (N_9121,N_8612,N_8529);
nand U9122 (N_9122,N_8862,N_8701);
xnor U9123 (N_9123,N_8394,N_8613);
or U9124 (N_9124,N_8370,N_8693);
nor U9125 (N_9125,N_8537,N_8250);
nor U9126 (N_9126,N_8330,N_8540);
and U9127 (N_9127,N_8401,N_8292);
xor U9128 (N_9128,N_8337,N_8444);
or U9129 (N_9129,N_8508,N_8586);
nand U9130 (N_9130,N_8744,N_8735);
or U9131 (N_9131,N_8621,N_8934);
xnor U9132 (N_9132,N_8360,N_8533);
and U9133 (N_9133,N_8986,N_8918);
nor U9134 (N_9134,N_8912,N_8737);
and U9135 (N_9135,N_8501,N_8658);
or U9136 (N_9136,N_8534,N_8255);
nor U9137 (N_9137,N_8410,N_8902);
nor U9138 (N_9138,N_8736,N_8985);
nor U9139 (N_9139,N_8903,N_8756);
or U9140 (N_9140,N_8547,N_8530);
xor U9141 (N_9141,N_8285,N_8590);
or U9142 (N_9142,N_8866,N_8935);
and U9143 (N_9143,N_8654,N_8624);
nor U9144 (N_9144,N_8667,N_8424);
and U9145 (N_9145,N_8931,N_8880);
nand U9146 (N_9146,N_8640,N_8487);
xnor U9147 (N_9147,N_8575,N_8818);
or U9148 (N_9148,N_8995,N_8346);
xnor U9149 (N_9149,N_8892,N_8314);
or U9150 (N_9150,N_8522,N_8889);
and U9151 (N_9151,N_8788,N_8984);
or U9152 (N_9152,N_8702,N_8719);
or U9153 (N_9153,N_8609,N_8926);
nand U9154 (N_9154,N_8518,N_8732);
nor U9155 (N_9155,N_8383,N_8299);
nand U9156 (N_9156,N_8676,N_8535);
nor U9157 (N_9157,N_8321,N_8704);
nor U9158 (N_9158,N_8821,N_8715);
nand U9159 (N_9159,N_8770,N_8544);
nor U9160 (N_9160,N_8284,N_8319);
and U9161 (N_9161,N_8531,N_8897);
xor U9162 (N_9162,N_8600,N_8388);
and U9163 (N_9163,N_8642,N_8979);
or U9164 (N_9164,N_8998,N_8291);
nor U9165 (N_9165,N_8422,N_8665);
nand U9166 (N_9166,N_8358,N_8447);
nor U9167 (N_9167,N_8891,N_8681);
and U9168 (N_9168,N_8964,N_8953);
xor U9169 (N_9169,N_8324,N_8656);
nor U9170 (N_9170,N_8272,N_8611);
nand U9171 (N_9171,N_8872,N_8606);
nand U9172 (N_9172,N_8721,N_8488);
or U9173 (N_9173,N_8955,N_8660);
xor U9174 (N_9174,N_8519,N_8502);
nand U9175 (N_9175,N_8812,N_8396);
nor U9176 (N_9176,N_8451,N_8908);
nand U9177 (N_9177,N_8283,N_8563);
xor U9178 (N_9178,N_8787,N_8414);
xnor U9179 (N_9179,N_8608,N_8747);
and U9180 (N_9180,N_8683,N_8515);
or U9181 (N_9181,N_8405,N_8970);
nor U9182 (N_9182,N_8824,N_8814);
or U9183 (N_9183,N_8420,N_8320);
nand U9184 (N_9184,N_8429,N_8589);
and U9185 (N_9185,N_8492,N_8753);
nand U9186 (N_9186,N_8620,N_8742);
nor U9187 (N_9187,N_8776,N_8362);
xor U9188 (N_9188,N_8876,N_8906);
or U9189 (N_9189,N_8466,N_8869);
nor U9190 (N_9190,N_8536,N_8432);
and U9191 (N_9191,N_8988,N_8649);
nand U9192 (N_9192,N_8905,N_8528);
or U9193 (N_9193,N_8622,N_8837);
or U9194 (N_9194,N_8762,N_8825);
and U9195 (N_9195,N_8381,N_8560);
or U9196 (N_9196,N_8707,N_8961);
nand U9197 (N_9197,N_8791,N_8936);
or U9198 (N_9198,N_8674,N_8720);
xnor U9199 (N_9199,N_8538,N_8810);
nand U9200 (N_9200,N_8943,N_8399);
nand U9201 (N_9201,N_8266,N_8679);
xnor U9202 (N_9202,N_8950,N_8443);
xor U9203 (N_9203,N_8476,N_8716);
nand U9204 (N_9204,N_8689,N_8697);
nand U9205 (N_9205,N_8713,N_8925);
or U9206 (N_9206,N_8603,N_8311);
and U9207 (N_9207,N_8890,N_8982);
nor U9208 (N_9208,N_8588,N_8694);
nor U9209 (N_9209,N_8461,N_8648);
and U9210 (N_9210,N_8879,N_8593);
or U9211 (N_9211,N_8328,N_8675);
xnor U9212 (N_9212,N_8511,N_8886);
nor U9213 (N_9213,N_8980,N_8740);
and U9214 (N_9214,N_8725,N_8738);
and U9215 (N_9215,N_8796,N_8809);
nand U9216 (N_9216,N_8469,N_8565);
nand U9217 (N_9217,N_8947,N_8597);
nand U9218 (N_9218,N_8789,N_8395);
nor U9219 (N_9219,N_8779,N_8981);
nor U9220 (N_9220,N_8576,N_8341);
or U9221 (N_9221,N_8343,N_8375);
and U9222 (N_9222,N_8552,N_8663);
and U9223 (N_9223,N_8570,N_8841);
nand U9224 (N_9224,N_8641,N_8415);
and U9225 (N_9225,N_8835,N_8965);
xnor U9226 (N_9226,N_8827,N_8962);
and U9227 (N_9227,N_8852,N_8604);
nand U9228 (N_9228,N_8927,N_8254);
or U9229 (N_9229,N_8499,N_8983);
xnor U9230 (N_9230,N_8384,N_8759);
nand U9231 (N_9231,N_8578,N_8748);
or U9232 (N_9232,N_8275,N_8755);
nor U9233 (N_9233,N_8619,N_8545);
nand U9234 (N_9234,N_8543,N_8795);
nand U9235 (N_9235,N_8417,N_8342);
nand U9236 (N_9236,N_8428,N_8915);
xor U9237 (N_9237,N_8573,N_8630);
or U9238 (N_9238,N_8668,N_8761);
nand U9239 (N_9239,N_8357,N_8493);
xnor U9240 (N_9240,N_8873,N_8561);
or U9241 (N_9241,N_8470,N_8364);
xnor U9242 (N_9242,N_8989,N_8267);
or U9243 (N_9243,N_8888,N_8386);
or U9244 (N_9244,N_8975,N_8557);
or U9245 (N_9245,N_8459,N_8411);
nor U9246 (N_9246,N_8752,N_8849);
and U9247 (N_9247,N_8808,N_8398);
nor U9248 (N_9248,N_8881,N_8378);
nor U9249 (N_9249,N_8497,N_8329);
nor U9250 (N_9250,N_8996,N_8295);
or U9251 (N_9251,N_8262,N_8938);
nand U9252 (N_9252,N_8577,N_8945);
or U9253 (N_9253,N_8458,N_8786);
or U9254 (N_9254,N_8867,N_8525);
and U9255 (N_9255,N_8870,N_8391);
and U9256 (N_9256,N_8664,N_8712);
nor U9257 (N_9257,N_8976,N_8857);
nor U9258 (N_9258,N_8313,N_8899);
xnor U9259 (N_9259,N_8541,N_8730);
or U9260 (N_9260,N_8999,N_8520);
nand U9261 (N_9261,N_8662,N_8971);
nand U9262 (N_9262,N_8929,N_8990);
nand U9263 (N_9263,N_8354,N_8706);
or U9264 (N_9264,N_8746,N_8854);
or U9265 (N_9265,N_8840,N_8859);
or U9266 (N_9266,N_8671,N_8433);
nor U9267 (N_9267,N_8403,N_8917);
and U9268 (N_9268,N_8498,N_8639);
xor U9269 (N_9269,N_8558,N_8766);
xor U9270 (N_9270,N_8412,N_8696);
and U9271 (N_9271,N_8626,N_8294);
and U9272 (N_9272,N_8963,N_8700);
or U9273 (N_9273,N_8489,N_8605);
nor U9274 (N_9274,N_8574,N_8949);
and U9275 (N_9275,N_8355,N_8647);
xor U9276 (N_9276,N_8436,N_8997);
xnor U9277 (N_9277,N_8828,N_8453);
and U9278 (N_9278,N_8910,N_8297);
nand U9279 (N_9279,N_8252,N_8941);
xor U9280 (N_9280,N_8479,N_8743);
or U9281 (N_9281,N_8505,N_8298);
xor U9282 (N_9282,N_8968,N_8751);
and U9283 (N_9283,N_8413,N_8450);
xnor U9284 (N_9284,N_8885,N_8802);
or U9285 (N_9285,N_8957,N_8365);
nor U9286 (N_9286,N_8439,N_8332);
xor U9287 (N_9287,N_8815,N_8509);
xnor U9288 (N_9288,N_8610,N_8421);
and U9289 (N_9289,N_8994,N_8666);
xnor U9290 (N_9290,N_8638,N_8780);
xor U9291 (N_9291,N_8921,N_8584);
nor U9292 (N_9292,N_8868,N_8596);
nand U9293 (N_9293,N_8952,N_8883);
xnor U9294 (N_9294,N_8306,N_8322);
nand U9295 (N_9295,N_8587,N_8367);
nand U9296 (N_9296,N_8829,N_8490);
or U9297 (N_9297,N_8404,N_8871);
xnor U9298 (N_9298,N_8733,N_8956);
xor U9299 (N_9299,N_8353,N_8655);
and U9300 (N_9300,N_8571,N_8644);
and U9301 (N_9301,N_8718,N_8374);
xnor U9302 (N_9302,N_8504,N_8408);
nand U9303 (N_9303,N_8803,N_8288);
or U9304 (N_9304,N_8758,N_8261);
or U9305 (N_9305,N_8898,N_8513);
and U9306 (N_9306,N_8823,N_8592);
nand U9307 (N_9307,N_8256,N_8598);
xor U9308 (N_9308,N_8582,N_8760);
nor U9309 (N_9309,N_8377,N_8463);
xnor U9310 (N_9310,N_8303,N_8928);
nor U9311 (N_9311,N_8904,N_8409);
or U9312 (N_9312,N_8564,N_8651);
xor U9313 (N_9313,N_8389,N_8581);
or U9314 (N_9314,N_8913,N_8820);
xnor U9315 (N_9315,N_8517,N_8514);
nor U9316 (N_9316,N_8555,N_8691);
xor U9317 (N_9317,N_8686,N_8833);
nor U9318 (N_9318,N_8617,N_8452);
xnor U9319 (N_9319,N_8954,N_8893);
and U9320 (N_9320,N_8754,N_8629);
and U9321 (N_9321,N_8838,N_8705);
and U9322 (N_9322,N_8289,N_8672);
xnor U9323 (N_9323,N_8524,N_8781);
and U9324 (N_9324,N_8804,N_8703);
xnor U9325 (N_9325,N_8274,N_8293);
and U9326 (N_9326,N_8481,N_8503);
xor U9327 (N_9327,N_8806,N_8282);
xor U9328 (N_9328,N_8562,N_8264);
nor U9329 (N_9329,N_8831,N_8659);
and U9330 (N_9330,N_8877,N_8722);
xnor U9331 (N_9331,N_8546,N_8969);
xnor U9332 (N_9332,N_8379,N_8670);
xor U9333 (N_9333,N_8708,N_8794);
nor U9334 (N_9334,N_8265,N_8767);
nor U9335 (N_9335,N_8260,N_8445);
nor U9336 (N_9336,N_8344,N_8277);
nor U9337 (N_9337,N_8465,N_8326);
and U9338 (N_9338,N_8438,N_8323);
nand U9339 (N_9339,N_8257,N_8494);
nor U9340 (N_9340,N_8734,N_8347);
or U9341 (N_9341,N_8930,N_8773);
or U9342 (N_9342,N_8652,N_8532);
nor U9343 (N_9343,N_8826,N_8521);
or U9344 (N_9344,N_8745,N_8281);
or U9345 (N_9345,N_8816,N_8625);
and U9346 (N_9346,N_8350,N_8567);
nand U9347 (N_9347,N_8483,N_8542);
nor U9348 (N_9348,N_8958,N_8307);
and U9349 (N_9349,N_8645,N_8966);
xor U9350 (N_9350,N_8846,N_8308);
xnor U9351 (N_9351,N_8848,N_8807);
nand U9352 (N_9352,N_8366,N_8677);
or U9353 (N_9353,N_8352,N_8387);
or U9354 (N_9354,N_8798,N_8843);
nand U9355 (N_9355,N_8757,N_8312);
nor U9356 (N_9356,N_8478,N_8426);
or U9357 (N_9357,N_8618,N_8419);
nand U9358 (N_9358,N_8485,N_8348);
and U9359 (N_9359,N_8475,N_8874);
xnor U9360 (N_9360,N_8797,N_8263);
nand U9361 (N_9361,N_8594,N_8680);
nand U9362 (N_9362,N_8599,N_8661);
xnor U9363 (N_9363,N_8397,N_8932);
or U9364 (N_9364,N_8380,N_8858);
xor U9365 (N_9365,N_8318,N_8477);
xnor U9366 (N_9366,N_8972,N_8632);
or U9367 (N_9367,N_8568,N_8431);
nor U9368 (N_9368,N_8987,N_8301);
nand U9369 (N_9369,N_8728,N_8359);
nor U9370 (N_9370,N_8682,N_8442);
and U9371 (N_9371,N_8948,N_8839);
nand U9372 (N_9372,N_8253,N_8960);
or U9373 (N_9373,N_8636,N_8920);
and U9374 (N_9374,N_8331,N_8548);
and U9375 (N_9375,N_8779,N_8436);
xor U9376 (N_9376,N_8430,N_8736);
nand U9377 (N_9377,N_8422,N_8372);
xor U9378 (N_9378,N_8486,N_8485);
and U9379 (N_9379,N_8652,N_8481);
xor U9380 (N_9380,N_8982,N_8789);
or U9381 (N_9381,N_8673,N_8490);
xor U9382 (N_9382,N_8646,N_8449);
nor U9383 (N_9383,N_8469,N_8490);
nand U9384 (N_9384,N_8366,N_8340);
and U9385 (N_9385,N_8360,N_8253);
nor U9386 (N_9386,N_8856,N_8908);
nor U9387 (N_9387,N_8961,N_8962);
or U9388 (N_9388,N_8423,N_8864);
or U9389 (N_9389,N_8338,N_8578);
xnor U9390 (N_9390,N_8945,N_8373);
xnor U9391 (N_9391,N_8718,N_8477);
nand U9392 (N_9392,N_8757,N_8742);
or U9393 (N_9393,N_8256,N_8487);
nand U9394 (N_9394,N_8518,N_8491);
or U9395 (N_9395,N_8839,N_8803);
nor U9396 (N_9396,N_8252,N_8884);
or U9397 (N_9397,N_8275,N_8439);
and U9398 (N_9398,N_8714,N_8395);
nand U9399 (N_9399,N_8806,N_8817);
and U9400 (N_9400,N_8929,N_8949);
xor U9401 (N_9401,N_8738,N_8485);
or U9402 (N_9402,N_8421,N_8873);
nand U9403 (N_9403,N_8723,N_8506);
xor U9404 (N_9404,N_8338,N_8266);
nor U9405 (N_9405,N_8602,N_8729);
nand U9406 (N_9406,N_8626,N_8434);
or U9407 (N_9407,N_8461,N_8811);
and U9408 (N_9408,N_8393,N_8376);
or U9409 (N_9409,N_8815,N_8320);
nand U9410 (N_9410,N_8499,N_8990);
nor U9411 (N_9411,N_8632,N_8661);
nand U9412 (N_9412,N_8925,N_8747);
nand U9413 (N_9413,N_8887,N_8727);
or U9414 (N_9414,N_8345,N_8349);
and U9415 (N_9415,N_8702,N_8316);
or U9416 (N_9416,N_8386,N_8409);
nor U9417 (N_9417,N_8265,N_8608);
nor U9418 (N_9418,N_8725,N_8862);
or U9419 (N_9419,N_8330,N_8274);
and U9420 (N_9420,N_8478,N_8339);
and U9421 (N_9421,N_8329,N_8969);
xor U9422 (N_9422,N_8577,N_8334);
or U9423 (N_9423,N_8981,N_8950);
or U9424 (N_9424,N_8927,N_8453);
xor U9425 (N_9425,N_8528,N_8968);
and U9426 (N_9426,N_8547,N_8927);
nand U9427 (N_9427,N_8423,N_8722);
nand U9428 (N_9428,N_8655,N_8860);
and U9429 (N_9429,N_8720,N_8275);
or U9430 (N_9430,N_8944,N_8688);
or U9431 (N_9431,N_8945,N_8972);
or U9432 (N_9432,N_8604,N_8463);
or U9433 (N_9433,N_8291,N_8316);
or U9434 (N_9434,N_8557,N_8349);
nor U9435 (N_9435,N_8324,N_8851);
xnor U9436 (N_9436,N_8626,N_8745);
or U9437 (N_9437,N_8352,N_8428);
nand U9438 (N_9438,N_8315,N_8881);
nor U9439 (N_9439,N_8358,N_8978);
and U9440 (N_9440,N_8647,N_8391);
nor U9441 (N_9441,N_8323,N_8318);
xor U9442 (N_9442,N_8933,N_8990);
nor U9443 (N_9443,N_8378,N_8825);
nand U9444 (N_9444,N_8746,N_8351);
nor U9445 (N_9445,N_8892,N_8260);
or U9446 (N_9446,N_8893,N_8299);
and U9447 (N_9447,N_8353,N_8859);
and U9448 (N_9448,N_8468,N_8851);
nand U9449 (N_9449,N_8446,N_8474);
xnor U9450 (N_9450,N_8500,N_8435);
nor U9451 (N_9451,N_8521,N_8734);
nor U9452 (N_9452,N_8342,N_8889);
xor U9453 (N_9453,N_8379,N_8604);
or U9454 (N_9454,N_8517,N_8815);
nand U9455 (N_9455,N_8592,N_8974);
xor U9456 (N_9456,N_8288,N_8350);
and U9457 (N_9457,N_8520,N_8732);
or U9458 (N_9458,N_8338,N_8661);
or U9459 (N_9459,N_8830,N_8576);
nand U9460 (N_9460,N_8829,N_8902);
nand U9461 (N_9461,N_8943,N_8697);
nor U9462 (N_9462,N_8357,N_8910);
and U9463 (N_9463,N_8376,N_8633);
nand U9464 (N_9464,N_8448,N_8489);
and U9465 (N_9465,N_8537,N_8476);
xnor U9466 (N_9466,N_8462,N_8491);
xnor U9467 (N_9467,N_8996,N_8466);
or U9468 (N_9468,N_8463,N_8305);
or U9469 (N_9469,N_8531,N_8735);
and U9470 (N_9470,N_8627,N_8669);
and U9471 (N_9471,N_8774,N_8355);
or U9472 (N_9472,N_8573,N_8932);
xor U9473 (N_9473,N_8737,N_8446);
nand U9474 (N_9474,N_8719,N_8438);
xor U9475 (N_9475,N_8445,N_8988);
or U9476 (N_9476,N_8749,N_8696);
xnor U9477 (N_9477,N_8341,N_8783);
nor U9478 (N_9478,N_8462,N_8946);
nand U9479 (N_9479,N_8561,N_8725);
xnor U9480 (N_9480,N_8665,N_8990);
nand U9481 (N_9481,N_8748,N_8472);
and U9482 (N_9482,N_8748,N_8774);
nor U9483 (N_9483,N_8957,N_8715);
and U9484 (N_9484,N_8332,N_8740);
xnor U9485 (N_9485,N_8869,N_8768);
and U9486 (N_9486,N_8266,N_8464);
or U9487 (N_9487,N_8692,N_8913);
nand U9488 (N_9488,N_8277,N_8364);
and U9489 (N_9489,N_8322,N_8520);
and U9490 (N_9490,N_8867,N_8431);
xnor U9491 (N_9491,N_8960,N_8654);
or U9492 (N_9492,N_8430,N_8873);
nor U9493 (N_9493,N_8936,N_8711);
xor U9494 (N_9494,N_8479,N_8288);
nor U9495 (N_9495,N_8960,N_8639);
nand U9496 (N_9496,N_8634,N_8775);
nor U9497 (N_9497,N_8301,N_8274);
xnor U9498 (N_9498,N_8475,N_8396);
and U9499 (N_9499,N_8488,N_8387);
xor U9500 (N_9500,N_8344,N_8267);
xor U9501 (N_9501,N_8407,N_8789);
or U9502 (N_9502,N_8655,N_8644);
and U9503 (N_9503,N_8570,N_8461);
and U9504 (N_9504,N_8980,N_8504);
nor U9505 (N_9505,N_8517,N_8921);
nor U9506 (N_9506,N_8979,N_8611);
xor U9507 (N_9507,N_8677,N_8273);
and U9508 (N_9508,N_8265,N_8307);
nor U9509 (N_9509,N_8417,N_8727);
and U9510 (N_9510,N_8765,N_8627);
nand U9511 (N_9511,N_8267,N_8376);
or U9512 (N_9512,N_8306,N_8780);
and U9513 (N_9513,N_8630,N_8739);
xor U9514 (N_9514,N_8380,N_8566);
xor U9515 (N_9515,N_8956,N_8439);
nor U9516 (N_9516,N_8723,N_8764);
xor U9517 (N_9517,N_8331,N_8635);
nand U9518 (N_9518,N_8448,N_8859);
xor U9519 (N_9519,N_8507,N_8777);
nor U9520 (N_9520,N_8325,N_8259);
nand U9521 (N_9521,N_8970,N_8917);
nor U9522 (N_9522,N_8418,N_8840);
nand U9523 (N_9523,N_8254,N_8387);
xnor U9524 (N_9524,N_8270,N_8815);
xor U9525 (N_9525,N_8767,N_8872);
xor U9526 (N_9526,N_8291,N_8769);
and U9527 (N_9527,N_8368,N_8650);
and U9528 (N_9528,N_8670,N_8316);
xnor U9529 (N_9529,N_8511,N_8329);
and U9530 (N_9530,N_8459,N_8549);
nor U9531 (N_9531,N_8346,N_8335);
or U9532 (N_9532,N_8482,N_8366);
and U9533 (N_9533,N_8958,N_8569);
nor U9534 (N_9534,N_8445,N_8474);
nor U9535 (N_9535,N_8564,N_8358);
or U9536 (N_9536,N_8562,N_8372);
and U9537 (N_9537,N_8678,N_8704);
or U9538 (N_9538,N_8568,N_8968);
or U9539 (N_9539,N_8402,N_8762);
xor U9540 (N_9540,N_8702,N_8657);
nor U9541 (N_9541,N_8609,N_8866);
nand U9542 (N_9542,N_8646,N_8454);
or U9543 (N_9543,N_8787,N_8688);
or U9544 (N_9544,N_8251,N_8371);
and U9545 (N_9545,N_8906,N_8690);
xor U9546 (N_9546,N_8742,N_8910);
nand U9547 (N_9547,N_8405,N_8871);
xor U9548 (N_9548,N_8632,N_8512);
or U9549 (N_9549,N_8946,N_8945);
xnor U9550 (N_9550,N_8794,N_8762);
and U9551 (N_9551,N_8259,N_8928);
or U9552 (N_9552,N_8869,N_8815);
or U9553 (N_9553,N_8579,N_8877);
nand U9554 (N_9554,N_8805,N_8886);
and U9555 (N_9555,N_8254,N_8662);
xnor U9556 (N_9556,N_8641,N_8284);
and U9557 (N_9557,N_8980,N_8669);
nor U9558 (N_9558,N_8561,N_8884);
nand U9559 (N_9559,N_8448,N_8499);
or U9560 (N_9560,N_8399,N_8385);
and U9561 (N_9561,N_8492,N_8766);
or U9562 (N_9562,N_8606,N_8317);
and U9563 (N_9563,N_8495,N_8640);
or U9564 (N_9564,N_8994,N_8423);
nor U9565 (N_9565,N_8308,N_8264);
nor U9566 (N_9566,N_8305,N_8565);
and U9567 (N_9567,N_8632,N_8859);
or U9568 (N_9568,N_8711,N_8331);
nor U9569 (N_9569,N_8993,N_8817);
nor U9570 (N_9570,N_8272,N_8977);
nand U9571 (N_9571,N_8702,N_8298);
and U9572 (N_9572,N_8456,N_8880);
and U9573 (N_9573,N_8507,N_8626);
nand U9574 (N_9574,N_8313,N_8440);
xor U9575 (N_9575,N_8773,N_8592);
nor U9576 (N_9576,N_8348,N_8593);
or U9577 (N_9577,N_8361,N_8445);
and U9578 (N_9578,N_8344,N_8834);
nor U9579 (N_9579,N_8345,N_8422);
and U9580 (N_9580,N_8583,N_8590);
xnor U9581 (N_9581,N_8427,N_8989);
nand U9582 (N_9582,N_8638,N_8868);
nand U9583 (N_9583,N_8617,N_8600);
or U9584 (N_9584,N_8600,N_8795);
nand U9585 (N_9585,N_8879,N_8490);
xnor U9586 (N_9586,N_8575,N_8319);
nand U9587 (N_9587,N_8500,N_8490);
or U9588 (N_9588,N_8977,N_8862);
and U9589 (N_9589,N_8654,N_8502);
or U9590 (N_9590,N_8773,N_8634);
or U9591 (N_9591,N_8340,N_8397);
or U9592 (N_9592,N_8875,N_8321);
or U9593 (N_9593,N_8328,N_8567);
and U9594 (N_9594,N_8449,N_8514);
xor U9595 (N_9595,N_8773,N_8934);
nor U9596 (N_9596,N_8364,N_8589);
or U9597 (N_9597,N_8294,N_8771);
or U9598 (N_9598,N_8582,N_8350);
nor U9599 (N_9599,N_8321,N_8296);
nand U9600 (N_9600,N_8410,N_8719);
and U9601 (N_9601,N_8594,N_8519);
xor U9602 (N_9602,N_8784,N_8637);
xor U9603 (N_9603,N_8758,N_8685);
nand U9604 (N_9604,N_8822,N_8793);
and U9605 (N_9605,N_8721,N_8996);
or U9606 (N_9606,N_8651,N_8837);
or U9607 (N_9607,N_8903,N_8623);
or U9608 (N_9608,N_8928,N_8521);
nand U9609 (N_9609,N_8456,N_8822);
xor U9610 (N_9610,N_8485,N_8819);
or U9611 (N_9611,N_8327,N_8412);
and U9612 (N_9612,N_8553,N_8574);
nor U9613 (N_9613,N_8693,N_8923);
and U9614 (N_9614,N_8424,N_8760);
and U9615 (N_9615,N_8609,N_8899);
and U9616 (N_9616,N_8291,N_8799);
or U9617 (N_9617,N_8607,N_8614);
xnor U9618 (N_9618,N_8508,N_8859);
or U9619 (N_9619,N_8813,N_8434);
nand U9620 (N_9620,N_8495,N_8284);
xor U9621 (N_9621,N_8361,N_8392);
and U9622 (N_9622,N_8320,N_8273);
or U9623 (N_9623,N_8462,N_8951);
or U9624 (N_9624,N_8635,N_8388);
and U9625 (N_9625,N_8314,N_8472);
or U9626 (N_9626,N_8848,N_8884);
or U9627 (N_9627,N_8345,N_8948);
nand U9628 (N_9628,N_8904,N_8391);
or U9629 (N_9629,N_8602,N_8636);
nor U9630 (N_9630,N_8578,N_8302);
xnor U9631 (N_9631,N_8704,N_8521);
xor U9632 (N_9632,N_8255,N_8791);
xnor U9633 (N_9633,N_8971,N_8569);
xor U9634 (N_9634,N_8460,N_8510);
or U9635 (N_9635,N_8712,N_8909);
xor U9636 (N_9636,N_8654,N_8797);
or U9637 (N_9637,N_8805,N_8952);
nor U9638 (N_9638,N_8327,N_8930);
or U9639 (N_9639,N_8810,N_8982);
and U9640 (N_9640,N_8326,N_8991);
nand U9641 (N_9641,N_8871,N_8361);
nand U9642 (N_9642,N_8478,N_8870);
or U9643 (N_9643,N_8861,N_8343);
or U9644 (N_9644,N_8656,N_8467);
xnor U9645 (N_9645,N_8583,N_8444);
nand U9646 (N_9646,N_8459,N_8641);
or U9647 (N_9647,N_8418,N_8348);
xnor U9648 (N_9648,N_8431,N_8416);
or U9649 (N_9649,N_8454,N_8935);
and U9650 (N_9650,N_8620,N_8288);
and U9651 (N_9651,N_8313,N_8278);
and U9652 (N_9652,N_8449,N_8747);
nand U9653 (N_9653,N_8782,N_8485);
and U9654 (N_9654,N_8927,N_8365);
nor U9655 (N_9655,N_8560,N_8344);
nand U9656 (N_9656,N_8466,N_8824);
xor U9657 (N_9657,N_8437,N_8526);
xor U9658 (N_9658,N_8543,N_8304);
nand U9659 (N_9659,N_8839,N_8445);
nand U9660 (N_9660,N_8766,N_8391);
xnor U9661 (N_9661,N_8854,N_8711);
nor U9662 (N_9662,N_8611,N_8439);
xor U9663 (N_9663,N_8442,N_8435);
or U9664 (N_9664,N_8376,N_8383);
and U9665 (N_9665,N_8795,N_8334);
nand U9666 (N_9666,N_8962,N_8525);
xnor U9667 (N_9667,N_8927,N_8320);
nand U9668 (N_9668,N_8761,N_8794);
or U9669 (N_9669,N_8785,N_8795);
xor U9670 (N_9670,N_8954,N_8845);
xnor U9671 (N_9671,N_8811,N_8720);
xnor U9672 (N_9672,N_8876,N_8337);
nor U9673 (N_9673,N_8414,N_8770);
xor U9674 (N_9674,N_8255,N_8427);
nor U9675 (N_9675,N_8945,N_8467);
xor U9676 (N_9676,N_8862,N_8876);
or U9677 (N_9677,N_8461,N_8251);
xor U9678 (N_9678,N_8768,N_8687);
or U9679 (N_9679,N_8874,N_8678);
or U9680 (N_9680,N_8798,N_8359);
xor U9681 (N_9681,N_8852,N_8349);
nor U9682 (N_9682,N_8533,N_8474);
and U9683 (N_9683,N_8710,N_8401);
nand U9684 (N_9684,N_8818,N_8676);
xnor U9685 (N_9685,N_8474,N_8866);
or U9686 (N_9686,N_8718,N_8826);
and U9687 (N_9687,N_8891,N_8500);
and U9688 (N_9688,N_8534,N_8297);
nand U9689 (N_9689,N_8933,N_8436);
nor U9690 (N_9690,N_8754,N_8536);
nor U9691 (N_9691,N_8831,N_8917);
xor U9692 (N_9692,N_8906,N_8934);
and U9693 (N_9693,N_8661,N_8648);
or U9694 (N_9694,N_8364,N_8250);
xnor U9695 (N_9695,N_8483,N_8864);
and U9696 (N_9696,N_8574,N_8795);
and U9697 (N_9697,N_8944,N_8296);
xor U9698 (N_9698,N_8715,N_8295);
and U9699 (N_9699,N_8955,N_8987);
and U9700 (N_9700,N_8740,N_8843);
nor U9701 (N_9701,N_8312,N_8281);
nand U9702 (N_9702,N_8364,N_8251);
nand U9703 (N_9703,N_8446,N_8309);
xnor U9704 (N_9704,N_8407,N_8898);
or U9705 (N_9705,N_8560,N_8320);
and U9706 (N_9706,N_8821,N_8745);
nor U9707 (N_9707,N_8966,N_8828);
nand U9708 (N_9708,N_8587,N_8938);
xnor U9709 (N_9709,N_8375,N_8336);
nor U9710 (N_9710,N_8307,N_8519);
or U9711 (N_9711,N_8652,N_8581);
nor U9712 (N_9712,N_8768,N_8903);
or U9713 (N_9713,N_8547,N_8649);
nor U9714 (N_9714,N_8748,N_8487);
or U9715 (N_9715,N_8529,N_8333);
nor U9716 (N_9716,N_8490,N_8667);
or U9717 (N_9717,N_8939,N_8539);
nor U9718 (N_9718,N_8293,N_8840);
or U9719 (N_9719,N_8924,N_8755);
and U9720 (N_9720,N_8939,N_8256);
nand U9721 (N_9721,N_8326,N_8762);
nor U9722 (N_9722,N_8671,N_8525);
or U9723 (N_9723,N_8672,N_8308);
and U9724 (N_9724,N_8977,N_8884);
nand U9725 (N_9725,N_8664,N_8336);
xor U9726 (N_9726,N_8263,N_8497);
and U9727 (N_9727,N_8818,N_8674);
nand U9728 (N_9728,N_8912,N_8926);
and U9729 (N_9729,N_8949,N_8852);
xor U9730 (N_9730,N_8816,N_8896);
nand U9731 (N_9731,N_8592,N_8955);
nor U9732 (N_9732,N_8414,N_8466);
and U9733 (N_9733,N_8621,N_8635);
nor U9734 (N_9734,N_8664,N_8733);
nor U9735 (N_9735,N_8840,N_8415);
nand U9736 (N_9736,N_8847,N_8540);
or U9737 (N_9737,N_8719,N_8588);
nand U9738 (N_9738,N_8429,N_8403);
or U9739 (N_9739,N_8414,N_8724);
xor U9740 (N_9740,N_8600,N_8281);
nor U9741 (N_9741,N_8310,N_8745);
xor U9742 (N_9742,N_8482,N_8480);
xnor U9743 (N_9743,N_8902,N_8344);
or U9744 (N_9744,N_8358,N_8441);
nand U9745 (N_9745,N_8743,N_8602);
and U9746 (N_9746,N_8940,N_8839);
nand U9747 (N_9747,N_8914,N_8582);
and U9748 (N_9748,N_8355,N_8562);
nand U9749 (N_9749,N_8541,N_8319);
and U9750 (N_9750,N_9556,N_9209);
or U9751 (N_9751,N_9561,N_9445);
and U9752 (N_9752,N_9048,N_9329);
and U9753 (N_9753,N_9088,N_9196);
xor U9754 (N_9754,N_9482,N_9373);
or U9755 (N_9755,N_9041,N_9162);
nor U9756 (N_9756,N_9706,N_9632);
xnor U9757 (N_9757,N_9524,N_9083);
and U9758 (N_9758,N_9584,N_9473);
and U9759 (N_9759,N_9058,N_9310);
nor U9760 (N_9760,N_9689,N_9281);
nand U9761 (N_9761,N_9105,N_9234);
nor U9762 (N_9762,N_9189,N_9344);
nand U9763 (N_9763,N_9051,N_9537);
xnor U9764 (N_9764,N_9271,N_9007);
nand U9765 (N_9765,N_9429,N_9486);
nor U9766 (N_9766,N_9700,N_9495);
nand U9767 (N_9767,N_9314,N_9625);
nor U9768 (N_9768,N_9669,N_9060);
nor U9769 (N_9769,N_9628,N_9484);
xor U9770 (N_9770,N_9559,N_9175);
and U9771 (N_9771,N_9572,N_9682);
nand U9772 (N_9772,N_9433,N_9115);
and U9773 (N_9773,N_9728,N_9404);
and U9774 (N_9774,N_9389,N_9139);
xor U9775 (N_9775,N_9457,N_9427);
nor U9776 (N_9776,N_9215,N_9423);
xnor U9777 (N_9777,N_9376,N_9093);
xnor U9778 (N_9778,N_9507,N_9421);
nand U9779 (N_9779,N_9574,N_9341);
or U9780 (N_9780,N_9532,N_9173);
or U9781 (N_9781,N_9049,N_9428);
nor U9782 (N_9782,N_9521,N_9040);
and U9783 (N_9783,N_9303,N_9431);
and U9784 (N_9784,N_9255,N_9006);
xor U9785 (N_9785,N_9459,N_9560);
xor U9786 (N_9786,N_9348,N_9265);
nor U9787 (N_9787,N_9074,N_9701);
or U9788 (N_9788,N_9541,N_9598);
and U9789 (N_9789,N_9177,N_9424);
nor U9790 (N_9790,N_9462,N_9277);
or U9791 (N_9791,N_9745,N_9050);
nand U9792 (N_9792,N_9213,N_9320);
nand U9793 (N_9793,N_9035,N_9061);
nand U9794 (N_9794,N_9515,N_9723);
nor U9795 (N_9795,N_9401,N_9097);
nand U9796 (N_9796,N_9544,N_9328);
xor U9797 (N_9797,N_9343,N_9152);
or U9798 (N_9798,N_9629,N_9678);
xnor U9799 (N_9799,N_9031,N_9090);
xnor U9800 (N_9800,N_9206,N_9695);
or U9801 (N_9801,N_9597,N_9295);
nor U9802 (N_9802,N_9370,N_9317);
nor U9803 (N_9803,N_9475,N_9354);
xor U9804 (N_9804,N_9523,N_9399);
or U9805 (N_9805,N_9141,N_9436);
nand U9806 (N_9806,N_9571,N_9359);
and U9807 (N_9807,N_9697,N_9346);
nor U9808 (N_9808,N_9202,N_9184);
nand U9809 (N_9809,N_9086,N_9166);
or U9810 (N_9810,N_9302,N_9722);
and U9811 (N_9811,N_9703,N_9052);
or U9812 (N_9812,N_9043,N_9583);
nor U9813 (N_9813,N_9749,N_9319);
nor U9814 (N_9814,N_9321,N_9670);
nand U9815 (N_9815,N_9621,N_9690);
nor U9816 (N_9816,N_9525,N_9563);
nand U9817 (N_9817,N_9084,N_9518);
or U9818 (N_9818,N_9407,N_9451);
or U9819 (N_9819,N_9594,N_9284);
or U9820 (N_9820,N_9642,N_9022);
and U9821 (N_9821,N_9668,N_9671);
or U9822 (N_9822,N_9080,N_9460);
and U9823 (N_9823,N_9365,N_9023);
nor U9824 (N_9824,N_9551,N_9120);
nor U9825 (N_9825,N_9600,N_9603);
or U9826 (N_9826,N_9536,N_9231);
xnor U9827 (N_9827,N_9463,N_9182);
xor U9828 (N_9828,N_9077,N_9245);
nand U9829 (N_9829,N_9230,N_9092);
and U9830 (N_9830,N_9241,N_9294);
nand U9831 (N_9831,N_9588,N_9510);
nand U9832 (N_9832,N_9480,N_9575);
xnor U9833 (N_9833,N_9454,N_9705);
nand U9834 (N_9834,N_9717,N_9117);
xor U9835 (N_9835,N_9103,N_9698);
nor U9836 (N_9836,N_9639,N_9727);
nand U9837 (N_9837,N_9154,N_9195);
xnor U9838 (N_9838,N_9529,N_9526);
xnor U9839 (N_9839,N_9025,N_9226);
nand U9840 (N_9840,N_9216,N_9297);
nand U9841 (N_9841,N_9334,N_9714);
nor U9842 (N_9842,N_9720,N_9742);
and U9843 (N_9843,N_9194,N_9548);
xor U9844 (N_9844,N_9638,N_9100);
nor U9845 (N_9845,N_9267,N_9176);
or U9846 (N_9846,N_9063,N_9251);
nand U9847 (N_9847,N_9223,N_9178);
nand U9848 (N_9848,N_9527,N_9019);
or U9849 (N_9849,N_9055,N_9726);
and U9850 (N_9850,N_9564,N_9264);
or U9851 (N_9851,N_9101,N_9474);
nand U9852 (N_9852,N_9448,N_9687);
nand U9853 (N_9853,N_9520,N_9640);
or U9854 (N_9854,N_9307,N_9498);
xor U9855 (N_9855,N_9693,N_9630);
nor U9856 (N_9856,N_9337,N_9624);
nand U9857 (N_9857,N_9153,N_9441);
xnor U9858 (N_9858,N_9374,N_9652);
and U9859 (N_9859,N_9593,N_9437);
xnor U9860 (N_9860,N_9067,N_9596);
or U9861 (N_9861,N_9609,N_9045);
or U9862 (N_9862,N_9469,N_9270);
xor U9863 (N_9863,N_9724,N_9165);
and U9864 (N_9864,N_9378,N_9410);
nand U9865 (N_9865,N_9253,N_9591);
and U9866 (N_9866,N_9535,N_9286);
xor U9867 (N_9867,N_9738,N_9491);
and U9868 (N_9868,N_9691,N_9179);
nor U9869 (N_9869,N_9029,N_9056);
nor U9870 (N_9870,N_9015,N_9237);
and U9871 (N_9871,N_9464,N_9085);
nand U9872 (N_9872,N_9138,N_9570);
or U9873 (N_9873,N_9707,N_9272);
nor U9874 (N_9874,N_9125,N_9538);
and U9875 (N_9875,N_9132,N_9409);
and U9876 (N_9876,N_9046,N_9108);
and U9877 (N_9877,N_9042,N_9386);
nand U9878 (N_9878,N_9499,N_9287);
nand U9879 (N_9879,N_9017,N_9361);
nor U9880 (N_9880,N_9497,N_9737);
xor U9881 (N_9881,N_9406,N_9371);
or U9882 (N_9882,N_9362,N_9512);
nor U9883 (N_9883,N_9010,N_9552);
and U9884 (N_9884,N_9385,N_9351);
or U9885 (N_9885,N_9211,N_9266);
or U9886 (N_9886,N_9496,N_9133);
and U9887 (N_9887,N_9034,N_9384);
nand U9888 (N_9888,N_9716,N_9543);
or U9889 (N_9889,N_9135,N_9679);
xor U9890 (N_9890,N_9070,N_9503);
nor U9891 (N_9891,N_9068,N_9109);
xnor U9892 (N_9892,N_9078,N_9350);
xor U9893 (N_9893,N_9533,N_9468);
xnor U9894 (N_9894,N_9592,N_9030);
nor U9895 (N_9895,N_9402,N_9147);
xor U9896 (N_9896,N_9220,N_9225);
or U9897 (N_9897,N_9653,N_9285);
or U9898 (N_9898,N_9106,N_9188);
xor U9899 (N_9899,N_9443,N_9089);
nand U9900 (N_9900,N_9504,N_9364);
xnor U9901 (N_9901,N_9259,N_9488);
xor U9902 (N_9902,N_9242,N_9221);
or U9903 (N_9903,N_9394,N_9203);
and U9904 (N_9904,N_9741,N_9479);
xor U9905 (N_9905,N_9201,N_9318);
or U9906 (N_9906,N_9467,N_9466);
xnor U9907 (N_9907,N_9210,N_9168);
nand U9908 (N_9908,N_9587,N_9159);
nand U9909 (N_9909,N_9744,N_9633);
xnor U9910 (N_9910,N_9011,N_9708);
nand U9911 (N_9911,N_9039,N_9390);
or U9912 (N_9912,N_9249,N_9155);
nor U9913 (N_9913,N_9069,N_9053);
nand U9914 (N_9914,N_9595,N_9037);
and U9915 (N_9915,N_9331,N_9094);
nor U9916 (N_9916,N_9477,N_9180);
nand U9917 (N_9917,N_9146,N_9440);
xnor U9918 (N_9918,N_9517,N_9143);
and U9919 (N_9919,N_9710,N_9696);
nor U9920 (N_9920,N_9313,N_9262);
xnor U9921 (N_9921,N_9719,N_9425);
nand U9922 (N_9922,N_9000,N_9128);
nor U9923 (N_9923,N_9065,N_9487);
or U9924 (N_9924,N_9227,N_9432);
and U9925 (N_9925,N_9008,N_9446);
nor U9926 (N_9926,N_9326,N_9016);
or U9927 (N_9927,N_9301,N_9157);
xnor U9928 (N_9928,N_9554,N_9415);
nand U9929 (N_9929,N_9660,N_9740);
and U9930 (N_9930,N_9347,N_9002);
nor U9931 (N_9931,N_9072,N_9131);
nand U9932 (N_9932,N_9528,N_9566);
nand U9933 (N_9933,N_9293,N_9263);
nor U9934 (N_9934,N_9243,N_9369);
xor U9935 (N_9935,N_9372,N_9485);
and U9936 (N_9936,N_9438,N_9082);
or U9937 (N_9937,N_9229,N_9519);
nor U9938 (N_9938,N_9033,N_9456);
nand U9939 (N_9939,N_9306,N_9662);
and U9940 (N_9940,N_9183,N_9481);
or U9941 (N_9941,N_9397,N_9119);
nor U9942 (N_9942,N_9309,N_9735);
nor U9943 (N_9943,N_9279,N_9611);
nor U9944 (N_9944,N_9127,N_9743);
and U9945 (N_9945,N_9140,N_9620);
and U9946 (N_9946,N_9686,N_9332);
nor U9947 (N_9947,N_9449,N_9396);
nand U9948 (N_9948,N_9324,N_9156);
and U9949 (N_9949,N_9607,N_9026);
or U9950 (N_9950,N_9066,N_9038);
and U9951 (N_9951,N_9569,N_9247);
xnor U9952 (N_9952,N_9470,N_9439);
nand U9953 (N_9953,N_9228,N_9192);
xnor U9954 (N_9954,N_9618,N_9167);
or U9955 (N_9955,N_9218,N_9236);
or U9956 (N_9956,N_9522,N_9126);
and U9957 (N_9957,N_9692,N_9096);
nand U9958 (N_9958,N_9557,N_9024);
and U9959 (N_9959,N_9114,N_9059);
nor U9960 (N_9960,N_9214,N_9158);
xnor U9961 (N_9961,N_9534,N_9455);
nand U9962 (N_9962,N_9204,N_9412);
xnor U9963 (N_9963,N_9684,N_9252);
nand U9964 (N_9964,N_9336,N_9208);
nor U9965 (N_9965,N_9680,N_9513);
and U9966 (N_9966,N_9617,N_9028);
nand U9967 (N_9967,N_9582,N_9161);
nand U9968 (N_9968,N_9516,N_9137);
or U9969 (N_9969,N_9663,N_9721);
and U9970 (N_9970,N_9036,N_9207);
and U9971 (N_9971,N_9296,N_9646);
xor U9972 (N_9972,N_9170,N_9258);
or U9973 (N_9973,N_9636,N_9657);
nand U9974 (N_9974,N_9327,N_9174);
and U9975 (N_9975,N_9076,N_9565);
xor U9976 (N_9976,N_9647,N_9338);
and U9977 (N_9977,N_9062,N_9257);
or U9978 (N_9978,N_9021,N_9379);
or U9979 (N_9979,N_9568,N_9136);
or U9980 (N_9980,N_9079,N_9553);
or U9981 (N_9981,N_9116,N_9308);
or U9982 (N_9982,N_9420,N_9240);
xor U9983 (N_9983,N_9368,N_9323);
nor U9984 (N_9984,N_9367,N_9181);
nand U9985 (N_9985,N_9057,N_9312);
xnor U9986 (N_9986,N_9643,N_9111);
nand U9987 (N_9987,N_9375,N_9278);
or U9988 (N_9988,N_9748,N_9577);
xor U9989 (N_9989,N_9235,N_9381);
xnor U9990 (N_9990,N_9704,N_9260);
or U9991 (N_9991,N_9222,N_9434);
nor U9992 (N_9992,N_9102,N_9465);
nand U9993 (N_9993,N_9458,N_9715);
nor U9994 (N_9994,N_9547,N_9442);
nand U9995 (N_9995,N_9567,N_9411);
nand U9996 (N_9996,N_9430,N_9349);
nand U9997 (N_9997,N_9492,N_9736);
and U9998 (N_9998,N_9601,N_9233);
nand U9999 (N_9999,N_9651,N_9185);
nand U10000 (N_10000,N_9667,N_9345);
nor U10001 (N_10001,N_9644,N_9305);
xnor U10002 (N_10002,N_9500,N_9112);
nor U10003 (N_10003,N_9164,N_9382);
nand U10004 (N_10004,N_9450,N_9675);
nand U10005 (N_10005,N_9316,N_9366);
and U10006 (N_10006,N_9353,N_9502);
and U10007 (N_10007,N_9713,N_9616);
xor U10008 (N_10008,N_9676,N_9032);
or U10009 (N_10009,N_9471,N_9254);
nand U10010 (N_10010,N_9580,N_9380);
nand U10011 (N_10011,N_9013,N_9645);
xnor U10012 (N_10012,N_9476,N_9699);
nor U10013 (N_10013,N_9613,N_9718);
and U10014 (N_10014,N_9299,N_9615);
xnor U10015 (N_10015,N_9709,N_9672);
or U10016 (N_10016,N_9405,N_9542);
nand U10017 (N_10017,N_9012,N_9198);
and U10018 (N_10018,N_9729,N_9095);
nor U10019 (N_10019,N_9360,N_9549);
or U10020 (N_10020,N_9483,N_9656);
nor U10021 (N_10021,N_9619,N_9416);
nand U10022 (N_10022,N_9268,N_9414);
nand U10023 (N_10023,N_9357,N_9356);
nand U10024 (N_10024,N_9732,N_9578);
or U10025 (N_10025,N_9586,N_9605);
and U10026 (N_10026,N_9001,N_9129);
and U10027 (N_10027,N_9702,N_9419);
xnor U10028 (N_10028,N_9163,N_9747);
and U10029 (N_10029,N_9661,N_9422);
and U10030 (N_10030,N_9355,N_9435);
xor U10031 (N_10031,N_9335,N_9623);
nand U10032 (N_10032,N_9004,N_9683);
nand U10033 (N_10033,N_9634,N_9725);
nand U10034 (N_10034,N_9280,N_9508);
xor U10035 (N_10035,N_9387,N_9674);
nand U10036 (N_10036,N_9217,N_9340);
nor U10037 (N_10037,N_9071,N_9232);
or U10038 (N_10038,N_9087,N_9694);
nand U10039 (N_10039,N_9734,N_9506);
nand U10040 (N_10040,N_9493,N_9191);
nand U10041 (N_10041,N_9169,N_9447);
or U10042 (N_10042,N_9148,N_9673);
and U10043 (N_10043,N_9681,N_9426);
and U10044 (N_10044,N_9107,N_9637);
xnor U10045 (N_10045,N_9635,N_9418);
and U10046 (N_10046,N_9339,N_9540);
or U10047 (N_10047,N_9144,N_9150);
and U10048 (N_10048,N_9124,N_9289);
nand U10049 (N_10049,N_9311,N_9205);
and U10050 (N_10050,N_9047,N_9453);
and U10051 (N_10051,N_9298,N_9461);
and U10052 (N_10052,N_9193,N_9573);
xor U10053 (N_10053,N_9711,N_9145);
and U10054 (N_10054,N_9160,N_9123);
xor U10055 (N_10055,N_9333,N_9490);
and U10056 (N_10056,N_9200,N_9290);
nand U10057 (N_10057,N_9283,N_9555);
nand U10058 (N_10058,N_9020,N_9562);
nand U10059 (N_10059,N_9315,N_9590);
or U10060 (N_10060,N_9186,N_9199);
nand U10061 (N_10061,N_9121,N_9505);
nand U10062 (N_10062,N_9091,N_9134);
and U10063 (N_10063,N_9395,N_9612);
or U10064 (N_10064,N_9014,N_9044);
or U10065 (N_10065,N_9608,N_9224);
nand U10066 (N_10066,N_9576,N_9585);
or U10067 (N_10067,N_9546,N_9610);
nand U10068 (N_10068,N_9300,N_9501);
xnor U10069 (N_10069,N_9392,N_9151);
nor U10070 (N_10070,N_9602,N_9444);
or U10071 (N_10071,N_9282,N_9212);
xnor U10072 (N_10072,N_9325,N_9400);
nor U10073 (N_10073,N_9452,N_9579);
xnor U10074 (N_10074,N_9739,N_9330);
nor U10075 (N_10075,N_9172,N_9531);
or U10076 (N_10076,N_9352,N_9027);
nor U10077 (N_10077,N_9322,N_9648);
nor U10078 (N_10078,N_9110,N_9604);
and U10079 (N_10079,N_9197,N_9246);
xnor U10080 (N_10080,N_9539,N_9417);
nor U10081 (N_10081,N_9403,N_9149);
and U10082 (N_10082,N_9276,N_9658);
or U10083 (N_10083,N_9666,N_9530);
xnor U10084 (N_10084,N_9275,N_9377);
or U10085 (N_10085,N_9187,N_9659);
or U10086 (N_10086,N_9599,N_9073);
and U10087 (N_10087,N_9269,N_9098);
xnor U10088 (N_10088,N_9730,N_9064);
or U10089 (N_10089,N_9514,N_9489);
xor U10090 (N_10090,N_9104,N_9472);
xnor U10091 (N_10091,N_9746,N_9654);
nor U10092 (N_10092,N_9494,N_9688);
nor U10093 (N_10093,N_9122,N_9250);
nand U10094 (N_10094,N_9009,N_9363);
xnor U10095 (N_10095,N_9342,N_9248);
or U10096 (N_10096,N_9550,N_9589);
or U10097 (N_10097,N_9075,N_9244);
xor U10098 (N_10098,N_9190,N_9358);
or U10099 (N_10099,N_9677,N_9731);
xnor U10100 (N_10100,N_9509,N_9099);
nand U10101 (N_10101,N_9622,N_9388);
and U10102 (N_10102,N_9408,N_9606);
or U10103 (N_10103,N_9398,N_9054);
nand U10104 (N_10104,N_9274,N_9413);
xnor U10105 (N_10105,N_9733,N_9511);
xnor U10106 (N_10106,N_9018,N_9558);
nor U10107 (N_10107,N_9614,N_9383);
and U10108 (N_10108,N_9256,N_9627);
and U10109 (N_10109,N_9081,N_9239);
nor U10110 (N_10110,N_9118,N_9664);
xnor U10111 (N_10111,N_9005,N_9685);
nor U10112 (N_10112,N_9665,N_9712);
or U10113 (N_10113,N_9238,N_9304);
xnor U10114 (N_10114,N_9581,N_9391);
nor U10115 (N_10115,N_9130,N_9626);
xnor U10116 (N_10116,N_9631,N_9142);
nand U10117 (N_10117,N_9650,N_9113);
nand U10118 (N_10118,N_9292,N_9393);
nor U10119 (N_10119,N_9273,N_9641);
nand U10120 (N_10120,N_9288,N_9655);
xor U10121 (N_10121,N_9171,N_9478);
xnor U10122 (N_10122,N_9261,N_9003);
or U10123 (N_10123,N_9649,N_9545);
and U10124 (N_10124,N_9291,N_9219);
or U10125 (N_10125,N_9211,N_9283);
nand U10126 (N_10126,N_9691,N_9079);
xor U10127 (N_10127,N_9301,N_9548);
nand U10128 (N_10128,N_9539,N_9205);
nand U10129 (N_10129,N_9186,N_9095);
or U10130 (N_10130,N_9289,N_9203);
and U10131 (N_10131,N_9685,N_9700);
and U10132 (N_10132,N_9233,N_9434);
or U10133 (N_10133,N_9592,N_9453);
and U10134 (N_10134,N_9078,N_9263);
nor U10135 (N_10135,N_9699,N_9161);
or U10136 (N_10136,N_9177,N_9184);
xor U10137 (N_10137,N_9638,N_9293);
xor U10138 (N_10138,N_9537,N_9456);
nor U10139 (N_10139,N_9733,N_9293);
nor U10140 (N_10140,N_9390,N_9541);
nand U10141 (N_10141,N_9644,N_9503);
and U10142 (N_10142,N_9173,N_9293);
nor U10143 (N_10143,N_9715,N_9126);
or U10144 (N_10144,N_9153,N_9563);
xor U10145 (N_10145,N_9093,N_9427);
nor U10146 (N_10146,N_9177,N_9613);
nand U10147 (N_10147,N_9322,N_9238);
nor U10148 (N_10148,N_9195,N_9462);
xor U10149 (N_10149,N_9180,N_9644);
or U10150 (N_10150,N_9079,N_9159);
nand U10151 (N_10151,N_9623,N_9221);
xnor U10152 (N_10152,N_9650,N_9338);
and U10153 (N_10153,N_9220,N_9517);
nor U10154 (N_10154,N_9473,N_9017);
or U10155 (N_10155,N_9435,N_9084);
or U10156 (N_10156,N_9316,N_9256);
and U10157 (N_10157,N_9551,N_9240);
and U10158 (N_10158,N_9433,N_9346);
xnor U10159 (N_10159,N_9552,N_9063);
and U10160 (N_10160,N_9634,N_9490);
and U10161 (N_10161,N_9275,N_9558);
and U10162 (N_10162,N_9116,N_9590);
xnor U10163 (N_10163,N_9135,N_9272);
nor U10164 (N_10164,N_9282,N_9442);
or U10165 (N_10165,N_9541,N_9497);
and U10166 (N_10166,N_9183,N_9530);
xor U10167 (N_10167,N_9037,N_9023);
or U10168 (N_10168,N_9640,N_9237);
nor U10169 (N_10169,N_9724,N_9521);
and U10170 (N_10170,N_9343,N_9675);
nor U10171 (N_10171,N_9725,N_9665);
and U10172 (N_10172,N_9127,N_9037);
and U10173 (N_10173,N_9021,N_9365);
nand U10174 (N_10174,N_9357,N_9603);
nand U10175 (N_10175,N_9441,N_9473);
nand U10176 (N_10176,N_9159,N_9234);
or U10177 (N_10177,N_9483,N_9115);
xor U10178 (N_10178,N_9591,N_9134);
nor U10179 (N_10179,N_9542,N_9300);
nand U10180 (N_10180,N_9583,N_9571);
or U10181 (N_10181,N_9709,N_9053);
or U10182 (N_10182,N_9670,N_9351);
or U10183 (N_10183,N_9465,N_9131);
xor U10184 (N_10184,N_9239,N_9506);
xor U10185 (N_10185,N_9580,N_9677);
and U10186 (N_10186,N_9438,N_9605);
xor U10187 (N_10187,N_9625,N_9147);
nor U10188 (N_10188,N_9476,N_9562);
nor U10189 (N_10189,N_9581,N_9512);
nor U10190 (N_10190,N_9044,N_9356);
nand U10191 (N_10191,N_9153,N_9606);
nor U10192 (N_10192,N_9659,N_9129);
or U10193 (N_10193,N_9474,N_9638);
or U10194 (N_10194,N_9311,N_9463);
nand U10195 (N_10195,N_9331,N_9349);
xor U10196 (N_10196,N_9339,N_9525);
nand U10197 (N_10197,N_9397,N_9174);
nand U10198 (N_10198,N_9563,N_9457);
and U10199 (N_10199,N_9304,N_9088);
or U10200 (N_10200,N_9491,N_9580);
xor U10201 (N_10201,N_9467,N_9612);
nand U10202 (N_10202,N_9213,N_9542);
nand U10203 (N_10203,N_9740,N_9299);
or U10204 (N_10204,N_9024,N_9158);
nand U10205 (N_10205,N_9163,N_9494);
or U10206 (N_10206,N_9582,N_9068);
xor U10207 (N_10207,N_9118,N_9197);
or U10208 (N_10208,N_9329,N_9226);
xnor U10209 (N_10209,N_9302,N_9099);
or U10210 (N_10210,N_9347,N_9015);
xor U10211 (N_10211,N_9310,N_9206);
or U10212 (N_10212,N_9147,N_9294);
or U10213 (N_10213,N_9576,N_9656);
nand U10214 (N_10214,N_9326,N_9122);
nand U10215 (N_10215,N_9458,N_9319);
nor U10216 (N_10216,N_9280,N_9336);
nand U10217 (N_10217,N_9472,N_9438);
and U10218 (N_10218,N_9222,N_9416);
nor U10219 (N_10219,N_9069,N_9649);
or U10220 (N_10220,N_9692,N_9052);
nand U10221 (N_10221,N_9031,N_9690);
nor U10222 (N_10222,N_9691,N_9109);
or U10223 (N_10223,N_9234,N_9422);
or U10224 (N_10224,N_9239,N_9708);
and U10225 (N_10225,N_9330,N_9511);
and U10226 (N_10226,N_9472,N_9591);
or U10227 (N_10227,N_9468,N_9027);
and U10228 (N_10228,N_9241,N_9523);
nand U10229 (N_10229,N_9744,N_9316);
and U10230 (N_10230,N_9392,N_9429);
xor U10231 (N_10231,N_9251,N_9149);
and U10232 (N_10232,N_9068,N_9092);
nor U10233 (N_10233,N_9061,N_9212);
nor U10234 (N_10234,N_9052,N_9151);
nand U10235 (N_10235,N_9673,N_9180);
nand U10236 (N_10236,N_9669,N_9074);
nand U10237 (N_10237,N_9486,N_9057);
or U10238 (N_10238,N_9630,N_9727);
nand U10239 (N_10239,N_9425,N_9524);
nand U10240 (N_10240,N_9277,N_9235);
xnor U10241 (N_10241,N_9390,N_9043);
xor U10242 (N_10242,N_9681,N_9238);
or U10243 (N_10243,N_9506,N_9659);
nor U10244 (N_10244,N_9261,N_9568);
nand U10245 (N_10245,N_9740,N_9628);
xor U10246 (N_10246,N_9269,N_9395);
nor U10247 (N_10247,N_9674,N_9646);
and U10248 (N_10248,N_9615,N_9533);
and U10249 (N_10249,N_9392,N_9051);
and U10250 (N_10250,N_9697,N_9194);
nor U10251 (N_10251,N_9424,N_9014);
nor U10252 (N_10252,N_9460,N_9591);
or U10253 (N_10253,N_9434,N_9433);
xnor U10254 (N_10254,N_9332,N_9370);
nor U10255 (N_10255,N_9717,N_9390);
nand U10256 (N_10256,N_9681,N_9409);
nand U10257 (N_10257,N_9734,N_9093);
or U10258 (N_10258,N_9348,N_9023);
nand U10259 (N_10259,N_9647,N_9545);
nand U10260 (N_10260,N_9001,N_9286);
and U10261 (N_10261,N_9322,N_9253);
or U10262 (N_10262,N_9739,N_9081);
nand U10263 (N_10263,N_9138,N_9121);
xnor U10264 (N_10264,N_9512,N_9532);
nand U10265 (N_10265,N_9535,N_9336);
and U10266 (N_10266,N_9011,N_9300);
or U10267 (N_10267,N_9563,N_9620);
or U10268 (N_10268,N_9727,N_9154);
or U10269 (N_10269,N_9033,N_9531);
nand U10270 (N_10270,N_9322,N_9397);
nand U10271 (N_10271,N_9232,N_9454);
nand U10272 (N_10272,N_9171,N_9346);
xnor U10273 (N_10273,N_9603,N_9000);
nand U10274 (N_10274,N_9038,N_9316);
xor U10275 (N_10275,N_9274,N_9080);
and U10276 (N_10276,N_9073,N_9466);
or U10277 (N_10277,N_9733,N_9439);
or U10278 (N_10278,N_9728,N_9381);
nor U10279 (N_10279,N_9335,N_9548);
or U10280 (N_10280,N_9075,N_9651);
or U10281 (N_10281,N_9293,N_9645);
and U10282 (N_10282,N_9133,N_9410);
xnor U10283 (N_10283,N_9085,N_9649);
nor U10284 (N_10284,N_9521,N_9281);
nor U10285 (N_10285,N_9120,N_9658);
nand U10286 (N_10286,N_9128,N_9240);
and U10287 (N_10287,N_9554,N_9419);
nor U10288 (N_10288,N_9227,N_9389);
xor U10289 (N_10289,N_9323,N_9194);
nor U10290 (N_10290,N_9718,N_9337);
xor U10291 (N_10291,N_9142,N_9717);
and U10292 (N_10292,N_9268,N_9749);
nand U10293 (N_10293,N_9621,N_9429);
nor U10294 (N_10294,N_9350,N_9708);
xnor U10295 (N_10295,N_9453,N_9213);
and U10296 (N_10296,N_9276,N_9181);
nand U10297 (N_10297,N_9196,N_9306);
or U10298 (N_10298,N_9121,N_9729);
or U10299 (N_10299,N_9278,N_9115);
nand U10300 (N_10300,N_9502,N_9485);
nor U10301 (N_10301,N_9277,N_9149);
xnor U10302 (N_10302,N_9323,N_9656);
nor U10303 (N_10303,N_9563,N_9658);
or U10304 (N_10304,N_9557,N_9230);
xor U10305 (N_10305,N_9633,N_9537);
nand U10306 (N_10306,N_9340,N_9331);
nand U10307 (N_10307,N_9716,N_9621);
nand U10308 (N_10308,N_9081,N_9460);
nand U10309 (N_10309,N_9024,N_9323);
or U10310 (N_10310,N_9388,N_9352);
nand U10311 (N_10311,N_9700,N_9439);
nor U10312 (N_10312,N_9139,N_9558);
or U10313 (N_10313,N_9544,N_9073);
and U10314 (N_10314,N_9655,N_9356);
and U10315 (N_10315,N_9281,N_9670);
xor U10316 (N_10316,N_9082,N_9527);
xnor U10317 (N_10317,N_9062,N_9693);
or U10318 (N_10318,N_9588,N_9400);
nand U10319 (N_10319,N_9695,N_9537);
and U10320 (N_10320,N_9495,N_9485);
nor U10321 (N_10321,N_9039,N_9163);
or U10322 (N_10322,N_9538,N_9685);
nand U10323 (N_10323,N_9100,N_9579);
nand U10324 (N_10324,N_9396,N_9515);
and U10325 (N_10325,N_9242,N_9104);
or U10326 (N_10326,N_9622,N_9139);
or U10327 (N_10327,N_9263,N_9616);
or U10328 (N_10328,N_9023,N_9382);
nor U10329 (N_10329,N_9469,N_9642);
nand U10330 (N_10330,N_9564,N_9406);
nor U10331 (N_10331,N_9311,N_9036);
xor U10332 (N_10332,N_9547,N_9024);
or U10333 (N_10333,N_9318,N_9465);
nor U10334 (N_10334,N_9037,N_9073);
or U10335 (N_10335,N_9041,N_9240);
nor U10336 (N_10336,N_9566,N_9233);
nand U10337 (N_10337,N_9260,N_9282);
nand U10338 (N_10338,N_9336,N_9705);
nand U10339 (N_10339,N_9347,N_9499);
nor U10340 (N_10340,N_9052,N_9092);
or U10341 (N_10341,N_9320,N_9492);
nor U10342 (N_10342,N_9244,N_9339);
and U10343 (N_10343,N_9127,N_9228);
xor U10344 (N_10344,N_9745,N_9503);
xor U10345 (N_10345,N_9320,N_9608);
xor U10346 (N_10346,N_9569,N_9708);
xnor U10347 (N_10347,N_9066,N_9122);
and U10348 (N_10348,N_9492,N_9486);
or U10349 (N_10349,N_9735,N_9668);
nand U10350 (N_10350,N_9371,N_9580);
and U10351 (N_10351,N_9352,N_9640);
nand U10352 (N_10352,N_9234,N_9319);
xor U10353 (N_10353,N_9560,N_9210);
xnor U10354 (N_10354,N_9640,N_9277);
xor U10355 (N_10355,N_9377,N_9058);
nor U10356 (N_10356,N_9328,N_9220);
nand U10357 (N_10357,N_9587,N_9577);
xor U10358 (N_10358,N_9123,N_9606);
or U10359 (N_10359,N_9499,N_9175);
or U10360 (N_10360,N_9102,N_9621);
and U10361 (N_10361,N_9695,N_9617);
and U10362 (N_10362,N_9181,N_9074);
and U10363 (N_10363,N_9708,N_9701);
and U10364 (N_10364,N_9526,N_9659);
and U10365 (N_10365,N_9518,N_9128);
and U10366 (N_10366,N_9180,N_9487);
and U10367 (N_10367,N_9286,N_9613);
or U10368 (N_10368,N_9009,N_9371);
nand U10369 (N_10369,N_9717,N_9701);
and U10370 (N_10370,N_9243,N_9241);
nor U10371 (N_10371,N_9077,N_9643);
and U10372 (N_10372,N_9424,N_9701);
and U10373 (N_10373,N_9320,N_9519);
xor U10374 (N_10374,N_9252,N_9494);
and U10375 (N_10375,N_9325,N_9609);
nand U10376 (N_10376,N_9587,N_9468);
xnor U10377 (N_10377,N_9299,N_9389);
nor U10378 (N_10378,N_9330,N_9408);
nor U10379 (N_10379,N_9187,N_9026);
and U10380 (N_10380,N_9220,N_9241);
xnor U10381 (N_10381,N_9181,N_9701);
xnor U10382 (N_10382,N_9091,N_9236);
nand U10383 (N_10383,N_9531,N_9225);
nand U10384 (N_10384,N_9190,N_9481);
or U10385 (N_10385,N_9702,N_9291);
or U10386 (N_10386,N_9460,N_9659);
xor U10387 (N_10387,N_9001,N_9676);
or U10388 (N_10388,N_9484,N_9266);
and U10389 (N_10389,N_9445,N_9714);
nand U10390 (N_10390,N_9346,N_9689);
nor U10391 (N_10391,N_9655,N_9565);
or U10392 (N_10392,N_9109,N_9240);
or U10393 (N_10393,N_9526,N_9148);
and U10394 (N_10394,N_9252,N_9566);
or U10395 (N_10395,N_9137,N_9148);
and U10396 (N_10396,N_9731,N_9578);
and U10397 (N_10397,N_9216,N_9643);
xnor U10398 (N_10398,N_9372,N_9645);
and U10399 (N_10399,N_9454,N_9448);
xnor U10400 (N_10400,N_9463,N_9485);
or U10401 (N_10401,N_9609,N_9511);
or U10402 (N_10402,N_9392,N_9434);
nor U10403 (N_10403,N_9287,N_9635);
xor U10404 (N_10404,N_9530,N_9591);
nor U10405 (N_10405,N_9638,N_9692);
or U10406 (N_10406,N_9086,N_9681);
nor U10407 (N_10407,N_9552,N_9067);
xor U10408 (N_10408,N_9303,N_9438);
nor U10409 (N_10409,N_9593,N_9479);
and U10410 (N_10410,N_9270,N_9131);
nor U10411 (N_10411,N_9039,N_9570);
and U10412 (N_10412,N_9309,N_9300);
nor U10413 (N_10413,N_9148,N_9572);
and U10414 (N_10414,N_9487,N_9251);
xnor U10415 (N_10415,N_9612,N_9550);
or U10416 (N_10416,N_9576,N_9579);
and U10417 (N_10417,N_9509,N_9263);
xnor U10418 (N_10418,N_9609,N_9449);
and U10419 (N_10419,N_9202,N_9175);
xnor U10420 (N_10420,N_9533,N_9134);
or U10421 (N_10421,N_9168,N_9299);
or U10422 (N_10422,N_9386,N_9191);
and U10423 (N_10423,N_9616,N_9509);
xnor U10424 (N_10424,N_9686,N_9314);
nor U10425 (N_10425,N_9096,N_9460);
xnor U10426 (N_10426,N_9512,N_9419);
nor U10427 (N_10427,N_9412,N_9059);
nor U10428 (N_10428,N_9171,N_9142);
or U10429 (N_10429,N_9333,N_9569);
or U10430 (N_10430,N_9642,N_9616);
nor U10431 (N_10431,N_9144,N_9570);
nand U10432 (N_10432,N_9124,N_9620);
nor U10433 (N_10433,N_9598,N_9238);
xnor U10434 (N_10434,N_9588,N_9305);
xnor U10435 (N_10435,N_9142,N_9330);
nand U10436 (N_10436,N_9352,N_9028);
and U10437 (N_10437,N_9747,N_9593);
or U10438 (N_10438,N_9731,N_9204);
and U10439 (N_10439,N_9702,N_9088);
or U10440 (N_10440,N_9315,N_9098);
and U10441 (N_10441,N_9014,N_9358);
nor U10442 (N_10442,N_9603,N_9574);
or U10443 (N_10443,N_9405,N_9658);
nand U10444 (N_10444,N_9088,N_9054);
and U10445 (N_10445,N_9382,N_9122);
xnor U10446 (N_10446,N_9075,N_9682);
xnor U10447 (N_10447,N_9008,N_9125);
nand U10448 (N_10448,N_9493,N_9039);
and U10449 (N_10449,N_9065,N_9650);
and U10450 (N_10450,N_9537,N_9606);
xor U10451 (N_10451,N_9689,N_9200);
xor U10452 (N_10452,N_9688,N_9720);
and U10453 (N_10453,N_9199,N_9446);
nor U10454 (N_10454,N_9731,N_9703);
nand U10455 (N_10455,N_9463,N_9071);
or U10456 (N_10456,N_9407,N_9265);
or U10457 (N_10457,N_9658,N_9535);
nor U10458 (N_10458,N_9436,N_9615);
nand U10459 (N_10459,N_9515,N_9478);
nor U10460 (N_10460,N_9651,N_9437);
nor U10461 (N_10461,N_9396,N_9416);
nor U10462 (N_10462,N_9325,N_9727);
nand U10463 (N_10463,N_9677,N_9736);
nor U10464 (N_10464,N_9499,N_9113);
xnor U10465 (N_10465,N_9276,N_9202);
nand U10466 (N_10466,N_9427,N_9304);
nand U10467 (N_10467,N_9002,N_9627);
or U10468 (N_10468,N_9226,N_9281);
xnor U10469 (N_10469,N_9491,N_9090);
and U10470 (N_10470,N_9655,N_9416);
nand U10471 (N_10471,N_9607,N_9639);
and U10472 (N_10472,N_9055,N_9097);
nor U10473 (N_10473,N_9625,N_9645);
and U10474 (N_10474,N_9722,N_9720);
xnor U10475 (N_10475,N_9437,N_9417);
nand U10476 (N_10476,N_9042,N_9662);
xnor U10477 (N_10477,N_9643,N_9686);
nor U10478 (N_10478,N_9684,N_9486);
or U10479 (N_10479,N_9394,N_9591);
nor U10480 (N_10480,N_9744,N_9088);
nand U10481 (N_10481,N_9628,N_9256);
nand U10482 (N_10482,N_9723,N_9299);
or U10483 (N_10483,N_9306,N_9366);
and U10484 (N_10484,N_9662,N_9050);
nor U10485 (N_10485,N_9374,N_9231);
nand U10486 (N_10486,N_9161,N_9602);
xor U10487 (N_10487,N_9569,N_9293);
and U10488 (N_10488,N_9541,N_9509);
xor U10489 (N_10489,N_9703,N_9005);
and U10490 (N_10490,N_9042,N_9467);
and U10491 (N_10491,N_9293,N_9086);
nor U10492 (N_10492,N_9136,N_9002);
nor U10493 (N_10493,N_9590,N_9051);
and U10494 (N_10494,N_9338,N_9708);
and U10495 (N_10495,N_9224,N_9321);
or U10496 (N_10496,N_9330,N_9179);
nor U10497 (N_10497,N_9557,N_9061);
xor U10498 (N_10498,N_9472,N_9338);
xnor U10499 (N_10499,N_9726,N_9400);
nand U10500 (N_10500,N_9929,N_10095);
nand U10501 (N_10501,N_10238,N_9939);
xor U10502 (N_10502,N_10053,N_10271);
and U10503 (N_10503,N_10291,N_9981);
and U10504 (N_10504,N_10314,N_10218);
nand U10505 (N_10505,N_10120,N_10299);
nand U10506 (N_10506,N_10436,N_10411);
nand U10507 (N_10507,N_9966,N_10270);
xnor U10508 (N_10508,N_10367,N_9935);
nor U10509 (N_10509,N_10173,N_10104);
and U10510 (N_10510,N_9821,N_9777);
and U10511 (N_10511,N_10319,N_10031);
nand U10512 (N_10512,N_9835,N_10106);
nor U10513 (N_10513,N_10161,N_10105);
nand U10514 (N_10514,N_10492,N_10004);
xor U10515 (N_10515,N_10341,N_9897);
and U10516 (N_10516,N_9754,N_10178);
nor U10517 (N_10517,N_10442,N_10060);
or U10518 (N_10518,N_9797,N_10466);
nor U10519 (N_10519,N_10136,N_10024);
xnor U10520 (N_10520,N_10322,N_10303);
nand U10521 (N_10521,N_10007,N_9758);
and U10522 (N_10522,N_10429,N_9903);
or U10523 (N_10523,N_10497,N_10108);
nand U10524 (N_10524,N_10203,N_9996);
nor U10525 (N_10525,N_10126,N_10052);
or U10526 (N_10526,N_10034,N_10254);
or U10527 (N_10527,N_9817,N_10283);
nand U10528 (N_10528,N_9948,N_10239);
nand U10529 (N_10529,N_9826,N_9963);
or U10530 (N_10530,N_9949,N_10424);
nor U10531 (N_10531,N_10428,N_10302);
and U10532 (N_10532,N_10490,N_9856);
nor U10533 (N_10533,N_10174,N_10018);
nand U10534 (N_10534,N_10032,N_10110);
and U10535 (N_10535,N_9863,N_9848);
xnor U10536 (N_10536,N_9904,N_10471);
and U10537 (N_10537,N_10495,N_10130);
xor U10538 (N_10538,N_10047,N_9831);
or U10539 (N_10539,N_9936,N_9919);
or U10540 (N_10540,N_10244,N_9973);
and U10541 (N_10541,N_10453,N_9778);
xnor U10542 (N_10542,N_10037,N_10125);
or U10543 (N_10543,N_10099,N_9887);
xnor U10544 (N_10544,N_10366,N_10134);
or U10545 (N_10545,N_10335,N_9814);
xor U10546 (N_10546,N_10012,N_10028);
or U10547 (N_10547,N_10340,N_10305);
or U10548 (N_10548,N_10432,N_9961);
xnor U10549 (N_10549,N_10371,N_9847);
and U10550 (N_10550,N_10059,N_10336);
nand U10551 (N_10551,N_10229,N_10222);
nand U10552 (N_10552,N_9783,N_9813);
nor U10553 (N_10553,N_10245,N_10397);
and U10554 (N_10554,N_10141,N_9909);
nand U10555 (N_10555,N_10478,N_9823);
and U10556 (N_10556,N_9871,N_10309);
nand U10557 (N_10557,N_10111,N_10073);
nor U10558 (N_10558,N_10396,N_10273);
xor U10559 (N_10559,N_10026,N_10035);
or U10560 (N_10560,N_9851,N_9832);
xor U10561 (N_10561,N_10437,N_9750);
or U10562 (N_10562,N_10472,N_9965);
or U10563 (N_10563,N_10454,N_10042);
or U10564 (N_10564,N_10065,N_10282);
nor U10565 (N_10565,N_10483,N_10040);
or U10566 (N_10566,N_10368,N_10008);
xnor U10567 (N_10567,N_9922,N_10207);
xnor U10568 (N_10568,N_10021,N_10473);
xnor U10569 (N_10569,N_10118,N_9938);
nand U10570 (N_10570,N_10150,N_10094);
nand U10571 (N_10571,N_9842,N_10285);
nor U10572 (N_10572,N_9877,N_10081);
nand U10573 (N_10573,N_10382,N_9769);
nor U10574 (N_10574,N_9844,N_10000);
and U10575 (N_10575,N_10117,N_10277);
or U10576 (N_10576,N_10410,N_10345);
and U10577 (N_10577,N_10433,N_9846);
nor U10578 (N_10578,N_10116,N_10370);
and U10579 (N_10579,N_9798,N_9980);
nor U10580 (N_10580,N_10189,N_10326);
nor U10581 (N_10581,N_9978,N_10082);
or U10582 (N_10582,N_9837,N_10164);
xnor U10583 (N_10583,N_9918,N_10499);
or U10584 (N_10584,N_9879,N_10293);
nor U10585 (N_10585,N_10360,N_10158);
and U10586 (N_10586,N_10405,N_10233);
nor U10587 (N_10587,N_10496,N_9959);
nand U10588 (N_10588,N_9776,N_10206);
xnor U10589 (N_10589,N_10331,N_10086);
or U10590 (N_10590,N_10284,N_9818);
nor U10591 (N_10591,N_10261,N_9943);
nor U10592 (N_10592,N_9795,N_9942);
nor U10593 (N_10593,N_10133,N_10043);
nand U10594 (N_10594,N_10482,N_10121);
and U10595 (N_10595,N_9977,N_9906);
or U10596 (N_10596,N_9808,N_9924);
or U10597 (N_10597,N_10249,N_10051);
and U10598 (N_10598,N_10219,N_9881);
or U10599 (N_10599,N_10132,N_10407);
nand U10600 (N_10600,N_10049,N_9820);
nand U10601 (N_10601,N_10301,N_10363);
nor U10602 (N_10602,N_10228,N_10395);
nor U10603 (N_10603,N_10276,N_10061);
and U10604 (N_10604,N_9896,N_10098);
xor U10605 (N_10605,N_9912,N_10379);
nor U10606 (N_10606,N_10421,N_10179);
nand U10607 (N_10607,N_10063,N_9993);
xor U10608 (N_10608,N_10115,N_10294);
nor U10609 (N_10609,N_9915,N_9945);
and U10610 (N_10610,N_10330,N_9852);
and U10611 (N_10611,N_10202,N_10055);
and U10612 (N_10612,N_10214,N_9811);
xor U10613 (N_10613,N_10237,N_10002);
nor U10614 (N_10614,N_10387,N_10304);
or U10615 (N_10615,N_10274,N_10071);
nor U10616 (N_10616,N_10427,N_9889);
or U10617 (N_10617,N_9792,N_9902);
nor U10618 (N_10618,N_10262,N_10474);
xor U10619 (N_10619,N_10230,N_10327);
nor U10620 (N_10620,N_9884,N_10090);
nor U10621 (N_10621,N_9999,N_10242);
xnor U10622 (N_10622,N_10259,N_10414);
nand U10623 (N_10623,N_10074,N_9766);
and U10624 (N_10624,N_9921,N_10165);
xnor U10625 (N_10625,N_9762,N_10250);
or U10626 (N_10626,N_9997,N_9885);
xnor U10627 (N_10627,N_9774,N_10441);
xor U10628 (N_10628,N_10143,N_9829);
nor U10629 (N_10629,N_9753,N_10085);
nand U10630 (N_10630,N_10374,N_9869);
nor U10631 (N_10631,N_10459,N_9974);
xor U10632 (N_10632,N_10257,N_9757);
xor U10633 (N_10633,N_9891,N_10413);
and U10634 (N_10634,N_10306,N_10369);
or U10635 (N_10635,N_10019,N_10344);
and U10636 (N_10636,N_10193,N_9895);
or U10637 (N_10637,N_10039,N_9971);
nand U10638 (N_10638,N_10223,N_10362);
nor U10639 (N_10639,N_10236,N_10464);
or U10640 (N_10640,N_9901,N_10440);
or U10641 (N_10641,N_10131,N_10080);
nor U10642 (N_10642,N_10321,N_10112);
nor U10643 (N_10643,N_10220,N_9861);
and U10644 (N_10644,N_10191,N_10253);
nor U10645 (N_10645,N_9953,N_10465);
nand U10646 (N_10646,N_10172,N_10169);
nand U10647 (N_10647,N_9952,N_9838);
and U10648 (N_10648,N_9768,N_10449);
xor U10649 (N_10649,N_9976,N_10353);
nor U10650 (N_10650,N_9812,N_10455);
nand U10651 (N_10651,N_9763,N_10408);
xor U10652 (N_10652,N_10488,N_9970);
xnor U10653 (N_10653,N_9770,N_10184);
and U10654 (N_10654,N_10114,N_10243);
nor U10655 (N_10655,N_10313,N_9805);
or U10656 (N_10656,N_9752,N_10025);
nand U10657 (N_10657,N_9911,N_9969);
xor U10658 (N_10658,N_10444,N_10481);
and U10659 (N_10659,N_10351,N_10287);
and U10660 (N_10660,N_9860,N_9800);
xor U10661 (N_10661,N_9975,N_9940);
and U10662 (N_10662,N_10016,N_10188);
nand U10663 (N_10663,N_9991,N_9850);
and U10664 (N_10664,N_9926,N_9866);
and U10665 (N_10665,N_9791,N_10140);
nand U10666 (N_10666,N_10477,N_10372);
nand U10667 (N_10667,N_10289,N_9986);
nor U10668 (N_10668,N_10102,N_10357);
or U10669 (N_10669,N_9937,N_9773);
nor U10670 (N_10670,N_10390,N_10339);
nand U10671 (N_10671,N_10355,N_10352);
xor U10672 (N_10672,N_9990,N_10247);
nand U10673 (N_10673,N_9873,N_9755);
xnor U10674 (N_10674,N_10167,N_10057);
xor U10675 (N_10675,N_9893,N_10468);
xor U10676 (N_10676,N_9931,N_9916);
nor U10677 (N_10677,N_10358,N_10388);
or U10678 (N_10678,N_9853,N_10045);
or U10679 (N_10679,N_9907,N_10297);
xnor U10680 (N_10680,N_10148,N_9886);
nor U10681 (N_10681,N_10423,N_10181);
or U10682 (N_10682,N_10248,N_9964);
and U10683 (N_10683,N_9992,N_10256);
nor U10684 (N_10684,N_9781,N_9767);
and U10685 (N_10685,N_10268,N_10011);
nand U10686 (N_10686,N_10146,N_9888);
or U10687 (N_10687,N_10347,N_10056);
nand U10688 (N_10688,N_10275,N_10486);
or U10689 (N_10689,N_10152,N_9958);
and U10690 (N_10690,N_9979,N_10175);
xnor U10691 (N_10691,N_9960,N_10232);
and U10692 (N_10692,N_9878,N_9804);
nor U10693 (N_10693,N_10216,N_9859);
nor U10694 (N_10694,N_9807,N_9787);
and U10695 (N_10695,N_10192,N_9932);
xnor U10696 (N_10696,N_9790,N_10231);
and U10697 (N_10697,N_10096,N_10354);
nor U10698 (N_10698,N_10068,N_10381);
xor U10699 (N_10699,N_9870,N_10348);
and U10700 (N_10700,N_10420,N_10097);
and U10701 (N_10701,N_9855,N_9782);
and U10702 (N_10702,N_10089,N_9968);
xnor U10703 (N_10703,N_10070,N_10211);
or U10704 (N_10704,N_10476,N_10401);
nor U10705 (N_10705,N_10320,N_10123);
nand U10706 (N_10706,N_10460,N_10194);
and U10707 (N_10707,N_9930,N_10365);
or U10708 (N_10708,N_10014,N_9925);
xor U10709 (N_10709,N_10196,N_10392);
or U10710 (N_10710,N_10448,N_10462);
and U10711 (N_10711,N_9756,N_10487);
xor U10712 (N_10712,N_10350,N_10258);
and U10713 (N_10713,N_10109,N_9772);
and U10714 (N_10714,N_10267,N_9786);
nand U10715 (N_10715,N_10463,N_9809);
nand U10716 (N_10716,N_9806,N_10139);
nand U10717 (N_10717,N_9857,N_10255);
and U10718 (N_10718,N_10416,N_10290);
and U10719 (N_10719,N_10318,N_10075);
or U10720 (N_10720,N_10198,N_9880);
xnor U10721 (N_10721,N_9882,N_9955);
nor U10722 (N_10722,N_10168,N_10020);
and U10723 (N_10723,N_10263,N_10295);
xnor U10724 (N_10724,N_10443,N_10447);
nand U10725 (N_10725,N_9956,N_9815);
xnor U10726 (N_10726,N_10226,N_9983);
and U10727 (N_10727,N_9914,N_10398);
and U10728 (N_10728,N_10457,N_10029);
and U10729 (N_10729,N_10378,N_10399);
nand U10730 (N_10730,N_10013,N_10338);
xnor U10731 (N_10731,N_10389,N_9894);
nand U10732 (N_10732,N_9876,N_9780);
nand U10733 (N_10733,N_10402,N_10485);
xnor U10734 (N_10734,N_10489,N_10186);
nor U10735 (N_10735,N_10006,N_10195);
nor U10736 (N_10736,N_9789,N_10434);
nand U10737 (N_10737,N_10093,N_9854);
and U10738 (N_10738,N_10470,N_9785);
nor U10739 (N_10739,N_10342,N_10252);
nor U10740 (N_10740,N_10323,N_10380);
nand U10741 (N_10741,N_10298,N_10145);
nand U10742 (N_10742,N_10494,N_10361);
or U10743 (N_10743,N_10113,N_10312);
and U10744 (N_10744,N_10182,N_9995);
and U10745 (N_10745,N_9927,N_10394);
or U10746 (N_10746,N_10062,N_10185);
nor U10747 (N_10747,N_10135,N_9984);
nor U10748 (N_10748,N_10155,N_10403);
nor U10749 (N_10749,N_10446,N_10337);
nand U10750 (N_10750,N_10176,N_9843);
nor U10751 (N_10751,N_9794,N_10425);
and U10752 (N_10752,N_10180,N_10046);
nor U10753 (N_10753,N_10419,N_9923);
or U10754 (N_10754,N_9827,N_10171);
xor U10755 (N_10755,N_10393,N_9788);
nor U10756 (N_10756,N_10159,N_10296);
nor U10757 (N_10757,N_9764,N_10439);
nand U10758 (N_10758,N_10023,N_9908);
nor U10759 (N_10759,N_10451,N_10151);
or U10760 (N_10760,N_10078,N_10484);
xnor U10761 (N_10761,N_10017,N_9849);
xnor U10762 (N_10762,N_9819,N_10156);
xor U10763 (N_10763,N_10149,N_10260);
nand U10764 (N_10764,N_10456,N_10069);
or U10765 (N_10765,N_9985,N_10406);
nor U10766 (N_10766,N_10317,N_9858);
and U10767 (N_10767,N_10376,N_10328);
or U10768 (N_10768,N_10458,N_10278);
and U10769 (N_10769,N_10409,N_9989);
or U10770 (N_10770,N_9839,N_10103);
xnor U10771 (N_10771,N_10137,N_9957);
or U10772 (N_10772,N_10050,N_10445);
nor U10773 (N_10773,N_10162,N_10072);
xor U10774 (N_10774,N_9962,N_10240);
nor U10775 (N_10775,N_9892,N_10225);
nor U10776 (N_10776,N_9913,N_9868);
and U10777 (N_10777,N_10087,N_10431);
nand U10778 (N_10778,N_9982,N_10030);
or U10779 (N_10779,N_10307,N_10166);
or U10780 (N_10780,N_9920,N_9988);
and U10781 (N_10781,N_10479,N_9874);
xor U10782 (N_10782,N_10221,N_10119);
and U10783 (N_10783,N_10038,N_10415);
and U10784 (N_10784,N_10329,N_10154);
nand U10785 (N_10785,N_9761,N_10153);
nor U10786 (N_10786,N_9900,N_9801);
or U10787 (N_10787,N_10107,N_10127);
or U10788 (N_10788,N_10215,N_9841);
nor U10789 (N_10789,N_9994,N_10187);
and U10790 (N_10790,N_10333,N_9875);
and U10791 (N_10791,N_10491,N_10067);
and U10792 (N_10792,N_10054,N_9824);
xor U10793 (N_10793,N_10022,N_9830);
and U10794 (N_10794,N_9898,N_9765);
or U10795 (N_10795,N_9917,N_10101);
nand U10796 (N_10796,N_10044,N_10292);
xnor U10797 (N_10797,N_10266,N_9864);
nand U10798 (N_10798,N_10197,N_10160);
or U10799 (N_10799,N_10005,N_10100);
nor U10800 (N_10800,N_9967,N_10404);
nand U10801 (N_10801,N_10058,N_10269);
nand U10802 (N_10802,N_10430,N_10264);
nor U10803 (N_10803,N_10426,N_10217);
and U10804 (N_10804,N_10009,N_9751);
nand U10805 (N_10805,N_9834,N_9796);
and U10806 (N_10806,N_10015,N_10480);
or U10807 (N_10807,N_10359,N_9828);
and U10808 (N_10808,N_10315,N_9934);
xnor U10809 (N_10809,N_9793,N_10373);
nand U10810 (N_10810,N_10375,N_10208);
nand U10811 (N_10811,N_10084,N_10467);
and U10812 (N_10812,N_10346,N_10079);
nand U10813 (N_10813,N_10204,N_9905);
xor U10814 (N_10814,N_10310,N_10205);
or U10815 (N_10815,N_10251,N_10241);
or U10816 (N_10816,N_10128,N_9810);
nor U10817 (N_10817,N_10147,N_10212);
and U10818 (N_10818,N_10001,N_9867);
xnor U10819 (N_10819,N_9872,N_10400);
xnor U10820 (N_10820,N_9803,N_10364);
or U10821 (N_10821,N_10036,N_10324);
or U10822 (N_10822,N_10234,N_10332);
or U10823 (N_10823,N_10209,N_9910);
or U10824 (N_10824,N_10163,N_9862);
nor U10825 (N_10825,N_9845,N_10475);
nand U10826 (N_10826,N_10048,N_10124);
xor U10827 (N_10827,N_10088,N_10138);
or U10828 (N_10828,N_10349,N_10300);
nand U10829 (N_10829,N_10201,N_10391);
xnor U10830 (N_10830,N_9775,N_9928);
or U10831 (N_10831,N_10077,N_10177);
nand U10832 (N_10832,N_10272,N_10418);
or U10833 (N_10833,N_9779,N_10385);
nand U10834 (N_10834,N_10157,N_10288);
xnor U10835 (N_10835,N_10386,N_10210);
or U10836 (N_10836,N_9816,N_9836);
nand U10837 (N_10837,N_9899,N_10311);
nor U10838 (N_10838,N_10450,N_9951);
nor U10839 (N_10839,N_10027,N_9771);
nand U10840 (N_10840,N_10199,N_9890);
nand U10841 (N_10841,N_10265,N_10384);
or U10842 (N_10842,N_10066,N_10200);
and U10843 (N_10843,N_9987,N_10417);
nand U10844 (N_10844,N_10144,N_9946);
xor U10845 (N_10845,N_9760,N_9883);
nand U10846 (N_10846,N_9933,N_10213);
or U10847 (N_10847,N_10003,N_10235);
and U10848 (N_10848,N_10325,N_10041);
nand U10849 (N_10849,N_10170,N_10076);
or U10850 (N_10850,N_9954,N_9825);
or U10851 (N_10851,N_10356,N_10122);
xor U10852 (N_10852,N_10308,N_9944);
or U10853 (N_10853,N_10142,N_10461);
or U10854 (N_10854,N_10227,N_10422);
and U10855 (N_10855,N_10190,N_9799);
or U10856 (N_10856,N_9865,N_10246);
and U10857 (N_10857,N_9947,N_10091);
nor U10858 (N_10858,N_10498,N_10435);
and U10859 (N_10859,N_10343,N_9802);
and U10860 (N_10860,N_10064,N_10183);
nor U10861 (N_10861,N_10224,N_10281);
xnor U10862 (N_10862,N_9941,N_10279);
nor U10863 (N_10863,N_9972,N_10493);
or U10864 (N_10864,N_10316,N_10377);
or U10865 (N_10865,N_9950,N_10469);
nor U10866 (N_10866,N_9840,N_10383);
nand U10867 (N_10867,N_10010,N_10280);
and U10868 (N_10868,N_10033,N_10412);
nand U10869 (N_10869,N_10092,N_9784);
nand U10870 (N_10870,N_9833,N_10129);
nand U10871 (N_10871,N_9998,N_9822);
xor U10872 (N_10872,N_10083,N_9759);
xnor U10873 (N_10873,N_10452,N_10334);
nor U10874 (N_10874,N_10286,N_10438);
nand U10875 (N_10875,N_10214,N_9999);
or U10876 (N_10876,N_10183,N_10090);
or U10877 (N_10877,N_10111,N_10080);
xor U10878 (N_10878,N_10066,N_10040);
or U10879 (N_10879,N_9787,N_10291);
xnor U10880 (N_10880,N_10410,N_9759);
nor U10881 (N_10881,N_10179,N_9986);
or U10882 (N_10882,N_9837,N_10470);
or U10883 (N_10883,N_9813,N_10372);
nor U10884 (N_10884,N_9861,N_9994);
and U10885 (N_10885,N_10138,N_10272);
nand U10886 (N_10886,N_9849,N_10163);
nor U10887 (N_10887,N_10358,N_10492);
and U10888 (N_10888,N_10093,N_10436);
and U10889 (N_10889,N_10342,N_10197);
xnor U10890 (N_10890,N_10195,N_10085);
xnor U10891 (N_10891,N_9950,N_10009);
nand U10892 (N_10892,N_9993,N_10279);
or U10893 (N_10893,N_9836,N_9838);
and U10894 (N_10894,N_10186,N_9841);
and U10895 (N_10895,N_10440,N_10005);
or U10896 (N_10896,N_10456,N_9755);
and U10897 (N_10897,N_10072,N_10300);
nor U10898 (N_10898,N_10341,N_10091);
nor U10899 (N_10899,N_10444,N_9928);
xnor U10900 (N_10900,N_9858,N_10159);
nor U10901 (N_10901,N_10435,N_10476);
nand U10902 (N_10902,N_10321,N_10361);
xor U10903 (N_10903,N_9766,N_10017);
nand U10904 (N_10904,N_10012,N_9818);
and U10905 (N_10905,N_10195,N_10429);
or U10906 (N_10906,N_10217,N_10338);
or U10907 (N_10907,N_10268,N_10384);
or U10908 (N_10908,N_10127,N_10405);
nand U10909 (N_10909,N_10424,N_10117);
nand U10910 (N_10910,N_9833,N_10394);
xor U10911 (N_10911,N_10204,N_10258);
and U10912 (N_10912,N_9859,N_10070);
nor U10913 (N_10913,N_10328,N_9944);
nor U10914 (N_10914,N_9790,N_10375);
xor U10915 (N_10915,N_9902,N_10326);
or U10916 (N_10916,N_9999,N_9894);
nand U10917 (N_10917,N_9875,N_10061);
or U10918 (N_10918,N_9852,N_10190);
or U10919 (N_10919,N_10006,N_10366);
nor U10920 (N_10920,N_9951,N_10339);
xnor U10921 (N_10921,N_10135,N_10109);
xnor U10922 (N_10922,N_10171,N_9896);
and U10923 (N_10923,N_10279,N_9940);
or U10924 (N_10924,N_10202,N_10424);
nand U10925 (N_10925,N_10216,N_9905);
xnor U10926 (N_10926,N_10161,N_10137);
or U10927 (N_10927,N_10132,N_10392);
or U10928 (N_10928,N_10211,N_9831);
nand U10929 (N_10929,N_10320,N_9954);
or U10930 (N_10930,N_10245,N_10384);
nor U10931 (N_10931,N_10325,N_10218);
and U10932 (N_10932,N_9973,N_9839);
and U10933 (N_10933,N_10119,N_10015);
xnor U10934 (N_10934,N_9804,N_10043);
nand U10935 (N_10935,N_9977,N_10386);
and U10936 (N_10936,N_9854,N_10201);
xor U10937 (N_10937,N_10153,N_10130);
nor U10938 (N_10938,N_10189,N_9766);
nand U10939 (N_10939,N_10261,N_10453);
xnor U10940 (N_10940,N_9876,N_9866);
and U10941 (N_10941,N_9775,N_10361);
and U10942 (N_10942,N_9886,N_10274);
nor U10943 (N_10943,N_9949,N_10481);
or U10944 (N_10944,N_10342,N_10322);
nand U10945 (N_10945,N_10247,N_9936);
or U10946 (N_10946,N_10189,N_10228);
nor U10947 (N_10947,N_9781,N_10467);
and U10948 (N_10948,N_10179,N_10103);
xnor U10949 (N_10949,N_9820,N_10318);
nor U10950 (N_10950,N_9798,N_10499);
nand U10951 (N_10951,N_10266,N_9887);
and U10952 (N_10952,N_9778,N_9827);
or U10953 (N_10953,N_10269,N_10053);
xnor U10954 (N_10954,N_9808,N_10440);
and U10955 (N_10955,N_9897,N_9789);
nand U10956 (N_10956,N_10054,N_10332);
nand U10957 (N_10957,N_10233,N_10092);
xnor U10958 (N_10958,N_9960,N_10367);
and U10959 (N_10959,N_10396,N_10193);
and U10960 (N_10960,N_10463,N_9817);
nor U10961 (N_10961,N_9842,N_10138);
and U10962 (N_10962,N_9831,N_10476);
nand U10963 (N_10963,N_10476,N_9843);
or U10964 (N_10964,N_10369,N_9975);
or U10965 (N_10965,N_10251,N_10143);
and U10966 (N_10966,N_9875,N_9825);
xor U10967 (N_10967,N_10429,N_10478);
and U10968 (N_10968,N_10183,N_9864);
and U10969 (N_10969,N_9865,N_10239);
or U10970 (N_10970,N_10490,N_9771);
or U10971 (N_10971,N_10057,N_10392);
xor U10972 (N_10972,N_9975,N_10395);
and U10973 (N_10973,N_9969,N_10372);
nor U10974 (N_10974,N_10498,N_9901);
xor U10975 (N_10975,N_9876,N_9760);
nand U10976 (N_10976,N_10080,N_10092);
nand U10977 (N_10977,N_9759,N_10440);
nand U10978 (N_10978,N_10021,N_10477);
xnor U10979 (N_10979,N_9824,N_10301);
nand U10980 (N_10980,N_10213,N_9786);
or U10981 (N_10981,N_10213,N_9973);
or U10982 (N_10982,N_10121,N_10053);
xnor U10983 (N_10983,N_9939,N_10274);
and U10984 (N_10984,N_10495,N_10499);
xor U10985 (N_10985,N_10076,N_10314);
xor U10986 (N_10986,N_10323,N_10319);
and U10987 (N_10987,N_10093,N_10328);
or U10988 (N_10988,N_10476,N_10266);
xnor U10989 (N_10989,N_10239,N_10037);
nand U10990 (N_10990,N_10435,N_10282);
nand U10991 (N_10991,N_9795,N_10061);
and U10992 (N_10992,N_9856,N_10431);
or U10993 (N_10993,N_10031,N_10132);
nand U10994 (N_10994,N_10271,N_10161);
or U10995 (N_10995,N_10292,N_9961);
nor U10996 (N_10996,N_10334,N_9976);
xnor U10997 (N_10997,N_10341,N_10335);
and U10998 (N_10998,N_10262,N_10000);
nor U10999 (N_10999,N_10222,N_9770);
nor U11000 (N_11000,N_10118,N_10158);
xnor U11001 (N_11001,N_10104,N_10444);
and U11002 (N_11002,N_10454,N_10397);
and U11003 (N_11003,N_10293,N_10260);
xor U11004 (N_11004,N_10301,N_10358);
nor U11005 (N_11005,N_10472,N_10386);
xnor U11006 (N_11006,N_9860,N_10067);
nor U11007 (N_11007,N_10057,N_10050);
or U11008 (N_11008,N_10382,N_10439);
and U11009 (N_11009,N_10389,N_10430);
xnor U11010 (N_11010,N_10379,N_10434);
nand U11011 (N_11011,N_9892,N_10240);
nor U11012 (N_11012,N_10030,N_10253);
nor U11013 (N_11013,N_10059,N_10368);
and U11014 (N_11014,N_10018,N_10325);
nand U11015 (N_11015,N_10234,N_10181);
and U11016 (N_11016,N_10067,N_10287);
and U11017 (N_11017,N_10314,N_10486);
xnor U11018 (N_11018,N_10314,N_10222);
nor U11019 (N_11019,N_10129,N_10406);
or U11020 (N_11020,N_10367,N_9916);
and U11021 (N_11021,N_10303,N_10030);
nand U11022 (N_11022,N_10145,N_10173);
and U11023 (N_11023,N_9891,N_10072);
nor U11024 (N_11024,N_10318,N_10280);
nand U11025 (N_11025,N_9989,N_10074);
or U11026 (N_11026,N_10139,N_9981);
and U11027 (N_11027,N_9787,N_10350);
or U11028 (N_11028,N_10359,N_10234);
nand U11029 (N_11029,N_10249,N_9807);
xnor U11030 (N_11030,N_9826,N_10185);
xnor U11031 (N_11031,N_10418,N_9780);
and U11032 (N_11032,N_10110,N_10475);
nand U11033 (N_11033,N_10291,N_10101);
nor U11034 (N_11034,N_10148,N_9788);
or U11035 (N_11035,N_10036,N_10071);
or U11036 (N_11036,N_10416,N_10085);
nand U11037 (N_11037,N_9923,N_9788);
xnor U11038 (N_11038,N_10458,N_9931);
and U11039 (N_11039,N_9972,N_10065);
xor U11040 (N_11040,N_9988,N_10011);
xor U11041 (N_11041,N_10200,N_9870);
nor U11042 (N_11042,N_10147,N_10406);
or U11043 (N_11043,N_9966,N_10097);
or U11044 (N_11044,N_10221,N_9940);
nand U11045 (N_11045,N_10304,N_10389);
nor U11046 (N_11046,N_9761,N_10486);
or U11047 (N_11047,N_10063,N_9840);
nand U11048 (N_11048,N_10107,N_9786);
or U11049 (N_11049,N_10214,N_9895);
nor U11050 (N_11050,N_10191,N_10283);
or U11051 (N_11051,N_10487,N_10486);
xor U11052 (N_11052,N_10170,N_9799);
or U11053 (N_11053,N_10324,N_10241);
nand U11054 (N_11054,N_10270,N_9812);
and U11055 (N_11055,N_10112,N_10464);
and U11056 (N_11056,N_10099,N_9949);
xor U11057 (N_11057,N_9960,N_10125);
xnor U11058 (N_11058,N_9800,N_10163);
or U11059 (N_11059,N_9820,N_9802);
or U11060 (N_11060,N_10084,N_9879);
and U11061 (N_11061,N_10247,N_9772);
or U11062 (N_11062,N_10216,N_10072);
nand U11063 (N_11063,N_10297,N_10429);
nor U11064 (N_11064,N_9959,N_9988);
and U11065 (N_11065,N_10264,N_10162);
nor U11066 (N_11066,N_10388,N_10265);
and U11067 (N_11067,N_9811,N_10235);
nand U11068 (N_11068,N_10112,N_9974);
xor U11069 (N_11069,N_10043,N_10134);
nor U11070 (N_11070,N_10066,N_9808);
nor U11071 (N_11071,N_10337,N_9845);
or U11072 (N_11072,N_9821,N_10319);
or U11073 (N_11073,N_10154,N_9806);
nand U11074 (N_11074,N_10190,N_9804);
nor U11075 (N_11075,N_10165,N_10429);
nand U11076 (N_11076,N_10111,N_10450);
and U11077 (N_11077,N_10413,N_10072);
nand U11078 (N_11078,N_9915,N_10393);
xnor U11079 (N_11079,N_9832,N_10454);
or U11080 (N_11080,N_10478,N_10165);
nand U11081 (N_11081,N_10229,N_10019);
nor U11082 (N_11082,N_10355,N_9805);
and U11083 (N_11083,N_9899,N_9883);
and U11084 (N_11084,N_10040,N_9773);
or U11085 (N_11085,N_9840,N_9914);
nor U11086 (N_11086,N_9970,N_10166);
nor U11087 (N_11087,N_9974,N_10078);
nor U11088 (N_11088,N_10477,N_10257);
nor U11089 (N_11089,N_9834,N_10188);
xnor U11090 (N_11090,N_10333,N_10298);
xor U11091 (N_11091,N_10318,N_10271);
and U11092 (N_11092,N_9788,N_9888);
and U11093 (N_11093,N_10408,N_10015);
and U11094 (N_11094,N_10412,N_10392);
xnor U11095 (N_11095,N_10386,N_10345);
nand U11096 (N_11096,N_10049,N_10494);
or U11097 (N_11097,N_10024,N_9765);
xnor U11098 (N_11098,N_10258,N_9854);
and U11099 (N_11099,N_9801,N_10389);
nor U11100 (N_11100,N_9786,N_10039);
and U11101 (N_11101,N_10190,N_10351);
nor U11102 (N_11102,N_9776,N_9945);
xor U11103 (N_11103,N_10321,N_9822);
xnor U11104 (N_11104,N_10071,N_10314);
and U11105 (N_11105,N_10406,N_10029);
and U11106 (N_11106,N_10019,N_9775);
and U11107 (N_11107,N_10112,N_9782);
nand U11108 (N_11108,N_9776,N_9789);
or U11109 (N_11109,N_10346,N_10212);
or U11110 (N_11110,N_9766,N_9774);
nand U11111 (N_11111,N_10302,N_10497);
xnor U11112 (N_11112,N_10096,N_10448);
nor U11113 (N_11113,N_10269,N_9818);
nand U11114 (N_11114,N_10310,N_9916);
and U11115 (N_11115,N_10342,N_9934);
and U11116 (N_11116,N_10072,N_10247);
xor U11117 (N_11117,N_10239,N_10251);
or U11118 (N_11118,N_10468,N_10156);
xnor U11119 (N_11119,N_9787,N_10233);
or U11120 (N_11120,N_9981,N_9907);
or U11121 (N_11121,N_10340,N_10210);
nand U11122 (N_11122,N_10394,N_10073);
or U11123 (N_11123,N_10492,N_10212);
or U11124 (N_11124,N_10004,N_10403);
nor U11125 (N_11125,N_10178,N_9841);
and U11126 (N_11126,N_9924,N_10060);
or U11127 (N_11127,N_10050,N_9966);
nand U11128 (N_11128,N_9926,N_10175);
or U11129 (N_11129,N_10104,N_9799);
and U11130 (N_11130,N_10370,N_10321);
nand U11131 (N_11131,N_9872,N_9837);
or U11132 (N_11132,N_9932,N_10137);
nor U11133 (N_11133,N_10069,N_10147);
nand U11134 (N_11134,N_10041,N_10479);
nand U11135 (N_11135,N_10073,N_9925);
and U11136 (N_11136,N_10219,N_10049);
xor U11137 (N_11137,N_10487,N_10342);
nand U11138 (N_11138,N_9966,N_10308);
nand U11139 (N_11139,N_9765,N_10016);
xnor U11140 (N_11140,N_10296,N_9814);
or U11141 (N_11141,N_10475,N_9823);
xnor U11142 (N_11142,N_10052,N_9943);
or U11143 (N_11143,N_9851,N_10223);
nand U11144 (N_11144,N_10144,N_10338);
nor U11145 (N_11145,N_10015,N_9825);
nor U11146 (N_11146,N_10433,N_10076);
xnor U11147 (N_11147,N_10145,N_10211);
nor U11148 (N_11148,N_10028,N_10003);
nand U11149 (N_11149,N_10085,N_10443);
or U11150 (N_11150,N_10389,N_9837);
and U11151 (N_11151,N_9789,N_10112);
xnor U11152 (N_11152,N_9941,N_10353);
and U11153 (N_11153,N_10202,N_10069);
nor U11154 (N_11154,N_9771,N_10077);
nor U11155 (N_11155,N_10084,N_10106);
or U11156 (N_11156,N_9961,N_10419);
xor U11157 (N_11157,N_9877,N_9768);
nand U11158 (N_11158,N_9819,N_10229);
nand U11159 (N_11159,N_9969,N_10104);
and U11160 (N_11160,N_10277,N_10301);
or U11161 (N_11161,N_9863,N_10026);
xor U11162 (N_11162,N_10368,N_9752);
or U11163 (N_11163,N_10188,N_10355);
and U11164 (N_11164,N_10195,N_9779);
or U11165 (N_11165,N_10168,N_9906);
nor U11166 (N_11166,N_10187,N_10430);
nor U11167 (N_11167,N_10491,N_10314);
xor U11168 (N_11168,N_10075,N_9917);
nand U11169 (N_11169,N_9937,N_10024);
xor U11170 (N_11170,N_10373,N_10213);
xnor U11171 (N_11171,N_9999,N_10198);
nand U11172 (N_11172,N_10340,N_10370);
xnor U11173 (N_11173,N_10130,N_10277);
nand U11174 (N_11174,N_10380,N_9898);
and U11175 (N_11175,N_10104,N_10411);
or U11176 (N_11176,N_9921,N_9791);
xor U11177 (N_11177,N_10434,N_10242);
and U11178 (N_11178,N_10429,N_10174);
xor U11179 (N_11179,N_10484,N_10188);
nand U11180 (N_11180,N_10411,N_10395);
nor U11181 (N_11181,N_9899,N_10101);
xor U11182 (N_11182,N_9868,N_10101);
or U11183 (N_11183,N_10156,N_10267);
xor U11184 (N_11184,N_10125,N_10425);
nor U11185 (N_11185,N_10121,N_9786);
nor U11186 (N_11186,N_10064,N_9756);
and U11187 (N_11187,N_9954,N_10190);
nand U11188 (N_11188,N_10047,N_9791);
xor U11189 (N_11189,N_10484,N_10091);
or U11190 (N_11190,N_10452,N_10418);
nand U11191 (N_11191,N_9772,N_10448);
or U11192 (N_11192,N_10287,N_10487);
and U11193 (N_11193,N_10005,N_9806);
or U11194 (N_11194,N_10103,N_9852);
xnor U11195 (N_11195,N_10040,N_10346);
and U11196 (N_11196,N_10192,N_10021);
or U11197 (N_11197,N_10308,N_10492);
nor U11198 (N_11198,N_10070,N_10084);
xor U11199 (N_11199,N_9912,N_10002);
xor U11200 (N_11200,N_9843,N_10484);
nor U11201 (N_11201,N_10307,N_10450);
xor U11202 (N_11202,N_10281,N_10279);
nor U11203 (N_11203,N_9891,N_9927);
and U11204 (N_11204,N_9887,N_10433);
and U11205 (N_11205,N_10476,N_10254);
nor U11206 (N_11206,N_9902,N_10402);
nor U11207 (N_11207,N_9930,N_10120);
and U11208 (N_11208,N_10267,N_10460);
or U11209 (N_11209,N_10392,N_10369);
nand U11210 (N_11210,N_10203,N_10233);
nand U11211 (N_11211,N_10137,N_9815);
xor U11212 (N_11212,N_9910,N_10296);
or U11213 (N_11213,N_9766,N_9930);
nand U11214 (N_11214,N_10172,N_10398);
and U11215 (N_11215,N_9857,N_9803);
xnor U11216 (N_11216,N_10388,N_9821);
nor U11217 (N_11217,N_10169,N_9945);
nand U11218 (N_11218,N_9845,N_10132);
xor U11219 (N_11219,N_10221,N_10367);
xor U11220 (N_11220,N_10081,N_10307);
and U11221 (N_11221,N_10294,N_10050);
and U11222 (N_11222,N_10029,N_10230);
nor U11223 (N_11223,N_10024,N_10213);
xnor U11224 (N_11224,N_9966,N_9904);
and U11225 (N_11225,N_10175,N_10251);
or U11226 (N_11226,N_10001,N_9927);
xnor U11227 (N_11227,N_9820,N_9882);
nand U11228 (N_11228,N_9816,N_9765);
xor U11229 (N_11229,N_10198,N_9781);
and U11230 (N_11230,N_10150,N_10057);
nand U11231 (N_11231,N_9827,N_10367);
and U11232 (N_11232,N_9859,N_10397);
xnor U11233 (N_11233,N_10369,N_9968);
nor U11234 (N_11234,N_10056,N_9805);
nor U11235 (N_11235,N_10082,N_10323);
xnor U11236 (N_11236,N_10174,N_10453);
nand U11237 (N_11237,N_10060,N_9949);
and U11238 (N_11238,N_10336,N_10320);
nand U11239 (N_11239,N_9996,N_10441);
nand U11240 (N_11240,N_10488,N_10341);
nor U11241 (N_11241,N_10199,N_10437);
and U11242 (N_11242,N_10365,N_10382);
or U11243 (N_11243,N_10345,N_10174);
or U11244 (N_11244,N_9759,N_10118);
nor U11245 (N_11245,N_10336,N_10096);
or U11246 (N_11246,N_10478,N_9936);
xnor U11247 (N_11247,N_10192,N_10481);
and U11248 (N_11248,N_10072,N_9991);
xnor U11249 (N_11249,N_10269,N_9910);
or U11250 (N_11250,N_11126,N_10977);
nand U11251 (N_11251,N_11131,N_10540);
xor U11252 (N_11252,N_10834,N_11199);
and U11253 (N_11253,N_11197,N_10951);
xor U11254 (N_11254,N_11025,N_11009);
nand U11255 (N_11255,N_11233,N_10684);
xor U11256 (N_11256,N_10722,N_11024);
and U11257 (N_11257,N_10967,N_10703);
xnor U11258 (N_11258,N_10856,N_10654);
xnor U11259 (N_11259,N_10509,N_11015);
xor U11260 (N_11260,N_11163,N_10518);
xor U11261 (N_11261,N_10646,N_10618);
or U11262 (N_11262,N_11210,N_11115);
nor U11263 (N_11263,N_11236,N_11152);
nor U11264 (N_11264,N_10903,N_10702);
or U11265 (N_11265,N_11171,N_10554);
and U11266 (N_11266,N_10689,N_11208);
or U11267 (N_11267,N_10687,N_10704);
nor U11268 (N_11268,N_10695,N_11005);
nor U11269 (N_11269,N_10806,N_10674);
and U11270 (N_11270,N_10517,N_10634);
nand U11271 (N_11271,N_10681,N_10602);
or U11272 (N_11272,N_10905,N_10897);
and U11273 (N_11273,N_10894,N_10755);
and U11274 (N_11274,N_11003,N_10958);
nor U11275 (N_11275,N_10882,N_10635);
and U11276 (N_11276,N_10948,N_11107);
or U11277 (N_11277,N_10575,N_10579);
nor U11278 (N_11278,N_11013,N_10623);
nand U11279 (N_11279,N_11190,N_10985);
nand U11280 (N_11280,N_10560,N_10547);
and U11281 (N_11281,N_10576,N_10523);
nor U11282 (N_11282,N_10633,N_10734);
nand U11283 (N_11283,N_11212,N_10921);
nor U11284 (N_11284,N_10876,N_10629);
and U11285 (N_11285,N_11019,N_10924);
xor U11286 (N_11286,N_11148,N_10655);
or U11287 (N_11287,N_10609,N_11004);
and U11288 (N_11288,N_11010,N_10658);
and U11289 (N_11289,N_10715,N_10556);
and U11290 (N_11290,N_11124,N_11158);
or U11291 (N_11291,N_10881,N_10991);
and U11292 (N_11292,N_10778,N_10521);
xor U11293 (N_11293,N_11247,N_10793);
and U11294 (N_11294,N_10960,N_10711);
nor U11295 (N_11295,N_11032,N_11156);
xnor U11296 (N_11296,N_10608,N_11240);
nor U11297 (N_11297,N_10616,N_10824);
xnor U11298 (N_11298,N_10796,N_11187);
or U11299 (N_11299,N_10961,N_11119);
xnor U11300 (N_11300,N_10808,N_10941);
xor U11301 (N_11301,N_10573,N_11087);
xor U11302 (N_11302,N_10879,N_10913);
nor U11303 (N_11303,N_10744,N_10762);
nor U11304 (N_11304,N_10822,N_10999);
nor U11305 (N_11305,N_11064,N_10752);
or U11306 (N_11306,N_10983,N_10639);
nor U11307 (N_11307,N_11023,N_10594);
nand U11308 (N_11308,N_11037,N_10982);
and U11309 (N_11309,N_10838,N_10846);
nor U11310 (N_11310,N_11214,N_10984);
or U11311 (N_11311,N_10500,N_11026);
nand U11312 (N_11312,N_11176,N_11061);
xnor U11313 (N_11313,N_10688,N_11222);
or U11314 (N_11314,N_10745,N_11196);
nand U11315 (N_11315,N_11194,N_11175);
xor U11316 (N_11316,N_10536,N_10835);
xnor U11317 (N_11317,N_10840,N_10945);
and U11318 (N_11318,N_10736,N_10511);
nor U11319 (N_11319,N_11067,N_10849);
xor U11320 (N_11320,N_10550,N_10767);
xor U11321 (N_11321,N_10875,N_10940);
or U11322 (N_11322,N_11213,N_11167);
nand U11323 (N_11323,N_11170,N_10901);
xor U11324 (N_11324,N_11077,N_10908);
xnor U11325 (N_11325,N_10836,N_10637);
nor U11326 (N_11326,N_10601,N_10993);
nand U11327 (N_11327,N_10775,N_11218);
nor U11328 (N_11328,N_11056,N_11044);
and U11329 (N_11329,N_10773,N_11092);
or U11330 (N_11330,N_10502,N_10530);
nand U11331 (N_11331,N_10677,N_10997);
and U11332 (N_11332,N_10870,N_10668);
and U11333 (N_11333,N_11122,N_10611);
and U11334 (N_11334,N_11052,N_10583);
xnor U11335 (N_11335,N_10662,N_10898);
and U11336 (N_11336,N_10992,N_11104);
nand U11337 (N_11337,N_11177,N_10785);
and U11338 (N_11338,N_11203,N_10770);
and U11339 (N_11339,N_11165,N_11215);
and U11340 (N_11340,N_11047,N_11138);
and U11341 (N_11341,N_10526,N_10569);
and U11342 (N_11342,N_11112,N_10878);
nor U11343 (N_11343,N_11111,N_11198);
or U11344 (N_11344,N_10725,N_10694);
xnor U11345 (N_11345,N_10619,N_10606);
nor U11346 (N_11346,N_10636,N_10890);
xor U11347 (N_11347,N_10656,N_10917);
nand U11348 (N_11348,N_10801,N_10508);
or U11349 (N_11349,N_10872,N_11065);
or U11350 (N_11350,N_11086,N_11183);
nand U11351 (N_11351,N_10645,N_10580);
xor U11352 (N_11352,N_10911,N_10716);
or U11353 (N_11353,N_10590,N_10818);
xnor U11354 (N_11354,N_10717,N_10631);
nand U11355 (N_11355,N_11185,N_10612);
nand U11356 (N_11356,N_11182,N_11181);
nand U11357 (N_11357,N_10915,N_10868);
nor U11358 (N_11358,N_11226,N_11029);
nand U11359 (N_11359,N_10589,N_10784);
nand U11360 (N_11360,N_10650,N_10730);
or U11361 (N_11361,N_10820,N_11098);
nor U11362 (N_11362,N_10975,N_11120);
or U11363 (N_11363,N_10859,N_10741);
nor U11364 (N_11364,N_10599,N_11193);
xor U11365 (N_11365,N_10931,N_10615);
xnor U11366 (N_11366,N_11143,N_11018);
xnor U11367 (N_11367,N_11231,N_10660);
nand U11368 (N_11368,N_10855,N_11160);
or U11369 (N_11369,N_10987,N_10877);
nand U11370 (N_11370,N_11083,N_10708);
and U11371 (N_11371,N_10976,N_10790);
and U11372 (N_11372,N_10647,N_10548);
nor U11373 (N_11373,N_11205,N_10735);
or U11374 (N_11374,N_11066,N_11162);
xor U11375 (N_11375,N_10544,N_11063);
nand U11376 (N_11376,N_10607,N_10821);
or U11377 (N_11377,N_10614,N_11166);
nand U11378 (N_11378,N_10567,N_10803);
nand U11379 (N_11379,N_10747,N_10728);
nor U11380 (N_11380,N_11238,N_10990);
nand U11381 (N_11381,N_11040,N_10974);
or U11382 (N_11382,N_10667,N_11225);
nand U11383 (N_11383,N_10831,N_11057);
nand U11384 (N_11384,N_11031,N_10817);
nor U11385 (N_11385,N_10857,N_10723);
or U11386 (N_11386,N_10542,N_10910);
xor U11387 (N_11387,N_11059,N_11128);
and U11388 (N_11388,N_11058,N_10553);
and U11389 (N_11389,N_11249,N_10693);
and U11390 (N_11390,N_10998,N_11036);
nor U11391 (N_11391,N_11189,N_10559);
and U11392 (N_11392,N_10659,N_10621);
nor U11393 (N_11393,N_10844,N_10680);
and U11394 (N_11394,N_10845,N_10597);
nor U11395 (N_11395,N_11123,N_10942);
xor U11396 (N_11396,N_10685,N_10783);
xor U11397 (N_11397,N_10833,N_11142);
or U11398 (N_11398,N_11050,N_11093);
nand U11399 (N_11399,N_11051,N_10832);
or U11400 (N_11400,N_11094,N_11114);
nand U11401 (N_11401,N_10925,N_11146);
xnor U11402 (N_11402,N_10740,N_10811);
xor U11403 (N_11403,N_11217,N_10828);
or U11404 (N_11404,N_10825,N_10651);
or U11405 (N_11405,N_11145,N_10810);
xnor U11406 (N_11406,N_11161,N_11125);
or U11407 (N_11407,N_10989,N_10871);
or U11408 (N_11408,N_10853,N_10779);
nand U11409 (N_11409,N_10952,N_11244);
or U11410 (N_11410,N_10527,N_10585);
nand U11411 (N_11411,N_11060,N_11076);
xor U11412 (N_11412,N_10776,N_10979);
nand U11413 (N_11413,N_10738,N_10813);
nor U11414 (N_11414,N_10698,N_10807);
nor U11415 (N_11415,N_11164,N_10938);
nand U11416 (N_11416,N_10692,N_11014);
xor U11417 (N_11417,N_10839,N_10522);
or U11418 (N_11418,N_11002,N_10787);
or U11419 (N_11419,N_11221,N_11246);
nor U11420 (N_11420,N_11000,N_10624);
and U11421 (N_11421,N_10653,N_10964);
nand U11422 (N_11422,N_11054,N_11006);
xnor U11423 (N_11423,N_10610,N_11016);
xnor U11424 (N_11424,N_11192,N_10678);
or U11425 (N_11425,N_11133,N_10541);
nand U11426 (N_11426,N_11089,N_10699);
or U11427 (N_11427,N_10705,N_10842);
nand U11428 (N_11428,N_10900,N_10549);
or U11429 (N_11429,N_10627,N_11074);
or U11430 (N_11430,N_11155,N_10710);
xor U11431 (N_11431,N_11021,N_11147);
and U11432 (N_11432,N_10850,N_11132);
and U11433 (N_11433,N_10848,N_11046);
or U11434 (N_11434,N_10919,N_11096);
nand U11435 (N_11435,N_10895,N_11140);
and U11436 (N_11436,N_10551,N_11038);
nor U11437 (N_11437,N_10843,N_10503);
nor U11438 (N_11438,N_10632,N_10706);
or U11439 (N_11439,N_11069,N_10869);
nor U11440 (N_11440,N_11184,N_11206);
or U11441 (N_11441,N_10930,N_10737);
xor U11442 (N_11442,N_10519,N_11118);
or U11443 (N_11443,N_10501,N_10746);
and U11444 (N_11444,N_10718,N_10622);
nand U11445 (N_11445,N_10804,N_10953);
and U11446 (N_11446,N_11109,N_10535);
nor U11447 (N_11447,N_10764,N_10972);
xor U11448 (N_11448,N_10934,N_10988);
nor U11449 (N_11449,N_10670,N_10754);
and U11450 (N_11450,N_10691,N_10543);
xnor U11451 (N_11451,N_11041,N_10928);
nor U11452 (N_11452,N_10907,N_10889);
or U11453 (N_11453,N_10739,N_10727);
nor U11454 (N_11454,N_10666,N_11039);
and U11455 (N_11455,N_10640,N_10920);
or U11456 (N_11456,N_11220,N_11135);
nand U11457 (N_11457,N_11027,N_10676);
or U11458 (N_11458,N_10969,N_10751);
xor U11459 (N_11459,N_10841,N_10593);
nand U11460 (N_11460,N_11117,N_10829);
or U11461 (N_11461,N_10625,N_10800);
xnor U11462 (N_11462,N_10719,N_11110);
and U11463 (N_11463,N_10798,N_10899);
and U11464 (N_11464,N_10863,N_10648);
xor U11465 (N_11465,N_11195,N_11127);
nand U11466 (N_11466,N_11049,N_10854);
nor U11467 (N_11467,N_11062,N_11099);
and U11468 (N_11468,N_11072,N_11073);
and U11469 (N_11469,N_11100,N_10709);
or U11470 (N_11470,N_11202,N_10732);
and U11471 (N_11471,N_10797,N_10902);
and U11472 (N_11472,N_10880,N_10552);
or U11473 (N_11473,N_10795,N_10534);
or U11474 (N_11474,N_10814,N_10760);
nand U11475 (N_11475,N_10944,N_10750);
xnor U11476 (N_11476,N_10954,N_11042);
or U11477 (N_11477,N_10891,N_10805);
or U11478 (N_11478,N_10690,N_10562);
xnor U11479 (N_11479,N_11200,N_10837);
or U11480 (N_11480,N_10520,N_11022);
nand U11481 (N_11481,N_10504,N_11033);
nor U11482 (N_11482,N_10957,N_10592);
nor U11483 (N_11483,N_10996,N_10799);
xor U11484 (N_11484,N_10682,N_10759);
or U11485 (N_11485,N_10577,N_11174);
nor U11486 (N_11486,N_11186,N_10596);
or U11487 (N_11487,N_11153,N_10909);
nand U11488 (N_11488,N_10932,N_11030);
xor U11489 (N_11489,N_10986,N_10701);
or U11490 (N_11490,N_11085,N_11237);
nand U11491 (N_11491,N_10620,N_10512);
or U11492 (N_11492,N_11154,N_11035);
nor U11493 (N_11493,N_10939,N_10851);
nor U11494 (N_11494,N_10978,N_11078);
nand U11495 (N_11495,N_11048,N_10545);
nor U11496 (N_11496,N_11180,N_10866);
or U11497 (N_11497,N_10756,N_10777);
or U11498 (N_11498,N_11017,N_10568);
and U11499 (N_11499,N_11075,N_11116);
nor U11500 (N_11500,N_10761,N_10574);
nand U11501 (N_11501,N_11082,N_10947);
nor U11502 (N_11502,N_10812,N_10586);
and U11503 (N_11503,N_11227,N_11071);
nand U11504 (N_11504,N_10792,N_10887);
nand U11505 (N_11505,N_11144,N_11008);
or U11506 (N_11506,N_10981,N_11216);
nand U11507 (N_11507,N_10883,N_11129);
and U11508 (N_11508,N_11151,N_10683);
xor U11509 (N_11509,N_11229,N_10714);
and U11510 (N_11510,N_10516,N_10628);
or U11511 (N_11511,N_10679,N_10864);
nand U11512 (N_11512,N_10906,N_10914);
xnor U11513 (N_11513,N_10571,N_10904);
xor U11514 (N_11514,N_11055,N_10994);
xor U11515 (N_11515,N_10507,N_11223);
xnor U11516 (N_11516,N_10697,N_10663);
or U11517 (N_11517,N_10918,N_10713);
nor U11518 (N_11518,N_10563,N_10995);
nand U11519 (N_11519,N_11159,N_11234);
xnor U11520 (N_11520,N_10661,N_10537);
nand U11521 (N_11521,N_10950,N_11178);
or U11522 (N_11522,N_10566,N_11053);
nand U11523 (N_11523,N_10962,N_10720);
nor U11524 (N_11524,N_11079,N_10561);
nor U11525 (N_11525,N_10643,N_11219);
or U11526 (N_11526,N_10587,N_10539);
or U11527 (N_11527,N_11102,N_11242);
nor U11528 (N_11528,N_10923,N_10827);
xnor U11529 (N_11529,N_10862,N_10927);
xor U11530 (N_11530,N_10686,N_11108);
or U11531 (N_11531,N_10772,N_10603);
xnor U11532 (N_11532,N_10700,N_10748);
and U11533 (N_11533,N_10933,N_10514);
and U11534 (N_11534,N_11106,N_10641);
nor U11535 (N_11535,N_10613,N_10652);
nand U11536 (N_11536,N_10830,N_10604);
nor U11537 (N_11537,N_11136,N_10823);
nand U11538 (N_11538,N_11139,N_11179);
xnor U11539 (N_11539,N_10861,N_10926);
or U11540 (N_11540,N_10729,N_10885);
or U11541 (N_11541,N_11043,N_10794);
or U11542 (N_11542,N_10766,N_10538);
nor U11543 (N_11543,N_11113,N_11137);
nor U11544 (N_11544,N_10753,N_11173);
nand U11545 (N_11545,N_11028,N_10768);
or U11546 (N_11546,N_10533,N_11070);
xor U11547 (N_11547,N_11134,N_11121);
and U11548 (N_11548,N_10578,N_10819);
or U11549 (N_11549,N_11091,N_10531);
nor U11550 (N_11550,N_10673,N_11149);
nor U11551 (N_11551,N_10546,N_11103);
and U11552 (N_11552,N_11239,N_10886);
nand U11553 (N_11553,N_10980,N_11095);
xnor U11554 (N_11554,N_10955,N_10749);
or U11555 (N_11555,N_11191,N_10581);
xnor U11556 (N_11556,N_10644,N_10721);
and U11557 (N_11557,N_11020,N_10630);
nor U11558 (N_11558,N_10584,N_11034);
nand U11559 (N_11559,N_10588,N_11235);
nor U11560 (N_11560,N_10565,N_11248);
and U11561 (N_11561,N_10815,N_10598);
nand U11562 (N_11562,N_11012,N_10963);
xor U11563 (N_11563,N_11068,N_10570);
nor U11564 (N_11564,N_10788,N_10860);
or U11565 (N_11565,N_10912,N_10858);
and U11566 (N_11566,N_10582,N_10742);
and U11567 (N_11567,N_10937,N_11101);
nor U11568 (N_11568,N_11243,N_11011);
nor U11569 (N_11569,N_10642,N_10600);
and U11570 (N_11570,N_10791,N_10675);
nand U11571 (N_11571,N_10672,N_11097);
xor U11572 (N_11572,N_10946,N_10956);
nor U11573 (N_11573,N_10771,N_10712);
nand U11574 (N_11574,N_10731,N_11207);
nor U11575 (N_11575,N_10893,N_11105);
nand U11576 (N_11576,N_10510,N_11230);
xor U11577 (N_11577,N_11150,N_10943);
or U11578 (N_11578,N_10626,N_11209);
and U11579 (N_11579,N_10555,N_10557);
nor U11580 (N_11580,N_10515,N_11157);
or U11581 (N_11581,N_10949,N_11084);
xor U11582 (N_11582,N_11204,N_11172);
nor U11583 (N_11583,N_10758,N_10780);
and U11584 (N_11584,N_11228,N_10595);
nor U11585 (N_11585,N_10696,N_10572);
nand U11586 (N_11586,N_11245,N_11001);
xor U11587 (N_11587,N_11224,N_10726);
xor U11588 (N_11588,N_11090,N_10782);
nand U11589 (N_11589,N_10707,N_10733);
xnor U11590 (N_11590,N_10916,N_11168);
or U11591 (N_11591,N_10524,N_10896);
and U11592 (N_11592,N_10671,N_11141);
nor U11593 (N_11593,N_10724,N_10852);
nand U11594 (N_11594,N_10506,N_11130);
xnor U11595 (N_11595,N_10781,N_10789);
or U11596 (N_11596,N_10922,N_10763);
or U11597 (N_11597,N_11188,N_10591);
and U11598 (N_11598,N_11169,N_10528);
nor U11599 (N_11599,N_10617,N_11045);
xor U11600 (N_11600,N_10867,N_11007);
xor U11601 (N_11601,N_10649,N_11232);
xor U11602 (N_11602,N_10786,N_10809);
and U11603 (N_11603,N_11211,N_10935);
and U11604 (N_11604,N_10765,N_11080);
and U11605 (N_11605,N_10874,N_10657);
and U11606 (N_11606,N_10558,N_10757);
nand U11607 (N_11607,N_10865,N_10529);
and U11608 (N_11608,N_10664,N_11081);
nor U11609 (N_11609,N_10959,N_10743);
nand U11610 (N_11610,N_10873,N_10826);
xnor U11611 (N_11611,N_10769,N_10605);
nor U11612 (N_11612,N_10816,N_10847);
nor U11613 (N_11613,N_10513,N_10532);
or U11614 (N_11614,N_11201,N_10638);
and U11615 (N_11615,N_10665,N_10936);
xnor U11616 (N_11616,N_10970,N_10966);
and U11617 (N_11617,N_10929,N_10892);
nand U11618 (N_11618,N_10525,N_10669);
nand U11619 (N_11619,N_11088,N_11241);
and U11620 (N_11620,N_10774,N_10973);
nand U11621 (N_11621,N_10884,N_10968);
nand U11622 (N_11622,N_10802,N_10971);
nand U11623 (N_11623,N_10965,N_10888);
nor U11624 (N_11624,N_10505,N_10564);
and U11625 (N_11625,N_10920,N_11080);
and U11626 (N_11626,N_10717,N_11112);
nor U11627 (N_11627,N_10675,N_11150);
nand U11628 (N_11628,N_11020,N_10604);
or U11629 (N_11629,N_10670,N_10664);
nand U11630 (N_11630,N_10503,N_10957);
xnor U11631 (N_11631,N_10994,N_11052);
xnor U11632 (N_11632,N_10700,N_11214);
and U11633 (N_11633,N_10793,N_10974);
or U11634 (N_11634,N_11228,N_10522);
and U11635 (N_11635,N_11047,N_10595);
nor U11636 (N_11636,N_11116,N_10593);
and U11637 (N_11637,N_10537,N_10539);
nor U11638 (N_11638,N_10593,N_10564);
nand U11639 (N_11639,N_10747,N_10959);
xor U11640 (N_11640,N_11188,N_10842);
and U11641 (N_11641,N_10998,N_11019);
and U11642 (N_11642,N_10530,N_11204);
nand U11643 (N_11643,N_11152,N_10634);
or U11644 (N_11644,N_11165,N_10624);
nor U11645 (N_11645,N_10503,N_10831);
nor U11646 (N_11646,N_11067,N_10828);
nor U11647 (N_11647,N_10722,N_10913);
xor U11648 (N_11648,N_10977,N_11094);
nand U11649 (N_11649,N_11057,N_11213);
nand U11650 (N_11650,N_11054,N_11131);
xnor U11651 (N_11651,N_11009,N_11185);
and U11652 (N_11652,N_11011,N_10548);
nor U11653 (N_11653,N_11149,N_10753);
or U11654 (N_11654,N_10667,N_10503);
and U11655 (N_11655,N_10971,N_10826);
or U11656 (N_11656,N_10870,N_11188);
nand U11657 (N_11657,N_10744,N_10917);
nand U11658 (N_11658,N_11147,N_10594);
and U11659 (N_11659,N_11054,N_10695);
nor U11660 (N_11660,N_10874,N_11113);
xor U11661 (N_11661,N_10718,N_10786);
xnor U11662 (N_11662,N_10576,N_11086);
nand U11663 (N_11663,N_11249,N_10569);
nor U11664 (N_11664,N_11238,N_11023);
or U11665 (N_11665,N_10875,N_11218);
xnor U11666 (N_11666,N_10648,N_10957);
nand U11667 (N_11667,N_10938,N_11036);
and U11668 (N_11668,N_10893,N_10745);
or U11669 (N_11669,N_11177,N_10744);
xnor U11670 (N_11670,N_10767,N_10590);
and U11671 (N_11671,N_10964,N_10825);
nor U11672 (N_11672,N_10707,N_10808);
and U11673 (N_11673,N_10993,N_10710);
and U11674 (N_11674,N_10563,N_10593);
and U11675 (N_11675,N_10868,N_10983);
nor U11676 (N_11676,N_11040,N_11077);
nor U11677 (N_11677,N_10925,N_11236);
and U11678 (N_11678,N_11192,N_10694);
nand U11679 (N_11679,N_10671,N_11033);
nand U11680 (N_11680,N_10687,N_10875);
or U11681 (N_11681,N_11146,N_11012);
and U11682 (N_11682,N_10966,N_10756);
or U11683 (N_11683,N_10934,N_11138);
or U11684 (N_11684,N_10919,N_11043);
or U11685 (N_11685,N_11121,N_11071);
nor U11686 (N_11686,N_10626,N_10866);
and U11687 (N_11687,N_11005,N_11176);
nor U11688 (N_11688,N_11040,N_11166);
nand U11689 (N_11689,N_10883,N_10956);
or U11690 (N_11690,N_11146,N_11200);
nand U11691 (N_11691,N_10637,N_11178);
nor U11692 (N_11692,N_10765,N_10769);
and U11693 (N_11693,N_10703,N_11089);
xor U11694 (N_11694,N_10549,N_10965);
and U11695 (N_11695,N_10623,N_11172);
nor U11696 (N_11696,N_10808,N_11022);
and U11697 (N_11697,N_10902,N_10653);
nor U11698 (N_11698,N_11240,N_10965);
nor U11699 (N_11699,N_11023,N_10579);
or U11700 (N_11700,N_10961,N_11248);
or U11701 (N_11701,N_10967,N_11231);
or U11702 (N_11702,N_11180,N_10729);
and U11703 (N_11703,N_11202,N_10599);
and U11704 (N_11704,N_11046,N_10951);
and U11705 (N_11705,N_10705,N_10693);
xor U11706 (N_11706,N_10887,N_11192);
and U11707 (N_11707,N_10744,N_10815);
or U11708 (N_11708,N_10900,N_10907);
xnor U11709 (N_11709,N_11225,N_11116);
nor U11710 (N_11710,N_10932,N_11080);
and U11711 (N_11711,N_11089,N_11192);
xnor U11712 (N_11712,N_11033,N_10580);
nor U11713 (N_11713,N_10675,N_10989);
nand U11714 (N_11714,N_10574,N_11015);
nand U11715 (N_11715,N_10915,N_10518);
nor U11716 (N_11716,N_10858,N_11220);
xnor U11717 (N_11717,N_10523,N_11165);
or U11718 (N_11718,N_10792,N_10946);
xor U11719 (N_11719,N_10980,N_10696);
or U11720 (N_11720,N_10687,N_10923);
nand U11721 (N_11721,N_10762,N_11035);
nand U11722 (N_11722,N_11157,N_10763);
nand U11723 (N_11723,N_10856,N_11191);
or U11724 (N_11724,N_11004,N_10935);
or U11725 (N_11725,N_11132,N_10693);
and U11726 (N_11726,N_10668,N_11098);
nor U11727 (N_11727,N_11042,N_11107);
xor U11728 (N_11728,N_10862,N_10565);
xor U11729 (N_11729,N_10828,N_11084);
nand U11730 (N_11730,N_10929,N_10796);
xnor U11731 (N_11731,N_10993,N_10981);
and U11732 (N_11732,N_11063,N_10509);
or U11733 (N_11733,N_10817,N_10629);
xor U11734 (N_11734,N_10651,N_10978);
xor U11735 (N_11735,N_11008,N_10814);
and U11736 (N_11736,N_11087,N_10577);
or U11737 (N_11737,N_11158,N_10652);
xnor U11738 (N_11738,N_11212,N_10685);
nor U11739 (N_11739,N_11200,N_10511);
nor U11740 (N_11740,N_10591,N_11039);
or U11741 (N_11741,N_10805,N_10788);
or U11742 (N_11742,N_10639,N_10535);
nand U11743 (N_11743,N_10872,N_10845);
nand U11744 (N_11744,N_10973,N_10628);
nand U11745 (N_11745,N_10676,N_11073);
nand U11746 (N_11746,N_10587,N_11189);
xnor U11747 (N_11747,N_10808,N_10533);
xor U11748 (N_11748,N_10748,N_10971);
nand U11749 (N_11749,N_10525,N_11168);
or U11750 (N_11750,N_10870,N_10636);
nor U11751 (N_11751,N_11038,N_10777);
and U11752 (N_11752,N_11200,N_10566);
and U11753 (N_11753,N_10877,N_10546);
nor U11754 (N_11754,N_10539,N_11043);
nand U11755 (N_11755,N_10701,N_10621);
or U11756 (N_11756,N_11008,N_10631);
nand U11757 (N_11757,N_10772,N_11003);
and U11758 (N_11758,N_10562,N_10555);
and U11759 (N_11759,N_11097,N_10703);
nor U11760 (N_11760,N_11143,N_10838);
or U11761 (N_11761,N_10665,N_10676);
nor U11762 (N_11762,N_11107,N_10905);
or U11763 (N_11763,N_10929,N_11094);
nand U11764 (N_11764,N_11119,N_10937);
and U11765 (N_11765,N_11154,N_11114);
or U11766 (N_11766,N_11002,N_10880);
and U11767 (N_11767,N_10919,N_10649);
nor U11768 (N_11768,N_11056,N_10576);
or U11769 (N_11769,N_10901,N_10740);
nand U11770 (N_11770,N_10714,N_11043);
and U11771 (N_11771,N_11219,N_10720);
or U11772 (N_11772,N_10957,N_11013);
or U11773 (N_11773,N_10587,N_10825);
and U11774 (N_11774,N_10523,N_10780);
xor U11775 (N_11775,N_10992,N_11123);
nand U11776 (N_11776,N_11126,N_11088);
and U11777 (N_11777,N_11244,N_10541);
and U11778 (N_11778,N_10903,N_10807);
xnor U11779 (N_11779,N_10596,N_10595);
or U11780 (N_11780,N_10726,N_10855);
and U11781 (N_11781,N_10589,N_10936);
and U11782 (N_11782,N_11034,N_10521);
and U11783 (N_11783,N_11152,N_10525);
and U11784 (N_11784,N_11001,N_10685);
nor U11785 (N_11785,N_10849,N_11058);
nand U11786 (N_11786,N_10869,N_10680);
nand U11787 (N_11787,N_11017,N_10777);
nor U11788 (N_11788,N_10941,N_10949);
or U11789 (N_11789,N_11105,N_10925);
nand U11790 (N_11790,N_10521,N_10937);
nor U11791 (N_11791,N_11041,N_10612);
and U11792 (N_11792,N_10965,N_10749);
nor U11793 (N_11793,N_10794,N_10646);
xnor U11794 (N_11794,N_11064,N_10677);
and U11795 (N_11795,N_10604,N_11144);
nor U11796 (N_11796,N_11009,N_10731);
nor U11797 (N_11797,N_10898,N_10782);
and U11798 (N_11798,N_11024,N_11147);
and U11799 (N_11799,N_10649,N_10627);
or U11800 (N_11800,N_11205,N_10951);
nand U11801 (N_11801,N_10600,N_11133);
nor U11802 (N_11802,N_10541,N_10826);
xor U11803 (N_11803,N_11132,N_11037);
xnor U11804 (N_11804,N_10683,N_10771);
xor U11805 (N_11805,N_11236,N_11108);
nand U11806 (N_11806,N_11163,N_10867);
or U11807 (N_11807,N_11248,N_10531);
or U11808 (N_11808,N_10900,N_10521);
nor U11809 (N_11809,N_11142,N_11244);
xor U11810 (N_11810,N_10549,N_10522);
xor U11811 (N_11811,N_10523,N_10996);
nand U11812 (N_11812,N_11195,N_10741);
nor U11813 (N_11813,N_10796,N_10558);
or U11814 (N_11814,N_10862,N_11155);
nand U11815 (N_11815,N_11130,N_10642);
and U11816 (N_11816,N_10857,N_10896);
or U11817 (N_11817,N_10698,N_10869);
nor U11818 (N_11818,N_10502,N_10536);
and U11819 (N_11819,N_10659,N_10845);
and U11820 (N_11820,N_10856,N_10833);
nand U11821 (N_11821,N_10748,N_10529);
and U11822 (N_11822,N_10515,N_11060);
or U11823 (N_11823,N_10558,N_11103);
xnor U11824 (N_11824,N_10933,N_11193);
or U11825 (N_11825,N_10881,N_10951);
nor U11826 (N_11826,N_11190,N_10824);
xor U11827 (N_11827,N_10831,N_10848);
nand U11828 (N_11828,N_10639,N_10604);
xnor U11829 (N_11829,N_11197,N_11135);
xor U11830 (N_11830,N_10527,N_11097);
and U11831 (N_11831,N_11003,N_10732);
or U11832 (N_11832,N_10887,N_11098);
xnor U11833 (N_11833,N_10526,N_10870);
or U11834 (N_11834,N_11119,N_11214);
xor U11835 (N_11835,N_10501,N_10824);
or U11836 (N_11836,N_10585,N_11129);
and U11837 (N_11837,N_10913,N_10554);
nand U11838 (N_11838,N_10720,N_11131);
or U11839 (N_11839,N_10781,N_10763);
xnor U11840 (N_11840,N_10568,N_10973);
nand U11841 (N_11841,N_10959,N_10775);
nor U11842 (N_11842,N_11196,N_11093);
nand U11843 (N_11843,N_10696,N_10567);
xor U11844 (N_11844,N_11059,N_10951);
nor U11845 (N_11845,N_10693,N_10856);
nor U11846 (N_11846,N_10591,N_10726);
or U11847 (N_11847,N_11150,N_10861);
nor U11848 (N_11848,N_11173,N_10810);
nor U11849 (N_11849,N_11042,N_10948);
xor U11850 (N_11850,N_11090,N_11239);
and U11851 (N_11851,N_11074,N_11106);
nor U11852 (N_11852,N_10709,N_10804);
xnor U11853 (N_11853,N_11054,N_11146);
and U11854 (N_11854,N_10948,N_11119);
nor U11855 (N_11855,N_10963,N_10520);
nand U11856 (N_11856,N_10613,N_10513);
or U11857 (N_11857,N_11232,N_10574);
and U11858 (N_11858,N_10597,N_10778);
and U11859 (N_11859,N_10618,N_10975);
xnor U11860 (N_11860,N_10670,N_10590);
nor U11861 (N_11861,N_11149,N_10734);
nor U11862 (N_11862,N_11118,N_10753);
nand U11863 (N_11863,N_11234,N_11209);
or U11864 (N_11864,N_10944,N_10694);
nor U11865 (N_11865,N_10701,N_10767);
xor U11866 (N_11866,N_11235,N_10672);
and U11867 (N_11867,N_10560,N_10908);
and U11868 (N_11868,N_10603,N_10675);
and U11869 (N_11869,N_11025,N_10599);
or U11870 (N_11870,N_10688,N_10508);
nor U11871 (N_11871,N_10581,N_11114);
or U11872 (N_11872,N_10682,N_10782);
xor U11873 (N_11873,N_10767,N_10633);
xor U11874 (N_11874,N_10541,N_10998);
xor U11875 (N_11875,N_11161,N_10892);
xor U11876 (N_11876,N_10656,N_10858);
or U11877 (N_11877,N_10727,N_10588);
and U11878 (N_11878,N_10605,N_11114);
xor U11879 (N_11879,N_11094,N_11245);
nand U11880 (N_11880,N_11094,N_11185);
nor U11881 (N_11881,N_10806,N_10691);
and U11882 (N_11882,N_11135,N_10896);
or U11883 (N_11883,N_11209,N_11222);
xor U11884 (N_11884,N_10572,N_10678);
nor U11885 (N_11885,N_10525,N_11119);
nand U11886 (N_11886,N_10875,N_11026);
nor U11887 (N_11887,N_11237,N_10890);
nand U11888 (N_11888,N_10526,N_10693);
nor U11889 (N_11889,N_10839,N_10586);
and U11890 (N_11890,N_11197,N_10743);
and U11891 (N_11891,N_10704,N_11084);
or U11892 (N_11892,N_10771,N_10538);
and U11893 (N_11893,N_11227,N_10895);
nor U11894 (N_11894,N_10742,N_10739);
or U11895 (N_11895,N_11056,N_10899);
and U11896 (N_11896,N_10610,N_10805);
or U11897 (N_11897,N_11046,N_10828);
nand U11898 (N_11898,N_11219,N_10880);
nand U11899 (N_11899,N_10887,N_11119);
and U11900 (N_11900,N_10599,N_10736);
xnor U11901 (N_11901,N_11190,N_10889);
nor U11902 (N_11902,N_11052,N_10623);
nand U11903 (N_11903,N_11015,N_11108);
nor U11904 (N_11904,N_10738,N_10526);
xnor U11905 (N_11905,N_10839,N_11201);
and U11906 (N_11906,N_10519,N_11179);
or U11907 (N_11907,N_10884,N_10835);
nand U11908 (N_11908,N_10744,N_10670);
xnor U11909 (N_11909,N_10853,N_10599);
nor U11910 (N_11910,N_11199,N_10853);
nand U11911 (N_11911,N_10777,N_10982);
nand U11912 (N_11912,N_10584,N_11014);
nor U11913 (N_11913,N_10755,N_11138);
nand U11914 (N_11914,N_10831,N_11005);
xnor U11915 (N_11915,N_10626,N_10759);
nand U11916 (N_11916,N_11069,N_11233);
nand U11917 (N_11917,N_10877,N_10798);
and U11918 (N_11918,N_10741,N_11050);
nor U11919 (N_11919,N_11215,N_10899);
xnor U11920 (N_11920,N_11243,N_10603);
xor U11921 (N_11921,N_11081,N_10754);
and U11922 (N_11922,N_11119,N_11184);
nand U11923 (N_11923,N_11065,N_10921);
xnor U11924 (N_11924,N_10956,N_11239);
nand U11925 (N_11925,N_11115,N_10588);
and U11926 (N_11926,N_11068,N_10908);
or U11927 (N_11927,N_10833,N_10823);
xor U11928 (N_11928,N_11120,N_10757);
xnor U11929 (N_11929,N_10957,N_10891);
xor U11930 (N_11930,N_11076,N_10804);
xnor U11931 (N_11931,N_11102,N_11002);
and U11932 (N_11932,N_10791,N_10606);
xor U11933 (N_11933,N_10889,N_10738);
nor U11934 (N_11934,N_11106,N_11199);
nand U11935 (N_11935,N_10800,N_11048);
xnor U11936 (N_11936,N_10899,N_11079);
or U11937 (N_11937,N_11121,N_11083);
xor U11938 (N_11938,N_11148,N_10810);
nor U11939 (N_11939,N_11010,N_11142);
nor U11940 (N_11940,N_10840,N_10508);
and U11941 (N_11941,N_10520,N_10756);
and U11942 (N_11942,N_10978,N_11015);
or U11943 (N_11943,N_10936,N_10840);
and U11944 (N_11944,N_11087,N_11216);
xor U11945 (N_11945,N_10892,N_10717);
nor U11946 (N_11946,N_10923,N_10882);
or U11947 (N_11947,N_10851,N_11118);
nand U11948 (N_11948,N_11206,N_10907);
xnor U11949 (N_11949,N_11114,N_11017);
xor U11950 (N_11950,N_10527,N_10919);
nor U11951 (N_11951,N_10721,N_10957);
and U11952 (N_11952,N_10678,N_11036);
and U11953 (N_11953,N_10924,N_11186);
and U11954 (N_11954,N_10797,N_10832);
or U11955 (N_11955,N_11197,N_10853);
and U11956 (N_11956,N_10556,N_10977);
xor U11957 (N_11957,N_11073,N_10594);
nand U11958 (N_11958,N_10901,N_10806);
and U11959 (N_11959,N_10802,N_10685);
xnor U11960 (N_11960,N_10890,N_11157);
xnor U11961 (N_11961,N_10689,N_10823);
xnor U11962 (N_11962,N_11113,N_10794);
and U11963 (N_11963,N_10654,N_10540);
and U11964 (N_11964,N_11076,N_10833);
xnor U11965 (N_11965,N_11034,N_10699);
xnor U11966 (N_11966,N_11162,N_10666);
xor U11967 (N_11967,N_10735,N_11175);
or U11968 (N_11968,N_10688,N_10875);
nor U11969 (N_11969,N_10966,N_10805);
xnor U11970 (N_11970,N_10604,N_10511);
or U11971 (N_11971,N_11077,N_10821);
or U11972 (N_11972,N_10609,N_10525);
nand U11973 (N_11973,N_10671,N_11107);
or U11974 (N_11974,N_10755,N_11175);
or U11975 (N_11975,N_11003,N_10525);
xnor U11976 (N_11976,N_10524,N_10621);
and U11977 (N_11977,N_10680,N_10820);
xnor U11978 (N_11978,N_10664,N_11039);
xnor U11979 (N_11979,N_11171,N_10536);
nand U11980 (N_11980,N_11180,N_10661);
and U11981 (N_11981,N_11106,N_10836);
nand U11982 (N_11982,N_10988,N_11240);
nand U11983 (N_11983,N_10520,N_10504);
and U11984 (N_11984,N_10598,N_10908);
xor U11985 (N_11985,N_11010,N_10597);
nor U11986 (N_11986,N_10931,N_10700);
nor U11987 (N_11987,N_11015,N_10723);
and U11988 (N_11988,N_10558,N_10691);
nand U11989 (N_11989,N_10648,N_10643);
nand U11990 (N_11990,N_10674,N_10562);
or U11991 (N_11991,N_10580,N_11045);
nor U11992 (N_11992,N_11019,N_10835);
nand U11993 (N_11993,N_10637,N_10855);
nand U11994 (N_11994,N_11051,N_10530);
and U11995 (N_11995,N_10915,N_11117);
and U11996 (N_11996,N_10817,N_10684);
and U11997 (N_11997,N_10505,N_10815);
xor U11998 (N_11998,N_10508,N_10912);
xnor U11999 (N_11999,N_11212,N_10870);
and U12000 (N_12000,N_11714,N_11991);
xor U12001 (N_12001,N_11726,N_11706);
xnor U12002 (N_12002,N_11792,N_11830);
or U12003 (N_12003,N_11552,N_11260);
xnor U12004 (N_12004,N_11691,N_11875);
xor U12005 (N_12005,N_11310,N_11938);
and U12006 (N_12006,N_11580,N_11890);
xor U12007 (N_12007,N_11320,N_11809);
xnor U12008 (N_12008,N_11453,N_11837);
or U12009 (N_12009,N_11971,N_11587);
nand U12010 (N_12010,N_11978,N_11669);
or U12011 (N_12011,N_11567,N_11914);
xnor U12012 (N_12012,N_11636,N_11266);
nor U12013 (N_12013,N_11823,N_11542);
xor U12014 (N_12014,N_11509,N_11425);
xnor U12015 (N_12015,N_11404,N_11607);
xnor U12016 (N_12016,N_11783,N_11822);
nor U12017 (N_12017,N_11810,N_11719);
and U12018 (N_12018,N_11947,N_11395);
or U12019 (N_12019,N_11759,N_11447);
or U12020 (N_12020,N_11250,N_11796);
nand U12021 (N_12021,N_11676,N_11570);
or U12022 (N_12022,N_11328,N_11268);
nand U12023 (N_12023,N_11274,N_11535);
nand U12024 (N_12024,N_11949,N_11973);
or U12025 (N_12025,N_11325,N_11708);
xnor U12026 (N_12026,N_11741,N_11705);
nor U12027 (N_12027,N_11743,N_11667);
nand U12028 (N_12028,N_11322,N_11637);
nor U12029 (N_12029,N_11370,N_11657);
and U12030 (N_12030,N_11256,N_11711);
xor U12031 (N_12031,N_11625,N_11794);
and U12032 (N_12032,N_11273,N_11656);
xor U12033 (N_12033,N_11617,N_11801);
nor U12034 (N_12034,N_11870,N_11622);
or U12035 (N_12035,N_11311,N_11684);
nand U12036 (N_12036,N_11892,N_11472);
nor U12037 (N_12037,N_11631,N_11730);
and U12038 (N_12038,N_11868,N_11886);
nor U12039 (N_12039,N_11693,N_11300);
xnor U12040 (N_12040,N_11884,N_11482);
nand U12041 (N_12041,N_11672,N_11775);
xnor U12042 (N_12042,N_11692,N_11508);
nand U12043 (N_12043,N_11519,N_11613);
and U12044 (N_12044,N_11731,N_11859);
and U12045 (N_12045,N_11873,N_11774);
xor U12046 (N_12046,N_11394,N_11764);
nor U12047 (N_12047,N_11770,N_11324);
nand U12048 (N_12048,N_11765,N_11299);
and U12049 (N_12049,N_11416,N_11514);
xor U12050 (N_12050,N_11757,N_11791);
nor U12051 (N_12051,N_11471,N_11318);
nor U12052 (N_12052,N_11339,N_11557);
nor U12053 (N_12053,N_11492,N_11965);
xnor U12054 (N_12054,N_11593,N_11660);
and U12055 (N_12055,N_11555,N_11422);
nor U12056 (N_12056,N_11553,N_11960);
nand U12057 (N_12057,N_11291,N_11819);
nor U12058 (N_12058,N_11288,N_11984);
nand U12059 (N_12059,N_11917,N_11866);
xnor U12060 (N_12060,N_11712,N_11369);
or U12061 (N_12061,N_11588,N_11350);
or U12062 (N_12062,N_11645,N_11487);
and U12063 (N_12063,N_11462,N_11372);
nor U12064 (N_12064,N_11280,N_11415);
and U12065 (N_12065,N_11477,N_11689);
nand U12066 (N_12066,N_11966,N_11451);
nor U12067 (N_12067,N_11643,N_11710);
nor U12068 (N_12068,N_11264,N_11448);
xnor U12069 (N_12069,N_11261,N_11897);
and U12070 (N_12070,N_11611,N_11827);
or U12071 (N_12071,N_11488,N_11305);
nor U12072 (N_12072,N_11768,N_11915);
and U12073 (N_12073,N_11423,N_11355);
xnor U12074 (N_12074,N_11387,N_11352);
nand U12075 (N_12075,N_11616,N_11308);
nor U12076 (N_12076,N_11847,N_11627);
and U12077 (N_12077,N_11539,N_11861);
xor U12078 (N_12078,N_11685,N_11327);
nor U12079 (N_12079,N_11826,N_11814);
xor U12080 (N_12080,N_11351,N_11494);
xnor U12081 (N_12081,N_11844,N_11358);
or U12082 (N_12082,N_11748,N_11278);
and U12083 (N_12083,N_11906,N_11835);
xor U12084 (N_12084,N_11834,N_11994);
xnor U12085 (N_12085,N_11377,N_11614);
nand U12086 (N_12086,N_11968,N_11756);
or U12087 (N_12087,N_11480,N_11362);
nor U12088 (N_12088,N_11463,N_11779);
and U12089 (N_12089,N_11259,N_11338);
nor U12090 (N_12090,N_11746,N_11346);
nand U12091 (N_12091,N_11615,N_11516);
xor U12092 (N_12092,N_11646,N_11301);
xor U12093 (N_12093,N_11518,N_11772);
nand U12094 (N_12094,N_11502,N_11406);
and U12095 (N_12095,N_11262,N_11703);
nor U12096 (N_12096,N_11862,N_11655);
and U12097 (N_12097,N_11523,N_11939);
nor U12098 (N_12098,N_11849,N_11610);
xor U12099 (N_12099,N_11590,N_11695);
xnor U12100 (N_12100,N_11344,N_11976);
or U12101 (N_12101,N_11806,N_11524);
xor U12102 (N_12102,N_11818,N_11589);
xor U12103 (N_12103,N_11688,N_11521);
nor U12104 (N_12104,N_11674,N_11990);
and U12105 (N_12105,N_11433,N_11332);
and U12106 (N_12106,N_11931,N_11825);
xnor U12107 (N_12107,N_11739,N_11538);
nor U12108 (N_12108,N_11568,N_11527);
nand U12109 (N_12109,N_11908,N_11981);
and U12110 (N_12110,N_11715,N_11493);
nand U12111 (N_12111,N_11501,N_11277);
nand U12112 (N_12112,N_11983,N_11969);
xor U12113 (N_12113,N_11479,N_11964);
and U12114 (N_12114,N_11998,N_11860);
nor U12115 (N_12115,N_11761,N_11558);
nor U12116 (N_12116,N_11373,N_11885);
nor U12117 (N_12117,N_11534,N_11331);
or U12118 (N_12118,N_11444,N_11769);
xor U12119 (N_12119,N_11388,N_11909);
xnor U12120 (N_12120,N_11435,N_11948);
xnor U12121 (N_12121,N_11854,N_11722);
and U12122 (N_12122,N_11773,N_11661);
or U12123 (N_12123,N_11564,N_11478);
xor U12124 (N_12124,N_11790,N_11785);
nand U12125 (N_12125,N_11620,N_11977);
xor U12126 (N_12126,N_11432,N_11512);
nor U12127 (N_12127,N_11881,N_11733);
nor U12128 (N_12128,N_11427,N_11363);
or U12129 (N_12129,N_11314,N_11694);
and U12130 (N_12130,N_11737,N_11591);
or U12131 (N_12131,N_11975,N_11982);
nand U12132 (N_12132,N_11323,N_11513);
xnor U12133 (N_12133,N_11955,N_11284);
xor U12134 (N_12134,N_11483,N_11727);
xnor U12135 (N_12135,N_11812,N_11348);
nor U12136 (N_12136,N_11343,N_11340);
xnor U12137 (N_12137,N_11953,N_11334);
and U12138 (N_12138,N_11988,N_11517);
or U12139 (N_12139,N_11896,N_11666);
and U12140 (N_12140,N_11414,N_11942);
nand U12141 (N_12141,N_11632,N_11441);
and U12142 (N_12142,N_11980,N_11495);
and U12143 (N_12143,N_11537,N_11560);
or U12144 (N_12144,N_11505,N_11578);
and U12145 (N_12145,N_11652,N_11718);
and U12146 (N_12146,N_11270,N_11381);
or U12147 (N_12147,N_11302,N_11816);
xnor U12148 (N_12148,N_11253,N_11397);
or U12149 (N_12149,N_11697,N_11724);
xnor U12150 (N_12150,N_11368,N_11698);
xor U12151 (N_12151,N_11475,N_11946);
nand U12152 (N_12152,N_11431,N_11439);
and U12153 (N_12153,N_11653,N_11460);
nand U12154 (N_12154,N_11329,N_11633);
and U12155 (N_12155,N_11569,N_11396);
nand U12156 (N_12156,N_11950,N_11876);
nor U12157 (N_12157,N_11913,N_11893);
or U12158 (N_12158,N_11638,N_11754);
nand U12159 (N_12159,N_11954,N_11670);
and U12160 (N_12160,N_11979,N_11490);
nand U12161 (N_12161,N_11421,N_11996);
and U12162 (N_12162,N_11356,N_11690);
and U12163 (N_12163,N_11753,N_11592);
nand U12164 (N_12164,N_11380,N_11292);
nor U12165 (N_12165,N_11842,N_11699);
or U12166 (N_12166,N_11675,N_11787);
xnor U12167 (N_12167,N_11738,N_11586);
or U12168 (N_12168,N_11936,N_11654);
or U12169 (N_12169,N_11997,N_11532);
xor U12170 (N_12170,N_11442,N_11829);
xor U12171 (N_12171,N_11347,N_11470);
nand U12172 (N_12172,N_11405,N_11579);
and U12173 (N_12173,N_11882,N_11788);
nor U12174 (N_12174,N_11776,N_11572);
xor U12175 (N_12175,N_11634,N_11336);
nand U12176 (N_12176,N_11918,N_11728);
nor U12177 (N_12177,N_11767,N_11455);
nor U12178 (N_12178,N_11600,N_11723);
xor U12179 (N_12179,N_11663,N_11604);
nand U12180 (N_12180,N_11596,N_11393);
xor U12181 (N_12181,N_11903,N_11598);
nand U12182 (N_12182,N_11258,N_11928);
and U12183 (N_12183,N_11530,N_11813);
nand U12184 (N_12184,N_11894,N_11798);
nor U12185 (N_12185,N_11856,N_11566);
or U12186 (N_12186,N_11644,N_11970);
nand U12187 (N_12187,N_11924,N_11576);
and U12188 (N_12188,N_11677,N_11398);
xor U12189 (N_12189,N_11929,N_11321);
or U12190 (N_12190,N_11251,N_11944);
nor U12191 (N_12191,N_11852,N_11536);
nor U12192 (N_12192,N_11824,N_11333);
and U12193 (N_12193,N_11295,N_11267);
nor U12194 (N_12194,N_11995,N_11382);
xnor U12195 (N_12195,N_11376,N_11476);
xnor U12196 (N_12196,N_11349,N_11879);
or U12197 (N_12197,N_11623,N_11507);
nor U12198 (N_12198,N_11371,N_11282);
nor U12199 (N_12199,N_11263,N_11606);
or U12200 (N_12200,N_11900,N_11777);
and U12201 (N_12201,N_11916,N_11602);
and U12202 (N_12202,N_11335,N_11491);
nor U12203 (N_12203,N_11951,N_11751);
xor U12204 (N_12204,N_11581,N_11989);
and U12205 (N_12205,N_11803,N_11497);
or U12206 (N_12206,N_11287,N_11681);
nor U12207 (N_12207,N_11889,N_11484);
and U12208 (N_12208,N_11912,N_11923);
or U12209 (N_12209,N_11506,N_11562);
xnor U12210 (N_12210,N_11863,N_11486);
and U12211 (N_12211,N_11888,N_11802);
nor U12212 (N_12212,N_11420,N_11639);
and U12213 (N_12213,N_11554,N_11353);
nand U12214 (N_12214,N_11467,N_11687);
nor U12215 (N_12215,N_11784,N_11342);
xor U12216 (N_12216,N_11281,N_11793);
nand U12217 (N_12217,N_11926,N_11940);
nand U12218 (N_12218,N_11437,N_11529);
xor U12219 (N_12219,N_11309,N_11504);
or U12220 (N_12220,N_11704,N_11528);
and U12221 (N_12221,N_11413,N_11808);
or U12222 (N_12222,N_11543,N_11755);
xor U12223 (N_12223,N_11402,N_11584);
nor U12224 (N_12224,N_11945,N_11533);
xnor U12225 (N_12225,N_11452,N_11804);
and U12226 (N_12226,N_11541,N_11780);
xor U12227 (N_12227,N_11845,N_11841);
xnor U12228 (N_12228,N_11461,N_11702);
nor U12229 (N_12229,N_11436,N_11817);
and U12230 (N_12230,N_11428,N_11474);
nor U12231 (N_12231,N_11609,N_11910);
nand U12232 (N_12232,N_11647,N_11659);
nand U12233 (N_12233,N_11498,N_11276);
and U12234 (N_12234,N_11409,N_11547);
or U12235 (N_12235,N_11489,N_11805);
nand U12236 (N_12236,N_11905,N_11904);
or U12237 (N_12237,N_11673,N_11701);
and U12238 (N_12238,N_11865,N_11550);
or U12239 (N_12239,N_11354,N_11599);
nor U12240 (N_12240,N_11855,N_11481);
or U12241 (N_12241,N_11390,N_11919);
or U12242 (N_12242,N_11771,N_11648);
nand U12243 (N_12243,N_11293,N_11716);
nand U12244 (N_12244,N_11385,N_11313);
nor U12245 (N_12245,N_11290,N_11265);
or U12246 (N_12246,N_11286,N_11389);
and U12247 (N_12247,N_11789,N_11400);
or U12248 (N_12248,N_11911,N_11608);
nand U12249 (N_12249,N_11575,N_11294);
nand U12250 (N_12250,N_11635,N_11871);
or U12251 (N_12251,N_11374,N_11583);
and U12252 (N_12252,N_11846,N_11443);
or U12253 (N_12253,N_11503,N_11306);
and U12254 (N_12254,N_11907,N_11927);
and U12255 (N_12255,N_11696,N_11843);
and U12256 (N_12256,N_11752,N_11665);
nand U12257 (N_12257,N_11811,N_11272);
xnor U12258 (N_12258,N_11499,N_11836);
nor U12259 (N_12259,N_11649,N_11678);
nand U12260 (N_12260,N_11386,N_11424);
nor U12261 (N_12261,N_11612,N_11500);
nor U12262 (N_12262,N_11720,N_11304);
nor U12263 (N_12263,N_11778,N_11736);
and U12264 (N_12264,N_11341,N_11820);
or U12265 (N_12265,N_11307,N_11937);
and U12266 (N_12266,N_11450,N_11878);
nor U12267 (N_12267,N_11797,N_11459);
xnor U12268 (N_12268,N_11540,N_11959);
or U12269 (N_12269,N_11709,N_11359);
xor U12270 (N_12270,N_11440,N_11650);
nand U12271 (N_12271,N_11967,N_11721);
and U12272 (N_12272,N_11867,N_11961);
xor U12273 (N_12273,N_11545,N_11618);
or U12274 (N_12274,N_11403,N_11807);
nor U12275 (N_12275,N_11430,N_11932);
or U12276 (N_12276,N_11594,N_11330);
and U12277 (N_12277,N_11434,N_11418);
nor U12278 (N_12278,N_11853,N_11901);
nand U12279 (N_12279,N_11619,N_11252);
and U12280 (N_12280,N_11367,N_11883);
or U12281 (N_12281,N_11851,N_11556);
nand U12282 (N_12282,N_11668,N_11360);
nand U12283 (N_12283,N_11269,N_11850);
and U12284 (N_12284,N_11515,N_11454);
nand U12285 (N_12285,N_11345,N_11925);
nor U12286 (N_12286,N_11456,N_11411);
and U12287 (N_12287,N_11510,N_11658);
nand U12288 (N_12288,N_11707,N_11601);
and U12289 (N_12289,N_11408,N_11285);
xor U12290 (N_12290,N_11429,N_11760);
nand U12291 (N_12291,N_11522,N_11315);
nand U12292 (N_12292,N_11375,N_11766);
xnor U12293 (N_12293,N_11999,N_11565);
nand U12294 (N_12294,N_11898,N_11457);
nand U12295 (N_12295,N_11603,N_11864);
and U12296 (N_12296,N_11952,N_11496);
or U12297 (N_12297,N_11520,N_11383);
xnor U12298 (N_12298,N_11935,N_11279);
or U12299 (N_12299,N_11464,N_11682);
or U12300 (N_12300,N_11546,N_11561);
or U12301 (N_12301,N_11511,N_11857);
nor U12302 (N_12302,N_11799,N_11891);
nor U12303 (N_12303,N_11605,N_11629);
nand U12304 (N_12304,N_11254,N_11366);
nand U12305 (N_12305,N_11683,N_11987);
nor U12306 (N_12306,N_11662,N_11921);
xor U12307 (N_12307,N_11582,N_11750);
nor U12308 (N_12308,N_11337,N_11763);
or U12309 (N_12309,N_11391,N_11934);
and U12310 (N_12310,N_11641,N_11680);
or U12311 (N_12311,N_11744,N_11958);
and U12312 (N_12312,N_11832,N_11933);
and U12313 (N_12313,N_11426,N_11762);
and U12314 (N_12314,N_11548,N_11974);
or U12315 (N_12315,N_11379,N_11563);
xor U12316 (N_12316,N_11742,N_11364);
nor U12317 (N_12317,N_11880,N_11595);
or U12318 (N_12318,N_11326,N_11992);
or U12319 (N_12319,N_11956,N_11401);
or U12320 (N_12320,N_11941,N_11255);
nor U12321 (N_12321,N_11957,N_11384);
and U12322 (N_12322,N_11419,N_11357);
xor U12323 (N_12323,N_11303,N_11630);
nor U12324 (N_12324,N_11271,N_11438);
and U12325 (N_12325,N_11734,N_11445);
nand U12326 (N_12326,N_11963,N_11275);
and U12327 (N_12327,N_11758,N_11840);
and U12328 (N_12328,N_11821,N_11626);
and U12329 (N_12329,N_11943,N_11671);
or U12330 (N_12330,N_11624,N_11729);
nor U12331 (N_12331,N_11316,N_11573);
and U12332 (N_12332,N_11747,N_11468);
and U12333 (N_12333,N_11986,N_11740);
nor U12334 (N_12334,N_11700,N_11686);
or U12335 (N_12335,N_11795,N_11781);
and U12336 (N_12336,N_11571,N_11257);
and U12337 (N_12337,N_11544,N_11392);
nor U12338 (N_12338,N_11902,N_11985);
xnor U12339 (N_12339,N_11839,N_11412);
nand U12340 (N_12340,N_11833,N_11887);
nor U12341 (N_12341,N_11782,N_11628);
or U12342 (N_12342,N_11800,N_11549);
and U12343 (N_12343,N_11828,N_11469);
and U12344 (N_12344,N_11574,N_11312);
and U12345 (N_12345,N_11621,N_11465);
xnor U12346 (N_12346,N_11449,N_11317);
nand U12347 (N_12347,N_11972,N_11526);
nor U12348 (N_12348,N_11319,N_11651);
nand U12349 (N_12349,N_11848,N_11597);
nor U12350 (N_12350,N_11877,N_11899);
nand U12351 (N_12351,N_11297,N_11531);
nor U12352 (N_12352,N_11399,N_11296);
or U12353 (N_12353,N_11838,N_11895);
and U12354 (N_12354,N_11446,N_11525);
nor U12355 (N_12355,N_11551,N_11664);
xor U12356 (N_12356,N_11713,N_11361);
or U12357 (N_12357,N_11869,N_11872);
or U12358 (N_12358,N_11485,N_11679);
xor U12359 (N_12359,N_11920,N_11642);
xnor U12360 (N_12360,N_11930,N_11831);
nand U12361 (N_12361,N_11585,N_11725);
or U12362 (N_12362,N_11473,N_11407);
xor U12363 (N_12363,N_11365,N_11749);
xnor U12364 (N_12364,N_11745,N_11417);
nor U12365 (N_12365,N_11289,N_11559);
or U12366 (N_12366,N_11815,N_11786);
and U12367 (N_12367,N_11962,N_11283);
xnor U12368 (N_12368,N_11410,N_11298);
nand U12369 (N_12369,N_11993,N_11466);
xor U12370 (N_12370,N_11858,N_11717);
xor U12371 (N_12371,N_11732,N_11922);
or U12372 (N_12372,N_11577,N_11458);
xor U12373 (N_12373,N_11378,N_11640);
or U12374 (N_12374,N_11874,N_11735);
nor U12375 (N_12375,N_11581,N_11749);
or U12376 (N_12376,N_11680,N_11277);
nor U12377 (N_12377,N_11909,N_11937);
and U12378 (N_12378,N_11309,N_11990);
xnor U12379 (N_12379,N_11441,N_11273);
or U12380 (N_12380,N_11928,N_11753);
or U12381 (N_12381,N_11608,N_11432);
nand U12382 (N_12382,N_11974,N_11557);
or U12383 (N_12383,N_11719,N_11412);
xor U12384 (N_12384,N_11822,N_11909);
xnor U12385 (N_12385,N_11531,N_11473);
and U12386 (N_12386,N_11875,N_11977);
nor U12387 (N_12387,N_11860,N_11816);
nor U12388 (N_12388,N_11585,N_11559);
nand U12389 (N_12389,N_11977,N_11798);
and U12390 (N_12390,N_11952,N_11846);
nor U12391 (N_12391,N_11954,N_11466);
nand U12392 (N_12392,N_11319,N_11720);
xor U12393 (N_12393,N_11445,N_11603);
nand U12394 (N_12394,N_11762,N_11371);
nor U12395 (N_12395,N_11722,N_11650);
nor U12396 (N_12396,N_11958,N_11437);
nor U12397 (N_12397,N_11497,N_11368);
nand U12398 (N_12398,N_11945,N_11540);
or U12399 (N_12399,N_11710,N_11338);
xnor U12400 (N_12400,N_11827,N_11256);
nand U12401 (N_12401,N_11633,N_11862);
nand U12402 (N_12402,N_11941,N_11418);
nand U12403 (N_12403,N_11283,N_11781);
or U12404 (N_12404,N_11544,N_11311);
or U12405 (N_12405,N_11965,N_11894);
xor U12406 (N_12406,N_11371,N_11890);
and U12407 (N_12407,N_11313,N_11586);
or U12408 (N_12408,N_11487,N_11472);
and U12409 (N_12409,N_11984,N_11359);
nor U12410 (N_12410,N_11954,N_11431);
xnor U12411 (N_12411,N_11390,N_11927);
and U12412 (N_12412,N_11575,N_11493);
or U12413 (N_12413,N_11945,N_11806);
nor U12414 (N_12414,N_11479,N_11922);
and U12415 (N_12415,N_11998,N_11445);
nor U12416 (N_12416,N_11751,N_11831);
nand U12417 (N_12417,N_11292,N_11776);
nor U12418 (N_12418,N_11567,N_11997);
nor U12419 (N_12419,N_11654,N_11937);
and U12420 (N_12420,N_11644,N_11713);
nor U12421 (N_12421,N_11659,N_11263);
and U12422 (N_12422,N_11369,N_11904);
xnor U12423 (N_12423,N_11780,N_11855);
nor U12424 (N_12424,N_11943,N_11544);
nand U12425 (N_12425,N_11324,N_11613);
or U12426 (N_12426,N_11586,N_11359);
nor U12427 (N_12427,N_11913,N_11658);
nor U12428 (N_12428,N_11772,N_11775);
and U12429 (N_12429,N_11710,N_11838);
or U12430 (N_12430,N_11502,N_11758);
or U12431 (N_12431,N_11544,N_11666);
nor U12432 (N_12432,N_11895,N_11503);
and U12433 (N_12433,N_11822,N_11387);
nor U12434 (N_12434,N_11910,N_11839);
nor U12435 (N_12435,N_11282,N_11410);
or U12436 (N_12436,N_11665,N_11849);
or U12437 (N_12437,N_11672,N_11417);
and U12438 (N_12438,N_11418,N_11857);
xnor U12439 (N_12439,N_11600,N_11576);
or U12440 (N_12440,N_11864,N_11360);
nand U12441 (N_12441,N_11817,N_11495);
nand U12442 (N_12442,N_11632,N_11994);
nand U12443 (N_12443,N_11951,N_11634);
or U12444 (N_12444,N_11884,N_11581);
nand U12445 (N_12445,N_11869,N_11892);
nand U12446 (N_12446,N_11946,N_11516);
xnor U12447 (N_12447,N_11544,N_11724);
xnor U12448 (N_12448,N_11604,N_11901);
and U12449 (N_12449,N_11801,N_11524);
nand U12450 (N_12450,N_11975,N_11515);
xnor U12451 (N_12451,N_11256,N_11284);
nor U12452 (N_12452,N_11409,N_11814);
xnor U12453 (N_12453,N_11262,N_11263);
xnor U12454 (N_12454,N_11383,N_11369);
nand U12455 (N_12455,N_11357,N_11408);
xnor U12456 (N_12456,N_11355,N_11986);
and U12457 (N_12457,N_11641,N_11400);
nor U12458 (N_12458,N_11900,N_11659);
and U12459 (N_12459,N_11902,N_11285);
and U12460 (N_12460,N_11618,N_11524);
and U12461 (N_12461,N_11868,N_11815);
nand U12462 (N_12462,N_11721,N_11813);
xnor U12463 (N_12463,N_11747,N_11899);
nand U12464 (N_12464,N_11992,N_11447);
nand U12465 (N_12465,N_11562,N_11920);
and U12466 (N_12466,N_11822,N_11958);
nand U12467 (N_12467,N_11608,N_11639);
xor U12468 (N_12468,N_11274,N_11278);
nor U12469 (N_12469,N_11273,N_11594);
nor U12470 (N_12470,N_11762,N_11573);
and U12471 (N_12471,N_11884,N_11817);
nor U12472 (N_12472,N_11739,N_11679);
nor U12473 (N_12473,N_11649,N_11689);
nand U12474 (N_12474,N_11821,N_11892);
nor U12475 (N_12475,N_11693,N_11661);
xor U12476 (N_12476,N_11513,N_11796);
and U12477 (N_12477,N_11868,N_11607);
nor U12478 (N_12478,N_11966,N_11625);
nor U12479 (N_12479,N_11301,N_11657);
nor U12480 (N_12480,N_11497,N_11462);
nor U12481 (N_12481,N_11773,N_11739);
xor U12482 (N_12482,N_11273,N_11847);
xnor U12483 (N_12483,N_11870,N_11352);
nor U12484 (N_12484,N_11673,N_11353);
and U12485 (N_12485,N_11852,N_11978);
and U12486 (N_12486,N_11256,N_11921);
and U12487 (N_12487,N_11871,N_11649);
and U12488 (N_12488,N_11967,N_11547);
and U12489 (N_12489,N_11593,N_11837);
xor U12490 (N_12490,N_11674,N_11738);
or U12491 (N_12491,N_11557,N_11497);
nor U12492 (N_12492,N_11499,N_11837);
and U12493 (N_12493,N_11381,N_11742);
xnor U12494 (N_12494,N_11530,N_11805);
xor U12495 (N_12495,N_11754,N_11597);
xor U12496 (N_12496,N_11482,N_11406);
and U12497 (N_12497,N_11808,N_11773);
xor U12498 (N_12498,N_11957,N_11577);
and U12499 (N_12499,N_11551,N_11810);
or U12500 (N_12500,N_11524,N_11729);
nand U12501 (N_12501,N_11415,N_11811);
and U12502 (N_12502,N_11448,N_11766);
nand U12503 (N_12503,N_11763,N_11779);
or U12504 (N_12504,N_11728,N_11433);
or U12505 (N_12505,N_11286,N_11571);
xor U12506 (N_12506,N_11612,N_11291);
nor U12507 (N_12507,N_11470,N_11671);
or U12508 (N_12508,N_11647,N_11702);
and U12509 (N_12509,N_11965,N_11706);
nand U12510 (N_12510,N_11253,N_11363);
or U12511 (N_12511,N_11618,N_11578);
nor U12512 (N_12512,N_11691,N_11827);
and U12513 (N_12513,N_11811,N_11994);
xnor U12514 (N_12514,N_11483,N_11825);
and U12515 (N_12515,N_11342,N_11652);
or U12516 (N_12516,N_11284,N_11675);
nor U12517 (N_12517,N_11658,N_11502);
or U12518 (N_12518,N_11417,N_11687);
xor U12519 (N_12519,N_11309,N_11973);
xor U12520 (N_12520,N_11705,N_11551);
nor U12521 (N_12521,N_11738,N_11679);
xnor U12522 (N_12522,N_11904,N_11842);
nor U12523 (N_12523,N_11541,N_11813);
and U12524 (N_12524,N_11466,N_11796);
and U12525 (N_12525,N_11615,N_11562);
and U12526 (N_12526,N_11301,N_11996);
nand U12527 (N_12527,N_11913,N_11451);
nand U12528 (N_12528,N_11589,N_11945);
xnor U12529 (N_12529,N_11306,N_11452);
or U12530 (N_12530,N_11842,N_11611);
xor U12531 (N_12531,N_11930,N_11296);
and U12532 (N_12532,N_11827,N_11366);
xnor U12533 (N_12533,N_11506,N_11551);
nor U12534 (N_12534,N_11353,N_11944);
and U12535 (N_12535,N_11985,N_11441);
and U12536 (N_12536,N_11313,N_11291);
or U12537 (N_12537,N_11991,N_11343);
and U12538 (N_12538,N_11685,N_11382);
nand U12539 (N_12539,N_11533,N_11582);
nand U12540 (N_12540,N_11374,N_11386);
xor U12541 (N_12541,N_11463,N_11869);
or U12542 (N_12542,N_11831,N_11426);
nand U12543 (N_12543,N_11996,N_11464);
nor U12544 (N_12544,N_11442,N_11260);
nand U12545 (N_12545,N_11765,N_11763);
and U12546 (N_12546,N_11840,N_11495);
nor U12547 (N_12547,N_11655,N_11347);
and U12548 (N_12548,N_11984,N_11754);
and U12549 (N_12549,N_11816,N_11790);
nor U12550 (N_12550,N_11522,N_11634);
or U12551 (N_12551,N_11293,N_11648);
or U12552 (N_12552,N_11542,N_11478);
nand U12553 (N_12553,N_11750,N_11958);
and U12554 (N_12554,N_11853,N_11679);
or U12555 (N_12555,N_11872,N_11903);
nand U12556 (N_12556,N_11666,N_11721);
nand U12557 (N_12557,N_11587,N_11755);
nand U12558 (N_12558,N_11447,N_11373);
and U12559 (N_12559,N_11564,N_11819);
or U12560 (N_12560,N_11735,N_11897);
and U12561 (N_12561,N_11543,N_11851);
or U12562 (N_12562,N_11923,N_11584);
nand U12563 (N_12563,N_11681,N_11312);
and U12564 (N_12564,N_11765,N_11869);
or U12565 (N_12565,N_11985,N_11603);
and U12566 (N_12566,N_11441,N_11394);
xor U12567 (N_12567,N_11818,N_11599);
xor U12568 (N_12568,N_11868,N_11584);
nor U12569 (N_12569,N_11717,N_11709);
nand U12570 (N_12570,N_11775,N_11475);
nor U12571 (N_12571,N_11925,N_11855);
or U12572 (N_12572,N_11470,N_11395);
nand U12573 (N_12573,N_11947,N_11817);
and U12574 (N_12574,N_11837,N_11599);
nor U12575 (N_12575,N_11863,N_11282);
and U12576 (N_12576,N_11764,N_11258);
nor U12577 (N_12577,N_11260,N_11504);
or U12578 (N_12578,N_11614,N_11806);
or U12579 (N_12579,N_11583,N_11561);
nor U12580 (N_12580,N_11569,N_11432);
xor U12581 (N_12581,N_11775,N_11675);
nand U12582 (N_12582,N_11329,N_11855);
or U12583 (N_12583,N_11333,N_11648);
or U12584 (N_12584,N_11973,N_11251);
or U12585 (N_12585,N_11786,N_11285);
xor U12586 (N_12586,N_11395,N_11489);
nand U12587 (N_12587,N_11685,N_11432);
and U12588 (N_12588,N_11849,N_11503);
or U12589 (N_12589,N_11856,N_11491);
and U12590 (N_12590,N_11517,N_11597);
and U12591 (N_12591,N_11739,N_11821);
and U12592 (N_12592,N_11872,N_11946);
and U12593 (N_12593,N_11701,N_11288);
nor U12594 (N_12594,N_11893,N_11664);
nand U12595 (N_12595,N_11581,N_11362);
nor U12596 (N_12596,N_11681,N_11373);
and U12597 (N_12597,N_11794,N_11806);
or U12598 (N_12598,N_11927,N_11584);
nor U12599 (N_12599,N_11680,N_11844);
nand U12600 (N_12600,N_11884,N_11349);
or U12601 (N_12601,N_11307,N_11408);
or U12602 (N_12602,N_11686,N_11837);
and U12603 (N_12603,N_11326,N_11296);
or U12604 (N_12604,N_11537,N_11675);
and U12605 (N_12605,N_11974,N_11354);
or U12606 (N_12606,N_11876,N_11327);
nor U12607 (N_12607,N_11929,N_11737);
or U12608 (N_12608,N_11836,N_11857);
or U12609 (N_12609,N_11987,N_11643);
nor U12610 (N_12610,N_11532,N_11821);
xor U12611 (N_12611,N_11967,N_11352);
and U12612 (N_12612,N_11893,N_11773);
xnor U12613 (N_12613,N_11551,N_11805);
or U12614 (N_12614,N_11295,N_11958);
nor U12615 (N_12615,N_11383,N_11921);
nor U12616 (N_12616,N_11413,N_11625);
or U12617 (N_12617,N_11861,N_11307);
nor U12618 (N_12618,N_11562,N_11832);
xor U12619 (N_12619,N_11555,N_11310);
xnor U12620 (N_12620,N_11732,N_11650);
nand U12621 (N_12621,N_11555,N_11510);
nand U12622 (N_12622,N_11325,N_11629);
and U12623 (N_12623,N_11374,N_11548);
xnor U12624 (N_12624,N_11866,N_11913);
xnor U12625 (N_12625,N_11923,N_11580);
or U12626 (N_12626,N_11737,N_11946);
nand U12627 (N_12627,N_11623,N_11406);
or U12628 (N_12628,N_11902,N_11983);
nor U12629 (N_12629,N_11763,N_11434);
and U12630 (N_12630,N_11334,N_11920);
nor U12631 (N_12631,N_11798,N_11275);
or U12632 (N_12632,N_11784,N_11462);
and U12633 (N_12633,N_11701,N_11916);
and U12634 (N_12634,N_11866,N_11556);
nor U12635 (N_12635,N_11601,N_11911);
and U12636 (N_12636,N_11624,N_11559);
or U12637 (N_12637,N_11961,N_11875);
nor U12638 (N_12638,N_11941,N_11665);
nor U12639 (N_12639,N_11922,N_11369);
nand U12640 (N_12640,N_11592,N_11815);
or U12641 (N_12641,N_11570,N_11913);
and U12642 (N_12642,N_11803,N_11568);
nor U12643 (N_12643,N_11271,N_11856);
nand U12644 (N_12644,N_11296,N_11791);
nor U12645 (N_12645,N_11530,N_11514);
nand U12646 (N_12646,N_11493,N_11785);
or U12647 (N_12647,N_11743,N_11438);
or U12648 (N_12648,N_11489,N_11809);
nor U12649 (N_12649,N_11624,N_11496);
nand U12650 (N_12650,N_11425,N_11934);
xor U12651 (N_12651,N_11617,N_11931);
xor U12652 (N_12652,N_11819,N_11451);
and U12653 (N_12653,N_11293,N_11852);
nand U12654 (N_12654,N_11325,N_11640);
nand U12655 (N_12655,N_11481,N_11863);
and U12656 (N_12656,N_11944,N_11923);
or U12657 (N_12657,N_11744,N_11691);
and U12658 (N_12658,N_11543,N_11614);
and U12659 (N_12659,N_11342,N_11448);
xor U12660 (N_12660,N_11434,N_11631);
or U12661 (N_12661,N_11913,N_11740);
and U12662 (N_12662,N_11835,N_11785);
or U12663 (N_12663,N_11707,N_11975);
nor U12664 (N_12664,N_11560,N_11900);
and U12665 (N_12665,N_11951,N_11510);
or U12666 (N_12666,N_11513,N_11673);
or U12667 (N_12667,N_11354,N_11271);
nor U12668 (N_12668,N_11701,N_11677);
or U12669 (N_12669,N_11795,N_11784);
nor U12670 (N_12670,N_11306,N_11844);
nor U12671 (N_12671,N_11664,N_11480);
or U12672 (N_12672,N_11454,N_11842);
xnor U12673 (N_12673,N_11831,N_11382);
xor U12674 (N_12674,N_11987,N_11831);
nand U12675 (N_12675,N_11654,N_11445);
or U12676 (N_12676,N_11683,N_11933);
nand U12677 (N_12677,N_11600,N_11480);
xnor U12678 (N_12678,N_11478,N_11331);
nor U12679 (N_12679,N_11927,N_11618);
or U12680 (N_12680,N_11370,N_11254);
and U12681 (N_12681,N_11589,N_11879);
and U12682 (N_12682,N_11733,N_11712);
xor U12683 (N_12683,N_11261,N_11451);
nor U12684 (N_12684,N_11732,N_11440);
nand U12685 (N_12685,N_11275,N_11988);
or U12686 (N_12686,N_11336,N_11986);
nor U12687 (N_12687,N_11909,N_11575);
and U12688 (N_12688,N_11270,N_11483);
nand U12689 (N_12689,N_11806,N_11569);
and U12690 (N_12690,N_11845,N_11935);
nand U12691 (N_12691,N_11953,N_11799);
or U12692 (N_12692,N_11456,N_11826);
xor U12693 (N_12693,N_11263,N_11971);
xnor U12694 (N_12694,N_11889,N_11589);
nor U12695 (N_12695,N_11837,N_11681);
or U12696 (N_12696,N_11365,N_11650);
xor U12697 (N_12697,N_11455,N_11954);
and U12698 (N_12698,N_11641,N_11872);
nor U12699 (N_12699,N_11715,N_11916);
nor U12700 (N_12700,N_11545,N_11626);
nand U12701 (N_12701,N_11466,N_11699);
xnor U12702 (N_12702,N_11289,N_11777);
or U12703 (N_12703,N_11990,N_11361);
nor U12704 (N_12704,N_11350,N_11766);
nor U12705 (N_12705,N_11768,N_11859);
or U12706 (N_12706,N_11988,N_11655);
or U12707 (N_12707,N_11464,N_11803);
nand U12708 (N_12708,N_11656,N_11655);
xnor U12709 (N_12709,N_11253,N_11358);
xnor U12710 (N_12710,N_11436,N_11294);
nor U12711 (N_12711,N_11393,N_11877);
or U12712 (N_12712,N_11738,N_11524);
xor U12713 (N_12713,N_11761,N_11491);
nand U12714 (N_12714,N_11811,N_11281);
xnor U12715 (N_12715,N_11448,N_11651);
xnor U12716 (N_12716,N_11651,N_11792);
or U12717 (N_12717,N_11478,N_11523);
nor U12718 (N_12718,N_11711,N_11951);
nand U12719 (N_12719,N_11694,N_11443);
nor U12720 (N_12720,N_11958,N_11612);
and U12721 (N_12721,N_11969,N_11621);
xnor U12722 (N_12722,N_11522,N_11842);
or U12723 (N_12723,N_11633,N_11898);
or U12724 (N_12724,N_11737,N_11559);
nor U12725 (N_12725,N_11869,N_11506);
nand U12726 (N_12726,N_11867,N_11694);
or U12727 (N_12727,N_11588,N_11946);
xor U12728 (N_12728,N_11962,N_11635);
or U12729 (N_12729,N_11800,N_11632);
or U12730 (N_12730,N_11741,N_11255);
xor U12731 (N_12731,N_11719,N_11883);
or U12732 (N_12732,N_11441,N_11872);
xor U12733 (N_12733,N_11806,N_11423);
nor U12734 (N_12734,N_11524,N_11955);
nor U12735 (N_12735,N_11512,N_11495);
and U12736 (N_12736,N_11792,N_11333);
xnor U12737 (N_12737,N_11874,N_11317);
or U12738 (N_12738,N_11284,N_11820);
nand U12739 (N_12739,N_11361,N_11297);
or U12740 (N_12740,N_11836,N_11270);
nor U12741 (N_12741,N_11665,N_11801);
nand U12742 (N_12742,N_11947,N_11316);
or U12743 (N_12743,N_11721,N_11587);
xnor U12744 (N_12744,N_11955,N_11892);
and U12745 (N_12745,N_11559,N_11388);
and U12746 (N_12746,N_11420,N_11584);
nor U12747 (N_12747,N_11479,N_11256);
and U12748 (N_12748,N_11370,N_11772);
and U12749 (N_12749,N_11496,N_11942);
and U12750 (N_12750,N_12173,N_12326);
and U12751 (N_12751,N_12148,N_12297);
xor U12752 (N_12752,N_12083,N_12645);
nor U12753 (N_12753,N_12348,N_12282);
or U12754 (N_12754,N_12335,N_12113);
and U12755 (N_12755,N_12685,N_12046);
or U12756 (N_12756,N_12548,N_12584);
or U12757 (N_12757,N_12712,N_12510);
or U12758 (N_12758,N_12183,N_12618);
nor U12759 (N_12759,N_12040,N_12306);
xor U12760 (N_12760,N_12150,N_12342);
and U12761 (N_12761,N_12216,N_12539);
nor U12762 (N_12762,N_12709,N_12707);
or U12763 (N_12763,N_12270,N_12341);
and U12764 (N_12764,N_12455,N_12069);
xor U12765 (N_12765,N_12118,N_12219);
nor U12766 (N_12766,N_12346,N_12401);
or U12767 (N_12767,N_12290,N_12375);
and U12768 (N_12768,N_12668,N_12655);
and U12769 (N_12769,N_12347,N_12314);
nand U12770 (N_12770,N_12543,N_12585);
xnor U12771 (N_12771,N_12280,N_12354);
nand U12772 (N_12772,N_12467,N_12649);
nand U12773 (N_12773,N_12312,N_12728);
nor U12774 (N_12774,N_12020,N_12513);
or U12775 (N_12775,N_12094,N_12378);
xnor U12776 (N_12776,N_12090,N_12582);
and U12777 (N_12777,N_12719,N_12405);
nand U12778 (N_12778,N_12363,N_12505);
or U12779 (N_12779,N_12286,N_12334);
or U12780 (N_12780,N_12576,N_12070);
xnor U12781 (N_12781,N_12678,N_12053);
or U12782 (N_12782,N_12367,N_12608);
xnor U12783 (N_12783,N_12450,N_12134);
or U12784 (N_12784,N_12005,N_12635);
nand U12785 (N_12785,N_12609,N_12267);
nand U12786 (N_12786,N_12708,N_12139);
xor U12787 (N_12787,N_12742,N_12396);
xnor U12788 (N_12788,N_12288,N_12079);
nor U12789 (N_12789,N_12594,N_12688);
xnor U12790 (N_12790,N_12397,N_12037);
or U12791 (N_12791,N_12032,N_12263);
or U12792 (N_12792,N_12460,N_12462);
or U12793 (N_12793,N_12366,N_12089);
nand U12794 (N_12794,N_12640,N_12222);
xnor U12795 (N_12795,N_12650,N_12019);
xnor U12796 (N_12796,N_12036,N_12107);
xnor U12797 (N_12797,N_12112,N_12411);
nand U12798 (N_12798,N_12319,N_12471);
xor U12799 (N_12799,N_12558,N_12238);
nor U12800 (N_12800,N_12181,N_12457);
and U12801 (N_12801,N_12295,N_12063);
xor U12802 (N_12802,N_12161,N_12338);
nor U12803 (N_12803,N_12591,N_12184);
nand U12804 (N_12804,N_12525,N_12500);
and U12805 (N_12805,N_12159,N_12062);
and U12806 (N_12806,N_12452,N_12209);
nor U12807 (N_12807,N_12430,N_12221);
nand U12808 (N_12808,N_12541,N_12661);
or U12809 (N_12809,N_12512,N_12377);
xor U12810 (N_12810,N_12738,N_12628);
nand U12811 (N_12811,N_12061,N_12516);
or U12812 (N_12812,N_12566,N_12615);
xnor U12813 (N_12813,N_12749,N_12489);
nand U12814 (N_12814,N_12553,N_12402);
or U12815 (N_12815,N_12469,N_12085);
nand U12816 (N_12816,N_12379,N_12514);
nor U12817 (N_12817,N_12440,N_12013);
and U12818 (N_12818,N_12117,N_12507);
nand U12819 (N_12819,N_12317,N_12185);
or U12820 (N_12820,N_12284,N_12435);
or U12821 (N_12821,N_12350,N_12621);
or U12822 (N_12822,N_12670,N_12413);
xor U12823 (N_12823,N_12601,N_12527);
and U12824 (N_12824,N_12333,N_12177);
nand U12825 (N_12825,N_12162,N_12357);
nand U12826 (N_12826,N_12307,N_12551);
or U12827 (N_12827,N_12245,N_12001);
or U12828 (N_12828,N_12065,N_12540);
nor U12829 (N_12829,N_12477,N_12081);
nor U12830 (N_12830,N_12140,N_12074);
and U12831 (N_12831,N_12138,N_12100);
or U12832 (N_12832,N_12508,N_12592);
nand U12833 (N_12833,N_12011,N_12544);
and U12834 (N_12834,N_12362,N_12538);
or U12835 (N_12835,N_12646,N_12017);
nor U12836 (N_12836,N_12250,N_12285);
nand U12837 (N_12837,N_12436,N_12213);
nor U12838 (N_12838,N_12547,N_12108);
nor U12839 (N_12839,N_12021,N_12671);
xnor U12840 (N_12840,N_12364,N_12748);
nor U12841 (N_12841,N_12648,N_12523);
xor U12842 (N_12842,N_12111,N_12724);
nor U12843 (N_12843,N_12515,N_12497);
xnor U12844 (N_12844,N_12392,N_12277);
and U12845 (N_12845,N_12071,N_12399);
nor U12846 (N_12846,N_12101,N_12410);
and U12847 (N_12847,N_12681,N_12394);
or U12848 (N_12848,N_12522,N_12642);
nor U12849 (N_12849,N_12320,N_12204);
nor U12850 (N_12850,N_12662,N_12116);
nand U12851 (N_12851,N_12234,N_12494);
nand U12852 (N_12852,N_12704,N_12199);
or U12853 (N_12853,N_12524,N_12043);
nor U12854 (N_12854,N_12291,N_12487);
or U12855 (N_12855,N_12151,N_12491);
nand U12856 (N_12856,N_12360,N_12745);
nand U12857 (N_12857,N_12192,N_12431);
xnor U12858 (N_12858,N_12137,N_12684);
xnor U12859 (N_12859,N_12387,N_12196);
xor U12860 (N_12860,N_12301,N_12128);
and U12861 (N_12861,N_12024,N_12673);
nor U12862 (N_12862,N_12235,N_12537);
nor U12863 (N_12863,N_12168,N_12262);
nor U12864 (N_12864,N_12230,N_12419);
and U12865 (N_12865,N_12501,N_12638);
nand U12866 (N_12866,N_12453,N_12389);
xnor U12867 (N_12867,N_12526,N_12122);
nand U12868 (N_12868,N_12374,N_12518);
or U12869 (N_12869,N_12143,N_12373);
xor U12870 (N_12870,N_12049,N_12265);
and U12871 (N_12871,N_12310,N_12266);
xor U12872 (N_12872,N_12016,N_12302);
xor U12873 (N_12873,N_12579,N_12602);
xnor U12874 (N_12874,N_12051,N_12495);
or U12875 (N_12875,N_12400,N_12075);
nor U12876 (N_12876,N_12099,N_12686);
nand U12877 (N_12877,N_12126,N_12597);
xnor U12878 (N_12878,N_12643,N_12690);
nor U12879 (N_12879,N_12329,N_12653);
nand U12880 (N_12880,N_12479,N_12569);
and U12881 (N_12881,N_12123,N_12251);
and U12882 (N_12882,N_12182,N_12422);
nand U12883 (N_12883,N_12004,N_12466);
and U12884 (N_12884,N_12458,N_12355);
and U12885 (N_12885,N_12088,N_12743);
or U12886 (N_12886,N_12395,N_12694);
xor U12887 (N_12887,N_12672,N_12322);
and U12888 (N_12888,N_12275,N_12598);
and U12889 (N_12889,N_12502,N_12141);
and U12890 (N_12890,N_12097,N_12664);
and U12891 (N_12891,N_12246,N_12571);
or U12892 (N_12892,N_12003,N_12142);
nand U12893 (N_12893,N_12157,N_12393);
or U12894 (N_12894,N_12178,N_12059);
nor U12895 (N_12895,N_12272,N_12388);
nor U12896 (N_12896,N_12381,N_12589);
nor U12897 (N_12897,N_12474,N_12189);
and U12898 (N_12898,N_12416,N_12084);
xor U12899 (N_12899,N_12736,N_12368);
or U12900 (N_12900,N_12190,N_12327);
nand U12901 (N_12901,N_12535,N_12560);
xnor U12902 (N_12902,N_12677,N_12703);
nor U12903 (N_12903,N_12220,N_12693);
and U12904 (N_12904,N_12146,N_12697);
or U12905 (N_12905,N_12133,N_12439);
or U12906 (N_12906,N_12232,N_12689);
and U12907 (N_12907,N_12634,N_12247);
and U12908 (N_12908,N_12441,N_12421);
and U12909 (N_12909,N_12570,N_12606);
and U12910 (N_12910,N_12531,N_12371);
nor U12911 (N_12911,N_12241,N_12418);
xnor U12912 (N_12912,N_12098,N_12057);
or U12913 (N_12913,N_12336,N_12666);
xnor U12914 (N_12914,N_12156,N_12580);
xnor U12915 (N_12915,N_12176,N_12136);
and U12916 (N_12916,N_12741,N_12563);
nand U12917 (N_12917,N_12587,N_12506);
xnor U12918 (N_12918,N_12659,N_12404);
or U12919 (N_12919,N_12055,N_12164);
nor U12920 (N_12920,N_12493,N_12415);
xor U12921 (N_12921,N_12165,N_12574);
nand U12922 (N_12922,N_12746,N_12554);
nand U12923 (N_12923,N_12242,N_12706);
nand U12924 (N_12924,N_12503,N_12729);
nand U12925 (N_12925,N_12412,N_12039);
nand U12926 (N_12926,N_12533,N_12682);
or U12927 (N_12927,N_12031,N_12068);
or U12928 (N_12928,N_12468,N_12044);
or U12929 (N_12929,N_12721,N_12244);
nor U12930 (N_12930,N_12391,N_12384);
xnor U12931 (N_12931,N_12720,N_12619);
xor U12932 (N_12932,N_12289,N_12734);
xnor U12933 (N_12933,N_12353,N_12432);
nor U12934 (N_12934,N_12376,N_12279);
xor U12935 (N_12935,N_12739,N_12253);
nand U12936 (N_12936,N_12683,N_12027);
or U12937 (N_12937,N_12517,N_12464);
nor U12938 (N_12938,N_12022,N_12331);
xor U12939 (N_12939,N_12237,N_12313);
nand U12940 (N_12940,N_12293,N_12488);
and U12941 (N_12941,N_12365,N_12713);
or U12942 (N_12942,N_12603,N_12008);
nand U12943 (N_12943,N_12042,N_12675);
and U12944 (N_12944,N_12731,N_12076);
and U12945 (N_12945,N_12700,N_12718);
and U12946 (N_12946,N_12604,N_12105);
or U12947 (N_12947,N_12264,N_12459);
or U12948 (N_12948,N_12425,N_12131);
or U12949 (N_12949,N_12552,N_12252);
nor U12950 (N_12950,N_12472,N_12239);
and U12951 (N_12951,N_12147,N_12740);
nand U12952 (N_12952,N_12733,N_12448);
xnor U12953 (N_12953,N_12248,N_12730);
or U12954 (N_12954,N_12722,N_12532);
and U12955 (N_12955,N_12296,N_12191);
nand U12956 (N_12956,N_12470,N_12260);
nor U12957 (N_12957,N_12723,N_12328);
and U12958 (N_12958,N_12186,N_12356);
or U12959 (N_12959,N_12417,N_12613);
xor U12960 (N_12960,N_12129,N_12298);
nand U12961 (N_12961,N_12054,N_12194);
nand U12962 (N_12962,N_12434,N_12485);
or U12963 (N_12963,N_12224,N_12406);
nand U12964 (N_12964,N_12195,N_12067);
nand U12965 (N_12965,N_12163,N_12386);
or U12966 (N_12966,N_12701,N_12259);
nor U12967 (N_12967,N_12599,N_12256);
and U12968 (N_12968,N_12035,N_12620);
nor U12969 (N_12969,N_12233,N_12398);
xor U12970 (N_12970,N_12261,N_12390);
nand U12971 (N_12971,N_12114,N_12130);
nand U12972 (N_12972,N_12145,N_12294);
or U12973 (N_12973,N_12581,N_12408);
nand U12974 (N_12974,N_12343,N_12271);
and U12975 (N_12975,N_12172,N_12211);
and U12976 (N_12976,N_12125,N_12546);
and U12977 (N_12977,N_12486,N_12476);
or U12978 (N_12978,N_12616,N_12166);
and U12979 (N_12979,N_12473,N_12499);
nand U12980 (N_12980,N_12443,N_12337);
nor U12981 (N_12981,N_12715,N_12567);
nor U12982 (N_12982,N_12498,N_12015);
and U12983 (N_12983,N_12292,N_12249);
or U12984 (N_12984,N_12636,N_12352);
nand U12985 (N_12985,N_12324,N_12660);
and U12986 (N_12986,N_12691,N_12323);
xor U12987 (N_12987,N_12197,N_12727);
xor U12988 (N_12988,N_12300,N_12456);
and U12989 (N_12989,N_12345,N_12573);
and U12990 (N_12990,N_12096,N_12536);
or U12991 (N_12991,N_12575,N_12451);
and U12992 (N_12992,N_12654,N_12236);
nand U12993 (N_12993,N_12315,N_12617);
or U12994 (N_12994,N_12429,N_12696);
xnor U12995 (N_12995,N_12454,N_12257);
nor U12996 (N_12996,N_12612,N_12283);
nand U12997 (N_12997,N_12590,N_12254);
and U12998 (N_12998,N_12647,N_12446);
xor U12999 (N_12999,N_12167,N_12577);
and U13000 (N_13000,N_12370,N_12680);
nor U13001 (N_13001,N_12534,N_12135);
nand U13002 (N_13002,N_12461,N_12086);
and U13003 (N_13003,N_12409,N_12308);
or U13004 (N_13004,N_12110,N_12311);
nand U13005 (N_13005,N_12465,N_12132);
xnor U13006 (N_13006,N_12622,N_12383);
and U13007 (N_13007,N_12009,N_12007);
and U13008 (N_13008,N_12578,N_12564);
nor U13009 (N_13009,N_12339,N_12644);
and U13010 (N_13010,N_12492,N_12205);
nand U13011 (N_13011,N_12714,N_12407);
nor U13012 (N_13012,N_12657,N_12447);
nor U13013 (N_13013,N_12332,N_12278);
and U13014 (N_13014,N_12705,N_12382);
nor U13015 (N_13015,N_12153,N_12014);
and U13016 (N_13016,N_12056,N_12632);
nor U13017 (N_13017,N_12509,N_12041);
xor U13018 (N_13018,N_12152,N_12426);
nor U13019 (N_13019,N_12025,N_12427);
or U13020 (N_13020,N_12633,N_12223);
or U13021 (N_13021,N_12218,N_12351);
or U13022 (N_13022,N_12530,N_12160);
and U13023 (N_13023,N_12193,N_12018);
nand U13024 (N_13024,N_12309,N_12208);
nand U13025 (N_13025,N_12607,N_12103);
or U13026 (N_13026,N_12428,N_12026);
xnor U13027 (N_13027,N_12542,N_12669);
nor U13028 (N_13028,N_12630,N_12318);
nand U13029 (N_13029,N_12087,N_12073);
xor U13030 (N_13030,N_12048,N_12359);
xor U13031 (N_13031,N_12414,N_12202);
and U13032 (N_13032,N_12325,N_12033);
xor U13033 (N_13033,N_12545,N_12679);
or U13034 (N_13034,N_12115,N_12529);
xor U13035 (N_13035,N_12699,N_12303);
nor U13036 (N_13036,N_12231,N_12735);
nor U13037 (N_13037,N_12212,N_12344);
and U13038 (N_13038,N_12268,N_12747);
and U13039 (N_13039,N_12188,N_12667);
nor U13040 (N_13040,N_12207,N_12000);
or U13041 (N_13041,N_12170,N_12050);
and U13042 (N_13042,N_12504,N_12002);
and U13043 (N_13043,N_12556,N_12559);
or U13044 (N_13044,N_12144,N_12445);
or U13045 (N_13045,N_12652,N_12555);
nor U13046 (N_13046,N_12586,N_12521);
xor U13047 (N_13047,N_12483,N_12732);
nor U13048 (N_13048,N_12561,N_12060);
and U13049 (N_13049,N_12120,N_12149);
nand U13050 (N_13050,N_12225,N_12449);
and U13051 (N_13051,N_12726,N_12091);
nor U13052 (N_13052,N_12478,N_12169);
nand U13053 (N_13053,N_12385,N_12519);
or U13054 (N_13054,N_12258,N_12358);
nand U13055 (N_13055,N_12692,N_12058);
nand U13056 (N_13056,N_12305,N_12716);
or U13057 (N_13057,N_12595,N_12281);
and U13058 (N_13058,N_12611,N_12361);
xnor U13059 (N_13059,N_12124,N_12349);
xor U13060 (N_13060,N_12201,N_12442);
xnor U13061 (N_13061,N_12121,N_12276);
xor U13062 (N_13062,N_12010,N_12217);
and U13063 (N_13063,N_12095,N_12102);
nor U13064 (N_13064,N_12064,N_12206);
or U13065 (N_13065,N_12629,N_12656);
and U13066 (N_13066,N_12484,N_12380);
or U13067 (N_13067,N_12226,N_12154);
and U13068 (N_13068,N_12725,N_12287);
and U13069 (N_13069,N_12463,N_12711);
nor U13070 (N_13070,N_12420,N_12127);
nor U13071 (N_13071,N_12610,N_12369);
xor U13072 (N_13072,N_12180,N_12623);
or U13073 (N_13073,N_12562,N_12593);
nor U13074 (N_13074,N_12023,N_12475);
nand U13075 (N_13075,N_12480,N_12304);
and U13076 (N_13076,N_12744,N_12274);
nor U13077 (N_13077,N_12424,N_12482);
and U13078 (N_13078,N_12078,N_12052);
xnor U13079 (N_13079,N_12109,N_12082);
xor U13080 (N_13080,N_12437,N_12717);
nor U13081 (N_13081,N_12549,N_12698);
or U13082 (N_13082,N_12030,N_12077);
and U13083 (N_13083,N_12340,N_12511);
xnor U13084 (N_13084,N_12588,N_12528);
or U13085 (N_13085,N_12203,N_12372);
nor U13086 (N_13086,N_12210,N_12158);
or U13087 (N_13087,N_12243,N_12229);
xor U13088 (N_13088,N_12093,N_12155);
nor U13089 (N_13089,N_12106,N_12423);
nor U13090 (N_13090,N_12737,N_12029);
nor U13091 (N_13091,N_12600,N_12045);
nand U13092 (N_13092,N_12072,N_12695);
xnor U13093 (N_13093,N_12012,N_12006);
or U13094 (N_13094,N_12174,N_12710);
and U13095 (N_13095,N_12625,N_12490);
and U13096 (N_13096,N_12641,N_12215);
xnor U13097 (N_13097,N_12066,N_12028);
and U13098 (N_13098,N_12572,N_12038);
nor U13099 (N_13099,N_12702,N_12631);
nor U13100 (N_13100,N_12047,N_12228);
and U13101 (N_13101,N_12321,N_12583);
xor U13102 (N_13102,N_12557,N_12674);
nand U13103 (N_13103,N_12624,N_12104);
nand U13104 (N_13104,N_12240,N_12676);
or U13105 (N_13105,N_12175,N_12651);
and U13106 (N_13106,N_12316,N_12269);
or U13107 (N_13107,N_12687,N_12626);
nor U13108 (N_13108,N_12171,N_12200);
nor U13109 (N_13109,N_12255,N_12214);
nor U13110 (N_13110,N_12568,N_12179);
and U13111 (N_13111,N_12614,N_12665);
xnor U13112 (N_13112,N_12119,N_12444);
and U13113 (N_13113,N_12627,N_12481);
xnor U13114 (N_13114,N_12187,N_12520);
nand U13115 (N_13115,N_12273,N_12330);
and U13116 (N_13116,N_12092,N_12080);
nor U13117 (N_13117,N_12639,N_12550);
nor U13118 (N_13118,N_12227,N_12565);
nand U13119 (N_13119,N_12198,N_12637);
nand U13120 (N_13120,N_12403,N_12605);
xor U13121 (N_13121,N_12034,N_12596);
or U13122 (N_13122,N_12496,N_12658);
xnor U13123 (N_13123,N_12438,N_12663);
and U13124 (N_13124,N_12299,N_12433);
or U13125 (N_13125,N_12447,N_12736);
xor U13126 (N_13126,N_12541,N_12697);
nand U13127 (N_13127,N_12587,N_12097);
nor U13128 (N_13128,N_12038,N_12183);
or U13129 (N_13129,N_12289,N_12355);
or U13130 (N_13130,N_12561,N_12305);
or U13131 (N_13131,N_12734,N_12381);
nand U13132 (N_13132,N_12491,N_12270);
nand U13133 (N_13133,N_12643,N_12414);
xnor U13134 (N_13134,N_12087,N_12216);
and U13135 (N_13135,N_12298,N_12438);
nand U13136 (N_13136,N_12367,N_12743);
and U13137 (N_13137,N_12290,N_12190);
xor U13138 (N_13138,N_12344,N_12071);
or U13139 (N_13139,N_12653,N_12555);
and U13140 (N_13140,N_12388,N_12697);
nor U13141 (N_13141,N_12001,N_12234);
xnor U13142 (N_13142,N_12090,N_12149);
nand U13143 (N_13143,N_12113,N_12656);
or U13144 (N_13144,N_12293,N_12662);
nand U13145 (N_13145,N_12010,N_12124);
xor U13146 (N_13146,N_12337,N_12012);
and U13147 (N_13147,N_12474,N_12608);
nand U13148 (N_13148,N_12171,N_12507);
nand U13149 (N_13149,N_12615,N_12339);
xnor U13150 (N_13150,N_12072,N_12223);
nor U13151 (N_13151,N_12518,N_12133);
nand U13152 (N_13152,N_12270,N_12726);
or U13153 (N_13153,N_12324,N_12458);
and U13154 (N_13154,N_12252,N_12215);
nand U13155 (N_13155,N_12286,N_12083);
xor U13156 (N_13156,N_12662,N_12604);
and U13157 (N_13157,N_12566,N_12118);
xor U13158 (N_13158,N_12182,N_12526);
and U13159 (N_13159,N_12605,N_12662);
nor U13160 (N_13160,N_12255,N_12239);
and U13161 (N_13161,N_12228,N_12029);
nand U13162 (N_13162,N_12450,N_12183);
and U13163 (N_13163,N_12293,N_12262);
xor U13164 (N_13164,N_12340,N_12570);
or U13165 (N_13165,N_12703,N_12625);
and U13166 (N_13166,N_12303,N_12701);
nor U13167 (N_13167,N_12442,N_12323);
xnor U13168 (N_13168,N_12207,N_12714);
xnor U13169 (N_13169,N_12380,N_12096);
nand U13170 (N_13170,N_12695,N_12369);
nor U13171 (N_13171,N_12150,N_12204);
nand U13172 (N_13172,N_12462,N_12556);
and U13173 (N_13173,N_12068,N_12369);
nor U13174 (N_13174,N_12466,N_12643);
and U13175 (N_13175,N_12229,N_12707);
or U13176 (N_13176,N_12437,N_12436);
nor U13177 (N_13177,N_12168,N_12428);
and U13178 (N_13178,N_12046,N_12578);
nand U13179 (N_13179,N_12682,N_12011);
and U13180 (N_13180,N_12727,N_12531);
xor U13181 (N_13181,N_12350,N_12630);
or U13182 (N_13182,N_12699,N_12508);
nor U13183 (N_13183,N_12482,N_12233);
xor U13184 (N_13184,N_12737,N_12309);
or U13185 (N_13185,N_12082,N_12674);
nor U13186 (N_13186,N_12485,N_12170);
xnor U13187 (N_13187,N_12240,N_12316);
nor U13188 (N_13188,N_12140,N_12410);
nand U13189 (N_13189,N_12464,N_12573);
nand U13190 (N_13190,N_12536,N_12685);
or U13191 (N_13191,N_12282,N_12675);
nor U13192 (N_13192,N_12289,N_12684);
nor U13193 (N_13193,N_12086,N_12400);
nor U13194 (N_13194,N_12203,N_12299);
xnor U13195 (N_13195,N_12670,N_12067);
and U13196 (N_13196,N_12593,N_12172);
xnor U13197 (N_13197,N_12460,N_12516);
or U13198 (N_13198,N_12677,N_12125);
and U13199 (N_13199,N_12538,N_12676);
or U13200 (N_13200,N_12199,N_12598);
nor U13201 (N_13201,N_12366,N_12254);
xnor U13202 (N_13202,N_12413,N_12152);
nand U13203 (N_13203,N_12399,N_12646);
and U13204 (N_13204,N_12097,N_12447);
xor U13205 (N_13205,N_12271,N_12577);
nor U13206 (N_13206,N_12574,N_12090);
and U13207 (N_13207,N_12046,N_12612);
xnor U13208 (N_13208,N_12295,N_12666);
nor U13209 (N_13209,N_12720,N_12402);
nor U13210 (N_13210,N_12383,N_12343);
or U13211 (N_13211,N_12707,N_12688);
and U13212 (N_13212,N_12120,N_12119);
and U13213 (N_13213,N_12047,N_12642);
and U13214 (N_13214,N_12113,N_12083);
nand U13215 (N_13215,N_12551,N_12036);
xor U13216 (N_13216,N_12124,N_12217);
nor U13217 (N_13217,N_12110,N_12255);
xor U13218 (N_13218,N_12328,N_12203);
or U13219 (N_13219,N_12632,N_12657);
nand U13220 (N_13220,N_12678,N_12509);
nand U13221 (N_13221,N_12073,N_12519);
xnor U13222 (N_13222,N_12178,N_12550);
xnor U13223 (N_13223,N_12147,N_12264);
or U13224 (N_13224,N_12263,N_12021);
or U13225 (N_13225,N_12546,N_12638);
nor U13226 (N_13226,N_12024,N_12430);
and U13227 (N_13227,N_12240,N_12112);
nor U13228 (N_13228,N_12020,N_12300);
xnor U13229 (N_13229,N_12415,N_12725);
and U13230 (N_13230,N_12572,N_12722);
nand U13231 (N_13231,N_12456,N_12003);
and U13232 (N_13232,N_12644,N_12262);
and U13233 (N_13233,N_12455,N_12397);
xor U13234 (N_13234,N_12385,N_12178);
nand U13235 (N_13235,N_12043,N_12222);
and U13236 (N_13236,N_12489,N_12105);
and U13237 (N_13237,N_12033,N_12268);
xor U13238 (N_13238,N_12595,N_12103);
nand U13239 (N_13239,N_12259,N_12571);
xor U13240 (N_13240,N_12172,N_12148);
xor U13241 (N_13241,N_12329,N_12665);
and U13242 (N_13242,N_12267,N_12725);
or U13243 (N_13243,N_12403,N_12292);
nand U13244 (N_13244,N_12687,N_12368);
xnor U13245 (N_13245,N_12664,N_12619);
nand U13246 (N_13246,N_12666,N_12072);
nor U13247 (N_13247,N_12288,N_12361);
and U13248 (N_13248,N_12359,N_12266);
nand U13249 (N_13249,N_12321,N_12460);
or U13250 (N_13250,N_12121,N_12716);
xor U13251 (N_13251,N_12636,N_12222);
xnor U13252 (N_13252,N_12367,N_12313);
nand U13253 (N_13253,N_12626,N_12412);
nand U13254 (N_13254,N_12086,N_12285);
xor U13255 (N_13255,N_12474,N_12618);
nor U13256 (N_13256,N_12067,N_12193);
or U13257 (N_13257,N_12204,N_12738);
xor U13258 (N_13258,N_12699,N_12467);
and U13259 (N_13259,N_12518,N_12150);
and U13260 (N_13260,N_12584,N_12708);
or U13261 (N_13261,N_12605,N_12352);
nor U13262 (N_13262,N_12190,N_12450);
xor U13263 (N_13263,N_12120,N_12037);
or U13264 (N_13264,N_12413,N_12102);
nand U13265 (N_13265,N_12160,N_12203);
nand U13266 (N_13266,N_12412,N_12365);
xor U13267 (N_13267,N_12629,N_12312);
nor U13268 (N_13268,N_12231,N_12285);
nand U13269 (N_13269,N_12687,N_12190);
or U13270 (N_13270,N_12266,N_12384);
xnor U13271 (N_13271,N_12729,N_12223);
or U13272 (N_13272,N_12485,N_12232);
or U13273 (N_13273,N_12208,N_12180);
or U13274 (N_13274,N_12006,N_12712);
xnor U13275 (N_13275,N_12542,N_12190);
nand U13276 (N_13276,N_12290,N_12457);
xnor U13277 (N_13277,N_12571,N_12359);
or U13278 (N_13278,N_12613,N_12747);
nor U13279 (N_13279,N_12088,N_12017);
nor U13280 (N_13280,N_12367,N_12620);
xor U13281 (N_13281,N_12548,N_12510);
or U13282 (N_13282,N_12656,N_12542);
xnor U13283 (N_13283,N_12222,N_12270);
nand U13284 (N_13284,N_12306,N_12178);
or U13285 (N_13285,N_12627,N_12384);
and U13286 (N_13286,N_12608,N_12137);
xnor U13287 (N_13287,N_12343,N_12700);
or U13288 (N_13288,N_12624,N_12364);
nand U13289 (N_13289,N_12222,N_12123);
and U13290 (N_13290,N_12536,N_12663);
nand U13291 (N_13291,N_12039,N_12667);
nor U13292 (N_13292,N_12522,N_12345);
nor U13293 (N_13293,N_12687,N_12254);
xnor U13294 (N_13294,N_12096,N_12533);
and U13295 (N_13295,N_12294,N_12326);
and U13296 (N_13296,N_12717,N_12323);
nand U13297 (N_13297,N_12651,N_12550);
nor U13298 (N_13298,N_12135,N_12568);
nand U13299 (N_13299,N_12571,N_12737);
and U13300 (N_13300,N_12074,N_12636);
or U13301 (N_13301,N_12333,N_12673);
or U13302 (N_13302,N_12081,N_12686);
and U13303 (N_13303,N_12223,N_12190);
nor U13304 (N_13304,N_12725,N_12601);
or U13305 (N_13305,N_12545,N_12138);
and U13306 (N_13306,N_12384,N_12005);
nand U13307 (N_13307,N_12579,N_12331);
xor U13308 (N_13308,N_12669,N_12251);
nand U13309 (N_13309,N_12318,N_12330);
and U13310 (N_13310,N_12028,N_12347);
xnor U13311 (N_13311,N_12709,N_12409);
xnor U13312 (N_13312,N_12042,N_12504);
and U13313 (N_13313,N_12639,N_12607);
and U13314 (N_13314,N_12590,N_12681);
nand U13315 (N_13315,N_12189,N_12106);
and U13316 (N_13316,N_12439,N_12362);
nor U13317 (N_13317,N_12424,N_12527);
or U13318 (N_13318,N_12590,N_12512);
nor U13319 (N_13319,N_12686,N_12633);
or U13320 (N_13320,N_12451,N_12109);
xor U13321 (N_13321,N_12049,N_12391);
xnor U13322 (N_13322,N_12292,N_12282);
xor U13323 (N_13323,N_12595,N_12394);
and U13324 (N_13324,N_12479,N_12113);
and U13325 (N_13325,N_12718,N_12419);
xnor U13326 (N_13326,N_12293,N_12206);
xnor U13327 (N_13327,N_12166,N_12178);
or U13328 (N_13328,N_12620,N_12428);
or U13329 (N_13329,N_12567,N_12014);
nor U13330 (N_13330,N_12163,N_12486);
and U13331 (N_13331,N_12160,N_12567);
nor U13332 (N_13332,N_12196,N_12309);
xnor U13333 (N_13333,N_12597,N_12627);
nand U13334 (N_13334,N_12184,N_12466);
xor U13335 (N_13335,N_12097,N_12478);
nand U13336 (N_13336,N_12708,N_12020);
xnor U13337 (N_13337,N_12183,N_12068);
nor U13338 (N_13338,N_12326,N_12045);
nand U13339 (N_13339,N_12557,N_12690);
xnor U13340 (N_13340,N_12734,N_12491);
xor U13341 (N_13341,N_12383,N_12665);
or U13342 (N_13342,N_12367,N_12451);
xor U13343 (N_13343,N_12543,N_12165);
nor U13344 (N_13344,N_12239,N_12627);
and U13345 (N_13345,N_12360,N_12620);
nor U13346 (N_13346,N_12654,N_12363);
xnor U13347 (N_13347,N_12449,N_12440);
nand U13348 (N_13348,N_12111,N_12338);
nor U13349 (N_13349,N_12026,N_12460);
or U13350 (N_13350,N_12316,N_12424);
xnor U13351 (N_13351,N_12489,N_12212);
and U13352 (N_13352,N_12382,N_12020);
nor U13353 (N_13353,N_12309,N_12681);
nand U13354 (N_13354,N_12562,N_12409);
and U13355 (N_13355,N_12409,N_12465);
xnor U13356 (N_13356,N_12288,N_12168);
or U13357 (N_13357,N_12211,N_12347);
nor U13358 (N_13358,N_12729,N_12060);
xor U13359 (N_13359,N_12407,N_12169);
or U13360 (N_13360,N_12513,N_12628);
or U13361 (N_13361,N_12469,N_12121);
nor U13362 (N_13362,N_12158,N_12122);
xnor U13363 (N_13363,N_12173,N_12380);
or U13364 (N_13364,N_12625,N_12274);
xnor U13365 (N_13365,N_12185,N_12426);
xor U13366 (N_13366,N_12148,N_12521);
and U13367 (N_13367,N_12185,N_12399);
nand U13368 (N_13368,N_12357,N_12481);
and U13369 (N_13369,N_12508,N_12312);
nor U13370 (N_13370,N_12654,N_12154);
nand U13371 (N_13371,N_12346,N_12483);
nand U13372 (N_13372,N_12430,N_12484);
or U13373 (N_13373,N_12718,N_12643);
xor U13374 (N_13374,N_12719,N_12654);
xnor U13375 (N_13375,N_12529,N_12132);
and U13376 (N_13376,N_12000,N_12124);
nand U13377 (N_13377,N_12525,N_12005);
xor U13378 (N_13378,N_12695,N_12187);
nor U13379 (N_13379,N_12488,N_12354);
nor U13380 (N_13380,N_12426,N_12468);
or U13381 (N_13381,N_12232,N_12712);
or U13382 (N_13382,N_12402,N_12347);
and U13383 (N_13383,N_12097,N_12388);
xor U13384 (N_13384,N_12413,N_12401);
or U13385 (N_13385,N_12421,N_12303);
nor U13386 (N_13386,N_12039,N_12114);
or U13387 (N_13387,N_12717,N_12289);
or U13388 (N_13388,N_12214,N_12077);
or U13389 (N_13389,N_12180,N_12414);
xor U13390 (N_13390,N_12622,N_12569);
nor U13391 (N_13391,N_12253,N_12481);
and U13392 (N_13392,N_12097,N_12663);
xnor U13393 (N_13393,N_12080,N_12045);
nand U13394 (N_13394,N_12616,N_12164);
and U13395 (N_13395,N_12683,N_12685);
nand U13396 (N_13396,N_12147,N_12418);
and U13397 (N_13397,N_12126,N_12653);
xnor U13398 (N_13398,N_12600,N_12354);
nand U13399 (N_13399,N_12117,N_12508);
xnor U13400 (N_13400,N_12670,N_12148);
xor U13401 (N_13401,N_12257,N_12477);
nor U13402 (N_13402,N_12502,N_12083);
nor U13403 (N_13403,N_12663,N_12570);
xnor U13404 (N_13404,N_12349,N_12646);
or U13405 (N_13405,N_12508,N_12310);
or U13406 (N_13406,N_12474,N_12550);
xnor U13407 (N_13407,N_12161,N_12593);
xnor U13408 (N_13408,N_12102,N_12657);
or U13409 (N_13409,N_12537,N_12108);
and U13410 (N_13410,N_12592,N_12306);
xor U13411 (N_13411,N_12160,N_12686);
and U13412 (N_13412,N_12468,N_12128);
or U13413 (N_13413,N_12640,N_12527);
xnor U13414 (N_13414,N_12506,N_12041);
xnor U13415 (N_13415,N_12395,N_12459);
and U13416 (N_13416,N_12492,N_12602);
or U13417 (N_13417,N_12041,N_12748);
xor U13418 (N_13418,N_12303,N_12131);
or U13419 (N_13419,N_12596,N_12520);
nand U13420 (N_13420,N_12282,N_12387);
and U13421 (N_13421,N_12263,N_12219);
or U13422 (N_13422,N_12174,N_12309);
nor U13423 (N_13423,N_12200,N_12076);
nor U13424 (N_13424,N_12113,N_12527);
or U13425 (N_13425,N_12615,N_12533);
nor U13426 (N_13426,N_12070,N_12469);
or U13427 (N_13427,N_12056,N_12231);
nand U13428 (N_13428,N_12091,N_12303);
nand U13429 (N_13429,N_12708,N_12186);
xnor U13430 (N_13430,N_12637,N_12317);
and U13431 (N_13431,N_12632,N_12212);
nand U13432 (N_13432,N_12353,N_12051);
nand U13433 (N_13433,N_12177,N_12006);
xnor U13434 (N_13434,N_12535,N_12120);
or U13435 (N_13435,N_12572,N_12263);
or U13436 (N_13436,N_12381,N_12104);
xnor U13437 (N_13437,N_12186,N_12380);
xor U13438 (N_13438,N_12080,N_12056);
xor U13439 (N_13439,N_12052,N_12664);
nand U13440 (N_13440,N_12584,N_12030);
xor U13441 (N_13441,N_12479,N_12520);
nand U13442 (N_13442,N_12593,N_12117);
xor U13443 (N_13443,N_12092,N_12144);
nand U13444 (N_13444,N_12102,N_12489);
or U13445 (N_13445,N_12749,N_12271);
xor U13446 (N_13446,N_12651,N_12717);
nand U13447 (N_13447,N_12486,N_12664);
nor U13448 (N_13448,N_12295,N_12270);
xnor U13449 (N_13449,N_12036,N_12657);
or U13450 (N_13450,N_12698,N_12275);
or U13451 (N_13451,N_12562,N_12553);
nand U13452 (N_13452,N_12283,N_12589);
or U13453 (N_13453,N_12682,N_12603);
xor U13454 (N_13454,N_12356,N_12525);
or U13455 (N_13455,N_12403,N_12097);
nor U13456 (N_13456,N_12331,N_12738);
nor U13457 (N_13457,N_12483,N_12038);
nand U13458 (N_13458,N_12418,N_12482);
and U13459 (N_13459,N_12443,N_12432);
nor U13460 (N_13460,N_12159,N_12412);
or U13461 (N_13461,N_12155,N_12275);
xnor U13462 (N_13462,N_12424,N_12274);
xnor U13463 (N_13463,N_12031,N_12084);
nand U13464 (N_13464,N_12277,N_12461);
xor U13465 (N_13465,N_12038,N_12515);
nand U13466 (N_13466,N_12050,N_12480);
or U13467 (N_13467,N_12562,N_12499);
or U13468 (N_13468,N_12733,N_12450);
nor U13469 (N_13469,N_12149,N_12489);
nor U13470 (N_13470,N_12303,N_12361);
nand U13471 (N_13471,N_12608,N_12435);
nor U13472 (N_13472,N_12667,N_12637);
nor U13473 (N_13473,N_12644,N_12030);
or U13474 (N_13474,N_12501,N_12738);
nand U13475 (N_13475,N_12007,N_12309);
xor U13476 (N_13476,N_12733,N_12515);
nand U13477 (N_13477,N_12098,N_12029);
nand U13478 (N_13478,N_12611,N_12299);
and U13479 (N_13479,N_12499,N_12395);
xor U13480 (N_13480,N_12546,N_12715);
nor U13481 (N_13481,N_12439,N_12435);
nor U13482 (N_13482,N_12574,N_12458);
and U13483 (N_13483,N_12082,N_12157);
nor U13484 (N_13484,N_12454,N_12508);
and U13485 (N_13485,N_12589,N_12141);
nand U13486 (N_13486,N_12392,N_12407);
nand U13487 (N_13487,N_12235,N_12530);
nand U13488 (N_13488,N_12460,N_12066);
or U13489 (N_13489,N_12578,N_12407);
nor U13490 (N_13490,N_12180,N_12063);
nand U13491 (N_13491,N_12637,N_12037);
nor U13492 (N_13492,N_12113,N_12012);
nor U13493 (N_13493,N_12737,N_12701);
and U13494 (N_13494,N_12535,N_12079);
and U13495 (N_13495,N_12627,N_12396);
xor U13496 (N_13496,N_12629,N_12619);
xor U13497 (N_13497,N_12046,N_12138);
nand U13498 (N_13498,N_12505,N_12287);
nand U13499 (N_13499,N_12680,N_12726);
and U13500 (N_13500,N_12859,N_13323);
or U13501 (N_13501,N_13066,N_13405);
xor U13502 (N_13502,N_13435,N_13302);
nor U13503 (N_13503,N_13313,N_12899);
nand U13504 (N_13504,N_12876,N_12932);
xnor U13505 (N_13505,N_13062,N_12926);
nand U13506 (N_13506,N_12917,N_12975);
xor U13507 (N_13507,N_12856,N_13085);
or U13508 (N_13508,N_12903,N_12817);
xor U13509 (N_13509,N_12776,N_12794);
xor U13510 (N_13510,N_13478,N_13188);
xor U13511 (N_13511,N_13342,N_12948);
nand U13512 (N_13512,N_12764,N_13238);
and U13513 (N_13513,N_13194,N_13002);
or U13514 (N_13514,N_12778,N_13232);
nand U13515 (N_13515,N_13437,N_13257);
xnor U13516 (N_13516,N_13226,N_13016);
or U13517 (N_13517,N_12964,N_13347);
nand U13518 (N_13518,N_12910,N_13420);
and U13519 (N_13519,N_13137,N_12960);
or U13520 (N_13520,N_13059,N_13281);
xor U13521 (N_13521,N_13297,N_13418);
or U13522 (N_13522,N_13190,N_13045);
or U13523 (N_13523,N_12968,N_12884);
or U13524 (N_13524,N_12814,N_13301);
nor U13525 (N_13525,N_13192,N_12797);
nor U13526 (N_13526,N_13357,N_13409);
nand U13527 (N_13527,N_13412,N_13125);
and U13528 (N_13528,N_12962,N_12923);
nor U13529 (N_13529,N_13097,N_13078);
nand U13530 (N_13530,N_13464,N_13497);
xor U13531 (N_13531,N_12961,N_13090);
nor U13532 (N_13532,N_12862,N_13024);
or U13533 (N_13533,N_13391,N_12750);
or U13534 (N_13534,N_13153,N_13132);
nor U13535 (N_13535,N_13161,N_13368);
xor U13536 (N_13536,N_13056,N_13375);
nand U13537 (N_13537,N_13414,N_13189);
and U13538 (N_13538,N_12878,N_12915);
or U13539 (N_13539,N_13385,N_13130);
nand U13540 (N_13540,N_13493,N_12763);
or U13541 (N_13541,N_13327,N_13254);
nor U13542 (N_13542,N_12938,N_12973);
or U13543 (N_13543,N_13366,N_13203);
xor U13544 (N_13544,N_13363,N_13263);
or U13545 (N_13545,N_12821,N_13422);
nor U13546 (N_13546,N_12805,N_13439);
or U13547 (N_13547,N_12992,N_12970);
and U13548 (N_13548,N_13111,N_12991);
nor U13549 (N_13549,N_12850,N_12993);
nor U13550 (N_13550,N_12790,N_13217);
nand U13551 (N_13551,N_13213,N_13040);
nor U13552 (N_13552,N_13228,N_13417);
or U13553 (N_13553,N_13241,N_12799);
or U13554 (N_13554,N_13429,N_12857);
and U13555 (N_13555,N_12870,N_13080);
xnor U13556 (N_13556,N_13096,N_12848);
nor U13557 (N_13557,N_13032,N_13242);
nand U13558 (N_13558,N_12858,N_13462);
or U13559 (N_13559,N_12809,N_13492);
or U13560 (N_13560,N_13403,N_13039);
nand U13561 (N_13561,N_13088,N_13460);
xnor U13562 (N_13562,N_12807,N_12869);
xor U13563 (N_13563,N_13127,N_13291);
nand U13564 (N_13564,N_13424,N_12902);
or U13565 (N_13565,N_13348,N_13124);
and U13566 (N_13566,N_12936,N_13000);
nor U13567 (N_13567,N_13370,N_13181);
xnor U13568 (N_13568,N_13411,N_13272);
xnor U13569 (N_13569,N_12772,N_13017);
or U13570 (N_13570,N_13459,N_13224);
or U13571 (N_13571,N_13237,N_13463);
and U13572 (N_13572,N_13221,N_12759);
and U13573 (N_13573,N_13148,N_13171);
nor U13574 (N_13574,N_13067,N_13210);
nor U13575 (N_13575,N_13372,N_13048);
nand U13576 (N_13576,N_12997,N_13406);
nand U13577 (N_13577,N_13036,N_13474);
nor U13578 (N_13578,N_13219,N_12958);
nand U13579 (N_13579,N_13072,N_13317);
and U13580 (N_13580,N_13456,N_12996);
nor U13581 (N_13581,N_13469,N_13328);
xnor U13582 (N_13582,N_13374,N_13471);
xnor U13583 (N_13583,N_13186,N_12933);
nor U13584 (N_13584,N_13094,N_12885);
xnor U13585 (N_13585,N_13329,N_12965);
nand U13586 (N_13586,N_13448,N_12985);
nand U13587 (N_13587,N_13477,N_12893);
and U13588 (N_13588,N_13173,N_13305);
and U13589 (N_13589,N_12909,N_13449);
or U13590 (N_13590,N_13271,N_13114);
and U13591 (N_13591,N_12868,N_13174);
nor U13592 (N_13592,N_13035,N_13454);
xnor U13593 (N_13593,N_13008,N_13335);
nor U13594 (N_13594,N_12877,N_12987);
nor U13595 (N_13595,N_12829,N_12911);
nand U13596 (N_13596,N_13319,N_13309);
nor U13597 (N_13597,N_13410,N_13350);
and U13598 (N_13598,N_12808,N_13012);
or U13599 (N_13599,N_12943,N_13250);
nor U13600 (N_13600,N_13499,N_13476);
nor U13601 (N_13601,N_13303,N_13240);
and U13602 (N_13602,N_12976,N_13280);
nor U13603 (N_13603,N_13438,N_13466);
and U13604 (N_13604,N_13491,N_12840);
xor U13605 (N_13605,N_13149,N_12952);
xor U13606 (N_13606,N_12752,N_12888);
nor U13607 (N_13607,N_13276,N_12802);
nand U13608 (N_13608,N_12875,N_13100);
or U13609 (N_13609,N_12828,N_12784);
xnor U13610 (N_13610,N_13294,N_13199);
or U13611 (N_13611,N_13255,N_13083);
and U13612 (N_13612,N_12963,N_13445);
or U13613 (N_13613,N_13296,N_13356);
or U13614 (N_13614,N_12955,N_13101);
xor U13615 (N_13615,N_13468,N_12783);
nor U13616 (N_13616,N_13396,N_13231);
nand U13617 (N_13617,N_12922,N_12937);
or U13618 (N_13618,N_13310,N_13156);
xnor U13619 (N_13619,N_13165,N_13209);
xor U13620 (N_13620,N_13371,N_12891);
xnor U13621 (N_13621,N_13482,N_13444);
or U13622 (N_13622,N_13401,N_13473);
xor U13623 (N_13623,N_13407,N_13277);
and U13624 (N_13624,N_13122,N_12836);
or U13625 (N_13625,N_13316,N_12981);
nand U13626 (N_13626,N_13047,N_13109);
nor U13627 (N_13627,N_13034,N_12780);
and U13628 (N_13628,N_13136,N_12754);
nand U13629 (N_13629,N_13239,N_12777);
xor U13630 (N_13630,N_13485,N_13106);
and U13631 (N_13631,N_12787,N_13431);
xnor U13632 (N_13632,N_12755,N_13398);
or U13633 (N_13633,N_12967,N_12804);
xnor U13634 (N_13634,N_12833,N_13113);
xnor U13635 (N_13635,N_13120,N_12806);
or U13636 (N_13636,N_13184,N_13353);
and U13637 (N_13637,N_13321,N_13457);
and U13638 (N_13638,N_13058,N_12920);
nand U13639 (N_13639,N_13021,N_13273);
nor U13640 (N_13640,N_12873,N_13107);
xnor U13641 (N_13641,N_13311,N_12871);
xor U13642 (N_13642,N_13404,N_13212);
and U13643 (N_13643,N_13290,N_13006);
nand U13644 (N_13644,N_13086,N_12818);
or U13645 (N_13645,N_13245,N_13177);
nand U13646 (N_13646,N_12944,N_13158);
nand U13647 (N_13647,N_12892,N_13200);
nor U13648 (N_13648,N_13247,N_12946);
nor U13649 (N_13649,N_13425,N_13386);
nor U13650 (N_13650,N_12872,N_13265);
nor U13651 (N_13651,N_13227,N_13128);
nand U13652 (N_13652,N_13175,N_12940);
xor U13653 (N_13653,N_13019,N_13266);
nor U13654 (N_13654,N_13160,N_12994);
and U13655 (N_13655,N_12798,N_12914);
nor U13656 (N_13656,N_12988,N_13395);
nand U13657 (N_13657,N_13269,N_13204);
or U13658 (N_13658,N_13044,N_13360);
and U13659 (N_13659,N_13258,N_13014);
xnor U13660 (N_13660,N_12830,N_13001);
nor U13661 (N_13661,N_12846,N_13421);
xor U13662 (N_13662,N_13381,N_12907);
or U13663 (N_13663,N_12852,N_12793);
nor U13664 (N_13664,N_12811,N_12900);
nor U13665 (N_13665,N_13487,N_13455);
and U13666 (N_13666,N_12919,N_13225);
nand U13667 (N_13667,N_12977,N_12820);
or U13668 (N_13668,N_13367,N_13236);
and U13669 (N_13669,N_13494,N_12894);
nand U13670 (N_13670,N_12950,N_12823);
xor U13671 (N_13671,N_13015,N_13157);
nor U13672 (N_13672,N_13139,N_13432);
nor U13673 (N_13673,N_12867,N_13261);
xnor U13674 (N_13674,N_13349,N_13207);
or U13675 (N_13675,N_13077,N_13314);
and U13676 (N_13676,N_13467,N_13134);
xnor U13677 (N_13677,N_13119,N_13223);
nand U13678 (N_13678,N_13193,N_12890);
and U13679 (N_13679,N_12978,N_13208);
xnor U13680 (N_13680,N_13075,N_13073);
xnor U13681 (N_13681,N_13135,N_13322);
nand U13682 (N_13682,N_13434,N_13027);
or U13683 (N_13683,N_13433,N_13144);
nand U13684 (N_13684,N_13098,N_12767);
xnor U13685 (N_13685,N_12782,N_12947);
xor U13686 (N_13686,N_13091,N_13095);
and U13687 (N_13687,N_13442,N_13352);
and U13688 (N_13688,N_13230,N_13140);
nor U13689 (N_13689,N_13343,N_13495);
nand U13690 (N_13690,N_12834,N_13079);
or U13691 (N_13691,N_13218,N_13436);
xor U13692 (N_13692,N_12801,N_13496);
xor U13693 (N_13693,N_13246,N_13292);
xor U13694 (N_13694,N_13214,N_12855);
or U13695 (N_13695,N_13441,N_13481);
or U13696 (N_13696,N_12774,N_12847);
nand U13697 (N_13697,N_13028,N_13064);
xnor U13698 (N_13698,N_13389,N_12785);
xor U13699 (N_13699,N_12971,N_13369);
xnor U13700 (N_13700,N_12974,N_12999);
or U13701 (N_13701,N_12864,N_12990);
nand U13702 (N_13702,N_12824,N_13452);
xnor U13703 (N_13703,N_13426,N_12881);
nand U13704 (N_13704,N_13065,N_12770);
nor U13705 (N_13705,N_12795,N_13390);
nand U13706 (N_13706,N_13050,N_13220);
nand U13707 (N_13707,N_13041,N_13279);
nand U13708 (N_13708,N_12916,N_13318);
or U13709 (N_13709,N_12898,N_12983);
or U13710 (N_13710,N_13117,N_13325);
nor U13711 (N_13711,N_12786,N_13176);
and U13712 (N_13712,N_12773,N_12865);
nor U13713 (N_13713,N_13253,N_12931);
and U13714 (N_13714,N_13112,N_12803);
nand U13715 (N_13715,N_13299,N_13326);
and U13716 (N_13716,N_12913,N_13102);
xnor U13717 (N_13717,N_13376,N_13498);
nand U13718 (N_13718,N_13345,N_12934);
xor U13719 (N_13719,N_13490,N_13206);
xnor U13720 (N_13720,N_12866,N_13118);
nand U13721 (N_13721,N_13105,N_13379);
nor U13722 (N_13722,N_13060,N_13116);
nor U13723 (N_13723,N_13092,N_13388);
and U13724 (N_13724,N_12906,N_13278);
and U13725 (N_13725,N_13408,N_13013);
xor U13726 (N_13726,N_13315,N_12941);
and U13727 (N_13727,N_12905,N_13307);
xor U13728 (N_13728,N_12880,N_12839);
or U13729 (N_13729,N_13289,N_13009);
xor U13730 (N_13730,N_12837,N_12788);
or U13731 (N_13731,N_13197,N_13355);
nor U13732 (N_13732,N_13215,N_12766);
nor U13733 (N_13733,N_13129,N_13488);
nand U13734 (N_13734,N_12854,N_13430);
nand U13735 (N_13735,N_13483,N_13196);
nand U13736 (N_13736,N_13152,N_13249);
or U13737 (N_13737,N_12860,N_13068);
nand U13738 (N_13738,N_13018,N_13071);
xor U13739 (N_13739,N_13010,N_13169);
and U13740 (N_13740,N_13030,N_13151);
nand U13741 (N_13741,N_13270,N_13378);
or U13742 (N_13742,N_12863,N_13423);
and U13743 (N_13743,N_12813,N_13133);
xor U13744 (N_13744,N_13033,N_13115);
nor U13745 (N_13745,N_13089,N_13063);
and U13746 (N_13746,N_13380,N_12969);
nand U13747 (N_13747,N_13282,N_13004);
nor U13748 (N_13748,N_13121,N_13055);
xor U13749 (N_13749,N_13243,N_12982);
nand U13750 (N_13750,N_12825,N_12851);
or U13751 (N_13751,N_12887,N_12816);
or U13752 (N_13752,N_12928,N_12949);
xnor U13753 (N_13753,N_13216,N_12954);
xnor U13754 (N_13754,N_12942,N_13126);
nor U13755 (N_13755,N_13264,N_12796);
xnor U13756 (N_13756,N_13146,N_12826);
nand U13757 (N_13757,N_12912,N_13087);
or U13758 (N_13758,N_13443,N_13359);
or U13759 (N_13759,N_13082,N_13489);
xnor U13760 (N_13760,N_12841,N_13362);
nor U13761 (N_13761,N_13451,N_13447);
or U13762 (N_13762,N_13052,N_13046);
or U13763 (N_13763,N_13402,N_13419);
nand U13764 (N_13764,N_13093,N_13320);
nor U13765 (N_13765,N_13170,N_13005);
and U13766 (N_13766,N_13003,N_13043);
nand U13767 (N_13767,N_13397,N_12889);
or U13768 (N_13768,N_13110,N_13286);
or U13769 (N_13769,N_13049,N_12897);
xnor U13770 (N_13770,N_12768,N_13150);
nor U13771 (N_13771,N_13399,N_13400);
nand U13772 (N_13772,N_12979,N_13167);
nor U13773 (N_13773,N_13069,N_13287);
nor U13774 (N_13774,N_12883,N_13479);
nor U13775 (N_13775,N_12953,N_12959);
or U13776 (N_13776,N_13031,N_13275);
nor U13777 (N_13777,N_12927,N_13344);
nand U13778 (N_13778,N_12822,N_13358);
xor U13779 (N_13779,N_13354,N_13026);
or U13780 (N_13780,N_13336,N_12879);
and U13781 (N_13781,N_13022,N_13029);
and U13782 (N_13782,N_13346,N_13159);
nand U13783 (N_13783,N_12957,N_12838);
xor U13784 (N_13784,N_13099,N_13284);
nand U13785 (N_13785,N_13274,N_13183);
and U13786 (N_13786,N_12800,N_13453);
and U13787 (N_13787,N_13377,N_13020);
and U13788 (N_13788,N_13195,N_13123);
nor U13789 (N_13789,N_13145,N_12843);
and U13790 (N_13790,N_13288,N_13306);
and U13791 (N_13791,N_13251,N_13178);
nand U13792 (N_13792,N_13285,N_13268);
or U13793 (N_13793,N_12901,N_13248);
or U13794 (N_13794,N_13382,N_12951);
nand U13795 (N_13795,N_12886,N_13053);
or U13796 (N_13796,N_12779,N_12835);
nand U13797 (N_13797,N_13138,N_12989);
and U13798 (N_13798,N_12935,N_13339);
nand U13799 (N_13799,N_13222,N_13384);
or U13800 (N_13800,N_13201,N_13179);
or U13801 (N_13801,N_12853,N_13440);
xnor U13802 (N_13802,N_13267,N_12908);
nand U13803 (N_13803,N_13233,N_12792);
nor U13804 (N_13804,N_13332,N_13262);
or U13805 (N_13805,N_13428,N_12819);
nor U13806 (N_13806,N_12918,N_13108);
xor U13807 (N_13807,N_13084,N_12832);
and U13808 (N_13808,N_13042,N_12753);
nand U13809 (N_13809,N_12980,N_13351);
xor U13810 (N_13810,N_12756,N_12831);
or U13811 (N_13811,N_12758,N_12861);
nor U13812 (N_13812,N_12815,N_13415);
nor U13813 (N_13813,N_12956,N_13484);
nor U13814 (N_13814,N_12930,N_12998);
nand U13815 (N_13815,N_13154,N_13365);
or U13816 (N_13816,N_12972,N_13427);
nand U13817 (N_13817,N_13180,N_13076);
and U13818 (N_13818,N_12769,N_12791);
and U13819 (N_13819,N_13187,N_13191);
and U13820 (N_13820,N_13283,N_12896);
xnor U13821 (N_13821,N_13155,N_12849);
or U13822 (N_13822,N_13131,N_13461);
and U13823 (N_13823,N_12812,N_13304);
nand U13824 (N_13824,N_13182,N_13054);
or U13825 (N_13825,N_13475,N_13324);
nor U13826 (N_13826,N_13185,N_13103);
or U13827 (N_13827,N_13162,N_12771);
or U13828 (N_13828,N_12789,N_13260);
nor U13829 (N_13829,N_13338,N_13166);
and U13830 (N_13830,N_13416,N_12904);
nand U13831 (N_13831,N_13331,N_13252);
nand U13832 (N_13832,N_12757,N_12929);
nor U13833 (N_13833,N_12827,N_13143);
xnor U13834 (N_13834,N_13472,N_13164);
nand U13835 (N_13835,N_12751,N_13298);
nand U13836 (N_13836,N_13259,N_13480);
nor U13837 (N_13837,N_12762,N_13142);
xnor U13838 (N_13838,N_13205,N_13458);
xor U13839 (N_13839,N_13011,N_12986);
nor U13840 (N_13840,N_12921,N_13337);
xor U13841 (N_13841,N_13234,N_12924);
nand U13842 (N_13842,N_13023,N_13392);
nand U13843 (N_13843,N_13334,N_12925);
nor U13844 (N_13844,N_13007,N_13373);
nor U13845 (N_13845,N_13037,N_13025);
nor U13846 (N_13846,N_13341,N_13312);
xor U13847 (N_13847,N_13300,N_13330);
nor U13848 (N_13848,N_13486,N_13364);
nand U13849 (N_13849,N_13446,N_13465);
nand U13850 (N_13850,N_13163,N_12761);
xnor U13851 (N_13851,N_13168,N_13383);
or U13852 (N_13852,N_12882,N_13070);
xor U13853 (N_13853,N_12810,N_13061);
or U13854 (N_13854,N_13244,N_13470);
nor U13855 (N_13855,N_12966,N_12842);
nor U13856 (N_13856,N_13229,N_13256);
nand U13857 (N_13857,N_13394,N_13295);
or U13858 (N_13858,N_13141,N_12995);
xor U13859 (N_13859,N_12760,N_12775);
nand U13860 (N_13860,N_13198,N_13393);
nor U13861 (N_13861,N_13172,N_13293);
nand U13862 (N_13862,N_13081,N_12939);
nor U13863 (N_13863,N_12844,N_13057);
or U13864 (N_13864,N_13051,N_12845);
xnor U13865 (N_13865,N_13387,N_13450);
and U13866 (N_13866,N_13308,N_13211);
nor U13867 (N_13867,N_13074,N_12874);
nand U13868 (N_13868,N_12895,N_13202);
and U13869 (N_13869,N_12781,N_13235);
nand U13870 (N_13870,N_12984,N_13038);
xor U13871 (N_13871,N_12765,N_13413);
or U13872 (N_13872,N_13361,N_12945);
and U13873 (N_13873,N_13333,N_13104);
xnor U13874 (N_13874,N_13147,N_13340);
or U13875 (N_13875,N_13329,N_13036);
and U13876 (N_13876,N_13311,N_12784);
or U13877 (N_13877,N_13258,N_13485);
and U13878 (N_13878,N_13464,N_13117);
and U13879 (N_13879,N_13471,N_13137);
xnor U13880 (N_13880,N_13278,N_13298);
nor U13881 (N_13881,N_12849,N_13223);
and U13882 (N_13882,N_13446,N_13039);
nand U13883 (N_13883,N_13228,N_12892);
or U13884 (N_13884,N_13141,N_12850);
and U13885 (N_13885,N_12821,N_13456);
or U13886 (N_13886,N_12872,N_12762);
or U13887 (N_13887,N_13314,N_13405);
nor U13888 (N_13888,N_12938,N_12949);
nand U13889 (N_13889,N_13399,N_13389);
or U13890 (N_13890,N_13301,N_12958);
nor U13891 (N_13891,N_12858,N_13372);
nor U13892 (N_13892,N_12864,N_13429);
xor U13893 (N_13893,N_13396,N_13426);
nor U13894 (N_13894,N_13082,N_13208);
nor U13895 (N_13895,N_13054,N_13074);
nor U13896 (N_13896,N_13264,N_13227);
and U13897 (N_13897,N_13400,N_13160);
nand U13898 (N_13898,N_13472,N_13414);
or U13899 (N_13899,N_13407,N_13225);
xnor U13900 (N_13900,N_13145,N_13470);
xnor U13901 (N_13901,N_12824,N_13432);
xnor U13902 (N_13902,N_13377,N_13188);
and U13903 (N_13903,N_13281,N_12824);
nand U13904 (N_13904,N_13408,N_12785);
xnor U13905 (N_13905,N_13044,N_13217);
or U13906 (N_13906,N_12892,N_13180);
xor U13907 (N_13907,N_13092,N_13031);
xnor U13908 (N_13908,N_13094,N_12838);
or U13909 (N_13909,N_13327,N_13126);
nand U13910 (N_13910,N_13346,N_12879);
nor U13911 (N_13911,N_12908,N_12966);
nor U13912 (N_13912,N_13186,N_13149);
nand U13913 (N_13913,N_13432,N_13189);
nor U13914 (N_13914,N_12831,N_13462);
or U13915 (N_13915,N_13203,N_13044);
and U13916 (N_13916,N_13468,N_13382);
and U13917 (N_13917,N_13064,N_13462);
and U13918 (N_13918,N_13446,N_13174);
nand U13919 (N_13919,N_12797,N_13376);
xnor U13920 (N_13920,N_13176,N_13396);
or U13921 (N_13921,N_13310,N_12806);
and U13922 (N_13922,N_13495,N_13243);
and U13923 (N_13923,N_13190,N_13256);
nand U13924 (N_13924,N_13456,N_13011);
xor U13925 (N_13925,N_12960,N_13233);
nor U13926 (N_13926,N_13246,N_13140);
xor U13927 (N_13927,N_13357,N_12771);
xnor U13928 (N_13928,N_12968,N_13192);
xor U13929 (N_13929,N_13099,N_12873);
and U13930 (N_13930,N_12790,N_12751);
or U13931 (N_13931,N_12972,N_13157);
and U13932 (N_13932,N_13450,N_13051);
and U13933 (N_13933,N_13455,N_13387);
or U13934 (N_13934,N_13071,N_12788);
or U13935 (N_13935,N_12772,N_13497);
xnor U13936 (N_13936,N_13347,N_12948);
nand U13937 (N_13937,N_13252,N_13251);
xor U13938 (N_13938,N_12961,N_13183);
xnor U13939 (N_13939,N_12836,N_13053);
or U13940 (N_13940,N_13277,N_13225);
or U13941 (N_13941,N_12974,N_12841);
or U13942 (N_13942,N_13385,N_13330);
or U13943 (N_13943,N_13300,N_12870);
nor U13944 (N_13944,N_12952,N_13446);
xnor U13945 (N_13945,N_13112,N_13093);
nand U13946 (N_13946,N_13310,N_13394);
and U13947 (N_13947,N_13007,N_13417);
xnor U13948 (N_13948,N_12789,N_12772);
or U13949 (N_13949,N_13386,N_12907);
nand U13950 (N_13950,N_13056,N_13331);
xor U13951 (N_13951,N_12899,N_12820);
and U13952 (N_13952,N_13431,N_13146);
or U13953 (N_13953,N_13344,N_12757);
nand U13954 (N_13954,N_13198,N_13226);
nor U13955 (N_13955,N_12836,N_12847);
xnor U13956 (N_13956,N_13188,N_12766);
or U13957 (N_13957,N_13225,N_13029);
xnor U13958 (N_13958,N_13295,N_13166);
and U13959 (N_13959,N_13189,N_13224);
xnor U13960 (N_13960,N_12842,N_12760);
xnor U13961 (N_13961,N_12751,N_13081);
nor U13962 (N_13962,N_13061,N_13215);
nor U13963 (N_13963,N_13001,N_13200);
and U13964 (N_13964,N_13234,N_13132);
and U13965 (N_13965,N_12891,N_13422);
or U13966 (N_13966,N_12996,N_13485);
or U13967 (N_13967,N_12876,N_12774);
and U13968 (N_13968,N_13236,N_13459);
and U13969 (N_13969,N_13099,N_12753);
nand U13970 (N_13970,N_12826,N_12850);
xnor U13971 (N_13971,N_12899,N_13475);
or U13972 (N_13972,N_13454,N_13011);
nand U13973 (N_13973,N_13146,N_13490);
nand U13974 (N_13974,N_13416,N_13125);
nand U13975 (N_13975,N_13349,N_13020);
nand U13976 (N_13976,N_13461,N_12862);
or U13977 (N_13977,N_13494,N_13389);
and U13978 (N_13978,N_12859,N_12864);
xor U13979 (N_13979,N_13026,N_12843);
and U13980 (N_13980,N_13412,N_13045);
and U13981 (N_13981,N_12860,N_12782);
and U13982 (N_13982,N_13018,N_13254);
nand U13983 (N_13983,N_13084,N_12914);
or U13984 (N_13984,N_13177,N_12790);
or U13985 (N_13985,N_13022,N_13360);
xor U13986 (N_13986,N_13195,N_12896);
nand U13987 (N_13987,N_13226,N_12977);
or U13988 (N_13988,N_13019,N_12948);
nor U13989 (N_13989,N_13026,N_13478);
nand U13990 (N_13990,N_12882,N_12913);
or U13991 (N_13991,N_13285,N_12777);
xor U13992 (N_13992,N_13462,N_13207);
xnor U13993 (N_13993,N_13057,N_13119);
xnor U13994 (N_13994,N_13204,N_12933);
or U13995 (N_13995,N_13034,N_12805);
or U13996 (N_13996,N_13252,N_13491);
or U13997 (N_13997,N_13086,N_13124);
nand U13998 (N_13998,N_12994,N_13017);
nand U13999 (N_13999,N_13384,N_13441);
or U14000 (N_14000,N_13037,N_12966);
and U14001 (N_14001,N_13038,N_12939);
or U14002 (N_14002,N_13423,N_13272);
or U14003 (N_14003,N_13271,N_12916);
nand U14004 (N_14004,N_13061,N_12798);
and U14005 (N_14005,N_13207,N_13389);
and U14006 (N_14006,N_13096,N_13281);
nor U14007 (N_14007,N_12752,N_12970);
or U14008 (N_14008,N_13114,N_13137);
nor U14009 (N_14009,N_13415,N_13017);
xnor U14010 (N_14010,N_13330,N_13254);
and U14011 (N_14011,N_13203,N_13131);
and U14012 (N_14012,N_13034,N_13025);
nand U14013 (N_14013,N_13491,N_12804);
nand U14014 (N_14014,N_12765,N_13441);
xnor U14015 (N_14015,N_13063,N_13342);
nand U14016 (N_14016,N_13055,N_12869);
and U14017 (N_14017,N_13387,N_13268);
nand U14018 (N_14018,N_13205,N_12989);
or U14019 (N_14019,N_13095,N_12818);
nand U14020 (N_14020,N_13359,N_13448);
nor U14021 (N_14021,N_12861,N_13334);
xnor U14022 (N_14022,N_13215,N_13031);
or U14023 (N_14023,N_13267,N_12937);
or U14024 (N_14024,N_12922,N_13235);
xor U14025 (N_14025,N_13027,N_12842);
nor U14026 (N_14026,N_13285,N_13468);
and U14027 (N_14027,N_13451,N_13370);
and U14028 (N_14028,N_13175,N_13090);
xnor U14029 (N_14029,N_13135,N_13334);
or U14030 (N_14030,N_12821,N_12956);
nor U14031 (N_14031,N_13274,N_13159);
nor U14032 (N_14032,N_12766,N_12962);
nand U14033 (N_14033,N_13409,N_12935);
and U14034 (N_14034,N_13238,N_13074);
or U14035 (N_14035,N_12896,N_13400);
and U14036 (N_14036,N_13207,N_13338);
or U14037 (N_14037,N_13270,N_13340);
nand U14038 (N_14038,N_13185,N_12990);
nor U14039 (N_14039,N_13266,N_13037);
and U14040 (N_14040,N_13453,N_13434);
or U14041 (N_14041,N_13340,N_13087);
xor U14042 (N_14042,N_13136,N_13465);
xnor U14043 (N_14043,N_13010,N_13287);
xor U14044 (N_14044,N_12855,N_13065);
or U14045 (N_14045,N_13002,N_12907);
and U14046 (N_14046,N_13493,N_13226);
nand U14047 (N_14047,N_12842,N_12938);
and U14048 (N_14048,N_12777,N_13462);
or U14049 (N_14049,N_13342,N_13414);
xor U14050 (N_14050,N_13136,N_13051);
nand U14051 (N_14051,N_13377,N_13457);
nand U14052 (N_14052,N_13197,N_13473);
nand U14053 (N_14053,N_13409,N_13375);
and U14054 (N_14054,N_12926,N_12809);
and U14055 (N_14055,N_13415,N_13343);
or U14056 (N_14056,N_13448,N_13250);
nand U14057 (N_14057,N_12815,N_12832);
and U14058 (N_14058,N_12920,N_13075);
nor U14059 (N_14059,N_12773,N_13101);
xnor U14060 (N_14060,N_13261,N_12938);
nand U14061 (N_14061,N_12853,N_13414);
and U14062 (N_14062,N_13428,N_13454);
and U14063 (N_14063,N_13439,N_12812);
nor U14064 (N_14064,N_13016,N_13038);
nor U14065 (N_14065,N_13432,N_13313);
nand U14066 (N_14066,N_12980,N_12795);
nand U14067 (N_14067,N_13242,N_13117);
and U14068 (N_14068,N_13220,N_13211);
nor U14069 (N_14069,N_12987,N_12835);
and U14070 (N_14070,N_13284,N_12995);
and U14071 (N_14071,N_13463,N_12895);
or U14072 (N_14072,N_13185,N_13428);
and U14073 (N_14073,N_13408,N_13311);
nand U14074 (N_14074,N_13466,N_13197);
xor U14075 (N_14075,N_13473,N_12825);
and U14076 (N_14076,N_13171,N_13495);
and U14077 (N_14077,N_13285,N_13391);
nor U14078 (N_14078,N_13312,N_13118);
xor U14079 (N_14079,N_12806,N_12850);
nor U14080 (N_14080,N_13131,N_13053);
xnor U14081 (N_14081,N_12973,N_13382);
nor U14082 (N_14082,N_13123,N_13482);
nor U14083 (N_14083,N_13093,N_13122);
nand U14084 (N_14084,N_13215,N_12911);
and U14085 (N_14085,N_13051,N_12808);
nor U14086 (N_14086,N_13323,N_13139);
nand U14087 (N_14087,N_12915,N_13422);
or U14088 (N_14088,N_12939,N_13089);
and U14089 (N_14089,N_13165,N_13241);
or U14090 (N_14090,N_13359,N_13223);
or U14091 (N_14091,N_12797,N_13371);
nand U14092 (N_14092,N_12926,N_12838);
nand U14093 (N_14093,N_13089,N_13339);
or U14094 (N_14094,N_12831,N_13330);
nand U14095 (N_14095,N_12939,N_12993);
and U14096 (N_14096,N_13383,N_13313);
or U14097 (N_14097,N_13093,N_13047);
xor U14098 (N_14098,N_13020,N_13338);
and U14099 (N_14099,N_13040,N_12953);
xnor U14100 (N_14100,N_13340,N_13390);
xor U14101 (N_14101,N_12820,N_13102);
nand U14102 (N_14102,N_13304,N_12833);
and U14103 (N_14103,N_12852,N_13348);
nand U14104 (N_14104,N_12907,N_13471);
xor U14105 (N_14105,N_13367,N_12886);
and U14106 (N_14106,N_12885,N_13374);
nand U14107 (N_14107,N_12919,N_12851);
xor U14108 (N_14108,N_12926,N_12853);
and U14109 (N_14109,N_12989,N_13481);
nor U14110 (N_14110,N_12814,N_13174);
nor U14111 (N_14111,N_12762,N_12966);
and U14112 (N_14112,N_12894,N_12999);
or U14113 (N_14113,N_12860,N_13291);
or U14114 (N_14114,N_13246,N_12887);
nor U14115 (N_14115,N_12797,N_13055);
nand U14116 (N_14116,N_13294,N_13137);
and U14117 (N_14117,N_13184,N_13201);
xnor U14118 (N_14118,N_13285,N_13371);
nor U14119 (N_14119,N_12991,N_12973);
nor U14120 (N_14120,N_13178,N_13321);
or U14121 (N_14121,N_12780,N_13301);
xnor U14122 (N_14122,N_13007,N_13049);
nor U14123 (N_14123,N_13487,N_13033);
or U14124 (N_14124,N_13174,N_13187);
or U14125 (N_14125,N_13081,N_13466);
and U14126 (N_14126,N_13212,N_12976);
nand U14127 (N_14127,N_13180,N_13397);
nor U14128 (N_14128,N_12824,N_12891);
nand U14129 (N_14129,N_12761,N_13305);
and U14130 (N_14130,N_13092,N_12861);
and U14131 (N_14131,N_13105,N_13146);
nor U14132 (N_14132,N_13224,N_13398);
nor U14133 (N_14133,N_12830,N_12923);
or U14134 (N_14134,N_12862,N_12757);
nor U14135 (N_14135,N_13206,N_13014);
nand U14136 (N_14136,N_12967,N_12884);
xnor U14137 (N_14137,N_13355,N_12807);
nand U14138 (N_14138,N_13293,N_13198);
and U14139 (N_14139,N_13132,N_13272);
nand U14140 (N_14140,N_12916,N_12921);
nor U14141 (N_14141,N_13032,N_13093);
nand U14142 (N_14142,N_13477,N_13495);
nor U14143 (N_14143,N_13025,N_12872);
and U14144 (N_14144,N_13389,N_13331);
xnor U14145 (N_14145,N_13271,N_12905);
and U14146 (N_14146,N_13429,N_13497);
and U14147 (N_14147,N_13340,N_13305);
nand U14148 (N_14148,N_13259,N_13088);
or U14149 (N_14149,N_13276,N_12948);
or U14150 (N_14150,N_12831,N_13312);
or U14151 (N_14151,N_13063,N_13008);
xor U14152 (N_14152,N_13040,N_13319);
and U14153 (N_14153,N_13362,N_13314);
xor U14154 (N_14154,N_12869,N_13344);
nand U14155 (N_14155,N_13373,N_12989);
xnor U14156 (N_14156,N_13359,N_13464);
nand U14157 (N_14157,N_12770,N_13132);
nor U14158 (N_14158,N_12777,N_13066);
and U14159 (N_14159,N_12815,N_13442);
or U14160 (N_14160,N_12767,N_13270);
nor U14161 (N_14161,N_13384,N_13168);
and U14162 (N_14162,N_13374,N_13263);
nor U14163 (N_14163,N_13127,N_12887);
nand U14164 (N_14164,N_12815,N_13438);
nand U14165 (N_14165,N_12851,N_13305);
nand U14166 (N_14166,N_12995,N_13070);
nand U14167 (N_14167,N_13304,N_13241);
nand U14168 (N_14168,N_13156,N_13317);
xnor U14169 (N_14169,N_13180,N_12845);
nor U14170 (N_14170,N_13417,N_12995);
and U14171 (N_14171,N_13496,N_13479);
nand U14172 (N_14172,N_13139,N_13083);
nand U14173 (N_14173,N_13443,N_12851);
xnor U14174 (N_14174,N_13372,N_13030);
nand U14175 (N_14175,N_13328,N_13198);
nor U14176 (N_14176,N_12953,N_12849);
nor U14177 (N_14177,N_12924,N_12770);
or U14178 (N_14178,N_13377,N_13140);
or U14179 (N_14179,N_13228,N_12781);
nand U14180 (N_14180,N_12851,N_12818);
or U14181 (N_14181,N_13361,N_13075);
nand U14182 (N_14182,N_13084,N_12993);
nor U14183 (N_14183,N_13109,N_12978);
xor U14184 (N_14184,N_12796,N_13218);
nand U14185 (N_14185,N_12785,N_13273);
and U14186 (N_14186,N_13380,N_13045);
nand U14187 (N_14187,N_13396,N_12758);
or U14188 (N_14188,N_13143,N_12801);
xnor U14189 (N_14189,N_12988,N_13282);
xor U14190 (N_14190,N_12898,N_13456);
and U14191 (N_14191,N_12942,N_13178);
nand U14192 (N_14192,N_12904,N_13437);
and U14193 (N_14193,N_12989,N_12974);
nor U14194 (N_14194,N_13271,N_12884);
xor U14195 (N_14195,N_13134,N_13334);
nor U14196 (N_14196,N_12866,N_13021);
and U14197 (N_14197,N_13489,N_13268);
nor U14198 (N_14198,N_13240,N_13181);
nand U14199 (N_14199,N_13149,N_13253);
and U14200 (N_14200,N_12923,N_12841);
nand U14201 (N_14201,N_12822,N_13261);
and U14202 (N_14202,N_12900,N_12772);
nand U14203 (N_14203,N_13351,N_13465);
xnor U14204 (N_14204,N_13170,N_13189);
nor U14205 (N_14205,N_13280,N_12960);
and U14206 (N_14206,N_13141,N_12811);
nand U14207 (N_14207,N_13098,N_13090);
nor U14208 (N_14208,N_13297,N_13272);
and U14209 (N_14209,N_13261,N_12811);
or U14210 (N_14210,N_13316,N_12761);
and U14211 (N_14211,N_13321,N_13381);
nand U14212 (N_14212,N_12921,N_13008);
or U14213 (N_14213,N_13256,N_13174);
xnor U14214 (N_14214,N_13472,N_12875);
and U14215 (N_14215,N_13437,N_13276);
and U14216 (N_14216,N_13188,N_12927);
and U14217 (N_14217,N_13087,N_12807);
and U14218 (N_14218,N_12889,N_13006);
nor U14219 (N_14219,N_13421,N_13378);
nor U14220 (N_14220,N_13074,N_13313);
nor U14221 (N_14221,N_13290,N_12944);
or U14222 (N_14222,N_13151,N_12946);
or U14223 (N_14223,N_13051,N_13367);
or U14224 (N_14224,N_13462,N_13194);
xor U14225 (N_14225,N_12962,N_13021);
nand U14226 (N_14226,N_13013,N_12917);
nor U14227 (N_14227,N_13048,N_13152);
and U14228 (N_14228,N_13376,N_13035);
nor U14229 (N_14229,N_13322,N_13228);
and U14230 (N_14230,N_13309,N_13355);
xor U14231 (N_14231,N_13004,N_13471);
or U14232 (N_14232,N_13069,N_12955);
and U14233 (N_14233,N_13225,N_13222);
or U14234 (N_14234,N_13230,N_12778);
or U14235 (N_14235,N_13445,N_12870);
nor U14236 (N_14236,N_12759,N_12926);
nor U14237 (N_14237,N_13488,N_13296);
nand U14238 (N_14238,N_13224,N_13150);
nor U14239 (N_14239,N_13025,N_13084);
or U14240 (N_14240,N_12961,N_12776);
or U14241 (N_14241,N_13284,N_13363);
or U14242 (N_14242,N_13108,N_13031);
nor U14243 (N_14243,N_13226,N_12756);
xnor U14244 (N_14244,N_13499,N_13069);
xnor U14245 (N_14245,N_13370,N_13315);
or U14246 (N_14246,N_13038,N_12886);
xor U14247 (N_14247,N_13369,N_13402);
or U14248 (N_14248,N_13089,N_13490);
xnor U14249 (N_14249,N_13086,N_13301);
xnor U14250 (N_14250,N_14161,N_14195);
and U14251 (N_14251,N_14077,N_13698);
or U14252 (N_14252,N_13574,N_14061);
nor U14253 (N_14253,N_13804,N_13676);
nor U14254 (N_14254,N_13796,N_13713);
nand U14255 (N_14255,N_13868,N_13779);
nand U14256 (N_14256,N_13542,N_13520);
or U14257 (N_14257,N_14145,N_13949);
or U14258 (N_14258,N_14014,N_13716);
nor U14259 (N_14259,N_13580,N_13819);
and U14260 (N_14260,N_13603,N_13971);
or U14261 (N_14261,N_13553,N_14187);
nand U14262 (N_14262,N_13906,N_13691);
nand U14263 (N_14263,N_14078,N_13701);
nor U14264 (N_14264,N_13623,N_14049);
nor U14265 (N_14265,N_14059,N_14073);
nor U14266 (N_14266,N_14227,N_13829);
and U14267 (N_14267,N_14041,N_13812);
nor U14268 (N_14268,N_13889,N_14178);
nand U14269 (N_14269,N_13552,N_13528);
nand U14270 (N_14270,N_13880,N_13831);
xor U14271 (N_14271,N_14221,N_13877);
nand U14272 (N_14272,N_13609,N_14232);
nor U14273 (N_14273,N_13665,N_13964);
and U14274 (N_14274,N_13758,N_14039);
xor U14275 (N_14275,N_13989,N_13718);
and U14276 (N_14276,N_14148,N_13882);
and U14277 (N_14277,N_13720,N_13611);
or U14278 (N_14278,N_13892,N_13821);
or U14279 (N_14279,N_13673,N_14057);
xnor U14280 (N_14280,N_14019,N_13905);
or U14281 (N_14281,N_13699,N_14036);
and U14282 (N_14282,N_14204,N_13715);
nor U14283 (N_14283,N_13567,N_14213);
or U14284 (N_14284,N_14099,N_13746);
nand U14285 (N_14285,N_14017,N_13709);
and U14286 (N_14286,N_14088,N_13823);
nand U14287 (N_14287,N_14132,N_14231);
or U14288 (N_14288,N_13937,N_13845);
xnor U14289 (N_14289,N_13932,N_14018);
xnor U14290 (N_14290,N_13785,N_13980);
nand U14291 (N_14291,N_13769,N_14079);
nor U14292 (N_14292,N_13621,N_14023);
nand U14293 (N_14293,N_13592,N_14081);
xnor U14294 (N_14294,N_13772,N_13667);
nand U14295 (N_14295,N_13873,N_13522);
and U14296 (N_14296,N_14159,N_13984);
nand U14297 (N_14297,N_13652,N_13942);
or U14298 (N_14298,N_13576,N_13900);
nand U14299 (N_14299,N_13885,N_14228);
or U14300 (N_14300,N_13757,N_14005);
xor U14301 (N_14301,N_13751,N_14022);
or U14302 (N_14302,N_14054,N_13695);
and U14303 (N_14303,N_13559,N_14163);
xor U14304 (N_14304,N_13705,N_13585);
xor U14305 (N_14305,N_13654,N_14175);
nand U14306 (N_14306,N_13678,N_13822);
or U14307 (N_14307,N_13756,N_14119);
xor U14308 (N_14308,N_14138,N_13643);
or U14309 (N_14309,N_13793,N_13935);
nand U14310 (N_14310,N_14208,N_14025);
nand U14311 (N_14311,N_14129,N_13943);
nor U14312 (N_14312,N_13683,N_13896);
nand U14313 (N_14313,N_14225,N_13597);
nor U14314 (N_14314,N_13607,N_13836);
xnor U14315 (N_14315,N_13930,N_13803);
nor U14316 (N_14316,N_13614,N_14033);
or U14317 (N_14317,N_14043,N_13696);
or U14318 (N_14318,N_13870,N_13961);
nor U14319 (N_14319,N_13968,N_13536);
nor U14320 (N_14320,N_13690,N_14080);
xnor U14321 (N_14321,N_13689,N_14071);
and U14322 (N_14322,N_13972,N_13507);
xnor U14323 (N_14323,N_13693,N_13620);
nand U14324 (N_14324,N_14108,N_13801);
and U14325 (N_14325,N_14157,N_13841);
nor U14326 (N_14326,N_14246,N_13837);
nor U14327 (N_14327,N_13915,N_13884);
nand U14328 (N_14328,N_13658,N_14144);
nand U14329 (N_14329,N_14124,N_13901);
or U14330 (N_14330,N_14001,N_13728);
nor U14331 (N_14331,N_13598,N_13749);
nor U14332 (N_14332,N_14141,N_14242);
or U14333 (N_14333,N_13876,N_13887);
xor U14334 (N_14334,N_14131,N_13869);
or U14335 (N_14335,N_14142,N_14083);
nor U14336 (N_14336,N_14021,N_14115);
xor U14337 (N_14337,N_13765,N_13920);
or U14338 (N_14338,N_14193,N_13578);
xor U14339 (N_14339,N_13988,N_14046);
nor U14340 (N_14340,N_13797,N_14037);
xor U14341 (N_14341,N_13685,N_13736);
or U14342 (N_14342,N_13927,N_13587);
nand U14343 (N_14343,N_13768,N_13719);
or U14344 (N_14344,N_14034,N_13677);
or U14345 (N_14345,N_13537,N_13790);
and U14346 (N_14346,N_13862,N_13526);
nor U14347 (N_14347,N_14137,N_13517);
xor U14348 (N_14348,N_14150,N_13997);
and U14349 (N_14349,N_13610,N_13558);
nor U14350 (N_14350,N_14009,N_13941);
nor U14351 (N_14351,N_13794,N_14184);
and U14352 (N_14352,N_14235,N_13962);
nor U14353 (N_14353,N_14245,N_13771);
xnor U14354 (N_14354,N_13764,N_14075);
nor U14355 (N_14355,N_13687,N_13702);
nand U14356 (N_14356,N_13748,N_13846);
and U14357 (N_14357,N_13516,N_13546);
or U14358 (N_14358,N_14210,N_14114);
xnor U14359 (N_14359,N_13508,N_13588);
xnor U14360 (N_14360,N_13886,N_13987);
nor U14361 (N_14361,N_13992,N_14062);
xnor U14362 (N_14362,N_13903,N_14024);
xor U14363 (N_14363,N_13878,N_13518);
xor U14364 (N_14364,N_14010,N_13531);
xor U14365 (N_14365,N_13525,N_14120);
and U14366 (N_14366,N_13619,N_13714);
or U14367 (N_14367,N_14020,N_13726);
and U14368 (N_14368,N_14205,N_13734);
nor U14369 (N_14369,N_14238,N_14133);
nand U14370 (N_14370,N_14042,N_14147);
nand U14371 (N_14371,N_14047,N_13505);
or U14372 (N_14372,N_14060,N_13830);
and U14373 (N_14373,N_13660,N_13636);
nand U14374 (N_14374,N_13991,N_14200);
or U14375 (N_14375,N_13629,N_13510);
nor U14376 (N_14376,N_13778,N_14089);
nand U14377 (N_14377,N_14202,N_13521);
xor U14378 (N_14378,N_13929,N_13659);
or U14379 (N_14379,N_13783,N_13564);
nand U14380 (N_14380,N_14165,N_14113);
or U14381 (N_14381,N_13630,N_13951);
or U14382 (N_14382,N_14031,N_13653);
xor U14383 (N_14383,N_14052,N_13979);
and U14384 (N_14384,N_13973,N_13589);
or U14385 (N_14385,N_14151,N_13849);
nor U14386 (N_14386,N_13923,N_14248);
and U14387 (N_14387,N_14215,N_14241);
xnor U14388 (N_14388,N_13515,N_14004);
nor U14389 (N_14389,N_13504,N_14162);
and U14390 (N_14390,N_13586,N_13600);
nor U14391 (N_14391,N_14007,N_14082);
nor U14392 (N_14392,N_13641,N_13635);
xor U14393 (N_14393,N_13717,N_13866);
nand U14394 (N_14394,N_13934,N_14068);
or U14395 (N_14395,N_13501,N_13550);
xor U14396 (N_14396,N_13514,N_14094);
nor U14397 (N_14397,N_14100,N_13787);
or U14398 (N_14398,N_13602,N_14140);
or U14399 (N_14399,N_14136,N_13897);
or U14400 (N_14400,N_13606,N_14169);
nand U14401 (N_14401,N_14026,N_14040);
and U14402 (N_14402,N_13612,N_13857);
nor U14403 (N_14403,N_13502,N_13985);
and U14404 (N_14404,N_13664,N_14234);
and U14405 (N_14405,N_13986,N_14000);
and U14406 (N_14406,N_13737,N_14174);
and U14407 (N_14407,N_13651,N_13670);
nor U14408 (N_14408,N_13860,N_13733);
nor U14409 (N_14409,N_13833,N_13631);
and U14410 (N_14410,N_14220,N_13573);
nor U14411 (N_14411,N_14110,N_14168);
or U14412 (N_14412,N_13952,N_13688);
and U14413 (N_14413,N_13560,N_13739);
and U14414 (N_14414,N_13792,N_13632);
nand U14415 (N_14415,N_13593,N_13815);
xor U14416 (N_14416,N_13963,N_13534);
nor U14417 (N_14417,N_13855,N_13890);
nand U14418 (N_14418,N_14015,N_13732);
xor U14419 (N_14419,N_13917,N_14192);
nand U14420 (N_14420,N_14167,N_13704);
nand U14421 (N_14421,N_13911,N_14172);
nor U14422 (N_14422,N_13908,N_14243);
xor U14423 (N_14423,N_13647,N_13864);
nand U14424 (N_14424,N_13512,N_14209);
nor U14425 (N_14425,N_14153,N_14112);
xnor U14426 (N_14426,N_14092,N_13582);
and U14427 (N_14427,N_13983,N_13770);
and U14428 (N_14428,N_13998,N_13538);
or U14429 (N_14429,N_14008,N_13777);
and U14430 (N_14430,N_14097,N_14139);
and U14431 (N_14431,N_13888,N_14029);
and U14432 (N_14432,N_13939,N_13711);
nor U14433 (N_14433,N_14011,N_13978);
and U14434 (N_14434,N_14158,N_13969);
and U14435 (N_14435,N_13825,N_13618);
and U14436 (N_14436,N_13729,N_13708);
nand U14437 (N_14437,N_14109,N_13549);
nand U14438 (N_14438,N_13958,N_13874);
nor U14439 (N_14439,N_14154,N_14096);
and U14440 (N_14440,N_14013,N_13852);
and U14441 (N_14441,N_14053,N_13996);
xor U14442 (N_14442,N_14105,N_14206);
nor U14443 (N_14443,N_14226,N_13858);
nor U14444 (N_14444,N_13506,N_13721);
and U14445 (N_14445,N_13990,N_13782);
nand U14446 (N_14446,N_13966,N_14072);
nor U14447 (N_14447,N_13671,N_14104);
xnor U14448 (N_14448,N_13854,N_13541);
nor U14449 (N_14449,N_13530,N_13839);
nor U14450 (N_14450,N_14098,N_13916);
and U14451 (N_14451,N_13832,N_14126);
or U14452 (N_14452,N_13881,N_14181);
or U14453 (N_14453,N_14035,N_14090);
and U14454 (N_14454,N_13680,N_13633);
nor U14455 (N_14455,N_14212,N_13738);
nor U14456 (N_14456,N_14064,N_13914);
or U14457 (N_14457,N_14125,N_13604);
nor U14458 (N_14458,N_14155,N_13752);
nand U14459 (N_14459,N_13959,N_13820);
nor U14460 (N_14460,N_14170,N_13807);
nor U14461 (N_14461,N_14171,N_13579);
nor U14462 (N_14462,N_14002,N_14050);
nand U14463 (N_14463,N_13981,N_13802);
nor U14464 (N_14464,N_13898,N_13856);
nand U14465 (N_14465,N_14128,N_14122);
or U14466 (N_14466,N_13925,N_13827);
nor U14467 (N_14467,N_14076,N_13760);
or U14468 (N_14468,N_13523,N_14111);
or U14469 (N_14469,N_13575,N_14087);
nor U14470 (N_14470,N_14230,N_13750);
nand U14471 (N_14471,N_14214,N_14030);
xor U14472 (N_14472,N_14045,N_14189);
or U14473 (N_14473,N_13735,N_13791);
or U14474 (N_14474,N_14190,N_13944);
xor U14475 (N_14475,N_13539,N_13977);
and U14476 (N_14476,N_13679,N_14067);
nor U14477 (N_14477,N_14146,N_13657);
nor U14478 (N_14478,N_13909,N_14084);
nor U14479 (N_14479,N_13840,N_13799);
nor U14480 (N_14480,N_14074,N_13809);
xnor U14481 (N_14481,N_14149,N_13544);
and U14482 (N_14482,N_13775,N_13590);
nor U14483 (N_14483,N_13712,N_13563);
xor U14484 (N_14484,N_13556,N_13511);
xor U14485 (N_14485,N_14222,N_13554);
or U14486 (N_14486,N_13875,N_13548);
nor U14487 (N_14487,N_13936,N_13668);
nor U14488 (N_14488,N_13828,N_13755);
and U14489 (N_14489,N_13813,N_14058);
xnor U14490 (N_14490,N_14207,N_14027);
and U14491 (N_14491,N_13814,N_14197);
or U14492 (N_14492,N_13761,N_14123);
nor U14493 (N_14493,N_13583,N_13891);
xnor U14494 (N_14494,N_13707,N_13817);
or U14495 (N_14495,N_13850,N_13919);
xnor U14496 (N_14496,N_13519,N_13859);
and U14497 (N_14497,N_13894,N_13599);
nand U14498 (N_14498,N_13835,N_13976);
nor U14499 (N_14499,N_13570,N_13646);
or U14500 (N_14500,N_14038,N_13524);
nand U14501 (N_14501,N_13644,N_14183);
nand U14502 (N_14502,N_13543,N_14185);
and U14503 (N_14503,N_14065,N_13741);
nand U14504 (N_14504,N_13781,N_13816);
xor U14505 (N_14505,N_13938,N_13767);
nand U14506 (N_14506,N_13591,N_13805);
xor U14507 (N_14507,N_13762,N_13622);
nor U14508 (N_14508,N_13710,N_14006);
nand U14509 (N_14509,N_14135,N_14166);
or U14510 (N_14510,N_13763,N_14176);
nor U14511 (N_14511,N_13669,N_13834);
xor U14512 (N_14512,N_13565,N_14249);
xor U14513 (N_14513,N_13865,N_14244);
and U14514 (N_14514,N_13753,N_13975);
nor U14515 (N_14515,N_13527,N_13773);
nand U14516 (N_14516,N_13686,N_13640);
and U14517 (N_14517,N_13581,N_13617);
xor U14518 (N_14518,N_13861,N_13557);
and U14519 (N_14519,N_13608,N_13532);
nor U14520 (N_14520,N_13744,N_13893);
xor U14521 (N_14521,N_13842,N_13745);
or U14522 (N_14522,N_13824,N_13933);
nand U14523 (N_14523,N_13547,N_13786);
or U14524 (N_14524,N_13743,N_13577);
nor U14525 (N_14525,N_13922,N_14003);
or U14526 (N_14526,N_13871,N_13649);
or U14527 (N_14527,N_14201,N_13533);
nand U14528 (N_14528,N_13626,N_13595);
nor U14529 (N_14529,N_14066,N_13867);
and U14530 (N_14530,N_13918,N_14095);
nand U14531 (N_14531,N_14199,N_14056);
nor U14532 (N_14532,N_14044,N_14032);
xnor U14533 (N_14533,N_13692,N_14203);
and U14534 (N_14534,N_13747,N_13954);
or U14535 (N_14535,N_14180,N_13910);
nor U14536 (N_14536,N_13742,N_13957);
and U14537 (N_14537,N_14102,N_14216);
nor U14538 (N_14538,N_14012,N_13895);
nand U14539 (N_14539,N_13883,N_13648);
and U14540 (N_14540,N_13672,N_13912);
xor U14541 (N_14541,N_13902,N_13926);
and U14542 (N_14542,N_13513,N_13784);
nor U14543 (N_14543,N_13843,N_13808);
and U14544 (N_14544,N_13965,N_13847);
and U14545 (N_14545,N_13555,N_14016);
nor U14546 (N_14546,N_13806,N_13788);
and U14547 (N_14547,N_13800,N_13945);
nand U14548 (N_14548,N_13970,N_14191);
nor U14549 (N_14549,N_14134,N_13562);
nor U14550 (N_14550,N_14164,N_13994);
and U14551 (N_14551,N_14179,N_13924);
nand U14552 (N_14552,N_14116,N_13638);
and U14553 (N_14553,N_13766,N_14229);
nor U14554 (N_14554,N_13624,N_13568);
xnor U14555 (N_14555,N_13650,N_14086);
or U14556 (N_14556,N_14063,N_13995);
nand U14557 (N_14557,N_14177,N_13613);
nor U14558 (N_14558,N_13956,N_13594);
nand U14559 (N_14559,N_14211,N_13662);
and U14560 (N_14560,N_13982,N_14070);
nand U14561 (N_14561,N_13872,N_13950);
nand U14562 (N_14562,N_13627,N_13851);
xor U14563 (N_14563,N_13904,N_13974);
xnor U14564 (N_14564,N_13913,N_13706);
or U14565 (N_14565,N_14224,N_13625);
nor U14566 (N_14566,N_14198,N_13725);
nor U14567 (N_14567,N_14236,N_13811);
nand U14568 (N_14568,N_13703,N_13535);
xnor U14569 (N_14569,N_14152,N_14091);
xor U14570 (N_14570,N_13838,N_13844);
and U14571 (N_14571,N_14118,N_13931);
and U14572 (N_14572,N_14093,N_14055);
xor U14573 (N_14573,N_14121,N_14117);
or U14574 (N_14574,N_14107,N_14069);
and U14575 (N_14575,N_14143,N_13545);
and U14576 (N_14576,N_13616,N_13960);
and U14577 (N_14577,N_14219,N_14196);
nand U14578 (N_14578,N_13947,N_13500);
xnor U14579 (N_14579,N_13666,N_13848);
nand U14580 (N_14580,N_14240,N_13571);
or U14581 (N_14581,N_13639,N_13637);
nor U14582 (N_14582,N_14186,N_14217);
or U14583 (N_14583,N_13697,N_13655);
or U14584 (N_14584,N_14237,N_13674);
nand U14585 (N_14585,N_13645,N_13681);
or U14586 (N_14586,N_13656,N_13700);
nand U14587 (N_14587,N_14223,N_13509);
or U14588 (N_14588,N_13967,N_14160);
nand U14589 (N_14589,N_13584,N_14103);
xor U14590 (N_14590,N_13551,N_13810);
or U14591 (N_14591,N_13675,N_13853);
nor U14592 (N_14592,N_13999,N_13730);
nand U14593 (N_14593,N_13795,N_13899);
nor U14594 (N_14594,N_13928,N_13601);
and U14595 (N_14595,N_14106,N_13798);
xnor U14596 (N_14596,N_13946,N_14239);
xnor U14597 (N_14597,N_13722,N_13754);
xnor U14598 (N_14598,N_14173,N_13642);
or U14599 (N_14599,N_13948,N_13789);
and U14600 (N_14600,N_14028,N_13940);
xnor U14601 (N_14601,N_13818,N_14194);
nand U14602 (N_14602,N_14085,N_13774);
and U14603 (N_14603,N_14188,N_13605);
or U14604 (N_14604,N_13684,N_13907);
nor U14605 (N_14605,N_14130,N_13993);
nor U14606 (N_14606,N_13723,N_14051);
nand U14607 (N_14607,N_13955,N_13780);
or U14608 (N_14608,N_13596,N_13682);
xnor U14609 (N_14609,N_13540,N_14233);
and U14610 (N_14610,N_14048,N_13776);
and U14611 (N_14611,N_13566,N_13628);
or U14612 (N_14612,N_13663,N_13953);
or U14613 (N_14613,N_14156,N_13503);
nand U14614 (N_14614,N_13826,N_13661);
or U14615 (N_14615,N_13572,N_13529);
nor U14616 (N_14616,N_13879,N_13731);
nor U14617 (N_14617,N_13569,N_13561);
and U14618 (N_14618,N_13921,N_14127);
nand U14619 (N_14619,N_13724,N_13759);
or U14620 (N_14620,N_13634,N_13727);
nor U14621 (N_14621,N_13863,N_13740);
and U14622 (N_14622,N_14218,N_14182);
and U14623 (N_14623,N_13615,N_14247);
nor U14624 (N_14624,N_13694,N_14101);
and U14625 (N_14625,N_14064,N_14043);
nor U14626 (N_14626,N_14116,N_13792);
nand U14627 (N_14627,N_13874,N_14155);
nor U14628 (N_14628,N_14084,N_14013);
or U14629 (N_14629,N_14161,N_14065);
and U14630 (N_14630,N_14246,N_13756);
nor U14631 (N_14631,N_13529,N_14210);
and U14632 (N_14632,N_13750,N_13765);
nor U14633 (N_14633,N_13559,N_13951);
nor U14634 (N_14634,N_13506,N_13580);
and U14635 (N_14635,N_13895,N_14153);
nor U14636 (N_14636,N_13751,N_13581);
nor U14637 (N_14637,N_13854,N_13702);
nand U14638 (N_14638,N_13826,N_13823);
nand U14639 (N_14639,N_13788,N_14146);
or U14640 (N_14640,N_13617,N_14074);
nor U14641 (N_14641,N_14104,N_13887);
nor U14642 (N_14642,N_13593,N_13980);
nor U14643 (N_14643,N_14157,N_13503);
or U14644 (N_14644,N_13924,N_14047);
nor U14645 (N_14645,N_13972,N_13710);
and U14646 (N_14646,N_13968,N_14031);
nand U14647 (N_14647,N_14175,N_14225);
nor U14648 (N_14648,N_13528,N_13730);
and U14649 (N_14649,N_13646,N_14078);
xnor U14650 (N_14650,N_13756,N_13573);
xor U14651 (N_14651,N_14181,N_14027);
xor U14652 (N_14652,N_13639,N_13892);
nand U14653 (N_14653,N_14228,N_13608);
nor U14654 (N_14654,N_14000,N_14161);
or U14655 (N_14655,N_13885,N_13964);
and U14656 (N_14656,N_13859,N_13567);
nand U14657 (N_14657,N_13981,N_13951);
and U14658 (N_14658,N_13749,N_13792);
or U14659 (N_14659,N_14124,N_13999);
and U14660 (N_14660,N_14227,N_13751);
nor U14661 (N_14661,N_14218,N_14029);
xor U14662 (N_14662,N_13747,N_13841);
nand U14663 (N_14663,N_13672,N_14091);
and U14664 (N_14664,N_13836,N_13557);
nand U14665 (N_14665,N_13895,N_13633);
or U14666 (N_14666,N_13627,N_14166);
or U14667 (N_14667,N_13897,N_13529);
xor U14668 (N_14668,N_14094,N_13591);
and U14669 (N_14669,N_14219,N_13574);
nand U14670 (N_14670,N_13800,N_13988);
nand U14671 (N_14671,N_13719,N_13838);
and U14672 (N_14672,N_13756,N_13843);
and U14673 (N_14673,N_13617,N_14046);
xor U14674 (N_14674,N_14015,N_13718);
nand U14675 (N_14675,N_13713,N_14106);
nor U14676 (N_14676,N_14220,N_14123);
nand U14677 (N_14677,N_13837,N_13763);
or U14678 (N_14678,N_13949,N_13903);
nor U14679 (N_14679,N_13714,N_13987);
and U14680 (N_14680,N_13747,N_13559);
or U14681 (N_14681,N_13572,N_13979);
or U14682 (N_14682,N_13645,N_13745);
xnor U14683 (N_14683,N_13697,N_13752);
or U14684 (N_14684,N_13904,N_13913);
nor U14685 (N_14685,N_13804,N_13632);
or U14686 (N_14686,N_13786,N_13706);
xnor U14687 (N_14687,N_13881,N_13639);
or U14688 (N_14688,N_13527,N_14175);
xnor U14689 (N_14689,N_13794,N_13997);
nor U14690 (N_14690,N_13615,N_14165);
and U14691 (N_14691,N_14160,N_13559);
xnor U14692 (N_14692,N_14055,N_13857);
nor U14693 (N_14693,N_14236,N_13553);
xor U14694 (N_14694,N_13895,N_13587);
and U14695 (N_14695,N_13964,N_13634);
and U14696 (N_14696,N_13827,N_13545);
xor U14697 (N_14697,N_14087,N_13767);
and U14698 (N_14698,N_13766,N_13725);
nor U14699 (N_14699,N_14126,N_13981);
and U14700 (N_14700,N_13817,N_14208);
or U14701 (N_14701,N_13667,N_14189);
and U14702 (N_14702,N_14071,N_14047);
xnor U14703 (N_14703,N_13535,N_14225);
xor U14704 (N_14704,N_14196,N_13926);
and U14705 (N_14705,N_13920,N_13621);
or U14706 (N_14706,N_14190,N_14174);
nor U14707 (N_14707,N_14146,N_14129);
or U14708 (N_14708,N_13864,N_14087);
or U14709 (N_14709,N_13643,N_13750);
xor U14710 (N_14710,N_13837,N_14203);
nor U14711 (N_14711,N_13952,N_14152);
xor U14712 (N_14712,N_13701,N_13939);
and U14713 (N_14713,N_14065,N_13844);
and U14714 (N_14714,N_13617,N_13921);
nor U14715 (N_14715,N_14027,N_14243);
or U14716 (N_14716,N_14001,N_13810);
or U14717 (N_14717,N_13677,N_13880);
xor U14718 (N_14718,N_14136,N_13594);
nor U14719 (N_14719,N_13885,N_13913);
or U14720 (N_14720,N_13920,N_14096);
or U14721 (N_14721,N_13604,N_13969);
xnor U14722 (N_14722,N_13852,N_14197);
nand U14723 (N_14723,N_13848,N_13975);
xor U14724 (N_14724,N_13640,N_13502);
or U14725 (N_14725,N_13962,N_13767);
xnor U14726 (N_14726,N_13833,N_14072);
nand U14727 (N_14727,N_13507,N_14122);
nand U14728 (N_14728,N_14136,N_13761);
nor U14729 (N_14729,N_14016,N_13786);
or U14730 (N_14730,N_14078,N_13993);
nor U14731 (N_14731,N_13529,N_13599);
nand U14732 (N_14732,N_13729,N_13894);
xnor U14733 (N_14733,N_13980,N_13544);
nand U14734 (N_14734,N_13922,N_14050);
or U14735 (N_14735,N_13674,N_14197);
or U14736 (N_14736,N_14055,N_13954);
nor U14737 (N_14737,N_14019,N_14015);
and U14738 (N_14738,N_13657,N_13865);
nor U14739 (N_14739,N_14102,N_13854);
xnor U14740 (N_14740,N_14023,N_13634);
xnor U14741 (N_14741,N_13561,N_13720);
or U14742 (N_14742,N_14122,N_14112);
nand U14743 (N_14743,N_13531,N_13933);
and U14744 (N_14744,N_13711,N_13855);
and U14745 (N_14745,N_13503,N_13905);
nor U14746 (N_14746,N_14115,N_13744);
and U14747 (N_14747,N_13599,N_14035);
nand U14748 (N_14748,N_13566,N_13661);
or U14749 (N_14749,N_13951,N_14074);
nor U14750 (N_14750,N_13519,N_14067);
nand U14751 (N_14751,N_14032,N_14134);
xnor U14752 (N_14752,N_14136,N_13871);
nand U14753 (N_14753,N_13918,N_13569);
and U14754 (N_14754,N_13925,N_13713);
and U14755 (N_14755,N_14247,N_14039);
xnor U14756 (N_14756,N_14061,N_14176);
xor U14757 (N_14757,N_14152,N_13679);
or U14758 (N_14758,N_14000,N_13915);
and U14759 (N_14759,N_13931,N_13878);
xnor U14760 (N_14760,N_13881,N_13633);
and U14761 (N_14761,N_13674,N_13587);
nor U14762 (N_14762,N_14194,N_14035);
nor U14763 (N_14763,N_13593,N_13882);
nor U14764 (N_14764,N_14037,N_13953);
or U14765 (N_14765,N_14126,N_13928);
xnor U14766 (N_14766,N_14247,N_13694);
nor U14767 (N_14767,N_13795,N_13501);
or U14768 (N_14768,N_13542,N_13530);
nand U14769 (N_14769,N_13855,N_13732);
nand U14770 (N_14770,N_13503,N_13666);
nor U14771 (N_14771,N_14064,N_13784);
and U14772 (N_14772,N_13783,N_13602);
nor U14773 (N_14773,N_14094,N_13773);
and U14774 (N_14774,N_13766,N_14107);
xor U14775 (N_14775,N_14097,N_13851);
nand U14776 (N_14776,N_13726,N_13761);
nor U14777 (N_14777,N_13646,N_13606);
and U14778 (N_14778,N_13745,N_13589);
nor U14779 (N_14779,N_13668,N_13860);
or U14780 (N_14780,N_13714,N_13997);
nand U14781 (N_14781,N_13581,N_14009);
and U14782 (N_14782,N_14171,N_13742);
and U14783 (N_14783,N_13876,N_14201);
nor U14784 (N_14784,N_13691,N_13782);
or U14785 (N_14785,N_13672,N_14171);
or U14786 (N_14786,N_14139,N_13781);
or U14787 (N_14787,N_13801,N_14013);
or U14788 (N_14788,N_13804,N_13641);
xor U14789 (N_14789,N_13639,N_13506);
nand U14790 (N_14790,N_13782,N_14232);
or U14791 (N_14791,N_14044,N_13641);
xnor U14792 (N_14792,N_13673,N_13818);
or U14793 (N_14793,N_13793,N_13574);
and U14794 (N_14794,N_13937,N_13572);
or U14795 (N_14795,N_14061,N_13753);
nand U14796 (N_14796,N_14021,N_13895);
nand U14797 (N_14797,N_13659,N_13900);
or U14798 (N_14798,N_13987,N_13522);
or U14799 (N_14799,N_13931,N_14070);
nor U14800 (N_14800,N_13628,N_13622);
or U14801 (N_14801,N_13553,N_13800);
nand U14802 (N_14802,N_13505,N_13538);
nand U14803 (N_14803,N_14047,N_14191);
or U14804 (N_14804,N_13885,N_13909);
nand U14805 (N_14805,N_14165,N_13620);
nor U14806 (N_14806,N_13621,N_13894);
xor U14807 (N_14807,N_13783,N_14135);
xnor U14808 (N_14808,N_13691,N_14213);
or U14809 (N_14809,N_13892,N_13605);
nor U14810 (N_14810,N_13881,N_14223);
xnor U14811 (N_14811,N_14223,N_14175);
and U14812 (N_14812,N_13621,N_13893);
and U14813 (N_14813,N_14063,N_13552);
or U14814 (N_14814,N_13824,N_13656);
nand U14815 (N_14815,N_13586,N_13735);
or U14816 (N_14816,N_13565,N_14211);
nand U14817 (N_14817,N_14220,N_14075);
or U14818 (N_14818,N_13816,N_13586);
or U14819 (N_14819,N_14147,N_13771);
nor U14820 (N_14820,N_13880,N_13878);
and U14821 (N_14821,N_13513,N_14220);
nand U14822 (N_14822,N_14203,N_13504);
xnor U14823 (N_14823,N_13936,N_13980);
or U14824 (N_14824,N_13777,N_13700);
nand U14825 (N_14825,N_13701,N_14168);
and U14826 (N_14826,N_14158,N_13636);
nand U14827 (N_14827,N_13590,N_13759);
nor U14828 (N_14828,N_13855,N_13938);
xor U14829 (N_14829,N_14246,N_14125);
xnor U14830 (N_14830,N_14126,N_14084);
nand U14831 (N_14831,N_14092,N_14089);
xnor U14832 (N_14832,N_13613,N_13692);
and U14833 (N_14833,N_14105,N_13926);
nor U14834 (N_14834,N_13830,N_13562);
or U14835 (N_14835,N_13940,N_14072);
and U14836 (N_14836,N_14117,N_13546);
or U14837 (N_14837,N_13650,N_13710);
xor U14838 (N_14838,N_14201,N_13729);
nand U14839 (N_14839,N_14076,N_13864);
nand U14840 (N_14840,N_14149,N_14237);
and U14841 (N_14841,N_13774,N_13582);
nand U14842 (N_14842,N_13809,N_14095);
nand U14843 (N_14843,N_14098,N_14058);
and U14844 (N_14844,N_13736,N_13847);
xor U14845 (N_14845,N_13544,N_13759);
nand U14846 (N_14846,N_13603,N_14181);
nor U14847 (N_14847,N_14020,N_13968);
xnor U14848 (N_14848,N_13735,N_13695);
nand U14849 (N_14849,N_13685,N_14168);
nand U14850 (N_14850,N_13504,N_13610);
nand U14851 (N_14851,N_14120,N_13937);
xnor U14852 (N_14852,N_14160,N_13710);
xnor U14853 (N_14853,N_13525,N_13846);
nand U14854 (N_14854,N_13622,N_13724);
nor U14855 (N_14855,N_13811,N_13689);
and U14856 (N_14856,N_13776,N_14116);
or U14857 (N_14857,N_13985,N_13512);
or U14858 (N_14858,N_13752,N_13993);
nand U14859 (N_14859,N_13871,N_13643);
or U14860 (N_14860,N_13703,N_13843);
xnor U14861 (N_14861,N_13643,N_13894);
nor U14862 (N_14862,N_13592,N_14239);
nand U14863 (N_14863,N_14086,N_14142);
xnor U14864 (N_14864,N_14161,N_13814);
or U14865 (N_14865,N_13963,N_13980);
nand U14866 (N_14866,N_13510,N_13560);
nor U14867 (N_14867,N_13518,N_13766);
nand U14868 (N_14868,N_13669,N_13596);
and U14869 (N_14869,N_13591,N_13717);
nor U14870 (N_14870,N_14157,N_14170);
nor U14871 (N_14871,N_14176,N_13966);
nor U14872 (N_14872,N_13669,N_14023);
nor U14873 (N_14873,N_14088,N_13782);
nor U14874 (N_14874,N_14245,N_13763);
nor U14875 (N_14875,N_14211,N_14120);
xor U14876 (N_14876,N_14245,N_13505);
nor U14877 (N_14877,N_13883,N_13622);
or U14878 (N_14878,N_13728,N_13782);
xnor U14879 (N_14879,N_13992,N_13840);
or U14880 (N_14880,N_13652,N_13901);
nand U14881 (N_14881,N_13571,N_14192);
or U14882 (N_14882,N_13555,N_13613);
xnor U14883 (N_14883,N_13572,N_13610);
and U14884 (N_14884,N_14100,N_14017);
or U14885 (N_14885,N_13787,N_14179);
or U14886 (N_14886,N_14197,N_13662);
nor U14887 (N_14887,N_13718,N_13594);
nor U14888 (N_14888,N_14196,N_13644);
or U14889 (N_14889,N_13955,N_14157);
nor U14890 (N_14890,N_14124,N_14115);
xor U14891 (N_14891,N_13713,N_14127);
and U14892 (N_14892,N_14135,N_14147);
and U14893 (N_14893,N_14127,N_14021);
and U14894 (N_14894,N_13738,N_13618);
nand U14895 (N_14895,N_13987,N_14005);
and U14896 (N_14896,N_13732,N_13712);
or U14897 (N_14897,N_14074,N_13664);
or U14898 (N_14898,N_14007,N_13506);
nor U14899 (N_14899,N_13751,N_13621);
xor U14900 (N_14900,N_13937,N_13711);
nor U14901 (N_14901,N_13773,N_13590);
nor U14902 (N_14902,N_14055,N_14056);
nor U14903 (N_14903,N_14096,N_14161);
or U14904 (N_14904,N_13779,N_13575);
xnor U14905 (N_14905,N_14002,N_13911);
nor U14906 (N_14906,N_14231,N_14173);
and U14907 (N_14907,N_14208,N_13987);
or U14908 (N_14908,N_13641,N_13928);
nand U14909 (N_14909,N_13859,N_13807);
xnor U14910 (N_14910,N_13733,N_14149);
and U14911 (N_14911,N_13675,N_13695);
nor U14912 (N_14912,N_14134,N_13607);
nor U14913 (N_14913,N_13544,N_13872);
nor U14914 (N_14914,N_14237,N_14102);
nor U14915 (N_14915,N_13779,N_13700);
or U14916 (N_14916,N_14043,N_13836);
nor U14917 (N_14917,N_13937,N_13908);
or U14918 (N_14918,N_14101,N_14172);
nor U14919 (N_14919,N_14233,N_13569);
nand U14920 (N_14920,N_13890,N_14149);
or U14921 (N_14921,N_13617,N_13618);
or U14922 (N_14922,N_14091,N_14241);
nor U14923 (N_14923,N_13975,N_14126);
nor U14924 (N_14924,N_13967,N_13644);
or U14925 (N_14925,N_14064,N_13573);
xnor U14926 (N_14926,N_13848,N_13993);
nand U14927 (N_14927,N_13644,N_14122);
nor U14928 (N_14928,N_14227,N_13528);
and U14929 (N_14929,N_13943,N_14215);
xnor U14930 (N_14930,N_14154,N_13633);
nor U14931 (N_14931,N_14037,N_13792);
nand U14932 (N_14932,N_13503,N_13898);
and U14933 (N_14933,N_13694,N_14080);
xnor U14934 (N_14934,N_14139,N_14055);
and U14935 (N_14935,N_13857,N_13931);
or U14936 (N_14936,N_13663,N_14119);
nor U14937 (N_14937,N_13860,N_13916);
xor U14938 (N_14938,N_13821,N_14198);
and U14939 (N_14939,N_13907,N_14037);
xor U14940 (N_14940,N_13897,N_13658);
nor U14941 (N_14941,N_13956,N_14025);
or U14942 (N_14942,N_14147,N_13769);
nand U14943 (N_14943,N_13617,N_14056);
nor U14944 (N_14944,N_13767,N_14085);
nor U14945 (N_14945,N_13672,N_13633);
nand U14946 (N_14946,N_13920,N_14198);
nor U14947 (N_14947,N_13836,N_14015);
xor U14948 (N_14948,N_14146,N_14060);
and U14949 (N_14949,N_13670,N_14230);
nand U14950 (N_14950,N_13925,N_14198);
nor U14951 (N_14951,N_13935,N_14213);
nor U14952 (N_14952,N_13622,N_13819);
nor U14953 (N_14953,N_14065,N_14196);
nor U14954 (N_14954,N_14117,N_14006);
and U14955 (N_14955,N_13660,N_13604);
and U14956 (N_14956,N_13807,N_13511);
xnor U14957 (N_14957,N_13977,N_13541);
nor U14958 (N_14958,N_13657,N_13611);
and U14959 (N_14959,N_14152,N_14025);
nand U14960 (N_14960,N_13965,N_13531);
nand U14961 (N_14961,N_13691,N_14090);
and U14962 (N_14962,N_13825,N_13680);
and U14963 (N_14963,N_14048,N_13597);
xnor U14964 (N_14964,N_14117,N_13803);
or U14965 (N_14965,N_13703,N_13890);
or U14966 (N_14966,N_13794,N_13915);
nor U14967 (N_14967,N_14154,N_14198);
nor U14968 (N_14968,N_13963,N_13776);
and U14969 (N_14969,N_14058,N_13647);
or U14970 (N_14970,N_13535,N_13928);
nand U14971 (N_14971,N_14040,N_13944);
and U14972 (N_14972,N_14144,N_13883);
nand U14973 (N_14973,N_14159,N_13962);
xnor U14974 (N_14974,N_13885,N_13687);
xor U14975 (N_14975,N_14010,N_13757);
nor U14976 (N_14976,N_13646,N_13694);
or U14977 (N_14977,N_13756,N_14020);
xnor U14978 (N_14978,N_14054,N_14172);
and U14979 (N_14979,N_14229,N_14118);
and U14980 (N_14980,N_14175,N_13758);
nor U14981 (N_14981,N_14151,N_13642);
and U14982 (N_14982,N_14089,N_13569);
and U14983 (N_14983,N_14023,N_14051);
nor U14984 (N_14984,N_13828,N_13991);
xor U14985 (N_14985,N_14241,N_14181);
nor U14986 (N_14986,N_14203,N_13841);
nand U14987 (N_14987,N_13904,N_14144);
and U14988 (N_14988,N_13591,N_14230);
nor U14989 (N_14989,N_14131,N_13698);
or U14990 (N_14990,N_13770,N_13616);
or U14991 (N_14991,N_14021,N_13968);
and U14992 (N_14992,N_13679,N_13620);
xnor U14993 (N_14993,N_13575,N_14106);
nor U14994 (N_14994,N_14163,N_13669);
xor U14995 (N_14995,N_14189,N_13956);
nor U14996 (N_14996,N_13565,N_13761);
nand U14997 (N_14997,N_13886,N_13883);
nor U14998 (N_14998,N_13591,N_13708);
nand U14999 (N_14999,N_14052,N_14140);
or UO_0 (O_0,N_14523,N_14925);
xor UO_1 (O_1,N_14595,N_14656);
nor UO_2 (O_2,N_14463,N_14291);
and UO_3 (O_3,N_14581,N_14750);
nand UO_4 (O_4,N_14794,N_14579);
xor UO_5 (O_5,N_14888,N_14279);
nand UO_6 (O_6,N_14639,N_14452);
and UO_7 (O_7,N_14479,N_14828);
xor UO_8 (O_8,N_14364,N_14937);
xor UO_9 (O_9,N_14459,N_14723);
nor UO_10 (O_10,N_14552,N_14576);
nand UO_11 (O_11,N_14757,N_14669);
nand UO_12 (O_12,N_14896,N_14301);
and UO_13 (O_13,N_14252,N_14319);
xor UO_14 (O_14,N_14497,N_14704);
or UO_15 (O_15,N_14522,N_14670);
and UO_16 (O_16,N_14601,N_14640);
xor UO_17 (O_17,N_14843,N_14393);
or UO_18 (O_18,N_14876,N_14920);
or UO_19 (O_19,N_14995,N_14535);
nor UO_20 (O_20,N_14842,N_14740);
nor UO_21 (O_21,N_14744,N_14310);
or UO_22 (O_22,N_14830,N_14858);
nand UO_23 (O_23,N_14651,N_14625);
xor UO_24 (O_24,N_14336,N_14353);
and UO_25 (O_25,N_14267,N_14617);
nand UO_26 (O_26,N_14682,N_14702);
xnor UO_27 (O_27,N_14966,N_14558);
nand UO_28 (O_28,N_14915,N_14761);
xor UO_29 (O_29,N_14976,N_14919);
and UO_30 (O_30,N_14324,N_14492);
and UO_31 (O_31,N_14981,N_14356);
nand UO_32 (O_32,N_14499,N_14574);
and UO_33 (O_33,N_14362,N_14904);
and UO_34 (O_34,N_14378,N_14436);
nor UO_35 (O_35,N_14433,N_14564);
and UO_36 (O_36,N_14638,N_14802);
nand UO_37 (O_37,N_14275,N_14594);
and UO_38 (O_38,N_14837,N_14658);
and UO_39 (O_39,N_14792,N_14456);
xnor UO_40 (O_40,N_14565,N_14939);
or UO_41 (O_41,N_14630,N_14829);
nor UO_42 (O_42,N_14690,N_14355);
nor UO_43 (O_43,N_14898,N_14671);
nand UO_44 (O_44,N_14278,N_14367);
nand UO_45 (O_45,N_14664,N_14569);
and UO_46 (O_46,N_14890,N_14851);
nand UO_47 (O_47,N_14610,N_14504);
and UO_48 (O_48,N_14276,N_14636);
and UO_49 (O_49,N_14906,N_14606);
nand UO_50 (O_50,N_14728,N_14972);
xnor UO_51 (O_51,N_14485,N_14668);
nand UO_52 (O_52,N_14371,N_14605);
and UO_53 (O_53,N_14910,N_14697);
and UO_54 (O_54,N_14866,N_14844);
and UO_55 (O_55,N_14883,N_14780);
nor UO_56 (O_56,N_14831,N_14999);
nand UO_57 (O_57,N_14855,N_14650);
nor UO_58 (O_58,N_14345,N_14985);
and UO_59 (O_59,N_14806,N_14982);
nor UO_60 (O_60,N_14694,N_14897);
xor UO_61 (O_61,N_14977,N_14381);
and UO_62 (O_62,N_14681,N_14462);
nand UO_63 (O_63,N_14513,N_14397);
xnor UO_64 (O_64,N_14363,N_14996);
or UO_65 (O_65,N_14621,N_14445);
or UO_66 (O_66,N_14812,N_14608);
xor UO_67 (O_67,N_14454,N_14495);
and UO_68 (O_68,N_14785,N_14955);
nor UO_69 (O_69,N_14517,N_14783);
nand UO_70 (O_70,N_14788,N_14340);
xor UO_71 (O_71,N_14335,N_14416);
and UO_72 (O_72,N_14734,N_14347);
or UO_73 (O_73,N_14631,N_14867);
nor UO_74 (O_74,N_14566,N_14434);
and UO_75 (O_75,N_14420,N_14696);
nand UO_76 (O_76,N_14551,N_14753);
nor UO_77 (O_77,N_14816,N_14731);
and UO_78 (O_78,N_14795,N_14747);
nor UO_79 (O_79,N_14468,N_14877);
xor UO_80 (O_80,N_14776,N_14333);
xnor UO_81 (O_81,N_14758,N_14674);
and UO_82 (O_82,N_14325,N_14732);
nand UO_83 (O_83,N_14321,N_14289);
nand UO_84 (O_84,N_14789,N_14916);
or UO_85 (O_85,N_14975,N_14864);
and UO_86 (O_86,N_14845,N_14719);
xnor UO_87 (O_87,N_14269,N_14743);
and UO_88 (O_88,N_14717,N_14527);
xnor UO_89 (O_89,N_14438,N_14318);
xnor UO_90 (O_90,N_14911,N_14821);
or UO_91 (O_91,N_14368,N_14528);
xnor UO_92 (O_92,N_14797,N_14895);
and UO_93 (O_93,N_14341,N_14796);
or UO_94 (O_94,N_14263,N_14339);
and UO_95 (O_95,N_14823,N_14516);
or UO_96 (O_96,N_14251,N_14414);
nor UO_97 (O_97,N_14315,N_14997);
or UO_98 (O_98,N_14729,N_14483);
nand UO_99 (O_99,N_14450,N_14913);
xnor UO_100 (O_100,N_14612,N_14798);
nand UO_101 (O_101,N_14469,N_14466);
nor UO_102 (O_102,N_14666,N_14947);
or UO_103 (O_103,N_14305,N_14411);
nand UO_104 (O_104,N_14693,N_14592);
xnor UO_105 (O_105,N_14948,N_14692);
or UO_106 (O_106,N_14404,N_14423);
xor UO_107 (O_107,N_14460,N_14358);
xnor UO_108 (O_108,N_14502,N_14375);
nand UO_109 (O_109,N_14933,N_14507);
and UO_110 (O_110,N_14735,N_14860);
or UO_111 (O_111,N_14649,N_14603);
nor UO_112 (O_112,N_14964,N_14993);
and UO_113 (O_113,N_14529,N_14779);
and UO_114 (O_114,N_14715,N_14775);
nor UO_115 (O_115,N_14559,N_14924);
nand UO_116 (O_116,N_14457,N_14292);
nand UO_117 (O_117,N_14818,N_14607);
nand UO_118 (O_118,N_14412,N_14677);
xor UO_119 (O_119,N_14880,N_14721);
or UO_120 (O_120,N_14361,N_14632);
nor UO_121 (O_121,N_14394,N_14846);
nand UO_122 (O_122,N_14689,N_14865);
xnor UO_123 (O_123,N_14872,N_14629);
or UO_124 (O_124,N_14951,N_14871);
nand UO_125 (O_125,N_14474,N_14600);
nand UO_126 (O_126,N_14524,N_14426);
nor UO_127 (O_127,N_14988,N_14921);
xnor UO_128 (O_128,N_14893,N_14688);
nor UO_129 (O_129,N_14583,N_14489);
nor UO_130 (O_130,N_14328,N_14745);
or UO_131 (O_131,N_14334,N_14998);
xnor UO_132 (O_132,N_14954,N_14862);
or UO_133 (O_133,N_14399,N_14493);
xnor UO_134 (O_134,N_14444,N_14590);
xnor UO_135 (O_135,N_14756,N_14365);
nand UO_136 (O_136,N_14902,N_14446);
xor UO_137 (O_137,N_14699,N_14622);
and UO_138 (O_138,N_14769,N_14733);
and UO_139 (O_139,N_14873,N_14965);
xor UO_140 (O_140,N_14679,N_14317);
xnor UO_141 (O_141,N_14967,N_14882);
nor UO_142 (O_142,N_14406,N_14531);
or UO_143 (O_143,N_14277,N_14620);
or UO_144 (O_144,N_14773,N_14593);
xnor UO_145 (O_145,N_14891,N_14912);
and UO_146 (O_146,N_14707,N_14657);
and UO_147 (O_147,N_14793,N_14413);
xnor UO_148 (O_148,N_14992,N_14514);
nor UO_149 (O_149,N_14974,N_14766);
nor UO_150 (O_150,N_14401,N_14491);
or UO_151 (O_151,N_14598,N_14979);
or UO_152 (O_152,N_14519,N_14332);
nor UO_153 (O_153,N_14791,N_14659);
or UO_154 (O_154,N_14685,N_14518);
and UO_155 (O_155,N_14970,N_14398);
xor UO_156 (O_156,N_14953,N_14989);
nand UO_157 (O_157,N_14448,N_14560);
nor UO_158 (O_158,N_14313,N_14626);
nand UO_159 (O_159,N_14295,N_14991);
or UO_160 (O_160,N_14755,N_14359);
nand UO_161 (O_161,N_14691,N_14616);
nand UO_162 (O_162,N_14892,N_14280);
xor UO_163 (O_163,N_14567,N_14490);
nor UO_164 (O_164,N_14928,N_14548);
nand UO_165 (O_165,N_14856,N_14738);
xor UO_166 (O_166,N_14400,N_14348);
nor UO_167 (O_167,N_14298,N_14311);
nand UO_168 (O_168,N_14494,N_14908);
and UO_169 (O_169,N_14570,N_14418);
or UO_170 (O_170,N_14587,N_14817);
xnor UO_171 (O_171,N_14557,N_14562);
and UO_172 (O_172,N_14575,N_14323);
and UO_173 (O_173,N_14498,N_14346);
xor UO_174 (O_174,N_14945,N_14962);
nor UO_175 (O_175,N_14405,N_14409);
nor UO_176 (O_176,N_14377,N_14961);
nor UO_177 (O_177,N_14875,N_14665);
or UO_178 (O_178,N_14260,N_14765);
or UO_179 (O_179,N_14396,N_14754);
nor UO_180 (O_180,N_14922,N_14472);
nor UO_181 (O_181,N_14386,N_14442);
nor UO_182 (O_182,N_14774,N_14857);
and UO_183 (O_183,N_14710,N_14708);
xnor UO_184 (O_184,N_14534,N_14627);
nor UO_185 (O_185,N_14487,N_14455);
nor UO_186 (O_186,N_14419,N_14441);
xnor UO_187 (O_187,N_14663,N_14628);
xor UO_188 (O_188,N_14960,N_14563);
nand UO_189 (O_189,N_14547,N_14672);
or UO_190 (O_190,N_14431,N_14784);
xor UO_191 (O_191,N_14770,N_14648);
nand UO_192 (O_192,N_14471,N_14422);
nand UO_193 (O_193,N_14737,N_14477);
xnor UO_194 (O_194,N_14272,N_14990);
xor UO_195 (O_195,N_14834,N_14500);
xor UO_196 (O_196,N_14329,N_14453);
nor UO_197 (O_197,N_14934,N_14521);
nor UO_198 (O_198,N_14464,N_14884);
or UO_199 (O_199,N_14449,N_14326);
xor UO_200 (O_200,N_14597,N_14488);
nor UO_201 (O_201,N_14503,N_14684);
nand UO_202 (O_202,N_14841,N_14287);
xnor UO_203 (O_203,N_14833,N_14421);
nand UO_204 (O_204,N_14591,N_14297);
or UO_205 (O_205,N_14635,N_14768);
and UO_206 (O_206,N_14678,N_14923);
xnor UO_207 (O_207,N_14762,N_14941);
and UO_208 (O_208,N_14615,N_14555);
xnor UO_209 (O_209,N_14458,N_14899);
and UO_210 (O_210,N_14388,N_14585);
xor UO_211 (O_211,N_14777,N_14501);
or UO_212 (O_212,N_14473,N_14808);
nand UO_213 (O_213,N_14294,N_14847);
xnor UO_214 (O_214,N_14701,N_14771);
xor UO_215 (O_215,N_14868,N_14786);
and UO_216 (O_216,N_14811,N_14814);
nor UO_217 (O_217,N_14506,N_14901);
or UO_218 (O_218,N_14342,N_14568);
or UO_219 (O_219,N_14714,N_14722);
nand UO_220 (O_220,N_14379,N_14308);
xnor UO_221 (O_221,N_14619,N_14720);
and UO_222 (O_222,N_14253,N_14312);
nor UO_223 (O_223,N_14695,N_14512);
nor UO_224 (O_224,N_14447,N_14480);
nand UO_225 (O_225,N_14268,N_14285);
nor UO_226 (O_226,N_14571,N_14589);
and UO_227 (O_227,N_14614,N_14599);
nor UO_228 (O_228,N_14742,N_14536);
or UO_229 (O_229,N_14509,N_14652);
nor UO_230 (O_230,N_14475,N_14337);
nand UO_231 (O_231,N_14711,N_14767);
and UO_232 (O_232,N_14357,N_14374);
and UO_233 (O_233,N_14705,N_14609);
xnor UO_234 (O_234,N_14261,N_14546);
or UO_235 (O_235,N_14533,N_14271);
nand UO_236 (O_236,N_14799,N_14344);
and UO_237 (O_237,N_14800,N_14573);
xnor UO_238 (O_238,N_14886,N_14662);
nand UO_239 (O_239,N_14741,N_14259);
nor UO_240 (O_240,N_14957,N_14293);
or UO_241 (O_241,N_14752,N_14417);
xnor UO_242 (O_242,N_14376,N_14646);
and UO_243 (O_243,N_14926,N_14820);
xor UO_244 (O_244,N_14712,N_14623);
xor UO_245 (O_245,N_14577,N_14827);
nand UO_246 (O_246,N_14541,N_14424);
or UO_247 (O_247,N_14706,N_14903);
or UO_248 (O_248,N_14936,N_14309);
or UO_249 (O_249,N_14410,N_14320);
xnor UO_250 (O_250,N_14935,N_14716);
nand UO_251 (O_251,N_14994,N_14437);
and UO_252 (O_252,N_14804,N_14661);
xor UO_253 (O_253,N_14853,N_14395);
xnor UO_254 (O_254,N_14726,N_14327);
and UO_255 (O_255,N_14680,N_14542);
xnor UO_256 (O_256,N_14403,N_14983);
nor UO_257 (O_257,N_14703,N_14254);
nand UO_258 (O_258,N_14366,N_14971);
and UO_259 (O_259,N_14316,N_14407);
or UO_260 (O_260,N_14805,N_14476);
or UO_261 (O_261,N_14307,N_14968);
nor UO_262 (O_262,N_14380,N_14869);
nor UO_263 (O_263,N_14894,N_14382);
nand UO_264 (O_264,N_14515,N_14586);
nor UO_265 (O_265,N_14950,N_14584);
or UO_266 (O_266,N_14544,N_14984);
nand UO_267 (O_267,N_14304,N_14824);
nor UO_268 (O_268,N_14350,N_14660);
nand UO_269 (O_269,N_14430,N_14675);
nor UO_270 (O_270,N_14718,N_14807);
and UO_271 (O_271,N_14637,N_14730);
and UO_272 (O_272,N_14510,N_14931);
and UO_273 (O_273,N_14943,N_14451);
nand UO_274 (O_274,N_14763,N_14553);
xnor UO_275 (O_275,N_14633,N_14545);
and UO_276 (O_276,N_14554,N_14525);
xnor UO_277 (O_277,N_14713,N_14496);
and UO_278 (O_278,N_14874,N_14641);
and UO_279 (O_279,N_14314,N_14687);
or UO_280 (O_280,N_14508,N_14940);
or UO_281 (O_281,N_14250,N_14643);
nand UO_282 (O_282,N_14854,N_14618);
nor UO_283 (O_283,N_14838,N_14288);
or UO_284 (O_284,N_14461,N_14372);
and UO_285 (O_285,N_14848,N_14602);
nor UO_286 (O_286,N_14914,N_14343);
xnor UO_287 (O_287,N_14826,N_14978);
and UO_288 (O_288,N_14482,N_14302);
or UO_289 (O_289,N_14810,N_14739);
nand UO_290 (O_290,N_14905,N_14836);
and UO_291 (O_291,N_14486,N_14764);
xor UO_292 (O_292,N_14647,N_14949);
nor UO_293 (O_293,N_14959,N_14642);
xnor UO_294 (O_294,N_14852,N_14303);
and UO_295 (O_295,N_14539,N_14580);
xor UO_296 (O_296,N_14526,N_14540);
and UO_297 (O_297,N_14700,N_14790);
xor UO_298 (O_298,N_14909,N_14440);
or UO_299 (O_299,N_14863,N_14676);
nor UO_300 (O_300,N_14255,N_14849);
xor UO_301 (O_301,N_14942,N_14385);
or UO_302 (O_302,N_14927,N_14443);
nor UO_303 (O_303,N_14907,N_14484);
nand UO_304 (O_304,N_14822,N_14408);
nand UO_305 (O_305,N_14813,N_14987);
xnor UO_306 (O_306,N_14383,N_14384);
or UO_307 (O_307,N_14969,N_14391);
or UO_308 (O_308,N_14655,N_14653);
or UO_309 (O_309,N_14556,N_14481);
xnor UO_310 (O_310,N_14296,N_14415);
xor UO_311 (O_311,N_14859,N_14351);
xnor UO_312 (O_312,N_14322,N_14432);
or UO_313 (O_313,N_14736,N_14938);
nor UO_314 (O_314,N_14809,N_14465);
nand UO_315 (O_315,N_14425,N_14698);
or UO_316 (O_316,N_14505,N_14781);
xnor UO_317 (O_317,N_14283,N_14604);
or UO_318 (O_318,N_14958,N_14338);
nand UO_319 (O_319,N_14530,N_14819);
and UO_320 (O_320,N_14264,N_14299);
nor UO_321 (O_321,N_14944,N_14511);
or UO_322 (O_322,N_14889,N_14667);
and UO_323 (O_323,N_14917,N_14349);
nand UO_324 (O_324,N_14686,N_14946);
nand UO_325 (O_325,N_14624,N_14803);
or UO_326 (O_326,N_14963,N_14256);
xnor UO_327 (O_327,N_14429,N_14532);
nor UO_328 (O_328,N_14727,N_14582);
nor UO_329 (O_329,N_14273,N_14932);
nor UO_330 (O_330,N_14815,N_14900);
nor UO_331 (O_331,N_14759,N_14772);
nor UO_332 (O_332,N_14282,N_14390);
and UO_333 (O_333,N_14879,N_14262);
and UO_334 (O_334,N_14370,N_14266);
and UO_335 (O_335,N_14360,N_14478);
nor UO_336 (O_336,N_14258,N_14986);
nand UO_337 (O_337,N_14683,N_14265);
and UO_338 (O_338,N_14634,N_14550);
xnor UO_339 (O_339,N_14439,N_14596);
nand UO_340 (O_340,N_14832,N_14787);
nor UO_341 (O_341,N_14929,N_14537);
and UO_342 (O_342,N_14835,N_14520);
xnor UO_343 (O_343,N_14290,N_14952);
nand UO_344 (O_344,N_14782,N_14428);
and UO_345 (O_345,N_14257,N_14801);
nand UO_346 (O_346,N_14850,N_14746);
nor UO_347 (O_347,N_14930,N_14839);
nor UO_348 (O_348,N_14588,N_14878);
nand UO_349 (O_349,N_14725,N_14274);
nand UO_350 (O_350,N_14644,N_14392);
xor UO_351 (O_351,N_14467,N_14435);
and UO_352 (O_352,N_14543,N_14956);
nor UO_353 (O_353,N_14331,N_14760);
and UO_354 (O_354,N_14709,N_14549);
and UO_355 (O_355,N_14270,N_14284);
and UO_356 (O_356,N_14611,N_14470);
nand UO_357 (O_357,N_14840,N_14724);
nor UO_358 (O_358,N_14306,N_14613);
nor UO_359 (O_359,N_14373,N_14881);
nor UO_360 (O_360,N_14300,N_14973);
nand UO_361 (O_361,N_14885,N_14748);
or UO_362 (O_362,N_14330,N_14354);
and UO_363 (O_363,N_14861,N_14572);
and UO_364 (O_364,N_14402,N_14281);
nor UO_365 (O_365,N_14749,N_14751);
or UO_366 (O_366,N_14578,N_14918);
nor UO_367 (O_367,N_14369,N_14778);
and UO_368 (O_368,N_14389,N_14887);
xor UO_369 (O_369,N_14870,N_14645);
or UO_370 (O_370,N_14387,N_14561);
xor UO_371 (O_371,N_14352,N_14427);
nand UO_372 (O_372,N_14673,N_14538);
nand UO_373 (O_373,N_14980,N_14286);
xor UO_374 (O_374,N_14825,N_14654);
xnor UO_375 (O_375,N_14365,N_14608);
nor UO_376 (O_376,N_14455,N_14788);
and UO_377 (O_377,N_14867,N_14550);
nor UO_378 (O_378,N_14743,N_14381);
and UO_379 (O_379,N_14820,N_14407);
nand UO_380 (O_380,N_14950,N_14903);
and UO_381 (O_381,N_14788,N_14892);
or UO_382 (O_382,N_14843,N_14825);
or UO_383 (O_383,N_14920,N_14380);
xor UO_384 (O_384,N_14962,N_14804);
nor UO_385 (O_385,N_14634,N_14658);
xor UO_386 (O_386,N_14923,N_14362);
and UO_387 (O_387,N_14885,N_14547);
and UO_388 (O_388,N_14401,N_14863);
nand UO_389 (O_389,N_14347,N_14852);
or UO_390 (O_390,N_14983,N_14858);
nand UO_391 (O_391,N_14913,N_14884);
and UO_392 (O_392,N_14476,N_14937);
and UO_393 (O_393,N_14889,N_14948);
or UO_394 (O_394,N_14357,N_14444);
nor UO_395 (O_395,N_14740,N_14554);
nand UO_396 (O_396,N_14406,N_14980);
xor UO_397 (O_397,N_14308,N_14301);
xor UO_398 (O_398,N_14396,N_14810);
xor UO_399 (O_399,N_14256,N_14634);
nor UO_400 (O_400,N_14570,N_14361);
nand UO_401 (O_401,N_14407,N_14627);
nand UO_402 (O_402,N_14558,N_14322);
or UO_403 (O_403,N_14817,N_14709);
and UO_404 (O_404,N_14470,N_14281);
nand UO_405 (O_405,N_14805,N_14500);
or UO_406 (O_406,N_14780,N_14471);
xor UO_407 (O_407,N_14778,N_14715);
and UO_408 (O_408,N_14617,N_14944);
nand UO_409 (O_409,N_14682,N_14840);
nand UO_410 (O_410,N_14338,N_14954);
and UO_411 (O_411,N_14902,N_14813);
and UO_412 (O_412,N_14885,N_14327);
or UO_413 (O_413,N_14685,N_14479);
nand UO_414 (O_414,N_14284,N_14652);
and UO_415 (O_415,N_14557,N_14350);
and UO_416 (O_416,N_14747,N_14634);
xnor UO_417 (O_417,N_14738,N_14665);
nand UO_418 (O_418,N_14714,N_14892);
nor UO_419 (O_419,N_14848,N_14790);
xor UO_420 (O_420,N_14573,N_14930);
xor UO_421 (O_421,N_14847,N_14957);
nand UO_422 (O_422,N_14684,N_14706);
or UO_423 (O_423,N_14633,N_14382);
xnor UO_424 (O_424,N_14666,N_14355);
nand UO_425 (O_425,N_14366,N_14541);
and UO_426 (O_426,N_14453,N_14509);
xnor UO_427 (O_427,N_14277,N_14701);
xor UO_428 (O_428,N_14854,N_14455);
and UO_429 (O_429,N_14580,N_14705);
xnor UO_430 (O_430,N_14829,N_14717);
nand UO_431 (O_431,N_14706,N_14397);
xor UO_432 (O_432,N_14806,N_14470);
nor UO_433 (O_433,N_14412,N_14888);
and UO_434 (O_434,N_14408,N_14646);
xnor UO_435 (O_435,N_14406,N_14635);
xor UO_436 (O_436,N_14853,N_14770);
and UO_437 (O_437,N_14623,N_14340);
and UO_438 (O_438,N_14453,N_14268);
nand UO_439 (O_439,N_14678,N_14672);
and UO_440 (O_440,N_14946,N_14901);
or UO_441 (O_441,N_14992,N_14904);
nand UO_442 (O_442,N_14704,N_14262);
and UO_443 (O_443,N_14360,N_14738);
nor UO_444 (O_444,N_14822,N_14678);
xor UO_445 (O_445,N_14295,N_14897);
xnor UO_446 (O_446,N_14697,N_14686);
nand UO_447 (O_447,N_14769,N_14512);
nand UO_448 (O_448,N_14590,N_14552);
and UO_449 (O_449,N_14434,N_14485);
and UO_450 (O_450,N_14813,N_14984);
nand UO_451 (O_451,N_14541,N_14370);
nand UO_452 (O_452,N_14926,N_14987);
or UO_453 (O_453,N_14531,N_14466);
and UO_454 (O_454,N_14710,N_14784);
nor UO_455 (O_455,N_14353,N_14824);
nand UO_456 (O_456,N_14557,N_14271);
and UO_457 (O_457,N_14606,N_14481);
and UO_458 (O_458,N_14432,N_14284);
or UO_459 (O_459,N_14771,N_14931);
xnor UO_460 (O_460,N_14833,N_14656);
nand UO_461 (O_461,N_14368,N_14443);
xnor UO_462 (O_462,N_14966,N_14547);
nor UO_463 (O_463,N_14881,N_14736);
or UO_464 (O_464,N_14922,N_14766);
nor UO_465 (O_465,N_14931,N_14386);
nor UO_466 (O_466,N_14848,N_14256);
and UO_467 (O_467,N_14445,N_14836);
and UO_468 (O_468,N_14308,N_14797);
xor UO_469 (O_469,N_14855,N_14545);
nor UO_470 (O_470,N_14943,N_14789);
xor UO_471 (O_471,N_14814,N_14392);
xor UO_472 (O_472,N_14629,N_14351);
nor UO_473 (O_473,N_14804,N_14959);
and UO_474 (O_474,N_14289,N_14904);
nor UO_475 (O_475,N_14343,N_14773);
nand UO_476 (O_476,N_14433,N_14451);
xor UO_477 (O_477,N_14800,N_14551);
xor UO_478 (O_478,N_14956,N_14729);
nor UO_479 (O_479,N_14649,N_14744);
or UO_480 (O_480,N_14559,N_14903);
and UO_481 (O_481,N_14488,N_14346);
nor UO_482 (O_482,N_14966,N_14278);
nor UO_483 (O_483,N_14621,N_14466);
and UO_484 (O_484,N_14562,N_14454);
xnor UO_485 (O_485,N_14775,N_14755);
xor UO_486 (O_486,N_14534,N_14433);
nor UO_487 (O_487,N_14298,N_14329);
nor UO_488 (O_488,N_14969,N_14813);
nor UO_489 (O_489,N_14412,N_14266);
xor UO_490 (O_490,N_14688,N_14509);
nand UO_491 (O_491,N_14992,N_14558);
and UO_492 (O_492,N_14931,N_14758);
nor UO_493 (O_493,N_14568,N_14992);
nor UO_494 (O_494,N_14505,N_14836);
or UO_495 (O_495,N_14627,N_14671);
and UO_496 (O_496,N_14420,N_14796);
and UO_497 (O_497,N_14365,N_14699);
nor UO_498 (O_498,N_14538,N_14398);
nand UO_499 (O_499,N_14632,N_14868);
nor UO_500 (O_500,N_14410,N_14716);
nor UO_501 (O_501,N_14879,N_14531);
xor UO_502 (O_502,N_14297,N_14843);
nor UO_503 (O_503,N_14929,N_14861);
or UO_504 (O_504,N_14518,N_14863);
nand UO_505 (O_505,N_14345,N_14796);
nor UO_506 (O_506,N_14611,N_14326);
xor UO_507 (O_507,N_14381,N_14945);
nor UO_508 (O_508,N_14997,N_14466);
xor UO_509 (O_509,N_14351,N_14330);
nand UO_510 (O_510,N_14923,N_14391);
and UO_511 (O_511,N_14720,N_14587);
and UO_512 (O_512,N_14831,N_14913);
nor UO_513 (O_513,N_14675,N_14582);
nor UO_514 (O_514,N_14791,N_14631);
nand UO_515 (O_515,N_14977,N_14820);
and UO_516 (O_516,N_14547,N_14637);
xnor UO_517 (O_517,N_14783,N_14635);
xor UO_518 (O_518,N_14368,N_14261);
xnor UO_519 (O_519,N_14617,N_14940);
and UO_520 (O_520,N_14745,N_14502);
or UO_521 (O_521,N_14858,N_14833);
nor UO_522 (O_522,N_14493,N_14419);
nor UO_523 (O_523,N_14752,N_14582);
xor UO_524 (O_524,N_14312,N_14303);
nor UO_525 (O_525,N_14948,N_14506);
or UO_526 (O_526,N_14317,N_14840);
nand UO_527 (O_527,N_14816,N_14854);
or UO_528 (O_528,N_14312,N_14752);
nand UO_529 (O_529,N_14509,N_14620);
nand UO_530 (O_530,N_14798,N_14630);
nand UO_531 (O_531,N_14595,N_14865);
or UO_532 (O_532,N_14941,N_14367);
nand UO_533 (O_533,N_14925,N_14345);
nor UO_534 (O_534,N_14475,N_14349);
nor UO_535 (O_535,N_14567,N_14383);
nor UO_536 (O_536,N_14314,N_14757);
nor UO_537 (O_537,N_14295,N_14697);
nand UO_538 (O_538,N_14879,N_14991);
nor UO_539 (O_539,N_14685,N_14640);
or UO_540 (O_540,N_14441,N_14990);
nor UO_541 (O_541,N_14673,N_14412);
and UO_542 (O_542,N_14553,N_14824);
nand UO_543 (O_543,N_14780,N_14483);
xnor UO_544 (O_544,N_14512,N_14670);
and UO_545 (O_545,N_14279,N_14532);
nor UO_546 (O_546,N_14348,N_14925);
and UO_547 (O_547,N_14310,N_14539);
nand UO_548 (O_548,N_14933,N_14783);
or UO_549 (O_549,N_14535,N_14496);
nor UO_550 (O_550,N_14541,N_14985);
xnor UO_551 (O_551,N_14872,N_14838);
or UO_552 (O_552,N_14321,N_14831);
nand UO_553 (O_553,N_14797,N_14301);
nand UO_554 (O_554,N_14663,N_14393);
and UO_555 (O_555,N_14814,N_14950);
nand UO_556 (O_556,N_14261,N_14924);
nand UO_557 (O_557,N_14474,N_14636);
nor UO_558 (O_558,N_14463,N_14425);
and UO_559 (O_559,N_14296,N_14307);
or UO_560 (O_560,N_14251,N_14538);
xor UO_561 (O_561,N_14699,N_14999);
and UO_562 (O_562,N_14476,N_14614);
nor UO_563 (O_563,N_14764,N_14636);
nand UO_564 (O_564,N_14947,N_14632);
nand UO_565 (O_565,N_14397,N_14630);
and UO_566 (O_566,N_14753,N_14303);
nor UO_567 (O_567,N_14666,N_14754);
nor UO_568 (O_568,N_14504,N_14528);
xnor UO_569 (O_569,N_14672,N_14542);
and UO_570 (O_570,N_14850,N_14622);
or UO_571 (O_571,N_14758,N_14688);
nand UO_572 (O_572,N_14309,N_14810);
and UO_573 (O_573,N_14748,N_14975);
xnor UO_574 (O_574,N_14719,N_14563);
nand UO_575 (O_575,N_14805,N_14416);
and UO_576 (O_576,N_14321,N_14371);
and UO_577 (O_577,N_14570,N_14387);
nand UO_578 (O_578,N_14251,N_14505);
and UO_579 (O_579,N_14444,N_14374);
nor UO_580 (O_580,N_14276,N_14544);
xnor UO_581 (O_581,N_14320,N_14352);
nand UO_582 (O_582,N_14510,N_14995);
or UO_583 (O_583,N_14446,N_14302);
xor UO_584 (O_584,N_14451,N_14679);
nor UO_585 (O_585,N_14545,N_14751);
nand UO_586 (O_586,N_14942,N_14909);
or UO_587 (O_587,N_14470,N_14544);
and UO_588 (O_588,N_14992,N_14691);
xnor UO_589 (O_589,N_14509,N_14322);
or UO_590 (O_590,N_14815,N_14275);
nor UO_591 (O_591,N_14897,N_14911);
nand UO_592 (O_592,N_14470,N_14722);
or UO_593 (O_593,N_14384,N_14619);
nor UO_594 (O_594,N_14702,N_14631);
nand UO_595 (O_595,N_14284,N_14843);
xor UO_596 (O_596,N_14643,N_14481);
nand UO_597 (O_597,N_14911,N_14398);
or UO_598 (O_598,N_14929,N_14382);
nor UO_599 (O_599,N_14756,N_14968);
or UO_600 (O_600,N_14578,N_14304);
xor UO_601 (O_601,N_14974,N_14308);
and UO_602 (O_602,N_14711,N_14808);
xor UO_603 (O_603,N_14591,N_14436);
or UO_604 (O_604,N_14502,N_14537);
xor UO_605 (O_605,N_14773,N_14703);
nand UO_606 (O_606,N_14380,N_14388);
nor UO_607 (O_607,N_14376,N_14487);
or UO_608 (O_608,N_14902,N_14456);
xnor UO_609 (O_609,N_14559,N_14681);
or UO_610 (O_610,N_14563,N_14690);
xnor UO_611 (O_611,N_14678,N_14899);
nand UO_612 (O_612,N_14448,N_14435);
nand UO_613 (O_613,N_14988,N_14464);
or UO_614 (O_614,N_14447,N_14679);
nor UO_615 (O_615,N_14305,N_14683);
nand UO_616 (O_616,N_14504,N_14622);
xnor UO_617 (O_617,N_14804,N_14315);
xor UO_618 (O_618,N_14990,N_14488);
and UO_619 (O_619,N_14361,N_14595);
or UO_620 (O_620,N_14343,N_14292);
or UO_621 (O_621,N_14851,N_14867);
and UO_622 (O_622,N_14421,N_14500);
nor UO_623 (O_623,N_14626,N_14847);
or UO_624 (O_624,N_14495,N_14499);
or UO_625 (O_625,N_14824,N_14749);
and UO_626 (O_626,N_14548,N_14933);
or UO_627 (O_627,N_14713,N_14286);
nor UO_628 (O_628,N_14552,N_14869);
or UO_629 (O_629,N_14542,N_14769);
and UO_630 (O_630,N_14488,N_14899);
xnor UO_631 (O_631,N_14463,N_14771);
nor UO_632 (O_632,N_14427,N_14287);
xor UO_633 (O_633,N_14737,N_14860);
and UO_634 (O_634,N_14426,N_14882);
nor UO_635 (O_635,N_14332,N_14280);
and UO_636 (O_636,N_14326,N_14491);
or UO_637 (O_637,N_14760,N_14470);
nand UO_638 (O_638,N_14600,N_14496);
nand UO_639 (O_639,N_14934,N_14816);
or UO_640 (O_640,N_14339,N_14259);
and UO_641 (O_641,N_14571,N_14369);
nor UO_642 (O_642,N_14311,N_14336);
nand UO_643 (O_643,N_14976,N_14273);
and UO_644 (O_644,N_14852,N_14743);
xor UO_645 (O_645,N_14738,N_14337);
and UO_646 (O_646,N_14397,N_14262);
nand UO_647 (O_647,N_14685,N_14629);
or UO_648 (O_648,N_14500,N_14671);
xnor UO_649 (O_649,N_14784,N_14940);
nor UO_650 (O_650,N_14687,N_14953);
xnor UO_651 (O_651,N_14286,N_14590);
nor UO_652 (O_652,N_14813,N_14630);
nand UO_653 (O_653,N_14412,N_14429);
xnor UO_654 (O_654,N_14884,N_14643);
nor UO_655 (O_655,N_14661,N_14757);
nand UO_656 (O_656,N_14430,N_14829);
nand UO_657 (O_657,N_14691,N_14572);
nor UO_658 (O_658,N_14854,N_14405);
or UO_659 (O_659,N_14467,N_14933);
nor UO_660 (O_660,N_14610,N_14934);
nand UO_661 (O_661,N_14259,N_14758);
or UO_662 (O_662,N_14826,N_14960);
nand UO_663 (O_663,N_14472,N_14338);
or UO_664 (O_664,N_14340,N_14592);
nor UO_665 (O_665,N_14512,N_14642);
nor UO_666 (O_666,N_14867,N_14293);
xor UO_667 (O_667,N_14309,N_14992);
nand UO_668 (O_668,N_14308,N_14536);
nand UO_669 (O_669,N_14927,N_14802);
xnor UO_670 (O_670,N_14276,N_14938);
and UO_671 (O_671,N_14460,N_14771);
nor UO_672 (O_672,N_14489,N_14760);
or UO_673 (O_673,N_14280,N_14775);
and UO_674 (O_674,N_14815,N_14551);
nand UO_675 (O_675,N_14442,N_14869);
nor UO_676 (O_676,N_14623,N_14601);
nor UO_677 (O_677,N_14983,N_14425);
xnor UO_678 (O_678,N_14955,N_14975);
and UO_679 (O_679,N_14454,N_14694);
nor UO_680 (O_680,N_14353,N_14345);
nand UO_681 (O_681,N_14515,N_14778);
nand UO_682 (O_682,N_14888,N_14663);
nor UO_683 (O_683,N_14444,N_14340);
nor UO_684 (O_684,N_14936,N_14713);
and UO_685 (O_685,N_14389,N_14953);
nand UO_686 (O_686,N_14615,N_14605);
and UO_687 (O_687,N_14482,N_14838);
or UO_688 (O_688,N_14725,N_14964);
nor UO_689 (O_689,N_14380,N_14773);
xnor UO_690 (O_690,N_14574,N_14930);
nor UO_691 (O_691,N_14908,N_14538);
nor UO_692 (O_692,N_14718,N_14505);
xor UO_693 (O_693,N_14951,N_14773);
or UO_694 (O_694,N_14558,N_14653);
or UO_695 (O_695,N_14393,N_14482);
nor UO_696 (O_696,N_14282,N_14584);
xnor UO_697 (O_697,N_14495,N_14915);
or UO_698 (O_698,N_14703,N_14628);
nand UO_699 (O_699,N_14417,N_14770);
nor UO_700 (O_700,N_14346,N_14378);
or UO_701 (O_701,N_14455,N_14291);
nor UO_702 (O_702,N_14405,N_14709);
nand UO_703 (O_703,N_14739,N_14987);
xor UO_704 (O_704,N_14319,N_14802);
xor UO_705 (O_705,N_14688,N_14456);
xor UO_706 (O_706,N_14646,N_14891);
nor UO_707 (O_707,N_14403,N_14961);
xnor UO_708 (O_708,N_14282,N_14436);
and UO_709 (O_709,N_14825,N_14525);
nand UO_710 (O_710,N_14642,N_14308);
nor UO_711 (O_711,N_14810,N_14627);
or UO_712 (O_712,N_14783,N_14950);
nand UO_713 (O_713,N_14989,N_14938);
nand UO_714 (O_714,N_14406,N_14615);
and UO_715 (O_715,N_14540,N_14270);
xor UO_716 (O_716,N_14507,N_14359);
or UO_717 (O_717,N_14803,N_14586);
and UO_718 (O_718,N_14683,N_14818);
nand UO_719 (O_719,N_14971,N_14621);
and UO_720 (O_720,N_14954,N_14799);
xor UO_721 (O_721,N_14494,N_14730);
or UO_722 (O_722,N_14387,N_14526);
nor UO_723 (O_723,N_14450,N_14369);
xor UO_724 (O_724,N_14823,N_14948);
xor UO_725 (O_725,N_14373,N_14640);
and UO_726 (O_726,N_14283,N_14560);
nand UO_727 (O_727,N_14515,N_14360);
and UO_728 (O_728,N_14583,N_14966);
nand UO_729 (O_729,N_14392,N_14414);
nand UO_730 (O_730,N_14317,N_14539);
and UO_731 (O_731,N_14356,N_14989);
xor UO_732 (O_732,N_14658,N_14959);
nor UO_733 (O_733,N_14806,N_14792);
nand UO_734 (O_734,N_14378,N_14696);
and UO_735 (O_735,N_14851,N_14706);
and UO_736 (O_736,N_14932,N_14356);
xnor UO_737 (O_737,N_14659,N_14809);
nand UO_738 (O_738,N_14549,N_14270);
xnor UO_739 (O_739,N_14878,N_14523);
nor UO_740 (O_740,N_14253,N_14894);
or UO_741 (O_741,N_14308,N_14467);
and UO_742 (O_742,N_14710,N_14855);
nand UO_743 (O_743,N_14568,N_14664);
nand UO_744 (O_744,N_14466,N_14947);
or UO_745 (O_745,N_14953,N_14836);
nand UO_746 (O_746,N_14281,N_14713);
nand UO_747 (O_747,N_14689,N_14952);
nand UO_748 (O_748,N_14319,N_14777);
or UO_749 (O_749,N_14796,N_14665);
or UO_750 (O_750,N_14544,N_14607);
and UO_751 (O_751,N_14774,N_14939);
nand UO_752 (O_752,N_14751,N_14484);
and UO_753 (O_753,N_14813,N_14814);
or UO_754 (O_754,N_14407,N_14611);
or UO_755 (O_755,N_14834,N_14563);
and UO_756 (O_756,N_14909,N_14438);
or UO_757 (O_757,N_14548,N_14772);
nand UO_758 (O_758,N_14485,N_14381);
or UO_759 (O_759,N_14498,N_14456);
nor UO_760 (O_760,N_14428,N_14795);
nand UO_761 (O_761,N_14380,N_14853);
or UO_762 (O_762,N_14949,N_14396);
nand UO_763 (O_763,N_14324,N_14419);
nand UO_764 (O_764,N_14525,N_14276);
or UO_765 (O_765,N_14612,N_14906);
and UO_766 (O_766,N_14626,N_14998);
and UO_767 (O_767,N_14433,N_14351);
nor UO_768 (O_768,N_14643,N_14489);
nand UO_769 (O_769,N_14590,N_14554);
and UO_770 (O_770,N_14482,N_14929);
nand UO_771 (O_771,N_14686,N_14714);
nor UO_772 (O_772,N_14821,N_14689);
or UO_773 (O_773,N_14337,N_14955);
or UO_774 (O_774,N_14761,N_14380);
or UO_775 (O_775,N_14823,N_14922);
nand UO_776 (O_776,N_14389,N_14444);
or UO_777 (O_777,N_14715,N_14253);
nor UO_778 (O_778,N_14549,N_14738);
and UO_779 (O_779,N_14852,N_14908);
nand UO_780 (O_780,N_14897,N_14472);
or UO_781 (O_781,N_14820,N_14348);
nor UO_782 (O_782,N_14737,N_14974);
and UO_783 (O_783,N_14913,N_14316);
nor UO_784 (O_784,N_14665,N_14834);
nand UO_785 (O_785,N_14319,N_14448);
nor UO_786 (O_786,N_14269,N_14457);
nor UO_787 (O_787,N_14699,N_14874);
nor UO_788 (O_788,N_14455,N_14960);
xor UO_789 (O_789,N_14362,N_14462);
xnor UO_790 (O_790,N_14494,N_14673);
xnor UO_791 (O_791,N_14535,N_14278);
or UO_792 (O_792,N_14970,N_14577);
or UO_793 (O_793,N_14853,N_14595);
nand UO_794 (O_794,N_14515,N_14651);
xnor UO_795 (O_795,N_14749,N_14921);
nor UO_796 (O_796,N_14980,N_14422);
nor UO_797 (O_797,N_14672,N_14960);
and UO_798 (O_798,N_14553,N_14973);
or UO_799 (O_799,N_14936,N_14280);
or UO_800 (O_800,N_14893,N_14697);
nand UO_801 (O_801,N_14726,N_14687);
nor UO_802 (O_802,N_14582,N_14571);
and UO_803 (O_803,N_14652,N_14303);
or UO_804 (O_804,N_14745,N_14558);
or UO_805 (O_805,N_14674,N_14975);
xor UO_806 (O_806,N_14679,N_14588);
nand UO_807 (O_807,N_14290,N_14423);
nand UO_808 (O_808,N_14506,N_14612);
nand UO_809 (O_809,N_14498,N_14823);
nor UO_810 (O_810,N_14628,N_14884);
nor UO_811 (O_811,N_14686,N_14663);
and UO_812 (O_812,N_14261,N_14271);
nand UO_813 (O_813,N_14373,N_14349);
nand UO_814 (O_814,N_14493,N_14327);
nand UO_815 (O_815,N_14970,N_14653);
xor UO_816 (O_816,N_14734,N_14687);
or UO_817 (O_817,N_14324,N_14989);
xnor UO_818 (O_818,N_14791,N_14688);
or UO_819 (O_819,N_14639,N_14367);
nand UO_820 (O_820,N_14808,N_14306);
nor UO_821 (O_821,N_14628,N_14742);
and UO_822 (O_822,N_14710,N_14990);
and UO_823 (O_823,N_14564,N_14510);
xor UO_824 (O_824,N_14486,N_14796);
nor UO_825 (O_825,N_14339,N_14880);
xor UO_826 (O_826,N_14267,N_14711);
nand UO_827 (O_827,N_14980,N_14862);
and UO_828 (O_828,N_14418,N_14486);
xor UO_829 (O_829,N_14298,N_14802);
and UO_830 (O_830,N_14957,N_14816);
nor UO_831 (O_831,N_14705,N_14781);
nor UO_832 (O_832,N_14386,N_14483);
and UO_833 (O_833,N_14316,N_14997);
xnor UO_834 (O_834,N_14920,N_14841);
and UO_835 (O_835,N_14883,N_14811);
xor UO_836 (O_836,N_14546,N_14370);
and UO_837 (O_837,N_14678,N_14384);
nor UO_838 (O_838,N_14525,N_14388);
xnor UO_839 (O_839,N_14395,N_14251);
and UO_840 (O_840,N_14430,N_14460);
nor UO_841 (O_841,N_14772,N_14326);
or UO_842 (O_842,N_14550,N_14332);
and UO_843 (O_843,N_14702,N_14412);
and UO_844 (O_844,N_14929,N_14579);
nand UO_845 (O_845,N_14421,N_14788);
and UO_846 (O_846,N_14518,N_14675);
or UO_847 (O_847,N_14723,N_14771);
and UO_848 (O_848,N_14606,N_14987);
nor UO_849 (O_849,N_14295,N_14501);
nand UO_850 (O_850,N_14518,N_14642);
nor UO_851 (O_851,N_14698,N_14545);
or UO_852 (O_852,N_14745,N_14459);
or UO_853 (O_853,N_14992,N_14687);
nand UO_854 (O_854,N_14572,N_14308);
and UO_855 (O_855,N_14457,N_14974);
and UO_856 (O_856,N_14861,N_14557);
and UO_857 (O_857,N_14418,N_14446);
nor UO_858 (O_858,N_14749,N_14566);
and UO_859 (O_859,N_14991,N_14943);
nor UO_860 (O_860,N_14409,N_14496);
or UO_861 (O_861,N_14541,N_14983);
nor UO_862 (O_862,N_14749,N_14442);
nand UO_863 (O_863,N_14454,N_14565);
nand UO_864 (O_864,N_14261,N_14512);
nor UO_865 (O_865,N_14921,N_14307);
nand UO_866 (O_866,N_14863,N_14283);
xnor UO_867 (O_867,N_14632,N_14608);
xor UO_868 (O_868,N_14840,N_14717);
xnor UO_869 (O_869,N_14496,N_14415);
xor UO_870 (O_870,N_14506,N_14895);
nand UO_871 (O_871,N_14270,N_14993);
xor UO_872 (O_872,N_14658,N_14570);
and UO_873 (O_873,N_14643,N_14579);
nor UO_874 (O_874,N_14286,N_14418);
xnor UO_875 (O_875,N_14294,N_14644);
xor UO_876 (O_876,N_14507,N_14470);
and UO_877 (O_877,N_14867,N_14619);
nor UO_878 (O_878,N_14661,N_14642);
nor UO_879 (O_879,N_14590,N_14737);
and UO_880 (O_880,N_14430,N_14975);
nand UO_881 (O_881,N_14466,N_14936);
or UO_882 (O_882,N_14669,N_14579);
or UO_883 (O_883,N_14776,N_14519);
and UO_884 (O_884,N_14931,N_14811);
or UO_885 (O_885,N_14755,N_14684);
and UO_886 (O_886,N_14540,N_14394);
or UO_887 (O_887,N_14669,N_14277);
or UO_888 (O_888,N_14280,N_14774);
or UO_889 (O_889,N_14386,N_14715);
nand UO_890 (O_890,N_14677,N_14263);
xnor UO_891 (O_891,N_14737,N_14383);
xor UO_892 (O_892,N_14590,N_14280);
or UO_893 (O_893,N_14690,N_14601);
nor UO_894 (O_894,N_14614,N_14792);
nand UO_895 (O_895,N_14978,N_14962);
nand UO_896 (O_896,N_14847,N_14701);
nor UO_897 (O_897,N_14322,N_14924);
xor UO_898 (O_898,N_14714,N_14349);
and UO_899 (O_899,N_14954,N_14335);
and UO_900 (O_900,N_14770,N_14858);
xnor UO_901 (O_901,N_14887,N_14729);
and UO_902 (O_902,N_14380,N_14631);
xnor UO_903 (O_903,N_14907,N_14540);
nor UO_904 (O_904,N_14446,N_14443);
xnor UO_905 (O_905,N_14706,N_14548);
xor UO_906 (O_906,N_14423,N_14646);
nor UO_907 (O_907,N_14514,N_14422);
and UO_908 (O_908,N_14432,N_14867);
xnor UO_909 (O_909,N_14692,N_14775);
or UO_910 (O_910,N_14896,N_14662);
nand UO_911 (O_911,N_14531,N_14250);
or UO_912 (O_912,N_14253,N_14460);
and UO_913 (O_913,N_14792,N_14677);
and UO_914 (O_914,N_14761,N_14394);
nor UO_915 (O_915,N_14485,N_14707);
nand UO_916 (O_916,N_14494,N_14331);
xnor UO_917 (O_917,N_14632,N_14428);
and UO_918 (O_918,N_14444,N_14332);
nand UO_919 (O_919,N_14694,N_14518);
nor UO_920 (O_920,N_14573,N_14658);
nand UO_921 (O_921,N_14943,N_14622);
xor UO_922 (O_922,N_14826,N_14401);
nor UO_923 (O_923,N_14845,N_14634);
nor UO_924 (O_924,N_14477,N_14265);
xor UO_925 (O_925,N_14551,N_14915);
nor UO_926 (O_926,N_14920,N_14523);
nand UO_927 (O_927,N_14626,N_14652);
nand UO_928 (O_928,N_14639,N_14670);
nand UO_929 (O_929,N_14959,N_14269);
xor UO_930 (O_930,N_14727,N_14938);
nand UO_931 (O_931,N_14464,N_14943);
and UO_932 (O_932,N_14328,N_14562);
or UO_933 (O_933,N_14520,N_14948);
xnor UO_934 (O_934,N_14451,N_14489);
nor UO_935 (O_935,N_14820,N_14821);
xor UO_936 (O_936,N_14664,N_14519);
nor UO_937 (O_937,N_14294,N_14727);
nor UO_938 (O_938,N_14394,N_14731);
nand UO_939 (O_939,N_14411,N_14307);
nor UO_940 (O_940,N_14255,N_14575);
nand UO_941 (O_941,N_14575,N_14689);
or UO_942 (O_942,N_14981,N_14749);
nor UO_943 (O_943,N_14838,N_14543);
nand UO_944 (O_944,N_14718,N_14306);
nand UO_945 (O_945,N_14641,N_14875);
xor UO_946 (O_946,N_14367,N_14747);
xnor UO_947 (O_947,N_14551,N_14715);
or UO_948 (O_948,N_14655,N_14866);
nor UO_949 (O_949,N_14806,N_14657);
nand UO_950 (O_950,N_14405,N_14634);
nand UO_951 (O_951,N_14489,N_14939);
xnor UO_952 (O_952,N_14581,N_14298);
or UO_953 (O_953,N_14381,N_14882);
xnor UO_954 (O_954,N_14366,N_14270);
and UO_955 (O_955,N_14414,N_14817);
xor UO_956 (O_956,N_14754,N_14367);
or UO_957 (O_957,N_14807,N_14770);
xnor UO_958 (O_958,N_14954,N_14453);
xnor UO_959 (O_959,N_14354,N_14895);
nand UO_960 (O_960,N_14625,N_14710);
and UO_961 (O_961,N_14747,N_14315);
or UO_962 (O_962,N_14445,N_14574);
xor UO_963 (O_963,N_14409,N_14569);
xor UO_964 (O_964,N_14341,N_14688);
nand UO_965 (O_965,N_14547,N_14422);
or UO_966 (O_966,N_14777,N_14591);
and UO_967 (O_967,N_14439,N_14503);
nor UO_968 (O_968,N_14699,N_14751);
nand UO_969 (O_969,N_14810,N_14853);
xnor UO_970 (O_970,N_14863,N_14673);
nor UO_971 (O_971,N_14997,N_14745);
nand UO_972 (O_972,N_14717,N_14431);
and UO_973 (O_973,N_14716,N_14512);
and UO_974 (O_974,N_14399,N_14255);
nor UO_975 (O_975,N_14994,N_14646);
nor UO_976 (O_976,N_14798,N_14268);
nand UO_977 (O_977,N_14275,N_14510);
nand UO_978 (O_978,N_14687,N_14740);
and UO_979 (O_979,N_14826,N_14643);
and UO_980 (O_980,N_14985,N_14858);
xor UO_981 (O_981,N_14353,N_14267);
xor UO_982 (O_982,N_14787,N_14259);
and UO_983 (O_983,N_14423,N_14730);
nor UO_984 (O_984,N_14782,N_14775);
or UO_985 (O_985,N_14386,N_14436);
nor UO_986 (O_986,N_14930,N_14684);
xnor UO_987 (O_987,N_14324,N_14893);
and UO_988 (O_988,N_14291,N_14384);
and UO_989 (O_989,N_14761,N_14665);
and UO_990 (O_990,N_14756,N_14459);
xnor UO_991 (O_991,N_14590,N_14521);
nand UO_992 (O_992,N_14832,N_14637);
xor UO_993 (O_993,N_14575,N_14875);
or UO_994 (O_994,N_14855,N_14937);
nand UO_995 (O_995,N_14303,N_14440);
or UO_996 (O_996,N_14830,N_14396);
or UO_997 (O_997,N_14709,N_14487);
xnor UO_998 (O_998,N_14460,N_14377);
or UO_999 (O_999,N_14639,N_14723);
or UO_1000 (O_1000,N_14894,N_14660);
and UO_1001 (O_1001,N_14311,N_14769);
and UO_1002 (O_1002,N_14895,N_14359);
xnor UO_1003 (O_1003,N_14940,N_14389);
or UO_1004 (O_1004,N_14269,N_14914);
xnor UO_1005 (O_1005,N_14492,N_14630);
nand UO_1006 (O_1006,N_14362,N_14836);
nand UO_1007 (O_1007,N_14574,N_14871);
nand UO_1008 (O_1008,N_14944,N_14760);
nor UO_1009 (O_1009,N_14901,N_14697);
xor UO_1010 (O_1010,N_14259,N_14526);
and UO_1011 (O_1011,N_14264,N_14501);
and UO_1012 (O_1012,N_14533,N_14463);
or UO_1013 (O_1013,N_14256,N_14929);
or UO_1014 (O_1014,N_14467,N_14708);
and UO_1015 (O_1015,N_14745,N_14430);
nand UO_1016 (O_1016,N_14906,N_14273);
nand UO_1017 (O_1017,N_14299,N_14753);
xnor UO_1018 (O_1018,N_14969,N_14637);
xnor UO_1019 (O_1019,N_14776,N_14259);
xor UO_1020 (O_1020,N_14983,N_14282);
or UO_1021 (O_1021,N_14434,N_14956);
nand UO_1022 (O_1022,N_14928,N_14938);
or UO_1023 (O_1023,N_14263,N_14368);
nand UO_1024 (O_1024,N_14897,N_14812);
xnor UO_1025 (O_1025,N_14723,N_14376);
xnor UO_1026 (O_1026,N_14418,N_14724);
or UO_1027 (O_1027,N_14641,N_14274);
nor UO_1028 (O_1028,N_14881,N_14448);
nor UO_1029 (O_1029,N_14972,N_14268);
or UO_1030 (O_1030,N_14532,N_14553);
xnor UO_1031 (O_1031,N_14367,N_14252);
nor UO_1032 (O_1032,N_14691,N_14410);
or UO_1033 (O_1033,N_14548,N_14286);
nor UO_1034 (O_1034,N_14886,N_14761);
or UO_1035 (O_1035,N_14495,N_14330);
nor UO_1036 (O_1036,N_14467,N_14456);
nor UO_1037 (O_1037,N_14358,N_14457);
or UO_1038 (O_1038,N_14669,N_14515);
nor UO_1039 (O_1039,N_14439,N_14835);
nand UO_1040 (O_1040,N_14275,N_14990);
nand UO_1041 (O_1041,N_14433,N_14865);
nor UO_1042 (O_1042,N_14457,N_14661);
xnor UO_1043 (O_1043,N_14536,N_14465);
and UO_1044 (O_1044,N_14527,N_14640);
and UO_1045 (O_1045,N_14265,N_14614);
or UO_1046 (O_1046,N_14612,N_14557);
nor UO_1047 (O_1047,N_14560,N_14524);
nor UO_1048 (O_1048,N_14780,N_14672);
nand UO_1049 (O_1049,N_14486,N_14364);
and UO_1050 (O_1050,N_14406,N_14640);
nor UO_1051 (O_1051,N_14288,N_14351);
or UO_1052 (O_1052,N_14735,N_14797);
or UO_1053 (O_1053,N_14980,N_14523);
xnor UO_1054 (O_1054,N_14467,N_14314);
nor UO_1055 (O_1055,N_14371,N_14781);
xor UO_1056 (O_1056,N_14996,N_14652);
or UO_1057 (O_1057,N_14850,N_14421);
or UO_1058 (O_1058,N_14566,N_14744);
xnor UO_1059 (O_1059,N_14836,N_14528);
and UO_1060 (O_1060,N_14561,N_14575);
nand UO_1061 (O_1061,N_14842,N_14255);
nor UO_1062 (O_1062,N_14896,N_14250);
nand UO_1063 (O_1063,N_14587,N_14651);
or UO_1064 (O_1064,N_14829,N_14501);
or UO_1065 (O_1065,N_14997,N_14593);
or UO_1066 (O_1066,N_14421,N_14916);
nand UO_1067 (O_1067,N_14723,N_14281);
nor UO_1068 (O_1068,N_14977,N_14279);
nand UO_1069 (O_1069,N_14598,N_14911);
and UO_1070 (O_1070,N_14957,N_14885);
or UO_1071 (O_1071,N_14908,N_14899);
and UO_1072 (O_1072,N_14883,N_14307);
nor UO_1073 (O_1073,N_14521,N_14764);
nand UO_1074 (O_1074,N_14332,N_14962);
nand UO_1075 (O_1075,N_14514,N_14634);
nor UO_1076 (O_1076,N_14627,N_14992);
and UO_1077 (O_1077,N_14910,N_14503);
nand UO_1078 (O_1078,N_14962,N_14750);
nor UO_1079 (O_1079,N_14657,N_14898);
xnor UO_1080 (O_1080,N_14253,N_14757);
nand UO_1081 (O_1081,N_14644,N_14942);
or UO_1082 (O_1082,N_14733,N_14286);
and UO_1083 (O_1083,N_14799,N_14690);
xor UO_1084 (O_1084,N_14467,N_14736);
and UO_1085 (O_1085,N_14613,N_14311);
nand UO_1086 (O_1086,N_14965,N_14424);
nor UO_1087 (O_1087,N_14980,N_14932);
and UO_1088 (O_1088,N_14496,N_14987);
nor UO_1089 (O_1089,N_14897,N_14847);
nand UO_1090 (O_1090,N_14767,N_14590);
xnor UO_1091 (O_1091,N_14928,N_14748);
or UO_1092 (O_1092,N_14462,N_14969);
or UO_1093 (O_1093,N_14287,N_14353);
or UO_1094 (O_1094,N_14815,N_14511);
or UO_1095 (O_1095,N_14647,N_14714);
xnor UO_1096 (O_1096,N_14440,N_14925);
xnor UO_1097 (O_1097,N_14611,N_14613);
and UO_1098 (O_1098,N_14501,N_14268);
nor UO_1099 (O_1099,N_14471,N_14415);
or UO_1100 (O_1100,N_14533,N_14493);
and UO_1101 (O_1101,N_14267,N_14499);
nand UO_1102 (O_1102,N_14946,N_14478);
xor UO_1103 (O_1103,N_14972,N_14464);
xnor UO_1104 (O_1104,N_14759,N_14871);
nand UO_1105 (O_1105,N_14883,N_14374);
nor UO_1106 (O_1106,N_14659,N_14824);
and UO_1107 (O_1107,N_14614,N_14520);
or UO_1108 (O_1108,N_14347,N_14311);
nor UO_1109 (O_1109,N_14656,N_14631);
xnor UO_1110 (O_1110,N_14703,N_14723);
or UO_1111 (O_1111,N_14794,N_14814);
nand UO_1112 (O_1112,N_14904,N_14471);
or UO_1113 (O_1113,N_14927,N_14459);
nand UO_1114 (O_1114,N_14815,N_14855);
nand UO_1115 (O_1115,N_14655,N_14621);
or UO_1116 (O_1116,N_14646,N_14318);
and UO_1117 (O_1117,N_14376,N_14278);
nand UO_1118 (O_1118,N_14447,N_14953);
nor UO_1119 (O_1119,N_14313,N_14406);
xnor UO_1120 (O_1120,N_14384,N_14789);
and UO_1121 (O_1121,N_14356,N_14312);
or UO_1122 (O_1122,N_14584,N_14295);
and UO_1123 (O_1123,N_14698,N_14459);
or UO_1124 (O_1124,N_14463,N_14614);
or UO_1125 (O_1125,N_14988,N_14743);
nand UO_1126 (O_1126,N_14816,N_14374);
xor UO_1127 (O_1127,N_14280,N_14677);
and UO_1128 (O_1128,N_14322,N_14680);
nand UO_1129 (O_1129,N_14686,N_14645);
and UO_1130 (O_1130,N_14833,N_14880);
or UO_1131 (O_1131,N_14277,N_14801);
and UO_1132 (O_1132,N_14922,N_14618);
and UO_1133 (O_1133,N_14636,N_14261);
nand UO_1134 (O_1134,N_14942,N_14303);
xnor UO_1135 (O_1135,N_14812,N_14625);
or UO_1136 (O_1136,N_14654,N_14675);
nor UO_1137 (O_1137,N_14545,N_14690);
xnor UO_1138 (O_1138,N_14941,N_14646);
and UO_1139 (O_1139,N_14539,N_14428);
xnor UO_1140 (O_1140,N_14863,N_14713);
nor UO_1141 (O_1141,N_14852,N_14975);
nor UO_1142 (O_1142,N_14418,N_14521);
nor UO_1143 (O_1143,N_14250,N_14999);
xor UO_1144 (O_1144,N_14447,N_14433);
or UO_1145 (O_1145,N_14539,N_14493);
nor UO_1146 (O_1146,N_14427,N_14536);
and UO_1147 (O_1147,N_14593,N_14465);
or UO_1148 (O_1148,N_14830,N_14652);
nor UO_1149 (O_1149,N_14417,N_14685);
and UO_1150 (O_1150,N_14736,N_14424);
nand UO_1151 (O_1151,N_14721,N_14987);
nand UO_1152 (O_1152,N_14818,N_14322);
nand UO_1153 (O_1153,N_14717,N_14554);
and UO_1154 (O_1154,N_14578,N_14889);
or UO_1155 (O_1155,N_14382,N_14990);
nand UO_1156 (O_1156,N_14388,N_14277);
nor UO_1157 (O_1157,N_14537,N_14525);
and UO_1158 (O_1158,N_14277,N_14412);
xnor UO_1159 (O_1159,N_14394,N_14770);
nor UO_1160 (O_1160,N_14865,N_14783);
nor UO_1161 (O_1161,N_14470,N_14803);
and UO_1162 (O_1162,N_14887,N_14274);
nor UO_1163 (O_1163,N_14772,N_14903);
nand UO_1164 (O_1164,N_14258,N_14288);
and UO_1165 (O_1165,N_14305,N_14999);
nor UO_1166 (O_1166,N_14335,N_14348);
or UO_1167 (O_1167,N_14593,N_14535);
xnor UO_1168 (O_1168,N_14456,N_14416);
or UO_1169 (O_1169,N_14371,N_14799);
and UO_1170 (O_1170,N_14849,N_14513);
nand UO_1171 (O_1171,N_14407,N_14281);
xnor UO_1172 (O_1172,N_14492,N_14723);
nand UO_1173 (O_1173,N_14882,N_14932);
xor UO_1174 (O_1174,N_14411,N_14470);
or UO_1175 (O_1175,N_14700,N_14455);
nand UO_1176 (O_1176,N_14439,N_14787);
nor UO_1177 (O_1177,N_14776,N_14623);
nand UO_1178 (O_1178,N_14780,N_14357);
nand UO_1179 (O_1179,N_14708,N_14548);
nand UO_1180 (O_1180,N_14585,N_14596);
and UO_1181 (O_1181,N_14483,N_14869);
or UO_1182 (O_1182,N_14982,N_14519);
xor UO_1183 (O_1183,N_14884,N_14331);
nor UO_1184 (O_1184,N_14336,N_14967);
xor UO_1185 (O_1185,N_14829,N_14681);
nor UO_1186 (O_1186,N_14656,N_14265);
nand UO_1187 (O_1187,N_14492,N_14485);
nor UO_1188 (O_1188,N_14717,N_14873);
xor UO_1189 (O_1189,N_14367,N_14616);
and UO_1190 (O_1190,N_14858,N_14757);
nor UO_1191 (O_1191,N_14358,N_14730);
nor UO_1192 (O_1192,N_14471,N_14891);
nand UO_1193 (O_1193,N_14933,N_14931);
or UO_1194 (O_1194,N_14959,N_14772);
and UO_1195 (O_1195,N_14799,N_14521);
nor UO_1196 (O_1196,N_14393,N_14530);
or UO_1197 (O_1197,N_14731,N_14704);
xor UO_1198 (O_1198,N_14491,N_14968);
xor UO_1199 (O_1199,N_14564,N_14763);
or UO_1200 (O_1200,N_14430,N_14328);
nor UO_1201 (O_1201,N_14874,N_14252);
nor UO_1202 (O_1202,N_14326,N_14934);
nand UO_1203 (O_1203,N_14479,N_14477);
nor UO_1204 (O_1204,N_14672,N_14947);
and UO_1205 (O_1205,N_14406,N_14948);
nand UO_1206 (O_1206,N_14566,N_14409);
or UO_1207 (O_1207,N_14978,N_14522);
and UO_1208 (O_1208,N_14569,N_14478);
nand UO_1209 (O_1209,N_14723,N_14958);
xor UO_1210 (O_1210,N_14453,N_14463);
nand UO_1211 (O_1211,N_14776,N_14861);
and UO_1212 (O_1212,N_14968,N_14262);
nor UO_1213 (O_1213,N_14792,N_14661);
xnor UO_1214 (O_1214,N_14722,N_14933);
and UO_1215 (O_1215,N_14552,N_14835);
nor UO_1216 (O_1216,N_14587,N_14254);
or UO_1217 (O_1217,N_14722,N_14475);
xnor UO_1218 (O_1218,N_14651,N_14596);
and UO_1219 (O_1219,N_14936,N_14786);
xnor UO_1220 (O_1220,N_14634,N_14294);
xnor UO_1221 (O_1221,N_14675,N_14944);
or UO_1222 (O_1222,N_14660,N_14519);
and UO_1223 (O_1223,N_14816,N_14602);
xnor UO_1224 (O_1224,N_14376,N_14804);
nor UO_1225 (O_1225,N_14470,N_14909);
nand UO_1226 (O_1226,N_14759,N_14946);
or UO_1227 (O_1227,N_14771,N_14753);
nor UO_1228 (O_1228,N_14514,N_14431);
xnor UO_1229 (O_1229,N_14819,N_14549);
or UO_1230 (O_1230,N_14947,N_14757);
and UO_1231 (O_1231,N_14597,N_14517);
nand UO_1232 (O_1232,N_14717,N_14471);
or UO_1233 (O_1233,N_14988,N_14683);
or UO_1234 (O_1234,N_14790,N_14720);
and UO_1235 (O_1235,N_14823,N_14666);
and UO_1236 (O_1236,N_14647,N_14815);
xnor UO_1237 (O_1237,N_14723,N_14853);
nor UO_1238 (O_1238,N_14402,N_14778);
or UO_1239 (O_1239,N_14533,N_14943);
nand UO_1240 (O_1240,N_14808,N_14913);
xnor UO_1241 (O_1241,N_14588,N_14478);
and UO_1242 (O_1242,N_14833,N_14785);
nand UO_1243 (O_1243,N_14635,N_14720);
and UO_1244 (O_1244,N_14364,N_14971);
xnor UO_1245 (O_1245,N_14788,N_14860);
and UO_1246 (O_1246,N_14687,N_14896);
nor UO_1247 (O_1247,N_14845,N_14469);
nand UO_1248 (O_1248,N_14633,N_14360);
or UO_1249 (O_1249,N_14430,N_14266);
and UO_1250 (O_1250,N_14737,N_14768);
nor UO_1251 (O_1251,N_14677,N_14498);
xor UO_1252 (O_1252,N_14969,N_14706);
or UO_1253 (O_1253,N_14620,N_14665);
and UO_1254 (O_1254,N_14499,N_14798);
nor UO_1255 (O_1255,N_14871,N_14263);
and UO_1256 (O_1256,N_14308,N_14626);
nand UO_1257 (O_1257,N_14306,N_14394);
or UO_1258 (O_1258,N_14409,N_14472);
nor UO_1259 (O_1259,N_14457,N_14674);
xor UO_1260 (O_1260,N_14563,N_14447);
and UO_1261 (O_1261,N_14782,N_14617);
and UO_1262 (O_1262,N_14367,N_14299);
nand UO_1263 (O_1263,N_14895,N_14326);
or UO_1264 (O_1264,N_14277,N_14302);
and UO_1265 (O_1265,N_14861,N_14962);
xnor UO_1266 (O_1266,N_14620,N_14698);
xnor UO_1267 (O_1267,N_14944,N_14319);
nor UO_1268 (O_1268,N_14564,N_14913);
xnor UO_1269 (O_1269,N_14286,N_14488);
or UO_1270 (O_1270,N_14933,N_14798);
and UO_1271 (O_1271,N_14875,N_14720);
or UO_1272 (O_1272,N_14474,N_14527);
xnor UO_1273 (O_1273,N_14668,N_14886);
xnor UO_1274 (O_1274,N_14907,N_14547);
nand UO_1275 (O_1275,N_14579,N_14746);
nand UO_1276 (O_1276,N_14958,N_14941);
nor UO_1277 (O_1277,N_14929,N_14481);
xor UO_1278 (O_1278,N_14418,N_14546);
or UO_1279 (O_1279,N_14533,N_14355);
or UO_1280 (O_1280,N_14716,N_14406);
xnor UO_1281 (O_1281,N_14633,N_14530);
nand UO_1282 (O_1282,N_14785,N_14439);
xor UO_1283 (O_1283,N_14775,N_14784);
nand UO_1284 (O_1284,N_14640,N_14519);
or UO_1285 (O_1285,N_14901,N_14257);
or UO_1286 (O_1286,N_14381,N_14484);
xor UO_1287 (O_1287,N_14301,N_14819);
xor UO_1288 (O_1288,N_14367,N_14322);
nor UO_1289 (O_1289,N_14308,N_14554);
or UO_1290 (O_1290,N_14801,N_14281);
nor UO_1291 (O_1291,N_14427,N_14765);
nor UO_1292 (O_1292,N_14346,N_14967);
nor UO_1293 (O_1293,N_14984,N_14961);
nor UO_1294 (O_1294,N_14565,N_14576);
and UO_1295 (O_1295,N_14652,N_14961);
nand UO_1296 (O_1296,N_14585,N_14616);
xnor UO_1297 (O_1297,N_14777,N_14935);
or UO_1298 (O_1298,N_14663,N_14724);
or UO_1299 (O_1299,N_14469,N_14532);
nor UO_1300 (O_1300,N_14309,N_14827);
nand UO_1301 (O_1301,N_14992,N_14807);
nor UO_1302 (O_1302,N_14488,N_14707);
or UO_1303 (O_1303,N_14423,N_14806);
nor UO_1304 (O_1304,N_14466,N_14478);
or UO_1305 (O_1305,N_14416,N_14437);
xnor UO_1306 (O_1306,N_14719,N_14931);
or UO_1307 (O_1307,N_14973,N_14772);
nor UO_1308 (O_1308,N_14867,N_14303);
or UO_1309 (O_1309,N_14928,N_14853);
and UO_1310 (O_1310,N_14484,N_14939);
nand UO_1311 (O_1311,N_14880,N_14602);
xnor UO_1312 (O_1312,N_14289,N_14485);
nand UO_1313 (O_1313,N_14407,N_14575);
or UO_1314 (O_1314,N_14362,N_14642);
nor UO_1315 (O_1315,N_14504,N_14755);
or UO_1316 (O_1316,N_14799,N_14919);
xnor UO_1317 (O_1317,N_14403,N_14661);
or UO_1318 (O_1318,N_14372,N_14438);
or UO_1319 (O_1319,N_14456,N_14841);
and UO_1320 (O_1320,N_14843,N_14732);
nor UO_1321 (O_1321,N_14954,N_14627);
nor UO_1322 (O_1322,N_14439,N_14563);
nand UO_1323 (O_1323,N_14257,N_14896);
and UO_1324 (O_1324,N_14721,N_14900);
xnor UO_1325 (O_1325,N_14264,N_14510);
nand UO_1326 (O_1326,N_14515,N_14250);
nand UO_1327 (O_1327,N_14702,N_14506);
or UO_1328 (O_1328,N_14688,N_14465);
xnor UO_1329 (O_1329,N_14929,N_14756);
nor UO_1330 (O_1330,N_14404,N_14762);
nor UO_1331 (O_1331,N_14377,N_14613);
xnor UO_1332 (O_1332,N_14451,N_14579);
or UO_1333 (O_1333,N_14927,N_14293);
nand UO_1334 (O_1334,N_14384,N_14410);
and UO_1335 (O_1335,N_14258,N_14570);
or UO_1336 (O_1336,N_14802,N_14294);
nor UO_1337 (O_1337,N_14641,N_14867);
or UO_1338 (O_1338,N_14704,N_14749);
nand UO_1339 (O_1339,N_14982,N_14406);
and UO_1340 (O_1340,N_14442,N_14976);
nor UO_1341 (O_1341,N_14607,N_14764);
and UO_1342 (O_1342,N_14636,N_14565);
or UO_1343 (O_1343,N_14381,N_14753);
or UO_1344 (O_1344,N_14490,N_14705);
nor UO_1345 (O_1345,N_14705,N_14944);
and UO_1346 (O_1346,N_14764,N_14930);
or UO_1347 (O_1347,N_14371,N_14484);
nor UO_1348 (O_1348,N_14557,N_14664);
and UO_1349 (O_1349,N_14663,N_14921);
nor UO_1350 (O_1350,N_14559,N_14968);
nand UO_1351 (O_1351,N_14647,N_14610);
nand UO_1352 (O_1352,N_14577,N_14869);
nand UO_1353 (O_1353,N_14997,N_14618);
or UO_1354 (O_1354,N_14470,N_14433);
xnor UO_1355 (O_1355,N_14584,N_14504);
or UO_1356 (O_1356,N_14677,N_14344);
nor UO_1357 (O_1357,N_14980,N_14797);
xnor UO_1358 (O_1358,N_14951,N_14936);
or UO_1359 (O_1359,N_14401,N_14758);
nor UO_1360 (O_1360,N_14917,N_14828);
nand UO_1361 (O_1361,N_14452,N_14581);
xnor UO_1362 (O_1362,N_14646,N_14717);
nor UO_1363 (O_1363,N_14805,N_14956);
or UO_1364 (O_1364,N_14701,N_14631);
xor UO_1365 (O_1365,N_14677,N_14511);
and UO_1366 (O_1366,N_14631,N_14816);
and UO_1367 (O_1367,N_14497,N_14926);
and UO_1368 (O_1368,N_14984,N_14442);
nor UO_1369 (O_1369,N_14606,N_14948);
xor UO_1370 (O_1370,N_14612,N_14708);
and UO_1371 (O_1371,N_14745,N_14254);
nor UO_1372 (O_1372,N_14739,N_14566);
xor UO_1373 (O_1373,N_14788,N_14322);
and UO_1374 (O_1374,N_14980,N_14965);
nand UO_1375 (O_1375,N_14596,N_14792);
and UO_1376 (O_1376,N_14496,N_14800);
or UO_1377 (O_1377,N_14415,N_14485);
nand UO_1378 (O_1378,N_14590,N_14582);
or UO_1379 (O_1379,N_14811,N_14927);
and UO_1380 (O_1380,N_14301,N_14849);
nor UO_1381 (O_1381,N_14569,N_14807);
xnor UO_1382 (O_1382,N_14814,N_14892);
nand UO_1383 (O_1383,N_14768,N_14295);
and UO_1384 (O_1384,N_14255,N_14526);
and UO_1385 (O_1385,N_14987,N_14310);
nor UO_1386 (O_1386,N_14843,N_14515);
nand UO_1387 (O_1387,N_14918,N_14936);
nand UO_1388 (O_1388,N_14505,N_14737);
and UO_1389 (O_1389,N_14959,N_14849);
nor UO_1390 (O_1390,N_14354,N_14421);
nand UO_1391 (O_1391,N_14903,N_14429);
or UO_1392 (O_1392,N_14880,N_14468);
xnor UO_1393 (O_1393,N_14800,N_14709);
nand UO_1394 (O_1394,N_14562,N_14754);
or UO_1395 (O_1395,N_14853,N_14484);
nor UO_1396 (O_1396,N_14305,N_14308);
or UO_1397 (O_1397,N_14515,N_14468);
nand UO_1398 (O_1398,N_14349,N_14735);
nand UO_1399 (O_1399,N_14703,N_14673);
and UO_1400 (O_1400,N_14905,N_14607);
and UO_1401 (O_1401,N_14460,N_14432);
xnor UO_1402 (O_1402,N_14828,N_14321);
nor UO_1403 (O_1403,N_14868,N_14452);
xnor UO_1404 (O_1404,N_14474,N_14442);
or UO_1405 (O_1405,N_14969,N_14614);
nor UO_1406 (O_1406,N_14790,N_14326);
and UO_1407 (O_1407,N_14958,N_14569);
and UO_1408 (O_1408,N_14503,N_14811);
nor UO_1409 (O_1409,N_14906,N_14487);
xnor UO_1410 (O_1410,N_14783,N_14728);
or UO_1411 (O_1411,N_14872,N_14733);
nor UO_1412 (O_1412,N_14802,N_14395);
and UO_1413 (O_1413,N_14912,N_14702);
or UO_1414 (O_1414,N_14688,N_14926);
nand UO_1415 (O_1415,N_14952,N_14745);
nor UO_1416 (O_1416,N_14398,N_14302);
and UO_1417 (O_1417,N_14572,N_14453);
and UO_1418 (O_1418,N_14623,N_14797);
xnor UO_1419 (O_1419,N_14815,N_14889);
or UO_1420 (O_1420,N_14372,N_14331);
or UO_1421 (O_1421,N_14734,N_14973);
or UO_1422 (O_1422,N_14291,N_14907);
nor UO_1423 (O_1423,N_14685,N_14929);
nand UO_1424 (O_1424,N_14535,N_14740);
nand UO_1425 (O_1425,N_14575,N_14858);
and UO_1426 (O_1426,N_14622,N_14732);
or UO_1427 (O_1427,N_14285,N_14683);
xor UO_1428 (O_1428,N_14634,N_14812);
and UO_1429 (O_1429,N_14826,N_14612);
xnor UO_1430 (O_1430,N_14860,N_14856);
and UO_1431 (O_1431,N_14692,N_14662);
and UO_1432 (O_1432,N_14783,N_14431);
and UO_1433 (O_1433,N_14286,N_14883);
nand UO_1434 (O_1434,N_14606,N_14501);
nand UO_1435 (O_1435,N_14456,N_14995);
and UO_1436 (O_1436,N_14907,N_14298);
xnor UO_1437 (O_1437,N_14285,N_14492);
or UO_1438 (O_1438,N_14471,N_14712);
and UO_1439 (O_1439,N_14927,N_14292);
nand UO_1440 (O_1440,N_14980,N_14897);
or UO_1441 (O_1441,N_14761,N_14481);
or UO_1442 (O_1442,N_14630,N_14560);
xnor UO_1443 (O_1443,N_14527,N_14948);
nand UO_1444 (O_1444,N_14864,N_14749);
or UO_1445 (O_1445,N_14567,N_14272);
xnor UO_1446 (O_1446,N_14276,N_14637);
nor UO_1447 (O_1447,N_14280,N_14605);
and UO_1448 (O_1448,N_14649,N_14259);
or UO_1449 (O_1449,N_14331,N_14604);
nor UO_1450 (O_1450,N_14862,N_14775);
nand UO_1451 (O_1451,N_14375,N_14738);
and UO_1452 (O_1452,N_14340,N_14380);
nand UO_1453 (O_1453,N_14950,N_14602);
nor UO_1454 (O_1454,N_14639,N_14708);
or UO_1455 (O_1455,N_14429,N_14402);
xnor UO_1456 (O_1456,N_14645,N_14783);
nor UO_1457 (O_1457,N_14677,N_14841);
nand UO_1458 (O_1458,N_14676,N_14324);
and UO_1459 (O_1459,N_14602,N_14846);
or UO_1460 (O_1460,N_14485,N_14895);
and UO_1461 (O_1461,N_14384,N_14849);
nand UO_1462 (O_1462,N_14380,N_14983);
or UO_1463 (O_1463,N_14684,N_14698);
xnor UO_1464 (O_1464,N_14498,N_14644);
and UO_1465 (O_1465,N_14935,N_14839);
xor UO_1466 (O_1466,N_14553,N_14501);
or UO_1467 (O_1467,N_14663,N_14795);
nor UO_1468 (O_1468,N_14716,N_14964);
xnor UO_1469 (O_1469,N_14871,N_14710);
nor UO_1470 (O_1470,N_14910,N_14703);
nor UO_1471 (O_1471,N_14686,N_14315);
nor UO_1472 (O_1472,N_14830,N_14536);
and UO_1473 (O_1473,N_14716,N_14993);
xnor UO_1474 (O_1474,N_14437,N_14604);
and UO_1475 (O_1475,N_14935,N_14275);
nor UO_1476 (O_1476,N_14606,N_14797);
nand UO_1477 (O_1477,N_14402,N_14881);
or UO_1478 (O_1478,N_14942,N_14673);
nand UO_1479 (O_1479,N_14669,N_14564);
or UO_1480 (O_1480,N_14391,N_14361);
nor UO_1481 (O_1481,N_14358,N_14411);
and UO_1482 (O_1482,N_14771,N_14486);
nand UO_1483 (O_1483,N_14500,N_14999);
nor UO_1484 (O_1484,N_14752,N_14436);
and UO_1485 (O_1485,N_14552,N_14652);
or UO_1486 (O_1486,N_14577,N_14329);
xor UO_1487 (O_1487,N_14916,N_14735);
nand UO_1488 (O_1488,N_14258,N_14813);
and UO_1489 (O_1489,N_14555,N_14730);
nor UO_1490 (O_1490,N_14784,N_14648);
xnor UO_1491 (O_1491,N_14261,N_14558);
xor UO_1492 (O_1492,N_14953,N_14403);
nand UO_1493 (O_1493,N_14859,N_14431);
xnor UO_1494 (O_1494,N_14792,N_14354);
or UO_1495 (O_1495,N_14563,N_14254);
xor UO_1496 (O_1496,N_14685,N_14638);
or UO_1497 (O_1497,N_14455,N_14727);
xor UO_1498 (O_1498,N_14527,N_14563);
and UO_1499 (O_1499,N_14441,N_14271);
or UO_1500 (O_1500,N_14889,N_14976);
xor UO_1501 (O_1501,N_14714,N_14491);
nand UO_1502 (O_1502,N_14630,N_14943);
xnor UO_1503 (O_1503,N_14344,N_14880);
nand UO_1504 (O_1504,N_14743,N_14874);
nor UO_1505 (O_1505,N_14977,N_14565);
or UO_1506 (O_1506,N_14308,N_14961);
nand UO_1507 (O_1507,N_14933,N_14681);
xor UO_1508 (O_1508,N_14443,N_14394);
or UO_1509 (O_1509,N_14813,N_14732);
nor UO_1510 (O_1510,N_14399,N_14530);
nand UO_1511 (O_1511,N_14705,N_14402);
nand UO_1512 (O_1512,N_14353,N_14724);
nand UO_1513 (O_1513,N_14410,N_14288);
xnor UO_1514 (O_1514,N_14444,N_14426);
and UO_1515 (O_1515,N_14318,N_14430);
nor UO_1516 (O_1516,N_14634,N_14710);
nor UO_1517 (O_1517,N_14756,N_14651);
and UO_1518 (O_1518,N_14749,N_14778);
xnor UO_1519 (O_1519,N_14607,N_14432);
nand UO_1520 (O_1520,N_14491,N_14408);
xnor UO_1521 (O_1521,N_14456,N_14551);
and UO_1522 (O_1522,N_14487,N_14744);
xnor UO_1523 (O_1523,N_14392,N_14977);
and UO_1524 (O_1524,N_14575,N_14482);
nand UO_1525 (O_1525,N_14373,N_14780);
nand UO_1526 (O_1526,N_14643,N_14668);
xnor UO_1527 (O_1527,N_14455,N_14944);
nand UO_1528 (O_1528,N_14263,N_14279);
nand UO_1529 (O_1529,N_14502,N_14563);
and UO_1530 (O_1530,N_14665,N_14395);
and UO_1531 (O_1531,N_14334,N_14488);
nor UO_1532 (O_1532,N_14729,N_14613);
nor UO_1533 (O_1533,N_14620,N_14585);
nand UO_1534 (O_1534,N_14797,N_14451);
nand UO_1535 (O_1535,N_14375,N_14980);
nand UO_1536 (O_1536,N_14886,N_14547);
and UO_1537 (O_1537,N_14665,N_14641);
or UO_1538 (O_1538,N_14529,N_14922);
nor UO_1539 (O_1539,N_14914,N_14304);
nor UO_1540 (O_1540,N_14817,N_14410);
nor UO_1541 (O_1541,N_14664,N_14773);
or UO_1542 (O_1542,N_14670,N_14857);
and UO_1543 (O_1543,N_14991,N_14841);
and UO_1544 (O_1544,N_14805,N_14320);
or UO_1545 (O_1545,N_14732,N_14424);
nand UO_1546 (O_1546,N_14814,N_14973);
xor UO_1547 (O_1547,N_14581,N_14916);
xnor UO_1548 (O_1548,N_14837,N_14359);
or UO_1549 (O_1549,N_14604,N_14910);
and UO_1550 (O_1550,N_14690,N_14663);
xor UO_1551 (O_1551,N_14895,N_14429);
or UO_1552 (O_1552,N_14642,N_14866);
xor UO_1553 (O_1553,N_14752,N_14653);
nor UO_1554 (O_1554,N_14510,N_14805);
or UO_1555 (O_1555,N_14263,N_14940);
nor UO_1556 (O_1556,N_14767,N_14604);
nor UO_1557 (O_1557,N_14788,N_14936);
xor UO_1558 (O_1558,N_14647,N_14434);
xnor UO_1559 (O_1559,N_14336,N_14983);
or UO_1560 (O_1560,N_14563,N_14583);
or UO_1561 (O_1561,N_14421,N_14892);
and UO_1562 (O_1562,N_14787,N_14827);
nand UO_1563 (O_1563,N_14928,N_14960);
nor UO_1564 (O_1564,N_14729,N_14487);
and UO_1565 (O_1565,N_14597,N_14444);
nand UO_1566 (O_1566,N_14898,N_14309);
xnor UO_1567 (O_1567,N_14340,N_14852);
xor UO_1568 (O_1568,N_14520,N_14344);
or UO_1569 (O_1569,N_14572,N_14669);
xnor UO_1570 (O_1570,N_14725,N_14548);
nand UO_1571 (O_1571,N_14567,N_14797);
or UO_1572 (O_1572,N_14320,N_14375);
or UO_1573 (O_1573,N_14968,N_14708);
and UO_1574 (O_1574,N_14276,N_14504);
and UO_1575 (O_1575,N_14700,N_14480);
nor UO_1576 (O_1576,N_14589,N_14608);
nor UO_1577 (O_1577,N_14773,N_14322);
nor UO_1578 (O_1578,N_14591,N_14811);
or UO_1579 (O_1579,N_14767,N_14902);
or UO_1580 (O_1580,N_14747,N_14944);
or UO_1581 (O_1581,N_14850,N_14578);
and UO_1582 (O_1582,N_14560,N_14405);
nand UO_1583 (O_1583,N_14884,N_14715);
nor UO_1584 (O_1584,N_14299,N_14383);
nor UO_1585 (O_1585,N_14415,N_14398);
xnor UO_1586 (O_1586,N_14664,N_14274);
and UO_1587 (O_1587,N_14362,N_14335);
or UO_1588 (O_1588,N_14543,N_14988);
nand UO_1589 (O_1589,N_14313,N_14974);
nor UO_1590 (O_1590,N_14359,N_14980);
nand UO_1591 (O_1591,N_14964,N_14691);
nand UO_1592 (O_1592,N_14293,N_14888);
xor UO_1593 (O_1593,N_14924,N_14579);
nor UO_1594 (O_1594,N_14359,N_14878);
or UO_1595 (O_1595,N_14998,N_14868);
nand UO_1596 (O_1596,N_14376,N_14747);
and UO_1597 (O_1597,N_14275,N_14898);
nand UO_1598 (O_1598,N_14553,N_14717);
xnor UO_1599 (O_1599,N_14344,N_14900);
xor UO_1600 (O_1600,N_14738,N_14653);
or UO_1601 (O_1601,N_14640,N_14739);
nand UO_1602 (O_1602,N_14518,N_14697);
nand UO_1603 (O_1603,N_14915,N_14346);
or UO_1604 (O_1604,N_14600,N_14934);
xnor UO_1605 (O_1605,N_14587,N_14322);
or UO_1606 (O_1606,N_14834,N_14932);
nand UO_1607 (O_1607,N_14728,N_14780);
nor UO_1608 (O_1608,N_14412,N_14524);
nor UO_1609 (O_1609,N_14497,N_14679);
or UO_1610 (O_1610,N_14369,N_14423);
xnor UO_1611 (O_1611,N_14351,N_14671);
and UO_1612 (O_1612,N_14455,N_14682);
nand UO_1613 (O_1613,N_14621,N_14867);
and UO_1614 (O_1614,N_14408,N_14778);
nor UO_1615 (O_1615,N_14985,N_14717);
xnor UO_1616 (O_1616,N_14840,N_14781);
nand UO_1617 (O_1617,N_14938,N_14826);
nand UO_1618 (O_1618,N_14893,N_14551);
or UO_1619 (O_1619,N_14276,N_14685);
nand UO_1620 (O_1620,N_14293,N_14304);
and UO_1621 (O_1621,N_14683,N_14567);
nand UO_1622 (O_1622,N_14806,N_14536);
nand UO_1623 (O_1623,N_14477,N_14955);
xnor UO_1624 (O_1624,N_14751,N_14520);
nand UO_1625 (O_1625,N_14371,N_14659);
or UO_1626 (O_1626,N_14390,N_14779);
nand UO_1627 (O_1627,N_14355,N_14682);
nand UO_1628 (O_1628,N_14782,N_14558);
nor UO_1629 (O_1629,N_14282,N_14975);
nor UO_1630 (O_1630,N_14421,N_14325);
or UO_1631 (O_1631,N_14376,N_14361);
xor UO_1632 (O_1632,N_14319,N_14715);
nand UO_1633 (O_1633,N_14620,N_14252);
xor UO_1634 (O_1634,N_14389,N_14643);
or UO_1635 (O_1635,N_14737,N_14932);
nand UO_1636 (O_1636,N_14734,N_14581);
nor UO_1637 (O_1637,N_14966,N_14331);
xnor UO_1638 (O_1638,N_14466,N_14676);
and UO_1639 (O_1639,N_14351,N_14652);
nor UO_1640 (O_1640,N_14353,N_14913);
xnor UO_1641 (O_1641,N_14792,N_14382);
xor UO_1642 (O_1642,N_14314,N_14915);
xnor UO_1643 (O_1643,N_14900,N_14652);
nor UO_1644 (O_1644,N_14443,N_14873);
and UO_1645 (O_1645,N_14984,N_14327);
nor UO_1646 (O_1646,N_14446,N_14267);
nand UO_1647 (O_1647,N_14812,N_14639);
xor UO_1648 (O_1648,N_14300,N_14466);
nand UO_1649 (O_1649,N_14648,N_14575);
or UO_1650 (O_1650,N_14310,N_14588);
xnor UO_1651 (O_1651,N_14967,N_14989);
xor UO_1652 (O_1652,N_14949,N_14353);
xnor UO_1653 (O_1653,N_14277,N_14667);
and UO_1654 (O_1654,N_14827,N_14867);
nor UO_1655 (O_1655,N_14394,N_14952);
nand UO_1656 (O_1656,N_14447,N_14428);
xnor UO_1657 (O_1657,N_14999,N_14268);
nor UO_1658 (O_1658,N_14358,N_14879);
or UO_1659 (O_1659,N_14950,N_14504);
or UO_1660 (O_1660,N_14801,N_14834);
and UO_1661 (O_1661,N_14976,N_14478);
nand UO_1662 (O_1662,N_14395,N_14636);
and UO_1663 (O_1663,N_14313,N_14827);
nand UO_1664 (O_1664,N_14640,N_14743);
nor UO_1665 (O_1665,N_14604,N_14958);
nand UO_1666 (O_1666,N_14777,N_14833);
and UO_1667 (O_1667,N_14520,N_14874);
xor UO_1668 (O_1668,N_14855,N_14575);
or UO_1669 (O_1669,N_14733,N_14310);
nor UO_1670 (O_1670,N_14631,N_14252);
and UO_1671 (O_1671,N_14565,N_14967);
xnor UO_1672 (O_1672,N_14776,N_14576);
and UO_1673 (O_1673,N_14624,N_14784);
xor UO_1674 (O_1674,N_14444,N_14572);
nand UO_1675 (O_1675,N_14517,N_14828);
nand UO_1676 (O_1676,N_14697,N_14441);
nand UO_1677 (O_1677,N_14606,N_14999);
nor UO_1678 (O_1678,N_14518,N_14893);
or UO_1679 (O_1679,N_14913,N_14858);
nor UO_1680 (O_1680,N_14915,N_14574);
or UO_1681 (O_1681,N_14590,N_14821);
nand UO_1682 (O_1682,N_14386,N_14709);
and UO_1683 (O_1683,N_14697,N_14326);
and UO_1684 (O_1684,N_14846,N_14385);
or UO_1685 (O_1685,N_14684,N_14508);
nor UO_1686 (O_1686,N_14717,N_14388);
nor UO_1687 (O_1687,N_14556,N_14483);
or UO_1688 (O_1688,N_14478,N_14396);
and UO_1689 (O_1689,N_14943,N_14820);
nor UO_1690 (O_1690,N_14384,N_14301);
nor UO_1691 (O_1691,N_14931,N_14892);
nand UO_1692 (O_1692,N_14540,N_14811);
nor UO_1693 (O_1693,N_14964,N_14327);
and UO_1694 (O_1694,N_14429,N_14597);
or UO_1695 (O_1695,N_14718,N_14507);
nor UO_1696 (O_1696,N_14734,N_14297);
nor UO_1697 (O_1697,N_14586,N_14827);
nand UO_1698 (O_1698,N_14915,N_14901);
nor UO_1699 (O_1699,N_14829,N_14882);
or UO_1700 (O_1700,N_14663,N_14390);
or UO_1701 (O_1701,N_14767,N_14692);
xnor UO_1702 (O_1702,N_14812,N_14535);
or UO_1703 (O_1703,N_14655,N_14346);
or UO_1704 (O_1704,N_14863,N_14811);
nor UO_1705 (O_1705,N_14707,N_14381);
nor UO_1706 (O_1706,N_14412,N_14447);
and UO_1707 (O_1707,N_14416,N_14594);
nor UO_1708 (O_1708,N_14472,N_14643);
nand UO_1709 (O_1709,N_14278,N_14696);
and UO_1710 (O_1710,N_14848,N_14629);
xnor UO_1711 (O_1711,N_14658,N_14272);
nor UO_1712 (O_1712,N_14988,N_14951);
xnor UO_1713 (O_1713,N_14472,N_14478);
nand UO_1714 (O_1714,N_14468,N_14584);
or UO_1715 (O_1715,N_14718,N_14423);
or UO_1716 (O_1716,N_14639,N_14542);
nor UO_1717 (O_1717,N_14641,N_14423);
xor UO_1718 (O_1718,N_14599,N_14736);
and UO_1719 (O_1719,N_14992,N_14547);
xnor UO_1720 (O_1720,N_14834,N_14504);
xnor UO_1721 (O_1721,N_14416,N_14504);
nand UO_1722 (O_1722,N_14344,N_14371);
or UO_1723 (O_1723,N_14938,N_14331);
and UO_1724 (O_1724,N_14326,N_14519);
xnor UO_1725 (O_1725,N_14617,N_14989);
nor UO_1726 (O_1726,N_14488,N_14497);
and UO_1727 (O_1727,N_14874,N_14721);
and UO_1728 (O_1728,N_14488,N_14293);
nor UO_1729 (O_1729,N_14754,N_14539);
nand UO_1730 (O_1730,N_14532,N_14870);
xor UO_1731 (O_1731,N_14307,N_14728);
or UO_1732 (O_1732,N_14286,N_14907);
nor UO_1733 (O_1733,N_14260,N_14648);
nor UO_1734 (O_1734,N_14612,N_14905);
nand UO_1735 (O_1735,N_14954,N_14607);
xor UO_1736 (O_1736,N_14749,N_14866);
xnor UO_1737 (O_1737,N_14300,N_14763);
and UO_1738 (O_1738,N_14827,N_14966);
nand UO_1739 (O_1739,N_14477,N_14425);
and UO_1740 (O_1740,N_14849,N_14626);
nor UO_1741 (O_1741,N_14512,N_14295);
xnor UO_1742 (O_1742,N_14409,N_14718);
xnor UO_1743 (O_1743,N_14469,N_14522);
nor UO_1744 (O_1744,N_14857,N_14486);
xnor UO_1745 (O_1745,N_14684,N_14999);
nor UO_1746 (O_1746,N_14833,N_14253);
or UO_1747 (O_1747,N_14620,N_14479);
or UO_1748 (O_1748,N_14776,N_14787);
and UO_1749 (O_1749,N_14473,N_14825);
xnor UO_1750 (O_1750,N_14876,N_14419);
nand UO_1751 (O_1751,N_14624,N_14806);
nand UO_1752 (O_1752,N_14376,N_14991);
nor UO_1753 (O_1753,N_14904,N_14439);
nand UO_1754 (O_1754,N_14933,N_14939);
nand UO_1755 (O_1755,N_14559,N_14562);
or UO_1756 (O_1756,N_14400,N_14974);
nor UO_1757 (O_1757,N_14572,N_14447);
nand UO_1758 (O_1758,N_14717,N_14669);
nand UO_1759 (O_1759,N_14653,N_14634);
or UO_1760 (O_1760,N_14687,N_14555);
nand UO_1761 (O_1761,N_14570,N_14424);
nand UO_1762 (O_1762,N_14513,N_14837);
nand UO_1763 (O_1763,N_14423,N_14720);
and UO_1764 (O_1764,N_14477,N_14892);
or UO_1765 (O_1765,N_14556,N_14456);
or UO_1766 (O_1766,N_14484,N_14776);
nor UO_1767 (O_1767,N_14560,N_14999);
or UO_1768 (O_1768,N_14752,N_14902);
nor UO_1769 (O_1769,N_14782,N_14985);
xor UO_1770 (O_1770,N_14636,N_14321);
xor UO_1771 (O_1771,N_14312,N_14690);
and UO_1772 (O_1772,N_14605,N_14342);
or UO_1773 (O_1773,N_14483,N_14893);
or UO_1774 (O_1774,N_14503,N_14312);
nand UO_1775 (O_1775,N_14811,N_14798);
or UO_1776 (O_1776,N_14421,N_14841);
and UO_1777 (O_1777,N_14273,N_14948);
nor UO_1778 (O_1778,N_14986,N_14267);
nand UO_1779 (O_1779,N_14822,N_14388);
xnor UO_1780 (O_1780,N_14875,N_14718);
and UO_1781 (O_1781,N_14401,N_14674);
or UO_1782 (O_1782,N_14537,N_14912);
nor UO_1783 (O_1783,N_14695,N_14390);
and UO_1784 (O_1784,N_14464,N_14999);
or UO_1785 (O_1785,N_14751,N_14269);
nand UO_1786 (O_1786,N_14322,N_14753);
or UO_1787 (O_1787,N_14307,N_14346);
or UO_1788 (O_1788,N_14585,N_14996);
nor UO_1789 (O_1789,N_14714,N_14860);
nor UO_1790 (O_1790,N_14419,N_14292);
nor UO_1791 (O_1791,N_14918,N_14514);
and UO_1792 (O_1792,N_14991,N_14431);
nor UO_1793 (O_1793,N_14465,N_14797);
and UO_1794 (O_1794,N_14264,N_14894);
or UO_1795 (O_1795,N_14696,N_14612);
xnor UO_1796 (O_1796,N_14368,N_14718);
and UO_1797 (O_1797,N_14982,N_14970);
nand UO_1798 (O_1798,N_14443,N_14385);
and UO_1799 (O_1799,N_14424,N_14730);
nor UO_1800 (O_1800,N_14903,N_14605);
or UO_1801 (O_1801,N_14691,N_14991);
or UO_1802 (O_1802,N_14863,N_14891);
xnor UO_1803 (O_1803,N_14453,N_14591);
or UO_1804 (O_1804,N_14703,N_14376);
or UO_1805 (O_1805,N_14734,N_14675);
xnor UO_1806 (O_1806,N_14874,N_14481);
nand UO_1807 (O_1807,N_14533,N_14422);
nand UO_1808 (O_1808,N_14305,N_14400);
xnor UO_1809 (O_1809,N_14437,N_14491);
nand UO_1810 (O_1810,N_14431,N_14571);
or UO_1811 (O_1811,N_14542,N_14813);
nand UO_1812 (O_1812,N_14351,N_14515);
nand UO_1813 (O_1813,N_14822,N_14856);
nor UO_1814 (O_1814,N_14329,N_14286);
nand UO_1815 (O_1815,N_14789,N_14457);
nand UO_1816 (O_1816,N_14400,N_14962);
or UO_1817 (O_1817,N_14807,N_14893);
nor UO_1818 (O_1818,N_14734,N_14591);
or UO_1819 (O_1819,N_14966,N_14852);
nor UO_1820 (O_1820,N_14455,N_14544);
xor UO_1821 (O_1821,N_14594,N_14332);
nand UO_1822 (O_1822,N_14278,N_14594);
xor UO_1823 (O_1823,N_14991,N_14502);
xor UO_1824 (O_1824,N_14391,N_14629);
xnor UO_1825 (O_1825,N_14613,N_14457);
or UO_1826 (O_1826,N_14890,N_14614);
and UO_1827 (O_1827,N_14975,N_14933);
and UO_1828 (O_1828,N_14919,N_14279);
nand UO_1829 (O_1829,N_14743,N_14879);
and UO_1830 (O_1830,N_14822,N_14998);
nor UO_1831 (O_1831,N_14484,N_14790);
and UO_1832 (O_1832,N_14324,N_14488);
nand UO_1833 (O_1833,N_14308,N_14600);
nand UO_1834 (O_1834,N_14513,N_14269);
or UO_1835 (O_1835,N_14685,N_14911);
or UO_1836 (O_1836,N_14742,N_14298);
xor UO_1837 (O_1837,N_14925,N_14791);
or UO_1838 (O_1838,N_14950,N_14878);
xor UO_1839 (O_1839,N_14888,N_14637);
nand UO_1840 (O_1840,N_14635,N_14926);
nand UO_1841 (O_1841,N_14604,N_14528);
xor UO_1842 (O_1842,N_14729,N_14641);
nand UO_1843 (O_1843,N_14336,N_14297);
or UO_1844 (O_1844,N_14712,N_14678);
and UO_1845 (O_1845,N_14602,N_14908);
nor UO_1846 (O_1846,N_14750,N_14598);
nor UO_1847 (O_1847,N_14934,N_14458);
nand UO_1848 (O_1848,N_14516,N_14655);
and UO_1849 (O_1849,N_14751,N_14490);
nand UO_1850 (O_1850,N_14655,N_14699);
xnor UO_1851 (O_1851,N_14628,N_14966);
and UO_1852 (O_1852,N_14255,N_14972);
and UO_1853 (O_1853,N_14990,N_14309);
nand UO_1854 (O_1854,N_14455,N_14669);
and UO_1855 (O_1855,N_14641,N_14781);
or UO_1856 (O_1856,N_14895,N_14551);
nand UO_1857 (O_1857,N_14272,N_14796);
nor UO_1858 (O_1858,N_14287,N_14545);
nand UO_1859 (O_1859,N_14334,N_14266);
nand UO_1860 (O_1860,N_14462,N_14913);
nand UO_1861 (O_1861,N_14314,N_14355);
nand UO_1862 (O_1862,N_14330,N_14462);
nand UO_1863 (O_1863,N_14901,N_14276);
nand UO_1864 (O_1864,N_14618,N_14259);
nand UO_1865 (O_1865,N_14722,N_14789);
and UO_1866 (O_1866,N_14756,N_14908);
xor UO_1867 (O_1867,N_14620,N_14424);
nor UO_1868 (O_1868,N_14345,N_14698);
or UO_1869 (O_1869,N_14373,N_14330);
or UO_1870 (O_1870,N_14712,N_14682);
nand UO_1871 (O_1871,N_14932,N_14257);
nor UO_1872 (O_1872,N_14336,N_14763);
xor UO_1873 (O_1873,N_14843,N_14661);
xnor UO_1874 (O_1874,N_14281,N_14921);
or UO_1875 (O_1875,N_14613,N_14560);
xnor UO_1876 (O_1876,N_14320,N_14466);
xnor UO_1877 (O_1877,N_14437,N_14273);
nand UO_1878 (O_1878,N_14744,N_14726);
or UO_1879 (O_1879,N_14253,N_14831);
xnor UO_1880 (O_1880,N_14854,N_14747);
and UO_1881 (O_1881,N_14625,N_14916);
nor UO_1882 (O_1882,N_14377,N_14746);
and UO_1883 (O_1883,N_14774,N_14802);
nor UO_1884 (O_1884,N_14432,N_14872);
xnor UO_1885 (O_1885,N_14841,N_14974);
or UO_1886 (O_1886,N_14296,N_14842);
nor UO_1887 (O_1887,N_14367,N_14458);
and UO_1888 (O_1888,N_14783,N_14724);
xor UO_1889 (O_1889,N_14767,N_14472);
and UO_1890 (O_1890,N_14526,N_14891);
xor UO_1891 (O_1891,N_14436,N_14986);
nand UO_1892 (O_1892,N_14540,N_14910);
xnor UO_1893 (O_1893,N_14985,N_14737);
xor UO_1894 (O_1894,N_14382,N_14819);
nand UO_1895 (O_1895,N_14780,N_14377);
nor UO_1896 (O_1896,N_14860,N_14740);
and UO_1897 (O_1897,N_14496,N_14443);
xnor UO_1898 (O_1898,N_14656,N_14353);
nand UO_1899 (O_1899,N_14293,N_14958);
nor UO_1900 (O_1900,N_14794,N_14887);
or UO_1901 (O_1901,N_14542,N_14653);
or UO_1902 (O_1902,N_14998,N_14903);
or UO_1903 (O_1903,N_14838,N_14520);
or UO_1904 (O_1904,N_14373,N_14730);
and UO_1905 (O_1905,N_14762,N_14642);
and UO_1906 (O_1906,N_14269,N_14741);
or UO_1907 (O_1907,N_14761,N_14504);
nor UO_1908 (O_1908,N_14428,N_14373);
nand UO_1909 (O_1909,N_14487,N_14657);
and UO_1910 (O_1910,N_14366,N_14355);
nor UO_1911 (O_1911,N_14797,N_14431);
and UO_1912 (O_1912,N_14452,N_14996);
nand UO_1913 (O_1913,N_14561,N_14892);
nor UO_1914 (O_1914,N_14735,N_14469);
nand UO_1915 (O_1915,N_14963,N_14774);
nor UO_1916 (O_1916,N_14434,N_14923);
nand UO_1917 (O_1917,N_14929,N_14327);
or UO_1918 (O_1918,N_14875,N_14501);
and UO_1919 (O_1919,N_14778,N_14993);
nor UO_1920 (O_1920,N_14624,N_14713);
nor UO_1921 (O_1921,N_14432,N_14710);
and UO_1922 (O_1922,N_14655,N_14685);
and UO_1923 (O_1923,N_14545,N_14819);
xor UO_1924 (O_1924,N_14369,N_14424);
and UO_1925 (O_1925,N_14799,N_14587);
xnor UO_1926 (O_1926,N_14816,N_14990);
nor UO_1927 (O_1927,N_14327,N_14595);
nor UO_1928 (O_1928,N_14935,N_14397);
nor UO_1929 (O_1929,N_14313,N_14870);
nor UO_1930 (O_1930,N_14641,N_14552);
nand UO_1931 (O_1931,N_14852,N_14513);
xor UO_1932 (O_1932,N_14655,N_14794);
nor UO_1933 (O_1933,N_14525,N_14812);
and UO_1934 (O_1934,N_14487,N_14769);
nor UO_1935 (O_1935,N_14525,N_14762);
and UO_1936 (O_1936,N_14404,N_14789);
and UO_1937 (O_1937,N_14725,N_14941);
and UO_1938 (O_1938,N_14863,N_14488);
and UO_1939 (O_1939,N_14310,N_14829);
xnor UO_1940 (O_1940,N_14947,N_14915);
nand UO_1941 (O_1941,N_14982,N_14555);
nor UO_1942 (O_1942,N_14931,N_14633);
nor UO_1943 (O_1943,N_14984,N_14413);
or UO_1944 (O_1944,N_14770,N_14339);
xor UO_1945 (O_1945,N_14666,N_14809);
nor UO_1946 (O_1946,N_14533,N_14958);
nand UO_1947 (O_1947,N_14761,N_14889);
nor UO_1948 (O_1948,N_14627,N_14894);
xor UO_1949 (O_1949,N_14604,N_14410);
xnor UO_1950 (O_1950,N_14835,N_14774);
or UO_1951 (O_1951,N_14970,N_14667);
and UO_1952 (O_1952,N_14453,N_14363);
and UO_1953 (O_1953,N_14321,N_14474);
or UO_1954 (O_1954,N_14892,N_14525);
nand UO_1955 (O_1955,N_14618,N_14390);
nand UO_1956 (O_1956,N_14604,N_14380);
and UO_1957 (O_1957,N_14303,N_14617);
xnor UO_1958 (O_1958,N_14332,N_14580);
xnor UO_1959 (O_1959,N_14435,N_14776);
nand UO_1960 (O_1960,N_14478,N_14995);
nand UO_1961 (O_1961,N_14582,N_14765);
xor UO_1962 (O_1962,N_14670,N_14840);
or UO_1963 (O_1963,N_14896,N_14357);
xor UO_1964 (O_1964,N_14686,N_14618);
and UO_1965 (O_1965,N_14423,N_14972);
nor UO_1966 (O_1966,N_14839,N_14999);
xnor UO_1967 (O_1967,N_14813,N_14864);
nand UO_1968 (O_1968,N_14463,N_14299);
nor UO_1969 (O_1969,N_14549,N_14376);
and UO_1970 (O_1970,N_14973,N_14461);
xnor UO_1971 (O_1971,N_14543,N_14487);
nor UO_1972 (O_1972,N_14821,N_14866);
nor UO_1973 (O_1973,N_14964,N_14548);
nor UO_1974 (O_1974,N_14854,N_14623);
xnor UO_1975 (O_1975,N_14265,N_14887);
nand UO_1976 (O_1976,N_14406,N_14896);
nand UO_1977 (O_1977,N_14880,N_14830);
and UO_1978 (O_1978,N_14363,N_14924);
nor UO_1979 (O_1979,N_14352,N_14512);
nand UO_1980 (O_1980,N_14648,N_14337);
xnor UO_1981 (O_1981,N_14667,N_14292);
nand UO_1982 (O_1982,N_14935,N_14430);
or UO_1983 (O_1983,N_14908,N_14842);
and UO_1984 (O_1984,N_14948,N_14858);
nor UO_1985 (O_1985,N_14893,N_14722);
xor UO_1986 (O_1986,N_14494,N_14328);
xnor UO_1987 (O_1987,N_14814,N_14391);
and UO_1988 (O_1988,N_14992,N_14696);
nor UO_1989 (O_1989,N_14640,N_14633);
and UO_1990 (O_1990,N_14456,N_14460);
xor UO_1991 (O_1991,N_14631,N_14493);
xor UO_1992 (O_1992,N_14261,N_14273);
xnor UO_1993 (O_1993,N_14752,N_14699);
or UO_1994 (O_1994,N_14438,N_14750);
nand UO_1995 (O_1995,N_14721,N_14676);
and UO_1996 (O_1996,N_14309,N_14513);
or UO_1997 (O_1997,N_14254,N_14406);
or UO_1998 (O_1998,N_14331,N_14353);
xnor UO_1999 (O_1999,N_14779,N_14617);
endmodule