module basic_2000_20000_2500_10_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_125,In_692);
xnor U1 (N_1,In_924,In_269);
nor U2 (N_2,In_528,In_214);
or U3 (N_3,In_1594,In_192);
nand U4 (N_4,In_1620,In_1913);
and U5 (N_5,In_249,In_978);
nor U6 (N_6,In_1250,In_1918);
xor U7 (N_7,In_478,In_1329);
nand U8 (N_8,In_1364,In_356);
or U9 (N_9,In_493,In_1551);
or U10 (N_10,In_1919,In_392);
nand U11 (N_11,In_1007,In_3);
or U12 (N_12,In_1129,In_1998);
and U13 (N_13,In_1018,In_1704);
and U14 (N_14,In_1385,In_626);
and U15 (N_15,In_284,In_487);
nor U16 (N_16,In_22,In_1033);
nand U17 (N_17,In_1167,In_762);
xnor U18 (N_18,In_189,In_1895);
nand U19 (N_19,In_1133,In_1082);
and U20 (N_20,In_530,In_208);
and U21 (N_21,In_275,In_691);
xor U22 (N_22,In_599,In_1684);
nor U23 (N_23,In_1685,In_1773);
xnor U24 (N_24,In_291,In_1572);
nand U25 (N_25,In_713,In_1553);
nor U26 (N_26,In_1219,In_1556);
nor U27 (N_27,In_245,In_1215);
xnor U28 (N_28,In_1228,In_1526);
nor U29 (N_29,In_93,In_130);
xnor U30 (N_30,In_974,In_1387);
nand U31 (N_31,In_748,In_433);
or U32 (N_32,In_1862,In_678);
or U33 (N_33,In_1593,In_1139);
or U34 (N_34,In_1410,In_413);
xnor U35 (N_35,In_1755,In_1398);
or U36 (N_36,In_8,In_285);
nand U37 (N_37,In_1058,In_1430);
nand U38 (N_38,In_467,In_496);
nor U39 (N_39,In_1798,In_188);
or U40 (N_40,In_1957,In_564);
nand U41 (N_41,In_650,In_602);
xor U42 (N_42,In_1948,In_568);
nand U43 (N_43,In_701,In_64);
and U44 (N_44,In_1667,In_169);
xor U45 (N_45,In_797,In_442);
and U46 (N_46,In_359,In_1887);
and U47 (N_47,In_1605,In_1561);
nor U48 (N_48,In_930,In_1305);
nor U49 (N_49,In_1189,In_981);
xnor U50 (N_50,In_1166,In_913);
or U51 (N_51,In_1448,In_1739);
and U52 (N_52,In_432,In_1666);
and U53 (N_53,In_1825,In_810);
or U54 (N_54,In_1193,In_1296);
xnor U55 (N_55,In_771,In_1021);
and U56 (N_56,In_1315,In_733);
nand U57 (N_57,In_1187,In_1506);
or U58 (N_58,In_166,In_314);
nor U59 (N_59,In_332,In_1105);
xnor U60 (N_60,In_997,In_1263);
xnor U61 (N_61,In_1920,In_440);
or U62 (N_62,In_301,In_1629);
nand U63 (N_63,In_403,In_1113);
and U64 (N_64,In_705,In_1603);
nand U65 (N_65,In_1851,In_1042);
nand U66 (N_66,In_1837,In_1447);
nand U67 (N_67,In_139,In_99);
nor U68 (N_68,In_644,In_1159);
xor U69 (N_69,In_1806,In_78);
and U70 (N_70,In_992,In_1345);
nand U71 (N_71,In_9,In_224);
nand U72 (N_72,In_370,In_711);
and U73 (N_73,In_1431,In_679);
nor U74 (N_74,In_1214,In_374);
nand U75 (N_75,In_182,In_1262);
xnor U76 (N_76,In_1707,In_829);
xor U77 (N_77,In_241,In_1403);
or U78 (N_78,In_1970,In_1184);
or U79 (N_79,In_1255,In_895);
and U80 (N_80,In_1376,In_1743);
xnor U81 (N_81,In_369,In_1468);
and U82 (N_82,In_686,In_546);
or U83 (N_83,In_460,In_1314);
nand U84 (N_84,In_1911,In_734);
or U85 (N_85,In_1891,In_943);
nor U86 (N_86,In_871,In_1952);
xnor U87 (N_87,In_716,In_1753);
or U88 (N_88,In_1587,In_71);
or U89 (N_89,In_240,In_647);
nand U90 (N_90,In_1404,In_97);
or U91 (N_91,In_915,In_671);
nand U92 (N_92,In_972,In_983);
and U93 (N_93,In_1897,In_1731);
xnor U94 (N_94,In_1246,In_796);
and U95 (N_95,In_280,In_1791);
xnor U96 (N_96,In_133,In_820);
and U97 (N_97,In_838,In_1446);
nor U98 (N_98,In_210,In_1053);
nand U99 (N_99,In_295,In_1232);
and U100 (N_100,In_1287,In_1720);
or U101 (N_101,In_819,In_1599);
nor U102 (N_102,In_1537,In_1118);
nor U103 (N_103,In_1420,In_1273);
xnor U104 (N_104,In_1521,In_916);
and U105 (N_105,In_1198,In_770);
and U106 (N_106,In_1630,In_890);
nand U107 (N_107,In_54,In_638);
and U108 (N_108,In_1585,In_402);
and U109 (N_109,In_150,In_1792);
xnor U110 (N_110,In_1407,In_1758);
xor U111 (N_111,In_1930,In_1369);
or U112 (N_112,In_357,In_1014);
and U113 (N_113,In_1213,In_62);
or U114 (N_114,In_1483,In_1516);
or U115 (N_115,In_126,In_1396);
and U116 (N_116,In_548,In_94);
xor U117 (N_117,In_324,In_1567);
nor U118 (N_118,In_724,In_1402);
nand U119 (N_119,In_756,In_1683);
xor U120 (N_120,In_1182,In_72);
and U121 (N_121,In_1705,In_289);
xnor U122 (N_122,In_929,In_113);
nor U123 (N_123,In_959,In_1881);
nor U124 (N_124,In_1669,In_798);
xnor U125 (N_125,In_1759,In_1375);
or U126 (N_126,In_216,In_1856);
and U127 (N_127,In_1980,In_793);
or U128 (N_128,In_761,In_254);
or U129 (N_129,In_988,In_366);
nor U130 (N_130,In_1966,In_1915);
nand U131 (N_131,In_1392,In_256);
and U132 (N_132,In_23,In_1833);
xnor U133 (N_133,In_1997,In_500);
xor U134 (N_134,In_1691,In_1717);
xnor U135 (N_135,In_1765,In_428);
xor U136 (N_136,In_937,In_164);
nor U137 (N_137,In_1672,In_741);
and U138 (N_138,In_754,In_140);
and U139 (N_139,In_555,In_1575);
or U140 (N_140,In_342,In_1342);
or U141 (N_141,In_1963,In_714);
and U142 (N_142,In_1044,In_887);
nor U143 (N_143,In_156,In_667);
nor U144 (N_144,In_1443,In_1240);
nor U145 (N_145,In_1648,In_654);
xnor U146 (N_146,In_1508,In_1172);
nor U147 (N_147,In_1015,In_207);
nand U148 (N_148,In_352,In_129);
and U149 (N_149,In_1584,In_1381);
xor U150 (N_150,In_149,In_196);
nor U151 (N_151,In_187,In_446);
nor U152 (N_152,In_1769,In_826);
or U153 (N_153,In_186,In_320);
xor U154 (N_154,In_1972,In_731);
nor U155 (N_155,In_749,In_185);
and U156 (N_156,In_6,In_1);
and U157 (N_157,In_326,In_950);
nor U158 (N_158,In_1652,In_1241);
and U159 (N_159,In_380,In_1680);
and U160 (N_160,In_1503,In_1030);
xnor U161 (N_161,In_1278,In_1094);
nor U162 (N_162,In_1389,In_1126);
nand U163 (N_163,In_600,In_1065);
nand U164 (N_164,In_98,In_376);
xnor U165 (N_165,In_1686,In_1211);
nor U166 (N_166,In_814,In_1764);
and U167 (N_167,In_1550,In_1912);
or U168 (N_168,In_1110,In_582);
and U169 (N_169,In_775,In_283);
and U170 (N_170,In_1128,In_1442);
and U171 (N_171,In_1380,In_1436);
or U172 (N_172,In_371,In_1892);
and U173 (N_173,In_390,In_1009);
and U174 (N_174,In_1327,In_1054);
xor U175 (N_175,In_1454,In_1064);
and U176 (N_176,In_253,In_1300);
nor U177 (N_177,In_844,In_355);
nand U178 (N_178,In_1037,In_1627);
or U179 (N_179,In_1861,In_1868);
xnor U180 (N_180,In_416,In_538);
xnor U181 (N_181,In_37,In_1253);
and U182 (N_182,In_1502,In_1543);
and U183 (N_183,In_795,In_891);
and U184 (N_184,In_1874,In_957);
nor U185 (N_185,In_222,In_1291);
nand U186 (N_186,In_459,In_411);
nor U187 (N_187,In_853,In_1153);
xor U188 (N_188,In_1060,In_1390);
or U189 (N_189,In_539,In_89);
xor U190 (N_190,In_1467,In_1086);
or U191 (N_191,In_281,In_1875);
or U192 (N_192,In_302,In_1069);
xor U193 (N_193,In_1104,In_1170);
nor U194 (N_194,In_1419,In_1738);
nand U195 (N_195,In_1274,In_1077);
or U196 (N_196,In_608,In_614);
xor U197 (N_197,In_1510,In_1025);
xor U198 (N_198,In_778,In_1746);
nand U199 (N_199,In_57,In_1281);
nand U200 (N_200,In_1247,In_1840);
nand U201 (N_201,In_1905,In_250);
xor U202 (N_202,In_938,In_1961);
nand U203 (N_203,In_1304,In_1264);
or U204 (N_204,In_1333,In_310);
nand U205 (N_205,In_1610,In_162);
nand U206 (N_206,In_1531,In_1761);
nor U207 (N_207,In_469,In_1100);
and U208 (N_208,In_1034,In_1774);
xor U209 (N_209,In_1070,In_334);
nand U210 (N_210,In_1067,In_958);
and U211 (N_211,In_1511,In_237);
nand U212 (N_212,In_225,In_272);
and U213 (N_213,In_1549,In_1618);
or U214 (N_214,In_1878,In_736);
nand U215 (N_215,In_1735,In_867);
or U216 (N_216,In_1899,In_846);
nor U217 (N_217,In_1482,In_1546);
and U218 (N_218,In_552,In_1950);
or U219 (N_219,In_521,In_1394);
xor U220 (N_220,In_834,In_1179);
nor U221 (N_221,In_1600,In_365);
or U222 (N_222,In_970,In_455);
nand U223 (N_223,In_1455,In_1309);
nor U224 (N_224,In_1284,In_1867);
or U225 (N_225,In_1324,In_852);
xor U226 (N_226,In_660,In_409);
and U227 (N_227,In_1290,In_1665);
xnor U228 (N_228,In_55,In_750);
or U229 (N_229,In_475,In_995);
and U230 (N_230,In_677,In_809);
nand U231 (N_231,In_1196,In_889);
nand U232 (N_232,In_1485,In_111);
nor U233 (N_233,In_1288,In_952);
nand U234 (N_234,In_1202,In_885);
nor U235 (N_235,In_1120,In_835);
nand U236 (N_236,In_1357,In_311);
nand U237 (N_237,In_699,In_1591);
and U238 (N_238,In_1525,In_554);
xnor U239 (N_239,In_1766,In_526);
and U240 (N_240,In_451,In_1882);
nand U241 (N_241,In_1953,In_1993);
xnor U242 (N_242,In_791,In_1257);
nor U243 (N_243,In_980,In_823);
and U244 (N_244,In_1098,In_1124);
nand U245 (N_245,In_1377,In_627);
or U246 (N_246,In_1566,In_640);
and U247 (N_247,In_5,In_1415);
xnor U248 (N_248,In_789,In_218);
nand U249 (N_249,In_1116,In_1624);
nand U250 (N_250,In_1902,In_518);
xor U251 (N_251,In_1180,In_193);
nor U252 (N_252,In_1023,In_1645);
and U253 (N_253,In_154,In_1076);
xnor U254 (N_254,In_1465,In_1272);
or U255 (N_255,In_238,In_1805);
and U256 (N_256,In_1718,In_1496);
nand U257 (N_257,In_934,In_1019);
nand U258 (N_258,In_1353,In_986);
nor U259 (N_259,In_309,In_1013);
nand U260 (N_260,In_1307,In_1249);
nand U261 (N_261,In_1744,In_529);
or U262 (N_262,In_148,In_109);
nand U263 (N_263,In_1760,In_361);
nor U264 (N_264,In_1035,In_211);
or U265 (N_265,In_523,In_41);
or U266 (N_266,In_1000,In_825);
xor U267 (N_267,In_739,In_923);
nor U268 (N_268,In_1108,In_124);
and U269 (N_269,In_421,In_1985);
xor U270 (N_270,In_1138,In_684);
nand U271 (N_271,In_1340,In_1716);
nor U272 (N_272,In_143,In_1971);
and U273 (N_273,In_197,In_501);
xnor U274 (N_274,In_486,In_118);
or U275 (N_275,In_1177,In_382);
xor U276 (N_276,In_345,In_1568);
xor U277 (N_277,In_1992,In_652);
or U278 (N_278,In_1259,In_1835);
xor U279 (N_279,In_690,In_1781);
nor U280 (N_280,In_1740,In_1382);
nor U281 (N_281,In_20,In_1414);
nand U282 (N_282,In_1337,In_525);
nand U283 (N_283,In_120,In_1767);
and U284 (N_284,In_1038,In_709);
and U285 (N_285,In_1097,In_40);
nor U286 (N_286,In_803,In_175);
nor U287 (N_287,In_674,In_1849);
xnor U288 (N_288,In_1909,In_848);
or U289 (N_289,In_1474,In_1723);
nand U290 (N_290,In_481,In_1800);
nor U291 (N_291,In_354,In_704);
xnor U292 (N_292,In_1268,In_331);
and U293 (N_293,In_1475,In_1432);
nor U294 (N_294,In_136,In_1884);
or U295 (N_295,In_611,In_1859);
nor U296 (N_296,In_1636,In_1662);
nor U297 (N_297,In_1362,In_742);
and U298 (N_298,In_948,In_1649);
nor U299 (N_299,In_1050,In_1960);
and U300 (N_300,In_651,In_1444);
nor U301 (N_301,In_910,In_1690);
nor U302 (N_302,In_772,In_812);
xnor U303 (N_303,In_1302,In_782);
nor U304 (N_304,In_753,In_1224);
nor U305 (N_305,In_1839,In_917);
or U306 (N_306,In_594,In_1320);
nor U307 (N_307,In_875,In_1200);
nor U308 (N_308,In_1005,In_1140);
and U309 (N_309,In_570,In_788);
nor U310 (N_310,In_708,In_1227);
nor U311 (N_311,In_512,In_381);
xor U312 (N_312,In_1999,In_505);
nor U313 (N_313,In_134,In_1338);
and U314 (N_314,In_595,In_1698);
nor U315 (N_315,In_1826,In_747);
nor U316 (N_316,In_404,In_1354);
or U317 (N_317,In_520,In_360);
and U318 (N_318,In_183,In_96);
nand U319 (N_319,In_776,In_944);
nand U320 (N_320,In_303,In_1079);
xor U321 (N_321,In_517,In_1470);
xnor U322 (N_322,In_1577,In_779);
or U323 (N_323,In_998,In_604);
or U324 (N_324,In_473,In_1433);
xor U325 (N_325,In_1570,In_1987);
nor U326 (N_326,In_964,In_1545);
or U327 (N_327,In_1907,In_1427);
xnor U328 (N_328,In_1087,In_1812);
xnor U329 (N_329,In_397,In_1528);
xor U330 (N_330,In_1039,In_883);
xor U331 (N_331,In_1693,In_1727);
nor U332 (N_332,In_804,In_45);
nor U333 (N_333,In_1583,In_760);
xnor U334 (N_334,In_1313,In_1519);
and U335 (N_335,In_1679,In_1445);
xor U336 (N_336,In_418,In_840);
xnor U337 (N_337,In_1544,In_907);
or U338 (N_338,In_1702,In_1940);
or U339 (N_339,In_230,In_991);
or U340 (N_340,In_854,In_398);
and U341 (N_341,In_1619,In_956);
xnor U342 (N_342,In_1956,In_1201);
or U343 (N_343,In_414,In_1609);
nor U344 (N_344,In_1616,In_329);
nor U345 (N_345,In_464,In_1135);
nand U346 (N_346,In_48,In_706);
nand U347 (N_347,In_252,In_267);
xnor U348 (N_348,In_79,In_902);
xor U349 (N_349,In_1106,In_1051);
nor U350 (N_350,In_1713,In_339);
nor U351 (N_351,In_1756,In_259);
or U352 (N_352,In_639,In_897);
or U353 (N_353,In_472,In_1834);
or U354 (N_354,In_653,In_1844);
or U355 (N_355,In_220,In_1994);
nor U356 (N_356,In_645,In_177);
nor U357 (N_357,In_349,In_1238);
or U358 (N_358,In_181,In_1355);
and U359 (N_359,In_247,In_86);
nand U360 (N_360,In_168,In_1843);
xor U361 (N_361,In_1149,In_680);
and U362 (N_362,In_458,In_591);
nor U363 (N_363,In_1171,In_1936);
or U364 (N_364,In_1046,In_908);
or U365 (N_365,In_946,In_817);
and U366 (N_366,In_634,In_617);
nor U367 (N_367,In_1922,In_180);
nor U368 (N_368,In_1697,In_971);
and U369 (N_369,In_687,In_531);
or U370 (N_370,In_1811,In_1931);
nor U371 (N_371,In_1157,In_1192);
nand U372 (N_372,In_1778,In_147);
nand U373 (N_373,In_822,In_1237);
nor U374 (N_374,In_1977,In_511);
or U375 (N_375,In_1770,In_426);
xor U376 (N_376,In_63,In_1933);
nor U377 (N_377,In_573,In_842);
and U378 (N_378,In_1661,In_491);
xnor U379 (N_379,In_1429,In_1654);
and U380 (N_380,In_1638,In_1775);
nor U381 (N_381,In_1395,In_1406);
or U382 (N_382,In_1117,In_1797);
nand U383 (N_383,In_315,In_21);
xor U384 (N_384,In_274,In_1486);
or U385 (N_385,In_1156,In_341);
or U386 (N_386,In_1162,In_781);
and U387 (N_387,In_1742,In_1949);
or U388 (N_388,In_1248,In_1823);
nor U389 (N_389,In_178,In_81);
nand U390 (N_390,In_430,In_1974);
nor U391 (N_391,In_194,In_1356);
and U392 (N_392,In_1601,In_1372);
and U393 (N_393,In_1500,In_1493);
nand U394 (N_394,In_15,In_1924);
nand U395 (N_395,In_450,In_88);
and U396 (N_396,In_1988,In_427);
nor U397 (N_397,In_1195,In_1900);
or U398 (N_398,In_277,In_758);
nor U399 (N_399,In_598,In_318);
and U400 (N_400,In_312,In_123);
nor U401 (N_401,In_1423,In_1440);
nand U402 (N_402,In_1650,In_802);
and U403 (N_403,In_642,In_1130);
or U404 (N_404,In_1242,In_1802);
or U405 (N_405,In_429,In_1150);
nand U406 (N_406,In_1653,In_1325);
nor U407 (N_407,In_1726,In_1488);
nor U408 (N_408,In_1499,In_921);
nand U409 (N_409,In_1318,In_1794);
xnor U410 (N_410,In_1265,In_1532);
and U411 (N_411,In_191,In_1628);
nor U412 (N_412,In_1724,In_489);
xor U413 (N_413,In_265,In_1548);
nand U414 (N_414,In_832,In_461);
and U415 (N_415,In_1206,In_290);
nand U416 (N_416,In_612,In_1854);
nor U417 (N_417,In_1494,In_386);
or U418 (N_418,In_1613,In_202);
xor U419 (N_419,In_135,In_410);
or U420 (N_420,In_547,In_358);
and U421 (N_421,In_939,In_1473);
and U422 (N_422,In_987,In_1449);
and U423 (N_423,In_1850,In_1643);
xnor U424 (N_424,In_394,In_85);
or U425 (N_425,In_813,In_715);
nor U426 (N_426,In_227,In_389);
nand U427 (N_427,In_1938,In_1010);
or U428 (N_428,In_1663,In_1527);
xor U429 (N_429,In_435,In_673);
xor U430 (N_430,In_495,In_1497);
nor U431 (N_431,In_170,In_933);
nand U432 (N_432,In_1687,In_1675);
or U433 (N_433,In_1815,In_82);
nand U434 (N_434,In_593,In_1975);
xnor U435 (N_435,In_534,In_84);
or U436 (N_436,In_1730,In_828);
and U437 (N_437,In_1973,In_385);
and U438 (N_438,In_1322,In_69);
nor U439 (N_439,In_1535,In_730);
xnor U440 (N_440,In_605,In_90);
and U441 (N_441,In_1022,In_1478);
or U442 (N_442,In_738,In_1459);
nor U443 (N_443,In_1490,In_966);
nor U444 (N_444,In_827,In_1602);
nor U445 (N_445,In_557,In_533);
nor U446 (N_446,In_1877,In_50);
nor U447 (N_447,In_1383,In_1990);
xnor U448 (N_448,In_1072,In_764);
nor U449 (N_449,In_655,In_1799);
nand U450 (N_450,In_378,In_1217);
or U451 (N_451,In_1016,In_551);
xnor U452 (N_452,In_367,In_1347);
and U453 (N_453,In_1306,In_1146);
or U454 (N_454,In_836,In_866);
and U455 (N_455,In_1359,In_438);
xor U456 (N_456,In_346,In_384);
and U457 (N_457,In_831,In_886);
nand U458 (N_458,In_117,In_17);
nor U459 (N_459,In_592,In_755);
nor U460 (N_460,In_1695,In_1308);
xor U461 (N_461,In_1608,In_1539);
and U462 (N_462,In_1463,In_1703);
or U463 (N_463,In_1185,In_1344);
xor U464 (N_464,In_1639,In_242);
and U465 (N_465,In_38,In_223);
and U466 (N_466,In_833,In_1123);
nor U467 (N_467,In_1209,In_1457);
and U468 (N_468,In_1137,In_879);
or U469 (N_469,In_1512,In_260);
and U470 (N_470,In_1323,In_586);
and U471 (N_471,In_251,In_1757);
xnor U472 (N_472,In_1745,In_1777);
nand U473 (N_473,In_919,In_115);
xnor U474 (N_474,In_783,In_279);
nand U475 (N_475,In_1635,In_1441);
and U476 (N_476,In_1080,In_1084);
nand U477 (N_477,In_1981,In_190);
or U478 (N_478,In_1131,In_1651);
xor U479 (N_479,In_1607,In_587);
and U480 (N_480,In_693,In_373);
and U481 (N_481,In_1634,In_1787);
and U482 (N_482,In_176,In_1173);
nand U483 (N_483,In_1728,In_712);
and U484 (N_484,In_851,In_728);
nand U485 (N_485,In_843,In_597);
xor U486 (N_486,In_172,In_1754);
xor U487 (N_487,In_463,In_1890);
xnor U488 (N_488,In_683,In_1095);
or U489 (N_489,In_928,In_1563);
nand U490 (N_490,In_1222,In_255);
and U491 (N_491,In_1828,In_273);
nand U492 (N_492,In_266,In_1929);
and U493 (N_493,In_492,In_1373);
nor U494 (N_494,In_559,In_1292);
or U495 (N_495,In_1295,In_1412);
nand U496 (N_496,In_982,In_1750);
and U497 (N_497,In_1709,In_296);
nand U498 (N_498,In_337,In_569);
or U499 (N_499,In_1578,In_839);
xor U500 (N_500,In_258,In_681);
nor U501 (N_501,In_906,In_572);
xor U502 (N_502,In_575,In_1996);
and U503 (N_503,In_110,In_695);
nand U504 (N_504,In_1059,In_226);
nor U505 (N_505,In_1071,In_863);
or U506 (N_506,In_1391,In_861);
nor U507 (N_507,In_646,In_1831);
and U508 (N_508,In_221,In_1942);
nor U509 (N_509,In_1784,In_590);
or U510 (N_510,In_1925,In_399);
xnor U511 (N_511,In_484,In_1043);
and U512 (N_512,In_1633,In_36);
xnor U513 (N_513,In_1564,In_567);
or U514 (N_514,In_1838,In_894);
nor U515 (N_515,In_1813,In_696);
or U516 (N_516,In_1484,In_13);
or U517 (N_517,In_1885,In_664);
nand U518 (N_518,In_16,In_960);
or U519 (N_519,In_514,In_616);
nand U520 (N_520,In_583,In_74);
and U521 (N_521,In_544,In_967);
xor U522 (N_522,In_278,In_1655);
or U523 (N_523,In_720,In_408);
nand U524 (N_524,In_316,In_794);
and U525 (N_525,In_707,In_1181);
nor U526 (N_526,In_522,In_1596);
nor U527 (N_527,In_1870,In_1085);
or U528 (N_528,In_619,In_532);
and U529 (N_529,In_1518,In_236);
nor U530 (N_530,In_1562,In_119);
nand U531 (N_531,In_574,In_1888);
nand U532 (N_532,In_1462,In_1533);
xor U533 (N_533,In_1509,In_1083);
or U534 (N_534,In_643,In_1221);
xnor U535 (N_535,In_976,In_1771);
and U536 (N_536,In_56,In_424);
nor U537 (N_537,In_1943,In_206);
nor U538 (N_538,In_669,In_1747);
or U539 (N_539,In_66,In_718);
or U540 (N_540,In_1598,In_1408);
and U541 (N_541,In_1959,In_784);
xnor U542 (N_542,In_479,In_1592);
nor U543 (N_543,In_1405,In_401);
nand U544 (N_544,In_1965,In_1491);
or U545 (N_545,In_1115,In_445);
or U546 (N_546,In_877,In_1132);
or U547 (N_547,In_884,In_1986);
and U548 (N_548,In_502,In_566);
nand U549 (N_549,In_51,In_1589);
and U550 (N_550,In_1254,In_179);
nand U551 (N_551,In_1542,In_945);
nor U552 (N_552,In_138,In_1848);
nor U553 (N_553,In_1872,In_1689);
xnor U554 (N_554,In_423,In_1623);
and U555 (N_555,In_1223,In_1896);
nor U556 (N_556,In_899,In_697);
nand U557 (N_557,In_388,In_1910);
xnor U558 (N_558,In_1810,In_1821);
and U559 (N_559,In_580,In_1939);
nand U560 (N_560,In_1658,In_1194);
and U561 (N_561,In_1260,In_1804);
nand U562 (N_562,In_792,In_1164);
and U563 (N_563,In_1571,In_1269);
xnor U564 (N_564,In_1341,In_335);
and U565 (N_565,In_1903,In_444);
nor U566 (N_566,In_1335,In_308);
or U567 (N_567,In_1277,In_299);
nor U568 (N_568,In_1934,In_1515);
xor U569 (N_569,In_1152,In_1579);
and U570 (N_570,In_321,In_122);
nor U571 (N_571,In_203,In_816);
nand U572 (N_572,In_1155,In_656);
nand U573 (N_573,In_200,In_1109);
nor U574 (N_574,In_92,In_1646);
and U575 (N_575,In_1091,In_918);
nor U576 (N_576,In_26,In_1946);
nand U577 (N_577,In_287,In_1458);
and U578 (N_578,In_1004,In_327);
or U579 (N_579,In_726,In_1671);
xor U580 (N_580,In_1954,In_1816);
or U581 (N_581,In_1147,In_83);
xor U582 (N_582,In_785,In_722);
nand U583 (N_583,In_878,In_1203);
nand U584 (N_584,In_1151,In_286);
nand U585 (N_585,In_173,In_698);
nor U586 (N_586,In_1827,In_1245);
xnor U587 (N_587,In_1074,In_1175);
xnor U588 (N_588,In_465,In_1006);
nor U589 (N_589,In_67,In_541);
nor U590 (N_590,In_1947,In_1513);
or U591 (N_591,In_1066,In_1029);
nand U592 (N_592,In_1048,In_1699);
or U593 (N_593,In_11,In_994);
nor U594 (N_594,In_1906,In_1197);
nor U595 (N_595,In_127,In_396);
nand U596 (N_596,In_1801,In_212);
or U597 (N_597,In_106,In_1845);
or U598 (N_598,In_1536,In_1090);
or U599 (N_599,In_364,In_305);
nand U600 (N_600,In_1439,In_1421);
xor U601 (N_601,In_563,In_1719);
nor U602 (N_602,In_558,In_1673);
or U603 (N_603,In_1127,In_1178);
nor U604 (N_604,In_131,In_18);
and U605 (N_605,In_700,In_1559);
and U606 (N_606,In_205,In_400);
nor U607 (N_607,In_233,In_14);
or U608 (N_608,In_1783,In_1818);
and U609 (N_609,In_1002,In_898);
or U610 (N_610,In_19,In_1514);
nand U611 (N_611,In_262,In_1088);
or U612 (N_612,In_1310,In_1472);
nand U613 (N_613,In_1154,In_1425);
nand U614 (N_614,In_1207,In_927);
nand U615 (N_615,In_1384,In_1822);
nor U616 (N_616,In_685,In_1122);
nand U617 (N_617,In_790,In_1889);
nand U618 (N_618,In_1779,In_1852);
and U619 (N_619,In_282,In_1976);
nand U620 (N_620,In_1158,In_33);
or U621 (N_621,In_49,In_271);
or U622 (N_622,In_1343,In_1893);
and U623 (N_623,In_1860,In_618);
and U624 (N_624,In_1012,In_632);
xnor U625 (N_625,In_1297,In_1517);
nand U626 (N_626,In_859,In_1932);
nand U627 (N_627,In_1908,In_1371);
xor U628 (N_628,In_1772,In_1230);
xnor U629 (N_629,In_101,In_1437);
nand U630 (N_630,In_1869,In_1729);
nor U631 (N_631,In_860,In_537);
nor U632 (N_632,In_1901,In_856);
and U633 (N_633,In_719,In_1275);
xor U634 (N_634,In_43,In_1637);
nor U635 (N_635,In_1400,In_1937);
nor U636 (N_636,In_1092,In_904);
xor U637 (N_637,In_1041,In_1858);
nor U638 (N_638,In_613,In_1417);
or U639 (N_639,In_1363,In_454);
and U640 (N_640,In_1857,In_1749);
nor U641 (N_641,In_457,In_25);
or U642 (N_642,In_1317,In_322);
nor U643 (N_643,In_830,In_1715);
xnor U644 (N_644,In_1967,In_1817);
xor U645 (N_645,In_1428,In_576);
nor U646 (N_646,In_556,In_805);
or U647 (N_647,In_1205,In_1656);
nor U648 (N_648,In_606,In_1422);
or U649 (N_649,In_1964,In_1968);
or U650 (N_650,In_1040,In_657);
nand U651 (N_651,In_737,In_1780);
or U652 (N_652,In_243,In_1886);
and U653 (N_653,In_1565,In_163);
nand U654 (N_654,In_1028,In_434);
nand U655 (N_655,In_1045,In_519);
or U656 (N_656,In_1134,In_1688);
nand U657 (N_657,In_1557,In_1732);
nand U658 (N_658,In_1547,In_1081);
nor U659 (N_659,In_849,In_1597);
or U660 (N_660,In_91,In_1504);
nor U661 (N_661,In_622,In_1832);
xnor U662 (N_662,In_1752,In_694);
and U663 (N_663,In_68,In_1216);
and U664 (N_664,In_1529,In_1068);
and U665 (N_665,In_246,In_615);
or U666 (N_666,In_1979,In_1714);
xnor U667 (N_667,In_1480,In_325);
nand U668 (N_668,In_419,In_24);
or U669 (N_669,In_447,In_1524);
nor U670 (N_670,In_1479,In_549);
and U671 (N_671,In_1853,In_1626);
xor U672 (N_672,In_1641,In_1461);
or U673 (N_673,In_768,In_330);
nor U674 (N_674,In_1814,In_34);
nor U675 (N_675,In_1020,In_1031);
xor U676 (N_676,In_824,In_46);
or U677 (N_677,In_102,In_969);
xnor U678 (N_678,In_1101,In_1489);
xnor U679 (N_679,In_609,In_1102);
and U680 (N_680,In_1921,In_1914);
or U681 (N_681,In_1312,In_1978);
nor U682 (N_682,In_841,In_767);
nor U683 (N_683,In_1736,In_348);
nand U684 (N_684,In_1476,In_935);
nor U685 (N_685,In_1190,In_383);
xor U686 (N_686,In_1962,In_132);
nand U687 (N_687,In_1424,In_1239);
nand U688 (N_688,In_39,In_490);
and U689 (N_689,In_471,In_732);
nand U690 (N_690,In_228,In_1604);
or U691 (N_691,In_759,In_155);
or U692 (N_692,In_506,In_1983);
xnor U693 (N_693,In_601,In_1199);
nand U694 (N_694,In_204,In_648);
xnor U695 (N_695,In_658,In_1505);
and U696 (N_696,In_1534,In_1836);
and U697 (N_697,In_436,In_483);
nand U698 (N_698,In_912,In_108);
nand U699 (N_699,In_585,In_633);
nor U700 (N_700,In_1668,In_1393);
nand U701 (N_701,In_1692,In_1582);
xor U702 (N_702,In_439,In_306);
and U703 (N_703,In_1279,In_488);
nand U704 (N_704,In_666,In_1366);
nand U705 (N_705,In_1346,In_276);
nor U706 (N_706,In_510,In_161);
and U707 (N_707,In_1552,In_914);
xor U708 (N_708,In_1617,In_1819);
or U709 (N_709,In_665,In_963);
xor U710 (N_710,In_1339,In_588);
nor U711 (N_711,In_350,In_882);
nor U712 (N_712,In_925,In_1451);
and U713 (N_713,In_456,In_1169);
nand U714 (N_714,In_1141,In_1710);
or U715 (N_715,In_1793,In_757);
and U716 (N_716,In_868,In_1958);
or U717 (N_717,In_1388,In_1829);
and U718 (N_718,In_1374,In_30);
and U719 (N_719,In_1052,In_1299);
and U720 (N_720,In_589,In_763);
nand U721 (N_721,In_1460,In_1841);
or U722 (N_722,In_4,In_880);
xor U723 (N_723,In_1748,In_1311);
nand U724 (N_724,In_1681,In_1569);
nand U725 (N_725,In_1574,In_103);
nand U726 (N_726,In_786,In_1235);
nand U727 (N_727,In_1350,In_1049);
nor U728 (N_728,In_375,In_468);
and U729 (N_729,In_1188,In_610);
xnor U730 (N_730,In_1492,In_1676);
nand U731 (N_731,In_319,In_53);
nand U732 (N_732,In_1762,In_1487);
and U733 (N_733,In_1879,In_231);
nand U734 (N_734,In_42,In_174);
or U735 (N_735,In_248,In_536);
and U736 (N_736,In_620,In_504);
nor U737 (N_737,In_323,In_961);
nand U738 (N_738,In_1163,In_905);
and U739 (N_739,In_932,In_1706);
or U740 (N_740,In_307,In_1657);
or U741 (N_741,In_372,In_818);
and U742 (N_742,In_920,In_1763);
and U743 (N_743,In_1625,In_239);
and U744 (N_744,In_293,In_288);
nand U745 (N_745,In_1276,In_1252);
or U746 (N_746,In_1267,In_1989);
nor U747 (N_747,In_393,In_1883);
or U748 (N_748,In_1615,In_1721);
nor U749 (N_749,In_1293,In_769);
nor U750 (N_750,In_1136,In_1894);
nand U751 (N_751,In_1846,In_1694);
or U752 (N_752,In_1904,In_32);
nor U753 (N_753,In_292,In_1119);
or U754 (N_754,In_328,In_1789);
nor U755 (N_755,In_993,In_1830);
and U756 (N_756,In_1334,In_107);
nor U757 (N_757,In_1397,In_1236);
nor U758 (N_758,In_773,In_903);
nand U759 (N_759,In_1271,In_77);
and U760 (N_760,In_745,In_420);
xnor U761 (N_761,In_70,In_1328);
nand U762 (N_762,In_422,In_184);
or U763 (N_763,In_1660,In_1664);
nand U764 (N_764,In_984,In_1786);
nand U765 (N_765,In_1855,In_470);
xor U766 (N_766,In_858,In_1165);
and U767 (N_767,In_508,In_629);
or U768 (N_768,In_850,In_721);
or U769 (N_769,In_201,In_1075);
nand U770 (N_770,In_343,In_1469);
nor U771 (N_771,In_881,In_1367);
or U772 (N_772,In_1036,In_1916);
and U773 (N_773,In_1640,In_338);
nand U774 (N_774,In_780,In_1229);
xnor U775 (N_775,In_1316,In_1477);
or U776 (N_776,In_65,In_1032);
nor U777 (N_777,In_232,In_1026);
nand U778 (N_778,In_462,In_1413);
nor U779 (N_779,In_1348,In_1298);
nor U780 (N_780,In_1399,In_387);
or U781 (N_781,In_146,In_953);
and U782 (N_782,In_304,In_942);
and U783 (N_783,In_1114,In_1808);
nand U784 (N_784,In_1183,In_1751);
or U785 (N_785,In_979,In_936);
nand U786 (N_786,In_167,In_1321);
nand U787 (N_787,In_497,In_1541);
or U788 (N_788,In_29,In_672);
nand U789 (N_789,In_909,In_498);
xor U790 (N_790,In_257,In_244);
and U791 (N_791,In_962,In_1011);
xor U792 (N_792,In_1554,In_1370);
and U793 (N_793,In_703,In_503);
xnor U794 (N_794,In_1847,In_1734);
nand U795 (N_795,In_1352,In_1790);
and U796 (N_796,In_553,In_1588);
xor U797 (N_797,In_740,In_300);
nand U798 (N_798,In_1294,In_1145);
nor U799 (N_799,In_527,In_80);
nand U800 (N_800,In_1700,In_931);
or U801 (N_801,In_10,In_847);
and U802 (N_802,In_1795,In_560);
nand U803 (N_803,In_417,In_1336);
and U804 (N_804,In_1453,In_141);
xnor U805 (N_805,In_58,In_1586);
nand U806 (N_806,In_294,In_1926);
xnor U807 (N_807,In_499,In_1056);
nor U808 (N_808,In_1142,In_1768);
xnor U809 (N_809,In_1522,In_1351);
nor U810 (N_810,In_857,In_1121);
or U811 (N_811,In_261,In_44);
and U812 (N_812,In_1995,In_1266);
nor U813 (N_813,In_75,In_542);
and U814 (N_814,In_636,In_1842);
nor U815 (N_815,In_1144,In_264);
xnor U816 (N_816,In_474,In_415);
nor U817 (N_817,In_1558,In_1951);
nor U818 (N_818,In_1434,In_1466);
xnor U819 (N_819,In_1401,In_1285);
nor U820 (N_820,In_571,In_151);
nand U821 (N_821,In_806,In_1174);
or U822 (N_822,In_452,In_7);
and U823 (N_823,In_229,In_340);
xor U824 (N_824,In_1456,In_893);
nor U825 (N_825,In_1330,In_837);
nand U826 (N_826,In_1411,In_524);
xnor U827 (N_827,In_1782,In_1573);
nor U828 (N_828,In_727,In_1176);
nor U829 (N_829,In_578,In_443);
xnor U830 (N_830,In_1523,In_1301);
xnor U831 (N_831,In_989,In_1210);
nor U832 (N_832,In_35,In_864);
nor U833 (N_833,In_1590,In_1796);
and U834 (N_834,In_213,In_774);
xnor U835 (N_835,In_717,In_160);
or U836 (N_836,In_1008,In_1733);
nor U837 (N_837,In_1452,In_751);
or U838 (N_838,In_1621,In_28);
nor U839 (N_839,In_577,In_112);
xor U840 (N_840,In_975,In_195);
and U841 (N_841,In_1280,In_158);
or U842 (N_842,In_47,In_870);
nor U843 (N_843,In_543,In_630);
nor U844 (N_844,In_807,In_1349);
nand U845 (N_845,In_821,In_682);
nor U846 (N_846,In_624,In_896);
and U847 (N_847,In_815,In_0);
nand U848 (N_848,In_453,In_1332);
nand U849 (N_849,In_1984,In_73);
nor U850 (N_850,In_1125,In_515);
xnor U851 (N_851,In_405,In_1898);
or U852 (N_852,In_1682,In_663);
and U853 (N_853,In_1611,In_128);
nand U854 (N_854,In_955,In_1982);
nand U855 (N_855,In_1809,In_702);
nor U856 (N_856,In_1435,In_76);
and U857 (N_857,In_1701,In_735);
nand U858 (N_858,In_1148,In_1530);
or U859 (N_859,In_152,In_1644);
xnor U860 (N_860,In_142,In_1001);
or U861 (N_861,In_215,In_1614);
or U862 (N_862,In_313,In_494);
nand U863 (N_863,In_95,In_1498);
nand U864 (N_864,In_1024,In_1233);
xor U865 (N_865,In_1111,In_808);
or U866 (N_866,In_1944,In_581);
and U867 (N_867,In_1632,In_235);
nor U868 (N_868,In_901,In_926);
nor U869 (N_869,In_1696,In_1923);
or U870 (N_870,In_1212,In_1928);
nor U871 (N_871,In_1319,In_353);
or U872 (N_872,In_977,In_1674);
nand U873 (N_873,In_441,In_985);
or U874 (N_874,In_752,In_973);
nor U875 (N_875,In_344,In_153);
nand U876 (N_876,In_1099,In_540);
or U877 (N_877,In_965,In_1581);
nor U878 (N_878,In_1941,In_1270);
nor U879 (N_879,In_1047,In_391);
xnor U880 (N_880,In_431,In_1208);
xor U881 (N_881,In_336,In_395);
and U882 (N_882,In_407,In_476);
and U883 (N_883,In_1945,In_1776);
and U884 (N_884,In_1450,In_765);
nand U885 (N_885,In_363,In_379);
or U886 (N_886,In_1256,In_729);
nand U887 (N_887,In_449,In_1204);
xor U888 (N_888,In_234,In_1251);
and U889 (N_889,In_1863,In_661);
or U890 (N_890,In_1820,In_217);
nor U891 (N_891,In_550,In_1379);
xnor U892 (N_892,In_1096,In_1331);
xor U893 (N_893,In_1712,In_477);
nand U894 (N_894,In_670,In_1803);
nand U895 (N_895,In_1606,In_507);
xnor U896 (N_896,In_892,In_1283);
and U897 (N_897,In_1168,In_333);
and U898 (N_898,In_607,In_31);
nor U899 (N_899,In_406,In_60);
nor U900 (N_900,In_1416,In_171);
xor U901 (N_901,In_1642,In_1143);
xnor U902 (N_902,In_888,In_1073);
nor U903 (N_903,In_27,In_1358);
nand U904 (N_904,In_941,In_545);
xor U905 (N_905,In_1711,In_1741);
nand U906 (N_906,In_999,In_351);
or U907 (N_907,In_1807,In_1880);
and U908 (N_908,In_377,In_1368);
nand U909 (N_909,In_947,In_480);
xor U910 (N_910,In_725,In_104);
nor U911 (N_911,In_1677,In_625);
nor U912 (N_912,In_584,In_1258);
xor U913 (N_913,In_535,In_1055);
or U914 (N_914,In_516,In_1161);
xnor U915 (N_915,In_1865,In_623);
xnor U916 (N_916,In_1871,In_219);
nand U917 (N_917,In_1580,In_1481);
nor U918 (N_918,In_412,In_263);
xor U919 (N_919,In_637,In_1360);
or U920 (N_920,In_872,In_1017);
xnor U921 (N_921,In_1386,In_1027);
or U922 (N_922,In_298,In_425);
xor U923 (N_923,In_676,In_1507);
or U924 (N_924,In_1670,In_513);
or U925 (N_925,In_144,In_1495);
or U926 (N_926,In_1220,In_1289);
xnor U927 (N_927,In_744,In_1612);
or U928 (N_928,In_922,In_199);
or U929 (N_929,In_1286,In_1057);
and U930 (N_930,In_1103,In_1659);
xor U931 (N_931,In_876,In_1464);
xor U932 (N_932,In_1873,In_1864);
or U933 (N_933,In_562,In_121);
nand U934 (N_934,In_485,In_347);
xnor U935 (N_935,In_1622,In_2);
nor U936 (N_936,In_688,In_579);
or U937 (N_937,In_603,In_466);
xnor U938 (N_938,In_869,In_743);
nand U939 (N_939,In_845,In_1955);
xor U940 (N_940,In_641,In_862);
nand U941 (N_941,In_746,In_949);
nand U942 (N_942,In_1540,In_1788);
nand U943 (N_943,In_900,In_116);
nor U944 (N_944,In_628,In_874);
nand U945 (N_945,In_1361,In_1303);
nor U946 (N_946,In_1365,In_1576);
xor U947 (N_947,In_270,In_437);
and U948 (N_948,In_1282,In_1538);
nand U949 (N_949,In_1722,In_362);
nand U950 (N_950,In_1231,In_1218);
nor U951 (N_951,In_1725,In_52);
xor U952 (N_952,In_1225,In_87);
nand U953 (N_953,In_1003,In_100);
nand U954 (N_954,In_198,In_317);
or U955 (N_955,In_561,In_105);
xor U956 (N_956,In_649,In_990);
and U957 (N_957,In_1078,In_631);
nor U958 (N_958,In_635,In_1866);
xor U959 (N_959,In_811,In_1226);
nor U960 (N_960,In_1326,In_1186);
and U961 (N_961,In_1063,In_1708);
or U962 (N_962,In_668,In_1555);
nor U963 (N_963,In_1935,In_621);
and U964 (N_964,In_137,In_145);
or U965 (N_965,In_1520,In_954);
and U966 (N_966,In_968,In_1824);
xor U967 (N_967,In_1560,In_1471);
and U968 (N_968,In_662,In_1991);
and U969 (N_969,In_1969,In_596);
xor U970 (N_970,In_59,In_157);
and U971 (N_971,In_1631,In_297);
nor U972 (N_972,In_165,In_787);
nand U973 (N_973,In_1678,In_766);
and U974 (N_974,In_1927,In_1438);
xor U975 (N_975,In_565,In_873);
xnor U976 (N_976,In_710,In_1191);
xor U977 (N_977,In_12,In_801);
xor U978 (N_978,In_675,In_1243);
and U979 (N_979,In_940,In_1418);
nand U980 (N_980,In_996,In_777);
nand U981 (N_981,In_1089,In_1062);
and U982 (N_982,In_951,In_448);
and U983 (N_983,In_114,In_1378);
xnor U984 (N_984,In_723,In_1244);
nor U985 (N_985,In_209,In_1785);
or U986 (N_986,In_865,In_1107);
nand U987 (N_987,In_159,In_1093);
and U988 (N_988,In_61,In_800);
xnor U989 (N_989,In_1595,In_1061);
or U990 (N_990,In_368,In_799);
nand U991 (N_991,In_1647,In_1501);
and U992 (N_992,In_911,In_509);
or U993 (N_993,In_482,In_1234);
or U994 (N_994,In_659,In_689);
or U995 (N_995,In_1737,In_1160);
or U996 (N_996,In_1112,In_1876);
xnor U997 (N_997,In_1409,In_855);
xnor U998 (N_998,In_1426,In_268);
nand U999 (N_999,In_1917,In_1261);
or U1000 (N_1000,In_489,In_1202);
nor U1001 (N_1001,In_1938,In_502);
or U1002 (N_1002,In_1984,In_480);
and U1003 (N_1003,In_531,In_65);
nand U1004 (N_1004,In_1734,In_1924);
nor U1005 (N_1005,In_1099,In_1318);
xnor U1006 (N_1006,In_600,In_1524);
xor U1007 (N_1007,In_1898,In_64);
xnor U1008 (N_1008,In_1315,In_249);
nand U1009 (N_1009,In_1695,In_1778);
xnor U1010 (N_1010,In_14,In_1042);
xnor U1011 (N_1011,In_201,In_1917);
nor U1012 (N_1012,In_958,In_452);
xor U1013 (N_1013,In_570,In_464);
or U1014 (N_1014,In_1438,In_1771);
or U1015 (N_1015,In_691,In_1080);
or U1016 (N_1016,In_1440,In_173);
nor U1017 (N_1017,In_1299,In_543);
nand U1018 (N_1018,In_1555,In_1860);
xnor U1019 (N_1019,In_1842,In_323);
nor U1020 (N_1020,In_344,In_1999);
xnor U1021 (N_1021,In_176,In_1890);
nand U1022 (N_1022,In_1040,In_1523);
nand U1023 (N_1023,In_306,In_732);
and U1024 (N_1024,In_620,In_505);
nor U1025 (N_1025,In_153,In_128);
and U1026 (N_1026,In_677,In_1213);
and U1027 (N_1027,In_1955,In_1087);
xnor U1028 (N_1028,In_1640,In_876);
or U1029 (N_1029,In_510,In_1387);
and U1030 (N_1030,In_589,In_1164);
nor U1031 (N_1031,In_1511,In_1167);
xor U1032 (N_1032,In_937,In_455);
nand U1033 (N_1033,In_49,In_902);
and U1034 (N_1034,In_929,In_1302);
nand U1035 (N_1035,In_1999,In_941);
or U1036 (N_1036,In_1808,In_41);
nor U1037 (N_1037,In_508,In_1649);
nand U1038 (N_1038,In_687,In_1012);
nor U1039 (N_1039,In_629,In_312);
or U1040 (N_1040,In_1939,In_1837);
nor U1041 (N_1041,In_714,In_862);
or U1042 (N_1042,In_1214,In_75);
nand U1043 (N_1043,In_1415,In_528);
or U1044 (N_1044,In_862,In_1786);
nor U1045 (N_1045,In_207,In_1430);
xnor U1046 (N_1046,In_168,In_852);
xnor U1047 (N_1047,In_1547,In_391);
nor U1048 (N_1048,In_1198,In_1487);
nand U1049 (N_1049,In_1659,In_1837);
nand U1050 (N_1050,In_943,In_1164);
xnor U1051 (N_1051,In_228,In_748);
nand U1052 (N_1052,In_1080,In_359);
nand U1053 (N_1053,In_1441,In_675);
xor U1054 (N_1054,In_215,In_1767);
xor U1055 (N_1055,In_1721,In_210);
xnor U1056 (N_1056,In_1873,In_579);
and U1057 (N_1057,In_1709,In_101);
nor U1058 (N_1058,In_1252,In_771);
nand U1059 (N_1059,In_1725,In_1445);
nor U1060 (N_1060,In_67,In_1040);
and U1061 (N_1061,In_1654,In_1246);
xnor U1062 (N_1062,In_813,In_1140);
nor U1063 (N_1063,In_1646,In_365);
xnor U1064 (N_1064,In_1336,In_1768);
and U1065 (N_1065,In_426,In_1265);
xnor U1066 (N_1066,In_1369,In_851);
nand U1067 (N_1067,In_143,In_756);
nor U1068 (N_1068,In_878,In_1225);
xnor U1069 (N_1069,In_1549,In_543);
nand U1070 (N_1070,In_1197,In_1861);
or U1071 (N_1071,In_1436,In_1424);
nand U1072 (N_1072,In_615,In_581);
nand U1073 (N_1073,In_1126,In_1915);
or U1074 (N_1074,In_1034,In_1135);
and U1075 (N_1075,In_1258,In_667);
and U1076 (N_1076,In_106,In_890);
and U1077 (N_1077,In_1164,In_762);
or U1078 (N_1078,In_1647,In_412);
xor U1079 (N_1079,In_1746,In_673);
nor U1080 (N_1080,In_828,In_607);
xor U1081 (N_1081,In_1831,In_546);
nand U1082 (N_1082,In_893,In_244);
and U1083 (N_1083,In_1133,In_1314);
nor U1084 (N_1084,In_1594,In_1819);
and U1085 (N_1085,In_1414,In_1365);
and U1086 (N_1086,In_147,In_618);
or U1087 (N_1087,In_1308,In_1253);
xor U1088 (N_1088,In_1766,In_1593);
nor U1089 (N_1089,In_563,In_1143);
or U1090 (N_1090,In_1365,In_441);
nand U1091 (N_1091,In_1993,In_222);
nor U1092 (N_1092,In_1574,In_1210);
xnor U1093 (N_1093,In_1732,In_496);
and U1094 (N_1094,In_948,In_909);
xor U1095 (N_1095,In_1030,In_929);
nor U1096 (N_1096,In_828,In_594);
or U1097 (N_1097,In_1005,In_975);
and U1098 (N_1098,In_336,In_872);
nand U1099 (N_1099,In_578,In_506);
and U1100 (N_1100,In_1085,In_1369);
and U1101 (N_1101,In_674,In_1054);
xor U1102 (N_1102,In_766,In_374);
xnor U1103 (N_1103,In_1689,In_1136);
nand U1104 (N_1104,In_1465,In_1622);
nor U1105 (N_1105,In_1911,In_807);
or U1106 (N_1106,In_30,In_1854);
and U1107 (N_1107,In_1342,In_1409);
xor U1108 (N_1108,In_279,In_1848);
or U1109 (N_1109,In_1971,In_410);
and U1110 (N_1110,In_258,In_109);
nor U1111 (N_1111,In_1936,In_1670);
nor U1112 (N_1112,In_485,In_1412);
nor U1113 (N_1113,In_81,In_517);
nand U1114 (N_1114,In_352,In_1019);
nor U1115 (N_1115,In_1721,In_1056);
xor U1116 (N_1116,In_330,In_1549);
or U1117 (N_1117,In_1787,In_1943);
xor U1118 (N_1118,In_1236,In_460);
nor U1119 (N_1119,In_557,In_808);
and U1120 (N_1120,In_891,In_20);
nor U1121 (N_1121,In_1948,In_78);
nor U1122 (N_1122,In_619,In_497);
nor U1123 (N_1123,In_1603,In_832);
and U1124 (N_1124,In_1220,In_1202);
nand U1125 (N_1125,In_602,In_1732);
xor U1126 (N_1126,In_357,In_6);
xnor U1127 (N_1127,In_1637,In_138);
nand U1128 (N_1128,In_697,In_302);
nand U1129 (N_1129,In_433,In_96);
and U1130 (N_1130,In_1803,In_240);
or U1131 (N_1131,In_125,In_841);
or U1132 (N_1132,In_104,In_1507);
or U1133 (N_1133,In_1037,In_274);
and U1134 (N_1134,In_944,In_401);
nor U1135 (N_1135,In_165,In_1453);
and U1136 (N_1136,In_855,In_1207);
xor U1137 (N_1137,In_408,In_178);
xnor U1138 (N_1138,In_347,In_1615);
or U1139 (N_1139,In_34,In_1705);
nand U1140 (N_1140,In_1333,In_139);
xnor U1141 (N_1141,In_1101,In_1831);
nor U1142 (N_1142,In_584,In_1798);
and U1143 (N_1143,In_1434,In_815);
and U1144 (N_1144,In_1781,In_724);
and U1145 (N_1145,In_434,In_1039);
and U1146 (N_1146,In_1603,In_1593);
nor U1147 (N_1147,In_1280,In_1433);
and U1148 (N_1148,In_945,In_482);
or U1149 (N_1149,In_216,In_912);
xor U1150 (N_1150,In_1486,In_1644);
and U1151 (N_1151,In_899,In_1473);
xnor U1152 (N_1152,In_391,In_1844);
nor U1153 (N_1153,In_271,In_1134);
nand U1154 (N_1154,In_298,In_1303);
xor U1155 (N_1155,In_1578,In_1060);
or U1156 (N_1156,In_1431,In_1591);
nand U1157 (N_1157,In_361,In_560);
nand U1158 (N_1158,In_87,In_387);
xor U1159 (N_1159,In_974,In_492);
nor U1160 (N_1160,In_1036,In_308);
xnor U1161 (N_1161,In_1338,In_1693);
and U1162 (N_1162,In_892,In_1782);
xor U1163 (N_1163,In_1018,In_394);
or U1164 (N_1164,In_1436,In_851);
and U1165 (N_1165,In_339,In_1397);
xor U1166 (N_1166,In_706,In_484);
or U1167 (N_1167,In_1204,In_1652);
or U1168 (N_1168,In_932,In_584);
nand U1169 (N_1169,In_1714,In_1489);
xnor U1170 (N_1170,In_441,In_547);
nor U1171 (N_1171,In_527,In_307);
or U1172 (N_1172,In_1697,In_1295);
nand U1173 (N_1173,In_1605,In_357);
or U1174 (N_1174,In_548,In_955);
and U1175 (N_1175,In_1213,In_1984);
and U1176 (N_1176,In_1928,In_498);
nor U1177 (N_1177,In_1620,In_865);
nor U1178 (N_1178,In_1172,In_1960);
or U1179 (N_1179,In_1113,In_870);
or U1180 (N_1180,In_1592,In_665);
nor U1181 (N_1181,In_65,In_1548);
xor U1182 (N_1182,In_1277,In_210);
and U1183 (N_1183,In_740,In_891);
nor U1184 (N_1184,In_1849,In_1161);
nor U1185 (N_1185,In_1743,In_800);
xor U1186 (N_1186,In_1519,In_661);
or U1187 (N_1187,In_706,In_225);
and U1188 (N_1188,In_1869,In_1632);
nand U1189 (N_1189,In_1745,In_1610);
nor U1190 (N_1190,In_568,In_939);
xnor U1191 (N_1191,In_1180,In_1369);
or U1192 (N_1192,In_593,In_649);
and U1193 (N_1193,In_1418,In_1460);
and U1194 (N_1194,In_1377,In_1001);
nor U1195 (N_1195,In_1888,In_1424);
nand U1196 (N_1196,In_1061,In_168);
nor U1197 (N_1197,In_1702,In_1010);
xnor U1198 (N_1198,In_1275,In_1284);
or U1199 (N_1199,In_39,In_1928);
nand U1200 (N_1200,In_1912,In_1088);
xnor U1201 (N_1201,In_923,In_1554);
or U1202 (N_1202,In_469,In_1718);
nor U1203 (N_1203,In_865,In_260);
xor U1204 (N_1204,In_1113,In_16);
and U1205 (N_1205,In_375,In_926);
nand U1206 (N_1206,In_1725,In_970);
nand U1207 (N_1207,In_330,In_645);
xor U1208 (N_1208,In_83,In_1552);
nand U1209 (N_1209,In_1501,In_20);
and U1210 (N_1210,In_21,In_965);
nor U1211 (N_1211,In_68,In_1835);
nor U1212 (N_1212,In_273,In_962);
nand U1213 (N_1213,In_80,In_1901);
and U1214 (N_1214,In_1089,In_414);
nand U1215 (N_1215,In_1568,In_256);
or U1216 (N_1216,In_1415,In_378);
xnor U1217 (N_1217,In_1841,In_1462);
or U1218 (N_1218,In_960,In_1745);
nand U1219 (N_1219,In_391,In_1619);
and U1220 (N_1220,In_1743,In_606);
nand U1221 (N_1221,In_1298,In_1327);
or U1222 (N_1222,In_325,In_25);
nor U1223 (N_1223,In_564,In_61);
xnor U1224 (N_1224,In_1263,In_1660);
nand U1225 (N_1225,In_1014,In_65);
xor U1226 (N_1226,In_451,In_623);
nor U1227 (N_1227,In_588,In_1810);
xor U1228 (N_1228,In_537,In_1673);
xor U1229 (N_1229,In_938,In_100);
xor U1230 (N_1230,In_82,In_1614);
or U1231 (N_1231,In_837,In_1759);
xor U1232 (N_1232,In_1633,In_763);
nand U1233 (N_1233,In_1363,In_1423);
nor U1234 (N_1234,In_736,In_1961);
and U1235 (N_1235,In_575,In_744);
xnor U1236 (N_1236,In_1371,In_372);
nand U1237 (N_1237,In_1944,In_720);
nand U1238 (N_1238,In_1073,In_1355);
xor U1239 (N_1239,In_36,In_535);
nor U1240 (N_1240,In_1640,In_1872);
xor U1241 (N_1241,In_1331,In_665);
nor U1242 (N_1242,In_1100,In_1668);
nand U1243 (N_1243,In_677,In_684);
nor U1244 (N_1244,In_1974,In_21);
nor U1245 (N_1245,In_797,In_231);
or U1246 (N_1246,In_416,In_377);
and U1247 (N_1247,In_274,In_1451);
nor U1248 (N_1248,In_580,In_95);
nor U1249 (N_1249,In_1259,In_441);
and U1250 (N_1250,In_10,In_372);
nor U1251 (N_1251,In_1508,In_1273);
xor U1252 (N_1252,In_343,In_1066);
nor U1253 (N_1253,In_1283,In_446);
nand U1254 (N_1254,In_702,In_1775);
or U1255 (N_1255,In_735,In_102);
nand U1256 (N_1256,In_1340,In_346);
nor U1257 (N_1257,In_1302,In_1325);
and U1258 (N_1258,In_893,In_1004);
and U1259 (N_1259,In_1870,In_589);
xnor U1260 (N_1260,In_1554,In_1231);
or U1261 (N_1261,In_909,In_189);
and U1262 (N_1262,In_564,In_1475);
and U1263 (N_1263,In_1908,In_1185);
nor U1264 (N_1264,In_531,In_972);
xnor U1265 (N_1265,In_608,In_1074);
or U1266 (N_1266,In_571,In_1028);
nand U1267 (N_1267,In_668,In_327);
or U1268 (N_1268,In_807,In_124);
or U1269 (N_1269,In_319,In_766);
nand U1270 (N_1270,In_1647,In_51);
xor U1271 (N_1271,In_688,In_1602);
nand U1272 (N_1272,In_704,In_1736);
or U1273 (N_1273,In_1353,In_570);
nor U1274 (N_1274,In_1479,In_760);
nand U1275 (N_1275,In_1626,In_682);
nor U1276 (N_1276,In_1258,In_1337);
xor U1277 (N_1277,In_1713,In_1625);
and U1278 (N_1278,In_460,In_1756);
xor U1279 (N_1279,In_1070,In_846);
xor U1280 (N_1280,In_1877,In_520);
and U1281 (N_1281,In_1469,In_1188);
or U1282 (N_1282,In_1889,In_583);
or U1283 (N_1283,In_1626,In_1866);
xor U1284 (N_1284,In_542,In_1364);
nor U1285 (N_1285,In_953,In_1595);
nor U1286 (N_1286,In_1402,In_1472);
or U1287 (N_1287,In_979,In_977);
nand U1288 (N_1288,In_1641,In_1655);
nor U1289 (N_1289,In_461,In_722);
and U1290 (N_1290,In_411,In_1729);
and U1291 (N_1291,In_1476,In_1621);
and U1292 (N_1292,In_1396,In_145);
nand U1293 (N_1293,In_737,In_151);
or U1294 (N_1294,In_1044,In_165);
nor U1295 (N_1295,In_1603,In_1264);
or U1296 (N_1296,In_909,In_1411);
nor U1297 (N_1297,In_624,In_1346);
nand U1298 (N_1298,In_926,In_1912);
or U1299 (N_1299,In_1211,In_927);
nand U1300 (N_1300,In_1256,In_829);
nand U1301 (N_1301,In_660,In_600);
nand U1302 (N_1302,In_1018,In_1006);
nor U1303 (N_1303,In_406,In_453);
nand U1304 (N_1304,In_297,In_1346);
xnor U1305 (N_1305,In_1745,In_1395);
nor U1306 (N_1306,In_1666,In_342);
or U1307 (N_1307,In_1553,In_1118);
and U1308 (N_1308,In_1014,In_696);
xnor U1309 (N_1309,In_1000,In_894);
or U1310 (N_1310,In_378,In_578);
nor U1311 (N_1311,In_1446,In_480);
and U1312 (N_1312,In_1097,In_860);
and U1313 (N_1313,In_314,In_30);
and U1314 (N_1314,In_581,In_1713);
or U1315 (N_1315,In_1660,In_468);
nand U1316 (N_1316,In_1524,In_651);
and U1317 (N_1317,In_1880,In_1636);
nor U1318 (N_1318,In_1637,In_1309);
or U1319 (N_1319,In_1195,In_945);
nand U1320 (N_1320,In_1304,In_318);
or U1321 (N_1321,In_1960,In_995);
nor U1322 (N_1322,In_1633,In_1625);
xor U1323 (N_1323,In_514,In_1946);
xor U1324 (N_1324,In_1668,In_1436);
nand U1325 (N_1325,In_871,In_1341);
nand U1326 (N_1326,In_1811,In_791);
xor U1327 (N_1327,In_1867,In_443);
or U1328 (N_1328,In_757,In_342);
nand U1329 (N_1329,In_1571,In_1746);
xor U1330 (N_1330,In_220,In_880);
nand U1331 (N_1331,In_610,In_914);
and U1332 (N_1332,In_309,In_1242);
nor U1333 (N_1333,In_1736,In_680);
nor U1334 (N_1334,In_873,In_1383);
xor U1335 (N_1335,In_664,In_358);
xor U1336 (N_1336,In_623,In_102);
nor U1337 (N_1337,In_1592,In_1400);
or U1338 (N_1338,In_1200,In_524);
nor U1339 (N_1339,In_1608,In_189);
and U1340 (N_1340,In_615,In_90);
xnor U1341 (N_1341,In_447,In_1788);
or U1342 (N_1342,In_1771,In_777);
nor U1343 (N_1343,In_880,In_826);
or U1344 (N_1344,In_968,In_1056);
nand U1345 (N_1345,In_732,In_891);
and U1346 (N_1346,In_1461,In_21);
nand U1347 (N_1347,In_1554,In_190);
nand U1348 (N_1348,In_1596,In_1227);
nand U1349 (N_1349,In_1331,In_699);
and U1350 (N_1350,In_1405,In_205);
nand U1351 (N_1351,In_1942,In_1523);
or U1352 (N_1352,In_1999,In_1792);
and U1353 (N_1353,In_1803,In_154);
and U1354 (N_1354,In_289,In_929);
xor U1355 (N_1355,In_1499,In_474);
and U1356 (N_1356,In_1580,In_1860);
nor U1357 (N_1357,In_1070,In_991);
and U1358 (N_1358,In_695,In_833);
xor U1359 (N_1359,In_576,In_550);
xor U1360 (N_1360,In_223,In_1000);
nand U1361 (N_1361,In_932,In_889);
and U1362 (N_1362,In_556,In_1414);
xor U1363 (N_1363,In_679,In_1833);
and U1364 (N_1364,In_549,In_960);
nor U1365 (N_1365,In_1685,In_756);
or U1366 (N_1366,In_385,In_1974);
xor U1367 (N_1367,In_1942,In_1317);
nand U1368 (N_1368,In_1161,In_599);
nor U1369 (N_1369,In_120,In_1865);
nor U1370 (N_1370,In_100,In_873);
xor U1371 (N_1371,In_1000,In_332);
nand U1372 (N_1372,In_793,In_727);
nor U1373 (N_1373,In_1322,In_1644);
xnor U1374 (N_1374,In_394,In_1285);
and U1375 (N_1375,In_1086,In_684);
and U1376 (N_1376,In_596,In_936);
or U1377 (N_1377,In_784,In_463);
xor U1378 (N_1378,In_1747,In_1190);
and U1379 (N_1379,In_758,In_1734);
and U1380 (N_1380,In_233,In_1071);
nor U1381 (N_1381,In_1305,In_1303);
and U1382 (N_1382,In_988,In_1252);
or U1383 (N_1383,In_1660,In_872);
nor U1384 (N_1384,In_1305,In_1969);
or U1385 (N_1385,In_735,In_1799);
xor U1386 (N_1386,In_1711,In_1514);
nor U1387 (N_1387,In_238,In_423);
or U1388 (N_1388,In_1126,In_616);
or U1389 (N_1389,In_632,In_1874);
nor U1390 (N_1390,In_684,In_296);
nand U1391 (N_1391,In_1574,In_1822);
or U1392 (N_1392,In_1679,In_1155);
or U1393 (N_1393,In_1008,In_1073);
or U1394 (N_1394,In_1744,In_404);
or U1395 (N_1395,In_898,In_279);
and U1396 (N_1396,In_628,In_384);
and U1397 (N_1397,In_1636,In_300);
nor U1398 (N_1398,In_1813,In_862);
and U1399 (N_1399,In_1751,In_330);
nand U1400 (N_1400,In_1277,In_432);
or U1401 (N_1401,In_1189,In_1148);
xor U1402 (N_1402,In_1992,In_885);
nand U1403 (N_1403,In_708,In_1566);
nand U1404 (N_1404,In_1470,In_672);
xnor U1405 (N_1405,In_1938,In_724);
xor U1406 (N_1406,In_1072,In_959);
and U1407 (N_1407,In_898,In_358);
xnor U1408 (N_1408,In_1250,In_1304);
nand U1409 (N_1409,In_1773,In_1167);
nor U1410 (N_1410,In_41,In_1002);
or U1411 (N_1411,In_1858,In_584);
or U1412 (N_1412,In_1905,In_1468);
or U1413 (N_1413,In_1424,In_246);
and U1414 (N_1414,In_1681,In_876);
nand U1415 (N_1415,In_1566,In_1774);
or U1416 (N_1416,In_721,In_1146);
and U1417 (N_1417,In_1097,In_1022);
and U1418 (N_1418,In_1449,In_645);
or U1419 (N_1419,In_504,In_1892);
nand U1420 (N_1420,In_158,In_269);
and U1421 (N_1421,In_1333,In_1749);
and U1422 (N_1422,In_1178,In_1829);
xor U1423 (N_1423,In_78,In_123);
and U1424 (N_1424,In_181,In_1670);
nor U1425 (N_1425,In_1271,In_1544);
xnor U1426 (N_1426,In_1398,In_1064);
xor U1427 (N_1427,In_1822,In_384);
xnor U1428 (N_1428,In_604,In_1149);
nor U1429 (N_1429,In_304,In_615);
nand U1430 (N_1430,In_926,In_531);
and U1431 (N_1431,In_1143,In_539);
xor U1432 (N_1432,In_258,In_1442);
and U1433 (N_1433,In_1261,In_242);
xor U1434 (N_1434,In_1216,In_991);
nand U1435 (N_1435,In_195,In_1977);
nor U1436 (N_1436,In_1594,In_636);
and U1437 (N_1437,In_958,In_899);
xnor U1438 (N_1438,In_391,In_1126);
nand U1439 (N_1439,In_730,In_390);
and U1440 (N_1440,In_15,In_226);
nor U1441 (N_1441,In_1733,In_616);
xor U1442 (N_1442,In_1079,In_919);
xor U1443 (N_1443,In_1432,In_1669);
and U1444 (N_1444,In_604,In_192);
xnor U1445 (N_1445,In_845,In_1737);
xnor U1446 (N_1446,In_1714,In_1766);
nand U1447 (N_1447,In_1178,In_1235);
xor U1448 (N_1448,In_1573,In_282);
nor U1449 (N_1449,In_629,In_1614);
and U1450 (N_1450,In_507,In_875);
xnor U1451 (N_1451,In_1373,In_866);
and U1452 (N_1452,In_851,In_231);
and U1453 (N_1453,In_1461,In_1651);
or U1454 (N_1454,In_656,In_1005);
and U1455 (N_1455,In_1537,In_343);
or U1456 (N_1456,In_1593,In_1373);
xnor U1457 (N_1457,In_1582,In_1455);
and U1458 (N_1458,In_718,In_1634);
nor U1459 (N_1459,In_1033,In_1287);
and U1460 (N_1460,In_297,In_180);
nor U1461 (N_1461,In_1490,In_1342);
or U1462 (N_1462,In_844,In_1226);
nand U1463 (N_1463,In_1480,In_1144);
nor U1464 (N_1464,In_642,In_1464);
and U1465 (N_1465,In_1498,In_1564);
xor U1466 (N_1466,In_1474,In_1495);
or U1467 (N_1467,In_1483,In_1627);
nand U1468 (N_1468,In_224,In_1618);
xor U1469 (N_1469,In_916,In_1541);
xnor U1470 (N_1470,In_416,In_772);
nand U1471 (N_1471,In_1936,In_426);
or U1472 (N_1472,In_1972,In_796);
or U1473 (N_1473,In_1347,In_668);
xor U1474 (N_1474,In_575,In_594);
nor U1475 (N_1475,In_1866,In_1996);
and U1476 (N_1476,In_339,In_1936);
xnor U1477 (N_1477,In_733,In_1327);
nor U1478 (N_1478,In_1187,In_1132);
nor U1479 (N_1479,In_1966,In_525);
nand U1480 (N_1480,In_343,In_1196);
xor U1481 (N_1481,In_1538,In_458);
nor U1482 (N_1482,In_1978,In_1336);
nand U1483 (N_1483,In_1208,In_1556);
nor U1484 (N_1484,In_600,In_555);
and U1485 (N_1485,In_793,In_896);
or U1486 (N_1486,In_1068,In_353);
or U1487 (N_1487,In_408,In_484);
nor U1488 (N_1488,In_696,In_299);
and U1489 (N_1489,In_1269,In_1804);
xor U1490 (N_1490,In_815,In_547);
or U1491 (N_1491,In_116,In_74);
or U1492 (N_1492,In_515,In_161);
and U1493 (N_1493,In_1728,In_42);
or U1494 (N_1494,In_1391,In_1362);
nand U1495 (N_1495,In_54,In_1559);
xnor U1496 (N_1496,In_1473,In_1837);
nand U1497 (N_1497,In_905,In_668);
or U1498 (N_1498,In_1734,In_1941);
or U1499 (N_1499,In_1283,In_373);
and U1500 (N_1500,In_411,In_207);
nor U1501 (N_1501,In_1032,In_1792);
and U1502 (N_1502,In_100,In_1918);
nor U1503 (N_1503,In_811,In_1540);
xor U1504 (N_1504,In_765,In_623);
and U1505 (N_1505,In_1469,In_324);
nand U1506 (N_1506,In_630,In_1591);
and U1507 (N_1507,In_1234,In_1837);
or U1508 (N_1508,In_279,In_1459);
nor U1509 (N_1509,In_1674,In_1040);
or U1510 (N_1510,In_1150,In_537);
xor U1511 (N_1511,In_276,In_1246);
xnor U1512 (N_1512,In_49,In_211);
or U1513 (N_1513,In_1862,In_1822);
or U1514 (N_1514,In_1479,In_1473);
or U1515 (N_1515,In_1290,In_1997);
xor U1516 (N_1516,In_1887,In_1572);
xor U1517 (N_1517,In_1460,In_5);
and U1518 (N_1518,In_493,In_499);
nand U1519 (N_1519,In_588,In_1265);
nor U1520 (N_1520,In_65,In_228);
nand U1521 (N_1521,In_234,In_1682);
nand U1522 (N_1522,In_1521,In_665);
nor U1523 (N_1523,In_1803,In_107);
nor U1524 (N_1524,In_1982,In_1459);
nor U1525 (N_1525,In_656,In_886);
or U1526 (N_1526,In_238,In_1990);
or U1527 (N_1527,In_471,In_855);
and U1528 (N_1528,In_1788,In_596);
nor U1529 (N_1529,In_1919,In_322);
nand U1530 (N_1530,In_663,In_754);
and U1531 (N_1531,In_1123,In_949);
nand U1532 (N_1532,In_150,In_503);
nor U1533 (N_1533,In_379,In_477);
nor U1534 (N_1534,In_1788,In_1688);
or U1535 (N_1535,In_1616,In_1040);
nand U1536 (N_1536,In_778,In_1970);
and U1537 (N_1537,In_1325,In_815);
or U1538 (N_1538,In_235,In_100);
nand U1539 (N_1539,In_1516,In_376);
nor U1540 (N_1540,In_1781,In_781);
and U1541 (N_1541,In_1932,In_1068);
or U1542 (N_1542,In_1606,In_864);
xor U1543 (N_1543,In_1540,In_1163);
nand U1544 (N_1544,In_1445,In_1578);
xnor U1545 (N_1545,In_472,In_1091);
nand U1546 (N_1546,In_933,In_1221);
and U1547 (N_1547,In_357,In_488);
and U1548 (N_1548,In_1493,In_967);
xor U1549 (N_1549,In_1580,In_26);
or U1550 (N_1550,In_1153,In_1788);
nor U1551 (N_1551,In_1234,In_41);
and U1552 (N_1552,In_1732,In_1137);
xnor U1553 (N_1553,In_1150,In_246);
nand U1554 (N_1554,In_1383,In_883);
or U1555 (N_1555,In_1358,In_907);
nand U1556 (N_1556,In_1693,In_1784);
xor U1557 (N_1557,In_1759,In_1694);
or U1558 (N_1558,In_1652,In_1888);
or U1559 (N_1559,In_1826,In_360);
nor U1560 (N_1560,In_1780,In_563);
nor U1561 (N_1561,In_326,In_19);
nand U1562 (N_1562,In_1212,In_355);
xnor U1563 (N_1563,In_1643,In_1903);
xor U1564 (N_1564,In_1811,In_1390);
nor U1565 (N_1565,In_543,In_589);
nand U1566 (N_1566,In_708,In_817);
or U1567 (N_1567,In_811,In_340);
xor U1568 (N_1568,In_1742,In_1944);
nor U1569 (N_1569,In_946,In_1203);
and U1570 (N_1570,In_1046,In_561);
or U1571 (N_1571,In_835,In_1734);
and U1572 (N_1572,In_1830,In_926);
or U1573 (N_1573,In_1828,In_1121);
nand U1574 (N_1574,In_575,In_630);
and U1575 (N_1575,In_1746,In_1995);
xnor U1576 (N_1576,In_1092,In_47);
nor U1577 (N_1577,In_475,In_176);
or U1578 (N_1578,In_694,In_1112);
nor U1579 (N_1579,In_189,In_73);
xor U1580 (N_1580,In_1303,In_895);
nand U1581 (N_1581,In_575,In_1138);
nor U1582 (N_1582,In_237,In_1538);
nor U1583 (N_1583,In_1716,In_593);
xnor U1584 (N_1584,In_947,In_881);
and U1585 (N_1585,In_135,In_1289);
xnor U1586 (N_1586,In_1310,In_727);
xor U1587 (N_1587,In_1762,In_1163);
and U1588 (N_1588,In_589,In_1736);
xnor U1589 (N_1589,In_695,In_506);
and U1590 (N_1590,In_1591,In_187);
xor U1591 (N_1591,In_920,In_549);
and U1592 (N_1592,In_1404,In_1850);
or U1593 (N_1593,In_547,In_294);
xnor U1594 (N_1594,In_1233,In_224);
or U1595 (N_1595,In_609,In_1809);
or U1596 (N_1596,In_521,In_1776);
nand U1597 (N_1597,In_630,In_512);
nor U1598 (N_1598,In_1544,In_540);
xor U1599 (N_1599,In_1647,In_216);
and U1600 (N_1600,In_954,In_419);
and U1601 (N_1601,In_1812,In_266);
and U1602 (N_1602,In_762,In_565);
nand U1603 (N_1603,In_898,In_1687);
and U1604 (N_1604,In_1555,In_93);
nand U1605 (N_1605,In_595,In_339);
and U1606 (N_1606,In_182,In_1025);
or U1607 (N_1607,In_1821,In_727);
or U1608 (N_1608,In_902,In_397);
xor U1609 (N_1609,In_1250,In_1220);
and U1610 (N_1610,In_1565,In_1007);
and U1611 (N_1611,In_1108,In_418);
xor U1612 (N_1612,In_157,In_975);
xnor U1613 (N_1613,In_1272,In_1779);
nor U1614 (N_1614,In_1239,In_716);
nor U1615 (N_1615,In_1721,In_1660);
xor U1616 (N_1616,In_237,In_413);
nor U1617 (N_1617,In_1398,In_540);
nor U1618 (N_1618,In_1771,In_1858);
or U1619 (N_1619,In_1118,In_1342);
nand U1620 (N_1620,In_927,In_1446);
or U1621 (N_1621,In_176,In_585);
or U1622 (N_1622,In_1468,In_396);
nor U1623 (N_1623,In_1239,In_1186);
nor U1624 (N_1624,In_310,In_758);
nand U1625 (N_1625,In_1418,In_933);
nand U1626 (N_1626,In_331,In_868);
xor U1627 (N_1627,In_114,In_1910);
and U1628 (N_1628,In_1275,In_1185);
nor U1629 (N_1629,In_1661,In_1260);
and U1630 (N_1630,In_1213,In_128);
and U1631 (N_1631,In_47,In_1066);
or U1632 (N_1632,In_1516,In_604);
and U1633 (N_1633,In_1585,In_1877);
nand U1634 (N_1634,In_196,In_1722);
or U1635 (N_1635,In_1373,In_708);
nor U1636 (N_1636,In_1720,In_608);
xnor U1637 (N_1637,In_958,In_245);
or U1638 (N_1638,In_446,In_1569);
and U1639 (N_1639,In_1886,In_451);
or U1640 (N_1640,In_1243,In_322);
nor U1641 (N_1641,In_893,In_1513);
and U1642 (N_1642,In_1333,In_1640);
or U1643 (N_1643,In_1789,In_809);
nand U1644 (N_1644,In_120,In_1704);
nor U1645 (N_1645,In_1191,In_448);
or U1646 (N_1646,In_1031,In_1603);
and U1647 (N_1647,In_686,In_636);
and U1648 (N_1648,In_775,In_940);
and U1649 (N_1649,In_1338,In_1676);
nor U1650 (N_1650,In_227,In_1535);
nand U1651 (N_1651,In_724,In_1399);
and U1652 (N_1652,In_1062,In_1016);
and U1653 (N_1653,In_179,In_550);
xor U1654 (N_1654,In_329,In_793);
xor U1655 (N_1655,In_921,In_1470);
and U1656 (N_1656,In_1353,In_1877);
and U1657 (N_1657,In_881,In_1429);
xor U1658 (N_1658,In_1762,In_856);
nor U1659 (N_1659,In_332,In_460);
and U1660 (N_1660,In_1517,In_891);
xnor U1661 (N_1661,In_688,In_1783);
or U1662 (N_1662,In_1188,In_526);
xor U1663 (N_1663,In_412,In_1156);
or U1664 (N_1664,In_1962,In_1035);
or U1665 (N_1665,In_1001,In_546);
nor U1666 (N_1666,In_444,In_168);
and U1667 (N_1667,In_1201,In_974);
nand U1668 (N_1668,In_954,In_97);
and U1669 (N_1669,In_1554,In_940);
xnor U1670 (N_1670,In_756,In_726);
nand U1671 (N_1671,In_30,In_246);
and U1672 (N_1672,In_384,In_916);
xor U1673 (N_1673,In_444,In_1342);
nor U1674 (N_1674,In_872,In_544);
or U1675 (N_1675,In_435,In_697);
nand U1676 (N_1676,In_1144,In_954);
or U1677 (N_1677,In_775,In_565);
and U1678 (N_1678,In_446,In_1808);
nand U1679 (N_1679,In_1017,In_365);
xnor U1680 (N_1680,In_688,In_1158);
nand U1681 (N_1681,In_793,In_0);
nor U1682 (N_1682,In_420,In_1771);
xnor U1683 (N_1683,In_1622,In_214);
or U1684 (N_1684,In_1171,In_281);
nor U1685 (N_1685,In_1970,In_1075);
nand U1686 (N_1686,In_789,In_1455);
or U1687 (N_1687,In_237,In_1751);
and U1688 (N_1688,In_916,In_1794);
or U1689 (N_1689,In_1152,In_1868);
nand U1690 (N_1690,In_205,In_526);
nand U1691 (N_1691,In_1634,In_662);
nand U1692 (N_1692,In_1475,In_892);
or U1693 (N_1693,In_40,In_1181);
and U1694 (N_1694,In_328,In_218);
nor U1695 (N_1695,In_1937,In_1250);
xnor U1696 (N_1696,In_1853,In_121);
and U1697 (N_1697,In_1619,In_657);
nand U1698 (N_1698,In_699,In_445);
and U1699 (N_1699,In_732,In_1423);
nand U1700 (N_1700,In_200,In_1839);
and U1701 (N_1701,In_1819,In_503);
xnor U1702 (N_1702,In_66,In_559);
and U1703 (N_1703,In_1977,In_1278);
and U1704 (N_1704,In_1678,In_1594);
nor U1705 (N_1705,In_373,In_1396);
nand U1706 (N_1706,In_1167,In_1358);
nand U1707 (N_1707,In_1239,In_821);
or U1708 (N_1708,In_177,In_1626);
or U1709 (N_1709,In_1357,In_1866);
xor U1710 (N_1710,In_349,In_38);
nand U1711 (N_1711,In_500,In_849);
or U1712 (N_1712,In_387,In_557);
nand U1713 (N_1713,In_1392,In_1363);
or U1714 (N_1714,In_1677,In_5);
xor U1715 (N_1715,In_753,In_1881);
nor U1716 (N_1716,In_912,In_1637);
and U1717 (N_1717,In_1638,In_267);
nand U1718 (N_1718,In_1607,In_433);
or U1719 (N_1719,In_204,In_257);
and U1720 (N_1720,In_1779,In_1672);
nand U1721 (N_1721,In_131,In_166);
and U1722 (N_1722,In_1643,In_1036);
xor U1723 (N_1723,In_1647,In_133);
nand U1724 (N_1724,In_1828,In_596);
or U1725 (N_1725,In_1127,In_1288);
nor U1726 (N_1726,In_1999,In_1716);
nand U1727 (N_1727,In_1823,In_990);
nor U1728 (N_1728,In_365,In_717);
nor U1729 (N_1729,In_99,In_1936);
and U1730 (N_1730,In_363,In_1215);
or U1731 (N_1731,In_1574,In_1976);
and U1732 (N_1732,In_1270,In_86);
and U1733 (N_1733,In_910,In_939);
or U1734 (N_1734,In_1454,In_1045);
xor U1735 (N_1735,In_1110,In_1538);
or U1736 (N_1736,In_1311,In_1192);
or U1737 (N_1737,In_702,In_954);
and U1738 (N_1738,In_1219,In_749);
and U1739 (N_1739,In_1518,In_1694);
and U1740 (N_1740,In_1140,In_373);
nand U1741 (N_1741,In_1737,In_405);
nor U1742 (N_1742,In_367,In_1050);
or U1743 (N_1743,In_1759,In_526);
or U1744 (N_1744,In_1035,In_1634);
nand U1745 (N_1745,In_366,In_464);
xor U1746 (N_1746,In_612,In_1641);
or U1747 (N_1747,In_1674,In_1894);
or U1748 (N_1748,In_140,In_1691);
and U1749 (N_1749,In_1622,In_1050);
or U1750 (N_1750,In_1764,In_1391);
or U1751 (N_1751,In_162,In_552);
nor U1752 (N_1752,In_1921,In_89);
nand U1753 (N_1753,In_1500,In_520);
nor U1754 (N_1754,In_185,In_1866);
xnor U1755 (N_1755,In_457,In_979);
xnor U1756 (N_1756,In_1930,In_951);
or U1757 (N_1757,In_748,In_931);
xor U1758 (N_1758,In_313,In_870);
and U1759 (N_1759,In_1221,In_1145);
or U1760 (N_1760,In_611,In_725);
or U1761 (N_1761,In_1571,In_1817);
or U1762 (N_1762,In_1895,In_933);
xor U1763 (N_1763,In_1297,In_210);
xnor U1764 (N_1764,In_780,In_205);
nand U1765 (N_1765,In_1459,In_687);
or U1766 (N_1766,In_1497,In_33);
xor U1767 (N_1767,In_559,In_879);
xnor U1768 (N_1768,In_1037,In_1392);
nand U1769 (N_1769,In_623,In_20);
or U1770 (N_1770,In_437,In_923);
nor U1771 (N_1771,In_158,In_446);
nor U1772 (N_1772,In_547,In_1345);
nand U1773 (N_1773,In_500,In_1571);
nand U1774 (N_1774,In_456,In_625);
nand U1775 (N_1775,In_1342,In_1548);
nand U1776 (N_1776,In_1040,In_1647);
nor U1777 (N_1777,In_1439,In_1730);
nand U1778 (N_1778,In_903,In_537);
xor U1779 (N_1779,In_791,In_627);
and U1780 (N_1780,In_1055,In_764);
or U1781 (N_1781,In_700,In_1765);
nor U1782 (N_1782,In_425,In_617);
or U1783 (N_1783,In_1969,In_1561);
nor U1784 (N_1784,In_209,In_1464);
nand U1785 (N_1785,In_1358,In_533);
nand U1786 (N_1786,In_742,In_1820);
nand U1787 (N_1787,In_290,In_1041);
xor U1788 (N_1788,In_1403,In_1828);
nand U1789 (N_1789,In_159,In_1952);
and U1790 (N_1790,In_299,In_925);
nor U1791 (N_1791,In_1605,In_23);
xnor U1792 (N_1792,In_598,In_1083);
nand U1793 (N_1793,In_1169,In_1116);
or U1794 (N_1794,In_1836,In_308);
nor U1795 (N_1795,In_1532,In_1005);
nor U1796 (N_1796,In_666,In_1551);
and U1797 (N_1797,In_474,In_315);
xnor U1798 (N_1798,In_706,In_1006);
nand U1799 (N_1799,In_625,In_304);
nor U1800 (N_1800,In_1543,In_1143);
or U1801 (N_1801,In_1796,In_352);
and U1802 (N_1802,In_1585,In_642);
or U1803 (N_1803,In_594,In_837);
and U1804 (N_1804,In_697,In_1032);
nor U1805 (N_1805,In_1546,In_1762);
xnor U1806 (N_1806,In_371,In_1247);
xnor U1807 (N_1807,In_1865,In_601);
nor U1808 (N_1808,In_667,In_1368);
nand U1809 (N_1809,In_505,In_47);
or U1810 (N_1810,In_516,In_1656);
nand U1811 (N_1811,In_1727,In_428);
nand U1812 (N_1812,In_434,In_1771);
nand U1813 (N_1813,In_338,In_732);
xnor U1814 (N_1814,In_877,In_675);
xnor U1815 (N_1815,In_696,In_152);
nor U1816 (N_1816,In_1392,In_1007);
nand U1817 (N_1817,In_1742,In_423);
and U1818 (N_1818,In_129,In_1610);
xor U1819 (N_1819,In_848,In_301);
nor U1820 (N_1820,In_919,In_1402);
nor U1821 (N_1821,In_1494,In_636);
and U1822 (N_1822,In_1254,In_977);
xor U1823 (N_1823,In_1383,In_1197);
nand U1824 (N_1824,In_1890,In_764);
xnor U1825 (N_1825,In_1987,In_1370);
nand U1826 (N_1826,In_1720,In_635);
or U1827 (N_1827,In_1938,In_1821);
nand U1828 (N_1828,In_701,In_616);
xnor U1829 (N_1829,In_246,In_1006);
or U1830 (N_1830,In_1263,In_1007);
nand U1831 (N_1831,In_1343,In_729);
xnor U1832 (N_1832,In_1457,In_66);
or U1833 (N_1833,In_263,In_994);
nand U1834 (N_1834,In_1390,In_326);
xnor U1835 (N_1835,In_1008,In_715);
nor U1836 (N_1836,In_159,In_989);
nand U1837 (N_1837,In_1583,In_1695);
nor U1838 (N_1838,In_1555,In_60);
nand U1839 (N_1839,In_1669,In_1581);
xor U1840 (N_1840,In_391,In_1111);
xor U1841 (N_1841,In_1050,In_217);
and U1842 (N_1842,In_1587,In_1898);
xor U1843 (N_1843,In_1989,In_1474);
nor U1844 (N_1844,In_1840,In_1356);
xor U1845 (N_1845,In_1485,In_693);
xor U1846 (N_1846,In_1082,In_1239);
nor U1847 (N_1847,In_1530,In_1283);
and U1848 (N_1848,In_1416,In_426);
xnor U1849 (N_1849,In_1688,In_780);
nand U1850 (N_1850,In_1357,In_1107);
xor U1851 (N_1851,In_890,In_711);
or U1852 (N_1852,In_765,In_1074);
nand U1853 (N_1853,In_1380,In_900);
xor U1854 (N_1854,In_1229,In_1837);
nor U1855 (N_1855,In_421,In_783);
or U1856 (N_1856,In_271,In_943);
or U1857 (N_1857,In_671,In_793);
nand U1858 (N_1858,In_1702,In_1048);
nor U1859 (N_1859,In_652,In_1404);
nor U1860 (N_1860,In_611,In_1122);
xnor U1861 (N_1861,In_1356,In_1842);
nand U1862 (N_1862,In_1855,In_1126);
nand U1863 (N_1863,In_1487,In_38);
nor U1864 (N_1864,In_1811,In_1208);
nor U1865 (N_1865,In_659,In_762);
and U1866 (N_1866,In_1083,In_794);
or U1867 (N_1867,In_883,In_1734);
nand U1868 (N_1868,In_64,In_933);
or U1869 (N_1869,In_1191,In_268);
or U1870 (N_1870,In_1332,In_1006);
xnor U1871 (N_1871,In_1103,In_416);
and U1872 (N_1872,In_1369,In_85);
and U1873 (N_1873,In_999,In_840);
xor U1874 (N_1874,In_888,In_932);
nor U1875 (N_1875,In_1413,In_1889);
nand U1876 (N_1876,In_686,In_1585);
and U1877 (N_1877,In_370,In_942);
and U1878 (N_1878,In_778,In_997);
nor U1879 (N_1879,In_1405,In_604);
and U1880 (N_1880,In_74,In_1531);
xnor U1881 (N_1881,In_1326,In_99);
nor U1882 (N_1882,In_1359,In_1553);
or U1883 (N_1883,In_1062,In_1349);
and U1884 (N_1884,In_627,In_460);
xor U1885 (N_1885,In_1379,In_1801);
and U1886 (N_1886,In_1171,In_1313);
or U1887 (N_1887,In_425,In_759);
or U1888 (N_1888,In_650,In_167);
nor U1889 (N_1889,In_1332,In_1234);
and U1890 (N_1890,In_286,In_310);
nor U1891 (N_1891,In_1363,In_769);
nor U1892 (N_1892,In_855,In_342);
nand U1893 (N_1893,In_91,In_1706);
nor U1894 (N_1894,In_1773,In_1705);
and U1895 (N_1895,In_1028,In_27);
and U1896 (N_1896,In_1179,In_1307);
xor U1897 (N_1897,In_1546,In_772);
nor U1898 (N_1898,In_434,In_1113);
nand U1899 (N_1899,In_1249,In_655);
nand U1900 (N_1900,In_1036,In_1930);
nor U1901 (N_1901,In_646,In_729);
xnor U1902 (N_1902,In_450,In_1639);
nand U1903 (N_1903,In_821,In_337);
and U1904 (N_1904,In_1150,In_1260);
nor U1905 (N_1905,In_56,In_560);
and U1906 (N_1906,In_537,In_287);
nand U1907 (N_1907,In_1198,In_41);
nor U1908 (N_1908,In_795,In_1740);
or U1909 (N_1909,In_599,In_1155);
or U1910 (N_1910,In_163,In_1862);
and U1911 (N_1911,In_525,In_758);
nor U1912 (N_1912,In_347,In_930);
or U1913 (N_1913,In_302,In_544);
and U1914 (N_1914,In_1261,In_153);
xor U1915 (N_1915,In_304,In_860);
nand U1916 (N_1916,In_753,In_1550);
nand U1917 (N_1917,In_54,In_1444);
or U1918 (N_1918,In_1,In_726);
nand U1919 (N_1919,In_61,In_685);
xor U1920 (N_1920,In_596,In_1986);
or U1921 (N_1921,In_1816,In_806);
and U1922 (N_1922,In_1931,In_461);
xnor U1923 (N_1923,In_447,In_971);
or U1924 (N_1924,In_672,In_166);
nand U1925 (N_1925,In_234,In_1621);
or U1926 (N_1926,In_41,In_813);
nand U1927 (N_1927,In_1354,In_97);
and U1928 (N_1928,In_1695,In_295);
nand U1929 (N_1929,In_1433,In_1254);
and U1930 (N_1930,In_1838,In_1378);
nand U1931 (N_1931,In_992,In_493);
xnor U1932 (N_1932,In_879,In_1861);
or U1933 (N_1933,In_917,In_168);
xnor U1934 (N_1934,In_1417,In_1437);
xnor U1935 (N_1935,In_1799,In_50);
xnor U1936 (N_1936,In_1260,In_268);
or U1937 (N_1937,In_1447,In_1636);
and U1938 (N_1938,In_370,In_1828);
xor U1939 (N_1939,In_522,In_49);
nor U1940 (N_1940,In_1735,In_1304);
xnor U1941 (N_1941,In_1710,In_1943);
nand U1942 (N_1942,In_1650,In_37);
nor U1943 (N_1943,In_662,In_1347);
xnor U1944 (N_1944,In_1660,In_1511);
nor U1945 (N_1945,In_1638,In_519);
nor U1946 (N_1946,In_1564,In_1417);
and U1947 (N_1947,In_471,In_1170);
nand U1948 (N_1948,In_382,In_764);
or U1949 (N_1949,In_1474,In_1882);
nor U1950 (N_1950,In_1575,In_923);
nor U1951 (N_1951,In_771,In_610);
nand U1952 (N_1952,In_1651,In_1906);
nor U1953 (N_1953,In_1704,In_521);
or U1954 (N_1954,In_598,In_190);
and U1955 (N_1955,In_1328,In_1114);
and U1956 (N_1956,In_1942,In_257);
nor U1957 (N_1957,In_537,In_1430);
and U1958 (N_1958,In_1403,In_1721);
and U1959 (N_1959,In_802,In_1116);
and U1960 (N_1960,In_1623,In_210);
and U1961 (N_1961,In_1406,In_1683);
nor U1962 (N_1962,In_1415,In_111);
xor U1963 (N_1963,In_1719,In_1251);
xor U1964 (N_1964,In_1383,In_1592);
nor U1965 (N_1965,In_1401,In_355);
nor U1966 (N_1966,In_1209,In_657);
xor U1967 (N_1967,In_1411,In_1953);
xor U1968 (N_1968,In_660,In_231);
nor U1969 (N_1969,In_1843,In_426);
nand U1970 (N_1970,In_1618,In_162);
and U1971 (N_1971,In_37,In_993);
nand U1972 (N_1972,In_9,In_1621);
and U1973 (N_1973,In_265,In_742);
nor U1974 (N_1974,In_1460,In_260);
and U1975 (N_1975,In_158,In_346);
and U1976 (N_1976,In_1139,In_153);
nor U1977 (N_1977,In_550,In_545);
xor U1978 (N_1978,In_1896,In_1976);
nor U1979 (N_1979,In_407,In_1282);
nor U1980 (N_1980,In_1362,In_1266);
or U1981 (N_1981,In_378,In_1676);
nor U1982 (N_1982,In_1578,In_777);
nand U1983 (N_1983,In_452,In_1386);
nor U1984 (N_1984,In_1992,In_613);
or U1985 (N_1985,In_1057,In_1186);
nor U1986 (N_1986,In_1104,In_277);
and U1987 (N_1987,In_1669,In_287);
and U1988 (N_1988,In_1821,In_1570);
nor U1989 (N_1989,In_1376,In_1842);
nor U1990 (N_1990,In_1356,In_554);
and U1991 (N_1991,In_1836,In_1466);
or U1992 (N_1992,In_462,In_1364);
nor U1993 (N_1993,In_1405,In_254);
or U1994 (N_1994,In_1888,In_1046);
xor U1995 (N_1995,In_270,In_145);
nor U1996 (N_1996,In_144,In_760);
nor U1997 (N_1997,In_1285,In_1679);
nand U1998 (N_1998,In_364,In_72);
and U1999 (N_1999,In_3,In_1613);
or U2000 (N_2000,N_1947,N_1538);
nor U2001 (N_2001,N_1184,N_1842);
and U2002 (N_2002,N_436,N_132);
xnor U2003 (N_2003,N_734,N_210);
xnor U2004 (N_2004,N_205,N_85);
nor U2005 (N_2005,N_74,N_1057);
nand U2006 (N_2006,N_684,N_474);
and U2007 (N_2007,N_1242,N_1784);
nand U2008 (N_2008,N_1767,N_772);
and U2009 (N_2009,N_1011,N_1162);
or U2010 (N_2010,N_1327,N_1083);
xnor U2011 (N_2011,N_1819,N_536);
xor U2012 (N_2012,N_135,N_1892);
and U2013 (N_2013,N_421,N_466);
and U2014 (N_2014,N_1497,N_953);
xnor U2015 (N_2015,N_549,N_1023);
and U2016 (N_2016,N_1448,N_1569);
nand U2017 (N_2017,N_1292,N_219);
nor U2018 (N_2018,N_1293,N_169);
nor U2019 (N_2019,N_996,N_1701);
nor U2020 (N_2020,N_444,N_1085);
and U2021 (N_2021,N_145,N_1194);
nor U2022 (N_2022,N_1126,N_1507);
and U2023 (N_2023,N_921,N_8);
and U2024 (N_2024,N_282,N_1676);
xnor U2025 (N_2025,N_1263,N_1181);
or U2026 (N_2026,N_1522,N_231);
nor U2027 (N_2027,N_284,N_906);
and U2028 (N_2028,N_1319,N_89);
and U2029 (N_2029,N_33,N_491);
nor U2030 (N_2030,N_1291,N_1087);
and U2031 (N_2031,N_1729,N_1749);
xnor U2032 (N_2032,N_1687,N_1314);
xor U2033 (N_2033,N_1330,N_472);
and U2034 (N_2034,N_236,N_27);
xor U2035 (N_2035,N_621,N_301);
nor U2036 (N_2036,N_930,N_1599);
nand U2037 (N_2037,N_1639,N_1220);
or U2038 (N_2038,N_1640,N_983);
or U2039 (N_2039,N_1421,N_887);
xnor U2040 (N_2040,N_702,N_1557);
and U2041 (N_2041,N_1902,N_1080);
xnor U2042 (N_2042,N_1521,N_718);
and U2043 (N_2043,N_1223,N_535);
nand U2044 (N_2044,N_1396,N_1843);
and U2045 (N_2045,N_923,N_1461);
nor U2046 (N_2046,N_753,N_67);
xnor U2047 (N_2047,N_1004,N_526);
nand U2048 (N_2048,N_1799,N_1611);
and U2049 (N_2049,N_489,N_1410);
nand U2050 (N_2050,N_1813,N_959);
nand U2051 (N_2051,N_835,N_192);
nand U2052 (N_2052,N_573,N_1680);
xor U2053 (N_2053,N_1688,N_1341);
nor U2054 (N_2054,N_517,N_409);
nor U2055 (N_2055,N_207,N_1622);
and U2056 (N_2056,N_1822,N_215);
and U2057 (N_2057,N_1187,N_1499);
nand U2058 (N_2058,N_309,N_877);
or U2059 (N_2059,N_1252,N_818);
and U2060 (N_2060,N_643,N_1417);
xor U2061 (N_2061,N_991,N_946);
xnor U2062 (N_2062,N_399,N_945);
nand U2063 (N_2063,N_1980,N_1884);
nor U2064 (N_2064,N_1322,N_1672);
or U2065 (N_2065,N_584,N_1130);
nor U2066 (N_2066,N_1608,N_1667);
and U2067 (N_2067,N_1695,N_1006);
nor U2068 (N_2068,N_555,N_1309);
nor U2069 (N_2069,N_1372,N_668);
and U2070 (N_2070,N_1214,N_63);
or U2071 (N_2071,N_253,N_1562);
nor U2072 (N_2072,N_171,N_1809);
or U2073 (N_2073,N_1794,N_128);
nand U2074 (N_2074,N_1956,N_334);
nor U2075 (N_2075,N_468,N_1266);
and U2076 (N_2076,N_755,N_62);
xnor U2077 (N_2077,N_430,N_1480);
or U2078 (N_2078,N_652,N_1171);
and U2079 (N_2079,N_1549,N_1803);
nand U2080 (N_2080,N_358,N_1906);
or U2081 (N_2081,N_434,N_1566);
and U2082 (N_2082,N_459,N_1312);
and U2083 (N_2083,N_361,N_703);
and U2084 (N_2084,N_800,N_515);
nor U2085 (N_2085,N_412,N_735);
and U2086 (N_2086,N_591,N_1539);
xnor U2087 (N_2087,N_1669,N_1017);
nand U2088 (N_2088,N_669,N_631);
xnor U2089 (N_2089,N_460,N_1240);
and U2090 (N_2090,N_495,N_1359);
nor U2091 (N_2091,N_1712,N_47);
nor U2092 (N_2092,N_408,N_1280);
and U2093 (N_2093,N_1820,N_1283);
nand U2094 (N_2094,N_262,N_342);
and U2095 (N_2095,N_298,N_469);
and U2096 (N_2096,N_752,N_1581);
nand U2097 (N_2097,N_929,N_245);
and U2098 (N_2098,N_1943,N_150);
xor U2099 (N_2099,N_485,N_1917);
xor U2100 (N_2100,N_314,N_1805);
xnor U2101 (N_2101,N_1908,N_498);
nand U2102 (N_2102,N_186,N_281);
nor U2103 (N_2103,N_1501,N_287);
and U2104 (N_2104,N_1453,N_891);
or U2105 (N_2105,N_1626,N_201);
nor U2106 (N_2106,N_1069,N_1321);
nand U2107 (N_2107,N_1300,N_327);
nand U2108 (N_2108,N_1728,N_1972);
and U2109 (N_2109,N_98,N_1132);
or U2110 (N_2110,N_54,N_636);
or U2111 (N_2111,N_1895,N_1962);
xor U2112 (N_2112,N_931,N_968);
nor U2113 (N_2113,N_1733,N_1441);
and U2114 (N_2114,N_994,N_1771);
or U2115 (N_2115,N_825,N_660);
nand U2116 (N_2116,N_689,N_1939);
nand U2117 (N_2117,N_1788,N_698);
nand U2118 (N_2118,N_1936,N_295);
xor U2119 (N_2119,N_1477,N_1624);
or U2120 (N_2120,N_1708,N_280);
nand U2121 (N_2121,N_1419,N_1804);
or U2122 (N_2122,N_263,N_830);
xnor U2123 (N_2123,N_293,N_1028);
nand U2124 (N_2124,N_570,N_502);
nor U2125 (N_2125,N_612,N_1574);
xnor U2126 (N_2126,N_1832,N_1153);
xor U2127 (N_2127,N_1655,N_94);
nor U2128 (N_2128,N_425,N_1550);
nand U2129 (N_2129,N_14,N_764);
and U2130 (N_2130,N_867,N_757);
or U2131 (N_2131,N_1157,N_1847);
nor U2132 (N_2132,N_710,N_1188);
or U2133 (N_2133,N_40,N_813);
nand U2134 (N_2134,N_1617,N_539);
and U2135 (N_2135,N_1165,N_1764);
and U2136 (N_2136,N_1005,N_714);
and U2137 (N_2137,N_101,N_1174);
and U2138 (N_2138,N_1484,N_1509);
xor U2139 (N_2139,N_801,N_1142);
or U2140 (N_2140,N_152,N_1294);
and U2141 (N_2141,N_1664,N_1816);
and U2142 (N_2142,N_1647,N_601);
nand U2143 (N_2143,N_1127,N_878);
xor U2144 (N_2144,N_1871,N_251);
xor U2145 (N_2145,N_908,N_274);
nor U2146 (N_2146,N_597,N_1725);
xor U2147 (N_2147,N_1631,N_695);
xnor U2148 (N_2148,N_1650,N_839);
xnor U2149 (N_2149,N_997,N_939);
and U2150 (N_2150,N_115,N_512);
nor U2151 (N_2151,N_1462,N_1244);
or U2152 (N_2152,N_1913,N_538);
nor U2153 (N_2153,N_1965,N_897);
and U2154 (N_2154,N_1144,N_943);
or U2155 (N_2155,N_1230,N_530);
and U2156 (N_2156,N_1348,N_1536);
and U2157 (N_2157,N_1047,N_427);
nor U2158 (N_2158,N_670,N_645);
or U2159 (N_2159,N_1323,N_879);
and U2160 (N_2160,N_154,N_1976);
or U2161 (N_2161,N_1637,N_1364);
and U2162 (N_2162,N_1973,N_844);
and U2163 (N_2163,N_556,N_1164);
or U2164 (N_2164,N_677,N_1352);
nor U2165 (N_2165,N_911,N_1945);
nor U2166 (N_2166,N_21,N_1675);
nand U2167 (N_2167,N_82,N_691);
nor U2168 (N_2168,N_582,N_1333);
xor U2169 (N_2169,N_1287,N_623);
or U2170 (N_2170,N_1585,N_1155);
or U2171 (N_2171,N_1591,N_1778);
xnor U2172 (N_2172,N_1114,N_1877);
or U2173 (N_2173,N_229,N_849);
nand U2174 (N_2174,N_1265,N_1548);
xnor U2175 (N_2175,N_949,N_671);
or U2176 (N_2176,N_1755,N_1935);
nand U2177 (N_2177,N_1679,N_1);
and U2178 (N_2178,N_365,N_178);
nor U2179 (N_2179,N_1633,N_130);
xnor U2180 (N_2180,N_34,N_1544);
nor U2181 (N_2181,N_833,N_264);
and U2182 (N_2182,N_1800,N_605);
nor U2183 (N_2183,N_1964,N_982);
or U2184 (N_2184,N_1859,N_497);
nor U2185 (N_2185,N_1700,N_1668);
xor U2186 (N_2186,N_1491,N_1339);
or U2187 (N_2187,N_1183,N_1024);
xnor U2188 (N_2188,N_1848,N_1075);
nand U2189 (N_2189,N_45,N_1344);
nand U2190 (N_2190,N_639,N_874);
nor U2191 (N_2191,N_450,N_1185);
and U2192 (N_2192,N_1367,N_1212);
xor U2193 (N_2193,N_276,N_1731);
and U2194 (N_2194,N_1008,N_259);
xnor U2195 (N_2195,N_1059,N_1002);
or U2196 (N_2196,N_1166,N_583);
or U2197 (N_2197,N_1863,N_815);
nand U2198 (N_2198,N_1105,N_824);
xnor U2199 (N_2199,N_1213,N_1559);
xor U2200 (N_2200,N_359,N_329);
and U2201 (N_2201,N_1878,N_315);
and U2202 (N_2202,N_12,N_509);
nor U2203 (N_2203,N_608,N_124);
nor U2204 (N_2204,N_1658,N_374);
nand U2205 (N_2205,N_37,N_1234);
or U2206 (N_2206,N_861,N_36);
and U2207 (N_2207,N_1723,N_1338);
or U2208 (N_2208,N_1691,N_248);
nand U2209 (N_2209,N_1613,N_95);
and U2210 (N_2210,N_795,N_1740);
nor U2211 (N_2211,N_1430,N_449);
and U2212 (N_2212,N_112,N_638);
nand U2213 (N_2213,N_537,N_1278);
nand U2214 (N_2214,N_888,N_222);
or U2215 (N_2215,N_750,N_564);
nor U2216 (N_2216,N_1190,N_125);
nand U2217 (N_2217,N_1385,N_954);
nor U2218 (N_2218,N_1091,N_1850);
nor U2219 (N_2219,N_1122,N_1136);
nand U2220 (N_2220,N_742,N_1706);
and U2221 (N_2221,N_1025,N_1058);
or U2222 (N_2222,N_1853,N_1405);
xor U2223 (N_2223,N_972,N_1587);
xnor U2224 (N_2224,N_1915,N_873);
and U2225 (N_2225,N_1382,N_751);
xor U2226 (N_2226,N_1232,N_72);
nor U2227 (N_2227,N_829,N_257);
nor U2228 (N_2228,N_50,N_307);
nand U2229 (N_2229,N_1420,N_938);
and U2230 (N_2230,N_744,N_736);
xnor U2231 (N_2231,N_1308,N_1032);
xnor U2232 (N_2232,N_181,N_1134);
nor U2233 (N_2233,N_1249,N_1224);
nand U2234 (N_2234,N_914,N_448);
nand U2235 (N_2235,N_807,N_133);
xor U2236 (N_2236,N_1838,N_1137);
or U2237 (N_2237,N_1148,N_1218);
or U2238 (N_2238,N_1227,N_320);
nor U2239 (N_2239,N_1496,N_1034);
or U2240 (N_2240,N_719,N_1851);
xor U2241 (N_2241,N_765,N_1900);
xnor U2242 (N_2242,N_892,N_1152);
nand U2243 (N_2243,N_981,N_1210);
xnor U2244 (N_2244,N_1404,N_1888);
or U2245 (N_2245,N_1773,N_453);
nor U2246 (N_2246,N_1628,N_581);
xnor U2247 (N_2247,N_855,N_603);
nor U2248 (N_2248,N_1845,N_16);
xnor U2249 (N_2249,N_1961,N_19);
nor U2250 (N_2250,N_596,N_1428);
or U2251 (N_2251,N_165,N_470);
nor U2252 (N_2252,N_26,N_1108);
nand U2253 (N_2253,N_1180,N_709);
and U2254 (N_2254,N_872,N_496);
nand U2255 (N_2255,N_1811,N_1135);
nor U2256 (N_2256,N_766,N_768);
nand U2257 (N_2257,N_452,N_1541);
or U2258 (N_2258,N_739,N_1744);
xor U2259 (N_2259,N_506,N_653);
nand U2260 (N_2260,N_1102,N_11);
and U2261 (N_2261,N_1674,N_167);
nand U2262 (N_2262,N_524,N_1128);
nand U2263 (N_2263,N_275,N_1437);
xnor U2264 (N_2264,N_978,N_73);
and U2265 (N_2265,N_79,N_1140);
nor U2266 (N_2266,N_482,N_553);
nor U2267 (N_2267,N_741,N_1609);
nand U2268 (N_2268,N_1960,N_121);
xor U2269 (N_2269,N_534,N_28);
nand U2270 (N_2270,N_1514,N_1802);
nor U2271 (N_2271,N_711,N_1656);
xnor U2272 (N_2272,N_1927,N_797);
nor U2273 (N_2273,N_111,N_679);
xnor U2274 (N_2274,N_883,N_1765);
nand U2275 (N_2275,N_565,N_722);
xnor U2276 (N_2276,N_1296,N_1388);
xnor U2277 (N_2277,N_1746,N_1928);
and U2278 (N_2278,N_1602,N_1350);
and U2279 (N_2279,N_1020,N_1736);
xnor U2280 (N_2280,N_558,N_937);
nand U2281 (N_2281,N_465,N_1243);
and U2282 (N_2282,N_446,N_1791);
nand U2283 (N_2283,N_182,N_893);
nor U2284 (N_2284,N_250,N_1365);
nand U2285 (N_2285,N_1525,N_662);
or U2286 (N_2286,N_410,N_1684);
or U2287 (N_2287,N_1654,N_1762);
or U2288 (N_2288,N_1310,N_965);
nand U2289 (N_2289,N_964,N_1440);
nand U2290 (N_2290,N_1923,N_1955);
or U2291 (N_2291,N_1959,N_1445);
or U2292 (N_2292,N_1376,N_1286);
and U2293 (N_2293,N_723,N_305);
nand U2294 (N_2294,N_1756,N_1763);
nor U2295 (N_2295,N_580,N_235);
nand U2296 (N_2296,N_1416,N_1619);
xor U2297 (N_2297,N_856,N_705);
nand U2298 (N_2298,N_1696,N_832);
nor U2299 (N_2299,N_303,N_649);
xor U2300 (N_2300,N_977,N_1209);
and U2301 (N_2301,N_1573,N_226);
xor U2302 (N_2302,N_337,N_999);
or U2303 (N_2303,N_1486,N_1125);
nand U2304 (N_2304,N_481,N_1439);
xnor U2305 (N_2305,N_778,N_1620);
and U2306 (N_2306,N_940,N_347);
nand U2307 (N_2307,N_1646,N_915);
or U2308 (N_2308,N_454,N_1922);
nand U2309 (N_2309,N_1475,N_1159);
xnor U2310 (N_2310,N_1315,N_58);
nor U2311 (N_2311,N_796,N_304);
nand U2312 (N_2312,N_1449,N_1178);
nor U2313 (N_2313,N_7,N_1035);
xnor U2314 (N_2314,N_858,N_1336);
nor U2315 (N_2315,N_1147,N_487);
xor U2316 (N_2316,N_1413,N_746);
xor U2317 (N_2317,N_1408,N_1123);
nor U2318 (N_2318,N_1219,N_1067);
or U2319 (N_2319,N_1909,N_1977);
or U2320 (N_2320,N_762,N_922);
or U2321 (N_2321,N_1288,N_1552);
xor U2322 (N_2322,N_1916,N_1828);
and U2323 (N_2323,N_1870,N_1891);
nand U2324 (N_2324,N_1070,N_1160);
and U2325 (N_2325,N_1446,N_221);
nand U2326 (N_2326,N_388,N_187);
xnor U2327 (N_2327,N_967,N_868);
and U2328 (N_2328,N_260,N_560);
nor U2329 (N_2329,N_1662,N_1375);
or U2330 (N_2330,N_1096,N_610);
nand U2331 (N_2331,N_149,N_158);
and U2332 (N_2332,N_1663,N_343);
or U2333 (N_2333,N_1919,N_1442);
nor U2334 (N_2334,N_341,N_1095);
and U2335 (N_2335,N_244,N_563);
nor U2336 (N_2336,N_414,N_590);
or U2337 (N_2337,N_1257,N_297);
or U2338 (N_2338,N_1896,N_435);
and U2339 (N_2339,N_1931,N_1279);
or U2340 (N_2340,N_234,N_1607);
xnor U2341 (N_2341,N_1406,N_732);
and U2342 (N_2342,N_1141,N_1215);
xnor U2343 (N_2343,N_831,N_693);
xor U2344 (N_2344,N_172,N_681);
nand U2345 (N_2345,N_974,N_385);
nand U2346 (N_2346,N_606,N_785);
or U2347 (N_2347,N_1389,N_1643);
or U2348 (N_2348,N_1056,N_212);
nor U2349 (N_2349,N_23,N_1920);
and U2350 (N_2350,N_1937,N_386);
nand U2351 (N_2351,N_673,N_932);
and U2352 (N_2352,N_1258,N_1197);
nor U2353 (N_2353,N_439,N_1652);
and U2354 (N_2354,N_1604,N_1303);
or U2355 (N_2355,N_1275,N_6);
or U2356 (N_2356,N_1869,N_352);
and U2357 (N_2357,N_1373,N_1248);
and U2358 (N_2358,N_1211,N_1858);
xnor U2359 (N_2359,N_696,N_655);
nand U2360 (N_2360,N_189,N_1206);
or U2361 (N_2361,N_958,N_697);
and U2362 (N_2362,N_242,N_1553);
nand U2363 (N_2363,N_1129,N_1738);
nor U2364 (N_2364,N_1576,N_1447);
nor U2365 (N_2365,N_389,N_475);
and U2366 (N_2366,N_22,N_1101);
and U2367 (N_2367,N_733,N_864);
nor U2368 (N_2368,N_1689,N_1259);
or U2369 (N_2369,N_339,N_1360);
nor U2370 (N_2370,N_700,N_973);
or U2371 (N_2371,N_398,N_65);
or U2372 (N_2372,N_381,N_18);
nand U2373 (N_2373,N_1526,N_1578);
xnor U2374 (N_2374,N_1739,N_87);
or U2375 (N_2375,N_781,N_1781);
or U2376 (N_2376,N_1632,N_1716);
nor U2377 (N_2377,N_947,N_379);
nor U2378 (N_2378,N_191,N_1175);
nor U2379 (N_2379,N_1084,N_1898);
nor U2380 (N_2380,N_935,N_1887);
nor U2381 (N_2381,N_300,N_882);
and U2382 (N_2382,N_1511,N_745);
xor U2383 (N_2383,N_1660,N_1495);
and U2384 (N_2384,N_531,N_1750);
xnor U2385 (N_2385,N_1369,N_1683);
and U2386 (N_2386,N_758,N_155);
nor U2387 (N_2387,N_426,N_1670);
nand U2388 (N_2388,N_1748,N_55);
or U2389 (N_2389,N_1795,N_1349);
and U2390 (N_2390,N_1216,N_321);
xnor U2391 (N_2391,N_1653,N_637);
xnor U2392 (N_2392,N_139,N_1598);
xnor U2393 (N_2393,N_1422,N_90);
xnor U2394 (N_2394,N_620,N_477);
xor U2395 (N_2395,N_1595,N_258);
nor U2396 (N_2396,N_917,N_1580);
nand U2397 (N_2397,N_69,N_1313);
or U2398 (N_2398,N_1434,N_979);
nor U2399 (N_2399,N_391,N_86);
nor U2400 (N_2400,N_195,N_1182);
and U2401 (N_2401,N_1474,N_1779);
nand U2402 (N_2402,N_1009,N_516);
and U2403 (N_2403,N_1985,N_646);
xnor U2404 (N_2404,N_395,N_1946);
and U2405 (N_2405,N_1872,N_756);
xnor U2406 (N_2406,N_328,N_862);
or U2407 (N_2407,N_1718,N_318);
or U2408 (N_2408,N_518,N_486);
and U2409 (N_2409,N_1110,N_1456);
xor U2410 (N_2410,N_1205,N_1370);
and U2411 (N_2411,N_1233,N_992);
xnor U2412 (N_2412,N_360,N_159);
or U2413 (N_2413,N_349,N_376);
and U2414 (N_2414,N_476,N_272);
nor U2415 (N_2415,N_607,N_134);
or U2416 (N_2416,N_206,N_179);
nor U2417 (N_2417,N_1302,N_420);
or U2418 (N_2418,N_729,N_1217);
or U2419 (N_2419,N_204,N_622);
xnor U2420 (N_2420,N_1307,N_1563);
nand U2421 (N_2421,N_1697,N_1742);
or U2422 (N_2422,N_1347,N_1827);
nor U2423 (N_2423,N_1846,N_310);
nor U2424 (N_2424,N_1013,N_323);
nand U2425 (N_2425,N_907,N_117);
and U2426 (N_2426,N_782,N_568);
nor U2427 (N_2427,N_404,N_820);
or U2428 (N_2428,N_1311,N_102);
nand U2429 (N_2429,N_851,N_1390);
and U2430 (N_2430,N_285,N_609);
xnor U2431 (N_2431,N_805,N_1362);
xor U2432 (N_2432,N_925,N_4);
nor U2433 (N_2433,N_579,N_1045);
and U2434 (N_2434,N_642,N_1203);
and U2435 (N_2435,N_1247,N_471);
xnor U2436 (N_2436,N_1316,N_1777);
and U2437 (N_2437,N_146,N_198);
or U2438 (N_2438,N_418,N_969);
and U2439 (N_2439,N_748,N_898);
nor U2440 (N_2440,N_961,N_1940);
and U2441 (N_2441,N_396,N_1849);
and U2442 (N_2442,N_1671,N_1571);
or U2443 (N_2443,N_483,N_811);
xor U2444 (N_2444,N_1699,N_103);
and U2445 (N_2445,N_1910,N_432);
and U2446 (N_2446,N_1320,N_1354);
and U2447 (N_2447,N_168,N_875);
and U2448 (N_2448,N_1177,N_611);
nor U2449 (N_2449,N_177,N_1812);
nand U2450 (N_2450,N_1455,N_1899);
or U2451 (N_2451,N_966,N_1570);
xor U2452 (N_2452,N_1596,N_927);
and U2453 (N_2453,N_1473,N_1545);
or U2454 (N_2454,N_208,N_626);
xor U2455 (N_2455,N_268,N_1926);
xor U2456 (N_2456,N_1090,N_896);
nor U2457 (N_2457,N_116,N_598);
nand U2458 (N_2458,N_1368,N_451);
nor U2459 (N_2459,N_895,N_827);
or U2460 (N_2460,N_241,N_1156);
or U2461 (N_2461,N_715,N_869);
nor U2462 (N_2462,N_1237,N_447);
nor U2463 (N_2463,N_1340,N_237);
xor U2464 (N_2464,N_663,N_213);
or U2465 (N_2465,N_1997,N_716);
nor U2466 (N_2466,N_1146,N_1060);
nor U2467 (N_2467,N_865,N_1904);
nor U2468 (N_2468,N_1659,N_1239);
nand U2469 (N_2469,N_249,N_157);
or U2470 (N_2470,N_1066,N_1111);
xor U2471 (N_2471,N_1505,N_1470);
nor U2472 (N_2472,N_76,N_1431);
and U2473 (N_2473,N_1094,N_1415);
or U2474 (N_2474,N_971,N_107);
nand U2475 (N_2475,N_202,N_789);
and U2476 (N_2476,N_325,N_1759);
xor U2477 (N_2477,N_1698,N_787);
nand U2478 (N_2478,N_1981,N_1010);
xor U2479 (N_2479,N_1577,N_1054);
and U2480 (N_2480,N_239,N_1107);
xnor U2481 (N_2481,N_1254,N_75);
xnor U2482 (N_2482,N_542,N_1030);
or U2483 (N_2483,N_488,N_1506);
and U2484 (N_2484,N_1709,N_1493);
xor U2485 (N_2485,N_1423,N_1579);
or U2486 (N_2486,N_1014,N_1821);
xor U2487 (N_2487,N_1774,N_1436);
and U2488 (N_2488,N_1754,N_5);
nand U2489 (N_2489,N_113,N_143);
and U2490 (N_2490,N_554,N_1605);
and U2491 (N_2491,N_1284,N_763);
and U2492 (N_2492,N_1377,N_233);
and U2493 (N_2493,N_1610,N_687);
nand U2494 (N_2494,N_1086,N_504);
nor U2495 (N_2495,N_578,N_1196);
nor U2496 (N_2496,N_1988,N_1814);
or U2497 (N_2497,N_217,N_1371);
and U2498 (N_2498,N_1905,N_1715);
and U2499 (N_2499,N_1963,N_885);
nand U2500 (N_2500,N_173,N_1554);
nor U2501 (N_2501,N_53,N_513);
and U2502 (N_2502,N_546,N_1494);
xnor U2503 (N_2503,N_559,N_1515);
nand U2504 (N_2504,N_1753,N_920);
xor U2505 (N_2505,N_599,N_951);
or U2506 (N_2506,N_1588,N_356);
or U2507 (N_2507,N_1702,N_100);
and U2508 (N_2508,N_1537,N_199);
nand U2509 (N_2509,N_1238,N_225);
nand U2510 (N_2510,N_1776,N_1261);
and U2511 (N_2511,N_256,N_1704);
and U2512 (N_2512,N_289,N_462);
xnor U2513 (N_2513,N_1524,N_1785);
and U2514 (N_2514,N_792,N_948);
xnor U2515 (N_2515,N_592,N_1407);
xor U2516 (N_2516,N_790,N_1864);
and U2517 (N_2517,N_1386,N_375);
nor U2518 (N_2518,N_1685,N_1876);
and U2519 (N_2519,N_680,N_1167);
and U2520 (N_2520,N_440,N_1944);
nand U2521 (N_2521,N_569,N_1881);
xnor U2522 (N_2522,N_43,N_333);
nor U2523 (N_2523,N_1374,N_1780);
or U2524 (N_2524,N_387,N_1115);
xor U2525 (N_2525,N_615,N_1564);
or U2526 (N_2526,N_99,N_1498);
or U2527 (N_2527,N_998,N_706);
or U2528 (N_2528,N_1714,N_905);
xnor U2529 (N_2529,N_1173,N_1169);
nand U2530 (N_2530,N_1277,N_1615);
nand U2531 (N_2531,N_480,N_644);
nand U2532 (N_2532,N_952,N_161);
nand U2533 (N_2533,N_1666,N_902);
xnor U2534 (N_2534,N_269,N_1022);
and U2535 (N_2535,N_984,N_871);
nand U2536 (N_2536,N_39,N_137);
and U2537 (N_2537,N_1970,N_988);
xor U2538 (N_2538,N_218,N_1427);
or U2539 (N_2539,N_1966,N_1299);
and U2540 (N_2540,N_628,N_1616);
xnor U2541 (N_2541,N_1366,N_42);
nor U2542 (N_2542,N_1317,N_1189);
xor U2543 (N_2543,N_313,N_793);
nand U2544 (N_2544,N_841,N_1730);
and U2545 (N_2545,N_316,N_846);
or U2546 (N_2546,N_1414,N_788);
nand U2547 (N_2547,N_666,N_1328);
nor U2548 (N_2548,N_493,N_1527);
xnor U2549 (N_2549,N_1276,N_25);
nand U2550 (N_2550,N_816,N_290);
nor U2551 (N_2551,N_1852,N_164);
nor U2552 (N_2552,N_1454,N_525);
nand U2553 (N_2553,N_336,N_311);
xnor U2554 (N_2554,N_1357,N_1271);
nand U2555 (N_2555,N_230,N_1384);
nand U2556 (N_2556,N_1121,N_13);
nor U2557 (N_2557,N_1953,N_151);
nor U2558 (N_2558,N_1590,N_1297);
and U2559 (N_2559,N_1879,N_1270);
xor U2560 (N_2560,N_1429,N_60);
and U2561 (N_2561,N_1079,N_340);
nand U2562 (N_2562,N_848,N_1179);
nor U2563 (N_2563,N_1465,N_747);
xor U2564 (N_2564,N_378,N_1775);
nor U2565 (N_2565,N_355,N_1099);
and U2566 (N_2566,N_1516,N_1737);
or U2567 (N_2567,N_1840,N_674);
or U2568 (N_2568,N_1751,N_1957);
nor U2569 (N_2569,N_1950,N_614);
nor U2570 (N_2570,N_1335,N_975);
nor U2571 (N_2571,N_769,N_1503);
nand U2572 (N_2572,N_624,N_129);
and U2573 (N_2573,N_544,N_717);
and U2574 (N_2574,N_1041,N_9);
or U2575 (N_2575,N_1508,N_24);
nand U2576 (N_2576,N_255,N_1792);
and U2577 (N_2577,N_411,N_59);
and U2578 (N_2578,N_174,N_1758);
and U2579 (N_2579,N_1063,N_1071);
nand U2580 (N_2580,N_1594,N_148);
xor U2581 (N_2581,N_1855,N_692);
nand U2582 (N_2582,N_458,N_803);
nor U2583 (N_2583,N_88,N_220);
and U2584 (N_2584,N_604,N_1593);
nand U2585 (N_2585,N_837,N_286);
xor U2586 (N_2586,N_322,N_203);
nor U2587 (N_2587,N_1500,N_1381);
nand U2588 (N_2588,N_791,N_1479);
nand U2589 (N_2589,N_812,N_901);
xnor U2590 (N_2590,N_1065,N_185);
nor U2591 (N_2591,N_1575,N_587);
xor U2592 (N_2592,N_97,N_550);
nand U2593 (N_2593,N_909,N_1889);
nor U2594 (N_2594,N_492,N_1100);
or U2595 (N_2595,N_728,N_1991);
and U2596 (N_2596,N_400,N_783);
xor U2597 (N_2597,N_1068,N_3);
xor U2598 (N_2598,N_1831,N_990);
or U2599 (N_2599,N_1395,N_1458);
and U2600 (N_2600,N_1150,N_1555);
nor U2601 (N_2601,N_989,N_1029);
nand U2602 (N_2602,N_1875,N_1411);
and U2603 (N_2603,N_804,N_1629);
nor U2604 (N_2604,N_588,N_678);
and U2605 (N_2605,N_1268,N_122);
xor U2606 (N_2606,N_1361,N_1409);
xnor U2607 (N_2607,N_1761,N_1546);
and U2608 (N_2608,N_1513,N_1894);
and U2609 (N_2609,N_886,N_1170);
xnor U2610 (N_2610,N_1636,N_523);
nor U2611 (N_2611,N_1686,N_1865);
nand U2612 (N_2612,N_522,N_1661);
nand U2613 (N_2613,N_648,N_478);
or U2614 (N_2614,N_1993,N_1112);
or U2615 (N_2615,N_131,N_1138);
xnor U2616 (N_2616,N_1012,N_1443);
xor U2617 (N_2617,N_1383,N_1710);
nand U2618 (N_2618,N_654,N_903);
nor U2619 (N_2619,N_330,N_1567);
nor U2620 (N_2620,N_1492,N_853);
or U2621 (N_2621,N_51,N_708);
and U2622 (N_2622,N_918,N_1088);
nor U2623 (N_2623,N_1472,N_726);
xor U2624 (N_2624,N_431,N_1235);
xor U2625 (N_2625,N_1880,N_1403);
or U2626 (N_2626,N_288,N_1379);
or U2627 (N_2627,N_1734,N_1064);
xnor U2628 (N_2628,N_57,N_380);
or U2629 (N_2629,N_1825,N_278);
nor U2630 (N_2630,N_1866,N_1269);
nand U2631 (N_2631,N_1721,N_657);
or U2632 (N_2632,N_392,N_780);
or U2633 (N_2633,N_66,N_1623);
and U2634 (N_2634,N_308,N_1113);
nand U2635 (N_2635,N_357,N_1703);
and U2636 (N_2636,N_1724,N_302);
xnor U2637 (N_2637,N_1817,N_1600);
nor U2638 (N_2638,N_338,N_913);
nor U2639 (N_2639,N_1092,N_1798);
xnor U2640 (N_2640,N_616,N_1830);
xor U2641 (N_2641,N_1984,N_428);
nor U2642 (N_2642,N_1195,N_1039);
nor U2643 (N_2643,N_720,N_600);
nand U2644 (N_2644,N_211,N_299);
and U2645 (N_2645,N_188,N_1941);
nor U2646 (N_2646,N_889,N_312);
and U2647 (N_2647,N_1044,N_1131);
and U2648 (N_2648,N_1531,N_1163);
xor U2649 (N_2649,N_1606,N_156);
xor U2650 (N_2650,N_1951,N_618);
or U2651 (N_2651,N_1603,N_1727);
nand U2652 (N_2652,N_986,N_423);
xnor U2653 (N_2653,N_941,N_699);
and U2654 (N_2654,N_438,N_919);
nand U2655 (N_2655,N_1118,N_725);
and U2656 (N_2656,N_1886,N_1690);
nor U2657 (N_2657,N_1996,N_348);
nor U2658 (N_2658,N_1907,N_1073);
and U2659 (N_2659,N_650,N_1986);
nor U2660 (N_2660,N_1289,N_1665);
nor U2661 (N_2661,N_704,N_508);
nor U2662 (N_2662,N_1186,N_324);
nand U2663 (N_2663,N_1285,N_1459);
and U2664 (N_2664,N_1914,N_774);
and U2665 (N_2665,N_1228,N_162);
nand U2666 (N_2666,N_296,N_1222);
nand U2667 (N_2667,N_1089,N_1720);
or U2668 (N_2668,N_1231,N_1717);
xor U2669 (N_2669,N_552,N_1104);
nor U2670 (N_2670,N_511,N_1452);
and U2671 (N_2671,N_1274,N_821);
or U2672 (N_2672,N_730,N_1324);
and U2673 (N_2673,N_1867,N_1050);
nand U2674 (N_2674,N_1363,N_17);
or U2675 (N_2675,N_214,N_1295);
or U2676 (N_2676,N_860,N_586);
nor U2677 (N_2677,N_1489,N_1201);
nor U2678 (N_2678,N_1597,N_955);
xor U2679 (N_2679,N_1673,N_283);
and U2680 (N_2680,N_1331,N_1797);
nor U2681 (N_2681,N_1994,N_589);
nor U2682 (N_2682,N_479,N_1768);
nand U2683 (N_2683,N_1948,N_1399);
or U2684 (N_2684,N_292,N_1974);
nand U2685 (N_2685,N_331,N_1560);
nand U2686 (N_2686,N_870,N_933);
or U2687 (N_2687,N_1808,N_640);
and U2688 (N_2688,N_880,N_1969);
nor U2689 (N_2689,N_1769,N_1529);
and U2690 (N_2690,N_433,N_20);
xnor U2691 (N_2691,N_779,N_463);
or U2692 (N_2692,N_993,N_1540);
nor U2693 (N_2693,N_1868,N_843);
xor U2694 (N_2694,N_521,N_494);
or U2695 (N_2695,N_1635,N_619);
xnor U2696 (N_2696,N_576,N_273);
xnor U2697 (N_2697,N_382,N_1893);
and U2698 (N_2698,N_1829,N_442);
xor U2699 (N_2699,N_547,N_183);
or U2700 (N_2700,N_894,N_1468);
nand U2701 (N_2701,N_1512,N_1649);
nand U2702 (N_2702,N_291,N_1478);
nand U2703 (N_2703,N_1942,N_936);
or U2704 (N_2704,N_770,N_859);
and U2705 (N_2705,N_1031,N_574);
or U2706 (N_2706,N_1707,N_876);
and U2707 (N_2707,N_1547,N_345);
and U2708 (N_2708,N_1933,N_1055);
and U2709 (N_2709,N_1490,N_175);
and U2710 (N_2710,N_1971,N_1770);
nand U2711 (N_2711,N_635,N_548);
nand U2712 (N_2712,N_1229,N_890);
xor U2713 (N_2713,N_985,N_667);
nand U2714 (N_2714,N_1949,N_659);
and U2715 (N_2715,N_144,N_585);
nor U2716 (N_2716,N_1398,N_802);
xor U2717 (N_2717,N_1823,N_1103);
nor U2718 (N_2718,N_1202,N_294);
xnor U2719 (N_2719,N_81,N_1983);
and U2720 (N_2720,N_1151,N_83);
nor U2721 (N_2721,N_528,N_270);
xnor U2722 (N_2722,N_545,N_1987);
and U2723 (N_2723,N_1760,N_625);
or U2724 (N_2724,N_928,N_176);
or U2725 (N_2725,N_1968,N_532);
and U2726 (N_2726,N_1938,N_1925);
xnor U2727 (N_2727,N_1337,N_647);
nand U2728 (N_2728,N_1345,N_519);
nor U2729 (N_2729,N_1614,N_737);
xor U2730 (N_2730,N_1199,N_1262);
and U2731 (N_2731,N_633,N_456);
nand U2732 (N_2732,N_56,N_277);
nor U2733 (N_2733,N_520,N_956);
nand U2734 (N_2734,N_1520,N_1790);
and U2735 (N_2735,N_1358,N_368);
nand U2736 (N_2736,N_1425,N_160);
and U2737 (N_2737,N_784,N_845);
nor U2738 (N_2738,N_490,N_963);
nor U2739 (N_2739,N_369,N_529);
nand U2740 (N_2740,N_1584,N_1168);
and U2741 (N_2741,N_962,N_1051);
nor U2742 (N_2742,N_1149,N_1824);
and U2743 (N_2743,N_142,N_806);
or U2744 (N_2744,N_507,N_406);
xor U2745 (N_2745,N_1193,N_1517);
and U2746 (N_2746,N_819,N_31);
nand U2747 (N_2747,N_197,N_394);
nand U2748 (N_2748,N_995,N_126);
nor U2749 (N_2749,N_1967,N_1583);
or U2750 (N_2750,N_857,N_1958);
xnor U2751 (N_2751,N_422,N_1326);
xor U2752 (N_2752,N_1934,N_319);
or U2753 (N_2753,N_1464,N_786);
xnor U2754 (N_2754,N_190,N_571);
nor U2755 (N_2755,N_1979,N_1978);
or U2756 (N_2756,N_724,N_1952);
xnor U2757 (N_2757,N_840,N_767);
nand U2758 (N_2758,N_838,N_665);
nand U2759 (N_2759,N_49,N_541);
or U2760 (N_2760,N_1975,N_1836);
xor U2761 (N_2761,N_279,N_1191);
and U2762 (N_2762,N_1139,N_46);
nor U2763 (N_2763,N_180,N_1841);
nor U2764 (N_2764,N_1911,N_1003);
nand U2765 (N_2765,N_1722,N_924);
nand U2766 (N_2766,N_1355,N_1873);
nand U2767 (N_2767,N_1677,N_1510);
and U2768 (N_2768,N_363,N_731);
xnor U2769 (N_2769,N_850,N_1634);
or U2770 (N_2770,N_1329,N_1154);
xnor U2771 (N_2771,N_1789,N_1380);
xor U2772 (N_2772,N_1402,N_1857);
and U2773 (N_2773,N_777,N_1450);
nor U2774 (N_2774,N_243,N_401);
nand U2775 (N_2775,N_1565,N_1543);
and U2776 (N_2776,N_685,N_759);
nor U2777 (N_2777,N_32,N_740);
xnor U2778 (N_2778,N_1882,N_1741);
nor U2779 (N_2779,N_1078,N_93);
xnor U2780 (N_2780,N_1158,N_900);
or U2781 (N_2781,N_712,N_127);
xor U2782 (N_2782,N_1693,N_346);
nand U2783 (N_2783,N_572,N_1460);
nand U2784 (N_2784,N_1834,N_1394);
nor U2785 (N_2785,N_1048,N_1612);
xor U2786 (N_2786,N_445,N_1267);
or U2787 (N_2787,N_372,N_1120);
nand U2788 (N_2788,N_630,N_817);
nor U2789 (N_2789,N_1124,N_1883);
or U2790 (N_2790,N_760,N_1890);
nand U2791 (N_2791,N_1786,N_1082);
or U2792 (N_2792,N_1097,N_1061);
xnor U2793 (N_2793,N_92,N_1982);
and U2794 (N_2794,N_1412,N_1535);
nand U2795 (N_2795,N_1255,N_415);
xor U2796 (N_2796,N_473,N_441);
xor U2797 (N_2797,N_863,N_166);
nand U2798 (N_2798,N_694,N_1998);
nand U2799 (N_2799,N_1176,N_1225);
nand U2800 (N_2800,N_1844,N_384);
or U2801 (N_2801,N_505,N_1648);
nand U2802 (N_2802,N_1485,N_960);
xor U2803 (N_2803,N_1192,N_271);
and U2804 (N_2804,N_934,N_1815);
xnor U2805 (N_2805,N_1007,N_1989);
nor U2806 (N_2806,N_106,N_1999);
and U2807 (N_2807,N_119,N_266);
xor U2808 (N_2808,N_1351,N_1040);
xor U2809 (N_2809,N_794,N_775);
nand U2810 (N_2810,N_1807,N_1332);
nor U2811 (N_2811,N_1469,N_834);
xor U2812 (N_2812,N_1618,N_1856);
or U2813 (N_2813,N_1990,N_809);
or U2814 (N_2814,N_140,N_84);
nor U2815 (N_2815,N_1837,N_1644);
nor U2816 (N_2816,N_1657,N_814);
nor U2817 (N_2817,N_836,N_503);
or U2818 (N_2818,N_543,N_1874);
xor U2819 (N_2819,N_1504,N_80);
and U2820 (N_2820,N_1053,N_527);
and U2821 (N_2821,N_1995,N_602);
or U2822 (N_2822,N_1476,N_1074);
and U2823 (N_2823,N_354,N_1826);
or U2824 (N_2824,N_464,N_1260);
and U2825 (N_2825,N_1133,N_1627);
nand U2826 (N_2826,N_682,N_1833);
nor U2827 (N_2827,N_1901,N_402);
nor U2828 (N_2828,N_1204,N_247);
and U2829 (N_2829,N_557,N_899);
or U2830 (N_2830,N_96,N_1273);
and U2831 (N_2831,N_1783,N_1451);
nor U2832 (N_2832,N_1793,N_1488);
nand U2833 (N_2833,N_64,N_118);
xnor U2834 (N_2834,N_904,N_196);
or U2835 (N_2835,N_1854,N_1921);
and U2836 (N_2836,N_1502,N_1281);
and U2837 (N_2837,N_417,N_823);
or U2838 (N_2838,N_1897,N_594);
and U2839 (N_2839,N_1713,N_1481);
nor U2840 (N_2840,N_170,N_1787);
xnor U2841 (N_2841,N_61,N_1912);
or U2842 (N_2842,N_629,N_1641);
and U2843 (N_2843,N_44,N_123);
nand U2844 (N_2844,N_1251,N_828);
nor U2845 (N_2845,N_1198,N_866);
and U2846 (N_2846,N_91,N_826);
nor U2847 (N_2847,N_1630,N_1726);
nor U2848 (N_2848,N_1444,N_593);
or U2849 (N_2849,N_1471,N_942);
xor U2850 (N_2850,N_1528,N_1642);
and U2851 (N_2851,N_1757,N_661);
nand U2852 (N_2852,N_1076,N_1860);
xor U2853 (N_2853,N_1052,N_1586);
or U2854 (N_2854,N_771,N_500);
nand U2855 (N_2855,N_656,N_424);
and U2856 (N_2856,N_727,N_443);
nor U2857 (N_2857,N_1172,N_1016);
or U2858 (N_2858,N_373,N_163);
and U2859 (N_2859,N_1743,N_1625);
and U2860 (N_2860,N_377,N_1342);
nand U2861 (N_2861,N_1226,N_847);
nand U2862 (N_2862,N_595,N_1221);
xor U2863 (N_2863,N_1861,N_1796);
xor U2864 (N_2864,N_1924,N_1397);
xor U2865 (N_2865,N_153,N_881);
nor U2866 (N_2866,N_252,N_30);
nand U2867 (N_2867,N_808,N_1918);
nor U2868 (N_2868,N_1015,N_1046);
nor U2869 (N_2869,N_1835,N_1601);
xnor U2870 (N_2870,N_1519,N_743);
nor U2871 (N_2871,N_77,N_916);
nand U2872 (N_2872,N_109,N_617);
nor U2873 (N_2873,N_1558,N_810);
nor U2874 (N_2874,N_749,N_754);
nor U2875 (N_2875,N_200,N_147);
and U2876 (N_2876,N_1457,N_232);
or U2877 (N_2877,N_238,N_690);
and U2878 (N_2878,N_1143,N_1810);
nor U2879 (N_2879,N_1885,N_267);
and U2880 (N_2880,N_78,N_1272);
nand U2881 (N_2881,N_1438,N_223);
xor U2882 (N_2882,N_1236,N_798);
and U2883 (N_2883,N_1747,N_1036);
xor U2884 (N_2884,N_1119,N_429);
nand U2885 (N_2885,N_701,N_1033);
nor U2886 (N_2886,N_353,N_1038);
nor U2887 (N_2887,N_926,N_0);
xor U2888 (N_2888,N_68,N_403);
nor U2889 (N_2889,N_1589,N_551);
nand U2890 (N_2890,N_1200,N_567);
nor U2891 (N_2891,N_738,N_664);
and U2892 (N_2892,N_1530,N_1534);
and U2893 (N_2893,N_397,N_1245);
nor U2894 (N_2894,N_683,N_38);
nor U2895 (N_2895,N_265,N_1435);
or U2896 (N_2896,N_976,N_437);
xnor U2897 (N_2897,N_1772,N_29);
nand U2898 (N_2898,N_1021,N_713);
nand U2899 (N_2899,N_371,N_110);
nor U2900 (N_2900,N_1930,N_1264);
nand U2901 (N_2901,N_1424,N_370);
nand U2902 (N_2902,N_1839,N_634);
xnor U2903 (N_2903,N_1711,N_484);
and U2904 (N_2904,N_675,N_1019);
xnor U2905 (N_2905,N_688,N_108);
nor U2906 (N_2906,N_1433,N_1694);
xnor U2907 (N_2907,N_1145,N_1745);
or U2908 (N_2908,N_970,N_912);
nand U2909 (N_2909,N_1645,N_1719);
and U2910 (N_2910,N_686,N_194);
or U2911 (N_2911,N_1042,N_261);
nand U2912 (N_2912,N_707,N_1542);
or U2913 (N_2913,N_980,N_71);
or U2914 (N_2914,N_1098,N_114);
and U2915 (N_2915,N_1378,N_910);
nand U2916 (N_2916,N_1561,N_2);
and U2917 (N_2917,N_1027,N_467);
nand U2918 (N_2918,N_48,N_1077);
xnor U2919 (N_2919,N_350,N_1568);
and U2920 (N_2920,N_367,N_658);
nand U2921 (N_2921,N_1401,N_1256);
xor U2922 (N_2922,N_1692,N_351);
nand U2923 (N_2923,N_70,N_15);
nand U2924 (N_2924,N_501,N_1318);
or U2925 (N_2925,N_240,N_216);
xnor U2926 (N_2926,N_1426,N_1732);
or U2927 (N_2927,N_1638,N_184);
or U2928 (N_2928,N_613,N_1681);
and U2929 (N_2929,N_1735,N_390);
nor U2930 (N_2930,N_1109,N_1026);
or U2931 (N_2931,N_52,N_407);
or U2932 (N_2932,N_1282,N_246);
xnor U2933 (N_2933,N_944,N_761);
or U2934 (N_2934,N_641,N_627);
and U2935 (N_2935,N_120,N_254);
nor U2936 (N_2936,N_1001,N_1072);
nand U2937 (N_2937,N_1093,N_393);
xor U2938 (N_2938,N_1592,N_1766);
and U2939 (N_2939,N_1306,N_1049);
nand U2940 (N_2940,N_455,N_1678);
or U2941 (N_2941,N_852,N_138);
xor U2942 (N_2942,N_514,N_822);
nor U2943 (N_2943,N_1393,N_1551);
xnor U2944 (N_2944,N_842,N_104);
or U2945 (N_2945,N_1705,N_1290);
xor U2946 (N_2946,N_561,N_364);
or U2947 (N_2947,N_1621,N_35);
and U2948 (N_2948,N_499,N_672);
or U2949 (N_2949,N_1518,N_1325);
and U2950 (N_2950,N_1353,N_1391);
nand U2951 (N_2951,N_1043,N_344);
and U2952 (N_2952,N_1387,N_141);
xnor U2953 (N_2953,N_228,N_1992);
nor U2954 (N_2954,N_457,N_510);
and U2955 (N_2955,N_957,N_1932);
and U2956 (N_2956,N_799,N_1356);
xnor U2957 (N_2957,N_1018,N_1482);
nand U2958 (N_2958,N_1466,N_1400);
and U2959 (N_2959,N_854,N_1903);
nor U2960 (N_2960,N_1343,N_1463);
xnor U2961 (N_2961,N_306,N_461);
nor U2962 (N_2962,N_632,N_1533);
and U2963 (N_2963,N_1106,N_1862);
xnor U2964 (N_2964,N_1682,N_332);
and U2965 (N_2965,N_105,N_419);
xor U2966 (N_2966,N_41,N_566);
nor U2967 (N_2967,N_1556,N_533);
or U2968 (N_2968,N_405,N_1305);
and U2969 (N_2969,N_1418,N_1483);
and U2970 (N_2970,N_776,N_1582);
xnor U2971 (N_2971,N_1116,N_562);
nand U2972 (N_2972,N_193,N_1161);
nand U2973 (N_2973,N_676,N_1062);
and U2974 (N_2974,N_1651,N_1346);
and U2975 (N_2975,N_1523,N_1487);
and U2976 (N_2976,N_1250,N_950);
xnor U2977 (N_2977,N_1037,N_540);
nand U2978 (N_2978,N_987,N_1253);
xnor U2979 (N_2979,N_383,N_10);
xor U2980 (N_2980,N_362,N_773);
or U2981 (N_2981,N_884,N_1246);
nor U2982 (N_2982,N_335,N_1532);
and U2983 (N_2983,N_1301,N_224);
nor U2984 (N_2984,N_326,N_1207);
and U2985 (N_2985,N_1117,N_1467);
nor U2986 (N_2986,N_1304,N_1208);
nand U2987 (N_2987,N_366,N_1000);
or U2988 (N_2988,N_577,N_721);
nand U2989 (N_2989,N_1392,N_416);
xor U2990 (N_2990,N_651,N_1929);
and U2991 (N_2991,N_1954,N_1298);
nand U2992 (N_2992,N_575,N_227);
nor U2993 (N_2993,N_1334,N_136);
nor U2994 (N_2994,N_209,N_1806);
nand U2995 (N_2995,N_1801,N_1752);
or U2996 (N_2996,N_1572,N_1432);
nand U2997 (N_2997,N_317,N_413);
and U2998 (N_2998,N_1782,N_1241);
or U2999 (N_2999,N_1081,N_1818);
or U3000 (N_3000,N_577,N_209);
nor U3001 (N_3001,N_1455,N_1537);
and U3002 (N_3002,N_1449,N_327);
or U3003 (N_3003,N_899,N_1617);
xnor U3004 (N_3004,N_1415,N_552);
or U3005 (N_3005,N_1222,N_1857);
or U3006 (N_3006,N_159,N_1288);
nor U3007 (N_3007,N_1189,N_1977);
nand U3008 (N_3008,N_585,N_1871);
and U3009 (N_3009,N_1555,N_951);
and U3010 (N_3010,N_1216,N_42);
or U3011 (N_3011,N_38,N_404);
nor U3012 (N_3012,N_1240,N_1525);
nand U3013 (N_3013,N_1080,N_1197);
nand U3014 (N_3014,N_44,N_65);
or U3015 (N_3015,N_1077,N_26);
and U3016 (N_3016,N_1277,N_1120);
and U3017 (N_3017,N_821,N_1050);
xnor U3018 (N_3018,N_323,N_593);
nand U3019 (N_3019,N_1942,N_884);
nor U3020 (N_3020,N_357,N_354);
xnor U3021 (N_3021,N_989,N_454);
and U3022 (N_3022,N_1767,N_1550);
xor U3023 (N_3023,N_468,N_1835);
or U3024 (N_3024,N_1307,N_1153);
or U3025 (N_3025,N_1313,N_410);
and U3026 (N_3026,N_1076,N_983);
xor U3027 (N_3027,N_5,N_1891);
nor U3028 (N_3028,N_1859,N_393);
or U3029 (N_3029,N_1961,N_1759);
or U3030 (N_3030,N_258,N_1658);
and U3031 (N_3031,N_1813,N_1786);
nor U3032 (N_3032,N_358,N_1503);
or U3033 (N_3033,N_951,N_103);
xnor U3034 (N_3034,N_311,N_279);
nor U3035 (N_3035,N_1033,N_546);
or U3036 (N_3036,N_227,N_745);
or U3037 (N_3037,N_1100,N_546);
xor U3038 (N_3038,N_157,N_148);
nor U3039 (N_3039,N_885,N_101);
or U3040 (N_3040,N_627,N_791);
xor U3041 (N_3041,N_1217,N_1369);
xnor U3042 (N_3042,N_1550,N_401);
nand U3043 (N_3043,N_729,N_1075);
xnor U3044 (N_3044,N_983,N_1564);
nor U3045 (N_3045,N_1565,N_1651);
and U3046 (N_3046,N_1152,N_210);
nor U3047 (N_3047,N_488,N_518);
nor U3048 (N_3048,N_612,N_882);
or U3049 (N_3049,N_374,N_1124);
or U3050 (N_3050,N_1801,N_111);
or U3051 (N_3051,N_1304,N_1210);
nand U3052 (N_3052,N_563,N_1564);
and U3053 (N_3053,N_871,N_1418);
xnor U3054 (N_3054,N_420,N_10);
nor U3055 (N_3055,N_737,N_371);
or U3056 (N_3056,N_1028,N_1904);
and U3057 (N_3057,N_1178,N_256);
nor U3058 (N_3058,N_418,N_1956);
nand U3059 (N_3059,N_1533,N_776);
nand U3060 (N_3060,N_1041,N_970);
or U3061 (N_3061,N_1872,N_582);
xnor U3062 (N_3062,N_650,N_579);
or U3063 (N_3063,N_1474,N_363);
xnor U3064 (N_3064,N_834,N_474);
xor U3065 (N_3065,N_1565,N_1155);
nand U3066 (N_3066,N_1688,N_1505);
and U3067 (N_3067,N_1690,N_335);
or U3068 (N_3068,N_1311,N_1639);
xor U3069 (N_3069,N_600,N_1907);
and U3070 (N_3070,N_1890,N_1558);
nand U3071 (N_3071,N_1579,N_99);
nor U3072 (N_3072,N_1988,N_246);
or U3073 (N_3073,N_188,N_877);
nand U3074 (N_3074,N_38,N_285);
nor U3075 (N_3075,N_40,N_1369);
xnor U3076 (N_3076,N_1693,N_153);
nand U3077 (N_3077,N_250,N_1380);
xnor U3078 (N_3078,N_1290,N_1199);
nand U3079 (N_3079,N_320,N_1899);
nand U3080 (N_3080,N_1163,N_1890);
or U3081 (N_3081,N_33,N_715);
xnor U3082 (N_3082,N_373,N_563);
xnor U3083 (N_3083,N_727,N_1595);
and U3084 (N_3084,N_1458,N_478);
and U3085 (N_3085,N_864,N_652);
or U3086 (N_3086,N_580,N_387);
nor U3087 (N_3087,N_1711,N_1145);
nor U3088 (N_3088,N_1215,N_787);
nor U3089 (N_3089,N_1418,N_1770);
xor U3090 (N_3090,N_1661,N_1616);
or U3091 (N_3091,N_1796,N_891);
and U3092 (N_3092,N_15,N_908);
and U3093 (N_3093,N_302,N_103);
xor U3094 (N_3094,N_1105,N_842);
and U3095 (N_3095,N_426,N_541);
nand U3096 (N_3096,N_322,N_412);
nor U3097 (N_3097,N_664,N_1750);
nor U3098 (N_3098,N_1172,N_595);
and U3099 (N_3099,N_1843,N_321);
nor U3100 (N_3100,N_224,N_1214);
nor U3101 (N_3101,N_423,N_686);
and U3102 (N_3102,N_322,N_75);
xor U3103 (N_3103,N_1044,N_301);
nand U3104 (N_3104,N_232,N_947);
nor U3105 (N_3105,N_1927,N_720);
nand U3106 (N_3106,N_1742,N_1127);
or U3107 (N_3107,N_1418,N_1684);
xnor U3108 (N_3108,N_1795,N_1133);
and U3109 (N_3109,N_708,N_1086);
nand U3110 (N_3110,N_774,N_767);
nand U3111 (N_3111,N_217,N_539);
nor U3112 (N_3112,N_1304,N_791);
xor U3113 (N_3113,N_1762,N_1233);
xor U3114 (N_3114,N_562,N_1601);
xnor U3115 (N_3115,N_1818,N_963);
nand U3116 (N_3116,N_189,N_1812);
nand U3117 (N_3117,N_429,N_1797);
xnor U3118 (N_3118,N_392,N_132);
and U3119 (N_3119,N_729,N_584);
or U3120 (N_3120,N_1430,N_107);
xor U3121 (N_3121,N_1164,N_440);
xnor U3122 (N_3122,N_214,N_421);
nand U3123 (N_3123,N_1147,N_1190);
and U3124 (N_3124,N_1811,N_821);
nand U3125 (N_3125,N_1028,N_276);
nand U3126 (N_3126,N_1404,N_1894);
nand U3127 (N_3127,N_1018,N_1410);
and U3128 (N_3128,N_1473,N_183);
nor U3129 (N_3129,N_1769,N_112);
and U3130 (N_3130,N_927,N_435);
nor U3131 (N_3131,N_94,N_414);
xor U3132 (N_3132,N_1439,N_769);
nor U3133 (N_3133,N_905,N_762);
nand U3134 (N_3134,N_796,N_1454);
xnor U3135 (N_3135,N_553,N_282);
or U3136 (N_3136,N_1364,N_1347);
xor U3137 (N_3137,N_1605,N_160);
nand U3138 (N_3138,N_661,N_152);
nor U3139 (N_3139,N_370,N_587);
nand U3140 (N_3140,N_1438,N_1667);
nand U3141 (N_3141,N_1486,N_715);
or U3142 (N_3142,N_104,N_527);
nand U3143 (N_3143,N_248,N_1711);
and U3144 (N_3144,N_1770,N_398);
or U3145 (N_3145,N_994,N_1389);
nor U3146 (N_3146,N_1650,N_201);
or U3147 (N_3147,N_1139,N_65);
xnor U3148 (N_3148,N_365,N_1962);
xnor U3149 (N_3149,N_672,N_1586);
nand U3150 (N_3150,N_13,N_159);
nor U3151 (N_3151,N_513,N_249);
or U3152 (N_3152,N_418,N_940);
nand U3153 (N_3153,N_793,N_1562);
or U3154 (N_3154,N_1286,N_1509);
xor U3155 (N_3155,N_733,N_20);
or U3156 (N_3156,N_1195,N_1079);
and U3157 (N_3157,N_1930,N_342);
or U3158 (N_3158,N_572,N_958);
nand U3159 (N_3159,N_35,N_1878);
nand U3160 (N_3160,N_1001,N_1650);
xnor U3161 (N_3161,N_98,N_625);
nor U3162 (N_3162,N_1785,N_1106);
and U3163 (N_3163,N_572,N_1913);
or U3164 (N_3164,N_1776,N_199);
and U3165 (N_3165,N_1203,N_425);
nor U3166 (N_3166,N_1914,N_375);
nor U3167 (N_3167,N_1678,N_1206);
or U3168 (N_3168,N_595,N_1968);
nand U3169 (N_3169,N_1645,N_500);
nor U3170 (N_3170,N_25,N_1532);
nor U3171 (N_3171,N_195,N_1510);
and U3172 (N_3172,N_476,N_1881);
and U3173 (N_3173,N_1856,N_276);
nor U3174 (N_3174,N_331,N_1834);
and U3175 (N_3175,N_1627,N_839);
or U3176 (N_3176,N_1005,N_263);
and U3177 (N_3177,N_608,N_1009);
nand U3178 (N_3178,N_1942,N_1050);
and U3179 (N_3179,N_1835,N_1460);
and U3180 (N_3180,N_1425,N_628);
xnor U3181 (N_3181,N_1712,N_757);
xnor U3182 (N_3182,N_1456,N_76);
nor U3183 (N_3183,N_447,N_489);
and U3184 (N_3184,N_1548,N_1664);
and U3185 (N_3185,N_893,N_38);
or U3186 (N_3186,N_656,N_434);
nor U3187 (N_3187,N_943,N_360);
and U3188 (N_3188,N_1531,N_1189);
nand U3189 (N_3189,N_1487,N_1409);
or U3190 (N_3190,N_1583,N_254);
nand U3191 (N_3191,N_273,N_708);
and U3192 (N_3192,N_1273,N_15);
nand U3193 (N_3193,N_1220,N_1598);
xnor U3194 (N_3194,N_1461,N_942);
or U3195 (N_3195,N_1133,N_906);
xnor U3196 (N_3196,N_935,N_70);
and U3197 (N_3197,N_1738,N_1656);
or U3198 (N_3198,N_1183,N_633);
or U3199 (N_3199,N_632,N_1324);
nor U3200 (N_3200,N_306,N_1019);
and U3201 (N_3201,N_287,N_443);
and U3202 (N_3202,N_1709,N_1968);
or U3203 (N_3203,N_654,N_99);
and U3204 (N_3204,N_1674,N_338);
nand U3205 (N_3205,N_1988,N_653);
xnor U3206 (N_3206,N_283,N_1316);
nand U3207 (N_3207,N_1574,N_1482);
or U3208 (N_3208,N_1293,N_1611);
or U3209 (N_3209,N_757,N_1803);
nor U3210 (N_3210,N_1433,N_1171);
nor U3211 (N_3211,N_1811,N_640);
nand U3212 (N_3212,N_1683,N_1864);
nor U3213 (N_3213,N_1714,N_1280);
nor U3214 (N_3214,N_239,N_1444);
nand U3215 (N_3215,N_1437,N_125);
nand U3216 (N_3216,N_1479,N_1475);
and U3217 (N_3217,N_1520,N_17);
nand U3218 (N_3218,N_639,N_497);
or U3219 (N_3219,N_1169,N_2);
or U3220 (N_3220,N_1178,N_1195);
nand U3221 (N_3221,N_290,N_1797);
nand U3222 (N_3222,N_1447,N_742);
xnor U3223 (N_3223,N_1873,N_992);
nor U3224 (N_3224,N_1059,N_134);
nand U3225 (N_3225,N_227,N_4);
nor U3226 (N_3226,N_1709,N_698);
nand U3227 (N_3227,N_678,N_1569);
nand U3228 (N_3228,N_19,N_1910);
nor U3229 (N_3229,N_771,N_1737);
or U3230 (N_3230,N_853,N_14);
or U3231 (N_3231,N_1922,N_1790);
nand U3232 (N_3232,N_828,N_365);
or U3233 (N_3233,N_857,N_1806);
xor U3234 (N_3234,N_320,N_1089);
nand U3235 (N_3235,N_982,N_701);
nand U3236 (N_3236,N_315,N_60);
or U3237 (N_3237,N_542,N_341);
and U3238 (N_3238,N_1531,N_1279);
and U3239 (N_3239,N_260,N_1208);
nand U3240 (N_3240,N_277,N_303);
and U3241 (N_3241,N_204,N_1352);
nand U3242 (N_3242,N_96,N_371);
xor U3243 (N_3243,N_616,N_467);
and U3244 (N_3244,N_1923,N_642);
xnor U3245 (N_3245,N_1361,N_1096);
nand U3246 (N_3246,N_1666,N_1809);
nand U3247 (N_3247,N_1260,N_522);
xor U3248 (N_3248,N_1199,N_983);
xnor U3249 (N_3249,N_451,N_1022);
and U3250 (N_3250,N_382,N_1804);
nand U3251 (N_3251,N_147,N_823);
nand U3252 (N_3252,N_810,N_875);
xor U3253 (N_3253,N_1847,N_1886);
and U3254 (N_3254,N_1558,N_110);
xor U3255 (N_3255,N_964,N_27);
and U3256 (N_3256,N_1385,N_409);
nor U3257 (N_3257,N_1785,N_371);
or U3258 (N_3258,N_810,N_1169);
xor U3259 (N_3259,N_286,N_853);
or U3260 (N_3260,N_926,N_406);
nand U3261 (N_3261,N_409,N_77);
and U3262 (N_3262,N_1736,N_1762);
xor U3263 (N_3263,N_150,N_30);
and U3264 (N_3264,N_1408,N_294);
nor U3265 (N_3265,N_1287,N_1163);
and U3266 (N_3266,N_259,N_1440);
or U3267 (N_3267,N_453,N_1497);
nor U3268 (N_3268,N_767,N_57);
or U3269 (N_3269,N_44,N_517);
and U3270 (N_3270,N_536,N_1789);
and U3271 (N_3271,N_699,N_1795);
and U3272 (N_3272,N_1851,N_768);
xor U3273 (N_3273,N_1048,N_142);
or U3274 (N_3274,N_345,N_1423);
or U3275 (N_3275,N_461,N_223);
xor U3276 (N_3276,N_1772,N_1228);
xnor U3277 (N_3277,N_134,N_171);
nor U3278 (N_3278,N_1607,N_1875);
nor U3279 (N_3279,N_836,N_1920);
and U3280 (N_3280,N_1642,N_1927);
or U3281 (N_3281,N_1615,N_560);
nand U3282 (N_3282,N_1716,N_1679);
xnor U3283 (N_3283,N_1519,N_752);
or U3284 (N_3284,N_873,N_777);
nand U3285 (N_3285,N_1168,N_259);
nor U3286 (N_3286,N_829,N_39);
nor U3287 (N_3287,N_53,N_1090);
or U3288 (N_3288,N_1577,N_1182);
and U3289 (N_3289,N_1286,N_1538);
and U3290 (N_3290,N_192,N_1119);
xnor U3291 (N_3291,N_1350,N_243);
nor U3292 (N_3292,N_1520,N_601);
xnor U3293 (N_3293,N_673,N_1783);
or U3294 (N_3294,N_1465,N_681);
xor U3295 (N_3295,N_761,N_691);
xor U3296 (N_3296,N_573,N_1575);
nor U3297 (N_3297,N_1298,N_736);
xnor U3298 (N_3298,N_1764,N_1213);
xnor U3299 (N_3299,N_1251,N_1368);
or U3300 (N_3300,N_1906,N_1311);
nand U3301 (N_3301,N_641,N_1827);
and U3302 (N_3302,N_107,N_335);
xnor U3303 (N_3303,N_1828,N_774);
and U3304 (N_3304,N_1085,N_127);
nand U3305 (N_3305,N_1707,N_1211);
or U3306 (N_3306,N_1170,N_401);
or U3307 (N_3307,N_536,N_247);
xnor U3308 (N_3308,N_1201,N_454);
nand U3309 (N_3309,N_78,N_1817);
or U3310 (N_3310,N_1682,N_1869);
nand U3311 (N_3311,N_785,N_1349);
nor U3312 (N_3312,N_283,N_908);
and U3313 (N_3313,N_1082,N_1787);
and U3314 (N_3314,N_1602,N_1383);
nand U3315 (N_3315,N_292,N_1573);
nand U3316 (N_3316,N_1620,N_1690);
and U3317 (N_3317,N_511,N_215);
xor U3318 (N_3318,N_64,N_55);
xnor U3319 (N_3319,N_1382,N_1880);
nor U3320 (N_3320,N_1415,N_1951);
or U3321 (N_3321,N_1418,N_1239);
and U3322 (N_3322,N_448,N_255);
xnor U3323 (N_3323,N_1604,N_1687);
nand U3324 (N_3324,N_255,N_92);
or U3325 (N_3325,N_1121,N_1056);
or U3326 (N_3326,N_1155,N_168);
xor U3327 (N_3327,N_1067,N_715);
xnor U3328 (N_3328,N_590,N_1804);
and U3329 (N_3329,N_1630,N_182);
xor U3330 (N_3330,N_1856,N_1707);
or U3331 (N_3331,N_1872,N_145);
nand U3332 (N_3332,N_1406,N_203);
and U3333 (N_3333,N_1944,N_851);
xor U3334 (N_3334,N_1664,N_580);
and U3335 (N_3335,N_1126,N_199);
and U3336 (N_3336,N_269,N_739);
xor U3337 (N_3337,N_594,N_1731);
nor U3338 (N_3338,N_642,N_54);
and U3339 (N_3339,N_1624,N_1381);
or U3340 (N_3340,N_1974,N_468);
nor U3341 (N_3341,N_1913,N_354);
nand U3342 (N_3342,N_1671,N_1154);
nor U3343 (N_3343,N_427,N_1217);
and U3344 (N_3344,N_198,N_1478);
nand U3345 (N_3345,N_1554,N_739);
and U3346 (N_3346,N_1275,N_1025);
nand U3347 (N_3347,N_1500,N_1269);
xor U3348 (N_3348,N_1456,N_635);
nand U3349 (N_3349,N_44,N_1809);
nand U3350 (N_3350,N_358,N_225);
nand U3351 (N_3351,N_437,N_1826);
xor U3352 (N_3352,N_309,N_1098);
xnor U3353 (N_3353,N_144,N_29);
nand U3354 (N_3354,N_1273,N_144);
xnor U3355 (N_3355,N_1045,N_1924);
nand U3356 (N_3356,N_1818,N_29);
nor U3357 (N_3357,N_1318,N_1808);
or U3358 (N_3358,N_315,N_804);
nand U3359 (N_3359,N_1013,N_1148);
or U3360 (N_3360,N_53,N_1322);
xnor U3361 (N_3361,N_1851,N_1742);
nor U3362 (N_3362,N_1434,N_719);
nor U3363 (N_3363,N_865,N_683);
and U3364 (N_3364,N_793,N_749);
nand U3365 (N_3365,N_1340,N_1503);
nor U3366 (N_3366,N_769,N_1033);
and U3367 (N_3367,N_242,N_1927);
and U3368 (N_3368,N_404,N_1069);
and U3369 (N_3369,N_1407,N_1114);
and U3370 (N_3370,N_1004,N_604);
nand U3371 (N_3371,N_272,N_1506);
xor U3372 (N_3372,N_821,N_1957);
xnor U3373 (N_3373,N_1415,N_1595);
nand U3374 (N_3374,N_657,N_1076);
xnor U3375 (N_3375,N_1146,N_295);
nor U3376 (N_3376,N_552,N_1676);
and U3377 (N_3377,N_218,N_140);
nor U3378 (N_3378,N_1225,N_714);
xnor U3379 (N_3379,N_458,N_1706);
nand U3380 (N_3380,N_715,N_1383);
nor U3381 (N_3381,N_1143,N_1282);
xor U3382 (N_3382,N_1610,N_728);
xnor U3383 (N_3383,N_1613,N_1569);
and U3384 (N_3384,N_1801,N_213);
and U3385 (N_3385,N_1924,N_608);
xnor U3386 (N_3386,N_1001,N_456);
nand U3387 (N_3387,N_936,N_1986);
and U3388 (N_3388,N_1065,N_734);
or U3389 (N_3389,N_1371,N_1667);
or U3390 (N_3390,N_1688,N_1043);
nand U3391 (N_3391,N_307,N_1656);
nand U3392 (N_3392,N_292,N_1681);
or U3393 (N_3393,N_1673,N_850);
nor U3394 (N_3394,N_762,N_589);
or U3395 (N_3395,N_845,N_1449);
nor U3396 (N_3396,N_826,N_603);
xnor U3397 (N_3397,N_557,N_333);
nand U3398 (N_3398,N_1880,N_1364);
nor U3399 (N_3399,N_1230,N_464);
xor U3400 (N_3400,N_25,N_757);
xor U3401 (N_3401,N_1150,N_1950);
or U3402 (N_3402,N_1075,N_1438);
or U3403 (N_3403,N_756,N_1952);
xnor U3404 (N_3404,N_1395,N_1841);
nand U3405 (N_3405,N_880,N_735);
xor U3406 (N_3406,N_378,N_861);
and U3407 (N_3407,N_1578,N_1822);
and U3408 (N_3408,N_1083,N_1293);
nand U3409 (N_3409,N_1438,N_542);
xnor U3410 (N_3410,N_620,N_1878);
and U3411 (N_3411,N_696,N_1697);
xnor U3412 (N_3412,N_192,N_1048);
xnor U3413 (N_3413,N_1905,N_727);
xor U3414 (N_3414,N_535,N_499);
xnor U3415 (N_3415,N_1832,N_1242);
nand U3416 (N_3416,N_970,N_1812);
nor U3417 (N_3417,N_269,N_1769);
xor U3418 (N_3418,N_440,N_803);
nor U3419 (N_3419,N_1283,N_1205);
or U3420 (N_3420,N_1920,N_1241);
or U3421 (N_3421,N_1057,N_993);
xor U3422 (N_3422,N_933,N_637);
or U3423 (N_3423,N_1122,N_821);
xor U3424 (N_3424,N_1732,N_915);
xnor U3425 (N_3425,N_359,N_1176);
or U3426 (N_3426,N_338,N_1878);
nand U3427 (N_3427,N_586,N_72);
or U3428 (N_3428,N_1291,N_924);
or U3429 (N_3429,N_1603,N_200);
nand U3430 (N_3430,N_69,N_1928);
or U3431 (N_3431,N_774,N_1559);
nor U3432 (N_3432,N_994,N_1349);
xor U3433 (N_3433,N_718,N_410);
and U3434 (N_3434,N_1530,N_635);
or U3435 (N_3435,N_110,N_982);
and U3436 (N_3436,N_211,N_1577);
xor U3437 (N_3437,N_710,N_426);
nand U3438 (N_3438,N_34,N_457);
or U3439 (N_3439,N_869,N_26);
nor U3440 (N_3440,N_466,N_995);
xor U3441 (N_3441,N_1414,N_909);
nor U3442 (N_3442,N_794,N_1447);
xnor U3443 (N_3443,N_1171,N_1583);
or U3444 (N_3444,N_1677,N_860);
and U3445 (N_3445,N_241,N_363);
nor U3446 (N_3446,N_720,N_341);
or U3447 (N_3447,N_134,N_1590);
or U3448 (N_3448,N_1545,N_1568);
nor U3449 (N_3449,N_723,N_984);
nand U3450 (N_3450,N_1450,N_487);
or U3451 (N_3451,N_1273,N_230);
nor U3452 (N_3452,N_437,N_1369);
xor U3453 (N_3453,N_1335,N_1892);
xnor U3454 (N_3454,N_1743,N_230);
nand U3455 (N_3455,N_665,N_1945);
nand U3456 (N_3456,N_1665,N_425);
nor U3457 (N_3457,N_1450,N_1213);
nor U3458 (N_3458,N_6,N_1777);
nor U3459 (N_3459,N_1466,N_711);
and U3460 (N_3460,N_320,N_250);
nand U3461 (N_3461,N_496,N_1335);
xor U3462 (N_3462,N_1996,N_541);
xor U3463 (N_3463,N_777,N_519);
and U3464 (N_3464,N_87,N_100);
and U3465 (N_3465,N_694,N_208);
nor U3466 (N_3466,N_195,N_781);
nor U3467 (N_3467,N_812,N_734);
xor U3468 (N_3468,N_531,N_877);
nand U3469 (N_3469,N_1975,N_1239);
xor U3470 (N_3470,N_384,N_1075);
xor U3471 (N_3471,N_970,N_183);
or U3472 (N_3472,N_1484,N_1022);
and U3473 (N_3473,N_1426,N_496);
nor U3474 (N_3474,N_1495,N_472);
nand U3475 (N_3475,N_237,N_1475);
nand U3476 (N_3476,N_708,N_1963);
nand U3477 (N_3477,N_1903,N_231);
xnor U3478 (N_3478,N_831,N_17);
nor U3479 (N_3479,N_154,N_1574);
nand U3480 (N_3480,N_177,N_1040);
and U3481 (N_3481,N_395,N_77);
xor U3482 (N_3482,N_1527,N_1524);
nor U3483 (N_3483,N_1957,N_614);
or U3484 (N_3484,N_664,N_905);
xnor U3485 (N_3485,N_1005,N_478);
nand U3486 (N_3486,N_1369,N_995);
nand U3487 (N_3487,N_965,N_1318);
and U3488 (N_3488,N_1013,N_1727);
or U3489 (N_3489,N_1990,N_442);
and U3490 (N_3490,N_1184,N_22);
xnor U3491 (N_3491,N_846,N_1534);
xnor U3492 (N_3492,N_208,N_1856);
xor U3493 (N_3493,N_392,N_1276);
nand U3494 (N_3494,N_944,N_161);
nor U3495 (N_3495,N_574,N_569);
nor U3496 (N_3496,N_828,N_469);
nand U3497 (N_3497,N_108,N_908);
or U3498 (N_3498,N_1464,N_871);
nand U3499 (N_3499,N_1791,N_1380);
xor U3500 (N_3500,N_1065,N_1567);
nor U3501 (N_3501,N_1010,N_1454);
nand U3502 (N_3502,N_1993,N_11);
xnor U3503 (N_3503,N_1246,N_1486);
nand U3504 (N_3504,N_1406,N_1148);
nor U3505 (N_3505,N_406,N_523);
xnor U3506 (N_3506,N_1775,N_69);
nand U3507 (N_3507,N_1896,N_1674);
and U3508 (N_3508,N_461,N_147);
nor U3509 (N_3509,N_1307,N_338);
or U3510 (N_3510,N_1139,N_239);
xor U3511 (N_3511,N_309,N_1983);
xnor U3512 (N_3512,N_1936,N_407);
nor U3513 (N_3513,N_953,N_1963);
and U3514 (N_3514,N_450,N_1310);
xor U3515 (N_3515,N_1501,N_1266);
or U3516 (N_3516,N_480,N_372);
nand U3517 (N_3517,N_717,N_107);
xnor U3518 (N_3518,N_1689,N_1904);
nor U3519 (N_3519,N_731,N_614);
or U3520 (N_3520,N_468,N_1100);
or U3521 (N_3521,N_241,N_1255);
or U3522 (N_3522,N_503,N_940);
and U3523 (N_3523,N_1024,N_1894);
nor U3524 (N_3524,N_1465,N_417);
xnor U3525 (N_3525,N_1590,N_807);
nor U3526 (N_3526,N_605,N_1483);
xor U3527 (N_3527,N_482,N_1084);
or U3528 (N_3528,N_502,N_1047);
xor U3529 (N_3529,N_1398,N_1224);
or U3530 (N_3530,N_1798,N_220);
xnor U3531 (N_3531,N_124,N_1705);
nand U3532 (N_3532,N_1421,N_1094);
or U3533 (N_3533,N_1782,N_1023);
or U3534 (N_3534,N_951,N_924);
and U3535 (N_3535,N_1520,N_1960);
xnor U3536 (N_3536,N_204,N_1324);
or U3537 (N_3537,N_1387,N_1835);
nor U3538 (N_3538,N_1360,N_1348);
and U3539 (N_3539,N_510,N_1016);
or U3540 (N_3540,N_1534,N_237);
nand U3541 (N_3541,N_861,N_263);
or U3542 (N_3542,N_623,N_835);
nor U3543 (N_3543,N_663,N_1148);
and U3544 (N_3544,N_1841,N_1982);
nand U3545 (N_3545,N_1281,N_1196);
nand U3546 (N_3546,N_1964,N_176);
and U3547 (N_3547,N_1026,N_812);
nand U3548 (N_3548,N_167,N_781);
xor U3549 (N_3549,N_1402,N_1976);
or U3550 (N_3550,N_1241,N_1661);
or U3551 (N_3551,N_327,N_1093);
xnor U3552 (N_3552,N_1377,N_1661);
nand U3553 (N_3553,N_547,N_1018);
or U3554 (N_3554,N_1532,N_1319);
xnor U3555 (N_3555,N_1135,N_436);
or U3556 (N_3556,N_1630,N_570);
or U3557 (N_3557,N_1111,N_1661);
nand U3558 (N_3558,N_46,N_128);
nand U3559 (N_3559,N_1306,N_1159);
and U3560 (N_3560,N_1378,N_1653);
nor U3561 (N_3561,N_1132,N_1810);
xor U3562 (N_3562,N_74,N_1669);
xnor U3563 (N_3563,N_219,N_324);
or U3564 (N_3564,N_188,N_1409);
nand U3565 (N_3565,N_57,N_146);
or U3566 (N_3566,N_915,N_1226);
nand U3567 (N_3567,N_1093,N_774);
xor U3568 (N_3568,N_1863,N_611);
nor U3569 (N_3569,N_792,N_523);
and U3570 (N_3570,N_1662,N_1540);
xor U3571 (N_3571,N_528,N_1148);
and U3572 (N_3572,N_1882,N_92);
nand U3573 (N_3573,N_987,N_407);
and U3574 (N_3574,N_1017,N_628);
xnor U3575 (N_3575,N_1614,N_527);
xor U3576 (N_3576,N_1505,N_465);
or U3577 (N_3577,N_1723,N_768);
and U3578 (N_3578,N_16,N_233);
nand U3579 (N_3579,N_1547,N_490);
and U3580 (N_3580,N_509,N_1083);
xnor U3581 (N_3581,N_1701,N_767);
nor U3582 (N_3582,N_1165,N_621);
nor U3583 (N_3583,N_1472,N_649);
and U3584 (N_3584,N_1739,N_1193);
and U3585 (N_3585,N_486,N_1752);
nand U3586 (N_3586,N_170,N_335);
or U3587 (N_3587,N_1829,N_1664);
nor U3588 (N_3588,N_256,N_939);
nand U3589 (N_3589,N_1737,N_1931);
nand U3590 (N_3590,N_1376,N_428);
nand U3591 (N_3591,N_1239,N_1680);
xnor U3592 (N_3592,N_1783,N_1484);
or U3593 (N_3593,N_1415,N_1557);
nor U3594 (N_3594,N_31,N_1091);
and U3595 (N_3595,N_1574,N_22);
nand U3596 (N_3596,N_924,N_393);
xor U3597 (N_3597,N_842,N_1326);
nor U3598 (N_3598,N_1532,N_1839);
or U3599 (N_3599,N_1901,N_1749);
or U3600 (N_3600,N_550,N_408);
xnor U3601 (N_3601,N_1732,N_1391);
and U3602 (N_3602,N_1829,N_1810);
nand U3603 (N_3603,N_1359,N_328);
or U3604 (N_3604,N_1458,N_1465);
nor U3605 (N_3605,N_64,N_249);
nor U3606 (N_3606,N_312,N_1453);
nor U3607 (N_3607,N_993,N_626);
or U3608 (N_3608,N_256,N_527);
nand U3609 (N_3609,N_90,N_1189);
nand U3610 (N_3610,N_581,N_1508);
and U3611 (N_3611,N_1935,N_1125);
or U3612 (N_3612,N_535,N_1929);
xor U3613 (N_3613,N_67,N_582);
or U3614 (N_3614,N_1216,N_1871);
and U3615 (N_3615,N_1846,N_1694);
and U3616 (N_3616,N_253,N_1959);
or U3617 (N_3617,N_1207,N_1686);
or U3618 (N_3618,N_1609,N_951);
nand U3619 (N_3619,N_1098,N_1688);
and U3620 (N_3620,N_1842,N_1757);
nand U3621 (N_3621,N_1061,N_802);
nand U3622 (N_3622,N_1770,N_809);
xor U3623 (N_3623,N_1039,N_1190);
nor U3624 (N_3624,N_779,N_1599);
nand U3625 (N_3625,N_1345,N_1840);
nand U3626 (N_3626,N_657,N_982);
and U3627 (N_3627,N_1151,N_1243);
nand U3628 (N_3628,N_1324,N_981);
or U3629 (N_3629,N_1353,N_930);
xnor U3630 (N_3630,N_1231,N_1182);
xor U3631 (N_3631,N_958,N_42);
nand U3632 (N_3632,N_1093,N_1003);
or U3633 (N_3633,N_7,N_912);
and U3634 (N_3634,N_668,N_542);
nand U3635 (N_3635,N_1116,N_1553);
and U3636 (N_3636,N_1690,N_1636);
nor U3637 (N_3637,N_1512,N_931);
and U3638 (N_3638,N_1033,N_441);
xnor U3639 (N_3639,N_913,N_901);
or U3640 (N_3640,N_1063,N_1443);
xor U3641 (N_3641,N_1758,N_1470);
or U3642 (N_3642,N_1674,N_1233);
xor U3643 (N_3643,N_293,N_691);
xor U3644 (N_3644,N_1120,N_1585);
nor U3645 (N_3645,N_1379,N_1099);
nor U3646 (N_3646,N_1436,N_66);
xor U3647 (N_3647,N_1482,N_1039);
xnor U3648 (N_3648,N_0,N_770);
or U3649 (N_3649,N_1219,N_1411);
xor U3650 (N_3650,N_1794,N_991);
xor U3651 (N_3651,N_139,N_1602);
xor U3652 (N_3652,N_478,N_990);
nand U3653 (N_3653,N_1069,N_527);
nor U3654 (N_3654,N_1209,N_1630);
nand U3655 (N_3655,N_1975,N_658);
or U3656 (N_3656,N_1664,N_661);
nor U3657 (N_3657,N_945,N_1317);
or U3658 (N_3658,N_1424,N_835);
or U3659 (N_3659,N_1657,N_1156);
nand U3660 (N_3660,N_1487,N_1397);
xnor U3661 (N_3661,N_1111,N_438);
nand U3662 (N_3662,N_1961,N_1356);
or U3663 (N_3663,N_400,N_1726);
nor U3664 (N_3664,N_1937,N_1479);
and U3665 (N_3665,N_1780,N_496);
or U3666 (N_3666,N_376,N_1788);
nor U3667 (N_3667,N_410,N_1719);
or U3668 (N_3668,N_581,N_950);
and U3669 (N_3669,N_1755,N_392);
or U3670 (N_3670,N_255,N_1385);
or U3671 (N_3671,N_919,N_483);
xnor U3672 (N_3672,N_707,N_359);
nand U3673 (N_3673,N_1536,N_1362);
and U3674 (N_3674,N_912,N_408);
xnor U3675 (N_3675,N_1307,N_920);
or U3676 (N_3676,N_1902,N_301);
nor U3677 (N_3677,N_1281,N_787);
nor U3678 (N_3678,N_1654,N_403);
nor U3679 (N_3679,N_1675,N_1169);
nor U3680 (N_3680,N_1783,N_516);
nand U3681 (N_3681,N_22,N_809);
nand U3682 (N_3682,N_235,N_524);
and U3683 (N_3683,N_652,N_456);
nor U3684 (N_3684,N_1654,N_1862);
or U3685 (N_3685,N_872,N_281);
or U3686 (N_3686,N_1770,N_425);
or U3687 (N_3687,N_1282,N_1844);
and U3688 (N_3688,N_1949,N_599);
nand U3689 (N_3689,N_32,N_1934);
and U3690 (N_3690,N_1469,N_1154);
nor U3691 (N_3691,N_1680,N_179);
xnor U3692 (N_3692,N_345,N_829);
or U3693 (N_3693,N_402,N_1961);
nand U3694 (N_3694,N_1847,N_300);
or U3695 (N_3695,N_475,N_1689);
xnor U3696 (N_3696,N_446,N_1865);
or U3697 (N_3697,N_362,N_1330);
or U3698 (N_3698,N_246,N_415);
or U3699 (N_3699,N_1063,N_669);
or U3700 (N_3700,N_187,N_474);
nand U3701 (N_3701,N_587,N_28);
and U3702 (N_3702,N_1835,N_776);
nand U3703 (N_3703,N_1471,N_364);
nand U3704 (N_3704,N_504,N_1727);
xnor U3705 (N_3705,N_366,N_1280);
nand U3706 (N_3706,N_1429,N_159);
or U3707 (N_3707,N_1079,N_415);
nand U3708 (N_3708,N_365,N_1092);
and U3709 (N_3709,N_428,N_259);
nand U3710 (N_3710,N_1552,N_1589);
or U3711 (N_3711,N_870,N_89);
nor U3712 (N_3712,N_1387,N_885);
or U3713 (N_3713,N_1270,N_1436);
xor U3714 (N_3714,N_745,N_302);
or U3715 (N_3715,N_1151,N_288);
nor U3716 (N_3716,N_1286,N_1578);
nor U3717 (N_3717,N_840,N_841);
nand U3718 (N_3718,N_149,N_1172);
and U3719 (N_3719,N_1201,N_1080);
or U3720 (N_3720,N_1698,N_248);
and U3721 (N_3721,N_1817,N_1149);
and U3722 (N_3722,N_678,N_355);
or U3723 (N_3723,N_310,N_628);
xnor U3724 (N_3724,N_418,N_1287);
nand U3725 (N_3725,N_1297,N_96);
and U3726 (N_3726,N_397,N_509);
or U3727 (N_3727,N_831,N_1869);
and U3728 (N_3728,N_1063,N_535);
nor U3729 (N_3729,N_202,N_899);
nor U3730 (N_3730,N_690,N_739);
or U3731 (N_3731,N_748,N_961);
or U3732 (N_3732,N_1278,N_1069);
nand U3733 (N_3733,N_1183,N_149);
nand U3734 (N_3734,N_1696,N_436);
xnor U3735 (N_3735,N_848,N_222);
xnor U3736 (N_3736,N_713,N_469);
nand U3737 (N_3737,N_329,N_928);
xor U3738 (N_3738,N_1720,N_342);
nand U3739 (N_3739,N_1901,N_796);
xnor U3740 (N_3740,N_1455,N_798);
and U3741 (N_3741,N_624,N_1891);
nor U3742 (N_3742,N_1825,N_1911);
and U3743 (N_3743,N_1927,N_1166);
nand U3744 (N_3744,N_790,N_507);
or U3745 (N_3745,N_1296,N_1939);
nand U3746 (N_3746,N_1941,N_1304);
nor U3747 (N_3747,N_489,N_1437);
nor U3748 (N_3748,N_1327,N_1734);
nor U3749 (N_3749,N_1354,N_1282);
or U3750 (N_3750,N_1575,N_1326);
nor U3751 (N_3751,N_1154,N_1354);
nor U3752 (N_3752,N_1018,N_1967);
nand U3753 (N_3753,N_1900,N_1887);
xor U3754 (N_3754,N_151,N_1867);
nand U3755 (N_3755,N_549,N_243);
nand U3756 (N_3756,N_1551,N_1282);
nor U3757 (N_3757,N_48,N_909);
nor U3758 (N_3758,N_63,N_45);
nand U3759 (N_3759,N_1874,N_1711);
xor U3760 (N_3760,N_807,N_311);
xnor U3761 (N_3761,N_1267,N_1669);
nor U3762 (N_3762,N_842,N_955);
xor U3763 (N_3763,N_1310,N_350);
xor U3764 (N_3764,N_1438,N_433);
xor U3765 (N_3765,N_425,N_184);
and U3766 (N_3766,N_752,N_1221);
nand U3767 (N_3767,N_1639,N_275);
and U3768 (N_3768,N_286,N_1586);
or U3769 (N_3769,N_814,N_1258);
nand U3770 (N_3770,N_1133,N_921);
and U3771 (N_3771,N_1192,N_734);
or U3772 (N_3772,N_813,N_165);
nor U3773 (N_3773,N_1448,N_1888);
or U3774 (N_3774,N_850,N_302);
or U3775 (N_3775,N_1072,N_560);
nand U3776 (N_3776,N_1981,N_811);
nand U3777 (N_3777,N_1106,N_145);
or U3778 (N_3778,N_1796,N_527);
nor U3779 (N_3779,N_1145,N_1207);
xnor U3780 (N_3780,N_1417,N_728);
or U3781 (N_3781,N_1486,N_635);
xnor U3782 (N_3782,N_594,N_72);
and U3783 (N_3783,N_1059,N_1945);
nand U3784 (N_3784,N_493,N_915);
nand U3785 (N_3785,N_652,N_1708);
xor U3786 (N_3786,N_1392,N_1208);
nor U3787 (N_3787,N_586,N_1320);
nand U3788 (N_3788,N_435,N_191);
or U3789 (N_3789,N_1438,N_1321);
and U3790 (N_3790,N_43,N_1680);
or U3791 (N_3791,N_1063,N_36);
nor U3792 (N_3792,N_1700,N_134);
or U3793 (N_3793,N_712,N_225);
or U3794 (N_3794,N_1632,N_1442);
and U3795 (N_3795,N_1258,N_538);
xor U3796 (N_3796,N_1585,N_119);
nand U3797 (N_3797,N_1304,N_760);
xnor U3798 (N_3798,N_47,N_1731);
and U3799 (N_3799,N_1736,N_1112);
xnor U3800 (N_3800,N_1603,N_1795);
xor U3801 (N_3801,N_1760,N_1156);
xnor U3802 (N_3802,N_1303,N_699);
nand U3803 (N_3803,N_1383,N_708);
nand U3804 (N_3804,N_1911,N_13);
xor U3805 (N_3805,N_953,N_1765);
xor U3806 (N_3806,N_1720,N_1152);
or U3807 (N_3807,N_458,N_1177);
xor U3808 (N_3808,N_1748,N_1004);
nor U3809 (N_3809,N_356,N_506);
nor U3810 (N_3810,N_1298,N_405);
xor U3811 (N_3811,N_187,N_85);
and U3812 (N_3812,N_1117,N_814);
xor U3813 (N_3813,N_1589,N_1100);
nor U3814 (N_3814,N_1605,N_1123);
nor U3815 (N_3815,N_940,N_556);
or U3816 (N_3816,N_999,N_155);
nand U3817 (N_3817,N_1294,N_763);
and U3818 (N_3818,N_1460,N_1626);
or U3819 (N_3819,N_997,N_1089);
xnor U3820 (N_3820,N_374,N_1882);
nor U3821 (N_3821,N_1944,N_401);
nand U3822 (N_3822,N_164,N_1055);
and U3823 (N_3823,N_1710,N_955);
nor U3824 (N_3824,N_1442,N_1658);
nor U3825 (N_3825,N_239,N_467);
nor U3826 (N_3826,N_880,N_366);
and U3827 (N_3827,N_141,N_1408);
nand U3828 (N_3828,N_182,N_30);
nor U3829 (N_3829,N_1363,N_1471);
nand U3830 (N_3830,N_921,N_1644);
nand U3831 (N_3831,N_273,N_303);
and U3832 (N_3832,N_1804,N_881);
or U3833 (N_3833,N_382,N_1452);
xor U3834 (N_3834,N_460,N_1791);
nor U3835 (N_3835,N_993,N_988);
nand U3836 (N_3836,N_1943,N_1565);
or U3837 (N_3837,N_1609,N_35);
xnor U3838 (N_3838,N_1958,N_949);
nand U3839 (N_3839,N_524,N_1112);
and U3840 (N_3840,N_1849,N_231);
xor U3841 (N_3841,N_855,N_1126);
xor U3842 (N_3842,N_1791,N_1955);
nand U3843 (N_3843,N_1900,N_522);
and U3844 (N_3844,N_1832,N_982);
nor U3845 (N_3845,N_376,N_32);
xor U3846 (N_3846,N_1479,N_1184);
or U3847 (N_3847,N_460,N_706);
and U3848 (N_3848,N_1244,N_510);
and U3849 (N_3849,N_67,N_1821);
xor U3850 (N_3850,N_1047,N_947);
nand U3851 (N_3851,N_898,N_571);
or U3852 (N_3852,N_542,N_460);
and U3853 (N_3853,N_929,N_1052);
or U3854 (N_3854,N_1917,N_1296);
xor U3855 (N_3855,N_1959,N_1972);
nor U3856 (N_3856,N_23,N_478);
xor U3857 (N_3857,N_484,N_508);
nand U3858 (N_3858,N_1018,N_1424);
xor U3859 (N_3859,N_1563,N_708);
nor U3860 (N_3860,N_1973,N_464);
xnor U3861 (N_3861,N_1172,N_1512);
nor U3862 (N_3862,N_460,N_1131);
nor U3863 (N_3863,N_111,N_1731);
nand U3864 (N_3864,N_69,N_1641);
and U3865 (N_3865,N_157,N_722);
xnor U3866 (N_3866,N_560,N_779);
and U3867 (N_3867,N_401,N_1617);
nand U3868 (N_3868,N_1122,N_1248);
nor U3869 (N_3869,N_677,N_792);
or U3870 (N_3870,N_1616,N_1671);
or U3871 (N_3871,N_1619,N_1426);
nand U3872 (N_3872,N_1400,N_1795);
or U3873 (N_3873,N_1807,N_1328);
or U3874 (N_3874,N_529,N_442);
and U3875 (N_3875,N_126,N_110);
nor U3876 (N_3876,N_365,N_872);
and U3877 (N_3877,N_559,N_791);
nand U3878 (N_3878,N_1906,N_728);
xor U3879 (N_3879,N_1809,N_540);
nand U3880 (N_3880,N_998,N_1696);
nor U3881 (N_3881,N_766,N_47);
or U3882 (N_3882,N_1810,N_1002);
nor U3883 (N_3883,N_655,N_1924);
nor U3884 (N_3884,N_941,N_1474);
nor U3885 (N_3885,N_1147,N_542);
or U3886 (N_3886,N_1885,N_124);
nand U3887 (N_3887,N_307,N_1131);
or U3888 (N_3888,N_946,N_1845);
and U3889 (N_3889,N_349,N_642);
nand U3890 (N_3890,N_131,N_1362);
nand U3891 (N_3891,N_1249,N_125);
or U3892 (N_3892,N_179,N_705);
or U3893 (N_3893,N_400,N_208);
or U3894 (N_3894,N_24,N_1868);
xor U3895 (N_3895,N_1753,N_1596);
or U3896 (N_3896,N_506,N_1447);
xnor U3897 (N_3897,N_1034,N_1673);
nand U3898 (N_3898,N_1738,N_1252);
nor U3899 (N_3899,N_420,N_1017);
nand U3900 (N_3900,N_1211,N_1203);
and U3901 (N_3901,N_1671,N_1018);
and U3902 (N_3902,N_8,N_1531);
nor U3903 (N_3903,N_293,N_468);
or U3904 (N_3904,N_68,N_1560);
nor U3905 (N_3905,N_1889,N_1193);
or U3906 (N_3906,N_1428,N_615);
nor U3907 (N_3907,N_751,N_776);
or U3908 (N_3908,N_1667,N_726);
xnor U3909 (N_3909,N_551,N_1139);
and U3910 (N_3910,N_744,N_1819);
nand U3911 (N_3911,N_279,N_1989);
or U3912 (N_3912,N_52,N_178);
or U3913 (N_3913,N_575,N_718);
and U3914 (N_3914,N_486,N_637);
and U3915 (N_3915,N_421,N_320);
nand U3916 (N_3916,N_83,N_1668);
and U3917 (N_3917,N_295,N_1551);
nand U3918 (N_3918,N_1682,N_1872);
and U3919 (N_3919,N_1167,N_804);
and U3920 (N_3920,N_981,N_605);
and U3921 (N_3921,N_341,N_1809);
and U3922 (N_3922,N_1055,N_1927);
nor U3923 (N_3923,N_38,N_1277);
and U3924 (N_3924,N_1103,N_1134);
xnor U3925 (N_3925,N_1122,N_373);
xnor U3926 (N_3926,N_995,N_762);
or U3927 (N_3927,N_470,N_1544);
and U3928 (N_3928,N_938,N_401);
and U3929 (N_3929,N_814,N_1907);
nand U3930 (N_3930,N_335,N_1334);
nor U3931 (N_3931,N_1679,N_1759);
xnor U3932 (N_3932,N_801,N_1586);
xnor U3933 (N_3933,N_860,N_395);
and U3934 (N_3934,N_1803,N_127);
nor U3935 (N_3935,N_1630,N_761);
xnor U3936 (N_3936,N_1334,N_1915);
and U3937 (N_3937,N_1134,N_1717);
xor U3938 (N_3938,N_1430,N_1714);
and U3939 (N_3939,N_1503,N_1307);
or U3940 (N_3940,N_1070,N_1851);
nor U3941 (N_3941,N_1768,N_1498);
nor U3942 (N_3942,N_1085,N_999);
and U3943 (N_3943,N_762,N_1337);
or U3944 (N_3944,N_939,N_1535);
xnor U3945 (N_3945,N_258,N_1032);
or U3946 (N_3946,N_31,N_167);
and U3947 (N_3947,N_459,N_1745);
and U3948 (N_3948,N_1227,N_1276);
or U3949 (N_3949,N_395,N_529);
or U3950 (N_3950,N_1855,N_588);
nor U3951 (N_3951,N_530,N_1668);
or U3952 (N_3952,N_562,N_1914);
and U3953 (N_3953,N_133,N_1986);
and U3954 (N_3954,N_1123,N_1524);
and U3955 (N_3955,N_674,N_396);
xor U3956 (N_3956,N_639,N_1199);
nand U3957 (N_3957,N_623,N_536);
or U3958 (N_3958,N_689,N_1815);
xnor U3959 (N_3959,N_1305,N_386);
nor U3960 (N_3960,N_893,N_310);
nand U3961 (N_3961,N_655,N_1044);
nor U3962 (N_3962,N_261,N_1131);
nor U3963 (N_3963,N_1739,N_428);
and U3964 (N_3964,N_1809,N_261);
nor U3965 (N_3965,N_1641,N_1279);
and U3966 (N_3966,N_1069,N_218);
nor U3967 (N_3967,N_933,N_868);
nand U3968 (N_3968,N_1747,N_1997);
nor U3969 (N_3969,N_883,N_1724);
nor U3970 (N_3970,N_886,N_535);
or U3971 (N_3971,N_1651,N_1294);
nand U3972 (N_3972,N_1522,N_1177);
nor U3973 (N_3973,N_762,N_28);
nor U3974 (N_3974,N_282,N_849);
nand U3975 (N_3975,N_1246,N_1997);
and U3976 (N_3976,N_1467,N_1692);
nand U3977 (N_3977,N_1760,N_1717);
xor U3978 (N_3978,N_851,N_411);
xnor U3979 (N_3979,N_1325,N_317);
xor U3980 (N_3980,N_1421,N_443);
nor U3981 (N_3981,N_419,N_52);
nor U3982 (N_3982,N_11,N_563);
nand U3983 (N_3983,N_1674,N_950);
nand U3984 (N_3984,N_167,N_1604);
and U3985 (N_3985,N_598,N_1959);
nand U3986 (N_3986,N_90,N_43);
xor U3987 (N_3987,N_1541,N_330);
or U3988 (N_3988,N_1380,N_1434);
xnor U3989 (N_3989,N_837,N_367);
or U3990 (N_3990,N_584,N_1199);
nand U3991 (N_3991,N_323,N_895);
xnor U3992 (N_3992,N_1315,N_1115);
nor U3993 (N_3993,N_803,N_633);
and U3994 (N_3994,N_349,N_1419);
nand U3995 (N_3995,N_1479,N_1306);
xor U3996 (N_3996,N_1411,N_747);
nor U3997 (N_3997,N_917,N_200);
or U3998 (N_3998,N_990,N_1469);
nand U3999 (N_3999,N_281,N_1281);
nor U4000 (N_4000,N_2645,N_3667);
nor U4001 (N_4001,N_3799,N_2700);
nor U4002 (N_4002,N_3991,N_2381);
nor U4003 (N_4003,N_2967,N_2701);
xnor U4004 (N_4004,N_3232,N_2254);
or U4005 (N_4005,N_2333,N_2594);
xor U4006 (N_4006,N_2162,N_2743);
nor U4007 (N_4007,N_3699,N_2454);
or U4008 (N_4008,N_2780,N_2834);
and U4009 (N_4009,N_2646,N_2145);
or U4010 (N_4010,N_3952,N_3826);
and U4011 (N_4011,N_2220,N_3139);
xnor U4012 (N_4012,N_3819,N_2112);
nand U4013 (N_4013,N_3481,N_3357);
xnor U4014 (N_4014,N_2833,N_2925);
xnor U4015 (N_4015,N_2434,N_3329);
nor U4016 (N_4016,N_3244,N_3393);
xor U4017 (N_4017,N_3445,N_3697);
and U4018 (N_4018,N_3479,N_3448);
nand U4019 (N_4019,N_2300,N_2073);
xor U4020 (N_4020,N_3258,N_3932);
xnor U4021 (N_4021,N_2379,N_3969);
xnor U4022 (N_4022,N_2561,N_2553);
xnor U4023 (N_4023,N_2596,N_2067);
and U4024 (N_4024,N_2005,N_2909);
or U4025 (N_4025,N_3511,N_3057);
xnor U4026 (N_4026,N_2931,N_3531);
or U4027 (N_4027,N_2643,N_2852);
xor U4028 (N_4028,N_3722,N_2471);
xor U4029 (N_4029,N_3761,N_3980);
nand U4030 (N_4030,N_2603,N_2205);
and U4031 (N_4031,N_2029,N_3065);
nor U4032 (N_4032,N_3256,N_3718);
and U4033 (N_4033,N_3178,N_2241);
xor U4034 (N_4034,N_2649,N_3430);
nand U4035 (N_4035,N_3536,N_2711);
and U4036 (N_4036,N_2707,N_3894);
xor U4037 (N_4037,N_3672,N_3276);
nand U4038 (N_4038,N_3294,N_2729);
and U4039 (N_4039,N_3158,N_2268);
nand U4040 (N_4040,N_2501,N_2634);
or U4041 (N_4041,N_3858,N_2447);
nand U4042 (N_4042,N_2330,N_2353);
or U4043 (N_4043,N_2320,N_2579);
and U4044 (N_4044,N_3459,N_2503);
xnor U4045 (N_4045,N_3746,N_3117);
nand U4046 (N_4046,N_2991,N_3328);
or U4047 (N_4047,N_3537,N_2010);
and U4048 (N_4048,N_3229,N_2824);
nand U4049 (N_4049,N_3671,N_3130);
and U4050 (N_4050,N_3175,N_3983);
xor U4051 (N_4051,N_3449,N_2635);
and U4052 (N_4052,N_3654,N_3008);
xor U4053 (N_4053,N_2375,N_3823);
nand U4054 (N_4054,N_2989,N_3047);
xnor U4055 (N_4055,N_3024,N_2959);
and U4056 (N_4056,N_3308,N_2715);
or U4057 (N_4057,N_2104,N_3153);
nor U4058 (N_4058,N_2150,N_2849);
xnor U4059 (N_4059,N_2633,N_2821);
nand U4060 (N_4060,N_2861,N_3595);
nand U4061 (N_4061,N_2516,N_3027);
and U4062 (N_4062,N_2489,N_3567);
or U4063 (N_4063,N_2250,N_3368);
nor U4064 (N_4064,N_2819,N_2283);
and U4065 (N_4065,N_3663,N_3520);
nor U4066 (N_4066,N_2227,N_2615);
xor U4067 (N_4067,N_3715,N_2483);
or U4068 (N_4068,N_3797,N_3001);
or U4069 (N_4069,N_3416,N_3780);
or U4070 (N_4070,N_3023,N_3404);
nor U4071 (N_4071,N_3634,N_2910);
xor U4072 (N_4072,N_3400,N_3255);
or U4073 (N_4073,N_3882,N_3740);
and U4074 (N_4074,N_3896,N_3542);
nand U4075 (N_4075,N_3769,N_3230);
nor U4076 (N_4076,N_2765,N_3692);
or U4077 (N_4077,N_2063,N_3381);
nand U4078 (N_4078,N_3086,N_3556);
nor U4079 (N_4079,N_2710,N_2725);
nor U4080 (N_4080,N_3380,N_3638);
nand U4081 (N_4081,N_2203,N_3909);
or U4082 (N_4082,N_3182,N_2284);
or U4083 (N_4083,N_2784,N_3745);
nand U4084 (N_4084,N_3719,N_3109);
xnor U4085 (N_4085,N_2424,N_3788);
and U4086 (N_4086,N_2787,N_2460);
nor U4087 (N_4087,N_2607,N_3660);
and U4088 (N_4088,N_3656,N_2046);
nand U4089 (N_4089,N_3790,N_3759);
and U4090 (N_4090,N_3734,N_3599);
xor U4091 (N_4091,N_3925,N_3825);
xor U4092 (N_4092,N_3437,N_3195);
nand U4093 (N_4093,N_3538,N_2000);
xor U4094 (N_4094,N_3604,N_3583);
or U4095 (N_4095,N_2986,N_2674);
nor U4096 (N_4096,N_3814,N_2409);
nor U4097 (N_4097,N_3771,N_3889);
nor U4098 (N_4098,N_2966,N_2900);
nor U4099 (N_4099,N_2221,N_3598);
or U4100 (N_4100,N_3326,N_2623);
xnor U4101 (N_4101,N_2100,N_3493);
or U4102 (N_4102,N_3074,N_2085);
nor U4103 (N_4103,N_3455,N_3702);
xor U4104 (N_4104,N_2259,N_2070);
xor U4105 (N_4105,N_3938,N_2621);
nand U4106 (N_4106,N_2593,N_3786);
and U4107 (N_4107,N_2987,N_3395);
nor U4108 (N_4108,N_2204,N_3714);
xnor U4109 (N_4109,N_2812,N_2018);
nor U4110 (N_4110,N_2288,N_3777);
xnor U4111 (N_4111,N_2979,N_2228);
nor U4112 (N_4112,N_2128,N_3042);
or U4113 (N_4113,N_2363,N_3475);
or U4114 (N_4114,N_2942,N_2573);
nand U4115 (N_4115,N_3054,N_3421);
nand U4116 (N_4116,N_3557,N_3774);
nor U4117 (N_4117,N_3364,N_2281);
nand U4118 (N_4118,N_2325,N_2659);
nor U4119 (N_4119,N_2164,N_3915);
or U4120 (N_4120,N_3624,N_2583);
nand U4121 (N_4121,N_3580,N_2044);
xor U4122 (N_4122,N_2897,N_3392);
nand U4123 (N_4123,N_3265,N_3432);
nand U4124 (N_4124,N_2420,N_3558);
nor U4125 (N_4125,N_2166,N_2341);
xor U4126 (N_4126,N_2226,N_2377);
nor U4127 (N_4127,N_3820,N_2832);
xor U4128 (N_4128,N_3176,N_2914);
nor U4129 (N_4129,N_2947,N_2212);
and U4130 (N_4130,N_2977,N_3010);
nor U4131 (N_4131,N_3462,N_2671);
xnor U4132 (N_4132,N_2704,N_3576);
nor U4133 (N_4133,N_3103,N_2862);
and U4134 (N_4134,N_3783,N_2415);
nor U4135 (N_4135,N_2136,N_3365);
xor U4136 (N_4136,N_2937,N_3457);
nand U4137 (N_4137,N_2586,N_2566);
nor U4138 (N_4138,N_3622,N_2169);
or U4139 (N_4139,N_3197,N_3907);
xor U4140 (N_4140,N_3278,N_2560);
nand U4141 (N_4141,N_2273,N_2094);
xnor U4142 (N_4142,N_3837,N_2695);
nand U4143 (N_4143,N_3353,N_3967);
nand U4144 (N_4144,N_2290,N_2324);
nand U4145 (N_4145,N_3424,N_2093);
nand U4146 (N_4146,N_2992,N_2518);
nor U4147 (N_4147,N_3245,N_3960);
xor U4148 (N_4148,N_3315,N_3497);
nand U4149 (N_4149,N_2080,N_3282);
or U4150 (N_4150,N_2151,N_2668);
nand U4151 (N_4151,N_2481,N_2514);
xnor U4152 (N_4152,N_3490,N_2177);
nand U4153 (N_4153,N_2970,N_3989);
xor U4154 (N_4154,N_3612,N_3770);
nand U4155 (N_4155,N_2801,N_2956);
or U4156 (N_4156,N_2337,N_3155);
or U4157 (N_4157,N_2686,N_3435);
or U4158 (N_4158,N_3933,N_2153);
nor U4159 (N_4159,N_2016,N_3104);
or U4160 (N_4160,N_3984,N_3854);
nor U4161 (N_4161,N_3091,N_3049);
nand U4162 (N_4162,N_2060,N_3690);
and U4163 (N_4163,N_3687,N_3524);
xor U4164 (N_4164,N_2474,N_3439);
or U4165 (N_4165,N_2476,N_2306);
nand U4166 (N_4166,N_2026,N_2215);
xnor U4167 (N_4167,N_2339,N_3693);
and U4168 (N_4168,N_2011,N_2039);
nor U4169 (N_4169,N_2143,N_3154);
or U4170 (N_4170,N_2554,N_2904);
nand U4171 (N_4171,N_3214,N_3478);
and U4172 (N_4172,N_2722,N_3762);
xnor U4173 (N_4173,N_2279,N_3354);
or U4174 (N_4174,N_3275,N_3089);
nor U4175 (N_4175,N_2015,N_2885);
nor U4176 (N_4176,N_3037,N_2628);
or U4177 (N_4177,N_3012,N_2282);
xor U4178 (N_4178,N_3829,N_2859);
xnor U4179 (N_4179,N_2437,N_2380);
nand U4180 (N_4180,N_3890,N_2269);
xor U4181 (N_4181,N_3375,N_3044);
nand U4182 (N_4182,N_2993,N_2693);
nor U4183 (N_4183,N_3846,N_2318);
nor U4184 (N_4184,N_3532,N_3813);
and U4185 (N_4185,N_3366,N_3434);
or U4186 (N_4186,N_3760,N_2493);
xor U4187 (N_4187,N_2135,N_2432);
and U4188 (N_4188,N_2488,N_2611);
or U4189 (N_4189,N_3540,N_3591);
xor U4190 (N_4190,N_3148,N_2097);
nand U4191 (N_4191,N_3233,N_2443);
nor U4192 (N_4192,N_3222,N_2519);
nand U4193 (N_4193,N_2877,N_2935);
xor U4194 (N_4194,N_3900,N_2562);
nand U4195 (N_4195,N_2405,N_3391);
nand U4196 (N_4196,N_3720,N_2004);
nor U4197 (N_4197,N_3845,N_2321);
xnor U4198 (N_4198,N_3076,N_2647);
nor U4199 (N_4199,N_2235,N_3396);
nor U4200 (N_4200,N_2124,N_3795);
xor U4201 (N_4201,N_2840,N_3464);
or U4202 (N_4202,N_3152,N_3655);
nand U4203 (N_4203,N_2602,N_2685);
nand U4204 (N_4204,N_3029,N_3322);
or U4205 (N_4205,N_3733,N_3847);
nor U4206 (N_4206,N_2720,N_3934);
or U4207 (N_4207,N_2193,N_2160);
nand U4208 (N_4208,N_2972,N_3281);
nand U4209 (N_4209,N_2034,N_2497);
xor U4210 (N_4210,N_3115,N_2800);
nand U4211 (N_4211,N_2247,N_3561);
nor U4212 (N_4212,N_3665,N_2081);
and U4213 (N_4213,N_2670,N_2983);
nand U4214 (N_4214,N_2737,N_3107);
nand U4215 (N_4215,N_2619,N_3552);
or U4216 (N_4216,N_2795,N_2390);
or U4217 (N_4217,N_2076,N_3048);
nor U4218 (N_4218,N_2901,N_2469);
or U4219 (N_4219,N_3530,N_2002);
nor U4220 (N_4220,N_3071,N_3249);
and U4221 (N_4221,N_2182,N_2786);
or U4222 (N_4222,N_2612,N_3879);
and U4223 (N_4223,N_2077,N_3463);
xor U4224 (N_4224,N_3600,N_2302);
xnor U4225 (N_4225,N_3905,N_3588);
nand U4226 (N_4226,N_3266,N_3191);
or U4227 (N_4227,N_2293,N_2650);
nor U4228 (N_4228,N_2708,N_2724);
nor U4229 (N_4229,N_3677,N_3767);
nand U4230 (N_4230,N_3941,N_3114);
nor U4231 (N_4231,N_2697,N_3261);
nand U4232 (N_4232,N_3043,N_3507);
nand U4233 (N_4233,N_2622,N_2492);
or U4234 (N_4234,N_2759,N_2731);
and U4235 (N_4235,N_3691,N_3857);
and U4236 (N_4236,N_3203,N_3053);
nand U4237 (N_4237,N_3956,N_2564);
or U4238 (N_4238,N_3628,N_3147);
or U4239 (N_4239,N_3781,N_2025);
xnor U4240 (N_4240,N_2892,N_2311);
or U4241 (N_4241,N_2091,N_2129);
nor U4242 (N_4242,N_2842,N_3725);
nand U4243 (N_4243,N_3413,N_2468);
xor U4244 (N_4244,N_3412,N_3943);
nor U4245 (N_4245,N_3264,N_3516);
or U4246 (N_4246,N_2933,N_2570);
xor U4247 (N_4247,N_3701,N_3986);
or U4248 (N_4248,N_2197,N_3133);
and U4249 (N_4249,N_3000,N_3397);
nand U4250 (N_4250,N_2482,N_3407);
nor U4251 (N_4251,N_3851,N_3417);
and U4252 (N_4252,N_2826,N_3917);
xnor U4253 (N_4253,N_3216,N_2827);
and U4254 (N_4254,N_2803,N_3243);
nor U4255 (N_4255,N_2639,N_2187);
and U4256 (N_4256,N_2682,N_2652);
and U4257 (N_4257,N_2716,N_3458);
or U4258 (N_4258,N_3190,N_2225);
xnor U4259 (N_4259,N_3274,N_3939);
nand U4260 (N_4260,N_2523,N_2581);
xnor U4261 (N_4261,N_2758,N_3776);
nor U4262 (N_4262,N_2352,N_3246);
nand U4263 (N_4263,N_3526,N_2176);
nand U4264 (N_4264,N_3288,N_3022);
nand U4265 (N_4265,N_2134,N_3514);
xnor U4266 (N_4266,N_2388,N_3834);
nor U4267 (N_4267,N_3059,N_3374);
nand U4268 (N_4268,N_3486,N_3100);
xor U4269 (N_4269,N_2510,N_2723);
or U4270 (N_4270,N_2732,N_3260);
or U4271 (N_4271,N_3642,N_2793);
nor U4272 (N_4272,N_3169,N_3961);
nand U4273 (N_4273,N_2750,N_2369);
xor U4274 (N_4274,N_2274,N_3267);
or U4275 (N_4275,N_2057,N_2557);
and U4276 (N_4276,N_2174,N_2576);
and U4277 (N_4277,N_2342,N_2442);
nand U4278 (N_4278,N_3904,N_3860);
and U4279 (N_4279,N_3948,N_3683);
or U4280 (N_4280,N_2955,N_3898);
xor U4281 (N_4281,N_3648,N_3348);
nand U4282 (N_4282,N_3192,N_3477);
xor U4283 (N_4283,N_2648,N_2994);
nand U4284 (N_4284,N_3843,N_3411);
xor U4285 (N_4285,N_3747,N_3379);
or U4286 (N_4286,N_3911,N_2421);
or U4287 (N_4287,N_2837,N_3436);
nor U4288 (N_4288,N_2272,N_2604);
xor U4289 (N_4289,N_3505,N_2184);
nor U4290 (N_4290,N_3138,N_2064);
nor U4291 (N_4291,N_2475,N_3386);
nand U4292 (N_4292,N_2637,N_3803);
and U4293 (N_4293,N_3174,N_2393);
nand U4294 (N_4294,N_2078,N_3808);
nand U4295 (N_4295,N_3739,N_3473);
nand U4296 (N_4296,N_3046,N_2059);
and U4297 (N_4297,N_3165,N_2003);
nor U4298 (N_4298,N_2445,N_3888);
or U4299 (N_4299,N_2350,N_2431);
nand U4300 (N_4300,N_3804,N_3822);
nor U4301 (N_4301,N_2111,N_3394);
nand U4302 (N_4302,N_3098,N_3212);
nor U4303 (N_4303,N_3559,N_2617);
or U4304 (N_4304,N_3962,N_3480);
or U4305 (N_4305,N_2001,N_3811);
xnor U4306 (N_4306,N_2446,N_2738);
and U4307 (N_4307,N_3077,N_3339);
or U4308 (N_4308,N_3242,N_3519);
xnor U4309 (N_4309,N_2858,N_3713);
nand U4310 (N_4310,N_3345,N_2061);
and U4311 (N_4311,N_2636,N_2303);
nand U4312 (N_4312,N_2895,N_3832);
nor U4313 (N_4313,N_3112,N_3867);
and U4314 (N_4314,N_2110,N_2130);
nand U4315 (N_4315,N_3425,N_3539);
or U4316 (N_4316,N_2349,N_2245);
and U4317 (N_4317,N_2630,N_2728);
and U4318 (N_4318,N_2556,N_2923);
or U4319 (N_4319,N_3387,N_3072);
nor U4320 (N_4320,N_2291,N_2665);
nor U4321 (N_4321,N_3703,N_3420);
nor U4322 (N_4322,N_2537,N_2857);
xnor U4323 (N_4323,N_2549,N_2797);
and U4324 (N_4324,N_3730,N_2748);
and U4325 (N_4325,N_2903,N_3597);
nand U4326 (N_4326,N_3555,N_3515);
xor U4327 (N_4327,N_3840,N_3185);
and U4328 (N_4328,N_2730,N_3087);
nor U4329 (N_4329,N_3501,N_3453);
and U4330 (N_4330,N_2717,N_2186);
xor U4331 (N_4331,N_3874,N_3675);
or U4332 (N_4332,N_2740,N_3290);
xnor U4333 (N_4333,N_3296,N_3650);
or U4334 (N_4334,N_3633,N_3172);
nor U4335 (N_4335,N_2920,N_2199);
or U4336 (N_4336,N_2037,N_3025);
and U4337 (N_4337,N_2936,N_2513);
xnor U4338 (N_4338,N_2908,N_2521);
nor U4339 (N_4339,N_3467,N_3224);
and U4340 (N_4340,N_3768,N_3880);
nor U4341 (N_4341,N_2323,N_2006);
nand U4342 (N_4342,N_2629,N_2132);
or U4343 (N_4343,N_2568,N_2036);
nor U4344 (N_4344,N_2411,N_3378);
or U4345 (N_4345,N_3712,N_3189);
and U4346 (N_4346,N_2660,N_3443);
xor U4347 (N_4347,N_2367,N_2326);
nor U4348 (N_4348,N_2175,N_2455);
xor U4349 (N_4349,N_3651,N_3050);
xor U4350 (N_4350,N_2981,N_3784);
and U4351 (N_4351,N_3965,N_3953);
xnor U4352 (N_4352,N_2504,N_2423);
nor U4353 (N_4353,N_2249,N_3283);
and U4354 (N_4354,N_2820,N_3085);
or U4355 (N_4355,N_2875,N_3094);
nand U4356 (N_4356,N_3553,N_2047);
or U4357 (N_4357,N_2571,N_2370);
xnor U4358 (N_4358,N_2741,N_3277);
nor U4359 (N_4359,N_3181,N_2086);
or U4360 (N_4360,N_3995,N_2438);
nor U4361 (N_4361,N_2314,N_3766);
and U4362 (N_4362,N_2307,N_2232);
nor U4363 (N_4363,N_3060,N_2789);
or U4364 (N_4364,N_3160,N_3541);
xor U4365 (N_4365,N_3234,N_2280);
nand U4366 (N_4366,N_3985,N_3645);
xor U4367 (N_4367,N_3491,N_3221);
nand U4368 (N_4368,N_2509,N_3157);
or U4369 (N_4369,N_3901,N_2627);
xor U4370 (N_4370,N_3543,N_2757);
and U4371 (N_4371,N_3056,N_2116);
and U4372 (N_4372,N_2694,N_2845);
nand U4373 (N_4373,N_2335,N_2574);
or U4374 (N_4374,N_3756,N_3004);
and U4375 (N_4375,N_3749,N_2102);
nor U4376 (N_4376,N_2939,N_3757);
nor U4377 (N_4377,N_2736,N_2090);
or U4378 (N_4378,N_2371,N_2746);
nand U4379 (N_4379,N_2552,N_2276);
nand U4380 (N_4380,N_2092,N_2703);
xor U4381 (N_4381,N_3796,N_2462);
nor U4382 (N_4382,N_3862,N_3990);
or U4383 (N_4383,N_2865,N_3061);
nand U4384 (N_4384,N_2683,N_2592);
xnor U4385 (N_4385,N_2915,N_2148);
xor U4386 (N_4386,N_2531,N_2426);
nand U4387 (N_4387,N_3325,N_3019);
or U4388 (N_4388,N_2285,N_3856);
nand U4389 (N_4389,N_2275,N_3226);
xnor U4390 (N_4390,N_3306,N_3723);
and U4391 (N_4391,N_3502,N_2218);
or U4392 (N_4392,N_2191,N_2927);
xnor U4393 (N_4393,N_3528,N_3918);
xor U4394 (N_4394,N_3332,N_3721);
nor U4395 (N_4395,N_3358,N_3498);
xnor U4396 (N_4396,N_2263,N_2133);
or U4397 (N_4397,N_3177,N_3922);
nand U4398 (N_4398,N_2329,N_2662);
nor U4399 (N_4399,N_3218,N_2163);
or U4400 (N_4400,N_3119,N_2040);
xor U4401 (N_4401,N_2995,N_2042);
nor U4402 (N_4402,N_2172,N_2769);
nand U4403 (N_4403,N_2261,N_2219);
xor U4404 (N_4404,N_3639,N_2068);
xor U4405 (N_4405,N_2798,N_3564);
nor U4406 (N_4406,N_3209,N_3549);
nor U4407 (N_4407,N_2173,N_2103);
nor U4408 (N_4408,N_2304,N_3159);
and U4409 (N_4409,N_2465,N_3465);
and U4410 (N_4410,N_3893,N_3083);
nand U4411 (N_4411,N_3641,N_2540);
nor U4412 (N_4412,N_3460,N_3668);
xnor U4413 (N_4413,N_3423,N_2580);
or U4414 (N_4414,N_2222,N_3142);
nor U4415 (N_4415,N_2257,N_2825);
or U4416 (N_4416,N_2921,N_3876);
nor U4417 (N_4417,N_2344,N_2971);
nand U4418 (N_4418,N_3335,N_3289);
nand U4419 (N_4419,N_2340,N_3311);
and U4420 (N_4420,N_2599,N_3513);
nand U4421 (N_4421,N_3207,N_2767);
and U4422 (N_4422,N_2528,N_3626);
nand U4423 (N_4423,N_2412,N_3533);
or U4424 (N_4424,N_2286,N_3593);
nor U4425 (N_4425,N_3180,N_3919);
xor U4426 (N_4426,N_2954,N_2463);
nor U4427 (N_4427,N_3954,N_3198);
xnor U4428 (N_4428,N_3162,N_2916);
or U4429 (N_4429,N_2013,N_3084);
and U4430 (N_4430,N_3807,N_3673);
nor U4431 (N_4431,N_3081,N_3979);
xnor U4432 (N_4432,N_3352,N_3875);
nand U4433 (N_4433,N_3447,N_2045);
or U4434 (N_4434,N_2591,N_3949);
or U4435 (N_4435,N_2651,N_2490);
xor U4436 (N_4436,N_2696,N_3710);
nor U4437 (N_4437,N_3067,N_3219);
xnor U4438 (N_4438,N_2520,N_2846);
xnor U4439 (N_4439,N_2030,N_3864);
and U4440 (N_4440,N_3284,N_2533);
and U4441 (N_4441,N_3619,N_2934);
and U4442 (N_4442,N_2456,N_2957);
and U4443 (N_4443,N_3116,N_3615);
or U4444 (N_4444,N_3126,N_3334);
or U4445 (N_4445,N_3011,N_2689);
xor U4446 (N_4446,N_2439,N_2802);
or U4447 (N_4447,N_3318,N_3350);
xnor U4448 (N_4448,N_3134,N_3020);
and U4449 (N_4449,N_2058,N_2677);
nor U4450 (N_4450,N_2601,N_3092);
or U4451 (N_4451,N_3279,N_3331);
nor U4452 (N_4452,N_3868,N_2973);
nor U4453 (N_4453,N_2383,N_2403);
xor U4454 (N_4454,N_2382,N_2451);
nor U4455 (N_4455,N_3271,N_3963);
and U4456 (N_4456,N_2113,N_2416);
nand U4457 (N_4457,N_2688,N_3577);
and U4458 (N_4458,N_3850,N_2347);
nand U4459 (N_4459,N_3844,N_2548);
xnor U4460 (N_4460,N_2019,N_2692);
or U4461 (N_4461,N_3323,N_2791);
nor U4462 (N_4462,N_3079,N_2588);
nand U4463 (N_4463,N_2753,N_2751);
xor U4464 (N_4464,N_3035,N_3006);
nor U4465 (N_4465,N_3484,N_2879);
and U4466 (N_4466,N_2433,N_3695);
nand U4467 (N_4467,N_2267,N_3285);
xnor U4468 (N_4468,N_3727,N_3483);
nor U4469 (N_4469,N_3349,N_2387);
xor U4470 (N_4470,N_2498,N_2642);
and U4471 (N_4471,N_2726,N_2190);
nand U4472 (N_4472,N_2213,N_2413);
and U4473 (N_4473,N_2679,N_3565);
nand U4474 (N_4474,N_3802,N_2401);
and U4475 (N_4475,N_3927,N_3653);
nand U4476 (N_4476,N_3187,N_2999);
nand U4477 (N_4477,N_2107,N_2126);
and U4478 (N_4478,N_2684,N_3976);
and U4479 (N_4479,N_3886,N_2464);
nor U4480 (N_4480,N_3183,N_2392);
and U4481 (N_4481,N_3509,N_3402);
or U4482 (N_4482,N_3631,N_3186);
or U4483 (N_4483,N_2891,N_2183);
nand U4484 (N_4484,N_3122,N_2527);
nand U4485 (N_4485,N_2022,N_2526);
or U4486 (N_4486,N_3623,N_3211);
xor U4487 (N_4487,N_3547,N_2362);
xnor U4488 (N_4488,N_3399,N_2161);
or U4489 (N_4489,N_2336,N_2843);
or U4490 (N_4490,N_2988,N_3821);
and U4491 (N_4491,N_2292,N_2886);
xnor U4492 (N_4492,N_2681,N_3450);
or U4493 (N_4493,N_2049,N_3908);
nor U4494 (N_4494,N_2760,N_2963);
nand U4495 (N_4495,N_3033,N_3923);
xnor U4496 (N_4496,N_3499,N_3069);
xor U4497 (N_4497,N_3582,N_2929);
nand U4498 (N_4498,N_3996,N_2799);
nand U4499 (N_4499,N_3128,N_3196);
and U4500 (N_4500,N_3500,N_2376);
or U4501 (N_4501,N_2754,N_3164);
xnor U4502 (N_4502,N_2354,N_2990);
xnor U4503 (N_4503,N_2185,N_2917);
and U4504 (N_4504,N_2962,N_2237);
or U4505 (N_4505,N_3131,N_2410);
and U4506 (N_4506,N_2719,N_3841);
nand U4507 (N_4507,N_2373,N_3300);
nor U4508 (N_4508,N_3034,N_2459);
and U4509 (N_4509,N_2663,N_3878);
and U4510 (N_4510,N_2976,N_2021);
nor U4511 (N_4511,N_2338,N_2295);
and U4512 (N_4512,N_2808,N_3657);
or U4513 (N_4513,N_2881,N_2785);
nand U4514 (N_4514,N_3835,N_2312);
xnor U4515 (N_4515,N_2969,N_3959);
xor U4516 (N_4516,N_2809,N_3356);
nor U4517 (N_4517,N_3247,N_2156);
nand U4518 (N_4518,N_2069,N_2202);
xnor U4519 (N_4519,N_2613,N_3666);
xnor U4520 (N_4520,N_2804,N_3609);
or U4521 (N_4521,N_3215,N_3563);
or U4522 (N_4522,N_2776,N_2610);
xor U4523 (N_4523,N_3248,N_3545);
nand U4524 (N_4524,N_2847,N_3385);
nand U4525 (N_4525,N_2631,N_2137);
and U4526 (N_4526,N_2582,N_3573);
nor U4527 (N_4527,N_2632,N_3062);
and U4528 (N_4528,N_3063,N_3744);
nor U4529 (N_4529,N_2031,N_3596);
or U4530 (N_4530,N_3101,N_3798);
nand U4531 (N_4531,N_2230,N_2502);
xor U4532 (N_4532,N_3441,N_3575);
xnor U4533 (N_4533,N_2384,N_2867);
and U4534 (N_4534,N_3026,N_3906);
xnor U4535 (N_4535,N_3369,N_3676);
xnor U4536 (N_4536,N_2609,N_2361);
nor U4537 (N_4537,N_2234,N_2691);
xor U4538 (N_4538,N_3066,N_2744);
nand U4539 (N_4539,N_2978,N_2958);
nor U4540 (N_4540,N_2258,N_3738);
xor U4541 (N_4541,N_2066,N_2322);
nor U4542 (N_4542,N_2868,N_2529);
nor U4543 (N_4543,N_3240,N_2790);
xnor U4544 (N_4544,N_2606,N_3970);
xor U4545 (N_4545,N_2075,N_2794);
nor U4546 (N_4546,N_2838,N_2654);
nor U4547 (N_4547,N_2214,N_3603);
nand U4548 (N_4548,N_3470,N_2425);
nand U4549 (N_4549,N_2051,N_2968);
or U4550 (N_4550,N_2813,N_2287);
nand U4551 (N_4551,N_2119,N_3250);
and U4552 (N_4552,N_3428,N_3293);
nand U4553 (N_4553,N_3370,N_2007);
or U4554 (N_4554,N_3041,N_2656);
and U4555 (N_4555,N_3403,N_3578);
nand U4556 (N_4556,N_2735,N_3073);
nand U4557 (N_4557,N_2171,N_2207);
xor U4558 (N_4558,N_3866,N_3377);
nor U4559 (N_4559,N_3316,N_2297);
or U4560 (N_4560,N_2653,N_2179);
xor U4561 (N_4561,N_2466,N_3589);
or U4562 (N_4562,N_3678,N_3307);
or U4563 (N_4563,N_3170,N_3075);
and U4564 (N_4564,N_3741,N_3251);
nor U4565 (N_4565,N_2524,N_2839);
nor U4566 (N_4566,N_2014,N_2511);
nor U4567 (N_4567,N_2907,N_2157);
nand U4568 (N_4568,N_3382,N_3398);
and U4569 (N_4569,N_2755,N_2035);
nor U4570 (N_4570,N_3030,N_2814);
and U4571 (N_4571,N_2188,N_3200);
or U4572 (N_4572,N_3885,N_3193);
nor U4573 (N_4573,N_2417,N_2569);
nand U4574 (N_4574,N_3964,N_2747);
or U4575 (N_4575,N_2099,N_2487);
or U4576 (N_4576,N_2690,N_3482);
xnor U4577 (N_4577,N_2898,N_2271);
nor U4578 (N_4578,N_3587,N_3751);
and U4579 (N_4579,N_2008,N_2578);
nor U4580 (N_4580,N_3168,N_3451);
or U4581 (N_4581,N_3914,N_3474);
nor U4582 (N_4582,N_3106,N_2948);
nor U4583 (N_4583,N_3728,N_2216);
nand U4584 (N_4584,N_2149,N_2138);
nand U4585 (N_4585,N_2638,N_3973);
xor U4586 (N_4586,N_3646,N_2082);
xnor U4587 (N_4587,N_3302,N_3338);
xor U4588 (N_4588,N_3494,N_3836);
xnor U4589 (N_4589,N_2980,N_3997);
xor U4590 (N_4590,N_3627,N_3684);
or U4591 (N_4591,N_3239,N_3805);
and U4592 (N_4592,N_3305,N_2399);
nand U4593 (N_4593,N_3504,N_2543);
xnor U4594 (N_4594,N_3883,N_3682);
nand U4595 (N_4595,N_3942,N_3958);
xor U4596 (N_4596,N_2248,N_3088);
or U4597 (N_4597,N_3038,N_2294);
nand U4598 (N_4598,N_3123,N_3611);
and U4599 (N_4599,N_3184,N_2450);
nand U4600 (N_4600,N_3390,N_3794);
xor U4601 (N_4601,N_2200,N_2419);
or U4602 (N_4602,N_2332,N_2127);
nand U4603 (N_4603,N_3070,N_2480);
xnor U4604 (N_4604,N_2938,N_3472);
nor U4605 (N_4605,N_2351,N_2189);
and U4606 (N_4606,N_2742,N_2851);
and U4607 (N_4607,N_3144,N_2308);
and U4608 (N_4608,N_3696,N_2033);
or U4609 (N_4609,N_3689,N_3848);
nor U4610 (N_4610,N_3367,N_2871);
and U4611 (N_4611,N_2998,N_2356);
nor U4612 (N_4612,N_2830,N_2953);
nor U4613 (N_4613,N_2745,N_2211);
nand U4614 (N_4614,N_3535,N_2547);
xor U4615 (N_4615,N_2309,N_2856);
and U4616 (N_4616,N_3488,N_3291);
nor U4617 (N_4617,N_3951,N_3686);
nand U4618 (N_4618,N_2178,N_2811);
and U4619 (N_4619,N_3227,N_3895);
and U4620 (N_4620,N_2810,N_2360);
or U4621 (N_4621,N_2277,N_3977);
or U4622 (N_4622,N_3418,N_3314);
nand U4623 (N_4623,N_3801,N_2734);
nor U4624 (N_4624,N_3869,N_2777);
or U4625 (N_4625,N_2605,N_3236);
and U4626 (N_4626,N_3806,N_3724);
or U4627 (N_4627,N_3912,N_2147);
nor U4628 (N_4628,N_2435,N_2641);
nor U4629 (N_4629,N_2964,N_3376);
or U4630 (N_4630,N_2544,N_2714);
nor U4631 (N_4631,N_3972,N_3974);
xnor U4632 (N_4632,N_2614,N_2142);
or U4633 (N_4633,N_3936,N_3787);
xnor U4634 (N_4634,N_3461,N_3231);
and U4635 (N_4635,N_2507,N_2244);
or U4636 (N_4636,N_2457,N_3940);
xnor U4637 (N_4637,N_2864,N_3419);
and U4638 (N_4638,N_2974,N_2778);
nor U4639 (N_4639,N_3815,N_2866);
nor U4640 (N_4640,N_3527,N_3617);
nor U4641 (N_4641,N_2158,N_2315);
nand U4642 (N_4642,N_3337,N_3852);
nor U4643 (N_4643,N_3865,N_3828);
and U4644 (N_4644,N_2334,N_3487);
or U4645 (N_4645,N_3892,N_3110);
nor U4646 (N_4646,N_3099,N_2698);
nor U4647 (N_4647,N_2783,N_3625);
nor U4648 (N_4648,N_2805,N_2944);
or U4649 (N_4649,N_2888,N_3992);
xor U4650 (N_4650,N_3015,N_3944);
or U4651 (N_4651,N_2661,N_3726);
nand U4652 (N_4652,N_2448,N_2499);
nand U4653 (N_4653,N_3643,N_3151);
and U4654 (N_4654,N_3204,N_3273);
or U4655 (N_4655,N_2587,N_2899);
nand U4656 (N_4656,N_2253,N_3095);
nand U4657 (N_4657,N_3661,N_2296);
and U4658 (N_4658,N_3145,N_2535);
xnor U4659 (N_4659,N_3090,N_2427);
nand U4660 (N_4660,N_3254,N_3485);
nand U4661 (N_4661,N_3743,N_3649);
xnor U4662 (N_4662,N_3208,N_2154);
xor U4663 (N_4663,N_3202,N_2874);
xnor U4664 (N_4664,N_3816,N_2771);
and U4665 (N_4665,N_3299,N_2125);
xnor U4666 (N_4666,N_3872,N_3993);
and U4667 (N_4667,N_3206,N_3446);
or U4668 (N_4668,N_3253,N_2123);
or U4669 (N_4669,N_2616,N_3605);
nor U4670 (N_4670,N_3966,N_2887);
or U4671 (N_4671,N_2705,N_2027);
or U4672 (N_4672,N_2088,N_3824);
and U4673 (N_4673,N_3055,N_2538);
xnor U4674 (N_4674,N_3606,N_2079);
nor U4675 (N_4675,N_2251,N_2246);
xnor U4676 (N_4676,N_3235,N_2709);
or U4677 (N_4677,N_2131,N_2152);
nand U4678 (N_4678,N_2041,N_3709);
or U4679 (N_4679,N_3877,N_3688);
nor U4680 (N_4680,N_2372,N_2928);
xor U4681 (N_4681,N_3201,N_2620);
nor U4682 (N_4682,N_3590,N_3842);
or U4683 (N_4683,N_3891,N_3809);
xnor U4684 (N_4684,N_2669,N_3735);
and U4685 (N_4685,N_2506,N_2749);
nor U4686 (N_4686,N_3704,N_2422);
and U4687 (N_4687,N_2368,N_2374);
xnor U4688 (N_4688,N_2243,N_2911);
xnor U4689 (N_4689,N_2301,N_3444);
nor U4690 (N_4690,N_3571,N_3102);
or U4691 (N_4691,N_2146,N_2389);
or U4692 (N_4692,N_2770,N_3135);
xnor U4693 (N_4693,N_3700,N_3789);
xnor U4694 (N_4694,N_3228,N_2270);
and U4695 (N_4695,N_3031,N_2555);
or U4696 (N_4696,N_3982,N_3257);
and U4697 (N_4697,N_2666,N_3705);
and U4698 (N_4698,N_3708,N_2658);
or U4699 (N_4699,N_2472,N_2238);
nand U4700 (N_4700,N_3928,N_3694);
xnor U4701 (N_4701,N_3736,N_2345);
and U4702 (N_4702,N_3161,N_2702);
nand U4703 (N_4703,N_3621,N_2121);
and U4704 (N_4704,N_2074,N_3988);
or U4705 (N_4705,N_2477,N_3268);
nor U4706 (N_4706,N_3669,N_2071);
or U4707 (N_4707,N_2919,N_2500);
xor U4708 (N_4708,N_2316,N_3476);
nor U4709 (N_4709,N_3213,N_3471);
nor U4710 (N_4710,N_2534,N_3658);
nand U4711 (N_4711,N_3120,N_2667);
or U4712 (N_4712,N_3156,N_3861);
or U4713 (N_4713,N_3389,N_2675);
nor U4714 (N_4714,N_3456,N_2120);
xnor U4715 (N_4715,N_3252,N_3884);
or U4716 (N_4716,N_3644,N_2260);
and U4717 (N_4717,N_2853,N_2926);
nand U4718 (N_4718,N_3833,N_3414);
nand U4719 (N_4719,N_3620,N_2065);
and U4720 (N_4720,N_2328,N_3068);
nor U4721 (N_4721,N_3737,N_2563);
or U4722 (N_4722,N_2313,N_3263);
or U4723 (N_4723,N_2050,N_3853);
or U4724 (N_4724,N_3550,N_3097);
nor U4725 (N_4725,N_2461,N_2101);
and U4726 (N_4726,N_2860,N_3931);
or U4727 (N_4727,N_3968,N_3401);
or U4728 (N_4728,N_3913,N_2585);
nand U4729 (N_4729,N_3469,N_2236);
nand U4730 (N_4730,N_3330,N_2884);
nand U4731 (N_4731,N_3987,N_2883);
nor U4732 (N_4732,N_2718,N_2083);
xor U4733 (N_4733,N_3647,N_3405);
nor U4734 (N_4734,N_3716,N_2657);
xor U4735 (N_4735,N_2348,N_3838);
or U4736 (N_4736,N_3945,N_2017);
xor U4737 (N_4737,N_2848,N_2949);
or U4738 (N_4738,N_3994,N_3150);
or U4739 (N_4739,N_2209,N_3298);
nand U4740 (N_4740,N_3362,N_3408);
or U4741 (N_4741,N_3924,N_3032);
or U4742 (N_4742,N_3748,N_2517);
or U4743 (N_4743,N_2298,N_2943);
nand U4744 (N_4744,N_3662,N_2397);
nor U4745 (N_4745,N_2817,N_2038);
or U4746 (N_4746,N_3132,N_2052);
nand U4747 (N_4747,N_3140,N_2484);
nand U4748 (N_4748,N_3111,N_2155);
and U4749 (N_4749,N_3706,N_2299);
nor U4750 (N_4750,N_3921,N_3618);
nor U4751 (N_4751,N_3568,N_3674);
xnor U4752 (N_4752,N_2766,N_2470);
xnor U4753 (N_4753,N_2626,N_2781);
or U4754 (N_4754,N_3632,N_3754);
and U4755 (N_4755,N_2062,N_2358);
nand U4756 (N_4756,N_2310,N_2841);
or U4757 (N_4757,N_2289,N_2597);
or U4758 (N_4758,N_2844,N_3863);
nor U4759 (N_4759,N_2491,N_2775);
and U4760 (N_4760,N_2266,N_2873);
nor U4761 (N_4761,N_3506,N_3262);
or U4762 (N_4762,N_2530,N_3764);
nand U4763 (N_4763,N_2109,N_3608);
nor U4764 (N_4764,N_3978,N_2404);
xor U4765 (N_4765,N_3319,N_2414);
nor U4766 (N_4766,N_3149,N_2224);
or U4767 (N_4767,N_2429,N_2053);
or U4768 (N_4768,N_2672,N_3426);
or U4769 (N_4769,N_2806,N_2252);
nand U4770 (N_4770,N_2201,N_2539);
and U4771 (N_4771,N_3778,N_3971);
or U4772 (N_4772,N_3388,N_3579);
nor U4773 (N_4773,N_2863,N_3188);
or U4774 (N_4774,N_3881,N_3827);
nor U4775 (N_4775,N_3926,N_3521);
nor U4776 (N_4776,N_2572,N_3523);
or U4777 (N_4777,N_3217,N_3946);
nand U4778 (N_4778,N_3742,N_2598);
nor U4779 (N_4779,N_3064,N_3007);
and U4780 (N_4780,N_2239,N_3327);
or U4781 (N_4781,N_3292,N_3546);
xor U4782 (N_4782,N_3309,N_3569);
and U4783 (N_4783,N_3586,N_2396);
and U4784 (N_4784,N_2317,N_3017);
or U4785 (N_4785,N_3998,N_2331);
nand U4786 (N_4786,N_3040,N_3259);
xnor U4787 (N_4787,N_2752,N_3146);
or U4788 (N_4788,N_2032,N_3343);
or U4789 (N_4789,N_3929,N_3910);
or U4790 (N_4790,N_3194,N_3551);
xor U4791 (N_4791,N_3018,N_2975);
nor U4792 (N_4792,N_2756,N_2400);
or U4793 (N_4793,N_2950,N_3468);
and U4794 (N_4794,N_2941,N_3503);
and U4795 (N_4795,N_3937,N_2357);
and U4796 (N_4796,N_3270,N_3082);
and U4797 (N_4797,N_2541,N_2418);
or U4798 (N_4798,N_3340,N_2020);
or U4799 (N_4799,N_3297,N_2905);
xor U4800 (N_4800,N_3849,N_2009);
and U4801 (N_4801,N_3359,N_2678);
nand U4802 (N_4802,N_3361,N_3080);
or U4803 (N_4803,N_3680,N_3096);
or U4804 (N_4804,N_2997,N_3594);
or U4805 (N_4805,N_3897,N_2792);
nor U4806 (N_4806,N_2878,N_3765);
xor U4807 (N_4807,N_2346,N_2105);
xor U4808 (N_4808,N_3630,N_3637);
and U4809 (N_4809,N_3859,N_2391);
or U4810 (N_4810,N_2996,N_2192);
nor U4811 (N_4811,N_2782,N_3752);
or U4812 (N_4812,N_3755,N_3711);
nor U4813 (N_4813,N_2512,N_2676);
or U4814 (N_4814,N_3916,N_3935);
and U4815 (N_4815,N_3887,N_2343);
nor U4816 (N_4816,N_3137,N_3344);
and U4817 (N_4817,N_2625,N_2365);
nand U4818 (N_4818,N_3014,N_3607);
nand U4819 (N_4819,N_3679,N_2772);
and U4820 (N_4820,N_2893,N_2436);
and U4821 (N_4821,N_2640,N_2788);
and U4822 (N_4822,N_3489,N_2012);
or U4823 (N_4823,N_3286,N_3830);
and U4824 (N_4824,N_2823,N_3930);
nand U4825 (N_4825,N_2816,N_2831);
and U4826 (N_4826,N_2319,N_3899);
or U4827 (N_4827,N_2600,N_2486);
and U4828 (N_4828,N_3782,N_2359);
nor U4829 (N_4829,N_2774,N_2855);
or U4830 (N_4830,N_2870,N_2932);
xor U4831 (N_4831,N_2089,N_2408);
and U4832 (N_4832,N_2761,N_3981);
or U4833 (N_4833,N_3051,N_2496);
and U4834 (N_4834,N_2876,N_2985);
or U4835 (N_4835,N_2869,N_3518);
nor U4836 (N_4836,N_3127,N_3529);
or U4837 (N_4837,N_2118,N_3548);
xnor U4838 (N_4838,N_2024,N_2198);
xnor U4839 (N_4839,N_2880,N_3433);
xnor U4840 (N_4840,N_2960,N_3601);
nand U4841 (N_4841,N_2961,N_3287);
nor U4842 (N_4842,N_2495,N_3036);
nand U4843 (N_4843,N_3199,N_2815);
and U4844 (N_4844,N_3124,N_3384);
or U4845 (N_4845,N_3812,N_2195);
and U4846 (N_4846,N_2624,N_3422);
nand U4847 (N_4847,N_2590,N_2940);
xnor U4848 (N_4848,N_3078,N_3902);
or U4849 (N_4849,N_3121,N_3205);
nor U4850 (N_4850,N_2930,N_2924);
nor U4851 (N_4851,N_3572,N_2278);
nor U4852 (N_4852,N_2558,N_2180);
and U4853 (N_4853,N_2918,N_2231);
nor U4854 (N_4854,N_3280,N_2796);
or U4855 (N_4855,N_2256,N_3818);
and U4856 (N_4856,N_3452,N_2072);
and U4857 (N_4857,N_2906,N_2449);
nor U4858 (N_4858,N_3903,N_3791);
nor U4859 (N_4859,N_3652,N_2458);
or U4860 (N_4860,N_3295,N_3021);
or U4861 (N_4861,N_3005,N_3415);
nor U4862 (N_4862,N_3955,N_2167);
nand U4863 (N_4863,N_2762,N_3241);
nand U4864 (N_4864,N_2551,N_3410);
or U4865 (N_4865,N_3574,N_3336);
nand U4866 (N_4866,N_2428,N_2850);
and U4867 (N_4867,N_2386,N_3303);
or U4868 (N_4868,N_2479,N_3492);
or U4869 (N_4869,N_3975,N_2223);
nand U4870 (N_4870,N_2054,N_2056);
nor U4871 (N_4871,N_3592,N_3758);
nor U4872 (N_4872,N_2194,N_2763);
xnor U4873 (N_4873,N_3118,N_3143);
or U4874 (N_4874,N_2913,N_2902);
and U4875 (N_4875,N_2467,N_2706);
or U4876 (N_4876,N_2768,N_3312);
nor U4877 (N_4877,N_2713,N_2106);
nor U4878 (N_4878,N_2922,N_2168);
nor U4879 (N_4879,N_3664,N_3341);
xnor U4880 (N_4880,N_2567,N_2140);
nand U4881 (N_4881,N_3510,N_2210);
and U4882 (N_4882,N_2452,N_3028);
xor U4883 (N_4883,N_3999,N_2687);
and U4884 (N_4884,N_3125,N_2208);
or U4885 (N_4885,N_2896,N_3581);
nand U4886 (N_4886,N_3610,N_2055);
nand U4887 (N_4887,N_3685,N_2087);
xor U4888 (N_4888,N_2508,N_3870);
xnor U4889 (N_4889,N_3640,N_3304);
xnor U4890 (N_4890,N_2525,N_3173);
and U4891 (N_4891,N_3052,N_3223);
and U4892 (N_4892,N_3950,N_2096);
and U4893 (N_4893,N_2882,N_2023);
xnor U4894 (N_4894,N_3636,N_3347);
nor U4895 (N_4895,N_3800,N_2721);
nand U4896 (N_4896,N_2965,N_3324);
nor U4897 (N_4897,N_2233,N_3957);
or U4898 (N_4898,N_2494,N_2394);
or U4899 (N_4899,N_2402,N_2043);
or U4900 (N_4900,N_3427,N_2265);
or U4901 (N_4901,N_3817,N_2440);
nor U4902 (N_4902,N_2536,N_3108);
nand U4903 (N_4903,N_2262,N_2395);
nor U4904 (N_4904,N_3810,N_3105);
and U4905 (N_4905,N_2206,N_2872);
or U4906 (N_4906,N_3495,N_3002);
xnor U4907 (N_4907,N_3167,N_2542);
or U4908 (N_4908,N_2305,N_2951);
nor U4909 (N_4909,N_3670,N_3317);
or U4910 (N_4910,N_3225,N_3466);
xnor U4911 (N_4911,N_3346,N_3792);
nand U4912 (N_4912,N_2577,N_2444);
or U4913 (N_4913,N_3429,N_3855);
xnor U4914 (N_4914,N_2589,N_2739);
or U4915 (N_4915,N_2122,N_2385);
and U4916 (N_4916,N_2378,N_2727);
or U4917 (N_4917,N_3372,N_3141);
or U4918 (N_4918,N_2522,N_2828);
nand U4919 (N_4919,N_3301,N_3873);
or U4920 (N_4920,N_3360,N_3313);
and U4921 (N_4921,N_3729,N_3237);
nor U4922 (N_4922,N_3272,N_2515);
or U4923 (N_4923,N_3775,N_3383);
nand U4924 (N_4924,N_2505,N_3442);
nand U4925 (N_4925,N_2829,N_3750);
or U4926 (N_4926,N_2165,N_2196);
xor U4927 (N_4927,N_2952,N_3584);
xor U4928 (N_4928,N_2644,N_2712);
xor U4929 (N_4929,N_3554,N_2836);
nand U4930 (N_4930,N_2699,N_2159);
nand U4931 (N_4931,N_2028,N_3566);
xor U4932 (N_4932,N_2355,N_2894);
or U4933 (N_4933,N_2559,N_3163);
nor U4934 (N_4934,N_2889,N_2764);
nor U4935 (N_4935,N_3570,N_2835);
or U4936 (N_4936,N_2144,N_3210);
and U4937 (N_4937,N_3717,N_2946);
nand U4938 (N_4938,N_2912,N_2807);
nand U4939 (N_4939,N_2565,N_3009);
nor U4940 (N_4940,N_2478,N_3659);
nand U4941 (N_4941,N_3136,N_3171);
nor U4942 (N_4942,N_3351,N_2114);
nand U4943 (N_4943,N_2673,N_3831);
and U4944 (N_4944,N_2406,N_2655);
xor U4945 (N_4945,N_3562,N_2264);
and U4946 (N_4946,N_3113,N_3522);
and U4947 (N_4947,N_3731,N_2818);
and U4948 (N_4948,N_2545,N_3373);
nand U4949 (N_4949,N_2115,N_3525);
and U4950 (N_4950,N_2441,N_3544);
nand U4951 (N_4951,N_2217,N_2984);
or U4952 (N_4952,N_3013,N_2550);
xnor U4953 (N_4953,N_2473,N_2822);
and U4954 (N_4954,N_2084,N_3496);
or U4955 (N_4955,N_3363,N_2255);
nand U4956 (N_4956,N_2664,N_2546);
and U4957 (N_4957,N_2733,N_3269);
nand U4958 (N_4958,N_3406,N_3045);
or U4959 (N_4959,N_3779,N_3793);
or U4960 (N_4960,N_2584,N_3371);
nor U4961 (N_4961,N_2170,N_2773);
nor U4962 (N_4962,N_2229,N_3517);
nor U4963 (N_4963,N_2854,N_2117);
nand U4964 (N_4964,N_2453,N_3635);
xor U4965 (N_4965,N_2364,N_3616);
or U4966 (N_4966,N_3772,N_3166);
nand U4967 (N_4967,N_3454,N_2608);
nor U4968 (N_4968,N_3058,N_2595);
or U4969 (N_4969,N_3039,N_3785);
nand U4970 (N_4970,N_3763,N_2430);
xor U4971 (N_4971,N_2095,N_3681);
or U4972 (N_4972,N_3602,N_2398);
nor U4973 (N_4973,N_3508,N_2242);
xnor U4974 (N_4974,N_3698,N_3016);
xor U4975 (N_4975,N_3534,N_3320);
nand U4976 (N_4976,N_3947,N_3179);
or U4977 (N_4977,N_3355,N_3560);
xnor U4978 (N_4978,N_3220,N_3512);
nand U4979 (N_4979,N_3129,N_2532);
or U4980 (N_4980,N_3839,N_2485);
nor U4981 (N_4981,N_3732,N_2048);
nand U4982 (N_4982,N_3871,N_2680);
and U4983 (N_4983,N_2327,N_2779);
nor U4984 (N_4984,N_3773,N_3438);
and U4985 (N_4985,N_2141,N_3614);
xor U4986 (N_4986,N_3920,N_3613);
nor U4987 (N_4987,N_3431,N_2108);
or U4988 (N_4988,N_3440,N_3333);
and U4989 (N_4989,N_3753,N_3409);
nor U4990 (N_4990,N_2407,N_3707);
nor U4991 (N_4991,N_2366,N_3342);
nor U4992 (N_4992,N_2098,N_3585);
and U4993 (N_4993,N_2181,N_2890);
and U4994 (N_4994,N_3093,N_2982);
and U4995 (N_4995,N_3238,N_2618);
nand U4996 (N_4996,N_2945,N_3321);
nor U4997 (N_4997,N_2575,N_3310);
xor U4998 (N_4998,N_3003,N_2240);
xor U4999 (N_4999,N_2139,N_3629);
and U5000 (N_5000,N_2240,N_2855);
nand U5001 (N_5001,N_2967,N_3486);
and U5002 (N_5002,N_2047,N_2346);
nor U5003 (N_5003,N_2050,N_3026);
nand U5004 (N_5004,N_2162,N_2033);
or U5005 (N_5005,N_2456,N_3687);
and U5006 (N_5006,N_3562,N_2626);
nand U5007 (N_5007,N_3963,N_2737);
nor U5008 (N_5008,N_2740,N_2504);
or U5009 (N_5009,N_2010,N_3842);
and U5010 (N_5010,N_3710,N_2501);
xnor U5011 (N_5011,N_2939,N_2468);
nor U5012 (N_5012,N_3162,N_2132);
nor U5013 (N_5013,N_2668,N_3973);
nand U5014 (N_5014,N_3160,N_3396);
or U5015 (N_5015,N_3275,N_2284);
nand U5016 (N_5016,N_2140,N_3433);
xnor U5017 (N_5017,N_2413,N_3090);
nor U5018 (N_5018,N_2202,N_3792);
nor U5019 (N_5019,N_3816,N_3985);
nor U5020 (N_5020,N_3093,N_2664);
nor U5021 (N_5021,N_3276,N_2925);
nor U5022 (N_5022,N_3049,N_3389);
xor U5023 (N_5023,N_2308,N_3377);
and U5024 (N_5024,N_3514,N_2233);
and U5025 (N_5025,N_3232,N_3658);
or U5026 (N_5026,N_3500,N_3900);
or U5027 (N_5027,N_3902,N_3882);
and U5028 (N_5028,N_2093,N_2246);
nand U5029 (N_5029,N_3132,N_2323);
nor U5030 (N_5030,N_2200,N_2929);
and U5031 (N_5031,N_2093,N_3092);
xnor U5032 (N_5032,N_3482,N_2849);
or U5033 (N_5033,N_3641,N_2098);
xnor U5034 (N_5034,N_3624,N_2931);
nor U5035 (N_5035,N_2069,N_3966);
xnor U5036 (N_5036,N_3745,N_2949);
nand U5037 (N_5037,N_3726,N_2519);
and U5038 (N_5038,N_3241,N_2317);
xnor U5039 (N_5039,N_3431,N_3018);
and U5040 (N_5040,N_2706,N_3027);
nand U5041 (N_5041,N_3148,N_3231);
nand U5042 (N_5042,N_2892,N_2972);
or U5043 (N_5043,N_3416,N_2376);
xor U5044 (N_5044,N_3612,N_2588);
nor U5045 (N_5045,N_3011,N_3932);
or U5046 (N_5046,N_2049,N_2959);
nor U5047 (N_5047,N_3682,N_3088);
nor U5048 (N_5048,N_3861,N_3519);
nand U5049 (N_5049,N_3941,N_3164);
and U5050 (N_5050,N_3856,N_2695);
and U5051 (N_5051,N_3008,N_3897);
nand U5052 (N_5052,N_2314,N_3901);
nor U5053 (N_5053,N_3857,N_3827);
and U5054 (N_5054,N_2294,N_3858);
nand U5055 (N_5055,N_3887,N_2111);
xnor U5056 (N_5056,N_3140,N_3829);
xnor U5057 (N_5057,N_3107,N_3228);
xnor U5058 (N_5058,N_3818,N_2711);
nor U5059 (N_5059,N_3700,N_3527);
or U5060 (N_5060,N_2666,N_2949);
and U5061 (N_5061,N_2095,N_2499);
or U5062 (N_5062,N_3151,N_2121);
or U5063 (N_5063,N_2953,N_3348);
or U5064 (N_5064,N_2995,N_3076);
nand U5065 (N_5065,N_2138,N_2193);
nand U5066 (N_5066,N_2239,N_2118);
nor U5067 (N_5067,N_2692,N_3865);
nor U5068 (N_5068,N_2437,N_2759);
and U5069 (N_5069,N_2154,N_3932);
and U5070 (N_5070,N_3971,N_2091);
and U5071 (N_5071,N_2802,N_2323);
nor U5072 (N_5072,N_2922,N_2320);
or U5073 (N_5073,N_2812,N_3853);
and U5074 (N_5074,N_3529,N_3133);
xor U5075 (N_5075,N_3583,N_3261);
xor U5076 (N_5076,N_2642,N_3005);
nand U5077 (N_5077,N_3704,N_2478);
nor U5078 (N_5078,N_3279,N_3451);
nor U5079 (N_5079,N_2000,N_2750);
and U5080 (N_5080,N_2233,N_2353);
nor U5081 (N_5081,N_3245,N_2527);
or U5082 (N_5082,N_2945,N_3930);
nand U5083 (N_5083,N_3725,N_2925);
nand U5084 (N_5084,N_2128,N_3849);
nand U5085 (N_5085,N_3817,N_2628);
and U5086 (N_5086,N_2591,N_3574);
xnor U5087 (N_5087,N_3562,N_2648);
nand U5088 (N_5088,N_2652,N_2686);
xor U5089 (N_5089,N_3920,N_3771);
or U5090 (N_5090,N_3193,N_3701);
or U5091 (N_5091,N_3339,N_2159);
and U5092 (N_5092,N_2897,N_3429);
xnor U5093 (N_5093,N_3028,N_2223);
and U5094 (N_5094,N_2598,N_3762);
nand U5095 (N_5095,N_3691,N_3271);
nand U5096 (N_5096,N_3480,N_2967);
xnor U5097 (N_5097,N_3198,N_2908);
xor U5098 (N_5098,N_2238,N_2819);
nand U5099 (N_5099,N_3522,N_3889);
nand U5100 (N_5100,N_3468,N_3842);
or U5101 (N_5101,N_2876,N_2076);
or U5102 (N_5102,N_2909,N_2298);
nand U5103 (N_5103,N_2848,N_3960);
nand U5104 (N_5104,N_2521,N_2958);
nor U5105 (N_5105,N_2854,N_3631);
xor U5106 (N_5106,N_2076,N_2158);
nor U5107 (N_5107,N_2612,N_3545);
xnor U5108 (N_5108,N_2192,N_3786);
xor U5109 (N_5109,N_3026,N_3809);
xnor U5110 (N_5110,N_2681,N_3562);
xnor U5111 (N_5111,N_3208,N_2197);
xnor U5112 (N_5112,N_2891,N_3923);
nand U5113 (N_5113,N_3764,N_2540);
xnor U5114 (N_5114,N_3166,N_2689);
nand U5115 (N_5115,N_2158,N_2776);
nand U5116 (N_5116,N_3900,N_3951);
and U5117 (N_5117,N_2749,N_3949);
xor U5118 (N_5118,N_2158,N_3122);
nor U5119 (N_5119,N_3997,N_2114);
nand U5120 (N_5120,N_2033,N_2412);
nand U5121 (N_5121,N_2556,N_3687);
xnor U5122 (N_5122,N_2573,N_2536);
nor U5123 (N_5123,N_3230,N_3546);
xor U5124 (N_5124,N_3642,N_3684);
and U5125 (N_5125,N_3487,N_2775);
xnor U5126 (N_5126,N_3274,N_2130);
nor U5127 (N_5127,N_2242,N_3259);
nor U5128 (N_5128,N_2358,N_3587);
or U5129 (N_5129,N_2969,N_3927);
nor U5130 (N_5130,N_2823,N_3534);
nand U5131 (N_5131,N_3615,N_3528);
and U5132 (N_5132,N_3634,N_3495);
nand U5133 (N_5133,N_2804,N_3049);
or U5134 (N_5134,N_2208,N_2333);
nand U5135 (N_5135,N_2249,N_3955);
nor U5136 (N_5136,N_3315,N_3540);
or U5137 (N_5137,N_3936,N_2611);
nand U5138 (N_5138,N_2085,N_2215);
and U5139 (N_5139,N_2870,N_3771);
and U5140 (N_5140,N_2840,N_3559);
nor U5141 (N_5141,N_2919,N_3527);
or U5142 (N_5142,N_3480,N_2129);
xnor U5143 (N_5143,N_2482,N_2553);
nor U5144 (N_5144,N_2491,N_3807);
and U5145 (N_5145,N_2870,N_2336);
and U5146 (N_5146,N_3754,N_3365);
nor U5147 (N_5147,N_3696,N_3901);
and U5148 (N_5148,N_2990,N_3119);
xor U5149 (N_5149,N_3448,N_3134);
xor U5150 (N_5150,N_3446,N_3172);
or U5151 (N_5151,N_2965,N_2534);
or U5152 (N_5152,N_3957,N_3927);
or U5153 (N_5153,N_2091,N_2534);
or U5154 (N_5154,N_3686,N_2035);
or U5155 (N_5155,N_2688,N_2194);
nand U5156 (N_5156,N_2559,N_2161);
or U5157 (N_5157,N_2270,N_3336);
or U5158 (N_5158,N_2633,N_2036);
or U5159 (N_5159,N_2987,N_3195);
nor U5160 (N_5160,N_3363,N_3896);
xnor U5161 (N_5161,N_2854,N_2258);
nand U5162 (N_5162,N_2712,N_2719);
nor U5163 (N_5163,N_3361,N_3774);
and U5164 (N_5164,N_2634,N_3576);
xor U5165 (N_5165,N_2459,N_3346);
nand U5166 (N_5166,N_3380,N_3924);
nor U5167 (N_5167,N_3401,N_2123);
or U5168 (N_5168,N_3284,N_3164);
nor U5169 (N_5169,N_2070,N_2856);
xor U5170 (N_5170,N_2635,N_2375);
and U5171 (N_5171,N_2106,N_3532);
nor U5172 (N_5172,N_3981,N_2952);
nor U5173 (N_5173,N_3628,N_2728);
xnor U5174 (N_5174,N_2441,N_2927);
xnor U5175 (N_5175,N_2760,N_3887);
xor U5176 (N_5176,N_2741,N_2795);
xor U5177 (N_5177,N_2703,N_2931);
xnor U5178 (N_5178,N_3673,N_2259);
nor U5179 (N_5179,N_2919,N_3019);
xnor U5180 (N_5180,N_2718,N_3605);
or U5181 (N_5181,N_3212,N_3167);
and U5182 (N_5182,N_2087,N_3915);
or U5183 (N_5183,N_3735,N_3368);
or U5184 (N_5184,N_2445,N_3065);
and U5185 (N_5185,N_3263,N_3672);
xnor U5186 (N_5186,N_3826,N_2307);
nor U5187 (N_5187,N_3043,N_2328);
xnor U5188 (N_5188,N_3649,N_2669);
nand U5189 (N_5189,N_2997,N_2462);
or U5190 (N_5190,N_2126,N_2416);
and U5191 (N_5191,N_2253,N_2175);
and U5192 (N_5192,N_3255,N_3994);
and U5193 (N_5193,N_3091,N_3534);
and U5194 (N_5194,N_3574,N_3486);
or U5195 (N_5195,N_3030,N_3098);
nor U5196 (N_5196,N_2905,N_2538);
or U5197 (N_5197,N_3982,N_2553);
xor U5198 (N_5198,N_3795,N_2925);
xor U5199 (N_5199,N_3416,N_3758);
or U5200 (N_5200,N_2499,N_2653);
xnor U5201 (N_5201,N_3250,N_2858);
nor U5202 (N_5202,N_3238,N_3030);
and U5203 (N_5203,N_3930,N_2820);
nand U5204 (N_5204,N_2834,N_3934);
or U5205 (N_5205,N_2386,N_2326);
or U5206 (N_5206,N_3864,N_3468);
and U5207 (N_5207,N_3378,N_3440);
xnor U5208 (N_5208,N_2917,N_3521);
nor U5209 (N_5209,N_2829,N_3593);
and U5210 (N_5210,N_3351,N_3287);
nand U5211 (N_5211,N_3178,N_2415);
nand U5212 (N_5212,N_2026,N_2746);
and U5213 (N_5213,N_3251,N_2312);
or U5214 (N_5214,N_2730,N_2143);
and U5215 (N_5215,N_2552,N_2423);
and U5216 (N_5216,N_3454,N_3249);
nor U5217 (N_5217,N_3796,N_2446);
or U5218 (N_5218,N_3146,N_2780);
or U5219 (N_5219,N_3296,N_3232);
or U5220 (N_5220,N_2170,N_3318);
xor U5221 (N_5221,N_2607,N_3374);
xor U5222 (N_5222,N_2275,N_3953);
and U5223 (N_5223,N_3390,N_3387);
nor U5224 (N_5224,N_2124,N_3959);
or U5225 (N_5225,N_2123,N_3544);
or U5226 (N_5226,N_2227,N_2995);
xnor U5227 (N_5227,N_3911,N_3217);
nor U5228 (N_5228,N_2722,N_2466);
nor U5229 (N_5229,N_3088,N_3994);
and U5230 (N_5230,N_2745,N_3228);
nor U5231 (N_5231,N_2393,N_3510);
xor U5232 (N_5232,N_2920,N_3614);
nand U5233 (N_5233,N_2247,N_3601);
or U5234 (N_5234,N_2395,N_2472);
nand U5235 (N_5235,N_3463,N_2196);
xor U5236 (N_5236,N_3815,N_3136);
and U5237 (N_5237,N_2429,N_2531);
nor U5238 (N_5238,N_2599,N_2678);
nor U5239 (N_5239,N_2867,N_2294);
nand U5240 (N_5240,N_3346,N_3193);
nor U5241 (N_5241,N_2667,N_3209);
and U5242 (N_5242,N_2147,N_2366);
or U5243 (N_5243,N_3907,N_2354);
nor U5244 (N_5244,N_2872,N_3972);
or U5245 (N_5245,N_2220,N_2011);
nor U5246 (N_5246,N_2850,N_3686);
xor U5247 (N_5247,N_3508,N_3904);
or U5248 (N_5248,N_2306,N_3304);
nand U5249 (N_5249,N_3367,N_2437);
nor U5250 (N_5250,N_2696,N_2386);
and U5251 (N_5251,N_2676,N_2659);
and U5252 (N_5252,N_2938,N_3102);
nand U5253 (N_5253,N_3732,N_2190);
nand U5254 (N_5254,N_2201,N_3380);
nand U5255 (N_5255,N_3682,N_3546);
xor U5256 (N_5256,N_3036,N_3983);
nand U5257 (N_5257,N_2859,N_2606);
or U5258 (N_5258,N_2596,N_3049);
xor U5259 (N_5259,N_3538,N_3877);
and U5260 (N_5260,N_3661,N_3187);
nand U5261 (N_5261,N_3332,N_2104);
nand U5262 (N_5262,N_3315,N_3896);
xor U5263 (N_5263,N_2560,N_2501);
nor U5264 (N_5264,N_2539,N_2955);
nor U5265 (N_5265,N_3145,N_3551);
or U5266 (N_5266,N_2952,N_3526);
nand U5267 (N_5267,N_2624,N_2569);
nor U5268 (N_5268,N_2710,N_3186);
and U5269 (N_5269,N_3208,N_3399);
and U5270 (N_5270,N_3121,N_3954);
or U5271 (N_5271,N_2378,N_2163);
and U5272 (N_5272,N_2513,N_3126);
and U5273 (N_5273,N_2009,N_3577);
or U5274 (N_5274,N_2254,N_3406);
nor U5275 (N_5275,N_3212,N_2674);
or U5276 (N_5276,N_2127,N_2764);
or U5277 (N_5277,N_3841,N_2742);
xor U5278 (N_5278,N_3512,N_2521);
or U5279 (N_5279,N_2738,N_2109);
and U5280 (N_5280,N_2423,N_3485);
nor U5281 (N_5281,N_2755,N_3585);
nand U5282 (N_5282,N_3154,N_3300);
nor U5283 (N_5283,N_2360,N_3089);
nor U5284 (N_5284,N_2189,N_2389);
nand U5285 (N_5285,N_2627,N_2953);
nor U5286 (N_5286,N_3807,N_2535);
or U5287 (N_5287,N_2610,N_3429);
nand U5288 (N_5288,N_3043,N_3258);
and U5289 (N_5289,N_2668,N_3130);
or U5290 (N_5290,N_3038,N_3961);
nor U5291 (N_5291,N_2110,N_2600);
or U5292 (N_5292,N_3086,N_2271);
or U5293 (N_5293,N_3459,N_2067);
and U5294 (N_5294,N_3918,N_2822);
xor U5295 (N_5295,N_2742,N_3611);
nor U5296 (N_5296,N_2659,N_3940);
xor U5297 (N_5297,N_3621,N_3511);
nand U5298 (N_5298,N_3292,N_3320);
xnor U5299 (N_5299,N_2998,N_2967);
nor U5300 (N_5300,N_2842,N_2986);
or U5301 (N_5301,N_3360,N_3441);
and U5302 (N_5302,N_3106,N_2472);
and U5303 (N_5303,N_3677,N_3488);
and U5304 (N_5304,N_2718,N_2490);
xnor U5305 (N_5305,N_3684,N_2952);
nand U5306 (N_5306,N_3529,N_3497);
xor U5307 (N_5307,N_3025,N_2167);
and U5308 (N_5308,N_3179,N_2110);
nand U5309 (N_5309,N_2093,N_3809);
nor U5310 (N_5310,N_2758,N_2742);
nand U5311 (N_5311,N_3819,N_2766);
or U5312 (N_5312,N_3603,N_2892);
and U5313 (N_5313,N_2735,N_2435);
nand U5314 (N_5314,N_2759,N_3071);
xor U5315 (N_5315,N_2192,N_3659);
or U5316 (N_5316,N_3360,N_3844);
nor U5317 (N_5317,N_2021,N_3047);
or U5318 (N_5318,N_3693,N_2702);
nand U5319 (N_5319,N_3054,N_2567);
xor U5320 (N_5320,N_3298,N_3549);
and U5321 (N_5321,N_2220,N_3453);
and U5322 (N_5322,N_3502,N_3014);
or U5323 (N_5323,N_2663,N_2485);
and U5324 (N_5324,N_2847,N_2047);
and U5325 (N_5325,N_3376,N_3270);
and U5326 (N_5326,N_2204,N_2380);
xor U5327 (N_5327,N_2199,N_2427);
nor U5328 (N_5328,N_3813,N_3140);
xnor U5329 (N_5329,N_3313,N_3781);
nand U5330 (N_5330,N_3602,N_2749);
or U5331 (N_5331,N_2642,N_2026);
nor U5332 (N_5332,N_2998,N_2124);
or U5333 (N_5333,N_3169,N_2107);
or U5334 (N_5334,N_3367,N_2835);
and U5335 (N_5335,N_2852,N_2224);
and U5336 (N_5336,N_2764,N_3250);
nand U5337 (N_5337,N_3221,N_2479);
xor U5338 (N_5338,N_3699,N_3642);
nand U5339 (N_5339,N_2144,N_2952);
and U5340 (N_5340,N_3281,N_3376);
and U5341 (N_5341,N_3254,N_3030);
nand U5342 (N_5342,N_2936,N_2710);
nor U5343 (N_5343,N_3236,N_2902);
nor U5344 (N_5344,N_3957,N_2613);
or U5345 (N_5345,N_3754,N_3459);
xnor U5346 (N_5346,N_3189,N_2077);
or U5347 (N_5347,N_2173,N_3816);
nand U5348 (N_5348,N_3893,N_2288);
nor U5349 (N_5349,N_2881,N_2988);
or U5350 (N_5350,N_3489,N_2593);
xnor U5351 (N_5351,N_2056,N_2093);
nor U5352 (N_5352,N_3157,N_3193);
and U5353 (N_5353,N_3521,N_3872);
and U5354 (N_5354,N_3985,N_3267);
nor U5355 (N_5355,N_3991,N_3781);
nand U5356 (N_5356,N_2849,N_2937);
and U5357 (N_5357,N_3561,N_2228);
or U5358 (N_5358,N_3642,N_3185);
nand U5359 (N_5359,N_2223,N_2836);
or U5360 (N_5360,N_3984,N_2181);
xnor U5361 (N_5361,N_2151,N_3387);
nor U5362 (N_5362,N_3813,N_3687);
nor U5363 (N_5363,N_3974,N_2401);
nand U5364 (N_5364,N_3151,N_2792);
and U5365 (N_5365,N_3303,N_3959);
and U5366 (N_5366,N_3303,N_2904);
nand U5367 (N_5367,N_2165,N_3756);
nand U5368 (N_5368,N_3722,N_3962);
nand U5369 (N_5369,N_3860,N_2680);
nand U5370 (N_5370,N_3503,N_3739);
nand U5371 (N_5371,N_3989,N_3763);
and U5372 (N_5372,N_2559,N_2943);
xor U5373 (N_5373,N_2601,N_2522);
nor U5374 (N_5374,N_3892,N_3837);
nand U5375 (N_5375,N_2974,N_3274);
nor U5376 (N_5376,N_2573,N_3994);
nor U5377 (N_5377,N_2383,N_3992);
xor U5378 (N_5378,N_2250,N_3344);
nand U5379 (N_5379,N_3953,N_3206);
nor U5380 (N_5380,N_3304,N_2584);
nor U5381 (N_5381,N_2554,N_3914);
and U5382 (N_5382,N_2599,N_2332);
and U5383 (N_5383,N_3239,N_2896);
or U5384 (N_5384,N_3012,N_3497);
nor U5385 (N_5385,N_2022,N_2622);
xor U5386 (N_5386,N_3577,N_2843);
xnor U5387 (N_5387,N_3864,N_3139);
and U5388 (N_5388,N_2984,N_2021);
nor U5389 (N_5389,N_2656,N_3896);
nand U5390 (N_5390,N_2073,N_2736);
nor U5391 (N_5391,N_2571,N_3777);
nand U5392 (N_5392,N_3526,N_3767);
nand U5393 (N_5393,N_3517,N_3189);
and U5394 (N_5394,N_3060,N_3154);
nor U5395 (N_5395,N_3312,N_2496);
nor U5396 (N_5396,N_2610,N_2265);
nor U5397 (N_5397,N_2887,N_2396);
nor U5398 (N_5398,N_2589,N_3477);
nand U5399 (N_5399,N_3595,N_3813);
and U5400 (N_5400,N_3002,N_2569);
and U5401 (N_5401,N_3869,N_2400);
and U5402 (N_5402,N_3294,N_2119);
xor U5403 (N_5403,N_3328,N_2231);
and U5404 (N_5404,N_3256,N_3413);
and U5405 (N_5405,N_2186,N_3620);
or U5406 (N_5406,N_3112,N_3422);
nor U5407 (N_5407,N_2398,N_2985);
xnor U5408 (N_5408,N_2979,N_2521);
and U5409 (N_5409,N_2402,N_2421);
xnor U5410 (N_5410,N_2042,N_2413);
or U5411 (N_5411,N_3776,N_2971);
and U5412 (N_5412,N_2851,N_3328);
nand U5413 (N_5413,N_2377,N_3961);
nor U5414 (N_5414,N_2378,N_3223);
and U5415 (N_5415,N_2487,N_2722);
xnor U5416 (N_5416,N_3445,N_2324);
or U5417 (N_5417,N_2575,N_2130);
nand U5418 (N_5418,N_2626,N_3122);
and U5419 (N_5419,N_3329,N_3458);
nor U5420 (N_5420,N_2148,N_3219);
xor U5421 (N_5421,N_2197,N_2812);
nand U5422 (N_5422,N_2729,N_2069);
and U5423 (N_5423,N_2744,N_2790);
nor U5424 (N_5424,N_3943,N_3683);
and U5425 (N_5425,N_2887,N_3226);
and U5426 (N_5426,N_2108,N_2671);
nand U5427 (N_5427,N_3567,N_2910);
or U5428 (N_5428,N_3365,N_2250);
nor U5429 (N_5429,N_3826,N_2141);
nor U5430 (N_5430,N_3994,N_2800);
xnor U5431 (N_5431,N_3977,N_2311);
nor U5432 (N_5432,N_3823,N_3612);
nor U5433 (N_5433,N_2491,N_3138);
and U5434 (N_5434,N_2825,N_2738);
xnor U5435 (N_5435,N_3332,N_2197);
xor U5436 (N_5436,N_3544,N_3117);
nor U5437 (N_5437,N_3157,N_2798);
or U5438 (N_5438,N_3962,N_2541);
nand U5439 (N_5439,N_2525,N_3567);
nor U5440 (N_5440,N_2495,N_3198);
nor U5441 (N_5441,N_2014,N_3323);
and U5442 (N_5442,N_2490,N_3692);
nor U5443 (N_5443,N_3295,N_3551);
and U5444 (N_5444,N_2291,N_2528);
or U5445 (N_5445,N_3513,N_3344);
nand U5446 (N_5446,N_3726,N_3309);
and U5447 (N_5447,N_3814,N_2368);
nor U5448 (N_5448,N_3074,N_3308);
xnor U5449 (N_5449,N_3784,N_2221);
nor U5450 (N_5450,N_2707,N_2574);
and U5451 (N_5451,N_3577,N_2361);
and U5452 (N_5452,N_2498,N_3875);
and U5453 (N_5453,N_2162,N_2736);
and U5454 (N_5454,N_2421,N_3867);
nand U5455 (N_5455,N_2593,N_3510);
xnor U5456 (N_5456,N_3965,N_2191);
and U5457 (N_5457,N_3526,N_3076);
nor U5458 (N_5458,N_3106,N_3245);
nor U5459 (N_5459,N_3009,N_2713);
xor U5460 (N_5460,N_2845,N_3226);
nand U5461 (N_5461,N_3998,N_3684);
or U5462 (N_5462,N_2248,N_3747);
nand U5463 (N_5463,N_3813,N_2690);
or U5464 (N_5464,N_2524,N_2301);
xor U5465 (N_5465,N_3288,N_2822);
or U5466 (N_5466,N_3430,N_3186);
and U5467 (N_5467,N_2345,N_3419);
nor U5468 (N_5468,N_3161,N_2645);
or U5469 (N_5469,N_3869,N_2271);
nor U5470 (N_5470,N_3290,N_2017);
nand U5471 (N_5471,N_2104,N_2510);
xnor U5472 (N_5472,N_2508,N_2449);
xor U5473 (N_5473,N_2896,N_2476);
xor U5474 (N_5474,N_2868,N_3365);
and U5475 (N_5475,N_2921,N_3333);
nand U5476 (N_5476,N_2820,N_3064);
xnor U5477 (N_5477,N_3035,N_3191);
and U5478 (N_5478,N_3266,N_3640);
nor U5479 (N_5479,N_2200,N_2646);
or U5480 (N_5480,N_2135,N_2946);
nand U5481 (N_5481,N_3465,N_2270);
or U5482 (N_5482,N_2665,N_3990);
or U5483 (N_5483,N_3690,N_3433);
or U5484 (N_5484,N_2383,N_3805);
or U5485 (N_5485,N_2129,N_3238);
nand U5486 (N_5486,N_2330,N_3549);
nor U5487 (N_5487,N_3138,N_3509);
and U5488 (N_5488,N_2528,N_2683);
and U5489 (N_5489,N_3159,N_3763);
and U5490 (N_5490,N_2110,N_2712);
or U5491 (N_5491,N_3298,N_3684);
or U5492 (N_5492,N_3642,N_3211);
nor U5493 (N_5493,N_3935,N_3876);
xor U5494 (N_5494,N_2854,N_3928);
nand U5495 (N_5495,N_2821,N_2327);
nor U5496 (N_5496,N_3324,N_3483);
nor U5497 (N_5497,N_3659,N_3853);
nand U5498 (N_5498,N_3792,N_3644);
nor U5499 (N_5499,N_3930,N_2843);
nor U5500 (N_5500,N_3389,N_2036);
nand U5501 (N_5501,N_2824,N_2066);
or U5502 (N_5502,N_2826,N_2110);
nand U5503 (N_5503,N_2331,N_3213);
xnor U5504 (N_5504,N_2907,N_3570);
nand U5505 (N_5505,N_3883,N_2125);
nor U5506 (N_5506,N_3348,N_3199);
xor U5507 (N_5507,N_3967,N_2670);
nand U5508 (N_5508,N_2427,N_2090);
and U5509 (N_5509,N_3065,N_3424);
nand U5510 (N_5510,N_2961,N_2307);
and U5511 (N_5511,N_3077,N_2825);
and U5512 (N_5512,N_2930,N_2961);
xnor U5513 (N_5513,N_2689,N_3852);
xnor U5514 (N_5514,N_2083,N_3558);
and U5515 (N_5515,N_2906,N_3244);
xnor U5516 (N_5516,N_3475,N_2460);
nor U5517 (N_5517,N_2200,N_3985);
xnor U5518 (N_5518,N_3657,N_2005);
and U5519 (N_5519,N_3462,N_2038);
nand U5520 (N_5520,N_2959,N_3903);
or U5521 (N_5521,N_2818,N_2298);
nand U5522 (N_5522,N_3362,N_2906);
nor U5523 (N_5523,N_3354,N_2169);
nand U5524 (N_5524,N_3588,N_3720);
nand U5525 (N_5525,N_3036,N_3078);
nand U5526 (N_5526,N_3663,N_3442);
nand U5527 (N_5527,N_3975,N_2109);
xor U5528 (N_5528,N_3967,N_2812);
xor U5529 (N_5529,N_3926,N_3262);
xnor U5530 (N_5530,N_2172,N_2804);
xnor U5531 (N_5531,N_2677,N_2119);
or U5532 (N_5532,N_3999,N_3136);
xor U5533 (N_5533,N_3984,N_2482);
nand U5534 (N_5534,N_3268,N_2177);
and U5535 (N_5535,N_2213,N_2772);
nand U5536 (N_5536,N_2495,N_2507);
and U5537 (N_5537,N_2211,N_3363);
nor U5538 (N_5538,N_3931,N_3881);
nand U5539 (N_5539,N_3499,N_2859);
nor U5540 (N_5540,N_2740,N_2584);
nand U5541 (N_5541,N_3239,N_3775);
nor U5542 (N_5542,N_3345,N_3826);
nand U5543 (N_5543,N_2355,N_3518);
and U5544 (N_5544,N_2040,N_2977);
and U5545 (N_5545,N_2202,N_2162);
nor U5546 (N_5546,N_3674,N_3039);
nand U5547 (N_5547,N_3313,N_3469);
nor U5548 (N_5548,N_3390,N_2925);
nor U5549 (N_5549,N_2970,N_2299);
nor U5550 (N_5550,N_2731,N_2204);
xnor U5551 (N_5551,N_2852,N_3773);
xor U5552 (N_5552,N_3470,N_3727);
or U5553 (N_5553,N_2709,N_3441);
and U5554 (N_5554,N_2015,N_2920);
or U5555 (N_5555,N_2009,N_2272);
nand U5556 (N_5556,N_2229,N_3845);
or U5557 (N_5557,N_3602,N_3347);
and U5558 (N_5558,N_3616,N_3066);
and U5559 (N_5559,N_2350,N_3960);
nor U5560 (N_5560,N_3181,N_2728);
nor U5561 (N_5561,N_2046,N_3029);
and U5562 (N_5562,N_2994,N_2256);
xnor U5563 (N_5563,N_3513,N_2950);
nor U5564 (N_5564,N_2931,N_3710);
or U5565 (N_5565,N_2787,N_2737);
or U5566 (N_5566,N_3822,N_2608);
nor U5567 (N_5567,N_3772,N_2752);
or U5568 (N_5568,N_3983,N_2068);
or U5569 (N_5569,N_3228,N_2305);
nor U5570 (N_5570,N_3549,N_2129);
nand U5571 (N_5571,N_3475,N_3707);
nand U5572 (N_5572,N_3933,N_3970);
or U5573 (N_5573,N_3195,N_2050);
xor U5574 (N_5574,N_3481,N_3807);
or U5575 (N_5575,N_2454,N_3387);
or U5576 (N_5576,N_2066,N_3554);
or U5577 (N_5577,N_3329,N_2830);
or U5578 (N_5578,N_2743,N_3670);
and U5579 (N_5579,N_3967,N_3236);
xnor U5580 (N_5580,N_3962,N_3785);
nand U5581 (N_5581,N_3948,N_3346);
nand U5582 (N_5582,N_2971,N_3868);
nand U5583 (N_5583,N_2045,N_2959);
nand U5584 (N_5584,N_2413,N_3416);
nand U5585 (N_5585,N_2381,N_3005);
nand U5586 (N_5586,N_3450,N_3608);
and U5587 (N_5587,N_3845,N_3126);
xnor U5588 (N_5588,N_2984,N_2389);
nor U5589 (N_5589,N_2940,N_2312);
xnor U5590 (N_5590,N_3085,N_2511);
xor U5591 (N_5591,N_3528,N_2293);
nor U5592 (N_5592,N_3933,N_2675);
or U5593 (N_5593,N_3525,N_2231);
xor U5594 (N_5594,N_3897,N_2151);
xnor U5595 (N_5595,N_3225,N_3940);
xnor U5596 (N_5596,N_3597,N_2596);
or U5597 (N_5597,N_2605,N_3631);
or U5598 (N_5598,N_2682,N_2904);
xnor U5599 (N_5599,N_2353,N_2060);
and U5600 (N_5600,N_3344,N_3201);
or U5601 (N_5601,N_3779,N_2979);
nand U5602 (N_5602,N_3337,N_2832);
or U5603 (N_5603,N_3842,N_3874);
xnor U5604 (N_5604,N_2171,N_2880);
and U5605 (N_5605,N_2380,N_2121);
nand U5606 (N_5606,N_3260,N_2194);
xnor U5607 (N_5607,N_2448,N_3973);
nor U5608 (N_5608,N_2369,N_3046);
or U5609 (N_5609,N_3618,N_2612);
and U5610 (N_5610,N_3223,N_2808);
nand U5611 (N_5611,N_3496,N_2464);
and U5612 (N_5612,N_3715,N_3197);
and U5613 (N_5613,N_3872,N_2375);
nand U5614 (N_5614,N_3810,N_2080);
or U5615 (N_5615,N_2675,N_2544);
nand U5616 (N_5616,N_2153,N_2234);
xor U5617 (N_5617,N_2579,N_3194);
and U5618 (N_5618,N_2584,N_3422);
and U5619 (N_5619,N_3091,N_3352);
or U5620 (N_5620,N_2787,N_2942);
xnor U5621 (N_5621,N_2805,N_3614);
nand U5622 (N_5622,N_2859,N_2783);
and U5623 (N_5623,N_3293,N_3244);
xor U5624 (N_5624,N_2992,N_2658);
nand U5625 (N_5625,N_2197,N_3236);
nor U5626 (N_5626,N_3818,N_2536);
and U5627 (N_5627,N_3151,N_2784);
nor U5628 (N_5628,N_2221,N_3171);
nor U5629 (N_5629,N_2005,N_2415);
xnor U5630 (N_5630,N_3240,N_3882);
nor U5631 (N_5631,N_3900,N_2403);
nor U5632 (N_5632,N_2548,N_3199);
nand U5633 (N_5633,N_3520,N_3310);
nor U5634 (N_5634,N_3400,N_3790);
or U5635 (N_5635,N_3613,N_3198);
nor U5636 (N_5636,N_3676,N_3417);
xnor U5637 (N_5637,N_2810,N_2553);
nand U5638 (N_5638,N_3401,N_2411);
nor U5639 (N_5639,N_2434,N_2510);
or U5640 (N_5640,N_2645,N_2914);
nand U5641 (N_5641,N_2721,N_3207);
or U5642 (N_5642,N_2754,N_3925);
nand U5643 (N_5643,N_2443,N_3912);
and U5644 (N_5644,N_3586,N_3380);
and U5645 (N_5645,N_2472,N_3687);
and U5646 (N_5646,N_3306,N_2542);
or U5647 (N_5647,N_3478,N_2639);
nor U5648 (N_5648,N_3947,N_3121);
or U5649 (N_5649,N_2727,N_2275);
xor U5650 (N_5650,N_2013,N_3750);
nand U5651 (N_5651,N_2002,N_2759);
and U5652 (N_5652,N_2327,N_3483);
and U5653 (N_5653,N_2591,N_3718);
and U5654 (N_5654,N_3075,N_2793);
xnor U5655 (N_5655,N_2406,N_3416);
or U5656 (N_5656,N_2824,N_2991);
xnor U5657 (N_5657,N_3346,N_2499);
or U5658 (N_5658,N_2897,N_3076);
or U5659 (N_5659,N_2494,N_2540);
or U5660 (N_5660,N_3190,N_2956);
nand U5661 (N_5661,N_2826,N_3805);
and U5662 (N_5662,N_2781,N_2040);
nor U5663 (N_5663,N_3126,N_3182);
nor U5664 (N_5664,N_3796,N_2212);
or U5665 (N_5665,N_2910,N_2256);
and U5666 (N_5666,N_2078,N_3470);
xnor U5667 (N_5667,N_2383,N_2459);
and U5668 (N_5668,N_2373,N_2209);
nand U5669 (N_5669,N_2997,N_3273);
and U5670 (N_5670,N_2305,N_2231);
xnor U5671 (N_5671,N_3877,N_3017);
nor U5672 (N_5672,N_2014,N_2621);
nor U5673 (N_5673,N_3918,N_2049);
and U5674 (N_5674,N_3693,N_2747);
and U5675 (N_5675,N_3660,N_3061);
or U5676 (N_5676,N_3765,N_3260);
nand U5677 (N_5677,N_3682,N_2027);
and U5678 (N_5678,N_3129,N_3496);
xnor U5679 (N_5679,N_3646,N_3267);
and U5680 (N_5680,N_3583,N_3384);
or U5681 (N_5681,N_3217,N_3052);
xnor U5682 (N_5682,N_3205,N_3582);
nor U5683 (N_5683,N_2241,N_3132);
xor U5684 (N_5684,N_3676,N_2055);
or U5685 (N_5685,N_2322,N_2957);
nor U5686 (N_5686,N_2171,N_2278);
or U5687 (N_5687,N_3342,N_2990);
nand U5688 (N_5688,N_2173,N_2993);
xnor U5689 (N_5689,N_3546,N_3235);
nand U5690 (N_5690,N_3874,N_2414);
and U5691 (N_5691,N_3936,N_3428);
nand U5692 (N_5692,N_2136,N_2790);
and U5693 (N_5693,N_2858,N_2044);
or U5694 (N_5694,N_3998,N_2103);
nor U5695 (N_5695,N_3942,N_2165);
nor U5696 (N_5696,N_2861,N_2050);
and U5697 (N_5697,N_3287,N_3378);
or U5698 (N_5698,N_2554,N_3521);
nand U5699 (N_5699,N_2027,N_2697);
nor U5700 (N_5700,N_3347,N_2041);
xor U5701 (N_5701,N_2858,N_2236);
nand U5702 (N_5702,N_2501,N_3702);
xnor U5703 (N_5703,N_2343,N_2876);
nor U5704 (N_5704,N_2918,N_3518);
or U5705 (N_5705,N_2938,N_2822);
and U5706 (N_5706,N_2366,N_2033);
or U5707 (N_5707,N_2195,N_3559);
nand U5708 (N_5708,N_3705,N_3779);
xor U5709 (N_5709,N_2227,N_3374);
nand U5710 (N_5710,N_3245,N_2011);
nor U5711 (N_5711,N_2329,N_2933);
and U5712 (N_5712,N_3032,N_3790);
and U5713 (N_5713,N_2249,N_2398);
xnor U5714 (N_5714,N_2011,N_2762);
or U5715 (N_5715,N_3963,N_2717);
and U5716 (N_5716,N_2837,N_3780);
and U5717 (N_5717,N_2660,N_3388);
nand U5718 (N_5718,N_2629,N_3771);
nand U5719 (N_5719,N_2359,N_3189);
nand U5720 (N_5720,N_2656,N_2563);
or U5721 (N_5721,N_3836,N_2499);
nor U5722 (N_5722,N_2982,N_3755);
nor U5723 (N_5723,N_2720,N_2557);
nand U5724 (N_5724,N_2907,N_2745);
nand U5725 (N_5725,N_2256,N_3931);
or U5726 (N_5726,N_3189,N_2209);
xnor U5727 (N_5727,N_2678,N_3830);
and U5728 (N_5728,N_3412,N_2120);
and U5729 (N_5729,N_2500,N_3447);
and U5730 (N_5730,N_2470,N_3956);
nor U5731 (N_5731,N_3820,N_2904);
xor U5732 (N_5732,N_3477,N_2496);
xnor U5733 (N_5733,N_3760,N_3308);
nand U5734 (N_5734,N_3825,N_2586);
and U5735 (N_5735,N_2774,N_2527);
and U5736 (N_5736,N_3644,N_2370);
nor U5737 (N_5737,N_3131,N_2397);
xor U5738 (N_5738,N_3244,N_3522);
and U5739 (N_5739,N_2750,N_3789);
or U5740 (N_5740,N_2731,N_3820);
or U5741 (N_5741,N_3007,N_2842);
nand U5742 (N_5742,N_3476,N_2212);
and U5743 (N_5743,N_3620,N_3761);
and U5744 (N_5744,N_3395,N_2343);
and U5745 (N_5745,N_3809,N_2761);
nor U5746 (N_5746,N_3187,N_3043);
nor U5747 (N_5747,N_3739,N_3959);
xnor U5748 (N_5748,N_2202,N_3938);
nor U5749 (N_5749,N_2033,N_2781);
or U5750 (N_5750,N_3476,N_2096);
xnor U5751 (N_5751,N_2184,N_3159);
nand U5752 (N_5752,N_2662,N_3844);
or U5753 (N_5753,N_3208,N_2406);
xnor U5754 (N_5754,N_3612,N_3920);
and U5755 (N_5755,N_2988,N_3045);
or U5756 (N_5756,N_3614,N_2219);
and U5757 (N_5757,N_2940,N_2755);
xor U5758 (N_5758,N_3069,N_2712);
xor U5759 (N_5759,N_3630,N_2699);
or U5760 (N_5760,N_3182,N_2037);
nor U5761 (N_5761,N_3731,N_3309);
or U5762 (N_5762,N_2395,N_2890);
or U5763 (N_5763,N_3365,N_2559);
and U5764 (N_5764,N_2427,N_2028);
nand U5765 (N_5765,N_2956,N_2957);
xor U5766 (N_5766,N_2161,N_3318);
nand U5767 (N_5767,N_3980,N_3875);
or U5768 (N_5768,N_2512,N_2008);
and U5769 (N_5769,N_3045,N_2545);
or U5770 (N_5770,N_2547,N_2271);
and U5771 (N_5771,N_3454,N_2028);
nor U5772 (N_5772,N_3747,N_2597);
nand U5773 (N_5773,N_3236,N_2778);
nand U5774 (N_5774,N_3671,N_3410);
or U5775 (N_5775,N_3094,N_2708);
nand U5776 (N_5776,N_3598,N_2466);
xnor U5777 (N_5777,N_3200,N_2720);
xnor U5778 (N_5778,N_2660,N_3207);
nor U5779 (N_5779,N_3392,N_3376);
nor U5780 (N_5780,N_3765,N_3936);
and U5781 (N_5781,N_3156,N_2864);
xor U5782 (N_5782,N_3745,N_2147);
nor U5783 (N_5783,N_3728,N_2509);
nand U5784 (N_5784,N_2172,N_3751);
nand U5785 (N_5785,N_2626,N_3262);
or U5786 (N_5786,N_2270,N_2759);
nor U5787 (N_5787,N_3990,N_2755);
xnor U5788 (N_5788,N_2886,N_3215);
xnor U5789 (N_5789,N_3569,N_2075);
nor U5790 (N_5790,N_2275,N_3343);
nand U5791 (N_5791,N_2563,N_3896);
and U5792 (N_5792,N_2961,N_2839);
nand U5793 (N_5793,N_2721,N_2193);
or U5794 (N_5794,N_2359,N_2902);
and U5795 (N_5795,N_3918,N_2613);
nor U5796 (N_5796,N_2380,N_3747);
or U5797 (N_5797,N_3927,N_2623);
nand U5798 (N_5798,N_3399,N_2704);
nor U5799 (N_5799,N_2291,N_3851);
or U5800 (N_5800,N_2091,N_3457);
and U5801 (N_5801,N_2879,N_3171);
and U5802 (N_5802,N_2910,N_2655);
or U5803 (N_5803,N_3696,N_2654);
and U5804 (N_5804,N_3824,N_3408);
nor U5805 (N_5805,N_2221,N_2159);
and U5806 (N_5806,N_2786,N_3805);
and U5807 (N_5807,N_2807,N_2419);
xnor U5808 (N_5808,N_2039,N_2613);
xor U5809 (N_5809,N_3318,N_2971);
xor U5810 (N_5810,N_3371,N_3339);
nor U5811 (N_5811,N_2548,N_2808);
xnor U5812 (N_5812,N_3286,N_3663);
and U5813 (N_5813,N_3124,N_3970);
nor U5814 (N_5814,N_2237,N_2652);
and U5815 (N_5815,N_2135,N_3533);
nor U5816 (N_5816,N_2778,N_2596);
nor U5817 (N_5817,N_2405,N_2050);
xor U5818 (N_5818,N_2286,N_2716);
or U5819 (N_5819,N_2246,N_2574);
and U5820 (N_5820,N_3022,N_3195);
nor U5821 (N_5821,N_3587,N_3290);
and U5822 (N_5822,N_2924,N_2083);
or U5823 (N_5823,N_2566,N_2850);
xor U5824 (N_5824,N_2652,N_3423);
nor U5825 (N_5825,N_3319,N_2243);
or U5826 (N_5826,N_3211,N_3867);
and U5827 (N_5827,N_3123,N_2787);
nor U5828 (N_5828,N_2997,N_2472);
xor U5829 (N_5829,N_2795,N_2833);
xnor U5830 (N_5830,N_3911,N_2174);
or U5831 (N_5831,N_3081,N_2047);
nand U5832 (N_5832,N_3359,N_3768);
and U5833 (N_5833,N_3060,N_3274);
nor U5834 (N_5834,N_3634,N_3577);
or U5835 (N_5835,N_2695,N_3936);
xnor U5836 (N_5836,N_3618,N_3526);
or U5837 (N_5837,N_2427,N_2983);
nand U5838 (N_5838,N_2901,N_2555);
and U5839 (N_5839,N_2980,N_3000);
and U5840 (N_5840,N_2525,N_2568);
or U5841 (N_5841,N_3562,N_2170);
nor U5842 (N_5842,N_3929,N_3510);
xor U5843 (N_5843,N_3974,N_2043);
xnor U5844 (N_5844,N_3702,N_3086);
xnor U5845 (N_5845,N_2699,N_2905);
nor U5846 (N_5846,N_3630,N_2122);
or U5847 (N_5847,N_2660,N_2620);
and U5848 (N_5848,N_2951,N_2435);
or U5849 (N_5849,N_3723,N_2727);
nand U5850 (N_5850,N_2196,N_3722);
and U5851 (N_5851,N_2065,N_3989);
nand U5852 (N_5852,N_3805,N_3195);
nand U5853 (N_5853,N_2000,N_3921);
nand U5854 (N_5854,N_2625,N_2464);
nand U5855 (N_5855,N_3320,N_3604);
nor U5856 (N_5856,N_2092,N_2696);
or U5857 (N_5857,N_3873,N_2423);
nor U5858 (N_5858,N_2625,N_2872);
or U5859 (N_5859,N_2657,N_2005);
or U5860 (N_5860,N_3835,N_2128);
nand U5861 (N_5861,N_2330,N_3415);
nor U5862 (N_5862,N_2989,N_2568);
nand U5863 (N_5863,N_3820,N_3342);
or U5864 (N_5864,N_3362,N_3236);
nand U5865 (N_5865,N_3666,N_3625);
nand U5866 (N_5866,N_3015,N_3651);
or U5867 (N_5867,N_3464,N_3933);
and U5868 (N_5868,N_3725,N_3927);
nor U5869 (N_5869,N_2293,N_2721);
nor U5870 (N_5870,N_2987,N_2459);
or U5871 (N_5871,N_3450,N_3766);
nor U5872 (N_5872,N_2201,N_3350);
or U5873 (N_5873,N_2465,N_2594);
and U5874 (N_5874,N_3952,N_2971);
nor U5875 (N_5875,N_3511,N_3323);
nand U5876 (N_5876,N_2739,N_2662);
nor U5877 (N_5877,N_2052,N_3680);
nor U5878 (N_5878,N_3130,N_3705);
and U5879 (N_5879,N_2482,N_2166);
nand U5880 (N_5880,N_2858,N_3003);
nand U5881 (N_5881,N_2746,N_2833);
xnor U5882 (N_5882,N_2676,N_2260);
or U5883 (N_5883,N_2322,N_3333);
nor U5884 (N_5884,N_2951,N_2889);
xor U5885 (N_5885,N_3632,N_2543);
nor U5886 (N_5886,N_3975,N_3883);
xnor U5887 (N_5887,N_3794,N_3978);
or U5888 (N_5888,N_3678,N_3688);
nand U5889 (N_5889,N_3934,N_3488);
or U5890 (N_5890,N_2077,N_3867);
xor U5891 (N_5891,N_3523,N_2245);
xnor U5892 (N_5892,N_3355,N_2161);
or U5893 (N_5893,N_3831,N_2893);
nand U5894 (N_5894,N_2754,N_3235);
xor U5895 (N_5895,N_2452,N_2102);
or U5896 (N_5896,N_2126,N_2901);
and U5897 (N_5897,N_2410,N_3652);
nor U5898 (N_5898,N_3420,N_3111);
and U5899 (N_5899,N_3021,N_3825);
nor U5900 (N_5900,N_2109,N_3206);
or U5901 (N_5901,N_3284,N_3215);
and U5902 (N_5902,N_3814,N_2830);
nor U5903 (N_5903,N_2025,N_3764);
nor U5904 (N_5904,N_3243,N_2357);
nand U5905 (N_5905,N_3449,N_2926);
nand U5906 (N_5906,N_3613,N_3636);
nand U5907 (N_5907,N_2481,N_3675);
and U5908 (N_5908,N_3215,N_2113);
or U5909 (N_5909,N_3472,N_3245);
xnor U5910 (N_5910,N_2360,N_2042);
nor U5911 (N_5911,N_2538,N_2888);
nor U5912 (N_5912,N_3025,N_2945);
and U5913 (N_5913,N_2747,N_2675);
nor U5914 (N_5914,N_3171,N_3006);
and U5915 (N_5915,N_3831,N_2662);
xnor U5916 (N_5916,N_3124,N_2327);
nor U5917 (N_5917,N_2883,N_2702);
and U5918 (N_5918,N_2858,N_3431);
or U5919 (N_5919,N_3770,N_3155);
and U5920 (N_5920,N_3735,N_2466);
xor U5921 (N_5921,N_3109,N_2276);
xor U5922 (N_5922,N_2734,N_3714);
and U5923 (N_5923,N_3023,N_3486);
and U5924 (N_5924,N_3765,N_3146);
xor U5925 (N_5925,N_3456,N_3658);
and U5926 (N_5926,N_3564,N_2203);
and U5927 (N_5927,N_3304,N_2407);
or U5928 (N_5928,N_2966,N_3728);
xnor U5929 (N_5929,N_2371,N_2218);
nor U5930 (N_5930,N_3228,N_3104);
or U5931 (N_5931,N_2804,N_2070);
nor U5932 (N_5932,N_3982,N_3674);
and U5933 (N_5933,N_2432,N_3444);
xor U5934 (N_5934,N_2854,N_2195);
nand U5935 (N_5935,N_3526,N_3939);
xnor U5936 (N_5936,N_3411,N_2603);
and U5937 (N_5937,N_3835,N_3478);
or U5938 (N_5938,N_3023,N_2679);
nor U5939 (N_5939,N_2754,N_2065);
and U5940 (N_5940,N_2038,N_3981);
xor U5941 (N_5941,N_3190,N_3586);
and U5942 (N_5942,N_2637,N_2595);
nor U5943 (N_5943,N_3953,N_3932);
or U5944 (N_5944,N_3920,N_2863);
or U5945 (N_5945,N_3238,N_2722);
or U5946 (N_5946,N_3867,N_3045);
nand U5947 (N_5947,N_2951,N_3963);
nand U5948 (N_5948,N_2688,N_2338);
xor U5949 (N_5949,N_2862,N_2249);
nand U5950 (N_5950,N_3936,N_2005);
and U5951 (N_5951,N_3838,N_2191);
nor U5952 (N_5952,N_3458,N_2400);
or U5953 (N_5953,N_3708,N_3566);
nand U5954 (N_5954,N_3309,N_3402);
xor U5955 (N_5955,N_3539,N_3808);
or U5956 (N_5956,N_2740,N_2505);
nor U5957 (N_5957,N_2825,N_3106);
nor U5958 (N_5958,N_2511,N_2883);
and U5959 (N_5959,N_3061,N_2167);
nand U5960 (N_5960,N_3398,N_3209);
and U5961 (N_5961,N_3560,N_2891);
and U5962 (N_5962,N_2171,N_2297);
nand U5963 (N_5963,N_3321,N_3473);
nor U5964 (N_5964,N_3302,N_2215);
or U5965 (N_5965,N_3795,N_3456);
nor U5966 (N_5966,N_2903,N_2183);
or U5967 (N_5967,N_2618,N_3201);
xor U5968 (N_5968,N_2471,N_2502);
and U5969 (N_5969,N_3466,N_2437);
and U5970 (N_5970,N_3526,N_3696);
and U5971 (N_5971,N_3870,N_2704);
nand U5972 (N_5972,N_3158,N_3549);
and U5973 (N_5973,N_3378,N_3392);
nand U5974 (N_5974,N_2464,N_3125);
nand U5975 (N_5975,N_2378,N_2277);
xor U5976 (N_5976,N_3641,N_2464);
nand U5977 (N_5977,N_3990,N_3435);
and U5978 (N_5978,N_2139,N_3238);
and U5979 (N_5979,N_2509,N_3090);
xor U5980 (N_5980,N_3802,N_3004);
xnor U5981 (N_5981,N_3486,N_2550);
and U5982 (N_5982,N_2972,N_2608);
nor U5983 (N_5983,N_3941,N_2541);
nand U5984 (N_5984,N_2073,N_3242);
nand U5985 (N_5985,N_2639,N_2992);
nand U5986 (N_5986,N_3802,N_3135);
xnor U5987 (N_5987,N_3295,N_2298);
nor U5988 (N_5988,N_2122,N_2999);
nor U5989 (N_5989,N_3995,N_3514);
or U5990 (N_5990,N_3353,N_3412);
or U5991 (N_5991,N_3769,N_3729);
and U5992 (N_5992,N_2220,N_3616);
and U5993 (N_5993,N_3841,N_2332);
nand U5994 (N_5994,N_2416,N_2873);
and U5995 (N_5995,N_2294,N_2811);
nor U5996 (N_5996,N_3498,N_3171);
nor U5997 (N_5997,N_3002,N_3018);
nor U5998 (N_5998,N_2915,N_3415);
and U5999 (N_5999,N_3896,N_3627);
and U6000 (N_6000,N_4828,N_4174);
or U6001 (N_6001,N_4794,N_5771);
or U6002 (N_6002,N_5868,N_4313);
and U6003 (N_6003,N_5361,N_4844);
nand U6004 (N_6004,N_5305,N_5393);
nand U6005 (N_6005,N_4860,N_5654);
or U6006 (N_6006,N_5022,N_4172);
and U6007 (N_6007,N_4231,N_5185);
or U6008 (N_6008,N_4964,N_4131);
nand U6009 (N_6009,N_5324,N_4102);
or U6010 (N_6010,N_5161,N_5245);
nand U6011 (N_6011,N_4729,N_5117);
nand U6012 (N_6012,N_5552,N_4104);
and U6013 (N_6013,N_5299,N_5559);
xor U6014 (N_6014,N_4521,N_4517);
and U6015 (N_6015,N_4795,N_4241);
nor U6016 (N_6016,N_4665,N_4380);
nand U6017 (N_6017,N_4444,N_5956);
nand U6018 (N_6018,N_5703,N_4190);
xor U6019 (N_6019,N_5809,N_5807);
and U6020 (N_6020,N_4976,N_5846);
xnor U6021 (N_6021,N_4737,N_5275);
and U6022 (N_6022,N_5668,N_4648);
nor U6023 (N_6023,N_5591,N_4660);
nand U6024 (N_6024,N_4759,N_4910);
nor U6025 (N_6025,N_5387,N_4146);
nor U6026 (N_6026,N_4956,N_4059);
nor U6027 (N_6027,N_4686,N_4462);
and U6028 (N_6028,N_5861,N_5561);
and U6029 (N_6029,N_4039,N_4314);
or U6030 (N_6030,N_5318,N_5611);
nor U6031 (N_6031,N_4381,N_5887);
nand U6032 (N_6032,N_4062,N_4012);
and U6033 (N_6033,N_5336,N_5996);
or U6034 (N_6034,N_5761,N_5293);
xnor U6035 (N_6035,N_5626,N_4133);
xnor U6036 (N_6036,N_4983,N_5939);
xor U6037 (N_6037,N_5075,N_4476);
nand U6038 (N_6038,N_5953,N_5995);
and U6039 (N_6039,N_4108,N_4985);
xnor U6040 (N_6040,N_4969,N_5148);
or U6041 (N_6041,N_4198,N_5268);
or U6042 (N_6042,N_4838,N_4638);
or U6043 (N_6043,N_4487,N_4590);
or U6044 (N_6044,N_4643,N_5532);
nor U6045 (N_6045,N_4178,N_5432);
nor U6046 (N_6046,N_5676,N_5090);
nand U6047 (N_6047,N_4689,N_5456);
or U6048 (N_6048,N_5933,N_4341);
nor U6049 (N_6049,N_4640,N_5620);
xor U6050 (N_6050,N_5854,N_4669);
xnor U6051 (N_6051,N_5828,N_5970);
or U6052 (N_6052,N_5764,N_4454);
xnor U6053 (N_6053,N_5327,N_5345);
nand U6054 (N_6054,N_5280,N_4701);
nand U6055 (N_6055,N_5758,N_4813);
nand U6056 (N_6056,N_5216,N_5859);
nor U6057 (N_6057,N_5811,N_4673);
and U6058 (N_6058,N_4988,N_5052);
and U6059 (N_6059,N_4322,N_4087);
and U6060 (N_6060,N_5012,N_4412);
nor U6061 (N_6061,N_5973,N_4579);
nor U6062 (N_6062,N_5094,N_4625);
xor U6063 (N_6063,N_5001,N_5158);
nand U6064 (N_6064,N_4365,N_5135);
and U6065 (N_6065,N_4709,N_4886);
xnor U6066 (N_6066,N_5834,N_5572);
or U6067 (N_6067,N_5778,N_5752);
nand U6068 (N_6068,N_4465,N_4175);
xor U6069 (N_6069,N_4327,N_4503);
and U6070 (N_6070,N_4748,N_5715);
nor U6071 (N_6071,N_5333,N_5139);
nand U6072 (N_6072,N_4716,N_5258);
nor U6073 (N_6073,N_5428,N_4698);
or U6074 (N_6074,N_4505,N_4280);
nor U6075 (N_6075,N_5741,N_4200);
nand U6076 (N_6076,N_4905,N_5013);
nand U6077 (N_6077,N_4741,N_5617);
nor U6078 (N_6078,N_5233,N_4552);
nor U6079 (N_6079,N_5922,N_5189);
xor U6080 (N_6080,N_5290,N_5507);
and U6081 (N_6081,N_5177,N_5994);
nand U6082 (N_6082,N_5365,N_5912);
or U6083 (N_6083,N_4491,N_4613);
nand U6084 (N_6084,N_5488,N_5546);
nor U6085 (N_6085,N_4308,N_5915);
or U6086 (N_6086,N_5307,N_5959);
and U6087 (N_6087,N_5653,N_5873);
nand U6088 (N_6088,N_4654,N_5621);
nor U6089 (N_6089,N_5081,N_5105);
or U6090 (N_6090,N_4268,N_4867);
and U6091 (N_6091,N_4077,N_4081);
xor U6092 (N_6092,N_5857,N_5501);
nand U6093 (N_6093,N_5582,N_5543);
and U6094 (N_6094,N_4763,N_5029);
and U6095 (N_6095,N_5150,N_5079);
or U6096 (N_6096,N_5864,N_5567);
and U6097 (N_6097,N_5844,N_5943);
and U6098 (N_6098,N_5792,N_5401);
or U6099 (N_6099,N_4255,N_5149);
or U6100 (N_6100,N_5242,N_4420);
nand U6101 (N_6101,N_4740,N_4697);
and U6102 (N_6102,N_5091,N_5418);
and U6103 (N_6103,N_4968,N_5250);
and U6104 (N_6104,N_4130,N_5583);
or U6105 (N_6105,N_5821,N_4219);
and U6106 (N_6106,N_5558,N_5948);
and U6107 (N_6107,N_5226,N_5754);
and U6108 (N_6108,N_5030,N_4150);
xor U6109 (N_6109,N_4068,N_5000);
or U6110 (N_6110,N_4941,N_5749);
nor U6111 (N_6111,N_4391,N_4815);
nor U6112 (N_6112,N_5313,N_5831);
nand U6113 (N_6113,N_4708,N_5151);
and U6114 (N_6114,N_4028,N_5795);
nand U6115 (N_6115,N_4728,N_5202);
nor U6116 (N_6116,N_5267,N_4591);
or U6117 (N_6117,N_4368,N_4753);
and U6118 (N_6118,N_5057,N_5731);
or U6119 (N_6119,N_4293,N_5332);
xor U6120 (N_6120,N_5717,N_5183);
or U6121 (N_6121,N_4540,N_5101);
nand U6122 (N_6122,N_5157,N_4967);
xnor U6123 (N_6123,N_4383,N_5706);
nor U6124 (N_6124,N_4186,N_5634);
xor U6125 (N_6125,N_5493,N_5092);
and U6126 (N_6126,N_5145,N_5722);
xnor U6127 (N_6127,N_4253,N_4713);
nor U6128 (N_6128,N_5503,N_5154);
or U6129 (N_6129,N_4113,N_4755);
xnor U6130 (N_6130,N_5575,N_5011);
and U6131 (N_6131,N_4156,N_4203);
and U6132 (N_6132,N_4467,N_4205);
or U6133 (N_6133,N_4548,N_4419);
or U6134 (N_6134,N_4774,N_4829);
nand U6135 (N_6135,N_4123,N_5460);
nand U6136 (N_6136,N_4916,N_4334);
and U6137 (N_6137,N_4263,N_4287);
nand U6138 (N_6138,N_5866,N_4355);
or U6139 (N_6139,N_4918,N_4496);
nor U6140 (N_6140,N_4023,N_4536);
xnor U6141 (N_6141,N_4196,N_5707);
or U6142 (N_6142,N_5407,N_4695);
and U6143 (N_6143,N_4047,N_5672);
and U6144 (N_6144,N_4237,N_4188);
nor U6145 (N_6145,N_5195,N_4637);
xor U6146 (N_6146,N_5627,N_4398);
or U6147 (N_6147,N_5952,N_5845);
nand U6148 (N_6148,N_5645,N_5006);
and U6149 (N_6149,N_4170,N_5727);
nand U6150 (N_6150,N_4276,N_4408);
or U6151 (N_6151,N_4064,N_5641);
nor U6152 (N_6152,N_5381,N_5783);
nand U6153 (N_6153,N_4471,N_4550);
nor U6154 (N_6154,N_4804,N_4187);
and U6155 (N_6155,N_4746,N_5466);
or U6156 (N_6156,N_5171,N_4776);
or U6157 (N_6157,N_4567,N_4778);
and U6158 (N_6158,N_4224,N_4635);
nand U6159 (N_6159,N_4636,N_5270);
nor U6160 (N_6160,N_5023,N_4814);
or U6161 (N_6161,N_5334,N_5093);
nor U6162 (N_6162,N_5298,N_5941);
nor U6163 (N_6163,N_4523,N_5056);
and U6164 (N_6164,N_5132,N_4090);
xnor U6165 (N_6165,N_4499,N_5253);
and U6166 (N_6166,N_4451,N_4406);
nand U6167 (N_6167,N_5455,N_4892);
and U6168 (N_6168,N_4769,N_5705);
nor U6169 (N_6169,N_5277,N_5820);
and U6170 (N_6170,N_5523,N_5475);
xor U6171 (N_6171,N_4456,N_4015);
xnor U6172 (N_6172,N_4250,N_5113);
nand U6173 (N_6173,N_4714,N_4233);
and U6174 (N_6174,N_4010,N_4859);
and U6175 (N_6175,N_4620,N_4576);
xor U6176 (N_6176,N_4880,N_4157);
and U6177 (N_6177,N_4630,N_4018);
xnor U6178 (N_6178,N_5659,N_4588);
nor U6179 (N_6179,N_4779,N_4899);
and U6180 (N_6180,N_4831,N_4928);
nor U6181 (N_6181,N_5977,N_4717);
xnor U6182 (N_6182,N_4390,N_4619);
xor U6183 (N_6183,N_5851,N_5812);
or U6184 (N_6184,N_4080,N_5961);
nor U6185 (N_6185,N_4480,N_5817);
xor U6186 (N_6186,N_5082,N_4682);
nand U6187 (N_6187,N_5457,N_4711);
and U6188 (N_6188,N_5062,N_4193);
nor U6189 (N_6189,N_4020,N_5289);
or U6190 (N_6190,N_5597,N_5096);
and U6191 (N_6191,N_4299,N_4938);
and U6192 (N_6192,N_4762,N_5147);
and U6193 (N_6193,N_4587,N_5286);
and U6194 (N_6194,N_4009,N_4306);
nand U6195 (N_6195,N_5719,N_4158);
xnor U6196 (N_6196,N_5010,N_5618);
nand U6197 (N_6197,N_4751,N_5122);
nand U6198 (N_6198,N_4050,N_4242);
xor U6199 (N_6199,N_5048,N_4977);
or U6200 (N_6200,N_4897,N_5037);
nor U6201 (N_6201,N_5784,N_5648);
and U6202 (N_6202,N_4783,N_5476);
or U6203 (N_6203,N_4288,N_4824);
or U6204 (N_6204,N_5398,N_4301);
xnor U6205 (N_6205,N_4626,N_5077);
nor U6206 (N_6206,N_5893,N_5038);
nand U6207 (N_6207,N_4633,N_5782);
and U6208 (N_6208,N_4091,N_4302);
xor U6209 (N_6209,N_5163,N_4519);
and U6210 (N_6210,N_5284,N_4315);
nand U6211 (N_6211,N_5197,N_4931);
nor U6212 (N_6212,N_4904,N_4307);
xnor U6213 (N_6213,N_4605,N_5599);
xor U6214 (N_6214,N_4166,N_4346);
nand U6215 (N_6215,N_4340,N_5003);
and U6216 (N_6216,N_5326,N_5569);
xnor U6217 (N_6217,N_4374,N_4128);
xnor U6218 (N_6218,N_5649,N_5292);
nand U6219 (N_6219,N_4442,N_4845);
nand U6220 (N_6220,N_4063,N_5067);
nor U6221 (N_6221,N_5716,N_4044);
xor U6222 (N_6222,N_4258,N_5417);
or U6223 (N_6223,N_4337,N_4092);
nor U6224 (N_6224,N_5076,N_4959);
nor U6225 (N_6225,N_5607,N_5487);
nor U6226 (N_6226,N_5913,N_5657);
xnor U6227 (N_6227,N_5423,N_4386);
and U6228 (N_6228,N_5304,N_4664);
xnor U6229 (N_6229,N_4864,N_5064);
nor U6230 (N_6230,N_4600,N_5872);
xor U6231 (N_6231,N_4275,N_4464);
xor U6232 (N_6232,N_5837,N_5108);
or U6233 (N_6233,N_4220,N_5232);
or U6234 (N_6234,N_5380,N_5917);
nand U6235 (N_6235,N_5880,N_4026);
and U6236 (N_6236,N_4019,N_4888);
xor U6237 (N_6237,N_5040,N_5496);
or U6238 (N_6238,N_5414,N_4396);
and U6239 (N_6239,N_5789,N_4411);
or U6240 (N_6240,N_5083,N_5505);
and U6241 (N_6241,N_4703,N_5200);
xnor U6242 (N_6242,N_5955,N_4097);
and U6243 (N_6243,N_5230,N_5842);
or U6244 (N_6244,N_4962,N_4216);
and U6245 (N_6245,N_5103,N_5684);
and U6246 (N_6246,N_4447,N_4428);
or U6247 (N_6247,N_5254,N_4176);
nor U6248 (N_6248,N_4681,N_4898);
xnor U6249 (N_6249,N_5279,N_5748);
xor U6250 (N_6250,N_4883,N_4184);
and U6251 (N_6251,N_5489,N_5060);
or U6252 (N_6252,N_4510,N_5382);
or U6253 (N_6253,N_5447,N_4940);
xor U6254 (N_6254,N_4564,N_5427);
xor U6255 (N_6255,N_4614,N_5848);
nor U6256 (N_6256,N_4971,N_4816);
nand U6257 (N_6257,N_5046,N_4434);
nor U6258 (N_6258,N_5322,N_4777);
nor U6259 (N_6259,N_4033,N_5220);
nand U6260 (N_6260,N_4954,N_5689);
and U6261 (N_6261,N_4259,N_4808);
nor U6262 (N_6262,N_5107,N_5840);
nor U6263 (N_6263,N_4734,N_4326);
or U6264 (N_6264,N_4827,N_5058);
xor U6265 (N_6265,N_4744,N_4901);
nor U6266 (N_6266,N_5796,N_5378);
or U6267 (N_6267,N_4129,N_5315);
nor U6268 (N_6268,N_4192,N_5188);
xor U6269 (N_6269,N_5517,N_4852);
nor U6270 (N_6270,N_4501,N_5947);
nand U6271 (N_6271,N_4295,N_4359);
and U6272 (N_6272,N_4754,N_4691);
and U6273 (N_6273,N_4209,N_4448);
or U6274 (N_6274,N_5997,N_5436);
or U6275 (N_6275,N_4520,N_4878);
and U6276 (N_6276,N_4847,N_5344);
nand U6277 (N_6277,N_5410,N_4425);
or U6278 (N_6278,N_5738,N_4376);
or U6279 (N_6279,N_5153,N_5445);
nor U6280 (N_6280,N_5622,N_4134);
nor U6281 (N_6281,N_4001,N_5078);
xor U6282 (N_6282,N_4538,N_5766);
or U6283 (N_6283,N_5337,N_4094);
and U6284 (N_6284,N_4054,N_5498);
or U6285 (N_6285,N_4357,N_5235);
and U6286 (N_6286,N_4082,N_5688);
nand U6287 (N_6287,N_5182,N_5041);
xnor U6288 (N_6288,N_5579,N_5699);
and U6289 (N_6289,N_4723,N_5679);
and U6290 (N_6290,N_4234,N_5463);
nor U6291 (N_6291,N_4707,N_5562);
and U6292 (N_6292,N_5349,N_5743);
nand U6293 (N_6293,N_5317,N_4950);
xnor U6294 (N_6294,N_4333,N_5372);
nor U6295 (N_6295,N_4668,N_4623);
and U6296 (N_6296,N_4830,N_5144);
nor U6297 (N_6297,N_4049,N_4811);
or U6298 (N_6298,N_4211,N_4949);
or U6299 (N_6299,N_4994,N_5736);
nor U6300 (N_6300,N_5850,N_5369);
or U6301 (N_6301,N_5063,N_5898);
nand U6302 (N_6302,N_4803,N_5394);
nand U6303 (N_6303,N_5824,N_4116);
xor U6304 (N_6304,N_4072,N_4217);
nand U6305 (N_6305,N_4181,N_4180);
nor U6306 (N_6306,N_5966,N_5187);
nor U6307 (N_6307,N_5097,N_5934);
and U6308 (N_6308,N_4126,N_4481);
nand U6309 (N_6309,N_5512,N_5020);
and U6310 (N_6310,N_5155,N_4733);
or U6311 (N_6311,N_5392,N_5734);
xnor U6312 (N_6312,N_4765,N_5390);
nor U6313 (N_6313,N_5021,N_4943);
nand U6314 (N_6314,N_5545,N_4992);
or U6315 (N_6315,N_5603,N_4749);
and U6316 (N_6316,N_4972,N_5613);
nor U6317 (N_6317,N_4036,N_4024);
and U6318 (N_6318,N_4432,N_5729);
nor U6319 (N_6319,N_5089,N_5890);
and U6320 (N_6320,N_5309,N_4244);
xnor U6321 (N_6321,N_4975,N_5350);
and U6322 (N_6322,N_4553,N_4747);
xnor U6323 (N_6323,N_5830,N_5160);
xor U6324 (N_6324,N_4926,N_4629);
xor U6325 (N_6325,N_5491,N_4479);
and U6326 (N_6326,N_4658,N_5801);
nor U6327 (N_6327,N_4163,N_4282);
xor U6328 (N_6328,N_5469,N_4011);
nand U6329 (N_6329,N_5112,N_5536);
or U6330 (N_6330,N_5711,N_4690);
or U6331 (N_6331,N_4861,N_4118);
xor U6332 (N_6332,N_4902,N_4602);
or U6333 (N_6333,N_5265,N_4284);
xnor U6334 (N_6334,N_4796,N_4822);
or U6335 (N_6335,N_4226,N_4378);
nor U6336 (N_6336,N_5847,N_4030);
nor U6337 (N_6337,N_4431,N_4850);
and U6338 (N_6338,N_4165,N_4497);
xor U6339 (N_6339,N_4109,N_5515);
nand U6340 (N_6340,N_4849,N_4727);
xnor U6341 (N_6341,N_5544,N_4397);
nor U6342 (N_6342,N_5207,N_4627);
or U6343 (N_6343,N_5798,N_4788);
nor U6344 (N_6344,N_5243,N_4305);
and U6345 (N_6345,N_5574,N_5992);
and U6346 (N_6346,N_4210,N_5281);
and U6347 (N_6347,N_5377,N_5643);
nand U6348 (N_6348,N_5363,N_5673);
nand U6349 (N_6349,N_4912,N_5896);
and U6350 (N_6350,N_4700,N_5629);
nand U6351 (N_6351,N_4580,N_5773);
nor U6352 (N_6352,N_4110,N_5500);
nand U6353 (N_6353,N_5573,N_4539);
xnor U6354 (N_6354,N_5533,N_5589);
or U6355 (N_6355,N_5215,N_4352);
xnor U6356 (N_6356,N_5271,N_4323);
nand U6357 (N_6357,N_5320,N_4865);
or U6358 (N_6358,N_4393,N_4141);
or U6359 (N_6359,N_5520,N_4167);
nor U6360 (N_6360,N_5009,N_4651);
xnor U6361 (N_6361,N_5780,N_4114);
or U6362 (N_6362,N_4093,N_4443);
xor U6363 (N_6363,N_5902,N_5329);
and U6364 (N_6364,N_5894,N_4269);
nand U6365 (N_6365,N_4429,N_4199);
nor U6366 (N_6366,N_4639,N_4834);
nand U6367 (N_6367,N_5221,N_4143);
xor U6368 (N_6368,N_4862,N_4485);
nand U6369 (N_6369,N_4595,N_4270);
nor U6370 (N_6370,N_4616,N_5695);
nor U6371 (N_6371,N_4688,N_4704);
nand U6372 (N_6372,N_5946,N_5762);
and U6373 (N_6373,N_4607,N_4421);
nor U6374 (N_6374,N_4678,N_4364);
and U6375 (N_6375,N_4601,N_5480);
and U6376 (N_6376,N_5296,N_5341);
xnor U6377 (N_6377,N_4369,N_5264);
xnor U6378 (N_6378,N_5087,N_5167);
and U6379 (N_6379,N_5192,N_4281);
nand U6380 (N_6380,N_4530,N_4122);
nand U6381 (N_6381,N_5528,N_4921);
or U6382 (N_6382,N_4649,N_4509);
or U6383 (N_6383,N_5218,N_5980);
xnor U6384 (N_6384,N_4201,N_4608);
xor U6385 (N_6385,N_4603,N_5450);
nor U6386 (N_6386,N_4162,N_4652);
or U6387 (N_6387,N_5301,N_4002);
nor U6388 (N_6388,N_5682,N_4215);
and U6389 (N_6389,N_5467,N_5303);
or U6390 (N_6390,N_5055,N_4449);
or U6391 (N_6391,N_5895,N_4872);
nor U6392 (N_6392,N_4913,N_5963);
or U6393 (N_6393,N_4631,N_5609);
and U6394 (N_6394,N_4998,N_5004);
nand U6395 (N_6395,N_5581,N_5359);
or U6396 (N_6396,N_5213,N_4854);
nor U6397 (N_6397,N_5026,N_5563);
or U6398 (N_6398,N_4379,N_4915);
nor U6399 (N_6399,N_5045,N_5708);
and U6400 (N_6400,N_4742,N_4303);
and U6401 (N_6401,N_5196,N_5273);
or U6402 (N_6402,N_4786,N_4088);
nand U6403 (N_6403,N_5179,N_5714);
xnor U6404 (N_6404,N_4646,N_5138);
and U6405 (N_6405,N_4570,N_4848);
xor U6406 (N_6406,N_5655,N_4535);
nand U6407 (N_6407,N_4653,N_5519);
nand U6408 (N_6408,N_5477,N_5863);
or U6409 (N_6409,N_4384,N_5767);
xnor U6410 (N_6410,N_4885,N_5400);
or U6411 (N_6411,N_4545,N_5663);
nor U6412 (N_6412,N_4936,N_4657);
or U6413 (N_6413,N_4490,N_4641);
or U6414 (N_6414,N_5162,N_5686);
and U6415 (N_6415,N_5355,N_5325);
nor U6416 (N_6416,N_4659,N_5884);
or U6417 (N_6417,N_4349,N_4843);
or U6418 (N_6418,N_4946,N_4264);
nand U6419 (N_6419,N_5808,N_5123);
and U6420 (N_6420,N_4581,N_5819);
nor U6421 (N_6421,N_5701,N_4136);
xnor U6422 (N_6422,N_4495,N_5619);
nand U6423 (N_6423,N_4556,N_5086);
or U6424 (N_6424,N_4524,N_5937);
xor U6425 (N_6425,N_5951,N_4450);
or U6426 (N_6426,N_5988,N_4817);
xor U6427 (N_6427,N_5343,N_4076);
xnor U6428 (N_6428,N_4922,N_5364);
and U6429 (N_6429,N_4267,N_5968);
nand U6430 (N_6430,N_4500,N_4621);
nor U6431 (N_6431,N_4101,N_5276);
or U6432 (N_6432,N_4870,N_4773);
or U6433 (N_6433,N_4182,N_4240);
and U6434 (N_6434,N_4189,N_4430);
or U6435 (N_6435,N_4532,N_5805);
or U6436 (N_6436,N_5257,N_4407);
or U6437 (N_6437,N_5669,N_4833);
nor U6438 (N_6438,N_5788,N_5438);
nor U6439 (N_6439,N_5239,N_5100);
and U6440 (N_6440,N_5206,N_5730);
and U6441 (N_6441,N_4324,N_4492);
or U6442 (N_6442,N_5005,N_5910);
or U6443 (N_6443,N_5786,N_4452);
and U6444 (N_6444,N_4161,N_5535);
or U6445 (N_6445,N_5129,N_4426);
and U6446 (N_6446,N_4212,N_4982);
and U6447 (N_6447,N_4331,N_4596);
or U6448 (N_6448,N_5357,N_5877);
nor U6449 (N_6449,N_5485,N_4266);
or U6450 (N_6450,N_4671,N_5605);
or U6451 (N_6451,N_4086,N_5111);
nand U6452 (N_6452,N_4153,N_5800);
and U6453 (N_6453,N_5482,N_4469);
nor U6454 (N_6454,N_4584,N_5667);
nand U6455 (N_6455,N_4067,N_5146);
nand U6456 (N_6456,N_5335,N_5990);
and U6457 (N_6457,N_4721,N_4821);
or U6458 (N_6458,N_4702,N_4385);
nor U6459 (N_6459,N_5744,N_4863);
nand U6460 (N_6460,N_4144,N_5550);
nand U6461 (N_6461,N_5537,N_4195);
and U6462 (N_6462,N_4223,N_5027);
and U6463 (N_6463,N_5640,N_5770);
nand U6464 (N_6464,N_5972,N_4835);
nor U6465 (N_6465,N_4243,N_4547);
xnor U6466 (N_6466,N_4502,N_5531);
and U6467 (N_6467,N_4100,N_5914);
or U6468 (N_6468,N_4705,N_5384);
nand U6469 (N_6469,N_4515,N_5449);
or U6470 (N_6470,N_5600,N_5924);
and U6471 (N_6471,N_4083,N_4839);
nor U6472 (N_6472,N_5652,N_5180);
and U6473 (N_6473,N_5577,N_5124);
xor U6474 (N_6474,N_5404,N_4750);
nor U6475 (N_6475,N_4731,N_5223);
nand U6476 (N_6476,N_4296,N_4000);
nand U6477 (N_6477,N_4789,N_4722);
xnor U6478 (N_6478,N_4504,N_4286);
or U6479 (N_6479,N_5746,N_4875);
or U6480 (N_6480,N_5069,N_5897);
and U6481 (N_6481,N_5492,N_5891);
xor U6482 (N_6482,N_5035,N_4055);
nor U6483 (N_6483,N_5745,N_4260);
xor U6484 (N_6484,N_4300,N_5201);
and U6485 (N_6485,N_4650,N_5495);
or U6486 (N_6486,N_4236,N_5047);
nor U6487 (N_6487,N_4472,N_5109);
or U6488 (N_6488,N_4712,N_5424);
and U6489 (N_6489,N_5367,N_5799);
nand U6490 (N_6490,N_4316,N_5718);
nand U6491 (N_6491,N_4057,N_5806);
xor U6492 (N_6492,N_4348,N_4842);
nand U6493 (N_6493,N_4404,N_5291);
nand U6494 (N_6494,N_5461,N_4311);
and U6495 (N_6495,N_4035,N_5302);
nor U6496 (N_6496,N_4433,N_5635);
xnor U6497 (N_6497,N_5539,N_5133);
xor U6498 (N_6498,N_4877,N_4785);
xnor U6499 (N_6499,N_4836,N_4760);
and U6500 (N_6500,N_5656,N_5288);
nand U6501 (N_6501,N_5373,N_4526);
xor U6502 (N_6502,N_4417,N_4693);
nor U6503 (N_6503,N_5921,N_5259);
or U6504 (N_6504,N_4642,N_4889);
nor U6505 (N_6505,N_4016,N_5590);
nor U6506 (N_6506,N_5043,N_4079);
or U6507 (N_6507,N_5940,N_5644);
xor U6508 (N_6508,N_5983,N_4792);
nor U6509 (N_6509,N_5838,N_5074);
xor U6510 (N_6510,N_5143,N_4154);
or U6511 (N_6511,N_4884,N_5646);
xor U6512 (N_6512,N_4818,N_5547);
nor U6513 (N_6513,N_4229,N_4272);
nor U6514 (N_6514,N_4251,N_5642);
nand U6515 (N_6515,N_5278,N_4837);
and U6516 (N_6516,N_4720,N_5905);
nand U6517 (N_6517,N_4078,N_4159);
nand U6518 (N_6518,N_5568,N_4249);
nor U6519 (N_6519,N_5464,N_4202);
nand U6520 (N_6520,N_4413,N_5785);
xor U6521 (N_6521,N_5042,N_4021);
xnor U6522 (N_6522,N_4445,N_4127);
xnor U6523 (N_6523,N_5319,N_4297);
nand U6524 (N_6524,N_4271,N_4670);
xor U6525 (N_6525,N_5237,N_4857);
and U6526 (N_6526,N_5680,N_4423);
and U6527 (N_6527,N_4074,N_4948);
xor U6528 (N_6528,N_5442,N_4981);
nand U6529 (N_6529,N_5169,N_5944);
and U6530 (N_6530,N_4978,N_5061);
and U6531 (N_6531,N_4806,N_4891);
xnor U6532 (N_6532,N_4377,N_5295);
and U6533 (N_6533,N_4684,N_4939);
xnor U6534 (N_6534,N_5370,N_4881);
or U6535 (N_6535,N_5751,N_4218);
and U6536 (N_6536,N_4562,N_4484);
or U6537 (N_6537,N_5231,N_5601);
and U6538 (N_6538,N_5712,N_5310);
or U6539 (N_6539,N_4148,N_4719);
and U6540 (N_6540,N_5612,N_4790);
and U6541 (N_6541,N_4610,N_4466);
and U6542 (N_6542,N_5433,N_5426);
and U6543 (N_6543,N_5697,N_5870);
or U6544 (N_6544,N_5402,N_4577);
nand U6545 (N_6545,N_5639,N_4594);
nor U6546 (N_6546,N_5224,N_4764);
or U6547 (N_6547,N_4132,N_5121);
or U6548 (N_6548,N_5175,N_5750);
or U6549 (N_6549,N_5836,N_5429);
and U6550 (N_6550,N_5678,N_4799);
and U6551 (N_6551,N_4053,N_5584);
xnor U6552 (N_6552,N_4470,N_4388);
or U6553 (N_6553,N_5416,N_4345);
and U6554 (N_6554,N_4565,N_5115);
nand U6555 (N_6555,N_5858,N_5835);
or U6556 (N_6556,N_5234,N_4221);
xnor U6557 (N_6557,N_5978,N_4265);
nand U6558 (N_6558,N_4963,N_4945);
xnor U6559 (N_6559,N_5548,N_5685);
xor U6560 (N_6560,N_5976,N_5514);
nand U6561 (N_6561,N_4771,N_5625);
xor U6562 (N_6562,N_4375,N_4598);
nand U6563 (N_6563,N_4096,N_5986);
nor U6564 (N_6564,N_5769,N_4732);
nor U6565 (N_6565,N_5610,N_4208);
and U6566 (N_6566,N_5159,N_5556);
or U6567 (N_6567,N_5173,N_4960);
xnor U6568 (N_6568,N_4304,N_4781);
nor U6569 (N_6569,N_5028,N_5797);
nand U6570 (N_6570,N_5802,N_4347);
or U6571 (N_6571,N_4791,N_5920);
or U6572 (N_6572,N_4527,N_5595);
nand U6573 (N_6573,N_5208,N_4868);
nand U6574 (N_6574,N_5184,N_5379);
nand U6575 (N_6575,N_5051,N_4599);
nand U6576 (N_6576,N_5238,N_4958);
nand U6577 (N_6577,N_5484,N_5904);
nor U6578 (N_6578,N_5636,N_4310);
nor U6579 (N_6579,N_4457,N_4458);
nand U6580 (N_6580,N_5841,N_5606);
xnor U6581 (N_6581,N_4534,N_4119);
or U6582 (N_6582,N_5521,N_5911);
and U6583 (N_6583,N_5958,N_4225);
nand U6584 (N_6584,N_5578,N_5901);
or U6585 (N_6585,N_4401,N_4593);
xor U6586 (N_6586,N_5790,N_4460);
xor U6587 (N_6587,N_5127,N_5892);
or U6588 (N_6588,N_5181,N_5867);
nor U6589 (N_6589,N_5490,N_5017);
nor U6590 (N_6590,N_4373,N_5486);
xor U6591 (N_6591,N_5389,N_5856);
nor U6592 (N_6592,N_5692,N_5628);
or U6593 (N_6593,N_5142,N_5925);
or U6594 (N_6594,N_4427,N_5479);
xor U6595 (N_6595,N_4046,N_5526);
or U6596 (N_6596,N_5662,N_5509);
xor U6597 (N_6597,N_4974,N_4923);
or U6598 (N_6598,N_4031,N_4952);
or U6599 (N_6599,N_4459,N_4805);
or U6600 (N_6600,N_5964,N_5614);
nand U6601 (N_6601,N_5204,N_5721);
nand U6602 (N_6602,N_5566,N_4061);
nand U6603 (N_6603,N_4784,N_4183);
or U6604 (N_6604,N_4052,N_5888);
and U6605 (N_6605,N_4512,N_4446);
or U6606 (N_6606,N_5677,N_5779);
or U6607 (N_6607,N_4812,N_4371);
xor U6608 (N_6608,N_5513,N_5664);
and U6609 (N_6609,N_5524,N_5282);
nand U6610 (N_6610,N_4647,N_5698);
and U6611 (N_6611,N_5338,N_5666);
nand U6612 (N_6612,N_4436,N_4735);
and U6613 (N_6613,N_5962,N_5598);
and U6614 (N_6614,N_4628,N_4152);
xor U6615 (N_6615,N_5508,N_5131);
and U6616 (N_6616,N_4354,N_5781);
and U6617 (N_6617,N_5979,N_4112);
xor U6618 (N_6618,N_4179,N_4027);
or U6619 (N_6619,N_5312,N_5451);
nor U6620 (N_6620,N_4572,N_5713);
nor U6621 (N_6621,N_5564,N_4489);
xnor U6622 (N_6622,N_4317,N_4770);
xor U6623 (N_6623,N_5272,N_5388);
nor U6624 (N_6624,N_4247,N_4105);
nor U6625 (N_6625,N_4775,N_5985);
and U6626 (N_6626,N_5816,N_4609);
xnor U6627 (N_6627,N_4929,N_4710);
or U6628 (N_6628,N_5459,N_5886);
xnor U6629 (N_6629,N_4394,N_4920);
and U6630 (N_6630,N_5737,N_5916);
xnor U6631 (N_6631,N_4807,N_4942);
xnor U6632 (N_6632,N_5827,N_4761);
and U6633 (N_6633,N_4312,N_5217);
xor U6634 (N_6634,N_4252,N_4586);
and U6635 (N_6635,N_4043,N_4273);
nand U6636 (N_6636,N_5879,N_4667);
nand U6637 (N_6637,N_5346,N_5931);
and U6638 (N_6638,N_4694,N_5554);
nand U6639 (N_6639,N_4900,N_5822);
and U6640 (N_6640,N_5068,N_4191);
nand U6641 (N_6641,N_4825,N_5118);
nand U6642 (N_6642,N_5421,N_4809);
and U6643 (N_6643,N_5395,N_5098);
nor U6644 (N_6644,N_4351,N_5453);
and U6645 (N_6645,N_4937,N_5088);
and U6646 (N_6646,N_5024,N_5425);
nand U6647 (N_6647,N_4544,N_5210);
nor U6648 (N_6648,N_5530,N_4568);
xor U6649 (N_6649,N_4248,N_4066);
nand U6650 (N_6650,N_4468,N_4995);
xnor U6651 (N_6651,N_4400,N_5252);
or U6652 (N_6652,N_5540,N_5529);
or U6653 (N_6653,N_5793,N_4542);
and U6654 (N_6654,N_5787,N_5803);
xnor U6655 (N_6655,N_5923,N_4797);
nor U6656 (N_6656,N_4493,N_4674);
nand U6657 (N_6657,N_4058,N_5441);
nand U6658 (N_6658,N_4506,N_4041);
nor U6659 (N_6659,N_4873,N_5984);
or U6660 (N_6660,N_5263,N_4917);
and U6661 (N_6661,N_4644,N_4463);
and U6662 (N_6662,N_4615,N_5647);
nor U6663 (N_6663,N_5141,N_4160);
or U6664 (N_6664,N_4336,N_5156);
nor U6665 (N_6665,N_5222,N_4283);
or U6666 (N_6666,N_5016,N_5174);
or U6667 (N_6667,N_4823,N_5371);
nor U6668 (N_6668,N_4006,N_5516);
nor U6669 (N_6669,N_4367,N_4793);
or U6670 (N_6670,N_4514,N_5739);
and U6671 (N_6671,N_5982,N_4961);
nand U6672 (N_6672,N_5938,N_4440);
or U6673 (N_6673,N_4947,N_5998);
nand U6674 (N_6674,N_5308,N_5406);
and U6675 (N_6675,N_5283,N_4230);
xor U6676 (N_6676,N_5971,N_5494);
or U6677 (N_6677,N_5732,N_5541);
nand U6678 (N_6678,N_5072,N_5130);
nand U6679 (N_6679,N_4924,N_4073);
or U6680 (N_6680,N_4543,N_5757);
or U6681 (N_6681,N_4679,N_4098);
or U6682 (N_6682,N_5176,N_5095);
or U6683 (N_6683,N_4569,N_5340);
xnor U6684 (N_6684,N_5247,N_4991);
nor U6685 (N_6685,N_5120,N_4048);
xnor U6686 (N_6686,N_5342,N_4895);
nand U6687 (N_6687,N_5229,N_5969);
xor U6688 (N_6688,N_5987,N_5906);
or U6689 (N_6689,N_5576,N_5675);
or U6690 (N_6690,N_4632,N_5033);
nor U6691 (N_6691,N_4139,N_4274);
and U6692 (N_6692,N_4533,N_5261);
nor U6693 (N_6693,N_4149,N_5862);
xnor U6694 (N_6694,N_5849,N_4120);
or U6695 (N_6695,N_5408,N_5919);
and U6696 (N_6696,N_4841,N_4893);
and U6697 (N_6697,N_5683,N_5604);
and U6698 (N_6698,N_5164,N_5899);
xnor U6699 (N_6699,N_4624,N_5632);
nor U6700 (N_6700,N_5869,N_5419);
and U6701 (N_6701,N_4585,N_5165);
nor U6702 (N_6702,N_5439,N_5412);
and U6703 (N_6703,N_4168,N_5518);
and U6704 (N_6704,N_5031,N_4996);
nand U6705 (N_6705,N_5137,N_5772);
nor U6706 (N_6706,N_4724,N_4685);
and U6707 (N_6707,N_4826,N_5823);
nand U6708 (N_6708,N_4339,N_4756);
or U6709 (N_6709,N_5104,N_4618);
xor U6710 (N_6710,N_4291,N_4592);
nand U6711 (N_6711,N_5386,N_4558);
nand U6712 (N_6712,N_5694,N_5960);
or U6713 (N_6713,N_4342,N_5140);
nand U6714 (N_6714,N_5084,N_5205);
nor U6715 (N_6715,N_5474,N_5443);
and U6716 (N_6716,N_4138,N_5360);
xor U6717 (N_6717,N_5383,N_5658);
nand U6718 (N_6718,N_4589,N_4017);
nand U6719 (N_6719,N_5878,N_5981);
and U6720 (N_6720,N_4004,N_5260);
xor U6721 (N_6721,N_5354,N_5759);
and U6722 (N_6722,N_4135,N_5592);
or U6723 (N_6723,N_4075,N_5631);
nor U6724 (N_6724,N_5511,N_4604);
nor U6725 (N_6725,N_5935,N_4987);
or U6726 (N_6726,N_4483,N_4566);
and U6727 (N_6727,N_4894,N_4551);
xnor U6728 (N_6728,N_4993,N_4069);
and U6729 (N_6729,N_4999,N_4245);
nor U6730 (N_6730,N_4951,N_4435);
xor U6731 (N_6731,N_5434,N_5471);
or U6732 (N_6732,N_4482,N_4772);
nor U6733 (N_6733,N_4478,N_5725);
nand U6734 (N_6734,N_4410,N_4403);
xnor U6735 (N_6735,N_4213,N_5316);
or U6736 (N_6736,N_5525,N_4508);
nor U6737 (N_6737,N_4169,N_5470);
or U6738 (N_6738,N_5102,N_5775);
or U6739 (N_6739,N_4855,N_4801);
or U6740 (N_6740,N_5244,N_5248);
xnor U6741 (N_6741,N_5472,N_5356);
and U6742 (N_6742,N_5853,N_4363);
nand U6743 (N_6743,N_5314,N_4925);
or U6744 (N_6744,N_5339,N_5080);
nor U6745 (N_6745,N_5166,N_5720);
and U6746 (N_6746,N_5918,N_4409);
or U6747 (N_6747,N_4738,N_4802);
or U6748 (N_6748,N_4051,N_5538);
nor U6749 (N_6749,N_4424,N_4879);
or U6750 (N_6750,N_4549,N_4798);
nand U6751 (N_6751,N_5852,N_5019);
nor U6752 (N_6752,N_4990,N_5615);
nor U6753 (N_6753,N_5065,N_4040);
nor U6754 (N_6754,N_5050,N_5454);
xnor U6755 (N_6755,N_5212,N_4617);
xnor U6756 (N_6756,N_5908,N_5700);
or U6757 (N_6757,N_5437,N_4869);
nand U6758 (N_6758,N_5693,N_4488);
nor U6759 (N_6759,N_5594,N_4140);
nand U6760 (N_6760,N_4757,N_4513);
nor U6761 (N_6761,N_4279,N_5623);
nand U6762 (N_6762,N_4541,N_5191);
nor U6763 (N_6763,N_5557,N_4656);
and U6764 (N_6764,N_4752,N_4914);
nor U6765 (N_6765,N_5624,N_5638);
or U6766 (N_6766,N_5251,N_5942);
nor U6767 (N_6767,N_4034,N_5882);
xnor U6768 (N_6768,N_5228,N_4405);
nand U6769 (N_6769,N_4362,N_5674);
and U6770 (N_6770,N_4522,N_4699);
nand U6771 (N_6771,N_5950,N_5214);
and U6772 (N_6772,N_5776,N_5194);
and U6773 (N_6773,N_5774,N_5691);
xnor U6774 (N_6774,N_4736,N_5114);
and U6775 (N_6775,N_4903,N_4008);
and U6776 (N_6776,N_4045,N_4121);
xnor U6777 (N_6777,N_5172,N_5285);
and U6778 (N_6778,N_5671,N_5328);
or U6779 (N_6779,N_5929,N_5034);
nor U6780 (N_6780,N_4142,N_5555);
and U6781 (N_6781,N_5499,N_5362);
or U6782 (N_6782,N_4574,N_5128);
or U6783 (N_6783,N_5735,N_4611);
nand U6784 (N_6784,N_4882,N_4655);
or U6785 (N_6785,N_5791,N_4934);
nor U6786 (N_6786,N_5765,N_5768);
xor U6787 (N_6787,N_5403,N_4858);
nor U6788 (N_6788,N_4422,N_5726);
xnor U6789 (N_6789,N_5397,N_5704);
and U6790 (N_6790,N_5932,N_4277);
nand U6791 (N_6791,N_4516,N_5755);
or U6792 (N_6792,N_4832,N_5126);
xor U6793 (N_6793,N_4908,N_4298);
nor U6794 (N_6794,N_4137,N_4453);
nand U6795 (N_6795,N_5763,N_4890);
nor U6796 (N_6796,N_4350,N_5865);
nor U6797 (N_6797,N_5723,N_4278);
xor U6798 (N_6798,N_5039,N_4666);
or U6799 (N_6799,N_5843,N_5875);
nand U6800 (N_6800,N_5287,N_5025);
and U6801 (N_6801,N_5670,N_4370);
nand U6802 (N_6802,N_5136,N_5415);
or U6803 (N_6803,N_5585,N_5637);
xor U6804 (N_6804,N_4787,N_4907);
and U6805 (N_6805,N_4554,N_4309);
xor U6806 (N_6806,N_5510,N_5936);
or U6807 (N_6807,N_4361,N_4856);
nor U6808 (N_6808,N_5049,N_4559);
xor U6809 (N_6809,N_4571,N_4989);
and U6810 (N_6810,N_5709,N_4851);
nand U6811 (N_6811,N_4935,N_5014);
xnor U6812 (N_6812,N_5193,N_5391);
and U6813 (N_6813,N_5269,N_5015);
and U6814 (N_6814,N_4155,N_5551);
xor U6815 (N_6815,N_4038,N_4416);
and U6816 (N_6816,N_4622,N_5889);
xor U6817 (N_6817,N_4529,N_5860);
nand U6818 (N_6818,N_4896,N_4563);
xor U6819 (N_6819,N_5991,N_4257);
and U6820 (N_6820,N_5262,N_4344);
nand U6821 (N_6821,N_4185,N_4005);
nand U6822 (N_6822,N_4227,N_5446);
nand U6823 (N_6823,N_4107,N_4768);
or U6824 (N_6824,N_4392,N_4800);
nand U6825 (N_6825,N_4612,N_4353);
or U6826 (N_6826,N_5256,N_5198);
nand U6827 (N_6827,N_4739,N_5957);
nor U6828 (N_6828,N_5903,N_5588);
and U6829 (N_6829,N_4321,N_4437);
and U6830 (N_6830,N_4261,N_5608);
and U6831 (N_6831,N_4840,N_5522);
nor U6832 (N_6832,N_5002,N_5431);
nand U6833 (N_6833,N_5814,N_4692);
nand U6834 (N_6834,N_4474,N_4661);
xnor U6835 (N_6835,N_5219,N_4095);
nor U6836 (N_6836,N_5211,N_5681);
and U6837 (N_6837,N_5071,N_5468);
and U6838 (N_6838,N_5753,N_5927);
nand U6839 (N_6839,N_4473,N_4932);
nand U6840 (N_6840,N_4944,N_5633);
or U6841 (N_6841,N_5651,N_4819);
nand U6842 (N_6842,N_5435,N_4575);
or U6843 (N_6843,N_4997,N_4239);
and U6844 (N_6844,N_5481,N_5826);
xnor U6845 (N_6845,N_4984,N_5855);
or U6846 (N_6846,N_4207,N_5527);
and U6847 (N_6847,N_4866,N_4876);
nor U6848 (N_6848,N_4725,N_4970);
nand U6849 (N_6849,N_5665,N_5266);
xnor U6850 (N_6850,N_5571,N_5881);
nor U6851 (N_6851,N_4662,N_4290);
nand U6852 (N_6852,N_4871,N_5876);
or U6853 (N_6853,N_5832,N_4518);
nand U6854 (N_6854,N_5465,N_5993);
nand U6855 (N_6855,N_5760,N_4111);
xnor U6856 (N_6856,N_4758,N_4356);
nor U6857 (N_6857,N_5661,N_4906);
nand U6858 (N_6858,N_5553,N_4966);
xor U6859 (N_6859,N_5549,N_5724);
nand U6860 (N_6860,N_4715,N_5225);
xor U6861 (N_6861,N_4103,N_4013);
nor U6862 (N_6862,N_4909,N_4582);
nor U6863 (N_6863,N_4953,N_4214);
nand U6864 (N_6864,N_4173,N_5255);
nor U6865 (N_6865,N_4194,N_5593);
or U6866 (N_6866,N_5396,N_4177);
nor U6867 (N_6867,N_5974,N_5190);
xor U6868 (N_6868,N_4125,N_4292);
and U6869 (N_6869,N_5422,N_4294);
or U6870 (N_6870,N_4680,N_4235);
xnor U6871 (N_6871,N_5321,N_5740);
or U6872 (N_6872,N_5965,N_4498);
and U6873 (N_6873,N_5587,N_5702);
xor U6874 (N_6874,N_4820,N_5909);
nand U6875 (N_6875,N_5756,N_5236);
nand U6876 (N_6876,N_5926,N_4486);
or U6877 (N_6877,N_4557,N_5246);
nand U6878 (N_6878,N_5616,N_5036);
nand U6879 (N_6879,N_4507,N_4767);
or U6880 (N_6880,N_4115,N_5358);
xor U6881 (N_6881,N_4070,N_4060);
and U6882 (N_6882,N_4343,N_5353);
nor U6883 (N_6883,N_4494,N_4743);
xor U6884 (N_6884,N_5241,N_5351);
and U6885 (N_6885,N_4511,N_5420);
nand U6886 (N_6886,N_4955,N_5444);
nor U6887 (N_6887,N_4730,N_5209);
or U6888 (N_6888,N_4042,N_4979);
xnor U6889 (N_6889,N_4147,N_5430);
and U6890 (N_6890,N_4810,N_4232);
and U6891 (N_6891,N_5804,N_5331);
and U6892 (N_6892,N_4415,N_5473);
nor U6893 (N_6893,N_4911,N_5580);
nor U6894 (N_6894,N_4887,N_5874);
and U6895 (N_6895,N_4246,N_5502);
nand U6896 (N_6896,N_4029,N_4106);
xnor U6897 (N_6897,N_4561,N_5810);
or U6898 (N_6898,N_4085,N_5650);
or U6899 (N_6899,N_4874,N_5199);
nand U6900 (N_6900,N_4846,N_4475);
nand U6901 (N_6901,N_5928,N_4007);
nor U6902 (N_6902,N_4382,N_4228);
nor U6903 (N_6903,N_5116,N_4645);
nor U6904 (N_6904,N_4056,N_4687);
nand U6905 (N_6905,N_4583,N_5409);
or U6906 (N_6906,N_5818,N_4285);
nor U6907 (N_6907,N_5945,N_4328);
and U6908 (N_6908,N_5497,N_5178);
nand U6909 (N_6909,N_4145,N_5742);
and U6910 (N_6910,N_5777,N_4117);
and U6911 (N_6911,N_5534,N_4606);
or U6912 (N_6912,N_4222,N_4525);
xor U6913 (N_6913,N_5170,N_4335);
or U6914 (N_6914,N_5306,N_5833);
xnor U6915 (N_6915,N_5374,N_5690);
or U6916 (N_6916,N_4455,N_5070);
nor U6917 (N_6917,N_5883,N_4766);
nor U6918 (N_6918,N_5602,N_5975);
or U6919 (N_6919,N_4675,N_5448);
nand U6920 (N_6920,N_5059,N_4531);
nor U6921 (N_6921,N_4171,N_4973);
nor U6922 (N_6922,N_4151,N_4395);
nor U6923 (N_6923,N_4289,N_4014);
nand U6924 (N_6924,N_5007,N_5954);
and U6925 (N_6925,N_5044,N_4065);
xnor U6926 (N_6926,N_5099,N_5825);
or U6927 (N_6927,N_4930,N_4927);
or U6928 (N_6928,N_5989,N_4124);
nor U6929 (N_6929,N_5504,N_4402);
xor U6930 (N_6930,N_4366,N_4238);
nand U6931 (N_6931,N_5687,N_5483);
and U6932 (N_6932,N_5066,N_5008);
nor U6933 (N_6933,N_5375,N_4262);
nor U6934 (N_6934,N_5186,N_5368);
nand U6935 (N_6935,N_4372,N_4254);
xnor U6936 (N_6936,N_4683,N_5733);
and U6937 (N_6937,N_5376,N_5399);
xor U6938 (N_6938,N_4438,N_5949);
nand U6939 (N_6939,N_5839,N_5110);
nand U6940 (N_6940,N_4360,N_5458);
nor U6941 (N_6941,N_5073,N_5134);
or U6942 (N_6942,N_4560,N_4853);
nor U6943 (N_6943,N_4780,N_5240);
xnor U6944 (N_6944,N_4980,N_4338);
nand U6945 (N_6945,N_5542,N_4461);
or U6946 (N_6946,N_5411,N_4676);
nand U6947 (N_6947,N_5297,N_4197);
and U6948 (N_6948,N_5119,N_5203);
xnor U6949 (N_6949,N_5565,N_5660);
or U6950 (N_6950,N_5506,N_4573);
or U6951 (N_6951,N_5152,N_4206);
or U6952 (N_6952,N_5560,N_4320);
xor U6953 (N_6953,N_5930,N_4672);
and U6954 (N_6954,N_5413,N_4957);
xnor U6955 (N_6955,N_4319,N_4986);
and U6956 (N_6956,N_4256,N_5054);
and U6957 (N_6957,N_4022,N_5967);
and U6958 (N_6958,N_4325,N_4389);
xor U6959 (N_6959,N_5366,N_5440);
nor U6960 (N_6960,N_4332,N_4477);
nor U6961 (N_6961,N_5300,N_4164);
and U6962 (N_6962,N_4318,N_4663);
or U6963 (N_6963,N_5323,N_5053);
nand U6964 (N_6964,N_4037,N_4528);
or U6965 (N_6965,N_5462,N_5125);
and U6966 (N_6966,N_5385,N_4330);
or U6967 (N_6967,N_5106,N_4677);
or U6968 (N_6968,N_4204,N_4084);
nor U6969 (N_6969,N_4546,N_5885);
nand U6970 (N_6970,N_5829,N_4597);
and U6971 (N_6971,N_5249,N_4555);
or U6972 (N_6972,N_4089,N_5999);
nor U6973 (N_6973,N_5596,N_4933);
xnor U6974 (N_6974,N_5747,N_4399);
and U6975 (N_6975,N_5018,N_4387);
xor U6976 (N_6976,N_5311,N_4696);
and U6977 (N_6977,N_4965,N_4919);
nand U6978 (N_6978,N_5794,N_5352);
nand U6979 (N_6979,N_5900,N_4358);
xnor U6980 (N_6980,N_5696,N_5405);
or U6981 (N_6981,N_5452,N_5032);
or U6982 (N_6982,N_4578,N_4418);
xor U6983 (N_6983,N_4718,N_4099);
xor U6984 (N_6984,N_4782,N_5227);
nand U6985 (N_6985,N_4745,N_4726);
nand U6986 (N_6986,N_4003,N_4634);
nand U6987 (N_6987,N_5728,N_4025);
and U6988 (N_6988,N_4537,N_5347);
nand U6989 (N_6989,N_4706,N_5813);
xnor U6990 (N_6990,N_5168,N_4414);
and U6991 (N_6991,N_5630,N_5570);
nand U6992 (N_6992,N_5085,N_5710);
xnor U6993 (N_6993,N_5274,N_5907);
or U6994 (N_6994,N_4329,N_5871);
nor U6995 (N_6995,N_5294,N_4439);
or U6996 (N_6996,N_5586,N_4071);
nor U6997 (N_6997,N_4032,N_4441);
nor U6998 (N_6998,N_5330,N_5478);
nor U6999 (N_6999,N_5815,N_5348);
or U7000 (N_7000,N_4345,N_4530);
xor U7001 (N_7001,N_5958,N_4356);
nor U7002 (N_7002,N_4553,N_5409);
or U7003 (N_7003,N_5973,N_5462);
and U7004 (N_7004,N_4043,N_5189);
or U7005 (N_7005,N_5685,N_4071);
xor U7006 (N_7006,N_5537,N_4444);
or U7007 (N_7007,N_4292,N_4967);
xor U7008 (N_7008,N_4963,N_4551);
nor U7009 (N_7009,N_4527,N_5643);
nor U7010 (N_7010,N_4123,N_4325);
and U7011 (N_7011,N_4157,N_4894);
or U7012 (N_7012,N_4903,N_4125);
nor U7013 (N_7013,N_4996,N_5842);
or U7014 (N_7014,N_5206,N_5068);
xnor U7015 (N_7015,N_5761,N_4890);
or U7016 (N_7016,N_4431,N_4052);
and U7017 (N_7017,N_4259,N_5452);
nand U7018 (N_7018,N_5643,N_4891);
xor U7019 (N_7019,N_5059,N_5124);
xor U7020 (N_7020,N_5901,N_5795);
xor U7021 (N_7021,N_4435,N_4457);
xor U7022 (N_7022,N_4839,N_4358);
nand U7023 (N_7023,N_4528,N_4330);
nor U7024 (N_7024,N_4102,N_4760);
and U7025 (N_7025,N_5959,N_4836);
nor U7026 (N_7026,N_5442,N_5947);
xor U7027 (N_7027,N_4852,N_4234);
xnor U7028 (N_7028,N_4039,N_4073);
nand U7029 (N_7029,N_4784,N_5463);
or U7030 (N_7030,N_4905,N_5190);
or U7031 (N_7031,N_4717,N_4231);
xnor U7032 (N_7032,N_4292,N_4968);
or U7033 (N_7033,N_4858,N_5158);
xnor U7034 (N_7034,N_4637,N_5544);
and U7035 (N_7035,N_4920,N_5286);
or U7036 (N_7036,N_5628,N_5968);
and U7037 (N_7037,N_4621,N_4457);
and U7038 (N_7038,N_5254,N_4250);
xor U7039 (N_7039,N_4743,N_5640);
and U7040 (N_7040,N_5299,N_4073);
nor U7041 (N_7041,N_4216,N_4129);
or U7042 (N_7042,N_4760,N_5825);
nand U7043 (N_7043,N_4216,N_4578);
nand U7044 (N_7044,N_4158,N_5526);
and U7045 (N_7045,N_5536,N_4522);
nand U7046 (N_7046,N_4060,N_5942);
and U7047 (N_7047,N_5660,N_5460);
xnor U7048 (N_7048,N_4413,N_4389);
nor U7049 (N_7049,N_5876,N_4410);
and U7050 (N_7050,N_4388,N_4747);
xor U7051 (N_7051,N_5610,N_5804);
nor U7052 (N_7052,N_5267,N_4577);
or U7053 (N_7053,N_5467,N_4323);
nor U7054 (N_7054,N_5733,N_4366);
and U7055 (N_7055,N_4918,N_4504);
nor U7056 (N_7056,N_5374,N_5229);
and U7057 (N_7057,N_5287,N_4657);
nand U7058 (N_7058,N_5702,N_4075);
or U7059 (N_7059,N_4586,N_5921);
xnor U7060 (N_7060,N_4454,N_5807);
xor U7061 (N_7061,N_5572,N_5406);
or U7062 (N_7062,N_4584,N_5433);
and U7063 (N_7063,N_5677,N_5368);
xor U7064 (N_7064,N_5966,N_4135);
nand U7065 (N_7065,N_5339,N_5861);
xnor U7066 (N_7066,N_5909,N_5818);
and U7067 (N_7067,N_5702,N_4335);
nor U7068 (N_7068,N_5134,N_4019);
or U7069 (N_7069,N_4228,N_4938);
nor U7070 (N_7070,N_4118,N_5780);
nand U7071 (N_7071,N_5747,N_4789);
or U7072 (N_7072,N_4071,N_5655);
or U7073 (N_7073,N_5072,N_4589);
xnor U7074 (N_7074,N_4115,N_4873);
and U7075 (N_7075,N_4416,N_5713);
and U7076 (N_7076,N_5161,N_4218);
or U7077 (N_7077,N_4965,N_5413);
nand U7078 (N_7078,N_5585,N_4652);
or U7079 (N_7079,N_4891,N_4371);
nand U7080 (N_7080,N_4784,N_5434);
or U7081 (N_7081,N_5489,N_5155);
and U7082 (N_7082,N_4778,N_5237);
nor U7083 (N_7083,N_4579,N_5944);
xnor U7084 (N_7084,N_4677,N_5868);
or U7085 (N_7085,N_5739,N_4426);
xor U7086 (N_7086,N_5750,N_4311);
or U7087 (N_7087,N_4587,N_4617);
and U7088 (N_7088,N_5178,N_5610);
nor U7089 (N_7089,N_4383,N_5601);
nand U7090 (N_7090,N_4259,N_4029);
xnor U7091 (N_7091,N_4086,N_4874);
xnor U7092 (N_7092,N_4749,N_4717);
and U7093 (N_7093,N_4328,N_5214);
nand U7094 (N_7094,N_5174,N_4258);
nand U7095 (N_7095,N_4927,N_5742);
nand U7096 (N_7096,N_4877,N_4587);
nor U7097 (N_7097,N_4583,N_5969);
nor U7098 (N_7098,N_5230,N_5849);
nor U7099 (N_7099,N_5281,N_4517);
nor U7100 (N_7100,N_4024,N_4941);
or U7101 (N_7101,N_5042,N_5585);
and U7102 (N_7102,N_4306,N_5208);
and U7103 (N_7103,N_5427,N_5181);
nor U7104 (N_7104,N_5616,N_5129);
or U7105 (N_7105,N_5785,N_4672);
nand U7106 (N_7106,N_4166,N_5135);
or U7107 (N_7107,N_4447,N_5938);
nand U7108 (N_7108,N_5849,N_4815);
nand U7109 (N_7109,N_5160,N_5548);
and U7110 (N_7110,N_4775,N_5239);
nor U7111 (N_7111,N_4804,N_5690);
and U7112 (N_7112,N_5458,N_4910);
nor U7113 (N_7113,N_4297,N_5681);
and U7114 (N_7114,N_4910,N_5059);
nand U7115 (N_7115,N_4325,N_5394);
nor U7116 (N_7116,N_4473,N_4891);
nor U7117 (N_7117,N_4008,N_5183);
nor U7118 (N_7118,N_5990,N_5475);
xor U7119 (N_7119,N_5110,N_5545);
or U7120 (N_7120,N_5869,N_5817);
xor U7121 (N_7121,N_5749,N_5529);
xnor U7122 (N_7122,N_4911,N_4966);
or U7123 (N_7123,N_4004,N_5967);
xor U7124 (N_7124,N_5811,N_4342);
nor U7125 (N_7125,N_5938,N_5162);
or U7126 (N_7126,N_4765,N_5680);
nor U7127 (N_7127,N_4808,N_5661);
and U7128 (N_7128,N_5845,N_5630);
nor U7129 (N_7129,N_4837,N_5011);
nand U7130 (N_7130,N_4136,N_5907);
xnor U7131 (N_7131,N_4431,N_5719);
or U7132 (N_7132,N_4294,N_4935);
and U7133 (N_7133,N_5684,N_4198);
xor U7134 (N_7134,N_4587,N_4538);
and U7135 (N_7135,N_5972,N_4192);
xor U7136 (N_7136,N_4739,N_4896);
and U7137 (N_7137,N_4719,N_5910);
and U7138 (N_7138,N_5636,N_5429);
nor U7139 (N_7139,N_5924,N_4890);
nor U7140 (N_7140,N_4636,N_4614);
nand U7141 (N_7141,N_4730,N_5140);
and U7142 (N_7142,N_5825,N_4828);
nor U7143 (N_7143,N_4759,N_5260);
nor U7144 (N_7144,N_5781,N_4466);
and U7145 (N_7145,N_4993,N_4028);
nand U7146 (N_7146,N_4579,N_4505);
or U7147 (N_7147,N_5406,N_4208);
xor U7148 (N_7148,N_5674,N_4992);
xor U7149 (N_7149,N_4059,N_4841);
and U7150 (N_7150,N_5760,N_4253);
and U7151 (N_7151,N_5211,N_5464);
or U7152 (N_7152,N_4804,N_5755);
xor U7153 (N_7153,N_5651,N_5711);
and U7154 (N_7154,N_5111,N_5131);
and U7155 (N_7155,N_4590,N_5115);
nor U7156 (N_7156,N_4535,N_4079);
xnor U7157 (N_7157,N_5821,N_5942);
xnor U7158 (N_7158,N_5448,N_4329);
nand U7159 (N_7159,N_4548,N_5812);
nand U7160 (N_7160,N_5355,N_5110);
or U7161 (N_7161,N_4859,N_5850);
nor U7162 (N_7162,N_4421,N_5820);
or U7163 (N_7163,N_4669,N_4056);
xnor U7164 (N_7164,N_5872,N_5154);
nand U7165 (N_7165,N_4032,N_5806);
nand U7166 (N_7166,N_4988,N_4251);
and U7167 (N_7167,N_4590,N_4948);
nor U7168 (N_7168,N_4369,N_4375);
xnor U7169 (N_7169,N_5271,N_5646);
nand U7170 (N_7170,N_5949,N_5284);
xor U7171 (N_7171,N_4799,N_5349);
or U7172 (N_7172,N_5994,N_5649);
nor U7173 (N_7173,N_4280,N_5909);
and U7174 (N_7174,N_4113,N_5578);
or U7175 (N_7175,N_4927,N_4925);
and U7176 (N_7176,N_4364,N_5450);
and U7177 (N_7177,N_5019,N_5926);
and U7178 (N_7178,N_5160,N_5724);
nand U7179 (N_7179,N_4378,N_5179);
and U7180 (N_7180,N_4049,N_4982);
nor U7181 (N_7181,N_5216,N_4373);
nand U7182 (N_7182,N_4485,N_5265);
or U7183 (N_7183,N_4112,N_5520);
nor U7184 (N_7184,N_5110,N_4639);
nand U7185 (N_7185,N_4849,N_4223);
or U7186 (N_7186,N_4504,N_4299);
nor U7187 (N_7187,N_5472,N_4544);
nor U7188 (N_7188,N_5741,N_4270);
and U7189 (N_7189,N_5407,N_4340);
xnor U7190 (N_7190,N_4281,N_5098);
nand U7191 (N_7191,N_5048,N_5141);
nor U7192 (N_7192,N_5358,N_4736);
and U7193 (N_7193,N_4721,N_4795);
xor U7194 (N_7194,N_4892,N_5898);
and U7195 (N_7195,N_5184,N_4310);
or U7196 (N_7196,N_5949,N_5982);
nand U7197 (N_7197,N_5364,N_5218);
or U7198 (N_7198,N_4843,N_4726);
nand U7199 (N_7199,N_4595,N_4451);
and U7200 (N_7200,N_5800,N_5251);
nand U7201 (N_7201,N_5757,N_4167);
and U7202 (N_7202,N_4355,N_4133);
nand U7203 (N_7203,N_4295,N_5472);
xnor U7204 (N_7204,N_5405,N_5207);
xnor U7205 (N_7205,N_4586,N_4748);
or U7206 (N_7206,N_4493,N_5994);
or U7207 (N_7207,N_5604,N_4061);
and U7208 (N_7208,N_4383,N_5503);
xor U7209 (N_7209,N_5330,N_5868);
xor U7210 (N_7210,N_4314,N_5614);
nand U7211 (N_7211,N_5909,N_4475);
and U7212 (N_7212,N_4434,N_5896);
or U7213 (N_7213,N_4701,N_4593);
nor U7214 (N_7214,N_5145,N_5602);
or U7215 (N_7215,N_4599,N_5805);
xor U7216 (N_7216,N_5937,N_5177);
nor U7217 (N_7217,N_5855,N_5798);
nand U7218 (N_7218,N_4965,N_5903);
nand U7219 (N_7219,N_5007,N_4192);
nor U7220 (N_7220,N_5815,N_5729);
or U7221 (N_7221,N_5284,N_5324);
and U7222 (N_7222,N_4561,N_5805);
nand U7223 (N_7223,N_5592,N_5765);
and U7224 (N_7224,N_4134,N_5186);
nand U7225 (N_7225,N_4288,N_5907);
nand U7226 (N_7226,N_4956,N_5267);
nor U7227 (N_7227,N_4703,N_5905);
and U7228 (N_7228,N_5016,N_5898);
nor U7229 (N_7229,N_4855,N_5730);
or U7230 (N_7230,N_4276,N_5181);
nand U7231 (N_7231,N_4619,N_5805);
or U7232 (N_7232,N_5651,N_4186);
nand U7233 (N_7233,N_4667,N_5210);
nand U7234 (N_7234,N_4426,N_4049);
and U7235 (N_7235,N_4498,N_4990);
nor U7236 (N_7236,N_5987,N_4509);
xnor U7237 (N_7237,N_5947,N_5096);
xnor U7238 (N_7238,N_4677,N_4476);
xor U7239 (N_7239,N_5564,N_5361);
xor U7240 (N_7240,N_4762,N_5795);
nor U7241 (N_7241,N_5868,N_4283);
nand U7242 (N_7242,N_4286,N_4826);
xor U7243 (N_7243,N_5832,N_4691);
nor U7244 (N_7244,N_4075,N_4311);
xnor U7245 (N_7245,N_4361,N_5694);
nand U7246 (N_7246,N_4110,N_5581);
and U7247 (N_7247,N_4675,N_4639);
and U7248 (N_7248,N_5460,N_5045);
xor U7249 (N_7249,N_5300,N_4099);
nand U7250 (N_7250,N_4615,N_4106);
or U7251 (N_7251,N_5216,N_5002);
and U7252 (N_7252,N_4026,N_4261);
and U7253 (N_7253,N_4055,N_4135);
nor U7254 (N_7254,N_4306,N_4061);
or U7255 (N_7255,N_4059,N_5681);
or U7256 (N_7256,N_5565,N_4174);
or U7257 (N_7257,N_5629,N_4100);
nand U7258 (N_7258,N_5221,N_4081);
or U7259 (N_7259,N_4552,N_5236);
xnor U7260 (N_7260,N_5978,N_4828);
xor U7261 (N_7261,N_5084,N_5075);
and U7262 (N_7262,N_4373,N_4919);
xor U7263 (N_7263,N_5173,N_4054);
nand U7264 (N_7264,N_4422,N_5601);
nand U7265 (N_7265,N_4537,N_5521);
xor U7266 (N_7266,N_4777,N_5864);
nor U7267 (N_7267,N_4061,N_4101);
and U7268 (N_7268,N_4092,N_5446);
nand U7269 (N_7269,N_5063,N_5188);
xor U7270 (N_7270,N_4871,N_5108);
nor U7271 (N_7271,N_4400,N_5747);
and U7272 (N_7272,N_5224,N_5325);
or U7273 (N_7273,N_4413,N_5031);
or U7274 (N_7274,N_4261,N_5372);
xnor U7275 (N_7275,N_5308,N_4084);
and U7276 (N_7276,N_5752,N_5440);
nand U7277 (N_7277,N_5066,N_5675);
nand U7278 (N_7278,N_5492,N_5286);
or U7279 (N_7279,N_5287,N_4545);
and U7280 (N_7280,N_5462,N_4279);
nand U7281 (N_7281,N_4100,N_4192);
and U7282 (N_7282,N_4772,N_4340);
nand U7283 (N_7283,N_5677,N_4579);
nand U7284 (N_7284,N_5917,N_5994);
nor U7285 (N_7285,N_5031,N_5897);
and U7286 (N_7286,N_5828,N_4134);
or U7287 (N_7287,N_4157,N_5451);
or U7288 (N_7288,N_4152,N_4183);
nor U7289 (N_7289,N_4896,N_5195);
nor U7290 (N_7290,N_5736,N_5615);
nor U7291 (N_7291,N_5957,N_4484);
nand U7292 (N_7292,N_4260,N_5343);
nand U7293 (N_7293,N_4817,N_5072);
nor U7294 (N_7294,N_4158,N_4331);
and U7295 (N_7295,N_4067,N_4567);
and U7296 (N_7296,N_5232,N_5235);
nor U7297 (N_7297,N_5519,N_5344);
nor U7298 (N_7298,N_5494,N_5711);
nor U7299 (N_7299,N_5027,N_5952);
nor U7300 (N_7300,N_5170,N_5656);
nor U7301 (N_7301,N_5001,N_4347);
and U7302 (N_7302,N_4518,N_4344);
nor U7303 (N_7303,N_4610,N_5170);
nor U7304 (N_7304,N_5003,N_4573);
and U7305 (N_7305,N_5094,N_5963);
or U7306 (N_7306,N_5783,N_4022);
xor U7307 (N_7307,N_4404,N_5036);
xnor U7308 (N_7308,N_5775,N_5760);
xor U7309 (N_7309,N_4862,N_4349);
and U7310 (N_7310,N_4143,N_4938);
xor U7311 (N_7311,N_5073,N_5747);
xnor U7312 (N_7312,N_5655,N_5522);
and U7313 (N_7313,N_5023,N_4654);
nor U7314 (N_7314,N_5164,N_5968);
nor U7315 (N_7315,N_5387,N_4456);
nand U7316 (N_7316,N_4909,N_5710);
and U7317 (N_7317,N_4742,N_4971);
nor U7318 (N_7318,N_5545,N_4122);
xnor U7319 (N_7319,N_4675,N_4257);
xnor U7320 (N_7320,N_5684,N_4211);
or U7321 (N_7321,N_5230,N_4906);
nor U7322 (N_7322,N_4507,N_4229);
nand U7323 (N_7323,N_5084,N_5363);
xnor U7324 (N_7324,N_5552,N_4156);
nand U7325 (N_7325,N_5059,N_4866);
or U7326 (N_7326,N_5820,N_5102);
nand U7327 (N_7327,N_5735,N_4460);
or U7328 (N_7328,N_5567,N_5732);
nand U7329 (N_7329,N_4940,N_4192);
nor U7330 (N_7330,N_5913,N_4931);
or U7331 (N_7331,N_5023,N_5733);
or U7332 (N_7332,N_4508,N_5857);
nor U7333 (N_7333,N_4559,N_4289);
or U7334 (N_7334,N_5472,N_4400);
xnor U7335 (N_7335,N_4071,N_5423);
and U7336 (N_7336,N_4255,N_4333);
nor U7337 (N_7337,N_5504,N_5849);
nor U7338 (N_7338,N_5125,N_5080);
and U7339 (N_7339,N_4309,N_4324);
nand U7340 (N_7340,N_4513,N_5867);
or U7341 (N_7341,N_4826,N_5826);
nand U7342 (N_7342,N_4740,N_4483);
and U7343 (N_7343,N_5333,N_5794);
nand U7344 (N_7344,N_4010,N_5590);
nand U7345 (N_7345,N_4768,N_4767);
or U7346 (N_7346,N_4357,N_4686);
xnor U7347 (N_7347,N_4290,N_5337);
or U7348 (N_7348,N_5404,N_4627);
or U7349 (N_7349,N_4273,N_4110);
xor U7350 (N_7350,N_4928,N_4262);
or U7351 (N_7351,N_5135,N_4367);
nor U7352 (N_7352,N_4046,N_4415);
nand U7353 (N_7353,N_4711,N_5193);
nor U7354 (N_7354,N_4748,N_5182);
nor U7355 (N_7355,N_5574,N_4008);
or U7356 (N_7356,N_4826,N_4994);
and U7357 (N_7357,N_4946,N_4556);
nand U7358 (N_7358,N_4451,N_4412);
nand U7359 (N_7359,N_5503,N_4942);
nand U7360 (N_7360,N_4304,N_5827);
and U7361 (N_7361,N_4608,N_5402);
or U7362 (N_7362,N_5593,N_5389);
xor U7363 (N_7363,N_5694,N_5201);
or U7364 (N_7364,N_5469,N_4610);
nor U7365 (N_7365,N_4968,N_4000);
nor U7366 (N_7366,N_5656,N_5380);
xnor U7367 (N_7367,N_4386,N_5713);
xor U7368 (N_7368,N_4372,N_5231);
nor U7369 (N_7369,N_4397,N_5391);
nand U7370 (N_7370,N_4511,N_4829);
nand U7371 (N_7371,N_5534,N_5139);
and U7372 (N_7372,N_4273,N_5715);
nor U7373 (N_7373,N_5158,N_4495);
or U7374 (N_7374,N_5161,N_5377);
xnor U7375 (N_7375,N_5333,N_4286);
and U7376 (N_7376,N_4435,N_5952);
xor U7377 (N_7377,N_4202,N_5720);
or U7378 (N_7378,N_5642,N_4039);
and U7379 (N_7379,N_4659,N_4699);
xnor U7380 (N_7380,N_5797,N_5078);
or U7381 (N_7381,N_5472,N_5463);
nand U7382 (N_7382,N_5172,N_4039);
and U7383 (N_7383,N_4425,N_5676);
nor U7384 (N_7384,N_5914,N_4038);
and U7385 (N_7385,N_4603,N_4783);
nand U7386 (N_7386,N_4078,N_4759);
xnor U7387 (N_7387,N_5070,N_4528);
and U7388 (N_7388,N_5741,N_5396);
xnor U7389 (N_7389,N_5191,N_5709);
nor U7390 (N_7390,N_4991,N_4196);
xor U7391 (N_7391,N_4981,N_5658);
xor U7392 (N_7392,N_4148,N_5859);
or U7393 (N_7393,N_5385,N_5529);
nor U7394 (N_7394,N_5852,N_5879);
xor U7395 (N_7395,N_5643,N_4850);
xor U7396 (N_7396,N_4692,N_4755);
nor U7397 (N_7397,N_5013,N_4603);
nand U7398 (N_7398,N_5477,N_5711);
nor U7399 (N_7399,N_5241,N_5305);
xor U7400 (N_7400,N_4070,N_4601);
nand U7401 (N_7401,N_5402,N_4004);
nand U7402 (N_7402,N_5747,N_5270);
nor U7403 (N_7403,N_4698,N_4344);
xnor U7404 (N_7404,N_5710,N_4942);
nand U7405 (N_7405,N_4157,N_4882);
or U7406 (N_7406,N_4614,N_5412);
xor U7407 (N_7407,N_5695,N_4676);
or U7408 (N_7408,N_5165,N_5132);
xor U7409 (N_7409,N_5625,N_5695);
and U7410 (N_7410,N_4290,N_4311);
and U7411 (N_7411,N_4525,N_4710);
or U7412 (N_7412,N_4431,N_4734);
xor U7413 (N_7413,N_5911,N_5617);
or U7414 (N_7414,N_5259,N_5283);
or U7415 (N_7415,N_5368,N_4660);
or U7416 (N_7416,N_5334,N_4969);
nor U7417 (N_7417,N_4418,N_5662);
xnor U7418 (N_7418,N_5282,N_5332);
or U7419 (N_7419,N_5640,N_5664);
xor U7420 (N_7420,N_5423,N_4121);
and U7421 (N_7421,N_5834,N_4738);
nor U7422 (N_7422,N_5181,N_4820);
xor U7423 (N_7423,N_5788,N_4002);
and U7424 (N_7424,N_5214,N_4158);
nor U7425 (N_7425,N_4764,N_4869);
and U7426 (N_7426,N_4435,N_5427);
and U7427 (N_7427,N_4140,N_4544);
xor U7428 (N_7428,N_5137,N_4794);
or U7429 (N_7429,N_5853,N_4021);
nand U7430 (N_7430,N_5690,N_4394);
nand U7431 (N_7431,N_5764,N_4208);
xor U7432 (N_7432,N_5806,N_5039);
nand U7433 (N_7433,N_4365,N_5253);
and U7434 (N_7434,N_5473,N_4731);
nor U7435 (N_7435,N_4493,N_4293);
or U7436 (N_7436,N_4570,N_4102);
xor U7437 (N_7437,N_5350,N_5988);
nor U7438 (N_7438,N_5302,N_5437);
and U7439 (N_7439,N_5797,N_4501);
and U7440 (N_7440,N_5548,N_5376);
or U7441 (N_7441,N_4150,N_4676);
nor U7442 (N_7442,N_4906,N_5232);
xor U7443 (N_7443,N_4220,N_5311);
nor U7444 (N_7444,N_5455,N_4682);
xor U7445 (N_7445,N_4076,N_4324);
or U7446 (N_7446,N_4447,N_4642);
or U7447 (N_7447,N_4775,N_5102);
nor U7448 (N_7448,N_4935,N_4564);
and U7449 (N_7449,N_5670,N_5060);
or U7450 (N_7450,N_5653,N_4163);
nand U7451 (N_7451,N_4183,N_4597);
or U7452 (N_7452,N_5534,N_5142);
nor U7453 (N_7453,N_5177,N_4769);
nand U7454 (N_7454,N_5380,N_4124);
nand U7455 (N_7455,N_5686,N_5367);
xor U7456 (N_7456,N_5561,N_5474);
nor U7457 (N_7457,N_5689,N_5821);
nand U7458 (N_7458,N_5104,N_5009);
nand U7459 (N_7459,N_4397,N_4317);
nand U7460 (N_7460,N_5856,N_5826);
nand U7461 (N_7461,N_5469,N_5623);
and U7462 (N_7462,N_5353,N_5042);
xor U7463 (N_7463,N_4334,N_5799);
or U7464 (N_7464,N_5413,N_4180);
and U7465 (N_7465,N_4014,N_5688);
xnor U7466 (N_7466,N_5125,N_4933);
nor U7467 (N_7467,N_4049,N_5784);
xor U7468 (N_7468,N_5650,N_4503);
nor U7469 (N_7469,N_5944,N_4606);
xnor U7470 (N_7470,N_4576,N_4787);
and U7471 (N_7471,N_5721,N_5122);
nand U7472 (N_7472,N_5213,N_4417);
nand U7473 (N_7473,N_5424,N_4639);
xor U7474 (N_7474,N_4492,N_4298);
and U7475 (N_7475,N_4074,N_4693);
xor U7476 (N_7476,N_4797,N_4287);
nor U7477 (N_7477,N_5573,N_5244);
or U7478 (N_7478,N_5800,N_5822);
nand U7479 (N_7479,N_4687,N_4084);
nand U7480 (N_7480,N_4381,N_5680);
nand U7481 (N_7481,N_4550,N_5998);
and U7482 (N_7482,N_5299,N_4455);
and U7483 (N_7483,N_5864,N_4921);
xnor U7484 (N_7484,N_5884,N_4530);
nand U7485 (N_7485,N_4830,N_5318);
xnor U7486 (N_7486,N_4942,N_5029);
and U7487 (N_7487,N_4098,N_5493);
and U7488 (N_7488,N_4183,N_5134);
xnor U7489 (N_7489,N_4337,N_4828);
nor U7490 (N_7490,N_5471,N_5444);
nand U7491 (N_7491,N_5466,N_5780);
or U7492 (N_7492,N_4356,N_4728);
nor U7493 (N_7493,N_4890,N_5220);
and U7494 (N_7494,N_5318,N_5732);
nor U7495 (N_7495,N_5911,N_5189);
xnor U7496 (N_7496,N_4159,N_4652);
and U7497 (N_7497,N_5990,N_4692);
nand U7498 (N_7498,N_4562,N_5555);
and U7499 (N_7499,N_4773,N_4020);
and U7500 (N_7500,N_4028,N_4046);
nand U7501 (N_7501,N_4985,N_5263);
xor U7502 (N_7502,N_4477,N_4089);
nand U7503 (N_7503,N_5692,N_5493);
nand U7504 (N_7504,N_5309,N_4098);
nand U7505 (N_7505,N_5907,N_4532);
xor U7506 (N_7506,N_4520,N_4860);
or U7507 (N_7507,N_4622,N_4804);
nand U7508 (N_7508,N_5494,N_5792);
and U7509 (N_7509,N_5558,N_5857);
nor U7510 (N_7510,N_4256,N_4550);
xor U7511 (N_7511,N_5126,N_4176);
xnor U7512 (N_7512,N_4097,N_5233);
xnor U7513 (N_7513,N_5463,N_5153);
or U7514 (N_7514,N_4136,N_4527);
nor U7515 (N_7515,N_5120,N_4612);
and U7516 (N_7516,N_5911,N_4279);
nor U7517 (N_7517,N_5539,N_5216);
or U7518 (N_7518,N_4800,N_4007);
xnor U7519 (N_7519,N_5597,N_4715);
nand U7520 (N_7520,N_4530,N_4650);
nand U7521 (N_7521,N_4168,N_4104);
xnor U7522 (N_7522,N_5733,N_4994);
nor U7523 (N_7523,N_5362,N_4699);
nor U7524 (N_7524,N_5074,N_4362);
or U7525 (N_7525,N_4023,N_4144);
and U7526 (N_7526,N_5009,N_5786);
and U7527 (N_7527,N_5468,N_5252);
and U7528 (N_7528,N_4806,N_4613);
and U7529 (N_7529,N_5182,N_5071);
and U7530 (N_7530,N_5804,N_4750);
xnor U7531 (N_7531,N_4787,N_5753);
or U7532 (N_7532,N_4290,N_5002);
or U7533 (N_7533,N_4256,N_4919);
nand U7534 (N_7534,N_4014,N_4570);
or U7535 (N_7535,N_5827,N_5924);
or U7536 (N_7536,N_5852,N_4727);
nor U7537 (N_7537,N_5430,N_5250);
nand U7538 (N_7538,N_4196,N_5310);
nand U7539 (N_7539,N_4068,N_5097);
nor U7540 (N_7540,N_4228,N_5912);
and U7541 (N_7541,N_4614,N_5081);
xnor U7542 (N_7542,N_4482,N_5651);
nand U7543 (N_7543,N_4629,N_5664);
nor U7544 (N_7544,N_5101,N_5796);
nand U7545 (N_7545,N_5933,N_4462);
xnor U7546 (N_7546,N_4123,N_5523);
nand U7547 (N_7547,N_4447,N_4448);
nor U7548 (N_7548,N_5128,N_4545);
nor U7549 (N_7549,N_4342,N_5860);
xor U7550 (N_7550,N_4196,N_4553);
nand U7551 (N_7551,N_4410,N_4814);
nor U7552 (N_7552,N_4502,N_4938);
xnor U7553 (N_7553,N_5514,N_4169);
or U7554 (N_7554,N_5493,N_5615);
xor U7555 (N_7555,N_4734,N_5902);
and U7556 (N_7556,N_4857,N_5680);
xnor U7557 (N_7557,N_4853,N_4146);
nor U7558 (N_7558,N_4696,N_4590);
nor U7559 (N_7559,N_5917,N_4723);
nand U7560 (N_7560,N_4301,N_4572);
nand U7561 (N_7561,N_5138,N_4315);
xor U7562 (N_7562,N_4873,N_4323);
xnor U7563 (N_7563,N_4930,N_5276);
and U7564 (N_7564,N_5682,N_4683);
xnor U7565 (N_7565,N_5462,N_4868);
and U7566 (N_7566,N_5535,N_4454);
nor U7567 (N_7567,N_4823,N_5291);
and U7568 (N_7568,N_5661,N_4284);
nor U7569 (N_7569,N_4929,N_5091);
nor U7570 (N_7570,N_5342,N_4962);
or U7571 (N_7571,N_4894,N_4408);
xnor U7572 (N_7572,N_5457,N_5580);
and U7573 (N_7573,N_5234,N_4478);
nand U7574 (N_7574,N_4593,N_5198);
and U7575 (N_7575,N_4987,N_4766);
nor U7576 (N_7576,N_5748,N_4050);
xor U7577 (N_7577,N_5838,N_5894);
nand U7578 (N_7578,N_5759,N_5326);
nor U7579 (N_7579,N_4639,N_5360);
xor U7580 (N_7580,N_5762,N_5362);
nor U7581 (N_7581,N_4810,N_4672);
or U7582 (N_7582,N_4263,N_5858);
or U7583 (N_7583,N_4263,N_4861);
nand U7584 (N_7584,N_5100,N_5904);
nor U7585 (N_7585,N_4624,N_4603);
xnor U7586 (N_7586,N_5104,N_5719);
xor U7587 (N_7587,N_4037,N_4029);
and U7588 (N_7588,N_5430,N_5899);
xor U7589 (N_7589,N_4121,N_5090);
xnor U7590 (N_7590,N_4924,N_5471);
nand U7591 (N_7591,N_5216,N_5076);
nor U7592 (N_7592,N_5851,N_5468);
nand U7593 (N_7593,N_5093,N_4189);
xor U7594 (N_7594,N_5599,N_5277);
nand U7595 (N_7595,N_4262,N_5117);
xnor U7596 (N_7596,N_5973,N_4836);
and U7597 (N_7597,N_4365,N_4110);
xor U7598 (N_7598,N_5899,N_4055);
or U7599 (N_7599,N_5184,N_4445);
xor U7600 (N_7600,N_4141,N_4851);
nand U7601 (N_7601,N_5412,N_4858);
nor U7602 (N_7602,N_4473,N_5832);
nor U7603 (N_7603,N_5645,N_5189);
nand U7604 (N_7604,N_4905,N_5690);
and U7605 (N_7605,N_5114,N_5560);
nand U7606 (N_7606,N_4478,N_5729);
or U7607 (N_7607,N_4907,N_4837);
or U7608 (N_7608,N_5997,N_5032);
and U7609 (N_7609,N_5686,N_5775);
xor U7610 (N_7610,N_4867,N_5442);
xnor U7611 (N_7611,N_4760,N_5700);
nor U7612 (N_7612,N_5974,N_5721);
nand U7613 (N_7613,N_5197,N_4029);
or U7614 (N_7614,N_4979,N_4085);
or U7615 (N_7615,N_5367,N_5724);
or U7616 (N_7616,N_5123,N_5097);
nand U7617 (N_7617,N_5575,N_4715);
xor U7618 (N_7618,N_5596,N_4015);
or U7619 (N_7619,N_5469,N_4202);
nand U7620 (N_7620,N_4294,N_4707);
or U7621 (N_7621,N_5393,N_5122);
xnor U7622 (N_7622,N_4322,N_4346);
xnor U7623 (N_7623,N_5634,N_5998);
and U7624 (N_7624,N_4263,N_4026);
or U7625 (N_7625,N_5442,N_4679);
and U7626 (N_7626,N_4631,N_5362);
nor U7627 (N_7627,N_4856,N_5817);
or U7628 (N_7628,N_4088,N_5258);
nor U7629 (N_7629,N_5149,N_4146);
xor U7630 (N_7630,N_5216,N_4871);
nand U7631 (N_7631,N_4798,N_4874);
xor U7632 (N_7632,N_4172,N_4845);
and U7633 (N_7633,N_4011,N_5108);
xor U7634 (N_7634,N_5712,N_4922);
nand U7635 (N_7635,N_5746,N_4170);
xnor U7636 (N_7636,N_4657,N_5570);
and U7637 (N_7637,N_4601,N_4981);
or U7638 (N_7638,N_5721,N_5737);
nor U7639 (N_7639,N_5330,N_5608);
or U7640 (N_7640,N_5700,N_4604);
or U7641 (N_7641,N_4006,N_5035);
nor U7642 (N_7642,N_5868,N_4332);
xnor U7643 (N_7643,N_5428,N_5712);
nand U7644 (N_7644,N_5522,N_4309);
or U7645 (N_7645,N_4817,N_5307);
nand U7646 (N_7646,N_5232,N_4128);
nor U7647 (N_7647,N_5958,N_5713);
xnor U7648 (N_7648,N_4308,N_5566);
nand U7649 (N_7649,N_5122,N_4360);
or U7650 (N_7650,N_5618,N_5797);
nand U7651 (N_7651,N_5214,N_4761);
nor U7652 (N_7652,N_4137,N_5551);
nand U7653 (N_7653,N_5998,N_5864);
and U7654 (N_7654,N_4784,N_4030);
xor U7655 (N_7655,N_5753,N_5161);
or U7656 (N_7656,N_4431,N_5281);
xor U7657 (N_7657,N_5524,N_4868);
and U7658 (N_7658,N_5465,N_4127);
and U7659 (N_7659,N_5947,N_4508);
nor U7660 (N_7660,N_5315,N_5084);
nand U7661 (N_7661,N_5307,N_5211);
or U7662 (N_7662,N_5451,N_4362);
nor U7663 (N_7663,N_4656,N_5060);
and U7664 (N_7664,N_4133,N_5113);
nand U7665 (N_7665,N_4369,N_5504);
or U7666 (N_7666,N_5633,N_4292);
and U7667 (N_7667,N_4932,N_4053);
nor U7668 (N_7668,N_4933,N_4052);
xor U7669 (N_7669,N_4498,N_5730);
or U7670 (N_7670,N_5362,N_5924);
xnor U7671 (N_7671,N_5427,N_4769);
nor U7672 (N_7672,N_5077,N_5013);
or U7673 (N_7673,N_5935,N_5327);
xor U7674 (N_7674,N_5983,N_4752);
xnor U7675 (N_7675,N_4513,N_4445);
or U7676 (N_7676,N_5494,N_5542);
and U7677 (N_7677,N_5202,N_5772);
xnor U7678 (N_7678,N_4612,N_4855);
or U7679 (N_7679,N_4162,N_4540);
nand U7680 (N_7680,N_4488,N_4357);
xnor U7681 (N_7681,N_4656,N_4218);
nor U7682 (N_7682,N_5845,N_5596);
or U7683 (N_7683,N_5484,N_5332);
and U7684 (N_7684,N_4779,N_5946);
nand U7685 (N_7685,N_5345,N_5803);
nor U7686 (N_7686,N_4315,N_5381);
nor U7687 (N_7687,N_5282,N_4386);
nor U7688 (N_7688,N_4500,N_5698);
and U7689 (N_7689,N_4252,N_5257);
or U7690 (N_7690,N_5225,N_5502);
and U7691 (N_7691,N_5898,N_5727);
nand U7692 (N_7692,N_5030,N_5082);
nand U7693 (N_7693,N_4724,N_4217);
or U7694 (N_7694,N_5323,N_4802);
and U7695 (N_7695,N_5931,N_4183);
xnor U7696 (N_7696,N_4487,N_5288);
nand U7697 (N_7697,N_5953,N_5459);
or U7698 (N_7698,N_5354,N_4150);
or U7699 (N_7699,N_4806,N_5257);
nand U7700 (N_7700,N_5259,N_4612);
or U7701 (N_7701,N_4627,N_5594);
nand U7702 (N_7702,N_5464,N_4677);
or U7703 (N_7703,N_5159,N_4478);
nand U7704 (N_7704,N_5544,N_5384);
and U7705 (N_7705,N_5742,N_4182);
or U7706 (N_7706,N_4981,N_5006);
xnor U7707 (N_7707,N_5800,N_5680);
nor U7708 (N_7708,N_4823,N_5323);
nand U7709 (N_7709,N_4998,N_4464);
nor U7710 (N_7710,N_4221,N_4216);
xnor U7711 (N_7711,N_5198,N_4932);
and U7712 (N_7712,N_4561,N_5815);
nor U7713 (N_7713,N_4593,N_4887);
and U7714 (N_7714,N_5864,N_5231);
or U7715 (N_7715,N_5589,N_5428);
nand U7716 (N_7716,N_5049,N_5105);
nor U7717 (N_7717,N_4159,N_5285);
xnor U7718 (N_7718,N_5978,N_5736);
xor U7719 (N_7719,N_5189,N_4896);
or U7720 (N_7720,N_4149,N_4023);
or U7721 (N_7721,N_4594,N_4009);
and U7722 (N_7722,N_5301,N_5067);
xnor U7723 (N_7723,N_5215,N_5139);
nand U7724 (N_7724,N_4837,N_5007);
or U7725 (N_7725,N_5814,N_4527);
nor U7726 (N_7726,N_4615,N_4748);
and U7727 (N_7727,N_4973,N_5170);
or U7728 (N_7728,N_4170,N_4064);
xnor U7729 (N_7729,N_5254,N_4105);
xnor U7730 (N_7730,N_5736,N_4082);
or U7731 (N_7731,N_5069,N_5013);
and U7732 (N_7732,N_5669,N_4335);
or U7733 (N_7733,N_5135,N_4583);
and U7734 (N_7734,N_4693,N_5004);
xnor U7735 (N_7735,N_4493,N_5884);
or U7736 (N_7736,N_4168,N_5050);
or U7737 (N_7737,N_5576,N_5712);
or U7738 (N_7738,N_5127,N_4597);
xor U7739 (N_7739,N_4889,N_4947);
nand U7740 (N_7740,N_4418,N_4498);
or U7741 (N_7741,N_4263,N_5921);
or U7742 (N_7742,N_4562,N_4825);
and U7743 (N_7743,N_4369,N_5304);
or U7744 (N_7744,N_4996,N_5611);
nor U7745 (N_7745,N_4259,N_4852);
nand U7746 (N_7746,N_5296,N_4297);
xnor U7747 (N_7747,N_5844,N_5124);
xor U7748 (N_7748,N_5026,N_4544);
nor U7749 (N_7749,N_4349,N_5827);
or U7750 (N_7750,N_5386,N_5281);
or U7751 (N_7751,N_4397,N_4587);
nand U7752 (N_7752,N_5484,N_4974);
and U7753 (N_7753,N_5101,N_4182);
and U7754 (N_7754,N_5153,N_4757);
nor U7755 (N_7755,N_5268,N_4806);
nand U7756 (N_7756,N_4441,N_4063);
xor U7757 (N_7757,N_4091,N_5091);
nor U7758 (N_7758,N_4331,N_5939);
or U7759 (N_7759,N_4859,N_5209);
nand U7760 (N_7760,N_4750,N_4213);
nand U7761 (N_7761,N_4253,N_4928);
and U7762 (N_7762,N_4286,N_4256);
nand U7763 (N_7763,N_4207,N_4472);
nor U7764 (N_7764,N_5453,N_5048);
or U7765 (N_7765,N_4126,N_4098);
nor U7766 (N_7766,N_5805,N_5342);
nand U7767 (N_7767,N_4407,N_5187);
nand U7768 (N_7768,N_4009,N_5996);
nor U7769 (N_7769,N_5675,N_5690);
and U7770 (N_7770,N_5495,N_5593);
xnor U7771 (N_7771,N_5323,N_5433);
nand U7772 (N_7772,N_5193,N_4412);
nor U7773 (N_7773,N_4069,N_5750);
or U7774 (N_7774,N_4958,N_5143);
or U7775 (N_7775,N_4196,N_5132);
xnor U7776 (N_7776,N_5982,N_5429);
nor U7777 (N_7777,N_5352,N_4237);
and U7778 (N_7778,N_5913,N_5167);
or U7779 (N_7779,N_5904,N_4966);
or U7780 (N_7780,N_4617,N_5174);
and U7781 (N_7781,N_4348,N_5416);
or U7782 (N_7782,N_4211,N_4321);
nand U7783 (N_7783,N_4073,N_4630);
nor U7784 (N_7784,N_5262,N_4411);
nor U7785 (N_7785,N_4486,N_5355);
nor U7786 (N_7786,N_5727,N_4864);
nor U7787 (N_7787,N_4396,N_5702);
and U7788 (N_7788,N_5995,N_5684);
and U7789 (N_7789,N_5211,N_4233);
nor U7790 (N_7790,N_4166,N_5422);
or U7791 (N_7791,N_4001,N_5472);
nor U7792 (N_7792,N_4442,N_4409);
or U7793 (N_7793,N_5845,N_5888);
xor U7794 (N_7794,N_5643,N_5648);
xor U7795 (N_7795,N_5003,N_5956);
nor U7796 (N_7796,N_5374,N_4311);
nand U7797 (N_7797,N_5323,N_4160);
or U7798 (N_7798,N_4116,N_5727);
xor U7799 (N_7799,N_4036,N_4971);
and U7800 (N_7800,N_4018,N_4888);
and U7801 (N_7801,N_4500,N_5006);
xnor U7802 (N_7802,N_4767,N_4224);
nor U7803 (N_7803,N_5915,N_4546);
xnor U7804 (N_7804,N_5997,N_5940);
nor U7805 (N_7805,N_4845,N_4638);
or U7806 (N_7806,N_5530,N_5206);
xor U7807 (N_7807,N_5821,N_4073);
or U7808 (N_7808,N_5230,N_5256);
nand U7809 (N_7809,N_4668,N_4378);
and U7810 (N_7810,N_5456,N_5712);
or U7811 (N_7811,N_4947,N_4801);
and U7812 (N_7812,N_4778,N_5319);
nand U7813 (N_7813,N_5337,N_5189);
nand U7814 (N_7814,N_4728,N_5057);
and U7815 (N_7815,N_5304,N_4469);
nand U7816 (N_7816,N_4975,N_4841);
xnor U7817 (N_7817,N_4022,N_4864);
or U7818 (N_7818,N_4982,N_4044);
or U7819 (N_7819,N_5710,N_4476);
and U7820 (N_7820,N_5995,N_5194);
and U7821 (N_7821,N_4212,N_4234);
nor U7822 (N_7822,N_5754,N_5520);
nand U7823 (N_7823,N_5965,N_5469);
nor U7824 (N_7824,N_5990,N_5159);
nor U7825 (N_7825,N_4089,N_5605);
or U7826 (N_7826,N_5758,N_4061);
and U7827 (N_7827,N_5189,N_5342);
nand U7828 (N_7828,N_5577,N_5966);
xor U7829 (N_7829,N_4031,N_4981);
nand U7830 (N_7830,N_4741,N_4957);
or U7831 (N_7831,N_4005,N_5063);
nor U7832 (N_7832,N_4689,N_4861);
nor U7833 (N_7833,N_5505,N_4554);
xnor U7834 (N_7834,N_5117,N_4307);
and U7835 (N_7835,N_5940,N_5626);
nor U7836 (N_7836,N_4644,N_5440);
xnor U7837 (N_7837,N_4223,N_4249);
nor U7838 (N_7838,N_4994,N_5582);
or U7839 (N_7839,N_5104,N_5992);
or U7840 (N_7840,N_5460,N_4203);
xnor U7841 (N_7841,N_4416,N_4373);
nor U7842 (N_7842,N_5560,N_4339);
xor U7843 (N_7843,N_5125,N_4191);
or U7844 (N_7844,N_4241,N_5292);
nand U7845 (N_7845,N_4366,N_4686);
nor U7846 (N_7846,N_5261,N_5648);
xnor U7847 (N_7847,N_5086,N_5885);
nor U7848 (N_7848,N_4864,N_4698);
and U7849 (N_7849,N_4955,N_4604);
nor U7850 (N_7850,N_5957,N_4913);
and U7851 (N_7851,N_4718,N_5258);
nor U7852 (N_7852,N_4662,N_5787);
nor U7853 (N_7853,N_5350,N_5241);
nand U7854 (N_7854,N_4141,N_4683);
and U7855 (N_7855,N_5202,N_4857);
nor U7856 (N_7856,N_5054,N_4163);
xnor U7857 (N_7857,N_5137,N_5378);
nand U7858 (N_7858,N_5936,N_4468);
nand U7859 (N_7859,N_5152,N_4617);
and U7860 (N_7860,N_5229,N_4306);
xor U7861 (N_7861,N_5331,N_5286);
xnor U7862 (N_7862,N_4327,N_4875);
and U7863 (N_7863,N_5367,N_5874);
or U7864 (N_7864,N_4921,N_4029);
xnor U7865 (N_7865,N_5246,N_5928);
nor U7866 (N_7866,N_4393,N_5547);
nor U7867 (N_7867,N_4163,N_5328);
and U7868 (N_7868,N_4643,N_5654);
xnor U7869 (N_7869,N_5199,N_4309);
nand U7870 (N_7870,N_4888,N_5505);
nor U7871 (N_7871,N_4287,N_4058);
xor U7872 (N_7872,N_5547,N_4477);
or U7873 (N_7873,N_5106,N_5936);
or U7874 (N_7874,N_4974,N_4544);
nand U7875 (N_7875,N_5120,N_5648);
or U7876 (N_7876,N_4125,N_5539);
xnor U7877 (N_7877,N_5282,N_4274);
and U7878 (N_7878,N_5100,N_5781);
and U7879 (N_7879,N_4433,N_4910);
nor U7880 (N_7880,N_5985,N_4466);
nor U7881 (N_7881,N_5313,N_4529);
nand U7882 (N_7882,N_4267,N_4473);
and U7883 (N_7883,N_4262,N_5427);
and U7884 (N_7884,N_5396,N_4046);
nand U7885 (N_7885,N_4006,N_4655);
nand U7886 (N_7886,N_4540,N_5154);
xor U7887 (N_7887,N_4121,N_5645);
nor U7888 (N_7888,N_5500,N_5685);
and U7889 (N_7889,N_4510,N_4850);
and U7890 (N_7890,N_5233,N_4208);
xor U7891 (N_7891,N_5213,N_5270);
xnor U7892 (N_7892,N_4245,N_4386);
or U7893 (N_7893,N_5811,N_4670);
nor U7894 (N_7894,N_5163,N_4505);
nor U7895 (N_7895,N_5747,N_5906);
or U7896 (N_7896,N_4902,N_4032);
nor U7897 (N_7897,N_5291,N_5529);
or U7898 (N_7898,N_4413,N_4205);
nand U7899 (N_7899,N_5497,N_4364);
and U7900 (N_7900,N_4727,N_5552);
xnor U7901 (N_7901,N_4630,N_5176);
nand U7902 (N_7902,N_5171,N_5209);
nand U7903 (N_7903,N_5218,N_4895);
nand U7904 (N_7904,N_4682,N_4579);
or U7905 (N_7905,N_4871,N_4993);
nand U7906 (N_7906,N_4604,N_4733);
and U7907 (N_7907,N_4080,N_5852);
or U7908 (N_7908,N_5112,N_4690);
or U7909 (N_7909,N_4164,N_5918);
nand U7910 (N_7910,N_5240,N_4699);
xnor U7911 (N_7911,N_4641,N_4433);
xnor U7912 (N_7912,N_5571,N_5883);
and U7913 (N_7913,N_4434,N_5202);
and U7914 (N_7914,N_5150,N_4334);
nand U7915 (N_7915,N_5777,N_4773);
nand U7916 (N_7916,N_5575,N_5206);
nand U7917 (N_7917,N_5757,N_4666);
nand U7918 (N_7918,N_5630,N_5414);
or U7919 (N_7919,N_4203,N_4611);
and U7920 (N_7920,N_5758,N_5321);
xor U7921 (N_7921,N_5599,N_4196);
xnor U7922 (N_7922,N_5883,N_5493);
or U7923 (N_7923,N_5400,N_5887);
xor U7924 (N_7924,N_5471,N_4724);
or U7925 (N_7925,N_5995,N_5196);
nor U7926 (N_7926,N_4199,N_4593);
or U7927 (N_7927,N_5248,N_5039);
nor U7928 (N_7928,N_5343,N_5913);
or U7929 (N_7929,N_5356,N_5428);
nand U7930 (N_7930,N_4794,N_5995);
or U7931 (N_7931,N_4373,N_5787);
nor U7932 (N_7932,N_5530,N_4479);
nand U7933 (N_7933,N_5736,N_5734);
xnor U7934 (N_7934,N_4338,N_5676);
and U7935 (N_7935,N_5851,N_4059);
xor U7936 (N_7936,N_4292,N_5306);
nand U7937 (N_7937,N_4759,N_5104);
or U7938 (N_7938,N_5672,N_5055);
or U7939 (N_7939,N_5383,N_4773);
and U7940 (N_7940,N_5340,N_4450);
or U7941 (N_7941,N_5730,N_4674);
or U7942 (N_7942,N_4208,N_4342);
and U7943 (N_7943,N_5876,N_4499);
or U7944 (N_7944,N_5316,N_5914);
or U7945 (N_7945,N_5660,N_4664);
nand U7946 (N_7946,N_4826,N_4965);
nand U7947 (N_7947,N_5781,N_5825);
and U7948 (N_7948,N_5047,N_5287);
and U7949 (N_7949,N_5648,N_5280);
and U7950 (N_7950,N_4439,N_5235);
xnor U7951 (N_7951,N_4535,N_4645);
nand U7952 (N_7952,N_4515,N_4707);
or U7953 (N_7953,N_4619,N_5814);
nand U7954 (N_7954,N_4360,N_5813);
nand U7955 (N_7955,N_4187,N_4924);
nand U7956 (N_7956,N_5501,N_4973);
xor U7957 (N_7957,N_4311,N_4971);
or U7958 (N_7958,N_5448,N_5511);
nand U7959 (N_7959,N_5681,N_5915);
xor U7960 (N_7960,N_5940,N_4699);
or U7961 (N_7961,N_5016,N_4271);
or U7962 (N_7962,N_4366,N_5754);
nand U7963 (N_7963,N_5331,N_4145);
xnor U7964 (N_7964,N_5542,N_5327);
or U7965 (N_7965,N_4097,N_4384);
nor U7966 (N_7966,N_4814,N_4268);
or U7967 (N_7967,N_5772,N_5349);
nand U7968 (N_7968,N_4858,N_4722);
nand U7969 (N_7969,N_4030,N_5504);
or U7970 (N_7970,N_5946,N_5694);
nand U7971 (N_7971,N_5065,N_5127);
xnor U7972 (N_7972,N_4110,N_5147);
or U7973 (N_7973,N_4702,N_4825);
or U7974 (N_7974,N_5233,N_4240);
nand U7975 (N_7975,N_4287,N_5247);
or U7976 (N_7976,N_5524,N_4398);
nand U7977 (N_7977,N_4109,N_5694);
and U7978 (N_7978,N_5724,N_4862);
nand U7979 (N_7979,N_5302,N_4675);
or U7980 (N_7980,N_4262,N_5691);
or U7981 (N_7981,N_5949,N_5942);
and U7982 (N_7982,N_5799,N_5020);
nor U7983 (N_7983,N_5835,N_5122);
nand U7984 (N_7984,N_4915,N_5321);
and U7985 (N_7985,N_4929,N_4008);
or U7986 (N_7986,N_5951,N_4006);
nand U7987 (N_7987,N_4732,N_5081);
nand U7988 (N_7988,N_4198,N_4377);
or U7989 (N_7989,N_5056,N_4247);
or U7990 (N_7990,N_4606,N_4521);
or U7991 (N_7991,N_4180,N_4001);
or U7992 (N_7992,N_5197,N_4771);
and U7993 (N_7993,N_4416,N_5099);
nand U7994 (N_7994,N_5589,N_4885);
xor U7995 (N_7995,N_4459,N_4922);
nand U7996 (N_7996,N_5190,N_5335);
and U7997 (N_7997,N_5765,N_5961);
nand U7998 (N_7998,N_4916,N_5955);
and U7999 (N_7999,N_4541,N_4558);
xor U8000 (N_8000,N_7925,N_7835);
xnor U8001 (N_8001,N_7732,N_6051);
nor U8002 (N_8002,N_7453,N_7298);
and U8003 (N_8003,N_6567,N_6751);
nor U8004 (N_8004,N_6017,N_7476);
nand U8005 (N_8005,N_7147,N_7444);
and U8006 (N_8006,N_6439,N_6163);
and U8007 (N_8007,N_7456,N_6294);
nor U8008 (N_8008,N_6870,N_7914);
xnor U8009 (N_8009,N_6280,N_7374);
or U8010 (N_8010,N_7826,N_7270);
nor U8011 (N_8011,N_6518,N_7040);
nand U8012 (N_8012,N_6995,N_6820);
and U8013 (N_8013,N_6049,N_6010);
nor U8014 (N_8014,N_7552,N_7803);
nor U8015 (N_8015,N_7322,N_6403);
nor U8016 (N_8016,N_6965,N_7787);
xnor U8017 (N_8017,N_6832,N_7435);
nor U8018 (N_8018,N_6967,N_7119);
xnor U8019 (N_8019,N_7655,N_6792);
nand U8020 (N_8020,N_6848,N_6709);
or U8021 (N_8021,N_7186,N_7929);
xnor U8022 (N_8022,N_6485,N_7267);
and U8023 (N_8023,N_6175,N_7092);
xor U8024 (N_8024,N_7184,N_6566);
or U8025 (N_8025,N_6934,N_6663);
nor U8026 (N_8026,N_6956,N_7100);
nor U8027 (N_8027,N_6152,N_7664);
nand U8028 (N_8028,N_6346,N_6464);
nand U8029 (N_8029,N_7897,N_7421);
nor U8030 (N_8030,N_6080,N_6739);
xor U8031 (N_8031,N_7351,N_7551);
nand U8032 (N_8032,N_7955,N_7229);
nor U8033 (N_8033,N_6826,N_6980);
and U8034 (N_8034,N_6181,N_7866);
and U8035 (N_8035,N_7341,N_6539);
and U8036 (N_8036,N_7534,N_6386);
nor U8037 (N_8037,N_6374,N_7556);
nor U8038 (N_8038,N_7756,N_7503);
xor U8039 (N_8039,N_7859,N_6332);
or U8040 (N_8040,N_7166,N_6930);
and U8041 (N_8041,N_7360,N_6693);
or U8042 (N_8042,N_7144,N_7523);
nor U8043 (N_8043,N_7297,N_7046);
and U8044 (N_8044,N_6284,N_6218);
xnor U8045 (N_8045,N_7012,N_7755);
and U8046 (N_8046,N_7057,N_6041);
and U8047 (N_8047,N_7437,N_6476);
nor U8048 (N_8048,N_7343,N_7828);
nor U8049 (N_8049,N_7068,N_6506);
nand U8050 (N_8050,N_6154,N_6846);
and U8051 (N_8051,N_6400,N_7804);
nor U8052 (N_8052,N_6678,N_7663);
or U8053 (N_8053,N_7284,N_6745);
xnor U8054 (N_8054,N_6918,N_7065);
and U8055 (N_8055,N_6653,N_6096);
nor U8056 (N_8056,N_7404,N_6406);
and U8057 (N_8057,N_7011,N_7299);
or U8058 (N_8058,N_7475,N_7987);
xnor U8059 (N_8059,N_6727,N_7561);
nand U8060 (N_8060,N_7771,N_7840);
nand U8061 (N_8061,N_7169,N_7443);
or U8062 (N_8062,N_6904,N_6951);
nor U8063 (N_8063,N_6587,N_6954);
xor U8064 (N_8064,N_7560,N_6033);
or U8065 (N_8065,N_6839,N_7362);
and U8066 (N_8066,N_6471,N_7954);
and U8067 (N_8067,N_6553,N_7191);
nor U8068 (N_8068,N_7535,N_6755);
and U8069 (N_8069,N_7539,N_7644);
and U8070 (N_8070,N_7668,N_7701);
nand U8071 (N_8071,N_7564,N_7905);
nand U8072 (N_8072,N_7164,N_7020);
xor U8073 (N_8073,N_6586,N_7146);
and U8074 (N_8074,N_6398,N_7510);
nand U8075 (N_8075,N_6185,N_7649);
xnor U8076 (N_8076,N_6793,N_6379);
nand U8077 (N_8077,N_6874,N_7818);
or U8078 (N_8078,N_6468,N_6768);
and U8079 (N_8079,N_6784,N_7530);
xnor U8080 (N_8080,N_7318,N_7436);
xor U8081 (N_8081,N_7139,N_6861);
nand U8082 (N_8082,N_7156,N_7347);
or U8083 (N_8083,N_6757,N_6859);
and U8084 (N_8084,N_6525,N_6533);
and U8085 (N_8085,N_7086,N_7189);
nand U8086 (N_8086,N_7201,N_7855);
nand U8087 (N_8087,N_7969,N_7354);
or U8088 (N_8088,N_7494,N_7747);
or U8089 (N_8089,N_6824,N_7678);
and U8090 (N_8090,N_6449,N_6576);
nand U8091 (N_8091,N_6221,N_6458);
xor U8092 (N_8092,N_7682,N_6062);
nand U8093 (N_8093,N_6548,N_6252);
nand U8094 (N_8094,N_6461,N_6531);
or U8095 (N_8095,N_7465,N_7231);
xnor U8096 (N_8096,N_7827,N_7137);
and U8097 (N_8097,N_6162,N_7010);
nand U8098 (N_8098,N_6882,N_6121);
and U8099 (N_8099,N_6030,N_6281);
xor U8100 (N_8100,N_7834,N_6949);
xnor U8101 (N_8101,N_7457,N_6027);
nand U8102 (N_8102,N_6470,N_7519);
or U8103 (N_8103,N_7087,N_6236);
xor U8104 (N_8104,N_7043,N_7016);
nor U8105 (N_8105,N_7735,N_7036);
and U8106 (N_8106,N_7285,N_7780);
nor U8107 (N_8107,N_7590,N_7625);
nand U8108 (N_8108,N_7965,N_6606);
or U8109 (N_8109,N_6306,N_6056);
xor U8110 (N_8110,N_6372,N_6927);
xor U8111 (N_8111,N_7513,N_6691);
xnor U8112 (N_8112,N_7093,N_6546);
nand U8113 (N_8113,N_6802,N_6625);
xnor U8114 (N_8114,N_6358,N_6766);
and U8115 (N_8115,N_7097,N_6047);
nand U8116 (N_8116,N_6535,N_7083);
nor U8117 (N_8117,N_7778,N_6872);
xnor U8118 (N_8118,N_7873,N_6522);
nor U8119 (N_8119,N_7366,N_7659);
nor U8120 (N_8120,N_6922,N_6735);
xor U8121 (N_8121,N_7788,N_6001);
nand U8122 (N_8122,N_6193,N_6662);
xor U8123 (N_8123,N_6925,N_7054);
or U8124 (N_8124,N_7143,N_7195);
nand U8125 (N_8125,N_6694,N_6437);
xnor U8126 (N_8126,N_7976,N_6078);
and U8127 (N_8127,N_6559,N_6367);
nor U8128 (N_8128,N_6058,N_7638);
or U8129 (N_8129,N_6699,N_6749);
or U8130 (N_8130,N_7240,N_6043);
nand U8131 (N_8131,N_7396,N_6005);
and U8132 (N_8132,N_6420,N_6720);
nand U8133 (N_8133,N_6417,N_6909);
nor U8134 (N_8134,N_6764,N_6838);
xnor U8135 (N_8135,N_7723,N_7591);
xor U8136 (N_8136,N_7041,N_7286);
and U8137 (N_8137,N_7142,N_6127);
nor U8138 (N_8138,N_6584,N_7162);
and U8139 (N_8139,N_7015,N_7709);
xor U8140 (N_8140,N_6459,N_7173);
or U8141 (N_8141,N_6184,N_7849);
or U8142 (N_8142,N_6462,N_7182);
and U8143 (N_8143,N_6232,N_7727);
nor U8144 (N_8144,N_7109,N_7848);
or U8145 (N_8145,N_7952,N_7931);
nor U8146 (N_8146,N_6677,N_7687);
xor U8147 (N_8147,N_7837,N_6512);
nand U8148 (N_8148,N_6300,N_7630);
or U8149 (N_8149,N_6270,N_6344);
or U8150 (N_8150,N_6960,N_7688);
xnor U8151 (N_8151,N_6979,N_6266);
and U8152 (N_8152,N_6151,N_6724);
nand U8153 (N_8153,N_7053,N_6167);
nand U8154 (N_8154,N_7488,N_7149);
or U8155 (N_8155,N_7052,N_7192);
nand U8156 (N_8156,N_7288,N_6070);
xor U8157 (N_8157,N_7992,N_7643);
or U8158 (N_8158,N_6238,N_6465);
or U8159 (N_8159,N_7814,N_7310);
xnor U8160 (N_8160,N_7907,N_6765);
or U8161 (N_8161,N_6276,N_7857);
and U8162 (N_8162,N_7593,N_6711);
nand U8163 (N_8163,N_6227,N_7677);
or U8164 (N_8164,N_7167,N_6338);
nor U8165 (N_8165,N_7268,N_7022);
xor U8166 (N_8166,N_6923,N_7283);
xor U8167 (N_8167,N_6165,N_6320);
and U8168 (N_8168,N_7380,N_7584);
or U8169 (N_8169,N_6000,N_7433);
and U8170 (N_8170,N_6953,N_7389);
and U8171 (N_8171,N_6989,N_7737);
or U8172 (N_8172,N_6640,N_6975);
xor U8173 (N_8173,N_6472,N_6772);
nand U8174 (N_8174,N_6095,N_6851);
nor U8175 (N_8175,N_6297,N_7988);
and U8176 (N_8176,N_6771,N_6575);
nor U8177 (N_8177,N_7572,N_7180);
nor U8178 (N_8178,N_7235,N_6208);
nor U8179 (N_8179,N_6326,N_7439);
or U8180 (N_8180,N_7023,N_7796);
nor U8181 (N_8181,N_7317,N_7027);
nor U8182 (N_8182,N_7750,N_7926);
or U8183 (N_8183,N_6288,N_6253);
and U8184 (N_8184,N_6045,N_6251);
or U8185 (N_8185,N_6776,N_7508);
and U8186 (N_8186,N_6378,N_6090);
nor U8187 (N_8187,N_7069,N_7853);
nor U8188 (N_8188,N_7058,N_7978);
or U8189 (N_8189,N_6307,N_7580);
and U8190 (N_8190,N_7882,N_7667);
and U8191 (N_8191,N_6556,N_6313);
xor U8192 (N_8192,N_6538,N_7919);
and U8193 (N_8193,N_7382,N_6170);
or U8194 (N_8194,N_7763,N_6550);
nor U8195 (N_8195,N_6250,N_7448);
nand U8196 (N_8196,N_7908,N_7281);
or U8197 (N_8197,N_7416,N_7953);
and U8198 (N_8198,N_6421,N_7924);
and U8199 (N_8199,N_7759,N_6490);
and U8200 (N_8200,N_6487,N_6209);
nand U8201 (N_8201,N_6079,N_7155);
nor U8202 (N_8202,N_6528,N_7685);
and U8203 (N_8203,N_6275,N_7589);
and U8204 (N_8204,N_7863,N_6274);
nand U8205 (N_8205,N_6039,N_6622);
xnor U8206 (N_8206,N_7632,N_6617);
and U8207 (N_8207,N_6428,N_6685);
and U8208 (N_8208,N_7316,N_6329);
or U8209 (N_8209,N_6671,N_6106);
or U8210 (N_8210,N_6945,N_7399);
and U8211 (N_8211,N_7761,N_6588);
nor U8212 (N_8212,N_7934,N_6876);
xor U8213 (N_8213,N_6821,N_6664);
and U8214 (N_8214,N_7883,N_6361);
xor U8215 (N_8215,N_6636,N_6524);
or U8216 (N_8216,N_6444,N_6124);
xor U8217 (N_8217,N_6189,N_6081);
nor U8218 (N_8218,N_6074,N_7912);
and U8219 (N_8219,N_6198,N_7946);
nor U8220 (N_8220,N_6686,N_6454);
xor U8221 (N_8221,N_7274,N_7982);
xor U8222 (N_8222,N_7466,N_7485);
nor U8223 (N_8223,N_6624,N_7082);
xnor U8224 (N_8224,N_6059,N_6534);
nand U8225 (N_8225,N_7636,N_7152);
or U8226 (N_8226,N_7333,N_7148);
xor U8227 (N_8227,N_7061,N_6948);
xor U8228 (N_8228,N_6635,N_6900);
nand U8229 (N_8229,N_6753,N_7246);
and U8230 (N_8230,N_7786,N_6407);
or U8231 (N_8231,N_6651,N_6639);
or U8232 (N_8232,N_7116,N_7626);
or U8233 (N_8233,N_7712,N_7260);
xor U8234 (N_8234,N_7656,N_7558);
nor U8235 (N_8235,N_7581,N_6111);
xnor U8236 (N_8236,N_7263,N_6705);
nor U8237 (N_8237,N_6133,N_7816);
xor U8238 (N_8238,N_7261,N_7356);
or U8239 (N_8239,N_7337,N_6268);
xnor U8240 (N_8240,N_6263,N_7095);
nand U8241 (N_8241,N_7110,N_6173);
and U8242 (N_8242,N_6940,N_7484);
or U8243 (N_8243,N_6865,N_7077);
and U8244 (N_8244,N_6259,N_6593);
or U8245 (N_8245,N_7008,N_7899);
nand U8246 (N_8246,N_7486,N_7205);
or U8247 (N_8247,N_6168,N_6473);
nor U8248 (N_8248,N_7579,N_7797);
and U8249 (N_8249,N_6537,N_6767);
or U8250 (N_8250,N_6012,N_6199);
nor U8251 (N_8251,N_7131,N_7567);
nor U8252 (N_8252,N_6893,N_6939);
nand U8253 (N_8253,N_6996,N_6862);
nor U8254 (N_8254,N_7798,N_6177);
nand U8255 (N_8255,N_7839,N_6648);
nor U8256 (N_8256,N_6710,N_7779);
xnor U8257 (N_8257,N_7895,N_6023);
nor U8258 (N_8258,N_6101,N_7107);
nand U8259 (N_8259,N_6069,N_7544);
and U8260 (N_8260,N_6613,N_7212);
nand U8261 (N_8261,N_7624,N_7427);
and U8262 (N_8262,N_6423,N_7614);
or U8263 (N_8263,N_6373,N_7699);
or U8264 (N_8264,N_7400,N_7193);
xor U8265 (N_8265,N_6126,N_7936);
or U8266 (N_8266,N_7860,N_7171);
nor U8267 (N_8267,N_6585,N_6176);
nor U8268 (N_8268,N_7277,N_7214);
nand U8269 (N_8269,N_7616,N_6331);
nand U8270 (N_8270,N_6670,N_6381);
or U8271 (N_8271,N_6321,N_7282);
xnor U8272 (N_8272,N_6333,N_7035);
and U8273 (N_8273,N_6169,N_6491);
xor U8274 (N_8274,N_7304,N_6216);
and U8275 (N_8275,N_7174,N_6630);
or U8276 (N_8276,N_7536,N_6246);
or U8277 (N_8277,N_6750,N_7696);
xnor U8278 (N_8278,N_6393,N_7017);
or U8279 (N_8279,N_7800,N_6103);
and U8280 (N_8280,N_6530,N_7940);
nand U8281 (N_8281,N_7592,N_7881);
or U8282 (N_8282,N_7241,N_6201);
nand U8283 (N_8283,N_6656,N_6702);
nor U8284 (N_8284,N_6409,N_6233);
nor U8285 (N_8285,N_7824,N_7722);
or U8286 (N_8286,N_7296,N_6113);
or U8287 (N_8287,N_7922,N_6130);
nor U8288 (N_8288,N_6489,N_6804);
xor U8289 (N_8289,N_7802,N_7669);
xor U8290 (N_8290,N_6778,N_6917);
nor U8291 (N_8291,N_7150,N_7204);
or U8292 (N_8292,N_6138,N_6797);
or U8293 (N_8293,N_6427,N_6657);
nor U8294 (N_8294,N_6944,N_6431);
or U8295 (N_8295,N_6695,N_7216);
nand U8296 (N_8296,N_6898,N_7398);
or U8297 (N_8297,N_7898,N_6053);
and U8298 (N_8298,N_6264,N_7305);
and U8299 (N_8299,N_6597,N_7122);
or U8300 (N_8300,N_7447,N_7179);
or U8301 (N_8301,N_6738,N_6370);
and U8302 (N_8302,N_7608,N_6383);
and U8303 (N_8303,N_7138,N_7446);
nor U8304 (N_8304,N_7689,N_6669);
xor U8305 (N_8305,N_7906,N_7408);
and U8306 (N_8306,N_7440,N_7702);
and U8307 (N_8307,N_6616,N_7477);
or U8308 (N_8308,N_6502,N_7495);
xor U8309 (N_8309,N_7734,N_6323);
nor U8310 (N_8310,N_7049,N_7044);
xnor U8311 (N_8311,N_6816,N_7964);
xor U8312 (N_8312,N_6615,N_7760);
nand U8313 (N_8313,N_7602,N_7887);
nor U8314 (N_8314,N_7118,N_7715);
or U8315 (N_8315,N_6610,N_6928);
or U8316 (N_8316,N_6048,N_7606);
nand U8317 (N_8317,N_6592,N_7540);
nand U8318 (N_8318,N_6318,N_6003);
and U8319 (N_8319,N_6481,N_6183);
xor U8320 (N_8320,N_7325,N_6661);
nor U8321 (N_8321,N_6384,N_7652);
nand U8322 (N_8322,N_7862,N_7245);
or U8323 (N_8323,N_7806,N_6414);
and U8324 (N_8324,N_7208,N_7514);
nand U8325 (N_8325,N_6571,N_7830);
nand U8326 (N_8326,N_7243,N_7583);
xor U8327 (N_8327,N_6204,N_6086);
nor U8328 (N_8328,N_7575,N_6132);
xor U8329 (N_8329,N_7313,N_6618);
nand U8330 (N_8330,N_7405,N_7612);
xnor U8331 (N_8331,N_6842,N_7418);
xnor U8332 (N_8332,N_7221,N_7364);
or U8333 (N_8333,N_7900,N_7845);
nand U8334 (N_8334,N_6484,N_7213);
xnor U8335 (N_8335,N_7550,N_6878);
nor U8336 (N_8336,N_7629,N_6194);
xor U8337 (N_8337,N_6296,N_7923);
xnor U8338 (N_8338,N_6408,N_7480);
and U8339 (N_8339,N_7868,N_6150);
or U8340 (N_8340,N_6544,N_7370);
xor U8341 (N_8341,N_6976,N_6557);
nand U8342 (N_8342,N_6445,N_7884);
nand U8343 (N_8343,N_6327,N_6603);
or U8344 (N_8344,N_7977,N_7279);
nand U8345 (N_8345,N_6231,N_7791);
or U8346 (N_8346,N_6104,N_7042);
nor U8347 (N_8347,N_6795,N_7153);
or U8348 (N_8348,N_6396,N_7991);
nand U8349 (N_8349,N_6054,N_6971);
nand U8350 (N_8350,N_7335,N_7501);
or U8351 (N_8351,N_7497,N_6282);
nand U8352 (N_8352,N_7258,N_7434);
or U8353 (N_8353,N_6763,N_7469);
or U8354 (N_8354,N_6981,N_7930);
and U8355 (N_8355,N_7247,N_6894);
or U8356 (N_8356,N_7547,N_7822);
or U8357 (N_8357,N_7117,N_7896);
nand U8358 (N_8358,N_6161,N_7273);
nand U8359 (N_8359,N_7995,N_7227);
nor U8360 (N_8360,N_7369,N_6834);
or U8361 (N_8361,N_7176,N_7134);
and U8362 (N_8362,N_6725,N_7031);
xor U8363 (N_8363,N_7030,N_6982);
or U8364 (N_8364,N_7290,N_7419);
and U8365 (N_8365,N_7680,N_7066);
nand U8366 (N_8366,N_7836,N_6600);
nand U8367 (N_8367,N_7817,N_7956);
or U8368 (N_8368,N_6360,N_7295);
xnor U8369 (N_8369,N_7397,N_7294);
or U8370 (N_8370,N_6867,N_6082);
xnor U8371 (N_8371,N_7331,N_6369);
or U8372 (N_8372,N_7051,N_7726);
or U8373 (N_8373,N_6906,N_6721);
nand U8374 (N_8374,N_7464,N_6311);
nor U8375 (N_8375,N_6692,N_6997);
nor U8376 (N_8376,N_6714,N_7459);
nor U8377 (N_8377,N_7971,N_7809);
xor U8378 (N_8378,N_7468,N_7743);
nand U8379 (N_8379,N_7864,N_6889);
and U8380 (N_8380,N_6272,N_7665);
nor U8381 (N_8381,N_7757,N_7232);
and U8382 (N_8382,N_6273,N_6769);
nor U8383 (N_8383,N_7423,N_6083);
nand U8384 (N_8384,N_7605,N_7917);
nor U8385 (N_8385,N_7344,N_6418);
xor U8386 (N_8386,N_7666,N_7002);
nand U8387 (N_8387,N_6959,N_6395);
xnor U8388 (N_8388,N_7504,N_6654);
nand U8389 (N_8389,N_6309,N_6741);
or U8390 (N_8390,N_6783,N_7951);
xor U8391 (N_8391,N_7811,N_7371);
nand U8392 (N_8392,N_7072,N_7937);
nor U8393 (N_8393,N_6827,N_7777);
nand U8394 (N_8394,N_7517,N_6277);
and U8395 (N_8395,N_7932,N_7808);
nand U8396 (N_8396,N_6747,N_7160);
nand U8397 (N_8397,N_6703,N_6697);
xor U8398 (N_8398,N_6479,N_6938);
nor U8399 (N_8399,N_7843,N_7562);
xnor U8400 (N_8400,N_6092,N_7559);
xor U8401 (N_8401,N_6496,N_6447);
nor U8402 (N_8402,N_7081,N_6153);
nand U8403 (N_8403,N_6060,N_6542);
and U8404 (N_8404,N_7493,N_6258);
nand U8405 (N_8405,N_7025,N_6052);
nor U8406 (N_8406,N_7675,N_6493);
nand U8407 (N_8407,N_6623,N_7377);
xor U8408 (N_8408,N_7319,N_7928);
xor U8409 (N_8409,N_7684,N_7762);
or U8410 (N_8410,N_6598,N_6290);
and U8411 (N_8411,N_7375,N_6279);
nor U8412 (N_8412,N_7901,N_7738);
nand U8413 (N_8413,N_7048,N_7425);
or U8414 (N_8414,N_7957,N_6093);
xnor U8415 (N_8415,N_7242,N_7455);
or U8416 (N_8416,N_7628,N_6128);
and U8417 (N_8417,N_7365,N_7121);
xnor U8418 (N_8418,N_7880,N_6990);
nor U8419 (N_8419,N_6164,N_7846);
xnor U8420 (N_8420,N_6422,N_7522);
nand U8421 (N_8421,N_6425,N_7067);
nand U8422 (N_8422,N_6336,N_6907);
and U8423 (N_8423,N_6419,N_7479);
or U8424 (N_8424,N_7753,N_7003);
nand U8425 (N_8425,N_6505,N_7553);
nor U8426 (N_8426,N_7251,N_6782);
xor U8427 (N_8427,N_7627,N_7617);
nand U8428 (N_8428,N_6740,N_6565);
and U8429 (N_8429,N_7733,N_6785);
and U8430 (N_8430,N_7461,N_6324);
xor U8431 (N_8431,N_6958,N_7491);
or U8432 (N_8432,N_7238,N_7289);
nand U8433 (N_8433,N_6174,N_6013);
nand U8434 (N_8434,N_6123,N_6415);
and U8435 (N_8435,N_6115,N_6364);
nor U8436 (N_8436,N_7492,N_6545);
and U8437 (N_8437,N_7115,N_7594);
and U8438 (N_8438,N_6140,N_6145);
or U8439 (N_8439,N_6105,N_7168);
or U8440 (N_8440,N_6845,N_7004);
nand U8441 (N_8441,N_7686,N_7228);
and U8442 (N_8442,N_7801,N_6511);
or U8443 (N_8443,N_6774,N_6760);
nand U8444 (N_8444,N_6143,N_6643);
xor U8445 (N_8445,N_6158,N_6914);
nand U8446 (N_8446,N_6915,N_6941);
and U8447 (N_8447,N_7740,N_6203);
nand U8448 (N_8448,N_7939,N_6682);
and U8449 (N_8449,N_6098,N_6837);
xor U8450 (N_8450,N_7783,N_7357);
and U8451 (N_8451,N_7555,N_6180);
xnor U8452 (N_8452,N_6399,N_7236);
xor U8453 (N_8453,N_6494,N_6166);
and U8454 (N_8454,N_6310,N_7890);
and U8455 (N_8455,N_6581,N_7332);
or U8456 (N_8456,N_7515,N_6637);
xnor U8457 (N_8457,N_6368,N_6513);
nand U8458 (N_8458,N_6933,N_7970);
nand U8459 (N_8459,N_6629,N_7078);
xor U8460 (N_8460,N_7714,N_7372);
nand U8461 (N_8461,N_7785,N_7154);
nand U8462 (N_8462,N_6810,N_6325);
and U8463 (N_8463,N_7639,N_6527);
nand U8464 (N_8464,N_6706,N_7615);
or U8465 (N_8465,N_7610,N_7949);
and U8466 (N_8466,N_7799,N_7063);
nand U8467 (N_8467,N_6228,N_6962);
or U8468 (N_8468,N_7032,N_7159);
or U8469 (N_8469,N_7451,N_7112);
nor U8470 (N_8470,N_6676,N_6002);
or U8471 (N_8471,N_6936,N_7691);
or U8472 (N_8472,N_7793,N_6988);
or U8473 (N_8473,N_7359,N_7108);
and U8474 (N_8474,N_7250,N_7026);
nor U8475 (N_8475,N_6813,N_6964);
nand U8476 (N_8476,N_7309,N_7865);
and U8477 (N_8477,N_7528,N_6110);
and U8478 (N_8478,N_7329,N_6032);
nor U8479 (N_8479,N_7631,N_6102);
and U8480 (N_8480,N_7473,N_6779);
and U8481 (N_8481,N_7720,N_7823);
xnor U8482 (N_8482,N_6847,N_6713);
xor U8483 (N_8483,N_7792,N_6883);
and U8484 (N_8484,N_7113,N_7367);
and U8485 (N_8485,N_7654,N_7033);
or U8486 (N_8486,N_7730,N_6224);
nand U8487 (N_8487,N_7203,N_6901);
or U8488 (N_8488,N_6477,N_7394);
nor U8489 (N_8489,N_7782,N_6257);
nor U8490 (N_8490,N_7573,N_7487);
xnor U8491 (N_8491,N_7124,N_7024);
or U8492 (N_8492,N_7234,N_6968);
xnor U8493 (N_8493,N_6343,N_6895);
or U8494 (N_8494,N_7123,N_7463);
xnor U8495 (N_8495,N_7472,N_7429);
nand U8496 (N_8496,N_7815,N_6881);
and U8497 (N_8497,N_7302,N_7140);
and U8498 (N_8498,N_7867,N_6135);
and U8499 (N_8499,N_7960,N_6737);
nand U8500 (N_8500,N_6911,N_7239);
and U8501 (N_8501,N_6025,N_6213);
nor U8502 (N_8502,N_6974,N_7128);
or U8503 (N_8503,N_7520,N_7697);
nand U8504 (N_8504,N_7904,N_6509);
or U8505 (N_8505,N_6404,N_6621);
nand U8506 (N_8506,N_6057,N_7545);
or U8507 (N_8507,N_6991,N_6107);
nor U8508 (N_8508,N_6563,N_6770);
xnor U8509 (N_8509,N_7151,N_6730);
nor U8510 (N_8510,N_7764,N_6903);
nand U8511 (N_8511,N_6902,N_7506);
or U8512 (N_8512,N_7481,N_7972);
or U8513 (N_8513,N_7449,N_6382);
or U8514 (N_8514,N_6411,N_7871);
nor U8515 (N_8515,N_6977,N_7458);
or U8516 (N_8516,N_6947,N_6365);
or U8517 (N_8517,N_6072,N_6202);
nand U8518 (N_8518,N_6410,N_6896);
and U8519 (N_8519,N_7178,N_6853);
or U8520 (N_8520,N_6674,N_7844);
nor U8521 (N_8521,N_6187,N_7407);
nor U8522 (N_8522,N_6608,N_7390);
or U8523 (N_8523,N_6389,N_7102);
and U8524 (N_8524,N_6337,N_6596);
nand U8525 (N_8525,N_6679,N_7266);
nand U8526 (N_8526,N_7974,N_7637);
xor U8527 (N_8527,N_7721,N_6986);
xor U8528 (N_8528,N_6942,N_7280);
and U8529 (N_8529,N_7819,N_6823);
nand U8530 (N_8530,N_6286,N_6743);
or U8531 (N_8531,N_6973,N_6350);
and U8532 (N_8532,N_6602,N_6950);
nand U8533 (N_8533,N_6362,N_6611);
and U8534 (N_8534,N_6214,N_6508);
or U8535 (N_8535,N_7533,N_7690);
nor U8536 (N_8536,N_7916,N_7725);
and U8537 (N_8537,N_6335,N_7876);
xor U8538 (N_8538,N_6808,N_7312);
nor U8539 (N_8539,N_7165,N_7877);
nand U8540 (N_8540,N_6854,N_6789);
nor U8541 (N_8541,N_6007,N_7328);
xnor U8542 (N_8542,N_7129,N_6811);
xor U8543 (N_8543,N_7724,N_6134);
nor U8544 (N_8544,N_6558,N_7420);
xnor U8545 (N_8545,N_6172,N_7450);
nand U8546 (N_8546,N_6469,N_7766);
xor U8547 (N_8547,N_6791,N_7708);
nand U8548 (N_8548,N_7776,N_6833);
and U8549 (N_8549,N_6355,N_7673);
nor U8550 (N_8550,N_6038,N_7271);
xnor U8551 (N_8551,N_6852,N_6429);
nor U8552 (N_8552,N_6044,N_6119);
nor U8553 (N_8553,N_7570,N_7339);
nand U8554 (N_8554,N_7224,N_7990);
nand U8555 (N_8555,N_6929,N_6742);
nand U8556 (N_8556,N_7774,N_7471);
nor U8557 (N_8557,N_6434,N_7368);
or U8558 (N_8558,N_7135,N_6190);
xor U8559 (N_8559,N_6684,N_6523);
xnor U8560 (N_8560,N_6579,N_7745);
nor U8561 (N_8561,N_7106,N_7767);
and U8562 (N_8562,N_6801,N_6295);
or U8563 (N_8563,N_7386,N_6207);
and U8564 (N_8564,N_7962,N_6572);
or U8565 (N_8565,N_6075,N_6131);
or U8566 (N_8566,N_6822,N_7543);
nand U8567 (N_8567,N_6492,N_6293);
nand U8568 (N_8568,N_7911,N_6397);
xnor U8569 (N_8569,N_6316,N_6825);
and U8570 (N_8570,N_7188,N_6435);
or U8571 (N_8571,N_6790,N_6254);
or U8572 (N_8572,N_7693,N_7557);
nand U8573 (N_8573,N_7330,N_6786);
and U8574 (N_8574,N_7829,N_7851);
nor U8575 (N_8575,N_6809,N_6849);
and U8576 (N_8576,N_7620,N_6526);
nor U8577 (N_8577,N_6037,N_6666);
xnor U8578 (N_8578,N_6348,N_6029);
or U8579 (N_8579,N_7085,N_7521);
and U8580 (N_8580,N_7062,N_6380);
nand U8581 (N_8581,N_7635,N_7326);
nor U8582 (N_8582,N_6245,N_6601);
nand U8583 (N_8583,N_6885,N_7736);
xor U8584 (N_8584,N_7483,N_7269);
and U8585 (N_8585,N_6552,N_7237);
nor U8586 (N_8586,N_7181,N_7264);
nor U8587 (N_8587,N_7379,N_6551);
and U8588 (N_8588,N_7327,N_7334);
nor U8589 (N_8589,N_6829,N_6024);
xnor U8590 (N_8590,N_7414,N_6888);
xnor U8591 (N_8591,N_6570,N_6482);
or U8592 (N_8592,N_7306,N_6510);
or U8593 (N_8593,N_7248,N_6803);
and U8594 (N_8594,N_6474,N_7648);
nor U8595 (N_8595,N_6631,N_6256);
nand U8596 (N_8596,N_6521,N_7498);
or U8597 (N_8597,N_6242,N_6599);
and U8598 (N_8598,N_6805,N_6800);
or U8599 (N_8599,N_6660,N_6815);
nand U8600 (N_8600,N_7713,N_7958);
or U8601 (N_8601,N_7099,N_7812);
and U8602 (N_8602,N_6376,N_6880);
xnor U8603 (N_8603,N_7661,N_7537);
nand U8604 (N_8604,N_7452,N_6658);
and U8605 (N_8605,N_6642,N_6718);
or U8606 (N_8606,N_6715,N_7933);
xor U8607 (N_8607,N_6097,N_7292);
nand U8608 (N_8608,N_7301,N_7349);
xnor U8609 (N_8609,N_7942,N_7211);
nor U8610 (N_8610,N_6495,N_7790);
and U8611 (N_8611,N_7833,N_6562);
nand U8612 (N_8612,N_6734,N_7999);
nor U8613 (N_8613,N_6351,N_6818);
nand U8614 (N_8614,N_6466,N_7249);
nand U8615 (N_8615,N_6723,N_7114);
nor U8616 (N_8616,N_6269,N_6887);
xnor U8617 (N_8617,N_6215,N_6301);
nand U8618 (N_8618,N_7910,N_7088);
and U8619 (N_8619,N_7554,N_6314);
and U8620 (N_8620,N_6432,N_6736);
nand U8621 (N_8621,N_7775,N_6205);
and U8622 (N_8622,N_7307,N_7676);
nand U8623 (N_8623,N_7163,N_7532);
or U8624 (N_8624,N_7968,N_6504);
nor U8625 (N_8625,N_6650,N_6347);
nand U8626 (N_8626,N_7096,N_7422);
and U8627 (N_8627,N_6220,N_7604);
xnor U8628 (N_8628,N_7711,N_7752);
or U8629 (N_8629,N_7718,N_6453);
or U8630 (N_8630,N_6334,N_6652);
xor U8631 (N_8631,N_7084,N_7470);
nand U8632 (N_8632,N_6698,N_6239);
and U8633 (N_8633,N_7185,N_7975);
xor U8634 (N_8634,N_6924,N_6704);
nor U8635 (N_8635,N_6392,N_6520);
nand U8636 (N_8636,N_6681,N_7810);
nor U8637 (N_8637,N_6063,N_7621);
xnor U8638 (N_8638,N_7230,N_7569);
xnor U8639 (N_8639,N_6436,N_7984);
and U8640 (N_8640,N_6483,N_7993);
nor U8641 (N_8641,N_6541,N_6019);
nor U8642 (N_8642,N_6433,N_7765);
or U8643 (N_8643,N_7768,N_7961);
nand U8644 (N_8644,N_6564,N_6317);
xor U8645 (N_8645,N_6787,N_6683);
nand U8646 (N_8646,N_6574,N_6514);
nand U8647 (N_8647,N_6758,N_6781);
xor U8648 (N_8648,N_6319,N_6993);
nor U8649 (N_8649,N_6076,N_6265);
or U8650 (N_8650,N_7411,N_6015);
xnor U8651 (N_8651,N_6345,N_7177);
nor U8652 (N_8652,N_6363,N_6426);
xor U8653 (N_8653,N_6619,N_6157);
nand U8654 (N_8654,N_6448,N_7308);
and U8655 (N_8655,N_7111,N_7609);
nand U8656 (N_8656,N_7640,N_7941);
or U8657 (N_8657,N_6773,N_7104);
nor U8658 (N_8658,N_6108,N_7293);
and U8659 (N_8659,N_7794,N_6497);
nor U8660 (N_8660,N_6645,N_6156);
and U8661 (N_8661,N_6831,N_6292);
xnor U8662 (N_8662,N_6775,N_7209);
nor U8663 (N_8663,N_6009,N_7076);
xor U8664 (N_8664,N_6424,N_6021);
and U8665 (N_8665,N_7623,N_6087);
nand U8666 (N_8666,N_6921,N_7145);
and U8667 (N_8667,N_7650,N_7391);
xnor U8668 (N_8668,N_6499,N_6708);
and U8669 (N_8669,N_6308,N_7474);
xnor U8670 (N_8670,N_7613,N_6614);
and U8671 (N_8671,N_6532,N_6966);
nand U8672 (N_8672,N_7413,N_7781);
nor U8673 (N_8673,N_7381,N_6594);
or U8674 (N_8674,N_6690,N_6142);
nand U8675 (N_8675,N_7320,N_6073);
and U8676 (N_8676,N_6726,N_6262);
or U8677 (N_8677,N_6315,N_6589);
nand U8678 (N_8678,N_7772,N_7705);
xor U8679 (N_8679,N_7499,N_6035);
or U8680 (N_8680,N_7383,N_7739);
nor U8681 (N_8681,N_6066,N_7402);
nor U8682 (N_8682,N_6020,N_6830);
xor U8683 (N_8683,N_6197,N_7921);
nand U8684 (N_8684,N_7662,N_7784);
and U8685 (N_8685,N_7651,N_7807);
and U8686 (N_8686,N_7409,N_6014);
or U8687 (N_8687,N_6632,N_6248);
and U8688 (N_8688,N_6696,N_6031);
and U8689 (N_8689,N_7222,N_6026);
xnor U8690 (N_8690,N_6910,N_7909);
nor U8691 (N_8691,N_6046,N_7658);
nor U8692 (N_8692,N_6112,N_6099);
and U8693 (N_8693,N_6109,N_6937);
xnor U8694 (N_8694,N_7039,N_6761);
and U8695 (N_8695,N_7983,N_7161);
nand U8696 (N_8696,N_6516,N_7524);
nand U8697 (N_8697,N_6646,N_7893);
or U8698 (N_8698,N_6884,N_6667);
nor U8699 (N_8699,N_7198,N_6578);
xor U8700 (N_8700,N_6328,N_6120);
nor U8701 (N_8701,N_6868,N_6627);
nor U8702 (N_8702,N_7415,N_7321);
and U8703 (N_8703,N_6788,N_7217);
xnor U8704 (N_8704,N_6247,N_7538);
nand U8705 (N_8705,N_7098,N_7707);
nor U8706 (N_8706,N_6759,N_7588);
and U8707 (N_8707,N_7692,N_7773);
and U8708 (N_8708,N_6628,N_7094);
and U8709 (N_8709,N_7090,N_7199);
nor U8710 (N_8710,N_6016,N_7529);
and U8711 (N_8711,N_7700,N_7585);
nor U8712 (N_8712,N_7598,N_6353);
and U8713 (N_8713,N_6171,N_7641);
or U8714 (N_8714,N_7353,N_7073);
and U8715 (N_8715,N_6515,N_7947);
or U8716 (N_8716,N_6507,N_6701);
xor U8717 (N_8717,N_7175,N_6899);
nand U8718 (N_8718,N_6871,N_6897);
and U8719 (N_8719,N_7315,N_7719);
nor U8720 (N_8720,N_7278,N_6304);
or U8721 (N_8721,N_7393,N_7432);
and U8722 (N_8722,N_6261,N_7006);
nor U8723 (N_8723,N_7670,N_7103);
or U8724 (N_8724,N_7125,N_6322);
and U8725 (N_8725,N_7546,N_7633);
xor U8726 (N_8726,N_6061,N_6855);
nor U8727 (N_8727,N_6129,N_7622);
xnor U8728 (N_8728,N_7080,N_6828);
nor U8729 (N_8729,N_7187,N_6680);
nand U8730 (N_8730,N_6412,N_7599);
xor U8731 (N_8731,N_6722,N_6998);
or U8732 (N_8732,N_6299,N_6034);
or U8733 (N_8733,N_6460,N_7060);
nand U8734 (N_8734,N_7821,N_7505);
nor U8735 (N_8735,N_6935,N_7496);
xor U8736 (N_8736,N_6463,N_7079);
nor U8737 (N_8737,N_7854,N_6573);
xnor U8738 (N_8738,N_7769,N_7028);
nor U8739 (N_8739,N_6040,N_7586);
or U8740 (N_8740,N_6480,N_6577);
xnor U8741 (N_8741,N_6452,N_7345);
xor U8742 (N_8742,N_6312,N_6569);
and U8743 (N_8743,N_6836,N_7417);
xnor U8744 (N_8744,N_6796,N_7348);
or U8745 (N_8745,N_6799,N_7619);
and U8746 (N_8746,N_6359,N_6926);
and U8747 (N_8747,N_7101,N_6712);
nor U8748 (N_8748,N_6707,N_7838);
or U8749 (N_8749,N_7220,N_6920);
nand U8750 (N_8750,N_6728,N_7703);
and U8751 (N_8751,N_6754,N_6777);
xor U8752 (N_8752,N_6285,N_6349);
or U8753 (N_8753,N_6283,N_6467);
nor U8754 (N_8754,N_7259,N_7568);
xor U8755 (N_8755,N_7945,N_6371);
xnor U8756 (N_8756,N_6992,N_7442);
nand U8757 (N_8757,N_7424,N_6241);
and U8758 (N_8758,N_6125,N_7548);
and U8759 (N_8759,N_7126,N_6561);
or U8760 (N_8760,N_7681,N_6401);
and U8761 (N_8761,N_7029,N_7172);
xor U8762 (N_8762,N_6094,N_7311);
nor U8763 (N_8763,N_6085,N_7431);
nand U8764 (N_8764,N_6912,N_7731);
and U8765 (N_8765,N_6554,N_6549);
or U8766 (N_8766,N_7257,N_7136);
or U8767 (N_8767,N_6195,N_7001);
or U8768 (N_8768,N_7218,N_6291);
xnor U8769 (N_8769,N_6441,N_7603);
xor U8770 (N_8770,N_6688,N_7358);
nor U8771 (N_8771,N_6717,N_6385);
nor U8772 (N_8772,N_6812,N_6488);
or U8773 (N_8773,N_6987,N_6858);
nor U8774 (N_8774,N_6857,N_6356);
nand U8775 (N_8775,N_6182,N_7710);
nor U8776 (N_8776,N_7997,N_7373);
nand U8777 (N_8777,N_6866,N_6647);
or U8778 (N_8778,N_7516,N_6687);
nor U8779 (N_8779,N_7482,N_7141);
and U8780 (N_8780,N_7478,N_7454);
or U8781 (N_8781,N_7226,N_7388);
and U8782 (N_8782,N_7075,N_7698);
xnor U8783 (N_8783,N_7938,N_7324);
xor U8784 (N_8784,N_6869,N_7225);
and U8785 (N_8785,N_6844,N_6729);
nor U8786 (N_8786,N_6141,N_7395);
xor U8787 (N_8787,N_7342,N_6873);
nor U8788 (N_8788,N_7361,N_6147);
xnor U8789 (N_8789,N_7255,N_7323);
or U8790 (N_8790,N_6088,N_6794);
nand U8791 (N_8791,N_7000,N_7338);
xnor U8792 (N_8792,N_7927,N_7994);
or U8793 (N_8793,N_7758,N_6230);
and U8794 (N_8794,N_6237,N_6416);
nor U8795 (N_8795,N_6984,N_6117);
nor U8796 (N_8796,N_6503,N_6583);
and U8797 (N_8797,N_6560,N_6387);
or U8798 (N_8798,N_7943,N_7314);
and U8799 (N_8799,N_7541,N_7518);
nand U8800 (N_8800,N_6890,N_6517);
xnor U8801 (N_8801,N_6994,N_7013);
or U8802 (N_8802,N_7852,N_6077);
and U8803 (N_8803,N_7130,N_7526);
nand U8804 (N_8804,N_7512,N_6580);
xor U8805 (N_8805,N_7445,N_7998);
nor U8806 (N_8806,N_7183,N_7950);
and U8807 (N_8807,N_7944,N_6036);
and U8808 (N_8808,N_6620,N_6856);
or U8809 (N_8809,N_6240,N_7694);
xnor U8810 (N_8810,N_6498,N_7647);
nand U8811 (N_8811,N_6908,N_7587);
xnor U8812 (N_8812,N_7384,N_6590);
and U8813 (N_8813,N_6957,N_6366);
xor U8814 (N_8814,N_7935,N_6442);
and U8815 (N_8815,N_6222,N_7207);
and U8816 (N_8816,N_7903,N_6609);
nor U8817 (N_8817,N_7754,N_6011);
xnor U8818 (N_8818,N_7695,N_6501);
nand U8819 (N_8819,N_6819,N_6970);
xnor U8820 (N_8820,N_6340,N_6733);
or U8821 (N_8821,N_6879,N_7287);
and U8822 (N_8822,N_7963,N_7262);
xor U8823 (N_8823,N_6210,N_6443);
nand U8824 (N_8824,N_6963,N_6260);
or U8825 (N_8825,N_6644,N_7387);
nor U8826 (N_8826,N_7894,N_7618);
and U8827 (N_8827,N_7200,N_6144);
or U8828 (N_8828,N_7120,N_6626);
and U8829 (N_8829,N_7653,N_7634);
nand U8830 (N_8830,N_6149,N_6303);
xor U8831 (N_8831,N_6234,N_6354);
xor U8832 (N_8832,N_6243,N_6298);
nor U8833 (N_8833,N_6972,N_6244);
or U8834 (N_8834,N_6302,N_7902);
xor U8835 (N_8835,N_6638,N_7219);
nor U8836 (N_8836,N_6634,N_6055);
xor U8837 (N_8837,N_6952,N_6943);
and U8838 (N_8838,N_7915,N_6071);
nand U8839 (N_8839,N_7070,N_7646);
nand U8840 (N_8840,N_7202,N_7600);
and U8841 (N_8841,N_6116,N_7276);
and U8842 (N_8842,N_7704,N_6519);
nand U8843 (N_8843,N_7132,N_6179);
nor U8844 (N_8844,N_7892,N_7059);
and U8845 (N_8845,N_6595,N_6067);
nand U8846 (N_8846,N_7056,N_7430);
or U8847 (N_8847,N_6716,N_6155);
xor U8848 (N_8848,N_6377,N_6341);
or U8849 (N_8849,N_6122,N_7350);
and U8850 (N_8850,N_6689,N_7795);
nor U8851 (N_8851,N_6840,N_6931);
and U8852 (N_8852,N_7047,N_7064);
and U8853 (N_8853,N_6969,N_7406);
or U8854 (N_8854,N_7215,N_6091);
xnor U8855 (N_8855,N_7741,N_7856);
nor U8856 (N_8856,N_6146,N_6352);
and U8857 (N_8857,N_6022,N_7577);
or U8858 (N_8858,N_7291,N_6089);
and U8859 (N_8859,N_7378,N_7578);
or U8860 (N_8860,N_7392,N_7412);
nor U8861 (N_8861,N_6719,N_6543);
xor U8862 (N_8862,N_7300,N_6136);
nand U8863 (N_8863,N_7352,N_6756);
xor U8864 (N_8864,N_7770,N_7210);
or U8865 (N_8865,N_6665,N_7748);
or U8866 (N_8866,N_7441,N_6006);
xnor U8867 (N_8867,N_7197,N_7460);
or U8868 (N_8868,N_6388,N_6863);
or U8869 (N_8869,N_6450,N_6675);
xor U8870 (N_8870,N_7566,N_6649);
nand U8871 (N_8871,N_6748,N_6438);
nor U8872 (N_8872,N_6065,N_7744);
nor U8873 (N_8873,N_6659,N_6955);
nand U8874 (N_8874,N_6339,N_7050);
nand U8875 (N_8875,N_7985,N_6673);
nor U8876 (N_8876,N_7746,N_7706);
or U8877 (N_8877,N_7595,N_6978);
nand U8878 (N_8878,N_7607,N_6841);
and U8879 (N_8879,N_6547,N_6008);
or U8880 (N_8880,N_6604,N_7716);
and U8881 (N_8881,N_6752,N_7565);
and U8882 (N_8882,N_7401,N_7847);
and U8883 (N_8883,N_6068,N_6289);
and U8884 (N_8884,N_6390,N_6402);
xor U8885 (N_8885,N_7525,N_7980);
and U8886 (N_8886,N_6860,N_7045);
and U8887 (N_8887,N_6500,N_6235);
xor U8888 (N_8888,N_6612,N_6798);
nor U8889 (N_8889,N_7527,N_6211);
xor U8890 (N_8890,N_7502,N_6780);
and U8891 (N_8891,N_6223,N_7645);
nand U8892 (N_8892,N_7071,N_6932);
and U8893 (N_8893,N_7363,N_6446);
nand U8894 (N_8894,N_7858,N_7355);
and U8895 (N_8895,N_7256,N_6225);
nor U8896 (N_8896,N_6864,N_7034);
and U8897 (N_8897,N_7385,N_6249);
or U8898 (N_8898,N_7832,N_7874);
and U8899 (N_8899,N_6486,N_7596);
and U8900 (N_8900,N_6137,N_7428);
xor U8901 (N_8901,N_7467,N_7671);
xor U8902 (N_8902,N_6191,N_7253);
and U8903 (N_8903,N_7410,N_6913);
and U8904 (N_8904,N_6961,N_6287);
xor U8905 (N_8905,N_6118,N_7018);
or U8906 (N_8906,N_7850,N_7376);
or U8907 (N_8907,N_7019,N_6814);
or U8908 (N_8908,N_6999,N_7679);
nand U8909 (N_8909,N_7005,N_7571);
xor U8910 (N_8910,N_6983,N_6641);
and U8911 (N_8911,N_7403,N_6018);
and U8912 (N_8912,N_7885,N_6278);
or U8913 (N_8913,N_6568,N_6391);
nor U8914 (N_8914,N_6892,N_6305);
and U8915 (N_8915,N_6455,N_6188);
xor U8916 (N_8916,N_6084,N_6064);
nor U8917 (N_8917,N_6148,N_7133);
nand U8918 (N_8918,N_7841,N_7601);
nor U8919 (N_8919,N_6050,N_7563);
nand U8920 (N_8920,N_6217,N_6114);
xor U8921 (N_8921,N_6028,N_6916);
and U8922 (N_8922,N_7966,N_6178);
or U8923 (N_8923,N_6139,N_7729);
and U8924 (N_8924,N_7891,N_7089);
and U8925 (N_8925,N_7789,N_7254);
xor U8926 (N_8926,N_6440,N_7886);
nor U8927 (N_8927,N_7438,N_7340);
nand U8928 (N_8928,N_6219,N_6605);
nand U8929 (N_8929,N_7660,N_7206);
and U8930 (N_8930,N_6817,N_7813);
nor U8931 (N_8931,N_6430,N_6746);
xor U8932 (N_8932,N_7683,N_7973);
nor U8933 (N_8933,N_7346,N_7913);
or U8934 (N_8934,N_6405,N_6229);
nand U8935 (N_8935,N_7959,N_7888);
nor U8936 (N_8936,N_7825,N_6744);
nor U8937 (N_8937,N_7672,N_6004);
or U8938 (N_8938,N_7542,N_7674);
and U8939 (N_8939,N_7996,N_7981);
xor U8940 (N_8940,N_6985,N_7918);
nand U8941 (N_8941,N_7531,N_7194);
nand U8942 (N_8942,N_6375,N_7157);
nor U8943 (N_8943,N_7265,N_6807);
and U8944 (N_8944,N_6226,N_6905);
xnor U8945 (N_8945,N_6342,N_7820);
or U8946 (N_8946,N_7091,N_7920);
or U8947 (N_8947,N_7549,N_6451);
xnor U8948 (N_8948,N_6330,N_7009);
xnor U8949 (N_8949,N_6200,N_6267);
nor U8950 (N_8950,N_7233,N_6529);
xnor U8951 (N_8951,N_6160,N_7127);
or U8952 (N_8952,N_6672,N_6875);
nor U8953 (N_8953,N_7879,N_6891);
nor U8954 (N_8954,N_6946,N_7055);
nand U8955 (N_8955,N_7511,N_7611);
nand U8956 (N_8956,N_6475,N_6877);
nor U8957 (N_8957,N_7831,N_7717);
or U8958 (N_8958,N_7507,N_7989);
nor U8959 (N_8959,N_6100,N_7170);
nand U8960 (N_8960,N_7986,N_6413);
nand U8961 (N_8961,N_6255,N_6835);
nand U8962 (N_8962,N_6850,N_7597);
nand U8963 (N_8963,N_6732,N_7336);
nand U8964 (N_8964,N_7272,N_7889);
nor U8965 (N_8965,N_6536,N_7728);
nand U8966 (N_8966,N_7500,N_7014);
and U8967 (N_8967,N_7869,N_7870);
nand U8968 (N_8968,N_6919,N_6456);
or U8969 (N_8969,N_6843,N_6192);
and U8970 (N_8970,N_7967,N_7244);
nand U8971 (N_8971,N_7105,N_7038);
xnor U8972 (N_8972,N_6159,N_7196);
nor U8973 (N_8973,N_6457,N_7872);
xnor U8974 (N_8974,N_7021,N_6582);
or U8975 (N_8975,N_7576,N_7074);
nand U8976 (N_8976,N_7642,N_7509);
or U8977 (N_8977,N_6271,N_7426);
nor U8978 (N_8978,N_6540,N_7582);
or U8979 (N_8979,N_7751,N_6212);
xor U8980 (N_8980,N_6886,N_7574);
nor U8981 (N_8981,N_6478,N_7037);
nor U8982 (N_8982,N_6607,N_7861);
nand U8983 (N_8983,N_7158,N_6633);
or U8984 (N_8984,N_6042,N_7462);
and U8985 (N_8985,N_6357,N_7979);
and U8986 (N_8986,N_6731,N_7490);
nor U8987 (N_8987,N_7875,N_7303);
or U8988 (N_8988,N_6806,N_7275);
nand U8989 (N_8989,N_7948,N_7878);
xnor U8990 (N_8990,N_7749,N_7805);
xor U8991 (N_8991,N_7489,N_6655);
and U8992 (N_8992,N_7742,N_6591);
and U8993 (N_8993,N_6668,N_6186);
xor U8994 (N_8994,N_6762,N_7007);
and U8995 (N_8995,N_6555,N_6196);
and U8996 (N_8996,N_6394,N_7842);
nand U8997 (N_8997,N_7190,N_7252);
and U8998 (N_8998,N_7223,N_6206);
xnor U8999 (N_8999,N_6700,N_7657);
xnor U9000 (N_9000,N_7592,N_7908);
xor U9001 (N_9001,N_7504,N_6433);
nand U9002 (N_9002,N_6085,N_6899);
nand U9003 (N_9003,N_6304,N_6727);
nand U9004 (N_9004,N_6032,N_6513);
nor U9005 (N_9005,N_7088,N_7403);
nor U9006 (N_9006,N_7737,N_7274);
nand U9007 (N_9007,N_6406,N_6046);
or U9008 (N_9008,N_7616,N_6109);
nor U9009 (N_9009,N_6300,N_7181);
nand U9010 (N_9010,N_6988,N_6476);
and U9011 (N_9011,N_7191,N_7812);
nand U9012 (N_9012,N_7571,N_7647);
and U9013 (N_9013,N_6273,N_6373);
and U9014 (N_9014,N_7768,N_6284);
nor U9015 (N_9015,N_7812,N_7124);
xnor U9016 (N_9016,N_7456,N_6103);
nor U9017 (N_9017,N_6858,N_7192);
and U9018 (N_9018,N_6294,N_6094);
nor U9019 (N_9019,N_6792,N_7287);
xor U9020 (N_9020,N_6414,N_6591);
nand U9021 (N_9021,N_7048,N_7785);
xor U9022 (N_9022,N_7873,N_6273);
xnor U9023 (N_9023,N_6282,N_6487);
nand U9024 (N_9024,N_7797,N_6925);
nand U9025 (N_9025,N_6656,N_7614);
or U9026 (N_9026,N_7275,N_7399);
nor U9027 (N_9027,N_6907,N_6532);
xnor U9028 (N_9028,N_7326,N_6882);
nor U9029 (N_9029,N_6356,N_6310);
or U9030 (N_9030,N_7287,N_6811);
xnor U9031 (N_9031,N_6199,N_6244);
xnor U9032 (N_9032,N_6542,N_7885);
and U9033 (N_9033,N_6069,N_6188);
nand U9034 (N_9034,N_6677,N_7373);
nand U9035 (N_9035,N_6466,N_6220);
nor U9036 (N_9036,N_6874,N_7420);
xnor U9037 (N_9037,N_7431,N_6707);
xor U9038 (N_9038,N_6787,N_7241);
or U9039 (N_9039,N_7813,N_6734);
and U9040 (N_9040,N_7157,N_7375);
nand U9041 (N_9041,N_6203,N_6808);
nand U9042 (N_9042,N_6191,N_7200);
nor U9043 (N_9043,N_6293,N_6360);
or U9044 (N_9044,N_7048,N_6749);
and U9045 (N_9045,N_6072,N_7999);
or U9046 (N_9046,N_7620,N_6207);
and U9047 (N_9047,N_6270,N_7801);
xnor U9048 (N_9048,N_6520,N_7719);
nor U9049 (N_9049,N_7908,N_6298);
nand U9050 (N_9050,N_6595,N_7276);
and U9051 (N_9051,N_7750,N_7385);
nand U9052 (N_9052,N_6770,N_6657);
xor U9053 (N_9053,N_7425,N_6164);
or U9054 (N_9054,N_7929,N_7592);
nor U9055 (N_9055,N_7966,N_6727);
and U9056 (N_9056,N_6981,N_6756);
xnor U9057 (N_9057,N_6949,N_7614);
nand U9058 (N_9058,N_7993,N_6607);
or U9059 (N_9059,N_6923,N_7671);
nand U9060 (N_9060,N_6567,N_7865);
or U9061 (N_9061,N_6136,N_6453);
or U9062 (N_9062,N_7945,N_6359);
nand U9063 (N_9063,N_7784,N_7989);
nor U9064 (N_9064,N_6241,N_7295);
xor U9065 (N_9065,N_7772,N_7662);
nand U9066 (N_9066,N_7423,N_6829);
and U9067 (N_9067,N_6290,N_7217);
and U9068 (N_9068,N_6129,N_7411);
xor U9069 (N_9069,N_7670,N_7441);
or U9070 (N_9070,N_6115,N_6459);
nand U9071 (N_9071,N_7575,N_6580);
nand U9072 (N_9072,N_6731,N_6660);
xnor U9073 (N_9073,N_6799,N_7323);
xor U9074 (N_9074,N_7429,N_7521);
xor U9075 (N_9075,N_6491,N_6157);
nor U9076 (N_9076,N_6430,N_7735);
nor U9077 (N_9077,N_7371,N_7524);
or U9078 (N_9078,N_6922,N_7442);
xnor U9079 (N_9079,N_7003,N_6853);
nand U9080 (N_9080,N_6703,N_7392);
nand U9081 (N_9081,N_7087,N_6985);
nand U9082 (N_9082,N_6355,N_7037);
nand U9083 (N_9083,N_6209,N_7236);
or U9084 (N_9084,N_6332,N_6280);
and U9085 (N_9085,N_6918,N_7086);
nor U9086 (N_9086,N_6962,N_6933);
nand U9087 (N_9087,N_7560,N_7796);
nand U9088 (N_9088,N_7136,N_6999);
and U9089 (N_9089,N_7108,N_6279);
or U9090 (N_9090,N_7191,N_6912);
or U9091 (N_9091,N_7948,N_7405);
nand U9092 (N_9092,N_7056,N_6833);
nor U9093 (N_9093,N_6333,N_6245);
nand U9094 (N_9094,N_6775,N_7560);
xor U9095 (N_9095,N_6920,N_6823);
and U9096 (N_9096,N_6281,N_6974);
xnor U9097 (N_9097,N_6255,N_6808);
nand U9098 (N_9098,N_7565,N_6185);
xnor U9099 (N_9099,N_6850,N_6322);
xor U9100 (N_9100,N_7535,N_7878);
nand U9101 (N_9101,N_6426,N_7158);
xnor U9102 (N_9102,N_6553,N_7926);
xnor U9103 (N_9103,N_7932,N_6612);
xor U9104 (N_9104,N_7412,N_6085);
nor U9105 (N_9105,N_7043,N_7692);
or U9106 (N_9106,N_6011,N_7400);
nor U9107 (N_9107,N_7006,N_6929);
and U9108 (N_9108,N_6029,N_6985);
or U9109 (N_9109,N_6234,N_6281);
nor U9110 (N_9110,N_6935,N_7781);
xor U9111 (N_9111,N_7337,N_7484);
nor U9112 (N_9112,N_7188,N_6812);
or U9113 (N_9113,N_6654,N_7846);
nor U9114 (N_9114,N_7083,N_6589);
or U9115 (N_9115,N_7621,N_6588);
xor U9116 (N_9116,N_6781,N_7799);
nand U9117 (N_9117,N_7810,N_7286);
or U9118 (N_9118,N_6365,N_6334);
xor U9119 (N_9119,N_6913,N_7842);
and U9120 (N_9120,N_7746,N_6020);
xor U9121 (N_9121,N_7720,N_6791);
nor U9122 (N_9122,N_7113,N_6400);
and U9123 (N_9123,N_6188,N_7515);
nor U9124 (N_9124,N_6229,N_6944);
nand U9125 (N_9125,N_6802,N_7803);
nor U9126 (N_9126,N_7630,N_7311);
nand U9127 (N_9127,N_7143,N_7640);
nand U9128 (N_9128,N_7376,N_7554);
and U9129 (N_9129,N_7025,N_7077);
and U9130 (N_9130,N_6453,N_7768);
nor U9131 (N_9131,N_7068,N_6513);
xor U9132 (N_9132,N_7323,N_6033);
xnor U9133 (N_9133,N_7927,N_7946);
or U9134 (N_9134,N_6068,N_6911);
nor U9135 (N_9135,N_6645,N_6579);
nor U9136 (N_9136,N_7103,N_7987);
and U9137 (N_9137,N_7835,N_6597);
nor U9138 (N_9138,N_6801,N_6034);
nand U9139 (N_9139,N_7957,N_7570);
and U9140 (N_9140,N_7036,N_7982);
nand U9141 (N_9141,N_6546,N_7225);
nor U9142 (N_9142,N_7794,N_7805);
and U9143 (N_9143,N_6049,N_6593);
and U9144 (N_9144,N_7458,N_6074);
and U9145 (N_9145,N_7300,N_6749);
nor U9146 (N_9146,N_7759,N_6420);
nand U9147 (N_9147,N_6977,N_7843);
nor U9148 (N_9148,N_6577,N_7536);
xnor U9149 (N_9149,N_6666,N_7247);
nor U9150 (N_9150,N_7292,N_6012);
and U9151 (N_9151,N_6546,N_6785);
or U9152 (N_9152,N_7150,N_6587);
nand U9153 (N_9153,N_6327,N_7609);
and U9154 (N_9154,N_6138,N_7137);
nor U9155 (N_9155,N_6465,N_7678);
and U9156 (N_9156,N_7865,N_7728);
nand U9157 (N_9157,N_6402,N_6910);
xor U9158 (N_9158,N_7803,N_6460);
nor U9159 (N_9159,N_6303,N_6420);
or U9160 (N_9160,N_7737,N_7119);
xnor U9161 (N_9161,N_7391,N_6044);
nor U9162 (N_9162,N_7970,N_7779);
nor U9163 (N_9163,N_6593,N_7731);
nor U9164 (N_9164,N_7183,N_7748);
xnor U9165 (N_9165,N_7805,N_6613);
xnor U9166 (N_9166,N_6146,N_6963);
xnor U9167 (N_9167,N_7732,N_6887);
xor U9168 (N_9168,N_7529,N_6071);
nor U9169 (N_9169,N_6477,N_6149);
nand U9170 (N_9170,N_6215,N_6286);
and U9171 (N_9171,N_7974,N_6037);
and U9172 (N_9172,N_7019,N_7567);
or U9173 (N_9173,N_7402,N_7522);
and U9174 (N_9174,N_7169,N_6080);
nor U9175 (N_9175,N_6554,N_6523);
nor U9176 (N_9176,N_6089,N_7672);
or U9177 (N_9177,N_7650,N_6826);
nand U9178 (N_9178,N_7076,N_7017);
and U9179 (N_9179,N_7444,N_6651);
xor U9180 (N_9180,N_7147,N_6435);
and U9181 (N_9181,N_6943,N_6638);
xnor U9182 (N_9182,N_7910,N_6752);
or U9183 (N_9183,N_6302,N_6267);
nor U9184 (N_9184,N_6396,N_7756);
nand U9185 (N_9185,N_6217,N_6739);
xor U9186 (N_9186,N_7954,N_6845);
nor U9187 (N_9187,N_6454,N_7326);
xnor U9188 (N_9188,N_7171,N_7588);
and U9189 (N_9189,N_7611,N_7381);
xnor U9190 (N_9190,N_7021,N_6604);
nor U9191 (N_9191,N_7942,N_6384);
nand U9192 (N_9192,N_7423,N_6440);
nor U9193 (N_9193,N_7516,N_7571);
nand U9194 (N_9194,N_6961,N_6519);
and U9195 (N_9195,N_7671,N_7746);
or U9196 (N_9196,N_7608,N_7389);
or U9197 (N_9197,N_7028,N_6828);
nand U9198 (N_9198,N_7392,N_6871);
xnor U9199 (N_9199,N_6154,N_6640);
or U9200 (N_9200,N_6251,N_6421);
or U9201 (N_9201,N_6063,N_6622);
nor U9202 (N_9202,N_6342,N_6977);
xnor U9203 (N_9203,N_6914,N_7832);
xnor U9204 (N_9204,N_7141,N_6080);
nor U9205 (N_9205,N_6804,N_7837);
and U9206 (N_9206,N_7383,N_6529);
nor U9207 (N_9207,N_6960,N_6422);
or U9208 (N_9208,N_7702,N_7650);
nor U9209 (N_9209,N_7307,N_6145);
and U9210 (N_9210,N_7649,N_6981);
or U9211 (N_9211,N_6870,N_6214);
nor U9212 (N_9212,N_6203,N_6834);
xor U9213 (N_9213,N_7858,N_6112);
xor U9214 (N_9214,N_6598,N_6684);
and U9215 (N_9215,N_6820,N_6886);
nor U9216 (N_9216,N_6021,N_7581);
or U9217 (N_9217,N_6361,N_6208);
or U9218 (N_9218,N_6448,N_6882);
or U9219 (N_9219,N_7817,N_7746);
nor U9220 (N_9220,N_7427,N_7108);
nand U9221 (N_9221,N_6319,N_7568);
and U9222 (N_9222,N_7969,N_7824);
and U9223 (N_9223,N_7628,N_6682);
and U9224 (N_9224,N_7831,N_7395);
and U9225 (N_9225,N_7169,N_7864);
or U9226 (N_9226,N_6813,N_6717);
nand U9227 (N_9227,N_6860,N_6889);
or U9228 (N_9228,N_7788,N_6590);
nand U9229 (N_9229,N_7612,N_6227);
nor U9230 (N_9230,N_7708,N_7413);
xnor U9231 (N_9231,N_7287,N_6087);
or U9232 (N_9232,N_7224,N_6827);
or U9233 (N_9233,N_6983,N_7661);
nor U9234 (N_9234,N_6202,N_7558);
xor U9235 (N_9235,N_6755,N_6509);
and U9236 (N_9236,N_6776,N_6578);
or U9237 (N_9237,N_7159,N_7337);
nor U9238 (N_9238,N_7585,N_6444);
and U9239 (N_9239,N_7738,N_6439);
nand U9240 (N_9240,N_6891,N_7564);
nor U9241 (N_9241,N_7341,N_6283);
nand U9242 (N_9242,N_7573,N_7713);
and U9243 (N_9243,N_7002,N_7890);
xor U9244 (N_9244,N_7704,N_6778);
xor U9245 (N_9245,N_6222,N_7460);
and U9246 (N_9246,N_6391,N_6907);
and U9247 (N_9247,N_6544,N_7294);
xnor U9248 (N_9248,N_7130,N_6186);
xnor U9249 (N_9249,N_7486,N_7586);
and U9250 (N_9250,N_7531,N_6784);
or U9251 (N_9251,N_6215,N_6316);
and U9252 (N_9252,N_6347,N_6490);
xnor U9253 (N_9253,N_6869,N_7525);
or U9254 (N_9254,N_6047,N_6348);
nand U9255 (N_9255,N_6210,N_7877);
and U9256 (N_9256,N_6678,N_6270);
nand U9257 (N_9257,N_6904,N_7272);
nand U9258 (N_9258,N_6272,N_6004);
nor U9259 (N_9259,N_6608,N_7417);
and U9260 (N_9260,N_7858,N_6092);
or U9261 (N_9261,N_6145,N_6933);
and U9262 (N_9262,N_7836,N_6544);
nor U9263 (N_9263,N_6173,N_6103);
and U9264 (N_9264,N_7892,N_6646);
xnor U9265 (N_9265,N_7693,N_7208);
or U9266 (N_9266,N_6216,N_7533);
xor U9267 (N_9267,N_7925,N_7728);
and U9268 (N_9268,N_6153,N_7492);
nor U9269 (N_9269,N_7307,N_6035);
nand U9270 (N_9270,N_7405,N_7560);
nor U9271 (N_9271,N_6350,N_6472);
or U9272 (N_9272,N_6775,N_7572);
nand U9273 (N_9273,N_6959,N_6882);
nand U9274 (N_9274,N_6523,N_7931);
xor U9275 (N_9275,N_6271,N_7870);
nor U9276 (N_9276,N_6746,N_7286);
or U9277 (N_9277,N_7791,N_7502);
and U9278 (N_9278,N_7302,N_6224);
nor U9279 (N_9279,N_7378,N_7167);
nor U9280 (N_9280,N_6576,N_7560);
and U9281 (N_9281,N_7805,N_7556);
and U9282 (N_9282,N_7757,N_6415);
nor U9283 (N_9283,N_7134,N_7012);
nand U9284 (N_9284,N_7193,N_7458);
xor U9285 (N_9285,N_7122,N_7599);
xor U9286 (N_9286,N_6525,N_6902);
xnor U9287 (N_9287,N_7705,N_7799);
nand U9288 (N_9288,N_7734,N_7953);
xor U9289 (N_9289,N_6937,N_6721);
nand U9290 (N_9290,N_6800,N_7118);
xnor U9291 (N_9291,N_7273,N_7056);
or U9292 (N_9292,N_7080,N_7414);
and U9293 (N_9293,N_6341,N_6135);
or U9294 (N_9294,N_6227,N_6148);
nor U9295 (N_9295,N_6363,N_7969);
nor U9296 (N_9296,N_6485,N_6120);
xor U9297 (N_9297,N_6859,N_7993);
nand U9298 (N_9298,N_6936,N_7251);
and U9299 (N_9299,N_7419,N_6122);
and U9300 (N_9300,N_7934,N_6624);
and U9301 (N_9301,N_6030,N_6261);
or U9302 (N_9302,N_7861,N_6284);
and U9303 (N_9303,N_6991,N_6378);
and U9304 (N_9304,N_6442,N_6646);
nand U9305 (N_9305,N_7393,N_6978);
nor U9306 (N_9306,N_7918,N_6009);
xor U9307 (N_9307,N_6123,N_6175);
or U9308 (N_9308,N_6951,N_6740);
xor U9309 (N_9309,N_6861,N_6458);
nand U9310 (N_9310,N_7006,N_7618);
nand U9311 (N_9311,N_6236,N_6866);
nand U9312 (N_9312,N_6429,N_7397);
and U9313 (N_9313,N_6898,N_6358);
xnor U9314 (N_9314,N_6324,N_7138);
or U9315 (N_9315,N_7493,N_6196);
xor U9316 (N_9316,N_6470,N_7931);
and U9317 (N_9317,N_7606,N_6954);
nand U9318 (N_9318,N_6845,N_7762);
nand U9319 (N_9319,N_6399,N_6872);
nor U9320 (N_9320,N_7685,N_7890);
or U9321 (N_9321,N_7983,N_7735);
and U9322 (N_9322,N_7530,N_6881);
nand U9323 (N_9323,N_6877,N_7496);
nor U9324 (N_9324,N_6088,N_7944);
and U9325 (N_9325,N_6932,N_6446);
and U9326 (N_9326,N_7142,N_7612);
xor U9327 (N_9327,N_6021,N_6653);
nor U9328 (N_9328,N_6352,N_6522);
and U9329 (N_9329,N_7778,N_6255);
or U9330 (N_9330,N_6816,N_7657);
or U9331 (N_9331,N_6914,N_7483);
or U9332 (N_9332,N_7267,N_6969);
and U9333 (N_9333,N_6573,N_6642);
nor U9334 (N_9334,N_7718,N_6825);
xnor U9335 (N_9335,N_6189,N_6810);
nor U9336 (N_9336,N_6149,N_7720);
and U9337 (N_9337,N_7532,N_6127);
nand U9338 (N_9338,N_7806,N_7246);
and U9339 (N_9339,N_6442,N_6616);
nand U9340 (N_9340,N_6791,N_6627);
nor U9341 (N_9341,N_7620,N_7109);
xor U9342 (N_9342,N_6144,N_6070);
xor U9343 (N_9343,N_7564,N_6319);
or U9344 (N_9344,N_7214,N_6461);
xnor U9345 (N_9345,N_6761,N_7347);
or U9346 (N_9346,N_6005,N_7105);
nor U9347 (N_9347,N_7703,N_7638);
and U9348 (N_9348,N_7041,N_7858);
and U9349 (N_9349,N_6388,N_7078);
nor U9350 (N_9350,N_6779,N_7725);
nand U9351 (N_9351,N_7624,N_7311);
xor U9352 (N_9352,N_6679,N_6238);
xnor U9353 (N_9353,N_6290,N_6554);
nor U9354 (N_9354,N_7024,N_6956);
xor U9355 (N_9355,N_7937,N_6623);
nor U9356 (N_9356,N_7876,N_6625);
and U9357 (N_9357,N_7308,N_7029);
nor U9358 (N_9358,N_7014,N_7523);
xor U9359 (N_9359,N_7163,N_7049);
xnor U9360 (N_9360,N_7882,N_6794);
nand U9361 (N_9361,N_7452,N_7303);
nor U9362 (N_9362,N_7111,N_7602);
nand U9363 (N_9363,N_7923,N_6022);
and U9364 (N_9364,N_6351,N_7947);
and U9365 (N_9365,N_6207,N_6894);
xnor U9366 (N_9366,N_7537,N_7351);
nand U9367 (N_9367,N_7819,N_6356);
and U9368 (N_9368,N_7195,N_7282);
or U9369 (N_9369,N_7257,N_6727);
nor U9370 (N_9370,N_6175,N_6941);
and U9371 (N_9371,N_7819,N_6648);
xor U9372 (N_9372,N_6218,N_6990);
or U9373 (N_9373,N_6139,N_7641);
xor U9374 (N_9374,N_6983,N_6049);
or U9375 (N_9375,N_6393,N_6908);
and U9376 (N_9376,N_7782,N_7264);
and U9377 (N_9377,N_7546,N_7829);
nand U9378 (N_9378,N_6226,N_7480);
nand U9379 (N_9379,N_7020,N_7035);
and U9380 (N_9380,N_6101,N_6462);
and U9381 (N_9381,N_7341,N_6291);
and U9382 (N_9382,N_7479,N_6135);
nor U9383 (N_9383,N_6674,N_7411);
nor U9384 (N_9384,N_7687,N_7834);
or U9385 (N_9385,N_6652,N_6705);
and U9386 (N_9386,N_6778,N_6820);
nor U9387 (N_9387,N_7777,N_6415);
nand U9388 (N_9388,N_7587,N_6992);
nor U9389 (N_9389,N_6726,N_7905);
and U9390 (N_9390,N_7506,N_6882);
xor U9391 (N_9391,N_7041,N_7488);
xnor U9392 (N_9392,N_6179,N_6414);
nor U9393 (N_9393,N_7011,N_6565);
nor U9394 (N_9394,N_7282,N_6450);
nand U9395 (N_9395,N_6926,N_7925);
xnor U9396 (N_9396,N_7917,N_7074);
or U9397 (N_9397,N_7276,N_6553);
nor U9398 (N_9398,N_6544,N_6903);
nor U9399 (N_9399,N_7145,N_7837);
and U9400 (N_9400,N_6240,N_7461);
or U9401 (N_9401,N_6607,N_7670);
nor U9402 (N_9402,N_6896,N_6259);
nor U9403 (N_9403,N_6477,N_7915);
nand U9404 (N_9404,N_7518,N_7020);
xor U9405 (N_9405,N_6223,N_7832);
nor U9406 (N_9406,N_6018,N_7726);
and U9407 (N_9407,N_7918,N_6311);
and U9408 (N_9408,N_6851,N_7291);
nand U9409 (N_9409,N_7504,N_7587);
or U9410 (N_9410,N_6721,N_7880);
xor U9411 (N_9411,N_6144,N_6800);
and U9412 (N_9412,N_7574,N_6985);
nand U9413 (N_9413,N_6031,N_6105);
nand U9414 (N_9414,N_6026,N_6746);
nand U9415 (N_9415,N_7492,N_6108);
or U9416 (N_9416,N_6753,N_7650);
nand U9417 (N_9417,N_6192,N_6520);
xor U9418 (N_9418,N_6191,N_7436);
xnor U9419 (N_9419,N_6474,N_7527);
nor U9420 (N_9420,N_6313,N_7715);
xor U9421 (N_9421,N_7396,N_7597);
and U9422 (N_9422,N_6021,N_7711);
or U9423 (N_9423,N_6909,N_7799);
or U9424 (N_9424,N_7626,N_7812);
and U9425 (N_9425,N_6965,N_6265);
xnor U9426 (N_9426,N_6085,N_7658);
nor U9427 (N_9427,N_7914,N_6242);
nand U9428 (N_9428,N_7246,N_6793);
xnor U9429 (N_9429,N_7914,N_7608);
and U9430 (N_9430,N_7265,N_7191);
nor U9431 (N_9431,N_6476,N_7592);
xor U9432 (N_9432,N_7016,N_7336);
or U9433 (N_9433,N_6628,N_6188);
nand U9434 (N_9434,N_7349,N_6511);
nor U9435 (N_9435,N_6060,N_6501);
or U9436 (N_9436,N_6276,N_7813);
or U9437 (N_9437,N_7708,N_7117);
or U9438 (N_9438,N_7539,N_6683);
nor U9439 (N_9439,N_6776,N_6891);
or U9440 (N_9440,N_6965,N_7631);
and U9441 (N_9441,N_6202,N_6682);
and U9442 (N_9442,N_7145,N_6721);
xnor U9443 (N_9443,N_7381,N_7983);
nand U9444 (N_9444,N_7533,N_6751);
and U9445 (N_9445,N_7213,N_6440);
xnor U9446 (N_9446,N_6161,N_7735);
nor U9447 (N_9447,N_6038,N_6495);
nand U9448 (N_9448,N_7860,N_6104);
and U9449 (N_9449,N_7014,N_6955);
nor U9450 (N_9450,N_6066,N_6609);
or U9451 (N_9451,N_7913,N_6011);
or U9452 (N_9452,N_7993,N_6083);
nor U9453 (N_9453,N_7633,N_7573);
nor U9454 (N_9454,N_7803,N_6536);
nand U9455 (N_9455,N_6441,N_7068);
xor U9456 (N_9456,N_7313,N_6559);
nand U9457 (N_9457,N_7000,N_6157);
or U9458 (N_9458,N_7237,N_6041);
and U9459 (N_9459,N_6287,N_6557);
nand U9460 (N_9460,N_6985,N_7838);
nor U9461 (N_9461,N_7945,N_6747);
nor U9462 (N_9462,N_7280,N_6302);
and U9463 (N_9463,N_6339,N_6327);
nor U9464 (N_9464,N_7881,N_6556);
nand U9465 (N_9465,N_6730,N_6408);
or U9466 (N_9466,N_6600,N_7959);
nor U9467 (N_9467,N_6182,N_6599);
or U9468 (N_9468,N_7224,N_7510);
or U9469 (N_9469,N_6174,N_6932);
nand U9470 (N_9470,N_7942,N_7423);
xnor U9471 (N_9471,N_6930,N_7994);
and U9472 (N_9472,N_6800,N_6719);
or U9473 (N_9473,N_6272,N_7129);
and U9474 (N_9474,N_7833,N_7287);
nand U9475 (N_9475,N_6685,N_6143);
nor U9476 (N_9476,N_6943,N_6178);
or U9477 (N_9477,N_6083,N_6509);
xor U9478 (N_9478,N_6981,N_6757);
xnor U9479 (N_9479,N_7851,N_6146);
nor U9480 (N_9480,N_6846,N_6239);
or U9481 (N_9481,N_6815,N_7158);
xnor U9482 (N_9482,N_6746,N_6290);
nor U9483 (N_9483,N_7398,N_7351);
nor U9484 (N_9484,N_6070,N_7660);
xnor U9485 (N_9485,N_7587,N_6431);
xor U9486 (N_9486,N_7015,N_7710);
and U9487 (N_9487,N_6861,N_6653);
and U9488 (N_9488,N_6692,N_7776);
and U9489 (N_9489,N_7526,N_6728);
and U9490 (N_9490,N_6839,N_6440);
nand U9491 (N_9491,N_6160,N_7529);
nor U9492 (N_9492,N_7760,N_6515);
nand U9493 (N_9493,N_7315,N_6924);
nand U9494 (N_9494,N_6584,N_6523);
nand U9495 (N_9495,N_6271,N_6652);
and U9496 (N_9496,N_7384,N_7967);
and U9497 (N_9497,N_7813,N_6881);
or U9498 (N_9498,N_7997,N_7303);
and U9499 (N_9499,N_6903,N_7270);
nor U9500 (N_9500,N_7742,N_7723);
nand U9501 (N_9501,N_7419,N_7811);
xnor U9502 (N_9502,N_6935,N_7105);
or U9503 (N_9503,N_6465,N_6986);
nor U9504 (N_9504,N_6182,N_7950);
and U9505 (N_9505,N_6475,N_6372);
or U9506 (N_9506,N_7766,N_7108);
xor U9507 (N_9507,N_7944,N_7590);
or U9508 (N_9508,N_7184,N_6604);
or U9509 (N_9509,N_6649,N_6311);
nor U9510 (N_9510,N_6913,N_6355);
nor U9511 (N_9511,N_6934,N_6095);
nor U9512 (N_9512,N_7085,N_6241);
and U9513 (N_9513,N_7953,N_6326);
nand U9514 (N_9514,N_6210,N_7261);
nor U9515 (N_9515,N_6581,N_7281);
nand U9516 (N_9516,N_6312,N_6718);
nor U9517 (N_9517,N_7983,N_6248);
or U9518 (N_9518,N_7670,N_7472);
or U9519 (N_9519,N_6680,N_6466);
or U9520 (N_9520,N_6177,N_7489);
xnor U9521 (N_9521,N_6911,N_6250);
nor U9522 (N_9522,N_6596,N_6906);
and U9523 (N_9523,N_6190,N_7352);
xnor U9524 (N_9524,N_7906,N_7521);
nand U9525 (N_9525,N_7034,N_7506);
xnor U9526 (N_9526,N_6384,N_6401);
nand U9527 (N_9527,N_7066,N_6190);
and U9528 (N_9528,N_6715,N_6447);
or U9529 (N_9529,N_6018,N_7678);
nor U9530 (N_9530,N_7169,N_7609);
and U9531 (N_9531,N_7867,N_7545);
and U9532 (N_9532,N_6533,N_6914);
xnor U9533 (N_9533,N_7786,N_7673);
and U9534 (N_9534,N_7926,N_7199);
and U9535 (N_9535,N_6276,N_7206);
and U9536 (N_9536,N_6261,N_6530);
and U9537 (N_9537,N_6141,N_6107);
and U9538 (N_9538,N_7632,N_6561);
xnor U9539 (N_9539,N_6236,N_6098);
nand U9540 (N_9540,N_6453,N_6248);
nand U9541 (N_9541,N_6521,N_7313);
and U9542 (N_9542,N_7586,N_6718);
nand U9543 (N_9543,N_7316,N_7597);
and U9544 (N_9544,N_6957,N_7626);
and U9545 (N_9545,N_6158,N_6341);
and U9546 (N_9546,N_6007,N_7836);
nor U9547 (N_9547,N_6681,N_6110);
or U9548 (N_9548,N_6870,N_6968);
or U9549 (N_9549,N_7816,N_6807);
xor U9550 (N_9550,N_7885,N_7206);
nand U9551 (N_9551,N_7416,N_7850);
or U9552 (N_9552,N_7972,N_6850);
and U9553 (N_9553,N_6687,N_7441);
nor U9554 (N_9554,N_7551,N_6167);
nand U9555 (N_9555,N_6660,N_6144);
and U9556 (N_9556,N_7968,N_7944);
nor U9557 (N_9557,N_6233,N_7304);
nor U9558 (N_9558,N_7833,N_6241);
nor U9559 (N_9559,N_7836,N_6651);
nor U9560 (N_9560,N_6428,N_7462);
nand U9561 (N_9561,N_7099,N_7671);
nor U9562 (N_9562,N_7947,N_6622);
and U9563 (N_9563,N_7587,N_7793);
or U9564 (N_9564,N_6660,N_6048);
nand U9565 (N_9565,N_7813,N_6638);
nor U9566 (N_9566,N_6039,N_7125);
or U9567 (N_9567,N_6856,N_7826);
and U9568 (N_9568,N_6009,N_6142);
nand U9569 (N_9569,N_6662,N_7283);
or U9570 (N_9570,N_7000,N_7640);
or U9571 (N_9571,N_7106,N_6564);
nor U9572 (N_9572,N_6730,N_7521);
or U9573 (N_9573,N_7514,N_7511);
nor U9574 (N_9574,N_7154,N_6351);
and U9575 (N_9575,N_7468,N_6918);
xnor U9576 (N_9576,N_6565,N_7005);
xor U9577 (N_9577,N_7409,N_6625);
nor U9578 (N_9578,N_6820,N_7621);
nor U9579 (N_9579,N_6727,N_7790);
or U9580 (N_9580,N_7822,N_7470);
and U9581 (N_9581,N_6125,N_6037);
xnor U9582 (N_9582,N_6380,N_6341);
nor U9583 (N_9583,N_6452,N_7973);
and U9584 (N_9584,N_6042,N_6869);
nor U9585 (N_9585,N_6557,N_6122);
nor U9586 (N_9586,N_6548,N_6609);
and U9587 (N_9587,N_7162,N_7322);
nor U9588 (N_9588,N_6029,N_6754);
and U9589 (N_9589,N_7370,N_7646);
or U9590 (N_9590,N_6712,N_6280);
and U9591 (N_9591,N_7119,N_6144);
and U9592 (N_9592,N_6932,N_7222);
xor U9593 (N_9593,N_6894,N_6242);
nor U9594 (N_9594,N_7102,N_7551);
and U9595 (N_9595,N_6807,N_6073);
or U9596 (N_9596,N_7857,N_6192);
xnor U9597 (N_9597,N_7873,N_7252);
nor U9598 (N_9598,N_7951,N_7338);
nand U9599 (N_9599,N_6716,N_7193);
nand U9600 (N_9600,N_6056,N_7164);
or U9601 (N_9601,N_7648,N_6360);
nand U9602 (N_9602,N_6281,N_7082);
or U9603 (N_9603,N_7431,N_6896);
xor U9604 (N_9604,N_7157,N_7042);
xnor U9605 (N_9605,N_6261,N_7573);
nand U9606 (N_9606,N_7307,N_6944);
or U9607 (N_9607,N_7299,N_7500);
nand U9608 (N_9608,N_6884,N_6920);
nor U9609 (N_9609,N_7817,N_6872);
xnor U9610 (N_9610,N_6946,N_6336);
or U9611 (N_9611,N_6690,N_6864);
and U9612 (N_9612,N_7191,N_7827);
or U9613 (N_9613,N_7125,N_6311);
nand U9614 (N_9614,N_6415,N_7554);
nand U9615 (N_9615,N_7608,N_7106);
nor U9616 (N_9616,N_6679,N_6242);
and U9617 (N_9617,N_6566,N_6076);
and U9618 (N_9618,N_7057,N_7894);
and U9619 (N_9619,N_6811,N_6836);
xnor U9620 (N_9620,N_7836,N_7998);
and U9621 (N_9621,N_6890,N_6322);
nand U9622 (N_9622,N_7261,N_7021);
nor U9623 (N_9623,N_6442,N_7274);
or U9624 (N_9624,N_6813,N_6982);
and U9625 (N_9625,N_6203,N_7047);
xnor U9626 (N_9626,N_7532,N_6990);
nand U9627 (N_9627,N_7628,N_6522);
nand U9628 (N_9628,N_7476,N_6999);
xor U9629 (N_9629,N_7176,N_7916);
nor U9630 (N_9630,N_7582,N_7493);
or U9631 (N_9631,N_6544,N_6510);
xnor U9632 (N_9632,N_6724,N_6859);
nor U9633 (N_9633,N_7678,N_7346);
or U9634 (N_9634,N_7140,N_6269);
xor U9635 (N_9635,N_6174,N_7707);
or U9636 (N_9636,N_7703,N_6013);
xnor U9637 (N_9637,N_7927,N_7366);
nand U9638 (N_9638,N_6890,N_6707);
and U9639 (N_9639,N_7836,N_6746);
or U9640 (N_9640,N_7180,N_7615);
nor U9641 (N_9641,N_6628,N_7149);
and U9642 (N_9642,N_7154,N_7227);
nand U9643 (N_9643,N_6655,N_6913);
or U9644 (N_9644,N_6729,N_7493);
xor U9645 (N_9645,N_7277,N_7958);
nand U9646 (N_9646,N_7111,N_7878);
nor U9647 (N_9647,N_7948,N_7197);
or U9648 (N_9648,N_6691,N_7538);
xor U9649 (N_9649,N_7001,N_6145);
and U9650 (N_9650,N_7190,N_7211);
and U9651 (N_9651,N_7493,N_7388);
nor U9652 (N_9652,N_7508,N_6686);
nand U9653 (N_9653,N_7835,N_6187);
or U9654 (N_9654,N_6256,N_7575);
nand U9655 (N_9655,N_6162,N_6255);
and U9656 (N_9656,N_7414,N_7802);
nand U9657 (N_9657,N_7281,N_7565);
or U9658 (N_9658,N_6004,N_6485);
and U9659 (N_9659,N_7919,N_6991);
xor U9660 (N_9660,N_7203,N_7940);
xor U9661 (N_9661,N_6519,N_6540);
xor U9662 (N_9662,N_7834,N_6754);
nand U9663 (N_9663,N_7085,N_7469);
and U9664 (N_9664,N_6139,N_7448);
nand U9665 (N_9665,N_7606,N_6541);
and U9666 (N_9666,N_6747,N_7152);
xnor U9667 (N_9667,N_7068,N_6095);
and U9668 (N_9668,N_6811,N_7066);
or U9669 (N_9669,N_7093,N_7272);
nor U9670 (N_9670,N_6052,N_7813);
nand U9671 (N_9671,N_7341,N_6932);
and U9672 (N_9672,N_7648,N_7518);
and U9673 (N_9673,N_7315,N_7430);
nor U9674 (N_9674,N_6167,N_6915);
nor U9675 (N_9675,N_6477,N_6892);
or U9676 (N_9676,N_6571,N_7818);
xor U9677 (N_9677,N_7929,N_6985);
xor U9678 (N_9678,N_6379,N_6443);
or U9679 (N_9679,N_7779,N_6771);
xor U9680 (N_9680,N_7324,N_6778);
or U9681 (N_9681,N_6204,N_7132);
nor U9682 (N_9682,N_7846,N_6764);
nor U9683 (N_9683,N_6692,N_7345);
or U9684 (N_9684,N_7568,N_7266);
xnor U9685 (N_9685,N_6587,N_6756);
xnor U9686 (N_9686,N_7467,N_6635);
nor U9687 (N_9687,N_6715,N_6051);
nand U9688 (N_9688,N_6041,N_6264);
or U9689 (N_9689,N_6958,N_6478);
nand U9690 (N_9690,N_7934,N_7440);
nand U9691 (N_9691,N_6491,N_6830);
and U9692 (N_9692,N_7932,N_7424);
xor U9693 (N_9693,N_7820,N_6232);
or U9694 (N_9694,N_6488,N_7457);
and U9695 (N_9695,N_6306,N_7948);
nor U9696 (N_9696,N_6419,N_7227);
and U9697 (N_9697,N_7068,N_6255);
nand U9698 (N_9698,N_6450,N_7368);
and U9699 (N_9699,N_6436,N_7283);
and U9700 (N_9700,N_7966,N_7559);
xnor U9701 (N_9701,N_7091,N_6929);
or U9702 (N_9702,N_6666,N_6670);
nor U9703 (N_9703,N_7478,N_6773);
nor U9704 (N_9704,N_6974,N_7014);
nor U9705 (N_9705,N_7568,N_7168);
nor U9706 (N_9706,N_7112,N_6454);
nor U9707 (N_9707,N_7374,N_7814);
xnor U9708 (N_9708,N_7514,N_6358);
and U9709 (N_9709,N_6575,N_7878);
xor U9710 (N_9710,N_6032,N_6728);
nor U9711 (N_9711,N_6099,N_7661);
nor U9712 (N_9712,N_7005,N_7454);
or U9713 (N_9713,N_7745,N_7111);
and U9714 (N_9714,N_6514,N_7477);
or U9715 (N_9715,N_6597,N_6793);
nand U9716 (N_9716,N_6400,N_6558);
nor U9717 (N_9717,N_7115,N_7249);
nor U9718 (N_9718,N_6689,N_7784);
nor U9719 (N_9719,N_7009,N_6745);
nand U9720 (N_9720,N_6016,N_6715);
and U9721 (N_9721,N_7845,N_6763);
and U9722 (N_9722,N_6107,N_7540);
or U9723 (N_9723,N_6966,N_6797);
and U9724 (N_9724,N_7049,N_6610);
xor U9725 (N_9725,N_7911,N_7243);
and U9726 (N_9726,N_7714,N_6685);
or U9727 (N_9727,N_7015,N_6788);
xor U9728 (N_9728,N_7184,N_7055);
xor U9729 (N_9729,N_6899,N_6494);
or U9730 (N_9730,N_7470,N_6095);
or U9731 (N_9731,N_6424,N_7986);
xor U9732 (N_9732,N_6526,N_6854);
and U9733 (N_9733,N_6653,N_7514);
xor U9734 (N_9734,N_6862,N_6857);
nor U9735 (N_9735,N_7990,N_6544);
nor U9736 (N_9736,N_6079,N_7837);
and U9737 (N_9737,N_7026,N_7077);
and U9738 (N_9738,N_6201,N_6138);
xnor U9739 (N_9739,N_6429,N_6062);
nor U9740 (N_9740,N_6113,N_7780);
and U9741 (N_9741,N_6627,N_6343);
or U9742 (N_9742,N_7814,N_7644);
or U9743 (N_9743,N_7995,N_7371);
or U9744 (N_9744,N_7957,N_6180);
xnor U9745 (N_9745,N_7288,N_6418);
nand U9746 (N_9746,N_7683,N_6600);
nand U9747 (N_9747,N_6951,N_6222);
nor U9748 (N_9748,N_6835,N_6659);
nor U9749 (N_9749,N_6866,N_6266);
xor U9750 (N_9750,N_7532,N_6691);
nand U9751 (N_9751,N_7626,N_7795);
and U9752 (N_9752,N_7249,N_6380);
nor U9753 (N_9753,N_6108,N_7113);
xnor U9754 (N_9754,N_6742,N_7854);
xnor U9755 (N_9755,N_6275,N_6786);
and U9756 (N_9756,N_7798,N_6553);
xor U9757 (N_9757,N_7769,N_7814);
or U9758 (N_9758,N_6896,N_7459);
nand U9759 (N_9759,N_7374,N_7461);
or U9760 (N_9760,N_7693,N_6963);
and U9761 (N_9761,N_6303,N_6491);
xor U9762 (N_9762,N_7572,N_6996);
nand U9763 (N_9763,N_6792,N_7050);
xnor U9764 (N_9764,N_7411,N_7023);
xor U9765 (N_9765,N_7219,N_6048);
nor U9766 (N_9766,N_7160,N_6329);
nand U9767 (N_9767,N_7683,N_7753);
nand U9768 (N_9768,N_6120,N_6322);
nor U9769 (N_9769,N_6022,N_6059);
xnor U9770 (N_9770,N_6130,N_6086);
nor U9771 (N_9771,N_7973,N_7075);
xnor U9772 (N_9772,N_7016,N_7463);
nand U9773 (N_9773,N_6118,N_7026);
nor U9774 (N_9774,N_6949,N_6609);
and U9775 (N_9775,N_6350,N_7553);
nand U9776 (N_9776,N_7870,N_7736);
nand U9777 (N_9777,N_7488,N_7910);
xnor U9778 (N_9778,N_6691,N_7012);
or U9779 (N_9779,N_6907,N_6950);
or U9780 (N_9780,N_6497,N_6844);
and U9781 (N_9781,N_6736,N_7227);
xnor U9782 (N_9782,N_7265,N_6458);
xnor U9783 (N_9783,N_6640,N_7507);
or U9784 (N_9784,N_7119,N_7268);
or U9785 (N_9785,N_7937,N_7227);
nand U9786 (N_9786,N_7203,N_7498);
nand U9787 (N_9787,N_6111,N_7632);
nand U9788 (N_9788,N_6163,N_7625);
nand U9789 (N_9789,N_7232,N_6487);
xor U9790 (N_9790,N_6475,N_7049);
or U9791 (N_9791,N_7048,N_6849);
or U9792 (N_9792,N_7652,N_7946);
or U9793 (N_9793,N_7623,N_7346);
xnor U9794 (N_9794,N_6575,N_6003);
or U9795 (N_9795,N_7145,N_6629);
or U9796 (N_9796,N_6175,N_6069);
or U9797 (N_9797,N_7473,N_6311);
nor U9798 (N_9798,N_6781,N_6521);
nor U9799 (N_9799,N_6840,N_6315);
nand U9800 (N_9800,N_6568,N_7496);
and U9801 (N_9801,N_7686,N_7326);
and U9802 (N_9802,N_6043,N_6730);
nor U9803 (N_9803,N_6088,N_7039);
or U9804 (N_9804,N_7063,N_7501);
and U9805 (N_9805,N_6353,N_7648);
nand U9806 (N_9806,N_7217,N_7701);
xnor U9807 (N_9807,N_7070,N_6035);
nand U9808 (N_9808,N_6644,N_7635);
or U9809 (N_9809,N_6717,N_6315);
or U9810 (N_9810,N_6324,N_6057);
xnor U9811 (N_9811,N_7703,N_7781);
nand U9812 (N_9812,N_6193,N_7391);
and U9813 (N_9813,N_6483,N_7376);
or U9814 (N_9814,N_6438,N_6270);
or U9815 (N_9815,N_7736,N_7965);
nor U9816 (N_9816,N_6644,N_7917);
or U9817 (N_9817,N_6209,N_7144);
or U9818 (N_9818,N_6615,N_6642);
or U9819 (N_9819,N_6912,N_6522);
nor U9820 (N_9820,N_7068,N_7740);
xor U9821 (N_9821,N_6182,N_6134);
or U9822 (N_9822,N_7469,N_7422);
nand U9823 (N_9823,N_6716,N_6143);
nand U9824 (N_9824,N_7809,N_7244);
xnor U9825 (N_9825,N_6819,N_7421);
and U9826 (N_9826,N_6921,N_6575);
xor U9827 (N_9827,N_6954,N_7910);
or U9828 (N_9828,N_7004,N_7650);
nand U9829 (N_9829,N_6576,N_6541);
nand U9830 (N_9830,N_7910,N_6422);
and U9831 (N_9831,N_6213,N_7095);
or U9832 (N_9832,N_7675,N_6358);
and U9833 (N_9833,N_7113,N_7012);
and U9834 (N_9834,N_7333,N_6137);
or U9835 (N_9835,N_6365,N_7903);
xor U9836 (N_9836,N_7459,N_6759);
nand U9837 (N_9837,N_6919,N_7796);
xor U9838 (N_9838,N_7785,N_7764);
nor U9839 (N_9839,N_7822,N_7483);
and U9840 (N_9840,N_6512,N_7143);
nor U9841 (N_9841,N_7699,N_7782);
and U9842 (N_9842,N_6167,N_7655);
or U9843 (N_9843,N_6634,N_6336);
nand U9844 (N_9844,N_6009,N_6072);
or U9845 (N_9845,N_6314,N_6139);
or U9846 (N_9846,N_6026,N_6819);
nor U9847 (N_9847,N_6176,N_6932);
nand U9848 (N_9848,N_6298,N_7718);
or U9849 (N_9849,N_6238,N_6036);
and U9850 (N_9850,N_6819,N_6294);
xnor U9851 (N_9851,N_7125,N_7252);
and U9852 (N_9852,N_6922,N_7264);
nand U9853 (N_9853,N_6032,N_6166);
nor U9854 (N_9854,N_6860,N_6699);
nor U9855 (N_9855,N_7412,N_7596);
xor U9856 (N_9856,N_7612,N_6869);
xor U9857 (N_9857,N_6014,N_6927);
xor U9858 (N_9858,N_6877,N_6075);
or U9859 (N_9859,N_6076,N_7600);
xor U9860 (N_9860,N_7126,N_7674);
and U9861 (N_9861,N_7070,N_7355);
and U9862 (N_9862,N_7961,N_6457);
xor U9863 (N_9863,N_7368,N_6417);
nor U9864 (N_9864,N_6406,N_6967);
and U9865 (N_9865,N_6773,N_7897);
or U9866 (N_9866,N_7664,N_7092);
and U9867 (N_9867,N_7262,N_7452);
nand U9868 (N_9868,N_6574,N_6266);
nor U9869 (N_9869,N_6497,N_6356);
nand U9870 (N_9870,N_7010,N_6993);
nor U9871 (N_9871,N_6034,N_7017);
nor U9872 (N_9872,N_6842,N_6237);
or U9873 (N_9873,N_6185,N_6799);
nand U9874 (N_9874,N_7000,N_6417);
nor U9875 (N_9875,N_7958,N_6112);
nand U9876 (N_9876,N_7882,N_7685);
xor U9877 (N_9877,N_6655,N_6759);
xnor U9878 (N_9878,N_6928,N_6912);
and U9879 (N_9879,N_7483,N_7588);
xnor U9880 (N_9880,N_6327,N_7252);
nor U9881 (N_9881,N_6220,N_7683);
nand U9882 (N_9882,N_6572,N_6930);
nor U9883 (N_9883,N_7382,N_7541);
and U9884 (N_9884,N_7845,N_7968);
nand U9885 (N_9885,N_6542,N_6317);
nand U9886 (N_9886,N_7210,N_6618);
xor U9887 (N_9887,N_7884,N_7606);
and U9888 (N_9888,N_6922,N_7613);
or U9889 (N_9889,N_7504,N_7575);
xnor U9890 (N_9890,N_7559,N_7452);
xnor U9891 (N_9891,N_6079,N_7657);
and U9892 (N_9892,N_7125,N_6665);
and U9893 (N_9893,N_6382,N_7347);
nor U9894 (N_9894,N_6505,N_7847);
xor U9895 (N_9895,N_6601,N_7597);
and U9896 (N_9896,N_7721,N_6710);
nor U9897 (N_9897,N_6089,N_6313);
nor U9898 (N_9898,N_7209,N_6346);
nand U9899 (N_9899,N_6428,N_6859);
nand U9900 (N_9900,N_7298,N_7101);
or U9901 (N_9901,N_6540,N_7547);
nor U9902 (N_9902,N_6880,N_7919);
xor U9903 (N_9903,N_6692,N_7786);
xnor U9904 (N_9904,N_6840,N_7331);
nor U9905 (N_9905,N_7661,N_7421);
and U9906 (N_9906,N_6773,N_7285);
and U9907 (N_9907,N_6675,N_7827);
nand U9908 (N_9908,N_7496,N_7109);
nor U9909 (N_9909,N_6054,N_7105);
and U9910 (N_9910,N_7246,N_7255);
and U9911 (N_9911,N_7646,N_7192);
nor U9912 (N_9912,N_6316,N_6918);
nor U9913 (N_9913,N_6577,N_7692);
nor U9914 (N_9914,N_6355,N_6887);
and U9915 (N_9915,N_7072,N_6796);
or U9916 (N_9916,N_6312,N_6965);
and U9917 (N_9917,N_6432,N_6054);
nor U9918 (N_9918,N_6244,N_7405);
xnor U9919 (N_9919,N_7165,N_7169);
or U9920 (N_9920,N_6528,N_7820);
or U9921 (N_9921,N_7892,N_7001);
or U9922 (N_9922,N_7599,N_6994);
xnor U9923 (N_9923,N_6140,N_7752);
or U9924 (N_9924,N_6150,N_7444);
and U9925 (N_9925,N_7745,N_6918);
and U9926 (N_9926,N_7090,N_7895);
xnor U9927 (N_9927,N_6202,N_7655);
and U9928 (N_9928,N_6635,N_6745);
nor U9929 (N_9929,N_7213,N_6734);
and U9930 (N_9930,N_6552,N_7267);
or U9931 (N_9931,N_7530,N_6412);
nand U9932 (N_9932,N_7709,N_6278);
or U9933 (N_9933,N_7421,N_7245);
or U9934 (N_9934,N_6720,N_7997);
nor U9935 (N_9935,N_6813,N_7486);
nor U9936 (N_9936,N_7592,N_7012);
nand U9937 (N_9937,N_6856,N_6733);
and U9938 (N_9938,N_7888,N_6526);
xor U9939 (N_9939,N_6412,N_6904);
and U9940 (N_9940,N_7626,N_6125);
nor U9941 (N_9941,N_6083,N_6201);
and U9942 (N_9942,N_7067,N_7936);
and U9943 (N_9943,N_6667,N_7277);
nor U9944 (N_9944,N_6135,N_7216);
nor U9945 (N_9945,N_6973,N_7044);
or U9946 (N_9946,N_6366,N_7630);
and U9947 (N_9947,N_6262,N_6985);
nand U9948 (N_9948,N_6105,N_6788);
nand U9949 (N_9949,N_7229,N_7242);
or U9950 (N_9950,N_7084,N_7083);
or U9951 (N_9951,N_7172,N_7022);
and U9952 (N_9952,N_7493,N_6830);
nor U9953 (N_9953,N_6910,N_6489);
and U9954 (N_9954,N_6119,N_6983);
nand U9955 (N_9955,N_7429,N_7460);
or U9956 (N_9956,N_7811,N_6796);
nor U9957 (N_9957,N_7753,N_6174);
nand U9958 (N_9958,N_6607,N_6482);
and U9959 (N_9959,N_6851,N_7013);
xor U9960 (N_9960,N_7739,N_7482);
xor U9961 (N_9961,N_6202,N_7789);
or U9962 (N_9962,N_6654,N_7100);
xnor U9963 (N_9963,N_6876,N_6423);
nor U9964 (N_9964,N_6794,N_7967);
or U9965 (N_9965,N_7865,N_7882);
nand U9966 (N_9966,N_7543,N_6633);
or U9967 (N_9967,N_6746,N_7965);
or U9968 (N_9968,N_6301,N_6425);
and U9969 (N_9969,N_6581,N_7571);
and U9970 (N_9970,N_7164,N_6757);
or U9971 (N_9971,N_7523,N_6347);
and U9972 (N_9972,N_6354,N_7184);
xnor U9973 (N_9973,N_7065,N_6236);
xor U9974 (N_9974,N_6692,N_7307);
and U9975 (N_9975,N_7871,N_7246);
xor U9976 (N_9976,N_6685,N_6224);
xnor U9977 (N_9977,N_6567,N_7858);
or U9978 (N_9978,N_6581,N_7544);
xnor U9979 (N_9979,N_7900,N_7619);
xnor U9980 (N_9980,N_6251,N_7650);
nor U9981 (N_9981,N_7917,N_7604);
nor U9982 (N_9982,N_7806,N_7140);
xnor U9983 (N_9983,N_6471,N_6003);
nand U9984 (N_9984,N_7701,N_6275);
and U9985 (N_9985,N_7906,N_7743);
or U9986 (N_9986,N_6127,N_6583);
nor U9987 (N_9987,N_7045,N_6784);
nor U9988 (N_9988,N_6522,N_6347);
xnor U9989 (N_9989,N_6344,N_6665);
nand U9990 (N_9990,N_6212,N_6884);
nor U9991 (N_9991,N_6314,N_6136);
or U9992 (N_9992,N_6341,N_6078);
or U9993 (N_9993,N_7608,N_7706);
nor U9994 (N_9994,N_6251,N_7605);
xnor U9995 (N_9995,N_7545,N_6384);
nand U9996 (N_9996,N_7957,N_7879);
nand U9997 (N_9997,N_7703,N_6235);
and U9998 (N_9998,N_6226,N_6507);
nand U9999 (N_9999,N_7558,N_7962);
nand U10000 (N_10000,N_9480,N_8890);
xnor U10001 (N_10001,N_9952,N_9324);
and U10002 (N_10002,N_8120,N_8446);
or U10003 (N_10003,N_8845,N_9907);
nor U10004 (N_10004,N_8458,N_9760);
xor U10005 (N_10005,N_8726,N_9006);
nor U10006 (N_10006,N_8755,N_9742);
nor U10007 (N_10007,N_8640,N_9404);
or U10008 (N_10008,N_8712,N_8113);
nor U10009 (N_10009,N_9401,N_8247);
nor U10010 (N_10010,N_9600,N_8613);
nor U10011 (N_10011,N_8894,N_8677);
nor U10012 (N_10012,N_9531,N_9367);
xnor U10013 (N_10013,N_8034,N_9921);
nand U10014 (N_10014,N_9008,N_9276);
nand U10015 (N_10015,N_9451,N_9486);
nand U10016 (N_10016,N_8339,N_9287);
nand U10017 (N_10017,N_9696,N_8630);
or U10018 (N_10018,N_9235,N_9745);
nor U10019 (N_10019,N_8179,N_8370);
or U10020 (N_10020,N_9337,N_8790);
or U10021 (N_10021,N_9091,N_9120);
or U10022 (N_10022,N_9378,N_9660);
nand U10023 (N_10023,N_8936,N_8468);
and U10024 (N_10024,N_9776,N_8929);
nand U10025 (N_10025,N_9520,N_8357);
nand U10026 (N_10026,N_8500,N_8607);
and U10027 (N_10027,N_9260,N_9042);
or U10028 (N_10028,N_9316,N_8896);
nor U10029 (N_10029,N_8056,N_8729);
nand U10030 (N_10030,N_8987,N_9107);
xnor U10031 (N_10031,N_9535,N_8157);
nor U10032 (N_10032,N_8307,N_9308);
or U10033 (N_10033,N_9695,N_8941);
nand U10034 (N_10034,N_9428,N_8840);
xnor U10035 (N_10035,N_8184,N_9497);
nand U10036 (N_10036,N_9547,N_9982);
xnor U10037 (N_10037,N_8895,N_9432);
xnor U10038 (N_10038,N_9821,N_8185);
and U10039 (N_10039,N_9593,N_8150);
nand U10040 (N_10040,N_9626,N_9927);
and U10041 (N_10041,N_8898,N_9291);
or U10042 (N_10042,N_8881,N_9941);
or U10043 (N_10043,N_8560,N_8750);
nand U10044 (N_10044,N_8336,N_9393);
and U10045 (N_10045,N_8545,N_9067);
nand U10046 (N_10046,N_8277,N_8624);
and U10047 (N_10047,N_9476,N_9686);
nor U10048 (N_10048,N_8988,N_9680);
nor U10049 (N_10049,N_9720,N_8015);
nand U10050 (N_10050,N_8550,N_8783);
nand U10051 (N_10051,N_8749,N_8200);
nand U10052 (N_10052,N_9346,N_9199);
xor U10053 (N_10053,N_8511,N_8576);
xor U10054 (N_10054,N_9658,N_9266);
and U10055 (N_10055,N_8662,N_9714);
and U10056 (N_10056,N_8658,N_8097);
and U10057 (N_10057,N_8258,N_9523);
or U10058 (N_10058,N_8009,N_8018);
nand U10059 (N_10059,N_8391,N_8463);
nand U10060 (N_10060,N_9074,N_8809);
xor U10061 (N_10061,N_9153,N_9043);
xnor U10062 (N_10062,N_8403,N_8163);
or U10063 (N_10063,N_8280,N_9784);
nor U10064 (N_10064,N_9648,N_8058);
xnor U10065 (N_10065,N_9550,N_9492);
xor U10066 (N_10066,N_9105,N_9746);
and U10067 (N_10067,N_9831,N_8700);
xor U10068 (N_10068,N_9450,N_8714);
or U10069 (N_10069,N_9127,N_9728);
or U10070 (N_10070,N_9464,N_9258);
nor U10071 (N_10071,N_8326,N_8919);
or U10072 (N_10072,N_9167,N_8615);
nand U10073 (N_10073,N_9394,N_8872);
nor U10074 (N_10074,N_9837,N_9479);
or U10075 (N_10075,N_9910,N_9913);
or U10076 (N_10076,N_9248,N_9779);
and U10077 (N_10077,N_9473,N_9937);
nand U10078 (N_10078,N_8868,N_9062);
nand U10079 (N_10079,N_8429,N_8693);
or U10080 (N_10080,N_9458,N_9433);
nand U10081 (N_10081,N_8186,N_8431);
xnor U10082 (N_10082,N_8367,N_8853);
nand U10083 (N_10083,N_8527,N_9577);
nand U10084 (N_10084,N_9771,N_8295);
and U10085 (N_10085,N_8273,N_9659);
or U10086 (N_10086,N_9886,N_9676);
and U10087 (N_10087,N_9007,N_9560);
nor U10088 (N_10088,N_9574,N_9059);
xor U10089 (N_10089,N_8368,N_9084);
or U10090 (N_10090,N_9970,N_9114);
nor U10091 (N_10091,N_9202,N_9440);
nand U10092 (N_10092,N_8333,N_9434);
and U10093 (N_10093,N_8785,N_8837);
nand U10094 (N_10094,N_9339,N_8535);
nand U10095 (N_10095,N_9573,N_9756);
or U10096 (N_10096,N_8397,N_8471);
or U10097 (N_10097,N_9549,N_9923);
or U10098 (N_10098,N_9809,N_9942);
nor U10099 (N_10099,N_8407,N_9160);
xnor U10100 (N_10100,N_8042,N_9350);
nand U10101 (N_10101,N_8452,N_9280);
and U10102 (N_10102,N_8180,N_8860);
and U10103 (N_10103,N_8760,N_9901);
nand U10104 (N_10104,N_8946,N_8032);
nand U10105 (N_10105,N_9027,N_9625);
or U10106 (N_10106,N_9786,N_9887);
nand U10107 (N_10107,N_9375,N_9187);
nor U10108 (N_10108,N_9704,N_8383);
nand U10109 (N_10109,N_9161,N_9524);
xnor U10110 (N_10110,N_8756,N_8076);
nor U10111 (N_10111,N_8008,N_9748);
nor U10112 (N_10112,N_8128,N_9672);
or U10113 (N_10113,N_8192,N_8718);
nor U10114 (N_10114,N_8181,N_8650);
xnor U10115 (N_10115,N_9169,N_8083);
nor U10116 (N_10116,N_8472,N_9788);
or U10117 (N_10117,N_9113,N_8591);
nand U10118 (N_10118,N_9782,N_8390);
xnor U10119 (N_10119,N_9493,N_9979);
nand U10120 (N_10120,N_9854,N_8546);
nand U10121 (N_10121,N_9569,N_8582);
xnor U10122 (N_10122,N_9594,N_9139);
nand U10123 (N_10123,N_9190,N_9866);
nand U10124 (N_10124,N_8937,N_8515);
or U10125 (N_10125,N_9500,N_8796);
nor U10126 (N_10126,N_8870,N_9320);
xor U10127 (N_10127,N_9951,N_8854);
or U10128 (N_10128,N_9206,N_8023);
and U10129 (N_10129,N_9912,N_8817);
xnor U10130 (N_10130,N_9013,N_8093);
nand U10131 (N_10131,N_9305,N_9331);
or U10132 (N_10132,N_8835,N_8909);
nand U10133 (N_10133,N_9508,N_9570);
or U10134 (N_10134,N_9616,N_8994);
xor U10135 (N_10135,N_8297,N_8969);
and U10136 (N_10136,N_9278,N_9752);
xor U10137 (N_10137,N_8255,N_9505);
nand U10138 (N_10138,N_9232,N_9640);
nor U10139 (N_10139,N_8141,N_9882);
and U10140 (N_10140,N_9985,N_9037);
or U10141 (N_10141,N_9210,N_9973);
xor U10142 (N_10142,N_8570,N_8622);
nand U10143 (N_10143,N_9471,N_8657);
nand U10144 (N_10144,N_9203,N_9922);
xor U10145 (N_10145,N_9368,N_8880);
nand U10146 (N_10146,N_8966,N_8938);
nor U10147 (N_10147,N_9272,N_8879);
or U10148 (N_10148,N_8884,N_8027);
xor U10149 (N_10149,N_9192,N_8832);
and U10150 (N_10150,N_8432,N_9030);
or U10151 (N_10151,N_9727,N_8174);
nand U10152 (N_10152,N_9466,N_8107);
and U10153 (N_10153,N_8318,N_9209);
nand U10154 (N_10154,N_9135,N_8112);
nand U10155 (N_10155,N_8782,N_9335);
xor U10156 (N_10156,N_9284,N_8285);
nor U10157 (N_10157,N_8968,N_8822);
nand U10158 (N_10158,N_8286,N_9805);
nor U10159 (N_10159,N_9313,N_9950);
nor U10160 (N_10160,N_8069,N_9358);
xor U10161 (N_10161,N_8469,N_8460);
nor U10162 (N_10162,N_9413,N_9140);
nor U10163 (N_10163,N_8340,N_8201);
or U10164 (N_10164,N_9935,N_9662);
nand U10165 (N_10165,N_8557,N_8897);
or U10166 (N_10166,N_9632,N_9986);
nand U10167 (N_10167,N_9802,N_9468);
nor U10168 (N_10168,N_8161,N_8971);
nand U10169 (N_10169,N_8239,N_8972);
xnor U10170 (N_10170,N_8165,N_8457);
or U10171 (N_10171,N_8648,N_8989);
and U10172 (N_10172,N_8135,N_9296);
or U10173 (N_10173,N_9005,N_9637);
nor U10174 (N_10174,N_9829,N_9791);
nand U10175 (N_10175,N_9281,N_9086);
xnor U10176 (N_10176,N_9900,N_9603);
nand U10177 (N_10177,N_8634,N_9615);
nor U10178 (N_10178,N_9124,N_8341);
nand U10179 (N_10179,N_8321,N_9863);
nand U10180 (N_10180,N_8730,N_9092);
xor U10181 (N_10181,N_8281,N_9373);
and U10182 (N_10182,N_8598,N_8133);
nand U10183 (N_10183,N_8825,N_8310);
nand U10184 (N_10184,N_8044,N_8385);
nand U10185 (N_10185,N_8268,N_9398);
and U10186 (N_10186,N_9799,N_8699);
or U10187 (N_10187,N_8587,N_8522);
nor U10188 (N_10188,N_8100,N_8625);
and U10189 (N_10189,N_8493,N_9944);
nor U10190 (N_10190,N_8621,N_8815);
or U10191 (N_10191,N_9587,N_8046);
xnor U10192 (N_10192,N_8057,N_8918);
nand U10193 (N_10193,N_9083,N_9638);
nand U10194 (N_10194,N_9933,N_9811);
and U10195 (N_10195,N_9087,N_8928);
or U10196 (N_10196,N_8529,N_8102);
and U10197 (N_10197,N_8156,N_8577);
or U10198 (N_10198,N_9909,N_8882);
or U10199 (N_10199,N_8002,N_9095);
nand U10200 (N_10200,N_8235,N_8272);
xor U10201 (N_10201,N_8911,N_8850);
xnor U10202 (N_10202,N_9691,N_8190);
nor U10203 (N_10203,N_9411,N_9274);
nand U10204 (N_10204,N_9804,N_9381);
and U10205 (N_10205,N_8505,N_9024);
or U10206 (N_10206,N_9624,N_8262);
nor U10207 (N_10207,N_8296,N_8148);
xor U10208 (N_10208,N_9732,N_9814);
or U10209 (N_10209,N_8199,N_9689);
xnor U10210 (N_10210,N_8082,N_8776);
xnor U10211 (N_10211,N_9004,N_8743);
or U10212 (N_10212,N_9726,N_9553);
nand U10213 (N_10213,N_9983,N_8438);
nand U10214 (N_10214,N_8865,N_8217);
xnor U10215 (N_10215,N_9038,N_9555);
xnor U10216 (N_10216,N_9009,N_8910);
xor U10217 (N_10217,N_9894,N_8487);
nand U10218 (N_10218,N_8606,N_8095);
xor U10219 (N_10219,N_8751,N_9302);
nor U10220 (N_10220,N_8701,N_8467);
nor U10221 (N_10221,N_8787,N_8584);
xnor U10222 (N_10222,N_9895,N_9967);
xor U10223 (N_10223,N_8494,N_8433);
nand U10224 (N_10224,N_8552,N_9045);
nor U10225 (N_10225,N_9976,N_9338);
nand U10226 (N_10226,N_8702,N_9818);
nand U10227 (N_10227,N_9562,N_8050);
nor U10228 (N_10228,N_8697,N_8033);
nand U10229 (N_10229,N_9864,N_9801);
nor U10230 (N_10230,N_9217,N_9988);
nand U10231 (N_10231,N_8228,N_9049);
nand U10232 (N_10232,N_8775,N_8167);
nand U10233 (N_10233,N_8293,N_9152);
nor U10234 (N_10234,N_9147,N_8883);
nor U10235 (N_10235,N_9806,N_9230);
xor U10236 (N_10236,N_9439,N_8921);
nand U10237 (N_10237,N_8792,N_9231);
nor U10238 (N_10238,N_9376,N_8311);
nor U10239 (N_10239,N_8427,N_9442);
and U10240 (N_10240,N_8331,N_9627);
or U10241 (N_10241,N_9684,N_9245);
nand U10242 (N_10242,N_8829,N_9077);
nand U10243 (N_10243,N_8684,N_8365);
nor U10244 (N_10244,N_8226,N_9993);
nand U10245 (N_10245,N_8520,N_8636);
or U10246 (N_10246,N_9034,N_8484);
xor U10247 (N_10247,N_9185,N_8253);
xnor U10248 (N_10248,N_9417,N_8745);
xor U10249 (N_10249,N_9852,N_8111);
and U10250 (N_10250,N_8735,N_8949);
or U10251 (N_10251,N_8134,N_9138);
xor U10252 (N_10252,N_8371,N_8542);
nor U10253 (N_10253,N_9292,N_9934);
nor U10254 (N_10254,N_9244,N_9054);
and U10255 (N_10255,N_8637,N_9406);
and U10256 (N_10256,N_8572,N_8764);
and U10257 (N_10257,N_8394,N_8816);
xnor U10258 (N_10258,N_8806,N_9265);
or U10259 (N_10259,N_8152,N_9995);
or U10260 (N_10260,N_8270,N_9136);
and U10261 (N_10261,N_9360,N_8302);
and U10262 (N_10262,N_8335,N_8079);
xnor U10263 (N_10263,N_9957,N_9867);
nor U10264 (N_10264,N_8000,N_9670);
nor U10265 (N_10265,N_9039,N_8222);
or U10266 (N_10266,N_8154,N_8106);
and U10267 (N_10267,N_8388,N_8182);
nor U10268 (N_10268,N_9298,N_9184);
xnor U10269 (N_10269,N_8599,N_9405);
and U10270 (N_10270,N_9908,N_8678);
nand U10271 (N_10271,N_8740,N_9762);
nand U10272 (N_10272,N_8935,N_9551);
nor U10273 (N_10273,N_9036,N_9869);
nor U10274 (N_10274,N_8719,N_8410);
nand U10275 (N_10275,N_8773,N_8260);
or U10276 (N_10276,N_8836,N_8225);
and U10277 (N_10277,N_8671,N_9647);
or U10278 (N_10278,N_9056,N_9905);
nor U10279 (N_10279,N_8830,N_9889);
nand U10280 (N_10280,N_8387,N_8944);
nor U10281 (N_10281,N_8954,N_8877);
and U10282 (N_10282,N_9507,N_8246);
nor U10283 (N_10283,N_8215,N_9702);
nand U10284 (N_10284,N_9117,N_8132);
or U10285 (N_10285,N_8705,N_9014);
nor U10286 (N_10286,N_8811,N_9962);
xnor U10287 (N_10287,N_9939,N_8384);
and U10288 (N_10288,N_8558,N_9467);
or U10289 (N_10289,N_8498,N_9607);
nor U10290 (N_10290,N_9755,N_8412);
or U10291 (N_10291,N_9736,N_9629);
and U10292 (N_10292,N_8805,N_8818);
nor U10293 (N_10293,N_8035,N_9477);
nor U10294 (N_10294,N_9264,N_8031);
xor U10295 (N_10295,N_8006,N_8103);
nand U10296 (N_10296,N_9588,N_8172);
nand U10297 (N_10297,N_9125,N_8011);
or U10298 (N_10298,N_9872,N_9242);
nor U10299 (N_10299,N_9424,N_8556);
xor U10300 (N_10300,N_9999,N_9875);
xnor U10301 (N_10301,N_9307,N_8202);
or U10302 (N_10302,N_8129,N_8820);
or U10303 (N_10303,N_8254,N_8999);
or U10304 (N_10304,N_8708,N_8916);
and U10305 (N_10305,N_9026,N_8908);
nor U10306 (N_10306,N_8761,N_9080);
and U10307 (N_10307,N_8862,N_9873);
xor U10308 (N_10308,N_9183,N_9142);
or U10309 (N_10309,N_9228,N_9494);
nand U10310 (N_10310,N_9787,N_9366);
xor U10311 (N_10311,N_8261,N_8278);
or U10312 (N_10312,N_8109,N_9475);
nor U10313 (N_10313,N_9633,N_9098);
nand U10314 (N_10314,N_9585,N_9552);
and U10315 (N_10315,N_8732,N_9137);
nor U10316 (N_10316,N_9019,N_9709);
nor U10317 (N_10317,N_8844,N_8642);
nor U10318 (N_10318,N_8716,N_9327);
nor U10319 (N_10319,N_9579,N_8171);
nand U10320 (N_10320,N_9711,N_8334);
nor U10321 (N_10321,N_8715,N_9251);
and U10322 (N_10322,N_9016,N_9953);
or U10323 (N_10323,N_9874,N_8950);
nand U10324 (N_10324,N_8401,N_9774);
xnor U10325 (N_10325,N_9017,N_8800);
nor U10326 (N_10326,N_8543,N_9075);
nor U10327 (N_10327,N_8052,N_9236);
nand U10328 (N_10328,N_9652,N_8160);
or U10329 (N_10329,N_8029,N_8823);
nor U10330 (N_10330,N_9273,N_8574);
nand U10331 (N_10331,N_8610,N_8985);
or U10332 (N_10332,N_8669,N_8026);
and U10333 (N_10333,N_9133,N_9385);
and U10334 (N_10334,N_9758,N_8110);
nor U10335 (N_10335,N_9041,N_9919);
nor U10336 (N_10336,N_9825,N_8963);
and U10337 (N_10337,N_9644,N_8528);
nand U10338 (N_10338,N_9241,N_9861);
nor U10339 (N_10339,N_9369,N_9845);
xor U10340 (N_10340,N_8428,N_8004);
and U10341 (N_10341,N_8580,N_8734);
nand U10342 (N_10342,N_8727,N_9753);
and U10343 (N_10343,N_9835,N_8514);
xor U10344 (N_10344,N_9741,N_9849);
nor U10345 (N_10345,N_9365,N_8967);
xor U10346 (N_10346,N_9182,N_9021);
nand U10347 (N_10347,N_8984,N_8548);
nand U10348 (N_10348,N_8763,N_8398);
xnor U10349 (N_10349,N_8549,N_8234);
xor U10350 (N_10350,N_8306,N_8858);
xnor U10351 (N_10351,N_8300,N_9194);
nand U10352 (N_10352,N_9955,N_9181);
xor U10353 (N_10353,N_8440,N_9673);
nand U10354 (N_10354,N_9700,N_9100);
or U10355 (N_10355,N_8218,N_9294);
nor U10356 (N_10356,N_9051,N_8094);
or U10357 (N_10357,N_8137,N_8435);
nor U10358 (N_10358,N_8481,N_8409);
nor U10359 (N_10359,N_8155,N_8633);
or U10360 (N_10360,N_9639,N_9154);
nand U10361 (N_10361,N_8583,N_9470);
and U10362 (N_10362,N_9390,N_9108);
xor U10363 (N_10363,N_8251,N_8197);
nor U10364 (N_10364,N_9800,N_8426);
nand U10365 (N_10365,N_8342,N_8758);
or U10366 (N_10366,N_8065,N_8242);
xor U10367 (N_10367,N_8245,N_9126);
nand U10368 (N_10368,N_8748,N_9364);
xor U10369 (N_10369,N_8329,N_9462);
nor U10370 (N_10370,N_8934,N_9881);
nand U10371 (N_10371,N_8126,N_8833);
nor U10372 (N_10372,N_8352,N_9506);
or U10373 (N_10373,N_8455,N_9106);
and U10374 (N_10374,N_8289,N_9430);
nor U10375 (N_10375,N_9383,N_8140);
or U10376 (N_10376,N_9511,N_9176);
nor U10377 (N_10377,N_8793,N_9556);
or U10378 (N_10378,N_9819,N_9522);
nand U10379 (N_10379,N_8090,N_9572);
nor U10380 (N_10380,N_8924,N_9698);
xor U10381 (N_10381,N_8096,N_8416);
or U10382 (N_10382,N_8831,N_8308);
or U10383 (N_10383,N_9645,N_9071);
or U10384 (N_10384,N_8964,N_8762);
or U10385 (N_10385,N_8495,N_9575);
nor U10386 (N_10386,N_9115,N_9839);
nand U10387 (N_10387,N_8283,N_9388);
and U10388 (N_10388,N_8153,N_8489);
nand U10389 (N_10389,N_8901,N_9205);
nand U10390 (N_10390,N_8864,N_8889);
or U10391 (N_10391,N_8169,N_9833);
or U10392 (N_10392,N_8077,N_8784);
and U10393 (N_10393,N_9767,N_8781);
nor U10394 (N_10394,N_8553,N_9218);
nand U10395 (N_10395,N_8942,N_8675);
or U10396 (N_10396,N_8539,N_9865);
nand U10397 (N_10397,N_8315,N_9254);
and U10398 (N_10398,N_9737,N_9420);
nor U10399 (N_10399,N_8476,N_8191);
nor U10400 (N_10400,N_9643,N_9286);
or U10401 (N_10401,N_9314,N_8485);
xnor U10402 (N_10402,N_9392,N_9893);
nand U10403 (N_10403,N_8064,N_9079);
nor U10404 (N_10404,N_9070,N_9333);
and U10405 (N_10405,N_8275,N_9116);
xnor U10406 (N_10406,N_8149,N_8744);
and U10407 (N_10407,N_8801,N_9850);
and U10408 (N_10408,N_8932,N_8389);
nand U10409 (N_10409,N_9978,N_8208);
xor U10410 (N_10410,N_8863,N_8089);
xor U10411 (N_10411,N_8562,N_9773);
nor U10412 (N_10412,N_9597,N_8777);
nor U10413 (N_10413,N_9224,N_9820);
nor U10414 (N_10414,N_9789,N_9938);
and U10415 (N_10415,N_8119,N_9992);
nand U10416 (N_10416,N_9884,N_9883);
and U10417 (N_10417,N_8256,N_8869);
nand U10418 (N_10418,N_8914,N_8211);
nor U10419 (N_10419,N_9452,N_9734);
and U10420 (N_10420,N_9422,N_9399);
nor U10421 (N_10421,N_9740,N_9816);
nor U10422 (N_10422,N_9055,N_9605);
xor U10423 (N_10423,N_9824,N_8224);
nand U10424 (N_10424,N_9453,N_9073);
xor U10425 (N_10425,N_9454,N_8014);
nand U10426 (N_10426,N_9403,N_9198);
xor U10427 (N_10427,N_9534,N_8561);
xnor U10428 (N_10428,N_8480,N_9924);
nand U10429 (N_10429,N_8961,N_8482);
nor U10430 (N_10430,N_9104,N_8417);
nor U10431 (N_10431,N_9196,N_8670);
or U10432 (N_10432,N_9018,N_9917);
or U10433 (N_10433,N_8206,N_9823);
and U10434 (N_10434,N_9757,N_8024);
nand U10435 (N_10435,N_8953,N_8330);
or U10436 (N_10436,N_8314,N_9357);
nand U10437 (N_10437,N_8673,N_8164);
nor U10438 (N_10438,N_9380,N_9926);
nand U10439 (N_10439,N_9118,N_9299);
nand U10440 (N_10440,N_9151,N_9620);
nand U10441 (N_10441,N_9020,N_9048);
or U10442 (N_10442,N_8531,N_8683);
xnor U10443 (N_10443,N_8720,N_9495);
and U10444 (N_10444,N_9925,N_9810);
or U10445 (N_10445,N_9966,N_9743);
nand U10446 (N_10446,N_8780,N_8223);
nand U10447 (N_10447,N_8080,N_8997);
nand U10448 (N_10448,N_9033,N_8054);
and U10449 (N_10449,N_8979,N_8204);
nor U10450 (N_10450,N_8986,N_8439);
nor U10451 (N_10451,N_8579,N_8687);
and U10452 (N_10452,N_8581,N_9148);
and U10453 (N_10453,N_9447,N_9396);
nand U10454 (N_10454,N_9311,N_8980);
xor U10455 (N_10455,N_9318,N_9253);
xor U10456 (N_10456,N_9304,N_8788);
xnor U10457 (N_10457,N_9397,N_9076);
nand U10458 (N_10458,N_8212,N_9469);
or U10459 (N_10459,N_8721,N_8361);
nand U10460 (N_10460,N_9733,N_8674);
and U10461 (N_10461,N_8958,N_8635);
nor U10462 (N_10462,N_8363,N_9418);
xor U10463 (N_10463,N_8876,N_8386);
xor U10464 (N_10464,N_9400,N_9631);
nand U10465 (N_10465,N_9618,N_9554);
nand U10466 (N_10466,N_9096,N_8643);
nor U10467 (N_10467,N_9915,N_9612);
or U10468 (N_10468,N_9681,N_8906);
or U10469 (N_10469,N_8526,N_8516);
nand U10470 (N_10470,N_8605,N_9227);
and U10471 (N_10471,N_9195,N_9427);
nand U10472 (N_10472,N_8162,N_9174);
or U10473 (N_10473,N_8436,N_9892);
xnor U10474 (N_10474,N_8940,N_8142);
and U10475 (N_10475,N_9948,N_8136);
nor U10476 (N_10476,N_8305,N_8652);
nor U10477 (N_10477,N_9436,N_8138);
or U10478 (N_10478,N_8519,N_9180);
xor U10479 (N_10479,N_9790,N_8873);
xnor U10480 (N_10480,N_9257,N_8866);
nor U10481 (N_10481,N_9330,N_9223);
xor U10482 (N_10482,N_9751,N_9353);
nand U10483 (N_10483,N_8437,N_8789);
xor U10484 (N_10484,N_8430,N_9409);
or U10485 (N_10485,N_8904,N_8473);
and U10486 (N_10486,N_8249,N_8448);
and U10487 (N_10487,N_8373,N_8317);
nor U10488 (N_10488,N_9536,N_8741);
or U10489 (N_10489,N_9035,N_9518);
and U10490 (N_10490,N_8183,N_9191);
and U10491 (N_10491,N_8538,N_8214);
nor U10492 (N_10492,N_9525,N_8379);
nor U10493 (N_10493,N_9391,N_9201);
nor U10494 (N_10494,N_8282,N_9310);
nand U10495 (N_10495,N_9031,N_8685);
or U10496 (N_10496,N_8074,N_8955);
nor U10497 (N_10497,N_9208,N_9300);
nor U10498 (N_10498,N_9984,N_8187);
xnor U10499 (N_10499,N_8450,N_9168);
nor U10500 (N_10500,N_9783,N_8803);
nor U10501 (N_10501,N_9747,N_9717);
or U10502 (N_10502,N_9628,N_8686);
nor U10503 (N_10503,N_9656,N_8252);
and U10504 (N_10504,N_9363,N_9694);
nor U10505 (N_10505,N_9954,N_8993);
xnor U10506 (N_10506,N_9876,N_9785);
xor U10507 (N_10507,N_9134,N_8992);
nand U10508 (N_10508,N_8654,N_9188);
or U10509 (N_10509,N_9541,N_8629);
xnor U10510 (N_10510,N_8604,N_9022);
or U10511 (N_10511,N_8325,N_9288);
and U10512 (N_10512,N_9220,N_9445);
xor U10513 (N_10513,N_8668,N_8888);
nor U10514 (N_10514,N_9646,N_9456);
xor U10515 (N_10515,N_9010,N_8062);
or U10516 (N_10516,N_9611,N_9384);
nand U10517 (N_10517,N_8488,N_9677);
nand U10518 (N_10518,N_9159,N_9249);
and U10519 (N_10519,N_8168,N_9794);
or U10520 (N_10520,N_8351,N_8619);
nor U10521 (N_10521,N_9444,N_9642);
and U10522 (N_10522,N_9141,N_9690);
or U10523 (N_10523,N_8738,N_9687);
and U10524 (N_10524,N_8952,N_8585);
or U10525 (N_10525,N_9455,N_8802);
nand U10526 (N_10526,N_9598,N_8828);
nor U10527 (N_10527,N_8616,N_9699);
nand U10528 (N_10528,N_9904,N_8360);
xor U10529 (N_10529,N_9465,N_8287);
and U10530 (N_10530,N_9057,N_9584);
and U10531 (N_10531,N_9827,N_8243);
nand U10532 (N_10532,N_8028,N_8358);
or U10533 (N_10533,N_9193,N_9571);
and U10534 (N_10534,N_9731,N_8834);
nand U10535 (N_10535,N_8125,N_8568);
or U10536 (N_10536,N_9047,N_8917);
nand U10537 (N_10537,N_9050,N_8981);
xnor U10538 (N_10538,N_8507,N_9998);
nor U10539 (N_10539,N_8976,N_9651);
nand U10540 (N_10540,N_8346,N_8170);
and U10541 (N_10541,N_9793,N_9359);
and U10542 (N_10542,N_8534,N_9341);
xnor U10543 (N_10543,N_9608,N_8478);
or U10544 (N_10544,N_8127,N_9247);
xnor U10545 (N_10545,N_8017,N_9374);
xor U10546 (N_10546,N_8399,N_8337);
and U10547 (N_10547,N_8878,N_8575);
and U10548 (N_10548,N_9132,N_9243);
xor U10549 (N_10549,N_8404,N_9501);
nand U10550 (N_10550,N_9060,N_9377);
xnor U10551 (N_10551,N_8824,N_8205);
xor U10552 (N_10552,N_8470,N_9943);
nand U10553 (N_10553,N_8752,N_8907);
xor U10554 (N_10554,N_9122,N_9896);
xor U10555 (N_10555,N_9309,N_9129);
or U10556 (N_10556,N_8930,N_8893);
xor U10557 (N_10557,N_8380,N_9303);
nor U10558 (N_10558,N_9530,N_8506);
xnor U10559 (N_10559,N_9974,N_9564);
nor U10560 (N_10560,N_8725,N_9968);
xor U10561 (N_10561,N_8962,N_9001);
xor U10562 (N_10562,N_9693,N_9617);
or U10563 (N_10563,N_9958,N_9226);
or U10564 (N_10564,N_8477,N_9581);
xor U10565 (N_10565,N_8679,N_8656);
nand U10566 (N_10566,N_8422,N_9482);
xnor U10567 (N_10567,N_8861,N_9128);
and U10568 (N_10568,N_8852,N_9634);
or U10569 (N_10569,N_9046,N_8343);
xnor U10570 (N_10570,N_9947,N_9319);
and U10571 (N_10571,N_8354,N_8257);
and U10572 (N_10572,N_8048,N_9880);
nor U10573 (N_10573,N_9931,N_8945);
nand U10574 (N_10574,N_9636,N_9754);
and U10575 (N_10575,N_8415,N_8681);
xnor U10576 (N_10576,N_8517,N_9622);
nand U10577 (N_10577,N_8933,N_9178);
and U10578 (N_10578,N_9352,N_9109);
or U10579 (N_10579,N_8563,N_8123);
and U10580 (N_10580,N_9940,N_8250);
or U10581 (N_10581,N_8382,N_8188);
or U10582 (N_10582,N_8723,N_9989);
and U10583 (N_10583,N_9110,N_8617);
nor U10584 (N_10584,N_8055,N_9685);
nor U10585 (N_10585,N_9580,N_8759);
xor U10586 (N_10586,N_8626,N_8101);
and U10587 (N_10587,N_9130,N_9498);
xnor U10588 (N_10588,N_9170,N_9526);
nor U10589 (N_10589,N_9813,N_9614);
nand U10590 (N_10590,N_9186,N_8791);
xnor U10591 (N_10591,N_8826,N_9537);
or U10592 (N_10592,N_8115,N_9932);
or U10593 (N_10593,N_9703,N_8856);
nand U10594 (N_10594,N_9715,N_9730);
and U10595 (N_10595,N_9355,N_9665);
or U10596 (N_10596,N_9271,N_9252);
nand U10597 (N_10597,N_8073,N_9343);
nand U10598 (N_10598,N_8586,N_8328);
or U10599 (N_10599,N_9275,N_8536);
xnor U10600 (N_10600,N_8421,N_8290);
or U10601 (N_10601,N_8362,N_9960);
or U10602 (N_10602,N_8765,N_8839);
or U10603 (N_10603,N_9844,N_8717);
xor U10604 (N_10604,N_8227,N_9173);
xnor U10605 (N_10605,N_8271,N_9015);
or U10606 (N_10606,N_9532,N_8923);
nor U10607 (N_10607,N_8886,N_8393);
nor U10608 (N_10608,N_8324,N_9514);
and U10609 (N_10609,N_9328,N_8418);
and U10610 (N_10610,N_8509,N_9279);
or U10611 (N_10611,N_9664,N_8045);
xnor U10612 (N_10612,N_9540,N_8219);
or U10613 (N_10613,N_8423,N_8742);
or U10614 (N_10614,N_8903,N_9078);
xor U10615 (N_10615,N_9956,N_9144);
and U10616 (N_10616,N_8647,N_8266);
xnor U10617 (N_10617,N_8644,N_9012);
xor U10618 (N_10618,N_8366,N_8118);
nand U10619 (N_10619,N_8594,N_8319);
nand U10620 (N_10620,N_9759,N_8178);
or U10621 (N_10621,N_8461,N_9166);
nand U10622 (N_10622,N_8099,N_8794);
or U10623 (N_10623,N_8757,N_8541);
nor U10624 (N_10624,N_8276,N_9661);
nor U10625 (N_10625,N_8036,N_8728);
or U10626 (N_10626,N_8263,N_8592);
nand U10627 (N_10627,N_8960,N_9165);
and U10628 (N_10628,N_9596,N_8338);
nor U10629 (N_10629,N_9697,N_8406);
xnor U10630 (N_10630,N_9312,N_9987);
nand U10631 (N_10631,N_9650,N_8849);
nand U10632 (N_10632,N_8060,N_9028);
nand U10633 (N_10633,N_9764,N_9234);
xor U10634 (N_10634,N_8667,N_9851);
and U10635 (N_10635,N_9065,N_9155);
nand U10636 (N_10636,N_9857,N_8661);
and U10637 (N_10637,N_8116,N_8207);
nor U10638 (N_10638,N_8301,N_8694);
xor U10639 (N_10639,N_8047,N_9345);
or U10640 (N_10640,N_9484,N_8198);
or U10641 (N_10641,N_9663,N_9214);
or U10642 (N_10642,N_9928,N_9542);
nand U10643 (N_10643,N_8075,N_9496);
and U10644 (N_10644,N_8259,N_8496);
or U10645 (N_10645,N_9326,N_9914);
or U10646 (N_10646,N_8827,N_8237);
or U10647 (N_10647,N_9334,N_9221);
and U10648 (N_10648,N_9847,N_8965);
nor U10649 (N_10649,N_9855,N_9842);
and U10650 (N_10650,N_8691,N_8887);
nor U10651 (N_10651,N_8072,N_8733);
nand U10652 (N_10652,N_8554,N_8808);
xnor U10653 (N_10653,N_8867,N_8139);
nor U10654 (N_10654,N_9807,N_8210);
and U10655 (N_10655,N_9163,N_8121);
xnor U10656 (N_10656,N_8040,N_8071);
nor U10657 (N_10657,N_8349,N_9053);
or U10658 (N_10658,N_8016,N_8532);
nor U10659 (N_10659,N_9735,N_9619);
and U10660 (N_10660,N_9654,N_9349);
and U10661 (N_10661,N_8544,N_9146);
and U10662 (N_10662,N_9121,N_8104);
nor U10663 (N_10663,N_9389,N_9063);
nand U10664 (N_10664,N_8372,N_9657);
xnor U10665 (N_10665,N_8920,N_8267);
nand U10666 (N_10666,N_9069,N_9692);
nand U10667 (N_10667,N_9961,N_8931);
nor U10668 (N_10668,N_9143,N_8597);
and U10669 (N_10669,N_8814,N_9315);
or U10670 (N_10670,N_8537,N_8736);
xor U10671 (N_10671,N_8709,N_9775);
nor U10672 (N_10672,N_8196,N_9348);
xnor U10673 (N_10673,N_8491,N_9538);
nand U10674 (N_10674,N_9623,N_8066);
and U10675 (N_10675,N_9578,N_8091);
and U10676 (N_10676,N_8996,N_8049);
xor U10677 (N_10677,N_9177,N_9599);
nor U10678 (N_10678,N_9860,N_8229);
and U10679 (N_10679,N_8070,N_9066);
or U10680 (N_10680,N_9289,N_8499);
xor U10681 (N_10681,N_8408,N_8799);
nor U10682 (N_10682,N_9959,N_8957);
or U10683 (N_10683,N_9808,N_8395);
xor U10684 (N_10684,N_9472,N_8521);
and U10685 (N_10685,N_9058,N_8021);
and U10686 (N_10686,N_8019,N_8475);
nand U10687 (N_10687,N_9739,N_8037);
or U10688 (N_10688,N_9102,N_9777);
xnor U10689 (N_10689,N_8353,N_8144);
nor U10690 (N_10690,N_8779,N_9601);
or U10691 (N_10691,N_9990,N_8216);
nor U10692 (N_10692,N_9641,N_8724);
nor U10693 (N_10693,N_8323,N_9002);
or U10694 (N_10694,N_8524,N_8947);
nor U10695 (N_10695,N_9103,N_8951);
xnor U10696 (N_10696,N_8664,N_9812);
nand U10697 (N_10697,N_9949,N_8807);
nor U10698 (N_10698,N_9513,N_9725);
nand U10699 (N_10699,N_8240,N_8983);
nor U10700 (N_10700,N_8443,N_9946);
and U10701 (N_10701,N_9483,N_8915);
xnor U10702 (N_10702,N_8939,N_9729);
or U10703 (N_10703,N_9981,N_9546);
xor U10704 (N_10704,N_9372,N_8977);
xnor U10705 (N_10705,N_8676,N_8754);
and U10706 (N_10706,N_8030,N_8689);
xor U10707 (N_10707,N_9438,N_9097);
and U10708 (N_10708,N_8639,N_9068);
xnor U10709 (N_10709,N_9040,N_8068);
or U10710 (N_10710,N_8176,N_8375);
nor U10711 (N_10711,N_9457,N_9576);
nand U10712 (N_10712,N_9621,N_9635);
nor U10713 (N_10713,N_8859,N_9888);
nor U10714 (N_10714,N_8722,N_8265);
xnor U10715 (N_10715,N_9408,N_8948);
xnor U10716 (N_10716,N_8810,N_9325);
nand U10717 (N_10717,N_8193,N_8451);
xor U10718 (N_10718,N_9277,N_9081);
nand U10719 (N_10719,N_9233,N_9474);
or U10720 (N_10720,N_8061,N_9268);
and U10721 (N_10721,N_9322,N_8269);
nor U10722 (N_10722,N_9682,N_8490);
and U10723 (N_10723,N_8659,N_9263);
and U10724 (N_10724,N_9290,N_9568);
xor U10725 (N_10725,N_9772,N_9175);
or U10726 (N_10726,N_8772,N_8838);
xnor U10727 (N_10727,N_8462,N_9528);
nor U10728 (N_10728,N_8348,N_8846);
xor U10729 (N_10729,N_8982,N_8233);
nor U10730 (N_10730,N_9936,N_8303);
and U10731 (N_10731,N_9963,N_9032);
xnor U10732 (N_10732,N_9158,N_9491);
nand U10733 (N_10733,N_9706,N_8847);
nand U10734 (N_10734,N_8925,N_8588);
xor U10735 (N_10735,N_9678,N_8851);
nor U10736 (N_10736,N_8177,N_9830);
and U10737 (N_10737,N_9061,N_8620);
or U10738 (N_10738,N_8819,N_9878);
xnor U10739 (N_10739,N_8885,N_9718);
or U10740 (N_10740,N_9256,N_9533);
nor U10741 (N_10741,N_8841,N_8359);
or U10742 (N_10742,N_8710,N_9200);
xor U10743 (N_10743,N_8145,N_8711);
and U10744 (N_10744,N_8612,N_8663);
xnor U10745 (N_10745,N_9387,N_8614);
nor U10746 (N_10746,N_9261,N_9920);
and U10747 (N_10747,N_8053,N_8771);
nor U10748 (N_10748,N_8611,N_8444);
nand U10749 (N_10749,N_8298,N_9997);
and U10750 (N_10750,N_9722,N_9485);
nor U10751 (N_10751,N_8645,N_9606);
xor U10752 (N_10752,N_9088,N_9082);
nor U10753 (N_10753,N_9171,N_8434);
xor U10754 (N_10754,N_9843,N_8264);
xnor U10755 (N_10755,N_8454,N_8892);
nand U10756 (N_10756,N_8848,N_8798);
xor U10757 (N_10757,N_9179,N_9971);
nor U10758 (N_10758,N_9443,N_8313);
and U10759 (N_10759,N_8973,N_8899);
or U10760 (N_10760,N_8631,N_9795);
and U10761 (N_10761,N_8778,N_9213);
xnor U10762 (N_10762,N_9262,N_9269);
xnor U10763 (N_10763,N_8975,N_9347);
xor U10764 (N_10764,N_8131,N_9897);
nand U10765 (N_10765,N_8632,N_8022);
nand U10766 (N_10766,N_8130,N_9463);
nand U10767 (N_10767,N_8396,N_8248);
nor U10768 (N_10768,N_8600,N_8766);
and U10769 (N_10769,N_8578,N_8565);
nor U10770 (N_10770,N_8194,N_8943);
and U10771 (N_10771,N_8857,N_8231);
and U10772 (N_10772,N_9838,N_9336);
and U10773 (N_10773,N_9449,N_9566);
or U10774 (N_10774,N_9649,N_8413);
or U10775 (N_10775,N_8912,N_9219);
nand U10776 (N_10776,N_8322,N_9796);
nand U10777 (N_10777,N_9023,N_9871);
and U10778 (N_10778,N_8649,N_9991);
nand U10779 (N_10779,N_8739,N_8213);
xor U10780 (N_10780,N_8274,N_9674);
nor U10781 (N_10781,N_9412,N_9204);
or U10782 (N_10782,N_9003,N_8875);
nand U10783 (N_10783,N_9770,N_9744);
or U10784 (N_10784,N_9846,N_8411);
and U10785 (N_10785,N_9094,N_9980);
nor U10786 (N_10786,N_9848,N_8345);
nand U10787 (N_10787,N_8414,N_9561);
xnor U10788 (N_10788,N_8402,N_8230);
nor U10789 (N_10789,N_8525,N_9899);
nor U10790 (N_10790,N_8555,N_8288);
xnor U10791 (N_10791,N_9089,N_9826);
or U10792 (N_10792,N_9011,N_9964);
nand U10793 (N_10793,N_9918,N_9448);
xor U10794 (N_10794,N_8666,N_8294);
nor U10795 (N_10795,N_9667,N_9655);
xnor U10796 (N_10796,N_9415,N_9255);
nand U10797 (N_10797,N_9025,N_8970);
and U10798 (N_10798,N_9543,N_9738);
and U10799 (N_10799,N_8173,N_9461);
and U10800 (N_10800,N_9712,N_9890);
xnor U10801 (N_10801,N_9996,N_9150);
nand U10802 (N_10802,N_8377,N_9815);
nor U10803 (N_10803,N_8453,N_9504);
or U10804 (N_10804,N_8232,N_9519);
nor U10805 (N_10805,N_9321,N_8569);
and U10806 (N_10806,N_8956,N_8020);
or U10807 (N_10807,N_8486,N_9604);
and U10808 (N_10808,N_9283,N_9342);
nand U10809 (N_10809,N_8312,N_9361);
nor U10810 (N_10810,N_9559,N_9583);
and U10811 (N_10811,N_8084,N_8902);
xnor U10812 (N_10812,N_8602,N_9306);
or U10813 (N_10813,N_8284,N_9421);
and U10814 (N_10814,N_8039,N_9488);
or U10815 (N_10815,N_8381,N_8279);
and U10816 (N_10816,N_9446,N_9856);
and U10817 (N_10817,N_9379,N_8812);
and U10818 (N_10818,N_9416,N_8672);
xnor U10819 (N_10819,N_9301,N_8508);
xnor U10820 (N_10820,N_8007,N_9172);
nand U10821 (N_10821,N_8122,N_9064);
nand U10822 (N_10822,N_9832,N_8813);
and U10823 (N_10823,N_9853,N_9512);
nand U10824 (N_10824,N_9666,N_9189);
or U10825 (N_10825,N_8593,N_8874);
nor U10826 (N_10826,N_9282,N_8051);
and U10827 (N_10827,N_8088,N_8355);
nor U10828 (N_10828,N_9072,N_8680);
nor U10829 (N_10829,N_9778,N_9090);
xor U10830 (N_10830,N_8067,N_9517);
nor U10831 (N_10831,N_9675,N_8746);
nand U10832 (N_10832,N_8041,N_8696);
nor U10833 (N_10833,N_9239,N_8795);
and U10834 (N_10834,N_8316,N_8087);
nor U10835 (N_10835,N_9769,N_8518);
and U10836 (N_10836,N_8523,N_9101);
xnor U10837 (N_10837,N_8483,N_9969);
nor U10838 (N_10838,N_9317,N_9765);
nor U10839 (N_10839,N_9929,N_9565);
and U10840 (N_10840,N_8424,N_9123);
or U10841 (N_10841,N_8456,N_8502);
nand U10842 (N_10842,N_9916,N_8105);
nor U10843 (N_10843,N_9828,N_9382);
or U10844 (N_10844,N_8513,N_8347);
nand U10845 (N_10845,N_9841,N_8005);
or U10846 (N_10846,N_8350,N_8698);
nand U10847 (N_10847,N_9763,N_8195);
or U10848 (N_10848,N_9460,N_9822);
and U10849 (N_10849,N_8786,N_9885);
nand U10850 (N_10850,N_9972,N_9431);
xnor U10851 (N_10851,N_8566,N_9761);
and U10852 (N_10852,N_8001,N_9766);
nor U10853 (N_10853,N_8114,N_8753);
and U10854 (N_10854,N_9548,N_8767);
nand U10855 (N_10855,N_9994,N_8025);
xor U10856 (N_10856,N_9225,N_8530);
or U10857 (N_10857,N_8147,N_8010);
xor U10858 (N_10858,N_9426,N_9903);
and U10859 (N_10859,N_8653,N_9419);
nand U10860 (N_10860,N_9589,N_9595);
nor U10861 (N_10861,N_8327,N_8459);
xor U10862 (N_10862,N_9930,N_8655);
or U10863 (N_10863,N_8175,N_8618);
or U10864 (N_10864,N_9544,N_9602);
nand U10865 (N_10865,N_9781,N_8332);
nor U10866 (N_10866,N_8665,N_9429);
or U10867 (N_10867,N_9499,N_9407);
and U10868 (N_10868,N_9351,N_9402);
xor U10869 (N_10869,N_8601,N_8774);
and U10870 (N_10870,N_8978,N_9229);
and U10871 (N_10871,N_9870,N_8369);
nand U10872 (N_10872,N_8503,N_9093);
nand U10873 (N_10873,N_8344,N_9246);
xnor U10874 (N_10874,N_8990,N_9817);
xnor U10875 (N_10875,N_9679,N_9653);
nor U10876 (N_10876,N_8166,N_8737);
or U10877 (N_10877,N_8151,N_9490);
xnor U10878 (N_10878,N_9798,N_8608);
xor U10879 (N_10879,N_8871,N_8304);
nand U10880 (N_10880,N_8804,N_9222);
or U10881 (N_10881,N_9840,N_8609);
or U10882 (N_10882,N_9119,N_8660);
xnor U10883 (N_10883,N_8533,N_8627);
xnor U10884 (N_10884,N_8512,N_8797);
or U10885 (N_10885,N_9323,N_8991);
nand U10886 (N_10886,N_8638,N_9582);
nand U10887 (N_10887,N_8564,N_8843);
and U10888 (N_10888,N_8567,N_8623);
and U10889 (N_10889,N_9688,N_8905);
and U10890 (N_10890,N_8241,N_8464);
nand U10891 (N_10891,N_9567,N_8747);
or U10892 (N_10892,N_8692,N_9197);
nand U10893 (N_10893,N_9724,N_9362);
and U10894 (N_10894,N_9052,N_8081);
nand U10895 (N_10895,N_9610,N_8146);
or U10896 (N_10896,N_9503,N_8445);
and U10897 (N_10897,N_9435,N_9332);
xor U10898 (N_10898,N_8510,N_9240);
xnor U10899 (N_10899,N_8707,N_9481);
nand U10900 (N_10900,N_8078,N_8378);
nand U10901 (N_10901,N_9719,N_8038);
or U10902 (N_10902,N_9721,N_8900);
or U10903 (N_10903,N_9112,N_8376);
nand U10904 (N_10904,N_8842,N_9509);
nor U10905 (N_10905,N_9898,N_9149);
or U10906 (N_10906,N_9586,N_9414);
nor U10907 (N_10907,N_8497,N_8143);
and U10908 (N_10908,N_9510,N_8641);
nand U10909 (N_10909,N_9502,N_9669);
and U10910 (N_10910,N_8595,N_9590);
nor U10911 (N_10911,N_9459,N_9212);
or U10912 (N_10912,N_9780,N_9267);
xor U10913 (N_10913,N_9527,N_8551);
nand U10914 (N_10914,N_8590,N_8236);
xor U10915 (N_10915,N_9216,N_9354);
nand U10916 (N_10916,N_9906,N_9370);
xnor U10917 (N_10917,N_9834,N_8821);
or U10918 (N_10918,N_9749,N_9705);
xnor U10919 (N_10919,N_8086,N_9259);
and U10920 (N_10920,N_9295,N_9423);
xnor U10921 (N_10921,N_8731,N_8221);
nor U10922 (N_10922,N_9156,N_8573);
or U10923 (N_10923,N_8646,N_9858);
xnor U10924 (N_10924,N_8559,N_8769);
and U10925 (N_10925,N_9516,N_8158);
or U10926 (N_10926,N_8013,N_9591);
and U10927 (N_10927,N_8425,N_8682);
or U10928 (N_10928,N_8466,N_8688);
and U10929 (N_10929,N_9131,N_9879);
or U10930 (N_10930,N_8492,N_9489);
and U10931 (N_10931,N_9708,N_9902);
xnor U10932 (N_10932,N_8124,N_8043);
or U10933 (N_10933,N_9563,N_9515);
xnor U10934 (N_10934,N_8995,N_9792);
xor U10935 (N_10935,N_8291,N_8420);
or U10936 (N_10936,N_8768,N_8695);
or U10937 (N_10937,N_9207,N_9356);
nor U10938 (N_10938,N_9099,N_8465);
nor U10939 (N_10939,N_8442,N_8540);
and U10940 (N_10940,N_9713,N_9029);
or U10941 (N_10941,N_9975,N_9145);
or U10942 (N_10942,N_9340,N_9111);
or U10943 (N_10943,N_8926,N_9750);
nor U10944 (N_10944,N_9250,N_8603);
nand U10945 (N_10945,N_8922,N_8108);
and U10946 (N_10946,N_9797,N_8405);
nand U10947 (N_10947,N_8547,N_8392);
or U10948 (N_10948,N_8974,N_9395);
nand U10949 (N_10949,N_8085,N_8891);
or U10950 (N_10950,N_8244,N_9085);
and U10951 (N_10951,N_9237,N_8959);
nand U10952 (N_10952,N_9545,N_9164);
or U10953 (N_10953,N_8441,N_8419);
nand U10954 (N_10954,N_9521,N_9613);
nor U10955 (N_10955,N_9701,N_9000);
xor U10956 (N_10956,N_9723,N_9529);
xnor U10957 (N_10957,N_8309,N_9487);
nand U10958 (N_10958,N_8209,N_8913);
or U10959 (N_10959,N_9965,N_8651);
xor U10960 (N_10960,N_8571,N_8690);
nor U10961 (N_10961,N_9592,N_9710);
nand U10962 (N_10962,N_8356,N_9371);
nor U10963 (N_10963,N_8713,N_9683);
nor U10964 (N_10964,N_9891,N_8704);
and U10965 (N_10965,N_9768,N_8447);
nor U10966 (N_10966,N_8292,N_9270);
xor U10967 (N_10967,N_8238,N_8364);
or U10968 (N_10968,N_9945,N_9707);
xnor U10969 (N_10969,N_8220,N_8092);
nor U10970 (N_10970,N_9162,N_9716);
and U10971 (N_10971,N_9386,N_9425);
or U10972 (N_10972,N_9558,N_8159);
and U10973 (N_10973,N_9836,N_8449);
or U10974 (N_10974,N_8003,N_8098);
or U10975 (N_10975,N_8479,N_8203);
nor U10976 (N_10976,N_8059,N_8998);
and U10977 (N_10977,N_8320,N_9977);
and U10978 (N_10978,N_8855,N_9293);
nand U10979 (N_10979,N_9630,N_9862);
xnor U10980 (N_10980,N_9211,N_8474);
nand U10981 (N_10981,N_9441,N_9609);
or U10982 (N_10982,N_8706,N_8374);
xor U10983 (N_10983,N_9044,N_9859);
nand U10984 (N_10984,N_8628,N_9215);
nor U10985 (N_10985,N_9877,N_9478);
nand U10986 (N_10986,N_9238,N_9911);
nor U10987 (N_10987,N_9285,N_8012);
xnor U10988 (N_10988,N_9671,N_8589);
nand U10989 (N_10989,N_9329,N_8703);
and U10990 (N_10990,N_9297,N_8927);
nand U10991 (N_10991,N_8770,N_8117);
nand U10992 (N_10992,N_9868,N_8299);
or U10993 (N_10993,N_9539,N_9557);
or U10994 (N_10994,N_8063,N_9410);
nor U10995 (N_10995,N_9668,N_8189);
xor U10996 (N_10996,N_8596,N_8501);
and U10997 (N_10997,N_9803,N_8400);
xor U10998 (N_10998,N_9344,N_9157);
nand U10999 (N_10999,N_8504,N_9437);
nor U11000 (N_11000,N_8530,N_8732);
and U11001 (N_11001,N_9660,N_8258);
and U11002 (N_11002,N_9464,N_8770);
and U11003 (N_11003,N_9470,N_9012);
or U11004 (N_11004,N_8974,N_8975);
nand U11005 (N_11005,N_8473,N_9618);
nand U11006 (N_11006,N_9166,N_9047);
or U11007 (N_11007,N_8517,N_8018);
and U11008 (N_11008,N_8737,N_8670);
and U11009 (N_11009,N_9411,N_8888);
and U11010 (N_11010,N_8393,N_9839);
nor U11011 (N_11011,N_9499,N_8759);
xor U11012 (N_11012,N_8432,N_9270);
nor U11013 (N_11013,N_8139,N_8000);
nand U11014 (N_11014,N_9707,N_9550);
and U11015 (N_11015,N_9347,N_9933);
and U11016 (N_11016,N_9656,N_8580);
xor U11017 (N_11017,N_9621,N_9536);
xnor U11018 (N_11018,N_9302,N_8582);
nand U11019 (N_11019,N_9790,N_9992);
and U11020 (N_11020,N_9852,N_8878);
nor U11021 (N_11021,N_8133,N_8181);
xor U11022 (N_11022,N_9701,N_9220);
nor U11023 (N_11023,N_9318,N_8544);
or U11024 (N_11024,N_9401,N_9975);
and U11025 (N_11025,N_9024,N_8135);
xor U11026 (N_11026,N_9874,N_8378);
and U11027 (N_11027,N_9452,N_9462);
nor U11028 (N_11028,N_8824,N_8731);
nor U11029 (N_11029,N_8992,N_9193);
nand U11030 (N_11030,N_9467,N_8798);
and U11031 (N_11031,N_9586,N_9940);
or U11032 (N_11032,N_8812,N_8330);
or U11033 (N_11033,N_8772,N_9658);
xnor U11034 (N_11034,N_8789,N_8990);
and U11035 (N_11035,N_8834,N_9591);
and U11036 (N_11036,N_9982,N_8943);
nand U11037 (N_11037,N_9545,N_8796);
nand U11038 (N_11038,N_9031,N_8947);
or U11039 (N_11039,N_9230,N_9292);
nor U11040 (N_11040,N_8290,N_9745);
nor U11041 (N_11041,N_9862,N_9086);
and U11042 (N_11042,N_9243,N_9440);
or U11043 (N_11043,N_9807,N_9801);
xor U11044 (N_11044,N_9104,N_8639);
xnor U11045 (N_11045,N_9490,N_8600);
or U11046 (N_11046,N_8092,N_8819);
nor U11047 (N_11047,N_9488,N_8209);
xor U11048 (N_11048,N_8607,N_9121);
and U11049 (N_11049,N_9524,N_9773);
and U11050 (N_11050,N_9614,N_9341);
nand U11051 (N_11051,N_8010,N_9686);
nor U11052 (N_11052,N_8213,N_9052);
nor U11053 (N_11053,N_8365,N_8868);
and U11054 (N_11054,N_9728,N_9579);
or U11055 (N_11055,N_9603,N_9421);
xor U11056 (N_11056,N_8561,N_8122);
or U11057 (N_11057,N_9486,N_9320);
nor U11058 (N_11058,N_9056,N_8232);
nor U11059 (N_11059,N_9008,N_8357);
and U11060 (N_11060,N_9643,N_8869);
nand U11061 (N_11061,N_9066,N_9980);
and U11062 (N_11062,N_8161,N_9160);
or U11063 (N_11063,N_9196,N_9957);
xor U11064 (N_11064,N_9146,N_8908);
and U11065 (N_11065,N_9905,N_9427);
nand U11066 (N_11066,N_8191,N_8662);
nand U11067 (N_11067,N_8111,N_8984);
and U11068 (N_11068,N_8754,N_9761);
or U11069 (N_11069,N_9514,N_8507);
or U11070 (N_11070,N_9604,N_8694);
or U11071 (N_11071,N_8477,N_9014);
nor U11072 (N_11072,N_8314,N_9236);
nor U11073 (N_11073,N_9088,N_9689);
nand U11074 (N_11074,N_9281,N_8688);
nand U11075 (N_11075,N_8789,N_8692);
xnor U11076 (N_11076,N_8875,N_9622);
or U11077 (N_11077,N_8722,N_9478);
xnor U11078 (N_11078,N_9265,N_8219);
and U11079 (N_11079,N_8400,N_8872);
nand U11080 (N_11080,N_9905,N_8804);
or U11081 (N_11081,N_9522,N_8431);
nor U11082 (N_11082,N_9281,N_9681);
or U11083 (N_11083,N_9753,N_8070);
nor U11084 (N_11084,N_8685,N_9342);
nand U11085 (N_11085,N_9733,N_8051);
xnor U11086 (N_11086,N_8704,N_8055);
xnor U11087 (N_11087,N_9734,N_9664);
xnor U11088 (N_11088,N_9786,N_8461);
nand U11089 (N_11089,N_8288,N_8208);
nor U11090 (N_11090,N_8509,N_9676);
nor U11091 (N_11091,N_9755,N_8293);
nor U11092 (N_11092,N_9276,N_9440);
nand U11093 (N_11093,N_8610,N_9181);
nand U11094 (N_11094,N_8006,N_8607);
or U11095 (N_11095,N_8903,N_9837);
or U11096 (N_11096,N_8506,N_8260);
nor U11097 (N_11097,N_9246,N_9268);
nor U11098 (N_11098,N_8831,N_9120);
or U11099 (N_11099,N_8375,N_9494);
xnor U11100 (N_11100,N_9903,N_9409);
nor U11101 (N_11101,N_8483,N_8234);
and U11102 (N_11102,N_9255,N_8440);
nor U11103 (N_11103,N_8321,N_8448);
and U11104 (N_11104,N_8015,N_8445);
and U11105 (N_11105,N_9810,N_9380);
and U11106 (N_11106,N_8059,N_8250);
or U11107 (N_11107,N_9621,N_9314);
nand U11108 (N_11108,N_9814,N_8070);
nand U11109 (N_11109,N_9266,N_9367);
or U11110 (N_11110,N_9971,N_9056);
nor U11111 (N_11111,N_9656,N_8885);
and U11112 (N_11112,N_9506,N_9643);
and U11113 (N_11113,N_9010,N_9380);
nand U11114 (N_11114,N_8172,N_8189);
nand U11115 (N_11115,N_8316,N_9522);
or U11116 (N_11116,N_9829,N_9254);
and U11117 (N_11117,N_8363,N_8961);
nor U11118 (N_11118,N_9343,N_8490);
xnor U11119 (N_11119,N_8467,N_8209);
nor U11120 (N_11120,N_9418,N_8389);
and U11121 (N_11121,N_9446,N_8451);
nor U11122 (N_11122,N_8301,N_8373);
xnor U11123 (N_11123,N_8560,N_9814);
nor U11124 (N_11124,N_9628,N_9432);
nand U11125 (N_11125,N_9530,N_9584);
and U11126 (N_11126,N_8918,N_9069);
xor U11127 (N_11127,N_8512,N_9168);
and U11128 (N_11128,N_9809,N_8559);
xor U11129 (N_11129,N_9556,N_9378);
nor U11130 (N_11130,N_9363,N_8281);
xnor U11131 (N_11131,N_9196,N_9150);
and U11132 (N_11132,N_8085,N_8993);
or U11133 (N_11133,N_8108,N_9691);
nor U11134 (N_11134,N_8449,N_9661);
nor U11135 (N_11135,N_8404,N_8884);
and U11136 (N_11136,N_8613,N_8133);
xnor U11137 (N_11137,N_9487,N_8856);
xnor U11138 (N_11138,N_8980,N_9490);
and U11139 (N_11139,N_8012,N_9924);
nor U11140 (N_11140,N_8308,N_9310);
nor U11141 (N_11141,N_9815,N_9313);
and U11142 (N_11142,N_9875,N_8653);
or U11143 (N_11143,N_9021,N_9713);
xnor U11144 (N_11144,N_8328,N_8545);
nand U11145 (N_11145,N_9272,N_8671);
xnor U11146 (N_11146,N_9715,N_9658);
or U11147 (N_11147,N_8013,N_8535);
and U11148 (N_11148,N_8710,N_8980);
nor U11149 (N_11149,N_9703,N_9532);
or U11150 (N_11150,N_8636,N_8547);
xor U11151 (N_11151,N_8126,N_8765);
xor U11152 (N_11152,N_8362,N_8998);
nor U11153 (N_11153,N_8560,N_9011);
and U11154 (N_11154,N_8212,N_9495);
or U11155 (N_11155,N_9720,N_8353);
nand U11156 (N_11156,N_8201,N_8110);
or U11157 (N_11157,N_8073,N_8575);
and U11158 (N_11158,N_8410,N_8305);
nor U11159 (N_11159,N_9242,N_9649);
xor U11160 (N_11160,N_8185,N_8743);
nor U11161 (N_11161,N_9734,N_8013);
nor U11162 (N_11162,N_8982,N_8091);
or U11163 (N_11163,N_8246,N_9466);
nor U11164 (N_11164,N_8540,N_8069);
xnor U11165 (N_11165,N_9623,N_8326);
and U11166 (N_11166,N_8376,N_8404);
and U11167 (N_11167,N_8404,N_8923);
or U11168 (N_11168,N_9009,N_9847);
xnor U11169 (N_11169,N_8791,N_9163);
xor U11170 (N_11170,N_9966,N_9701);
and U11171 (N_11171,N_8190,N_8055);
nor U11172 (N_11172,N_8434,N_9321);
and U11173 (N_11173,N_8900,N_9530);
or U11174 (N_11174,N_9527,N_9747);
nand U11175 (N_11175,N_8127,N_9089);
nor U11176 (N_11176,N_8250,N_8201);
nand U11177 (N_11177,N_9182,N_9177);
nor U11178 (N_11178,N_9559,N_9526);
nand U11179 (N_11179,N_9081,N_9900);
xnor U11180 (N_11180,N_8956,N_8318);
nor U11181 (N_11181,N_8626,N_8682);
nor U11182 (N_11182,N_8059,N_9814);
nor U11183 (N_11183,N_9422,N_9921);
nor U11184 (N_11184,N_9648,N_8316);
xor U11185 (N_11185,N_8573,N_9349);
and U11186 (N_11186,N_9023,N_8885);
or U11187 (N_11187,N_8727,N_8267);
and U11188 (N_11188,N_8243,N_9679);
and U11189 (N_11189,N_9365,N_8265);
nand U11190 (N_11190,N_9327,N_8665);
or U11191 (N_11191,N_8628,N_9156);
or U11192 (N_11192,N_9060,N_9580);
nor U11193 (N_11193,N_9904,N_9930);
nand U11194 (N_11194,N_8166,N_8852);
nand U11195 (N_11195,N_8398,N_8422);
nor U11196 (N_11196,N_8351,N_9785);
or U11197 (N_11197,N_8759,N_8142);
nor U11198 (N_11198,N_8635,N_9778);
xnor U11199 (N_11199,N_8803,N_9271);
and U11200 (N_11200,N_9771,N_9145);
and U11201 (N_11201,N_9369,N_9921);
xor U11202 (N_11202,N_8669,N_9979);
or U11203 (N_11203,N_9704,N_9631);
nand U11204 (N_11204,N_9669,N_8179);
xor U11205 (N_11205,N_9768,N_8825);
or U11206 (N_11206,N_9576,N_9946);
and U11207 (N_11207,N_8045,N_8881);
nor U11208 (N_11208,N_8464,N_9700);
nor U11209 (N_11209,N_8465,N_8377);
or U11210 (N_11210,N_8544,N_9651);
and U11211 (N_11211,N_8092,N_9702);
or U11212 (N_11212,N_9504,N_8333);
nor U11213 (N_11213,N_8262,N_9299);
and U11214 (N_11214,N_8142,N_9550);
nand U11215 (N_11215,N_9627,N_9686);
or U11216 (N_11216,N_8614,N_8410);
and U11217 (N_11217,N_8733,N_9838);
nor U11218 (N_11218,N_9334,N_9121);
nor U11219 (N_11219,N_8254,N_8883);
nor U11220 (N_11220,N_9145,N_9011);
xor U11221 (N_11221,N_9516,N_9073);
and U11222 (N_11222,N_8696,N_9192);
and U11223 (N_11223,N_9690,N_8779);
and U11224 (N_11224,N_9449,N_9286);
and U11225 (N_11225,N_8903,N_8468);
or U11226 (N_11226,N_8173,N_8500);
nand U11227 (N_11227,N_9162,N_9720);
and U11228 (N_11228,N_8366,N_8943);
and U11229 (N_11229,N_9940,N_9937);
xor U11230 (N_11230,N_8827,N_8099);
nand U11231 (N_11231,N_8511,N_9276);
and U11232 (N_11232,N_9732,N_8636);
and U11233 (N_11233,N_9873,N_9305);
and U11234 (N_11234,N_9181,N_9031);
xnor U11235 (N_11235,N_9375,N_8967);
nor U11236 (N_11236,N_9742,N_8191);
xor U11237 (N_11237,N_9976,N_9231);
xor U11238 (N_11238,N_8924,N_8588);
nor U11239 (N_11239,N_8839,N_8505);
nand U11240 (N_11240,N_9616,N_8606);
xnor U11241 (N_11241,N_8384,N_9503);
nor U11242 (N_11242,N_8422,N_9199);
nor U11243 (N_11243,N_8702,N_9518);
xnor U11244 (N_11244,N_8812,N_8584);
or U11245 (N_11245,N_8115,N_9397);
and U11246 (N_11246,N_9321,N_9642);
nand U11247 (N_11247,N_8258,N_8521);
and U11248 (N_11248,N_8705,N_8685);
or U11249 (N_11249,N_8156,N_9504);
nor U11250 (N_11250,N_8716,N_8519);
and U11251 (N_11251,N_8940,N_9283);
nor U11252 (N_11252,N_9261,N_8445);
and U11253 (N_11253,N_8671,N_8050);
xnor U11254 (N_11254,N_9000,N_9452);
or U11255 (N_11255,N_8293,N_9959);
or U11256 (N_11256,N_8918,N_9525);
or U11257 (N_11257,N_8794,N_9827);
xnor U11258 (N_11258,N_9504,N_9304);
xnor U11259 (N_11259,N_9965,N_9349);
nor U11260 (N_11260,N_9046,N_8319);
and U11261 (N_11261,N_9006,N_8444);
and U11262 (N_11262,N_8695,N_9539);
and U11263 (N_11263,N_9400,N_8085);
nand U11264 (N_11264,N_9553,N_9588);
nor U11265 (N_11265,N_8403,N_8297);
xor U11266 (N_11266,N_8546,N_9374);
nor U11267 (N_11267,N_8917,N_9721);
nand U11268 (N_11268,N_9200,N_9352);
or U11269 (N_11269,N_9928,N_9078);
nor U11270 (N_11270,N_9538,N_9757);
nor U11271 (N_11271,N_8618,N_8811);
nor U11272 (N_11272,N_9446,N_8377);
nor U11273 (N_11273,N_9853,N_9115);
nor U11274 (N_11274,N_8277,N_9046);
nor U11275 (N_11275,N_8690,N_8496);
nand U11276 (N_11276,N_9559,N_9201);
nand U11277 (N_11277,N_9849,N_8001);
nand U11278 (N_11278,N_8748,N_8282);
and U11279 (N_11279,N_8616,N_8544);
or U11280 (N_11280,N_8197,N_8352);
nor U11281 (N_11281,N_9197,N_8568);
or U11282 (N_11282,N_8731,N_8359);
nand U11283 (N_11283,N_8283,N_8396);
and U11284 (N_11284,N_9680,N_9439);
xnor U11285 (N_11285,N_8168,N_9494);
nor U11286 (N_11286,N_9361,N_8826);
nor U11287 (N_11287,N_8660,N_8510);
and U11288 (N_11288,N_8614,N_8848);
xnor U11289 (N_11289,N_8706,N_8289);
or U11290 (N_11290,N_8738,N_9676);
nor U11291 (N_11291,N_8556,N_9410);
and U11292 (N_11292,N_8118,N_8405);
and U11293 (N_11293,N_9136,N_8897);
nor U11294 (N_11294,N_9105,N_8657);
or U11295 (N_11295,N_9613,N_9549);
or U11296 (N_11296,N_9716,N_9505);
or U11297 (N_11297,N_9574,N_9847);
nand U11298 (N_11298,N_9813,N_8087);
and U11299 (N_11299,N_8895,N_8566);
nor U11300 (N_11300,N_9708,N_8492);
nand U11301 (N_11301,N_9846,N_8048);
or U11302 (N_11302,N_9341,N_9855);
and U11303 (N_11303,N_9648,N_8943);
and U11304 (N_11304,N_9850,N_8343);
or U11305 (N_11305,N_8939,N_9781);
nand U11306 (N_11306,N_9447,N_9310);
or U11307 (N_11307,N_8702,N_8221);
or U11308 (N_11308,N_8399,N_9286);
and U11309 (N_11309,N_8904,N_8872);
nor U11310 (N_11310,N_9127,N_9853);
or U11311 (N_11311,N_9029,N_8853);
nand U11312 (N_11312,N_9948,N_9906);
and U11313 (N_11313,N_9742,N_9430);
nand U11314 (N_11314,N_9063,N_8380);
xnor U11315 (N_11315,N_9135,N_8743);
xnor U11316 (N_11316,N_8347,N_9183);
nor U11317 (N_11317,N_8211,N_8786);
or U11318 (N_11318,N_8060,N_9306);
xnor U11319 (N_11319,N_9787,N_8898);
and U11320 (N_11320,N_9808,N_9346);
and U11321 (N_11321,N_8916,N_8903);
nor U11322 (N_11322,N_8346,N_8947);
or U11323 (N_11323,N_8916,N_8148);
nand U11324 (N_11324,N_8943,N_9305);
nor U11325 (N_11325,N_8480,N_8962);
nor U11326 (N_11326,N_9222,N_8078);
or U11327 (N_11327,N_9994,N_8623);
or U11328 (N_11328,N_9936,N_8985);
xnor U11329 (N_11329,N_9327,N_8924);
nor U11330 (N_11330,N_8628,N_9095);
or U11331 (N_11331,N_8749,N_8953);
and U11332 (N_11332,N_8571,N_9891);
xnor U11333 (N_11333,N_8857,N_8239);
or U11334 (N_11334,N_9560,N_8611);
nor U11335 (N_11335,N_8424,N_9050);
xor U11336 (N_11336,N_9660,N_9110);
nor U11337 (N_11337,N_9904,N_9085);
nand U11338 (N_11338,N_9104,N_9764);
nand U11339 (N_11339,N_9919,N_9988);
nand U11340 (N_11340,N_8704,N_8527);
and U11341 (N_11341,N_8806,N_9380);
or U11342 (N_11342,N_9448,N_8238);
nor U11343 (N_11343,N_9012,N_9477);
or U11344 (N_11344,N_9929,N_8274);
nand U11345 (N_11345,N_8698,N_9543);
and U11346 (N_11346,N_9929,N_9073);
xnor U11347 (N_11347,N_9072,N_8844);
and U11348 (N_11348,N_9416,N_9829);
or U11349 (N_11349,N_8537,N_8109);
nor U11350 (N_11350,N_8087,N_8878);
and U11351 (N_11351,N_9380,N_8098);
nor U11352 (N_11352,N_9127,N_9774);
or U11353 (N_11353,N_9972,N_8841);
nor U11354 (N_11354,N_8470,N_9225);
nor U11355 (N_11355,N_9086,N_9951);
nor U11356 (N_11356,N_8895,N_9211);
and U11357 (N_11357,N_8144,N_8491);
nor U11358 (N_11358,N_8112,N_8946);
or U11359 (N_11359,N_9230,N_9378);
xor U11360 (N_11360,N_8266,N_9544);
xnor U11361 (N_11361,N_9391,N_9720);
xor U11362 (N_11362,N_8906,N_9165);
and U11363 (N_11363,N_9641,N_9955);
nand U11364 (N_11364,N_9026,N_8470);
and U11365 (N_11365,N_9122,N_8613);
xnor U11366 (N_11366,N_9370,N_9474);
nor U11367 (N_11367,N_9391,N_9529);
xnor U11368 (N_11368,N_9370,N_9549);
or U11369 (N_11369,N_8092,N_9439);
nand U11370 (N_11370,N_9399,N_8144);
nand U11371 (N_11371,N_9347,N_8130);
and U11372 (N_11372,N_8967,N_9579);
nand U11373 (N_11373,N_8349,N_9228);
and U11374 (N_11374,N_9019,N_9738);
nand U11375 (N_11375,N_9282,N_8077);
xor U11376 (N_11376,N_9330,N_9951);
and U11377 (N_11377,N_8853,N_8313);
xnor U11378 (N_11378,N_8886,N_9956);
and U11379 (N_11379,N_8575,N_8559);
and U11380 (N_11380,N_8480,N_8045);
or U11381 (N_11381,N_9724,N_9772);
nor U11382 (N_11382,N_8030,N_8477);
and U11383 (N_11383,N_8095,N_9604);
xnor U11384 (N_11384,N_9174,N_9201);
and U11385 (N_11385,N_8312,N_9251);
nor U11386 (N_11386,N_9149,N_8698);
nor U11387 (N_11387,N_9469,N_9438);
xor U11388 (N_11388,N_8917,N_9285);
nand U11389 (N_11389,N_9882,N_9434);
nor U11390 (N_11390,N_9926,N_8809);
or U11391 (N_11391,N_9657,N_8257);
and U11392 (N_11392,N_8291,N_8247);
nand U11393 (N_11393,N_9877,N_9997);
and U11394 (N_11394,N_9467,N_9055);
and U11395 (N_11395,N_9163,N_8306);
and U11396 (N_11396,N_8575,N_9590);
and U11397 (N_11397,N_8392,N_8505);
or U11398 (N_11398,N_9400,N_8802);
nand U11399 (N_11399,N_8414,N_8764);
and U11400 (N_11400,N_9585,N_9990);
xor U11401 (N_11401,N_9067,N_9859);
or U11402 (N_11402,N_8837,N_9936);
xnor U11403 (N_11403,N_8872,N_8456);
and U11404 (N_11404,N_8932,N_9076);
nand U11405 (N_11405,N_8720,N_8481);
nand U11406 (N_11406,N_8116,N_9637);
xnor U11407 (N_11407,N_8203,N_9370);
nand U11408 (N_11408,N_9254,N_8611);
or U11409 (N_11409,N_8325,N_8599);
or U11410 (N_11410,N_9485,N_9867);
nor U11411 (N_11411,N_8912,N_8618);
and U11412 (N_11412,N_9011,N_8991);
nor U11413 (N_11413,N_9284,N_9851);
or U11414 (N_11414,N_8256,N_9624);
nor U11415 (N_11415,N_8079,N_9608);
nor U11416 (N_11416,N_8723,N_9979);
nor U11417 (N_11417,N_8603,N_9127);
xor U11418 (N_11418,N_8559,N_8458);
xnor U11419 (N_11419,N_8259,N_9755);
nor U11420 (N_11420,N_9437,N_8005);
or U11421 (N_11421,N_9011,N_9420);
nand U11422 (N_11422,N_9922,N_9183);
and U11423 (N_11423,N_9102,N_9321);
xnor U11424 (N_11424,N_8853,N_9043);
nor U11425 (N_11425,N_9926,N_9562);
nor U11426 (N_11426,N_8137,N_9749);
nand U11427 (N_11427,N_8346,N_9721);
nor U11428 (N_11428,N_9718,N_9527);
or U11429 (N_11429,N_8165,N_9042);
nor U11430 (N_11430,N_9543,N_9989);
xor U11431 (N_11431,N_9200,N_9424);
nand U11432 (N_11432,N_9237,N_8692);
xor U11433 (N_11433,N_8446,N_9715);
nor U11434 (N_11434,N_9282,N_8180);
or U11435 (N_11435,N_8588,N_9437);
nor U11436 (N_11436,N_8382,N_9199);
or U11437 (N_11437,N_9963,N_8926);
nand U11438 (N_11438,N_8674,N_8259);
xor U11439 (N_11439,N_9849,N_9408);
xnor U11440 (N_11440,N_9110,N_8807);
xnor U11441 (N_11441,N_9513,N_9160);
nor U11442 (N_11442,N_8123,N_8679);
xnor U11443 (N_11443,N_8089,N_9528);
nor U11444 (N_11444,N_8305,N_8408);
xor U11445 (N_11445,N_9099,N_9835);
nand U11446 (N_11446,N_9779,N_9113);
nor U11447 (N_11447,N_8754,N_8272);
xnor U11448 (N_11448,N_9152,N_9491);
nor U11449 (N_11449,N_9128,N_8622);
and U11450 (N_11450,N_8230,N_9202);
xnor U11451 (N_11451,N_8976,N_9125);
xnor U11452 (N_11452,N_8860,N_9595);
nor U11453 (N_11453,N_9607,N_8241);
nor U11454 (N_11454,N_9859,N_9228);
or U11455 (N_11455,N_9442,N_9407);
and U11456 (N_11456,N_9336,N_8423);
nor U11457 (N_11457,N_9677,N_9642);
nand U11458 (N_11458,N_8553,N_9244);
or U11459 (N_11459,N_8537,N_8925);
nor U11460 (N_11460,N_8628,N_9528);
and U11461 (N_11461,N_8040,N_9733);
nand U11462 (N_11462,N_9452,N_9235);
or U11463 (N_11463,N_9600,N_8915);
xnor U11464 (N_11464,N_9096,N_8709);
nand U11465 (N_11465,N_8324,N_9823);
nand U11466 (N_11466,N_8869,N_8237);
or U11467 (N_11467,N_9690,N_8273);
or U11468 (N_11468,N_8192,N_9959);
or U11469 (N_11469,N_8200,N_8476);
nand U11470 (N_11470,N_8833,N_9487);
or U11471 (N_11471,N_9210,N_8151);
xnor U11472 (N_11472,N_8160,N_8625);
nor U11473 (N_11473,N_8939,N_9201);
nand U11474 (N_11474,N_8014,N_9714);
and U11475 (N_11475,N_9781,N_8255);
nor U11476 (N_11476,N_8136,N_9290);
and U11477 (N_11477,N_8938,N_9235);
and U11478 (N_11478,N_8633,N_9448);
and U11479 (N_11479,N_9305,N_9516);
nand U11480 (N_11480,N_8714,N_9749);
xnor U11481 (N_11481,N_9380,N_8517);
xor U11482 (N_11482,N_9854,N_9907);
or U11483 (N_11483,N_8019,N_9748);
or U11484 (N_11484,N_8403,N_9472);
nand U11485 (N_11485,N_9468,N_9153);
and U11486 (N_11486,N_9294,N_9174);
and U11487 (N_11487,N_8037,N_9507);
and U11488 (N_11488,N_8219,N_9395);
nand U11489 (N_11489,N_8343,N_9440);
and U11490 (N_11490,N_9056,N_8894);
xnor U11491 (N_11491,N_9746,N_8013);
and U11492 (N_11492,N_9383,N_8222);
or U11493 (N_11493,N_8052,N_9493);
and U11494 (N_11494,N_9187,N_9976);
xor U11495 (N_11495,N_8622,N_9864);
nand U11496 (N_11496,N_8275,N_9515);
or U11497 (N_11497,N_9082,N_9714);
or U11498 (N_11498,N_9211,N_8125);
xor U11499 (N_11499,N_8650,N_8242);
and U11500 (N_11500,N_9181,N_9771);
nor U11501 (N_11501,N_8292,N_8488);
nor U11502 (N_11502,N_8315,N_9408);
and U11503 (N_11503,N_8876,N_9913);
nor U11504 (N_11504,N_8392,N_8681);
or U11505 (N_11505,N_9392,N_9912);
and U11506 (N_11506,N_8676,N_8790);
and U11507 (N_11507,N_8047,N_8812);
or U11508 (N_11508,N_9317,N_8354);
xnor U11509 (N_11509,N_9728,N_8161);
xor U11510 (N_11510,N_8248,N_9477);
nand U11511 (N_11511,N_9805,N_8086);
and U11512 (N_11512,N_9449,N_9443);
xor U11513 (N_11513,N_9428,N_9058);
nand U11514 (N_11514,N_9663,N_9378);
nand U11515 (N_11515,N_8869,N_8749);
or U11516 (N_11516,N_8798,N_9570);
xnor U11517 (N_11517,N_9490,N_8882);
and U11518 (N_11518,N_8612,N_9634);
xor U11519 (N_11519,N_8776,N_8731);
nor U11520 (N_11520,N_9011,N_9472);
or U11521 (N_11521,N_9236,N_9850);
or U11522 (N_11522,N_9599,N_9232);
nand U11523 (N_11523,N_9177,N_8797);
nor U11524 (N_11524,N_9911,N_8606);
xnor U11525 (N_11525,N_8624,N_8026);
and U11526 (N_11526,N_8860,N_9314);
or U11527 (N_11527,N_9718,N_8307);
or U11528 (N_11528,N_8864,N_9912);
or U11529 (N_11529,N_9426,N_8630);
nand U11530 (N_11530,N_9104,N_9994);
xnor U11531 (N_11531,N_9811,N_9415);
nand U11532 (N_11532,N_8269,N_9250);
or U11533 (N_11533,N_8484,N_9690);
xnor U11534 (N_11534,N_8380,N_8850);
xor U11535 (N_11535,N_9688,N_8293);
xnor U11536 (N_11536,N_8503,N_9639);
nand U11537 (N_11537,N_9212,N_8433);
xor U11538 (N_11538,N_8558,N_8854);
nand U11539 (N_11539,N_8818,N_8276);
xnor U11540 (N_11540,N_9238,N_9000);
or U11541 (N_11541,N_9508,N_9377);
and U11542 (N_11542,N_9468,N_9897);
and U11543 (N_11543,N_8198,N_9651);
nand U11544 (N_11544,N_9768,N_8826);
and U11545 (N_11545,N_8955,N_8170);
or U11546 (N_11546,N_9062,N_8884);
xnor U11547 (N_11547,N_9670,N_9634);
or U11548 (N_11548,N_9493,N_9731);
nor U11549 (N_11549,N_8562,N_9235);
nand U11550 (N_11550,N_8954,N_9072);
nand U11551 (N_11551,N_8501,N_8647);
nand U11552 (N_11552,N_8043,N_8064);
or U11553 (N_11553,N_9045,N_9078);
nand U11554 (N_11554,N_8732,N_8791);
and U11555 (N_11555,N_9368,N_8893);
nand U11556 (N_11556,N_9351,N_8079);
nand U11557 (N_11557,N_9995,N_8670);
nand U11558 (N_11558,N_8959,N_9094);
or U11559 (N_11559,N_9721,N_9230);
and U11560 (N_11560,N_8385,N_9668);
nand U11561 (N_11561,N_9660,N_9313);
or U11562 (N_11562,N_9789,N_9342);
or U11563 (N_11563,N_8192,N_8110);
or U11564 (N_11564,N_9118,N_8982);
and U11565 (N_11565,N_8767,N_9651);
xor U11566 (N_11566,N_8609,N_9876);
xnor U11567 (N_11567,N_8139,N_8849);
xor U11568 (N_11568,N_9085,N_9209);
nand U11569 (N_11569,N_8484,N_9917);
nand U11570 (N_11570,N_8028,N_9137);
nand U11571 (N_11571,N_9715,N_8582);
and U11572 (N_11572,N_8488,N_9544);
or U11573 (N_11573,N_9219,N_9533);
nor U11574 (N_11574,N_8454,N_8250);
or U11575 (N_11575,N_8781,N_8393);
and U11576 (N_11576,N_9046,N_9392);
nand U11577 (N_11577,N_9265,N_9887);
nand U11578 (N_11578,N_9254,N_8127);
nand U11579 (N_11579,N_8762,N_9802);
xnor U11580 (N_11580,N_9141,N_9574);
nand U11581 (N_11581,N_8554,N_9026);
or U11582 (N_11582,N_9921,N_8461);
xor U11583 (N_11583,N_9564,N_8698);
nand U11584 (N_11584,N_8403,N_8811);
nor U11585 (N_11585,N_8478,N_9385);
xnor U11586 (N_11586,N_8386,N_8740);
nand U11587 (N_11587,N_8825,N_8553);
nor U11588 (N_11588,N_9071,N_9798);
nor U11589 (N_11589,N_8622,N_9848);
or U11590 (N_11590,N_8075,N_8168);
and U11591 (N_11591,N_8861,N_9819);
and U11592 (N_11592,N_9861,N_9937);
or U11593 (N_11593,N_9241,N_8774);
or U11594 (N_11594,N_8314,N_8850);
nand U11595 (N_11595,N_9117,N_8093);
or U11596 (N_11596,N_9808,N_8897);
nor U11597 (N_11597,N_9175,N_9407);
nor U11598 (N_11598,N_9067,N_8421);
xor U11599 (N_11599,N_8125,N_8420);
or U11600 (N_11600,N_8745,N_8696);
or U11601 (N_11601,N_9053,N_8539);
and U11602 (N_11602,N_8188,N_9389);
nor U11603 (N_11603,N_8570,N_8916);
nor U11604 (N_11604,N_9837,N_8802);
xnor U11605 (N_11605,N_8339,N_9129);
nor U11606 (N_11606,N_9602,N_9825);
nand U11607 (N_11607,N_9111,N_8239);
nand U11608 (N_11608,N_8446,N_8465);
or U11609 (N_11609,N_8236,N_9717);
and U11610 (N_11610,N_9789,N_8758);
nand U11611 (N_11611,N_8641,N_8051);
nor U11612 (N_11612,N_8449,N_9290);
and U11613 (N_11613,N_9600,N_8768);
xor U11614 (N_11614,N_8327,N_8643);
xor U11615 (N_11615,N_9796,N_9459);
or U11616 (N_11616,N_9973,N_9504);
or U11617 (N_11617,N_8936,N_8767);
xor U11618 (N_11618,N_9373,N_9635);
nor U11619 (N_11619,N_9017,N_8825);
nor U11620 (N_11620,N_8364,N_9346);
or U11621 (N_11621,N_9339,N_9126);
nand U11622 (N_11622,N_8535,N_8078);
nand U11623 (N_11623,N_9944,N_9049);
nor U11624 (N_11624,N_8460,N_9409);
nor U11625 (N_11625,N_9883,N_8820);
and U11626 (N_11626,N_9830,N_8877);
xor U11627 (N_11627,N_8845,N_9474);
xor U11628 (N_11628,N_8628,N_9767);
nor U11629 (N_11629,N_9083,N_9959);
nand U11630 (N_11630,N_8853,N_8964);
or U11631 (N_11631,N_9535,N_8752);
nand U11632 (N_11632,N_8933,N_8970);
or U11633 (N_11633,N_8236,N_9683);
or U11634 (N_11634,N_8069,N_8364);
nand U11635 (N_11635,N_8699,N_8100);
or U11636 (N_11636,N_8421,N_9056);
nand U11637 (N_11637,N_9164,N_9918);
xor U11638 (N_11638,N_9802,N_9996);
and U11639 (N_11639,N_9388,N_9881);
nor U11640 (N_11640,N_9344,N_8806);
and U11641 (N_11641,N_9596,N_9567);
nand U11642 (N_11642,N_8206,N_8511);
xnor U11643 (N_11643,N_9507,N_9081);
or U11644 (N_11644,N_9321,N_9742);
xnor U11645 (N_11645,N_9170,N_8298);
nor U11646 (N_11646,N_8605,N_8896);
or U11647 (N_11647,N_9669,N_8308);
nor U11648 (N_11648,N_9086,N_9114);
xor U11649 (N_11649,N_8098,N_8007);
nand U11650 (N_11650,N_8679,N_9641);
xnor U11651 (N_11651,N_8490,N_8374);
xor U11652 (N_11652,N_9241,N_8643);
or U11653 (N_11653,N_8038,N_9914);
nand U11654 (N_11654,N_8290,N_8259);
nand U11655 (N_11655,N_8328,N_8800);
xor U11656 (N_11656,N_8613,N_9642);
nand U11657 (N_11657,N_8848,N_8166);
or U11658 (N_11658,N_8926,N_8479);
and U11659 (N_11659,N_8478,N_8130);
xor U11660 (N_11660,N_8757,N_8570);
nor U11661 (N_11661,N_9729,N_8345);
xor U11662 (N_11662,N_9431,N_9954);
or U11663 (N_11663,N_9131,N_9802);
or U11664 (N_11664,N_9606,N_9419);
nand U11665 (N_11665,N_8268,N_8685);
or U11666 (N_11666,N_9430,N_9789);
nor U11667 (N_11667,N_9716,N_9221);
xor U11668 (N_11668,N_9109,N_9970);
xnor U11669 (N_11669,N_9630,N_9472);
xnor U11670 (N_11670,N_8228,N_8018);
and U11671 (N_11671,N_8751,N_8863);
nor U11672 (N_11672,N_8076,N_9777);
or U11673 (N_11673,N_9565,N_8906);
xor U11674 (N_11674,N_9129,N_8611);
nand U11675 (N_11675,N_8406,N_9127);
xor U11676 (N_11676,N_9931,N_8782);
nand U11677 (N_11677,N_8651,N_8248);
and U11678 (N_11678,N_9633,N_8312);
nand U11679 (N_11679,N_9208,N_8302);
and U11680 (N_11680,N_9745,N_9032);
xor U11681 (N_11681,N_9655,N_8452);
nor U11682 (N_11682,N_8610,N_9287);
nand U11683 (N_11683,N_9238,N_8038);
or U11684 (N_11684,N_8201,N_8991);
nor U11685 (N_11685,N_9916,N_8595);
nand U11686 (N_11686,N_8708,N_9479);
nand U11687 (N_11687,N_9884,N_9537);
nor U11688 (N_11688,N_8816,N_8484);
nand U11689 (N_11689,N_9167,N_9845);
and U11690 (N_11690,N_9027,N_9414);
xnor U11691 (N_11691,N_9837,N_8507);
nor U11692 (N_11692,N_9765,N_9384);
xor U11693 (N_11693,N_9908,N_8995);
nor U11694 (N_11694,N_9265,N_9633);
and U11695 (N_11695,N_9267,N_9282);
and U11696 (N_11696,N_9502,N_8104);
nand U11697 (N_11697,N_8980,N_8706);
or U11698 (N_11698,N_8147,N_8588);
xnor U11699 (N_11699,N_9720,N_8445);
xor U11700 (N_11700,N_9922,N_8651);
and U11701 (N_11701,N_9844,N_9876);
nand U11702 (N_11702,N_8104,N_8678);
xor U11703 (N_11703,N_9501,N_9505);
xnor U11704 (N_11704,N_9507,N_8563);
nand U11705 (N_11705,N_9381,N_8727);
and U11706 (N_11706,N_8738,N_8454);
nand U11707 (N_11707,N_8010,N_9173);
and U11708 (N_11708,N_8583,N_9479);
xnor U11709 (N_11709,N_8342,N_8211);
xor U11710 (N_11710,N_9505,N_8270);
nor U11711 (N_11711,N_8416,N_8606);
or U11712 (N_11712,N_8909,N_8684);
nand U11713 (N_11713,N_9683,N_9674);
or U11714 (N_11714,N_9930,N_8028);
and U11715 (N_11715,N_8590,N_8209);
and U11716 (N_11716,N_8717,N_8040);
nand U11717 (N_11717,N_8012,N_8505);
xnor U11718 (N_11718,N_9603,N_8653);
or U11719 (N_11719,N_8985,N_8159);
and U11720 (N_11720,N_8078,N_9724);
or U11721 (N_11721,N_9786,N_8404);
nand U11722 (N_11722,N_8798,N_9947);
nand U11723 (N_11723,N_9427,N_9709);
xor U11724 (N_11724,N_9301,N_9889);
or U11725 (N_11725,N_9046,N_9476);
nor U11726 (N_11726,N_8783,N_9870);
nand U11727 (N_11727,N_9750,N_9582);
xnor U11728 (N_11728,N_8404,N_8184);
or U11729 (N_11729,N_8263,N_8647);
xor U11730 (N_11730,N_8636,N_8922);
or U11731 (N_11731,N_9089,N_9696);
nor U11732 (N_11732,N_8348,N_9096);
nand U11733 (N_11733,N_9065,N_8808);
and U11734 (N_11734,N_8118,N_9014);
xor U11735 (N_11735,N_9933,N_8154);
nand U11736 (N_11736,N_9887,N_9340);
nand U11737 (N_11737,N_9909,N_8165);
nand U11738 (N_11738,N_9721,N_9060);
or U11739 (N_11739,N_9444,N_8438);
nand U11740 (N_11740,N_8435,N_9436);
and U11741 (N_11741,N_9474,N_9256);
xor U11742 (N_11742,N_9154,N_9722);
or U11743 (N_11743,N_8365,N_9009);
and U11744 (N_11744,N_9965,N_9619);
xnor U11745 (N_11745,N_9935,N_9726);
and U11746 (N_11746,N_9253,N_9471);
and U11747 (N_11747,N_8395,N_9762);
nor U11748 (N_11748,N_8521,N_8397);
nor U11749 (N_11749,N_9845,N_8473);
nand U11750 (N_11750,N_9579,N_8396);
or U11751 (N_11751,N_8804,N_8101);
or U11752 (N_11752,N_9262,N_9552);
and U11753 (N_11753,N_8884,N_8098);
or U11754 (N_11754,N_8820,N_9435);
or U11755 (N_11755,N_8605,N_9205);
or U11756 (N_11756,N_8876,N_9133);
nor U11757 (N_11757,N_9373,N_9424);
nand U11758 (N_11758,N_9949,N_8231);
nor U11759 (N_11759,N_9886,N_8390);
and U11760 (N_11760,N_8655,N_8664);
xor U11761 (N_11761,N_9828,N_9226);
xnor U11762 (N_11762,N_9710,N_9990);
and U11763 (N_11763,N_8552,N_9483);
or U11764 (N_11764,N_8120,N_9901);
nor U11765 (N_11765,N_9299,N_8437);
or U11766 (N_11766,N_9263,N_8714);
nand U11767 (N_11767,N_9682,N_8409);
nand U11768 (N_11768,N_8707,N_9281);
nand U11769 (N_11769,N_8640,N_8525);
xnor U11770 (N_11770,N_8538,N_9731);
and U11771 (N_11771,N_8329,N_8164);
xor U11772 (N_11772,N_9275,N_8406);
nand U11773 (N_11773,N_8923,N_8418);
or U11774 (N_11774,N_8583,N_9554);
xor U11775 (N_11775,N_9070,N_9002);
and U11776 (N_11776,N_8404,N_8865);
nand U11777 (N_11777,N_8148,N_8396);
and U11778 (N_11778,N_8079,N_9309);
nor U11779 (N_11779,N_9672,N_9060);
or U11780 (N_11780,N_8404,N_9787);
nand U11781 (N_11781,N_9683,N_9500);
or U11782 (N_11782,N_8197,N_9285);
and U11783 (N_11783,N_9853,N_8550);
or U11784 (N_11784,N_8437,N_8221);
or U11785 (N_11785,N_9611,N_8150);
and U11786 (N_11786,N_9910,N_8191);
or U11787 (N_11787,N_8103,N_8310);
nand U11788 (N_11788,N_9711,N_9877);
nor U11789 (N_11789,N_9706,N_9675);
nor U11790 (N_11790,N_8781,N_8523);
xor U11791 (N_11791,N_9827,N_8088);
or U11792 (N_11792,N_9858,N_8531);
or U11793 (N_11793,N_8829,N_9437);
or U11794 (N_11794,N_8435,N_9141);
or U11795 (N_11795,N_9865,N_8242);
or U11796 (N_11796,N_8243,N_9113);
xor U11797 (N_11797,N_9563,N_8288);
nand U11798 (N_11798,N_8078,N_8263);
nand U11799 (N_11799,N_8505,N_8211);
or U11800 (N_11800,N_8176,N_9569);
xor U11801 (N_11801,N_8252,N_9421);
or U11802 (N_11802,N_8013,N_8128);
nand U11803 (N_11803,N_9133,N_8537);
xor U11804 (N_11804,N_8504,N_9474);
xnor U11805 (N_11805,N_9609,N_8572);
xor U11806 (N_11806,N_9173,N_8147);
nand U11807 (N_11807,N_9211,N_9889);
or U11808 (N_11808,N_8534,N_9918);
or U11809 (N_11809,N_8905,N_8594);
or U11810 (N_11810,N_8954,N_8555);
nand U11811 (N_11811,N_8319,N_8005);
or U11812 (N_11812,N_9000,N_8732);
nand U11813 (N_11813,N_8689,N_9014);
or U11814 (N_11814,N_8224,N_9283);
and U11815 (N_11815,N_8566,N_8129);
nor U11816 (N_11816,N_8929,N_9735);
nor U11817 (N_11817,N_9278,N_8364);
nor U11818 (N_11818,N_8397,N_9001);
xnor U11819 (N_11819,N_9708,N_8082);
xor U11820 (N_11820,N_9998,N_8995);
nor U11821 (N_11821,N_8266,N_8626);
and U11822 (N_11822,N_8570,N_8960);
xor U11823 (N_11823,N_8722,N_9056);
and U11824 (N_11824,N_8484,N_9535);
or U11825 (N_11825,N_9884,N_8320);
nor U11826 (N_11826,N_8975,N_8942);
nand U11827 (N_11827,N_8331,N_8315);
nand U11828 (N_11828,N_9070,N_8642);
or U11829 (N_11829,N_9041,N_8633);
and U11830 (N_11830,N_8629,N_8734);
or U11831 (N_11831,N_9995,N_9194);
or U11832 (N_11832,N_8480,N_8973);
and U11833 (N_11833,N_9408,N_8042);
nand U11834 (N_11834,N_8309,N_8423);
nor U11835 (N_11835,N_8054,N_8781);
or U11836 (N_11836,N_9769,N_9251);
nor U11837 (N_11837,N_9828,N_9107);
or U11838 (N_11838,N_8451,N_9774);
nand U11839 (N_11839,N_9002,N_9656);
and U11840 (N_11840,N_8389,N_8783);
nand U11841 (N_11841,N_8519,N_8053);
or U11842 (N_11842,N_9373,N_9924);
nor U11843 (N_11843,N_9193,N_8670);
xor U11844 (N_11844,N_9297,N_8513);
and U11845 (N_11845,N_8419,N_8450);
nor U11846 (N_11846,N_8162,N_8605);
or U11847 (N_11847,N_9615,N_9187);
nor U11848 (N_11848,N_9088,N_8474);
or U11849 (N_11849,N_8156,N_9342);
and U11850 (N_11850,N_9682,N_8051);
nor U11851 (N_11851,N_8197,N_9741);
or U11852 (N_11852,N_8108,N_8390);
and U11853 (N_11853,N_9666,N_9507);
nand U11854 (N_11854,N_9364,N_8589);
nand U11855 (N_11855,N_8658,N_8223);
nand U11856 (N_11856,N_8061,N_8766);
and U11857 (N_11857,N_9811,N_8202);
and U11858 (N_11858,N_9520,N_9949);
nand U11859 (N_11859,N_8424,N_9538);
and U11860 (N_11860,N_9324,N_8528);
nor U11861 (N_11861,N_9323,N_8301);
xnor U11862 (N_11862,N_9459,N_8069);
or U11863 (N_11863,N_8783,N_8175);
or U11864 (N_11864,N_9380,N_8465);
nand U11865 (N_11865,N_9975,N_8925);
xor U11866 (N_11866,N_8889,N_8614);
nor U11867 (N_11867,N_9202,N_8492);
xor U11868 (N_11868,N_8175,N_9066);
nand U11869 (N_11869,N_8169,N_8780);
xnor U11870 (N_11870,N_8540,N_8505);
and U11871 (N_11871,N_8653,N_8929);
xnor U11872 (N_11872,N_8660,N_8337);
nor U11873 (N_11873,N_8571,N_8270);
or U11874 (N_11874,N_8153,N_8169);
nand U11875 (N_11875,N_9358,N_9081);
or U11876 (N_11876,N_9309,N_9299);
or U11877 (N_11877,N_9651,N_9076);
and U11878 (N_11878,N_9682,N_8633);
and U11879 (N_11879,N_8625,N_9941);
xor U11880 (N_11880,N_9621,N_8217);
nor U11881 (N_11881,N_8143,N_8002);
and U11882 (N_11882,N_9131,N_9738);
xor U11883 (N_11883,N_8645,N_8079);
or U11884 (N_11884,N_9914,N_8472);
nor U11885 (N_11885,N_9499,N_9176);
xnor U11886 (N_11886,N_9342,N_9436);
or U11887 (N_11887,N_8289,N_9806);
xnor U11888 (N_11888,N_9745,N_9345);
and U11889 (N_11889,N_8319,N_8833);
nand U11890 (N_11890,N_8198,N_8456);
and U11891 (N_11891,N_9467,N_9210);
or U11892 (N_11892,N_8935,N_9998);
nand U11893 (N_11893,N_8083,N_8598);
nor U11894 (N_11894,N_8594,N_9122);
and U11895 (N_11895,N_8327,N_9891);
xnor U11896 (N_11896,N_8298,N_8974);
and U11897 (N_11897,N_8990,N_8533);
xnor U11898 (N_11898,N_8836,N_9191);
nor U11899 (N_11899,N_9440,N_8422);
xnor U11900 (N_11900,N_9224,N_8383);
and U11901 (N_11901,N_9221,N_9599);
nand U11902 (N_11902,N_9614,N_8736);
or U11903 (N_11903,N_8474,N_9892);
nand U11904 (N_11904,N_9620,N_9078);
and U11905 (N_11905,N_9964,N_8551);
nor U11906 (N_11906,N_9930,N_9643);
nor U11907 (N_11907,N_9413,N_8963);
nor U11908 (N_11908,N_9763,N_9071);
nor U11909 (N_11909,N_8432,N_8214);
or U11910 (N_11910,N_9742,N_9259);
and U11911 (N_11911,N_8771,N_8122);
and U11912 (N_11912,N_9947,N_9257);
or U11913 (N_11913,N_8187,N_9889);
and U11914 (N_11914,N_9730,N_9719);
nand U11915 (N_11915,N_8237,N_8583);
and U11916 (N_11916,N_8195,N_9709);
xor U11917 (N_11917,N_8858,N_9789);
xor U11918 (N_11918,N_9085,N_8440);
xnor U11919 (N_11919,N_8390,N_9081);
nand U11920 (N_11920,N_9151,N_8255);
or U11921 (N_11921,N_9596,N_9971);
nand U11922 (N_11922,N_9603,N_8303);
and U11923 (N_11923,N_9777,N_9056);
and U11924 (N_11924,N_8148,N_9868);
xnor U11925 (N_11925,N_8308,N_9168);
nand U11926 (N_11926,N_9183,N_9736);
nand U11927 (N_11927,N_9065,N_8211);
and U11928 (N_11928,N_9349,N_9402);
nand U11929 (N_11929,N_9408,N_9735);
nor U11930 (N_11930,N_9151,N_8798);
nand U11931 (N_11931,N_8425,N_9893);
nand U11932 (N_11932,N_9899,N_8991);
nand U11933 (N_11933,N_9020,N_9603);
or U11934 (N_11934,N_9923,N_9264);
or U11935 (N_11935,N_9019,N_9375);
xor U11936 (N_11936,N_9270,N_8088);
nor U11937 (N_11937,N_8437,N_9596);
nand U11938 (N_11938,N_8262,N_8801);
and U11939 (N_11939,N_8043,N_8909);
xnor U11940 (N_11940,N_8619,N_8485);
nand U11941 (N_11941,N_8413,N_8219);
nor U11942 (N_11942,N_9243,N_8675);
nor U11943 (N_11943,N_9151,N_9627);
nor U11944 (N_11944,N_9552,N_8241);
and U11945 (N_11945,N_9969,N_8936);
xor U11946 (N_11946,N_8699,N_9547);
nand U11947 (N_11947,N_8790,N_8914);
nor U11948 (N_11948,N_8970,N_8064);
nand U11949 (N_11949,N_8585,N_9458);
nand U11950 (N_11950,N_8178,N_9497);
nand U11951 (N_11951,N_9430,N_8280);
nand U11952 (N_11952,N_9437,N_8321);
nor U11953 (N_11953,N_9286,N_9771);
and U11954 (N_11954,N_9473,N_8000);
and U11955 (N_11955,N_9517,N_8749);
or U11956 (N_11956,N_9419,N_8387);
nand U11957 (N_11957,N_9464,N_9627);
nand U11958 (N_11958,N_8004,N_8540);
or U11959 (N_11959,N_9105,N_8034);
xnor U11960 (N_11960,N_8105,N_9935);
nor U11961 (N_11961,N_8267,N_9599);
nor U11962 (N_11962,N_9631,N_9880);
or U11963 (N_11963,N_9375,N_9563);
and U11964 (N_11964,N_9663,N_9645);
xor U11965 (N_11965,N_8882,N_8973);
or U11966 (N_11966,N_9029,N_9521);
and U11967 (N_11967,N_9528,N_8111);
or U11968 (N_11968,N_9665,N_8778);
nand U11969 (N_11969,N_8705,N_8102);
xor U11970 (N_11970,N_8284,N_9157);
xnor U11971 (N_11971,N_9196,N_9393);
nor U11972 (N_11972,N_8410,N_9983);
and U11973 (N_11973,N_9534,N_8904);
nor U11974 (N_11974,N_9258,N_8082);
or U11975 (N_11975,N_8170,N_9036);
nor U11976 (N_11976,N_9038,N_8945);
and U11977 (N_11977,N_8924,N_9055);
and U11978 (N_11978,N_9159,N_8296);
or U11979 (N_11979,N_8412,N_8710);
xor U11980 (N_11980,N_8477,N_8262);
or U11981 (N_11981,N_8325,N_8239);
xnor U11982 (N_11982,N_8795,N_8004);
and U11983 (N_11983,N_8984,N_9106);
or U11984 (N_11984,N_8876,N_8472);
and U11985 (N_11985,N_9113,N_9835);
xnor U11986 (N_11986,N_8015,N_8913);
nand U11987 (N_11987,N_8007,N_8447);
nor U11988 (N_11988,N_8945,N_9661);
and U11989 (N_11989,N_9200,N_9426);
nand U11990 (N_11990,N_8898,N_9103);
xor U11991 (N_11991,N_9614,N_8404);
and U11992 (N_11992,N_9638,N_8423);
and U11993 (N_11993,N_9634,N_8426);
or U11994 (N_11994,N_8920,N_9281);
and U11995 (N_11995,N_8678,N_9773);
xor U11996 (N_11996,N_9566,N_8050);
nor U11997 (N_11997,N_8081,N_8813);
nand U11998 (N_11998,N_9371,N_8242);
or U11999 (N_11999,N_9640,N_9179);
xnor U12000 (N_12000,N_10297,N_10129);
nor U12001 (N_12001,N_10197,N_10811);
nor U12002 (N_12002,N_11592,N_11244);
nand U12003 (N_12003,N_11327,N_11863);
and U12004 (N_12004,N_11835,N_10694);
xor U12005 (N_12005,N_11583,N_10348);
nor U12006 (N_12006,N_11738,N_11257);
xnor U12007 (N_12007,N_10661,N_11542);
xnor U12008 (N_12008,N_11306,N_10123);
nor U12009 (N_12009,N_11288,N_11567);
or U12010 (N_12010,N_10116,N_11816);
and U12011 (N_12011,N_10070,N_10687);
nand U12012 (N_12012,N_11154,N_11869);
xor U12013 (N_12013,N_11871,N_11423);
and U12014 (N_12014,N_11468,N_10863);
and U12015 (N_12015,N_10463,N_10994);
nor U12016 (N_12016,N_10496,N_11409);
xnor U12017 (N_12017,N_10349,N_10991);
nor U12018 (N_12018,N_10585,N_11575);
nor U12019 (N_12019,N_11482,N_10645);
xnor U12020 (N_12020,N_11351,N_11969);
and U12021 (N_12021,N_11611,N_10933);
or U12022 (N_12022,N_11456,N_10640);
or U12023 (N_12023,N_10621,N_10708);
and U12024 (N_12024,N_11204,N_10968);
nor U12025 (N_12025,N_11493,N_10534);
nand U12026 (N_12026,N_10013,N_10178);
or U12027 (N_12027,N_10165,N_10320);
or U12028 (N_12028,N_11067,N_11130);
or U12029 (N_12029,N_10336,N_11431);
nor U12030 (N_12030,N_11903,N_11939);
xor U12031 (N_12031,N_10308,N_10728);
and U12032 (N_12032,N_11776,N_10975);
or U12033 (N_12033,N_11931,N_10170);
xor U12034 (N_12034,N_11698,N_10449);
nor U12035 (N_12035,N_11398,N_10145);
xnor U12036 (N_12036,N_10515,N_10839);
xor U12037 (N_12037,N_11201,N_10138);
and U12038 (N_12038,N_10808,N_10806);
or U12039 (N_12039,N_11087,N_11368);
nand U12040 (N_12040,N_11483,N_10216);
and U12041 (N_12041,N_10048,N_11068);
xor U12042 (N_12042,N_11720,N_10797);
nand U12043 (N_12043,N_11677,N_10142);
nor U12044 (N_12044,N_10199,N_10194);
nor U12045 (N_12045,N_11660,N_11047);
nor U12046 (N_12046,N_11000,N_11739);
xnor U12047 (N_12047,N_10281,N_10539);
nor U12048 (N_12048,N_11301,N_10397);
and U12049 (N_12049,N_10732,N_10247);
xnor U12050 (N_12050,N_10664,N_10931);
xor U12051 (N_12051,N_10094,N_11976);
nor U12052 (N_12052,N_11399,N_10924);
or U12053 (N_12053,N_10869,N_11641);
or U12054 (N_12054,N_11491,N_10286);
nor U12055 (N_12055,N_11282,N_10840);
xor U12056 (N_12056,N_10493,N_11184);
nor U12057 (N_12057,N_10024,N_11454);
nand U12058 (N_12058,N_11403,N_10686);
nor U12059 (N_12059,N_11653,N_10327);
or U12060 (N_12060,N_11235,N_11886);
nand U12061 (N_12061,N_11316,N_11138);
nand U12062 (N_12062,N_10544,N_10101);
nand U12063 (N_12063,N_11508,N_10910);
nor U12064 (N_12064,N_10016,N_11794);
nand U12065 (N_12065,N_10230,N_10789);
xnor U12066 (N_12066,N_10002,N_10542);
nand U12067 (N_12067,N_11561,N_10020);
and U12068 (N_12068,N_11158,N_10115);
xor U12069 (N_12069,N_10607,N_11674);
nor U12070 (N_12070,N_11919,N_10632);
or U12071 (N_12071,N_11766,N_10273);
or U12072 (N_12072,N_11751,N_11092);
and U12073 (N_12073,N_11627,N_10543);
nand U12074 (N_12074,N_11029,N_10844);
nand U12075 (N_12075,N_11271,N_10492);
and U12076 (N_12076,N_11962,N_11484);
or U12077 (N_12077,N_11986,N_11361);
and U12078 (N_12078,N_11094,N_11145);
nand U12079 (N_12079,N_11810,N_11421);
xor U12080 (N_12080,N_10989,N_10724);
xor U12081 (N_12081,N_11336,N_11198);
nor U12082 (N_12082,N_11551,N_11830);
and U12083 (N_12083,N_11540,N_11314);
or U12084 (N_12084,N_10679,N_11658);
nor U12085 (N_12085,N_10856,N_11119);
nor U12086 (N_12086,N_11297,N_10395);
and U12087 (N_12087,N_11851,N_10814);
or U12088 (N_12088,N_11408,N_11412);
and U12089 (N_12089,N_11817,N_11234);
nand U12090 (N_12090,N_11868,N_11501);
nand U12091 (N_12091,N_10313,N_11917);
xnor U12092 (N_12092,N_10122,N_11189);
nor U12093 (N_12093,N_11418,N_10915);
or U12094 (N_12094,N_11113,N_11550);
xor U12095 (N_12095,N_10654,N_11425);
or U12096 (N_12096,N_11394,N_11120);
xnor U12097 (N_12097,N_11742,N_10793);
or U12098 (N_12098,N_10435,N_10173);
nor U12099 (N_12099,N_10124,N_11325);
and U12100 (N_12100,N_11709,N_10353);
nand U12101 (N_12101,N_10689,N_10064);
nor U12102 (N_12102,N_10053,N_11734);
xor U12103 (N_12103,N_11950,N_10849);
or U12104 (N_12104,N_10825,N_10331);
and U12105 (N_12105,N_11849,N_10155);
nand U12106 (N_12106,N_10545,N_11016);
nand U12107 (N_12107,N_10663,N_10943);
nor U12108 (N_12108,N_10438,N_10057);
xnor U12109 (N_12109,N_10881,N_11285);
nand U12110 (N_12110,N_10316,N_10083);
nor U12111 (N_12111,N_10383,N_10695);
nand U12112 (N_12112,N_11884,N_10425);
nor U12113 (N_12113,N_10309,N_11481);
nor U12114 (N_12114,N_11988,N_10282);
nor U12115 (N_12115,N_10995,N_11356);
nand U12116 (N_12116,N_11892,N_10426);
nor U12117 (N_12117,N_10219,N_11888);
xnor U12118 (N_12118,N_11636,N_10710);
nand U12119 (N_12119,N_11073,N_11977);
xnor U12120 (N_12120,N_11384,N_10890);
nand U12121 (N_12121,N_11944,N_10163);
xnor U12122 (N_12122,N_10831,N_11031);
nand U12123 (N_12123,N_10117,N_10809);
or U12124 (N_12124,N_10030,N_10522);
nor U12125 (N_12125,N_11125,N_10445);
nor U12126 (N_12126,N_10940,N_11993);
nor U12127 (N_12127,N_11935,N_10011);
nand U12128 (N_12128,N_10558,N_10867);
xor U12129 (N_12129,N_10152,N_10644);
or U12130 (N_12130,N_11217,N_11467);
and U12131 (N_12131,N_10935,N_10277);
or U12132 (N_12132,N_10690,N_10485);
or U12133 (N_12133,N_10780,N_11556);
or U12134 (N_12134,N_11172,N_11793);
nor U12135 (N_12135,N_11140,N_11060);
nor U12136 (N_12136,N_11365,N_11442);
or U12137 (N_12137,N_10568,N_11401);
or U12138 (N_12138,N_11630,N_11552);
nand U12139 (N_12139,N_11599,N_10625);
xnor U12140 (N_12140,N_10414,N_11787);
or U12141 (N_12141,N_10424,N_10382);
nand U12142 (N_12142,N_11227,N_10528);
nor U12143 (N_12143,N_11497,N_11203);
nor U12144 (N_12144,N_11461,N_11153);
or U12145 (N_12145,N_10720,N_11434);
or U12146 (N_12146,N_10437,N_10206);
and U12147 (N_12147,N_10893,N_10469);
xor U12148 (N_12148,N_10174,N_10734);
nand U12149 (N_12149,N_10619,N_10352);
nand U12150 (N_12150,N_11837,N_10176);
nand U12151 (N_12151,N_11949,N_11155);
nor U12152 (N_12152,N_11238,N_11232);
and U12153 (N_12153,N_11182,N_10718);
nor U12154 (N_12154,N_11961,N_10570);
xnor U12155 (N_12155,N_11918,N_11545);
and U12156 (N_12156,N_11608,N_11323);
or U12157 (N_12157,N_10314,N_10949);
and U12158 (N_12158,N_10028,N_11001);
xor U12159 (N_12159,N_11331,N_11359);
nor U12160 (N_12160,N_10051,N_10032);
nor U12161 (N_12161,N_10879,N_11514);
or U12162 (N_12162,N_10676,N_11870);
nor U12163 (N_12163,N_11874,N_10618);
xor U12164 (N_12164,N_10378,N_11017);
or U12165 (N_12165,N_11433,N_10604);
nor U12166 (N_12166,N_11825,N_10345);
nor U12167 (N_12167,N_11737,N_10614);
nand U12168 (N_12168,N_11322,N_11829);
and U12169 (N_12169,N_10201,N_11444);
nor U12170 (N_12170,N_11333,N_10322);
nor U12171 (N_12171,N_10250,N_10396);
nand U12172 (N_12172,N_10193,N_11929);
and U12173 (N_12173,N_10525,N_10491);
nand U12174 (N_12174,N_10261,N_10310);
nand U12175 (N_12175,N_10393,N_10775);
xor U12176 (N_12176,N_10498,N_11528);
xnor U12177 (N_12177,N_11590,N_10805);
nand U12178 (N_12178,N_11752,N_10911);
or U12179 (N_12179,N_11048,N_10186);
nor U12180 (N_12180,N_11725,N_11971);
nand U12181 (N_12181,N_10954,N_11866);
or U12182 (N_12182,N_11251,N_10785);
nor U12183 (N_12183,N_11748,N_11254);
and U12184 (N_12184,N_10118,N_11273);
and U12185 (N_12185,N_11202,N_10610);
nor U12186 (N_12186,N_10191,N_10370);
and U12187 (N_12187,N_11972,N_10705);
or U12188 (N_12188,N_10932,N_11978);
xnor U12189 (N_12189,N_10787,N_10183);
or U12190 (N_12190,N_11591,N_10360);
and U12191 (N_12191,N_10877,N_10829);
xor U12192 (N_12192,N_11982,N_11136);
or U12193 (N_12193,N_11774,N_11649);
nand U12194 (N_12194,N_11249,N_10305);
nand U12195 (N_12195,N_11526,N_10486);
nor U12196 (N_12196,N_11762,N_10826);
and U12197 (N_12197,N_11956,N_11521);
xnor U12198 (N_12198,N_10088,N_10634);
nor U12199 (N_12199,N_11926,N_10537);
nand U12200 (N_12200,N_10605,N_10448);
and U12201 (N_12201,N_11936,N_11267);
and U12202 (N_12202,N_10533,N_11360);
nor U12203 (N_12203,N_11631,N_11382);
and U12204 (N_12204,N_10341,N_10796);
xor U12205 (N_12205,N_11906,N_11300);
nand U12206 (N_12206,N_11848,N_10977);
and U12207 (N_12207,N_10195,N_10476);
nand U12208 (N_12208,N_10730,N_11453);
nand U12209 (N_12209,N_11287,N_11879);
xnor U12210 (N_12210,N_10726,N_11838);
nor U12211 (N_12211,N_10630,N_11696);
and U12212 (N_12212,N_10133,N_10015);
xor U12213 (N_12213,N_10008,N_10800);
or U12214 (N_12214,N_11381,N_10266);
nand U12215 (N_12215,N_11240,N_10081);
and U12216 (N_12216,N_11389,N_10578);
nand U12217 (N_12217,N_10061,N_10085);
or U12218 (N_12218,N_10407,N_11124);
nand U12219 (N_12219,N_11842,N_11350);
nor U12220 (N_12220,N_11312,N_11248);
xnor U12221 (N_12221,N_11999,N_11554);
or U12222 (N_12222,N_10420,N_11543);
xor U12223 (N_12223,N_10421,N_10125);
nand U12224 (N_12224,N_10955,N_10459);
nor U12225 (N_12225,N_10357,N_10577);
or U12226 (N_12226,N_10287,N_11980);
and U12227 (N_12227,N_10590,N_10801);
nor U12228 (N_12228,N_10272,N_10752);
and U12229 (N_12229,N_10523,N_11134);
nor U12230 (N_12230,N_11618,N_10819);
nor U12231 (N_12231,N_10538,N_10703);
xor U12232 (N_12232,N_11471,N_11144);
nor U12233 (N_12233,N_10184,N_11662);
or U12234 (N_12234,N_10518,N_10936);
xnor U12235 (N_12235,N_10299,N_11317);
nand U12236 (N_12236,N_11974,N_11353);
xor U12237 (N_12237,N_10300,N_10602);
nand U12238 (N_12238,N_11901,N_10573);
nand U12239 (N_12239,N_10376,N_11400);
nor U12240 (N_12240,N_11688,N_10059);
and U12241 (N_12241,N_10156,N_10942);
nand U12242 (N_12242,N_10624,N_10891);
nand U12243 (N_12243,N_11754,N_10700);
xor U12244 (N_12244,N_10228,N_10744);
and U12245 (N_12245,N_10406,N_11815);
nand U12246 (N_12246,N_10136,N_10919);
nand U12247 (N_12247,N_10803,N_10761);
xor U12248 (N_12248,N_11429,N_11318);
nor U12249 (N_12249,N_11535,N_10892);
nor U12250 (N_12250,N_11195,N_11715);
and U12251 (N_12251,N_11231,N_10569);
and U12252 (N_12252,N_11236,N_11560);
nor U12253 (N_12253,N_10749,N_10777);
xnor U12254 (N_12254,N_11369,N_11455);
and U12255 (N_12255,N_11650,N_10220);
and U12256 (N_12256,N_10470,N_11387);
and U12257 (N_12257,N_11527,N_11756);
nor U12258 (N_12258,N_10641,N_11812);
and U12259 (N_12259,N_11302,N_10662);
or U12260 (N_12260,N_11348,N_11020);
xnor U12261 (N_12261,N_10431,N_11504);
nand U12262 (N_12262,N_11018,N_10853);
or U12263 (N_12263,N_10337,N_11450);
nand U12264 (N_12264,N_10714,N_10212);
and U12265 (N_12265,N_11494,N_11176);
xor U12266 (N_12266,N_11188,N_10458);
nor U12267 (N_12267,N_11907,N_11206);
nand U12268 (N_12268,N_11954,N_10271);
and U12269 (N_12269,N_10131,N_10189);
nor U12270 (N_12270,N_10409,N_11654);
and U12271 (N_12271,N_11833,N_10897);
and U12272 (N_12272,N_10601,N_11072);
xnor U12273 (N_12273,N_11857,N_11127);
nand U12274 (N_12274,N_11637,N_11354);
xor U12275 (N_12275,N_10984,N_11162);
nor U12276 (N_12276,N_10465,N_11487);
xor U12277 (N_12277,N_11479,N_10790);
nand U12278 (N_12278,N_10638,N_10180);
and U12279 (N_12279,N_11564,N_11395);
or U12280 (N_12280,N_11711,N_11924);
xor U12281 (N_12281,N_10121,N_10633);
xor U12282 (N_12282,N_11308,N_11058);
nor U12283 (N_12283,N_11622,N_11506);
or U12284 (N_12284,N_10862,N_11809);
nor U12285 (N_12285,N_11372,N_11490);
xor U12286 (N_12286,N_10683,N_10966);
or U12287 (N_12287,N_10557,N_10597);
or U12288 (N_12288,N_11876,N_10227);
or U12289 (N_12289,N_11781,N_10304);
nand U12290 (N_12290,N_10511,N_10482);
xor U12291 (N_12291,N_10340,N_11729);
and U12292 (N_12292,N_11464,N_10017);
nand U12293 (N_12293,N_11533,N_10914);
nand U12294 (N_12294,N_11411,N_11451);
and U12295 (N_12295,N_10697,N_11726);
nor U12296 (N_12296,N_10467,N_10794);
or U12297 (N_12297,N_10411,N_10643);
nor U12298 (N_12298,N_11164,N_11856);
and U12299 (N_12299,N_11413,N_10530);
nand U12300 (N_12300,N_10161,N_10418);
and U12301 (N_12301,N_11963,N_10905);
nor U12302 (N_12302,N_11790,N_10574);
nand U12303 (N_12303,N_10205,N_10218);
nand U12304 (N_12304,N_11003,N_10450);
nor U12305 (N_12305,N_10549,N_10288);
xor U12306 (N_12306,N_11960,N_10364);
and U12307 (N_12307,N_11771,N_11416);
xor U12308 (N_12308,N_11078,N_10715);
nor U12309 (N_12309,N_10179,N_10665);
nand U12310 (N_12310,N_11463,N_11516);
xnor U12311 (N_12311,N_10381,N_10973);
nand U12312 (N_12312,N_11272,N_10615);
nand U12313 (N_12313,N_10307,N_10894);
xnor U12314 (N_12314,N_11968,N_11958);
or U12315 (N_12315,N_11743,N_10938);
nor U12316 (N_12316,N_10102,N_11230);
nor U12317 (N_12317,N_11131,N_11759);
or U12318 (N_12318,N_11205,N_10846);
nand U12319 (N_12319,N_11761,N_11459);
and U12320 (N_12320,N_11358,N_10251);
and U12321 (N_12321,N_10171,N_11967);
and U12322 (N_12322,N_11652,N_10965);
and U12323 (N_12323,N_11745,N_10739);
nor U12324 (N_12324,N_10899,N_11981);
xnor U12325 (N_12325,N_10267,N_11557);
nand U12326 (N_12326,N_10592,N_11510);
xor U12327 (N_12327,N_11022,N_10875);
xor U12328 (N_12328,N_10012,N_10754);
xor U12329 (N_12329,N_10816,N_10154);
and U12330 (N_12330,N_10146,N_10392);
or U12331 (N_12331,N_11605,N_11079);
and U12332 (N_12332,N_10471,N_11841);
nand U12333 (N_12333,N_10084,N_11375);
or U12334 (N_12334,N_10810,N_10818);
and U12335 (N_12335,N_11291,N_11645);
xnor U12336 (N_12336,N_11639,N_11495);
and U12337 (N_12337,N_11702,N_10361);
xnor U12338 (N_12338,N_10512,N_11789);
or U12339 (N_12339,N_10692,N_11229);
nor U12340 (N_12340,N_10139,N_10007);
xnor U12341 (N_12341,N_11405,N_10872);
nor U12342 (N_12342,N_10150,N_10572);
and U12343 (N_12343,N_10652,N_11749);
nand U12344 (N_12344,N_10385,N_10743);
xnor U12345 (N_12345,N_11763,N_11985);
nand U12346 (N_12346,N_11224,N_10058);
and U12347 (N_12347,N_11635,N_11335);
nor U12348 (N_12348,N_11824,N_11397);
nand U12349 (N_12349,N_11277,N_10760);
nand U12350 (N_12350,N_11573,N_11965);
or U12351 (N_12351,N_10095,N_11678);
and U12352 (N_12352,N_11443,N_10507);
and U12353 (N_12353,N_11607,N_10656);
nor U12354 (N_12354,N_11097,N_11035);
nor U12355 (N_12355,N_10490,N_10258);
nand U12356 (N_12356,N_10778,N_11713);
nand U12357 (N_12357,N_11476,N_10434);
nand U12358 (N_12358,N_10895,N_10182);
nand U12359 (N_12359,N_11160,N_10584);
nor U12360 (N_12360,N_11885,N_11860);
xnor U12361 (N_12361,N_10209,N_10443);
xnor U12362 (N_12362,N_11983,N_11899);
xor U12363 (N_12363,N_10772,N_10576);
xor U12364 (N_12364,N_10120,N_10859);
xor U12365 (N_12365,N_10706,N_11165);
nand U12366 (N_12366,N_10992,N_11428);
and U12367 (N_12367,N_10041,N_11009);
nor U12368 (N_12368,N_11013,N_10413);
or U12369 (N_12369,N_11038,N_11213);
and U12370 (N_12370,N_11284,N_11724);
or U12371 (N_12371,N_11534,N_11243);
nand U12372 (N_12372,N_10091,N_11150);
xor U12373 (N_12373,N_10480,N_11264);
nor U12374 (N_12374,N_10845,N_11680);
and U12375 (N_12375,N_10318,N_11448);
nor U12376 (N_12376,N_11700,N_11077);
and U12377 (N_12377,N_11502,N_10046);
or U12378 (N_12378,N_10215,N_11915);
nor U12379 (N_12379,N_10946,N_10976);
xnor U12380 (N_12380,N_10750,N_10517);
or U12381 (N_12381,N_10903,N_11818);
nand U12382 (N_12382,N_11286,N_10781);
nor U12383 (N_12383,N_10211,N_11030);
nand U12384 (N_12384,N_10255,N_10035);
xnor U12385 (N_12385,N_10527,N_11994);
and U12386 (N_12386,N_11190,N_11209);
nor U12387 (N_12387,N_11952,N_10256);
xnor U12388 (N_12388,N_11595,N_10196);
or U12389 (N_12389,N_11299,N_10702);
or U12390 (N_12390,N_11666,N_10958);
xor U12391 (N_12391,N_11033,N_10359);
nand U12392 (N_12392,N_11692,N_10725);
or U12393 (N_12393,N_11719,N_10505);
nand U12394 (N_12394,N_11933,N_10389);
nor U12395 (N_12395,N_11991,N_11755);
nor U12396 (N_12396,N_10036,N_10850);
or U12397 (N_12397,N_11619,N_10329);
and U12398 (N_12398,N_11806,N_10044);
or U12399 (N_12399,N_10843,N_11191);
and U12400 (N_12400,N_11007,N_11861);
or U12401 (N_12401,N_11383,N_10295);
nor U12402 (N_12402,N_10873,N_11912);
or U12403 (N_12403,N_10321,N_10052);
xnor U12404 (N_12404,N_10637,N_11701);
xnor U12405 (N_12405,N_10766,N_11095);
nor U12406 (N_12406,N_11538,N_11081);
nand U12407 (N_12407,N_10080,N_11161);
or U12408 (N_12408,N_10157,N_11945);
or U12409 (N_12409,N_11558,N_10334);
xnor U12410 (N_12410,N_10144,N_10647);
xor U12411 (N_12411,N_10575,N_10929);
nand U12412 (N_12412,N_10999,N_10099);
nand U12413 (N_12413,N_11430,N_11539);
and U12414 (N_12414,N_10468,N_10009);
or U12415 (N_12415,N_10148,N_10830);
nand U12416 (N_12416,N_11122,N_11565);
nor U12417 (N_12417,N_11684,N_10489);
or U12418 (N_12418,N_11681,N_11946);
nand U12419 (N_12419,N_11782,N_10200);
or U12420 (N_12420,N_11295,N_10065);
nand U12421 (N_12421,N_10520,N_11061);
xnor U12422 (N_12422,N_11574,N_10678);
or U12423 (N_12423,N_11458,N_11208);
xnor U12424 (N_12424,N_10552,N_11625);
and U12425 (N_12425,N_10472,N_11750);
and U12426 (N_12426,N_10242,N_11883);
xor U12427 (N_12427,N_11324,N_10848);
or U12428 (N_12428,N_10087,N_10909);
and U12429 (N_12429,N_11406,N_10698);
and U12430 (N_12430,N_10140,N_11044);
nor U12431 (N_12431,N_10763,N_11727);
xor U12432 (N_12432,N_11050,N_11435);
and U12433 (N_12433,N_10865,N_10113);
xor U12434 (N_12434,N_11896,N_10603);
or U12435 (N_12435,N_10067,N_11315);
xor U12436 (N_12436,N_10040,N_11041);
or U12437 (N_12437,N_10651,N_10926);
or U12438 (N_12438,N_10741,N_10107);
nor U12439 (N_12439,N_11632,N_11832);
and U12440 (N_12440,N_10753,N_11518);
and U12441 (N_12441,N_11052,N_10723);
xnor U12442 (N_12442,N_11364,N_10745);
and U12443 (N_12443,N_11672,N_11005);
nand U12444 (N_12444,N_11588,N_11987);
xor U12445 (N_12445,N_11875,N_11194);
or U12446 (N_12446,N_11347,N_10996);
nor U12447 (N_12447,N_11548,N_11858);
and U12448 (N_12448,N_10442,N_10177);
and U12449 (N_12449,N_10068,N_10038);
nand U12450 (N_12450,N_10917,N_11332);
and U12451 (N_12451,N_11133,N_10868);
xnor U12452 (N_12452,N_10137,N_10422);
xnor U12453 (N_12453,N_11800,N_10278);
nand U12454 (N_12454,N_11321,N_11791);
nand U12455 (N_12455,N_10834,N_11811);
and U12456 (N_12456,N_11717,N_11010);
and U12457 (N_12457,N_10981,N_11582);
xor U12458 (N_12458,N_11853,N_11862);
or U12459 (N_12459,N_11388,N_11784);
and U12460 (N_12460,N_10681,N_11640);
nand U12461 (N_12461,N_11283,N_11820);
nand U12462 (N_12462,N_10003,N_11174);
and U12463 (N_12463,N_10713,N_10263);
nor U12464 (N_12464,N_10755,N_10606);
nor U12465 (N_12465,N_10284,N_11266);
nand U12466 (N_12466,N_11269,N_11687);
xor U12467 (N_12467,N_10925,N_10055);
xnor U12468 (N_12468,N_11628,N_10112);
nand U12469 (N_12469,N_10870,N_10060);
nand U12470 (N_12470,N_10639,N_11722);
nor U12471 (N_12471,N_11085,N_11123);
nor U12472 (N_12472,N_10784,N_11589);
and U12473 (N_12473,N_10985,N_11686);
nor U12474 (N_12474,N_10000,N_11247);
nor U12475 (N_12475,N_11909,N_10786);
xor U12476 (N_12476,N_10792,N_11753);
nand U12477 (N_12477,N_11877,N_10956);
xnor U12478 (N_12478,N_11452,N_10682);
xor U12479 (N_12479,N_11307,N_10338);
or U12480 (N_12480,N_10172,N_10961);
nand U12481 (N_12481,N_10026,N_10312);
nor U12482 (N_12482,N_10583,N_11777);
nor U12483 (N_12483,N_10223,N_10855);
nand U12484 (N_12484,N_11096,N_11051);
or U12485 (N_12485,N_11002,N_10900);
nor U12486 (N_12486,N_10440,N_10626);
and U12487 (N_12487,N_11345,N_11855);
nand U12488 (N_12488,N_10769,N_10904);
and U12489 (N_12489,N_11643,N_11404);
and U12490 (N_12490,N_11177,N_11225);
xnor U12491 (N_12491,N_10423,N_10335);
xnor U12492 (N_12492,N_10368,N_10073);
or U12493 (N_12493,N_11889,N_10560);
or U12494 (N_12494,N_10444,N_10119);
and U12495 (N_12495,N_11326,N_10462);
nor U12496 (N_12496,N_10246,N_10798);
nor U12497 (N_12497,N_11596,N_11319);
nand U12498 (N_12498,N_10709,N_11407);
and U12499 (N_12499,N_11775,N_11865);
xor U12500 (N_12500,N_10387,N_10841);
or U12501 (N_12501,N_11904,N_11769);
xnor U12502 (N_12502,N_11708,N_10232);
nand U12503 (N_12503,N_10021,N_11902);
and U12504 (N_12504,N_11187,N_10497);
or U12505 (N_12505,N_10913,N_10236);
or U12506 (N_12506,N_11910,N_10369);
nor U12507 (N_12507,N_10071,N_11274);
xor U12508 (N_12508,N_10934,N_10210);
nor U12509 (N_12509,N_11004,N_11091);
nand U12510 (N_12510,N_10132,N_11069);
nand U12511 (N_12511,N_10226,N_11669);
and U12512 (N_12512,N_11059,N_11612);
or U12513 (N_12513,N_10078,N_10567);
or U12514 (N_12514,N_11419,N_10054);
or U12515 (N_12515,N_10100,N_11587);
and U12516 (N_12516,N_11895,N_10436);
and U12517 (N_12517,N_11925,N_11152);
xor U12518 (N_12518,N_10483,N_11996);
nor U12519 (N_12519,N_11292,N_11928);
xnor U12520 (N_12520,N_11167,N_10719);
and U12521 (N_12521,N_10631,N_11488);
nand U12522 (N_12522,N_11329,N_11617);
or U12523 (N_12523,N_10898,N_11379);
nand U12524 (N_12524,N_10532,N_10531);
nor U12525 (N_12525,N_11168,N_10430);
xnor U12526 (N_12526,N_10441,N_11241);
or U12527 (N_12527,N_11932,N_10185);
or U12528 (N_12528,N_11898,N_10487);
nor U12529 (N_12529,N_11100,N_10283);
nor U12530 (N_12530,N_10742,N_10330);
and U12531 (N_12531,N_11569,N_11173);
xor U12532 (N_12532,N_10758,N_10599);
xor U12533 (N_12533,N_10390,N_11673);
or U12534 (N_12534,N_11088,N_10043);
xor U12535 (N_12535,N_10550,N_11716);
and U12536 (N_12536,N_11549,N_11114);
xnor U12537 (N_12537,N_11328,N_11485);
nor U12538 (N_12538,N_10428,N_11601);
nor U12539 (N_12539,N_11655,N_10162);
xor U12540 (N_12540,N_10159,N_11070);
nor U12541 (N_12541,N_11378,N_10817);
and U12542 (N_12542,N_10764,N_11822);
xnor U12543 (N_12543,N_11998,N_11391);
nor U12544 (N_12544,N_11341,N_10229);
and U12545 (N_12545,N_10835,N_11511);
xnor U12546 (N_12546,N_11562,N_10241);
and U12547 (N_12547,N_10883,N_10669);
or U12548 (N_12548,N_10788,N_10104);
nor U12549 (N_12549,N_10866,N_11112);
or U12550 (N_12550,N_10579,N_10668);
nor U12551 (N_12551,N_10405,N_10871);
nor U12552 (N_12552,N_10291,N_11836);
and U12553 (N_12553,N_10264,N_11199);
nand U12554 (N_12554,N_11572,N_11330);
and U12555 (N_12555,N_11371,N_11663);
or U12556 (N_12556,N_10791,N_10453);
and U12557 (N_12557,N_10022,N_10105);
xnor U12558 (N_12558,N_11420,N_10696);
nor U12559 (N_12559,N_11480,N_10783);
and U12560 (N_12560,N_11275,N_11175);
nor U12561 (N_12561,N_11289,N_10111);
nand U12562 (N_12562,N_11278,N_10004);
or U12563 (N_12563,N_11449,N_10260);
nand U12564 (N_12564,N_11024,N_10774);
xnor U12565 (N_12565,N_10716,N_11422);
nor U12566 (N_12566,N_10066,N_11108);
xor U12567 (N_12567,N_11474,N_10037);
nor U12568 (N_12568,N_11656,N_10356);
nand U12569 (N_12569,N_11731,N_11957);
nor U12570 (N_12570,N_11415,N_10233);
nand U12571 (N_12571,N_11566,N_11616);
nand U12572 (N_12572,N_11803,N_11911);
nand U12573 (N_12573,N_10311,N_11357);
xnor U12574 (N_12574,N_10562,N_10417);
xnor U12575 (N_12575,N_11268,N_11814);
nor U12576 (N_12576,N_11697,N_10988);
nand U12577 (N_12577,N_10275,N_11647);
nor U12578 (N_12578,N_10541,N_10751);
nor U12579 (N_12579,N_10874,N_11143);
nand U12580 (N_12580,N_10930,N_11417);
nor U12581 (N_12581,N_11186,N_10265);
nand U12582 (N_12582,N_11057,N_10446);
or U12583 (N_12583,N_10388,N_11008);
nand U12584 (N_12584,N_11989,N_11252);
nand U12585 (N_12585,N_10143,N_10722);
nor U12586 (N_12586,N_11163,N_10198);
and U12587 (N_12587,N_11804,N_10049);
nor U12588 (N_12588,N_11294,N_10027);
or U12589 (N_12589,N_11137,N_10433);
and U12590 (N_12590,N_11828,N_10659);
nand U12591 (N_12591,N_10135,N_11496);
nor U12592 (N_12592,N_10882,N_11126);
nor U12593 (N_12593,N_10069,N_10386);
xor U12594 (N_12594,N_11920,N_11393);
xnor U12595 (N_12595,N_10031,N_11513);
or U12596 (N_12596,N_11212,N_10106);
nand U12597 (N_12597,N_11642,N_11042);
nor U12598 (N_12598,N_10896,N_10595);
xnor U12599 (N_12599,N_10168,N_11802);
nand U12600 (N_12600,N_11099,N_11930);
xnor U12601 (N_12601,N_10025,N_10323);
and U12602 (N_12602,N_11975,N_11772);
and U12603 (N_12603,N_11465,N_10548);
nor U12604 (N_12604,N_10253,N_11532);
xnor U12605 (N_12605,N_11064,N_11216);
and U12606 (N_12606,N_10776,N_10375);
nand U12607 (N_12607,N_11259,N_11390);
nand U12608 (N_12608,N_11142,N_11492);
and U12609 (N_12609,N_11169,N_10589);
nor U12610 (N_12610,N_11805,N_11279);
and U12611 (N_12611,N_10367,N_11436);
nor U12612 (N_12612,N_11166,N_11524);
xnor U12613 (N_12613,N_11466,N_10842);
nor U12614 (N_12614,N_11066,N_10677);
xnor U12615 (N_12615,N_10547,N_10508);
nand U12616 (N_12616,N_11437,N_10296);
nor U12617 (N_12617,N_10673,N_11603);
and U12618 (N_12618,N_10324,N_11115);
nand U12619 (N_12619,N_10333,N_10366);
and U12620 (N_12620,N_10707,N_10464);
nor U12621 (N_12621,N_10408,N_11116);
xor U12622 (N_12622,N_10902,N_11585);
nand U12623 (N_12623,N_10456,N_11427);
xnor U12624 (N_12624,N_10952,N_10907);
nand U12625 (N_12625,N_11355,N_11872);
and U12626 (N_12626,N_11544,N_10555);
or U12627 (N_12627,N_11614,N_11139);
xnor U12628 (N_12628,N_10350,N_11222);
nand U12629 (N_12629,N_10114,N_10948);
xnor U12630 (N_12630,N_11036,N_10006);
and U12631 (N_12631,N_11489,N_11445);
or U12632 (N_12632,N_11012,N_10290);
and U12633 (N_12633,N_11149,N_11973);
xnor U12634 (N_12634,N_11082,N_10941);
nand U12635 (N_12635,N_10243,N_11736);
nor U12636 (N_12636,N_10029,N_10513);
nand U12637 (N_12637,N_11414,N_10622);
and U12638 (N_12638,N_11089,N_11531);
and U12639 (N_12639,N_10586,N_10649);
or U12640 (N_12640,N_11880,N_11179);
nor U12641 (N_12641,N_11555,N_10317);
xor U12642 (N_12642,N_11280,N_10292);
nand U12643 (N_12643,N_10151,N_10158);
and U12644 (N_12644,N_11522,N_10454);
and U12645 (N_12645,N_11764,N_11290);
nor U12646 (N_12646,N_10225,N_11921);
xor U12647 (N_12647,N_11563,N_10221);
nand U12648 (N_12648,N_11185,N_11576);
nor U12649 (N_12649,N_11053,N_11626);
nor U12650 (N_12650,N_11103,N_11104);
nand U12651 (N_12651,N_10711,N_11062);
nand U12652 (N_12652,N_11740,N_11797);
or U12653 (N_12653,N_11032,N_10691);
nor U12654 (N_12654,N_10153,N_10684);
or U12655 (N_12655,N_10737,N_10611);
nor U12656 (N_12656,N_11695,N_11801);
or U12657 (N_12657,N_11597,N_11065);
nand U12658 (N_12658,N_11512,N_11786);
nand U12659 (N_12659,N_10072,N_10108);
or U12660 (N_12660,N_10010,N_11546);
xor U12661 (N_12661,N_11303,N_11530);
and U12662 (N_12662,N_11859,N_11349);
xnor U12663 (N_12663,N_11043,N_11634);
nor U12664 (N_12664,N_11440,N_10276);
or U12665 (N_12665,N_10033,N_11233);
and U12666 (N_12666,N_11362,N_11151);
xnor U12667 (N_12667,N_11304,N_10192);
xnor U12668 (N_12668,N_11439,N_11844);
or U12669 (N_12669,N_11083,N_11712);
nand U12670 (N_12670,N_11373,N_10280);
xnor U12671 (N_12671,N_10160,N_10526);
and U12672 (N_12672,N_11964,N_11938);
nor U12673 (N_12673,N_10937,N_11410);
nor U12674 (N_12674,N_10768,N_10514);
nor U12675 (N_12675,N_10947,N_10415);
nor U12676 (N_12676,N_10499,N_11117);
and U12677 (N_12677,N_11226,N_11651);
nor U12678 (N_12678,N_11659,N_10213);
nand U12679 (N_12679,N_10886,N_10922);
nor U12680 (N_12680,N_10852,N_10346);
and U12681 (N_12681,N_11180,N_10807);
nand U12682 (N_12682,N_10452,N_10014);
and U12683 (N_12683,N_10927,N_11034);
xnor U12684 (N_12684,N_11261,N_11721);
and U12685 (N_12685,N_11086,N_11577);
nand U12686 (N_12686,N_11311,N_10556);
and U12687 (N_12687,N_11025,N_10190);
and U12688 (N_12688,N_10403,N_11046);
nand U12689 (N_12689,N_11109,N_11693);
xor U12690 (N_12690,N_10918,N_10203);
nor U12691 (N_12691,N_10983,N_10097);
nand U12692 (N_12692,N_10920,N_10939);
nand U12693 (N_12693,N_11947,N_11867);
xnor U12694 (N_12694,N_11507,N_11878);
nand U12695 (N_12695,N_10916,N_10636);
nor U12696 (N_12696,N_11320,N_10398);
and U12697 (N_12697,N_10371,N_11951);
nand U12698 (N_12698,N_11881,N_10347);
xnor U12699 (N_12699,N_11598,N_10986);
nand U12700 (N_12700,N_11106,N_10928);
nor U12701 (N_12701,N_10325,N_10249);
or U12702 (N_12702,N_11827,N_11110);
nor U12703 (N_12703,N_11783,N_10399);
nand U12704 (N_12704,N_11352,N_10328);
or U12705 (N_12705,N_10379,N_10524);
xor U12706 (N_12706,N_11900,N_11940);
and U12707 (N_12707,N_11380,N_11568);
and U12708 (N_12708,N_11937,N_11309);
or U12709 (N_12709,N_10001,N_11682);
xor U12710 (N_12710,N_11027,N_11258);
nand U12711 (N_12711,N_11733,N_11758);
and U12712 (N_12712,N_11170,N_10957);
nand U12713 (N_12713,N_11679,N_10169);
and U12714 (N_12714,N_11220,N_11779);
and U12715 (N_12715,N_11157,N_10980);
or U12716 (N_12716,N_10503,N_11665);
and U12717 (N_12717,N_10298,N_10623);
or U12718 (N_12718,N_10731,N_11438);
xnor U12719 (N_12719,N_11840,N_11646);
and U12720 (N_12720,N_10535,N_10901);
nor U12721 (N_12721,N_11891,N_11313);
nand U12722 (N_12722,N_10969,N_10217);
nand U12723 (N_12723,N_10092,N_10738);
nor U12724 (N_12724,N_11683,N_10740);
nor U12725 (N_12725,N_10460,N_10762);
nor U12726 (N_12726,N_10813,N_10735);
or U12727 (N_12727,N_10979,N_11218);
xnor U12728 (N_12728,N_11525,N_10238);
and U12729 (N_12729,N_11246,N_10756);
and U12730 (N_12730,N_10821,N_11193);
nand U12731 (N_12731,N_11023,N_11037);
and U12732 (N_12732,N_11823,N_10953);
or U12733 (N_12733,N_11953,N_11593);
nor U12734 (N_12734,N_11090,N_11704);
and U12735 (N_12735,N_10770,N_10642);
nor U12736 (N_12736,N_10596,N_10090);
nor U12737 (N_12737,N_10248,N_11211);
xor U12738 (N_12738,N_10098,N_10086);
nor U12739 (N_12739,N_11770,N_11080);
nor U12740 (N_12740,N_10571,N_10455);
nand U12741 (N_12741,N_11922,N_11342);
xor U12742 (N_12742,N_10546,N_11256);
xnor U12743 (N_12743,N_10224,N_10259);
and U12744 (N_12744,N_10509,N_10502);
nor U12745 (N_12745,N_11509,N_10134);
nor U12746 (N_12746,N_11821,N_10302);
xor U12747 (N_12747,N_11916,N_11897);
nand U12748 (N_12748,N_10293,N_11948);
xnor U12749 (N_12749,N_10050,N_11765);
and U12750 (N_12750,N_11367,N_10593);
nand U12751 (N_12751,N_11093,N_11098);
nand U12752 (N_12752,N_11621,N_10301);
nor U12753 (N_12753,N_11071,N_10401);
or U12754 (N_12754,N_11344,N_10771);
and U12755 (N_12755,N_11056,N_10987);
xor U12756 (N_12756,N_11699,N_11873);
nor U12757 (N_12757,N_10609,N_10967);
nor U12758 (N_12758,N_10993,N_11028);
or U12759 (N_12759,N_10245,N_11768);
xnor U12760 (N_12760,N_10062,N_10876);
or U12761 (N_12761,N_10594,N_10795);
nor U12762 (N_12762,N_11559,N_11586);
nor U12763 (N_12763,N_10019,N_10110);
nand U12764 (N_12764,N_11475,N_10374);
or U12765 (N_12765,N_10627,N_11536);
xor U12766 (N_12766,N_11970,N_11281);
or U12767 (N_12767,N_11118,N_11214);
xor U12768 (N_12768,N_11276,N_10563);
xor U12769 (N_12769,N_11741,N_11260);
xor U12770 (N_12770,N_11541,N_11718);
xnor U12771 (N_12771,N_10478,N_11245);
nor U12772 (N_12772,N_11006,N_10082);
xnor U12773 (N_12773,N_10721,N_10675);
or U12774 (N_12774,N_10056,N_11197);
nor U12775 (N_12775,N_10519,N_11606);
or U12776 (N_12776,N_10885,N_11959);
nor U12777 (N_12777,N_11021,N_10473);
and U12778 (N_12778,N_10103,N_11594);
xor U12779 (N_12779,N_10457,N_11200);
nand U12780 (N_12780,N_10342,N_10598);
and U12781 (N_12781,N_10704,N_10884);
or U12782 (N_12782,N_11570,N_11305);
xor U12783 (N_12783,N_11602,N_10391);
xor U12784 (N_12784,N_11171,N_11376);
xnor U12785 (N_12785,N_11584,N_11529);
xor U12786 (N_12786,N_11045,N_10832);
or U12787 (N_12787,N_10912,N_11600);
nand U12788 (N_12788,N_11610,N_10944);
nor U12789 (N_12789,N_10650,N_10181);
nor U12790 (N_12790,N_10773,N_11890);
or U12791 (N_12791,N_11746,N_11730);
xor U12792 (N_12792,N_10733,N_11792);
nor U12793 (N_12793,N_10660,N_11210);
nor U12794 (N_12794,N_11128,N_10306);
and U12795 (N_12795,N_10962,N_10998);
or U12796 (N_12796,N_10824,N_10477);
nand U12797 (N_12797,N_11995,N_11923);
and U12798 (N_12798,N_10963,N_10591);
nand U12799 (N_12799,N_10466,N_11706);
xnor U12800 (N_12800,N_11181,N_11691);
xnor U12801 (N_12801,N_10657,N_11159);
xnor U12802 (N_12802,N_11148,N_10906);
nor U12803 (N_12803,N_10214,N_10628);
or U12804 (N_12804,N_10339,N_10419);
nor U12805 (N_12805,N_11049,N_10351);
nand U12806 (N_12806,N_10951,N_10354);
or U12807 (N_12807,N_11338,N_10187);
nand U12808 (N_12808,N_10802,N_11773);
xor U12809 (N_12809,N_10175,N_11934);
or U12810 (N_12810,N_10074,N_11633);
and U12811 (N_12811,N_10667,N_11638);
or U12812 (N_12812,N_11386,N_11242);
and U12813 (N_12813,N_10270,N_11629);
and U12814 (N_12814,N_11263,N_11788);
or U12815 (N_12815,N_10608,N_11547);
xnor U12816 (N_12816,N_10655,N_11334);
and U12817 (N_12817,N_10268,N_11457);
nor U12818 (N_12818,N_11984,N_11845);
nand U12819 (N_12819,N_11441,N_10565);
xor U12820 (N_12820,N_10561,N_10959);
and U12821 (N_12821,N_11723,N_11505);
nand U12822 (N_12822,N_10447,N_10076);
nand U12823 (N_12823,N_11799,N_10377);
xnor U12824 (N_12824,N_11239,N_11310);
nand U12825 (N_12825,N_11571,N_10712);
nor U12826 (N_12826,N_10096,N_10945);
nand U12827 (N_12827,N_11908,N_11396);
xnor U12828 (N_12828,N_11343,N_11694);
nand U12829 (N_12829,N_10727,N_11648);
and U12830 (N_12830,N_10045,N_10729);
or U12831 (N_12831,N_10495,N_10416);
or U12832 (N_12832,N_11997,N_10504);
nand U12833 (N_12833,N_11374,N_10332);
nor U12834 (N_12834,N_10612,N_10285);
nor U12835 (N_12835,N_10373,N_11615);
and U12836 (N_12836,N_10147,N_10484);
xor U12837 (N_12837,N_11675,N_11850);
xnor U12838 (N_12838,N_11146,N_10252);
and U12839 (N_12839,N_11503,N_10587);
nor U12840 (N_12840,N_10553,N_10208);
nand U12841 (N_12841,N_10130,N_11893);
and U12842 (N_12842,N_11298,N_11979);
nand U12843 (N_12843,N_10782,N_10580);
nor U12844 (N_12844,N_11613,N_11486);
or U12845 (N_12845,N_11670,N_10566);
and U12846 (N_12846,N_10997,N_10648);
nand U12847 (N_12847,N_10394,N_10889);
nor U12848 (N_12848,N_10990,N_10362);
xnor U12849 (N_12849,N_11667,N_10439);
and U12850 (N_12850,N_11432,N_11255);
nand U12851 (N_12851,N_10551,N_11894);
xnor U12852 (N_12852,N_11671,N_11074);
nor U12853 (N_12853,N_11664,N_11472);
nor U12854 (N_12854,N_10974,N_11966);
nand U12855 (N_12855,N_11366,N_10620);
nand U12856 (N_12856,N_10757,N_10950);
nor U12857 (N_12857,N_11927,N_10257);
xor U12858 (N_12858,N_10262,N_10854);
and U12859 (N_12859,N_11253,N_11778);
nor U12860 (N_12860,N_10141,N_10613);
and U12861 (N_12861,N_10582,N_11111);
or U12862 (N_12862,N_11377,N_10289);
xnor U12863 (N_12863,N_11499,N_10670);
nand U12864 (N_12864,N_10748,N_10581);
and U12865 (N_12865,N_11839,N_11500);
nand U12866 (N_12866,N_11796,N_10326);
nor U12867 (N_12867,N_11831,N_11446);
nand U12868 (N_12868,N_11846,N_11676);
xor U12869 (N_12869,N_11129,N_11337);
or U12870 (N_12870,N_11462,N_10204);
nand U12871 (N_12871,N_10564,N_10034);
and U12872 (N_12872,N_11864,N_10126);
xor U12873 (N_12873,N_11011,N_10501);
nand U12874 (N_12874,N_11798,N_11780);
and U12875 (N_12875,N_10837,N_10653);
nand U12876 (N_12876,N_10964,N_11402);
nand U12877 (N_12877,N_10923,N_11760);
xnor U12878 (N_12878,N_11147,N_10747);
and U12879 (N_12879,N_10828,N_11478);
xnor U12880 (N_12880,N_10510,N_10838);
nand U12881 (N_12881,N_11015,N_11262);
nand U12882 (N_12882,N_11992,N_10432);
nor U12883 (N_12883,N_11523,N_11955);
nor U12884 (N_12884,N_10671,N_10294);
or U12885 (N_12885,N_11265,N_10759);
nand U12886 (N_12886,N_11470,N_11942);
xor U12887 (N_12887,N_11914,N_10075);
nand U12888 (N_12888,N_11834,N_11537);
and U12889 (N_12889,N_10488,N_10355);
and U12890 (N_12890,N_11105,N_10908);
nand U12891 (N_12891,N_10921,N_11102);
and U12892 (N_12892,N_11517,N_10982);
xor U12893 (N_12893,N_11196,N_10479);
or U12894 (N_12894,N_11943,N_10254);
xor U12895 (N_12895,N_11941,N_11370);
and U12896 (N_12896,N_10972,N_11757);
xnor U12897 (N_12897,N_11101,N_10812);
xor U12898 (N_12898,N_11447,N_10063);
nor U12899 (N_12899,N_11580,N_10617);
xor U12900 (N_12900,N_11620,N_10978);
and U12901 (N_12901,N_11250,N_11339);
xnor U12902 (N_12902,N_11014,N_10864);
or U12903 (N_12903,N_10860,N_10023);
nand U12904 (N_12904,N_11515,N_10164);
or U12905 (N_12905,N_10365,N_11767);
xnor U12906 (N_12906,N_11135,N_11689);
and U12907 (N_12907,N_10481,N_10018);
and U12908 (N_12908,N_10799,N_10400);
xor U12909 (N_12909,N_10412,N_10274);
nand U12910 (N_12910,N_11221,N_11084);
nor U12911 (N_12911,N_11228,N_11623);
or U12912 (N_12912,N_11207,N_10128);
or U12913 (N_12913,N_11477,N_11270);
xor U12914 (N_12914,N_10222,N_10005);
or U12915 (N_12915,N_10540,N_11847);
xnor U12916 (N_12916,N_11661,N_10207);
and U12917 (N_12917,N_10358,N_11690);
xor U12918 (N_12918,N_10858,N_10319);
or U12919 (N_12919,N_11520,N_11710);
nand U12920 (N_12920,N_11604,N_10240);
nor U12921 (N_12921,N_11121,N_11107);
nand U12922 (N_12922,N_11826,N_11747);
xnor U12923 (N_12923,N_10878,N_10736);
or U12924 (N_12924,N_10475,N_10861);
nor U12925 (N_12925,N_10079,N_11019);
or U12926 (N_12926,N_10559,N_10166);
nor U12927 (N_12927,N_11714,N_10688);
or U12928 (N_12928,N_11178,N_11054);
or U12929 (N_12929,N_10685,N_11237);
nand U12930 (N_12930,N_10461,N_11039);
nor U12931 (N_12931,N_10093,N_10516);
or U12932 (N_12932,N_10077,N_11293);
nand U12933 (N_12933,N_11219,N_10380);
xnor U12934 (N_12934,N_11852,N_10888);
or U12935 (N_12935,N_10042,N_11887);
nand U12936 (N_12936,N_10244,N_11609);
or U12937 (N_12937,N_11913,N_11657);
and U12938 (N_12938,N_10089,N_11905);
and U12939 (N_12939,N_11819,N_11703);
nand U12940 (N_12940,N_11026,N_11141);
nor U12941 (N_12941,N_11579,N_11685);
nor U12942 (N_12942,N_10279,N_10629);
xor U12943 (N_12943,N_11075,N_10410);
xor U12944 (N_12944,N_10109,N_10616);
xnor U12945 (N_12945,N_11990,N_10536);
and U12946 (N_12946,N_10451,N_11795);
nand U12947 (N_12947,N_10344,N_11040);
nor U12948 (N_12948,N_10384,N_11807);
xor U12949 (N_12949,N_11183,N_11705);
and U12950 (N_12950,N_11426,N_11424);
nand U12951 (N_12951,N_11498,N_10674);
xor U12952 (N_12952,N_10717,N_11785);
or U12953 (N_12953,N_11132,N_10746);
nor U12954 (N_12954,N_10970,N_10646);
or U12955 (N_12955,N_10823,N_10847);
and U12956 (N_12956,N_11063,N_11460);
nor U12957 (N_12957,N_10474,N_10600);
xor U12958 (N_12958,N_11578,N_10779);
or U12959 (N_12959,N_11156,N_10149);
and U12960 (N_12960,N_11519,N_10857);
nor U12961 (N_12961,N_11346,N_10822);
and U12962 (N_12962,N_11644,N_10960);
or U12963 (N_12963,N_10237,N_10851);
nor U12964 (N_12964,N_10635,N_10363);
nand U12965 (N_12965,N_10235,N_11854);
or U12966 (N_12966,N_10833,N_11581);
and U12967 (N_12967,N_10521,N_10827);
or U12968 (N_12968,N_10767,N_11808);
nor U12969 (N_12969,N_11223,N_11392);
nand U12970 (N_12970,N_10239,N_10404);
nand U12971 (N_12971,N_11192,N_10500);
and U12972 (N_12972,N_10372,N_10836);
and U12973 (N_12973,N_10887,N_11340);
nor U12974 (N_12974,N_10303,N_11296);
nand U12975 (N_12975,N_10554,N_11624);
and U12976 (N_12976,N_11363,N_11385);
or U12977 (N_12977,N_10680,N_11882);
and U12978 (N_12978,N_10658,N_11813);
or U12979 (N_12979,N_11728,N_10699);
nand U12980 (N_12980,N_10880,N_10815);
nand U12981 (N_12981,N_11735,N_10127);
xnor U12982 (N_12982,N_10269,N_10529);
or U12983 (N_12983,N_11473,N_10666);
xnor U12984 (N_12984,N_10202,N_10693);
nand U12985 (N_12985,N_10402,N_10804);
nor U12986 (N_12986,N_11469,N_11055);
and U12987 (N_12987,N_11215,N_10506);
nand U12988 (N_12988,N_11843,N_10971);
nor U12989 (N_12989,N_11744,N_10343);
xor U12990 (N_12990,N_11668,N_11553);
or U12991 (N_12991,N_11076,N_10701);
nor U12992 (N_12992,N_11707,N_10039);
nand U12993 (N_12993,N_10188,N_10234);
or U12994 (N_12994,N_10427,N_10765);
and U12995 (N_12995,N_10672,N_10820);
xnor U12996 (N_12996,N_10231,N_11732);
xnor U12997 (N_12997,N_10047,N_10494);
nand U12998 (N_12998,N_10429,N_10588);
xor U12999 (N_12999,N_10315,N_10167);
nor U13000 (N_13000,N_11458,N_10820);
xor U13001 (N_13001,N_10275,N_11676);
or U13002 (N_13002,N_10190,N_11692);
nor U13003 (N_13003,N_10635,N_11725);
nand U13004 (N_13004,N_10154,N_11556);
and U13005 (N_13005,N_11485,N_10581);
or U13006 (N_13006,N_10899,N_10761);
nand U13007 (N_13007,N_10987,N_10893);
or U13008 (N_13008,N_10858,N_11894);
xnor U13009 (N_13009,N_11691,N_11453);
xor U13010 (N_13010,N_10316,N_11704);
nor U13011 (N_13011,N_10805,N_11018);
nand U13012 (N_13012,N_10475,N_10272);
nand U13013 (N_13013,N_10088,N_11956);
nor U13014 (N_13014,N_10242,N_11526);
or U13015 (N_13015,N_10247,N_10634);
or U13016 (N_13016,N_10028,N_11232);
or U13017 (N_13017,N_11223,N_11467);
or U13018 (N_13018,N_11793,N_10625);
nand U13019 (N_13019,N_10076,N_11257);
and U13020 (N_13020,N_10700,N_11431);
nor U13021 (N_13021,N_11579,N_11867);
xor U13022 (N_13022,N_11904,N_11053);
nand U13023 (N_13023,N_11743,N_11430);
or U13024 (N_13024,N_10598,N_10682);
xnor U13025 (N_13025,N_11470,N_11889);
and U13026 (N_13026,N_10389,N_10436);
or U13027 (N_13027,N_11014,N_11651);
nand U13028 (N_13028,N_11817,N_10060);
nor U13029 (N_13029,N_11651,N_11946);
or U13030 (N_13030,N_11005,N_11462);
and U13031 (N_13031,N_10806,N_10326);
nor U13032 (N_13032,N_11415,N_11408);
and U13033 (N_13033,N_10681,N_10866);
xor U13034 (N_13034,N_11348,N_11559);
nor U13035 (N_13035,N_10096,N_10955);
xor U13036 (N_13036,N_10133,N_10329);
nor U13037 (N_13037,N_11874,N_10799);
nand U13038 (N_13038,N_11500,N_10733);
and U13039 (N_13039,N_10851,N_11892);
xnor U13040 (N_13040,N_10822,N_11459);
or U13041 (N_13041,N_11586,N_10961);
and U13042 (N_13042,N_11091,N_11751);
xnor U13043 (N_13043,N_11928,N_10349);
and U13044 (N_13044,N_11158,N_11517);
or U13045 (N_13045,N_11050,N_11017);
nand U13046 (N_13046,N_11536,N_10101);
and U13047 (N_13047,N_10155,N_11383);
nand U13048 (N_13048,N_11353,N_10586);
and U13049 (N_13049,N_10402,N_10641);
or U13050 (N_13050,N_11896,N_11666);
nor U13051 (N_13051,N_10921,N_11163);
and U13052 (N_13052,N_10750,N_10243);
nand U13053 (N_13053,N_10135,N_10969);
nand U13054 (N_13054,N_11101,N_10613);
nor U13055 (N_13055,N_11665,N_11678);
and U13056 (N_13056,N_10891,N_11916);
or U13057 (N_13057,N_10897,N_11301);
nor U13058 (N_13058,N_11835,N_11108);
nand U13059 (N_13059,N_10495,N_11552);
nor U13060 (N_13060,N_11382,N_10112);
and U13061 (N_13061,N_11835,N_10200);
xnor U13062 (N_13062,N_10343,N_11393);
and U13063 (N_13063,N_10724,N_10553);
and U13064 (N_13064,N_11909,N_10807);
nand U13065 (N_13065,N_10303,N_10901);
and U13066 (N_13066,N_11142,N_10303);
xnor U13067 (N_13067,N_10620,N_10441);
and U13068 (N_13068,N_10877,N_11549);
and U13069 (N_13069,N_10646,N_10710);
nand U13070 (N_13070,N_10359,N_10191);
or U13071 (N_13071,N_10139,N_11806);
and U13072 (N_13072,N_11340,N_11585);
xor U13073 (N_13073,N_11427,N_10639);
xnor U13074 (N_13074,N_10925,N_10403);
nor U13075 (N_13075,N_11903,N_11563);
nand U13076 (N_13076,N_10557,N_10057);
and U13077 (N_13077,N_10050,N_11607);
nand U13078 (N_13078,N_10538,N_10506);
nor U13079 (N_13079,N_10273,N_11193);
nand U13080 (N_13080,N_10568,N_11738);
or U13081 (N_13081,N_11291,N_10364);
and U13082 (N_13082,N_10094,N_11102);
nand U13083 (N_13083,N_11917,N_11569);
nor U13084 (N_13084,N_10542,N_11250);
or U13085 (N_13085,N_10887,N_11577);
nor U13086 (N_13086,N_10646,N_10827);
nor U13087 (N_13087,N_11589,N_11441);
nand U13088 (N_13088,N_10295,N_10148);
or U13089 (N_13089,N_10508,N_11497);
nor U13090 (N_13090,N_11097,N_11397);
nand U13091 (N_13091,N_10621,N_11855);
and U13092 (N_13092,N_10451,N_11878);
xor U13093 (N_13093,N_10633,N_10934);
xor U13094 (N_13094,N_10400,N_11748);
and U13095 (N_13095,N_11638,N_10789);
or U13096 (N_13096,N_11981,N_10252);
xnor U13097 (N_13097,N_10124,N_11000);
nand U13098 (N_13098,N_11165,N_11574);
nand U13099 (N_13099,N_10997,N_10542);
or U13100 (N_13100,N_11611,N_10167);
and U13101 (N_13101,N_10447,N_10376);
and U13102 (N_13102,N_10771,N_11166);
or U13103 (N_13103,N_10942,N_10748);
nor U13104 (N_13104,N_10366,N_11136);
xnor U13105 (N_13105,N_10896,N_11961);
and U13106 (N_13106,N_10913,N_11549);
nor U13107 (N_13107,N_11108,N_10462);
nand U13108 (N_13108,N_11745,N_11452);
or U13109 (N_13109,N_11478,N_11192);
nor U13110 (N_13110,N_11880,N_11059);
nor U13111 (N_13111,N_10810,N_11208);
nor U13112 (N_13112,N_10344,N_11973);
nand U13113 (N_13113,N_11677,N_11900);
and U13114 (N_13114,N_10542,N_11792);
nor U13115 (N_13115,N_10381,N_11523);
or U13116 (N_13116,N_11485,N_10363);
or U13117 (N_13117,N_10902,N_10037);
nor U13118 (N_13118,N_11111,N_11493);
xor U13119 (N_13119,N_11614,N_10592);
or U13120 (N_13120,N_10628,N_10783);
or U13121 (N_13121,N_11563,N_11041);
xor U13122 (N_13122,N_10961,N_10860);
and U13123 (N_13123,N_11785,N_10351);
or U13124 (N_13124,N_11163,N_11063);
or U13125 (N_13125,N_10785,N_11302);
nand U13126 (N_13126,N_10249,N_10877);
nand U13127 (N_13127,N_11223,N_11500);
or U13128 (N_13128,N_11658,N_10753);
xnor U13129 (N_13129,N_11657,N_11058);
and U13130 (N_13130,N_11827,N_11256);
or U13131 (N_13131,N_11568,N_11127);
and U13132 (N_13132,N_11523,N_10454);
or U13133 (N_13133,N_11834,N_10867);
and U13134 (N_13134,N_10606,N_10320);
nand U13135 (N_13135,N_10860,N_11612);
or U13136 (N_13136,N_11476,N_10946);
nand U13137 (N_13137,N_10194,N_11934);
xnor U13138 (N_13138,N_11829,N_11962);
xor U13139 (N_13139,N_11030,N_10190);
xor U13140 (N_13140,N_10282,N_10061);
or U13141 (N_13141,N_10141,N_11050);
xnor U13142 (N_13142,N_10158,N_11663);
xor U13143 (N_13143,N_10107,N_11375);
xnor U13144 (N_13144,N_10568,N_11314);
or U13145 (N_13145,N_11233,N_10577);
and U13146 (N_13146,N_11634,N_11567);
xor U13147 (N_13147,N_10657,N_10968);
nor U13148 (N_13148,N_10194,N_10995);
or U13149 (N_13149,N_10448,N_10593);
nor U13150 (N_13150,N_11551,N_10138);
nand U13151 (N_13151,N_11551,N_11443);
or U13152 (N_13152,N_11483,N_10954);
nor U13153 (N_13153,N_10709,N_11586);
and U13154 (N_13154,N_10288,N_11953);
nor U13155 (N_13155,N_11614,N_10403);
or U13156 (N_13156,N_10247,N_10714);
xnor U13157 (N_13157,N_10177,N_11162);
nor U13158 (N_13158,N_10417,N_10619);
nor U13159 (N_13159,N_11673,N_10262);
or U13160 (N_13160,N_11157,N_11325);
xor U13161 (N_13161,N_11375,N_10980);
nand U13162 (N_13162,N_10547,N_10010);
nand U13163 (N_13163,N_11532,N_11331);
or U13164 (N_13164,N_11022,N_11267);
nand U13165 (N_13165,N_11954,N_11136);
xor U13166 (N_13166,N_11064,N_11193);
nor U13167 (N_13167,N_11345,N_11580);
and U13168 (N_13168,N_11800,N_11224);
xnor U13169 (N_13169,N_10145,N_11518);
nor U13170 (N_13170,N_10684,N_10210);
or U13171 (N_13171,N_10162,N_11019);
and U13172 (N_13172,N_10624,N_10303);
xnor U13173 (N_13173,N_10095,N_11833);
or U13174 (N_13174,N_10222,N_11320);
nand U13175 (N_13175,N_10126,N_11732);
nand U13176 (N_13176,N_11268,N_11387);
nand U13177 (N_13177,N_10655,N_10567);
nand U13178 (N_13178,N_11202,N_11272);
nand U13179 (N_13179,N_10551,N_11193);
xor U13180 (N_13180,N_10628,N_11111);
nand U13181 (N_13181,N_11126,N_11050);
nor U13182 (N_13182,N_11588,N_11926);
and U13183 (N_13183,N_10720,N_11229);
and U13184 (N_13184,N_10711,N_10649);
and U13185 (N_13185,N_11280,N_11366);
nor U13186 (N_13186,N_10155,N_11937);
and U13187 (N_13187,N_10343,N_10708);
and U13188 (N_13188,N_10843,N_10624);
or U13189 (N_13189,N_10110,N_11675);
and U13190 (N_13190,N_10265,N_11436);
nand U13191 (N_13191,N_10277,N_10889);
nor U13192 (N_13192,N_11217,N_10230);
and U13193 (N_13193,N_10577,N_10565);
nor U13194 (N_13194,N_10659,N_10848);
nor U13195 (N_13195,N_10647,N_10460);
nand U13196 (N_13196,N_10316,N_11702);
and U13197 (N_13197,N_10278,N_10992);
and U13198 (N_13198,N_10825,N_11381);
and U13199 (N_13199,N_11626,N_11831);
or U13200 (N_13200,N_10430,N_10926);
nor U13201 (N_13201,N_11109,N_11826);
nor U13202 (N_13202,N_10979,N_10031);
nand U13203 (N_13203,N_11466,N_10276);
or U13204 (N_13204,N_10326,N_11931);
nor U13205 (N_13205,N_10028,N_10389);
nor U13206 (N_13206,N_10587,N_10924);
and U13207 (N_13207,N_10125,N_10023);
and U13208 (N_13208,N_10079,N_11084);
or U13209 (N_13209,N_11215,N_10171);
nand U13210 (N_13210,N_10630,N_11000);
xnor U13211 (N_13211,N_10925,N_11254);
nand U13212 (N_13212,N_10496,N_10529);
and U13213 (N_13213,N_11475,N_11257);
nor U13214 (N_13214,N_10266,N_10090);
nor U13215 (N_13215,N_10501,N_11300);
nand U13216 (N_13216,N_11988,N_10002);
or U13217 (N_13217,N_11472,N_11893);
nand U13218 (N_13218,N_11337,N_10603);
nor U13219 (N_13219,N_11901,N_11087);
xor U13220 (N_13220,N_11456,N_10456);
or U13221 (N_13221,N_10841,N_11597);
nand U13222 (N_13222,N_11335,N_11460);
and U13223 (N_13223,N_11805,N_10047);
xnor U13224 (N_13224,N_11593,N_11553);
nand U13225 (N_13225,N_10900,N_10385);
or U13226 (N_13226,N_10619,N_10677);
xnor U13227 (N_13227,N_11669,N_11747);
or U13228 (N_13228,N_10678,N_11795);
nor U13229 (N_13229,N_10275,N_11080);
nand U13230 (N_13230,N_11258,N_10160);
nor U13231 (N_13231,N_10432,N_11582);
xnor U13232 (N_13232,N_10342,N_10204);
nand U13233 (N_13233,N_11434,N_10122);
nand U13234 (N_13234,N_11447,N_11405);
nor U13235 (N_13235,N_11711,N_10455);
xor U13236 (N_13236,N_10407,N_11043);
xnor U13237 (N_13237,N_10505,N_11457);
and U13238 (N_13238,N_10483,N_10983);
nor U13239 (N_13239,N_10649,N_11206);
nand U13240 (N_13240,N_10058,N_11517);
xor U13241 (N_13241,N_11570,N_10570);
or U13242 (N_13242,N_11624,N_10273);
and U13243 (N_13243,N_11905,N_10643);
nor U13244 (N_13244,N_11386,N_11756);
xnor U13245 (N_13245,N_11092,N_11325);
or U13246 (N_13246,N_10614,N_10228);
xnor U13247 (N_13247,N_11397,N_10639);
and U13248 (N_13248,N_10188,N_11389);
nand U13249 (N_13249,N_11792,N_10833);
and U13250 (N_13250,N_11679,N_11803);
nand U13251 (N_13251,N_11691,N_10470);
nor U13252 (N_13252,N_10223,N_10279);
nor U13253 (N_13253,N_11175,N_11751);
and U13254 (N_13254,N_11038,N_11004);
and U13255 (N_13255,N_10008,N_11156);
nand U13256 (N_13256,N_10256,N_11951);
or U13257 (N_13257,N_10222,N_10096);
nand U13258 (N_13258,N_11358,N_11799);
or U13259 (N_13259,N_10950,N_10867);
xor U13260 (N_13260,N_10267,N_11282);
or U13261 (N_13261,N_10883,N_11677);
xor U13262 (N_13262,N_11569,N_11426);
and U13263 (N_13263,N_11640,N_11120);
or U13264 (N_13264,N_11528,N_10127);
xor U13265 (N_13265,N_10299,N_10616);
and U13266 (N_13266,N_10960,N_10362);
or U13267 (N_13267,N_11670,N_11622);
xor U13268 (N_13268,N_10276,N_11260);
and U13269 (N_13269,N_10311,N_10817);
or U13270 (N_13270,N_10975,N_10789);
xor U13271 (N_13271,N_11469,N_11356);
nor U13272 (N_13272,N_10634,N_10632);
nor U13273 (N_13273,N_11788,N_10432);
nand U13274 (N_13274,N_10792,N_11304);
or U13275 (N_13275,N_10873,N_11259);
nor U13276 (N_13276,N_10457,N_11323);
xnor U13277 (N_13277,N_11355,N_11309);
xnor U13278 (N_13278,N_11272,N_11362);
or U13279 (N_13279,N_10117,N_11638);
xor U13280 (N_13280,N_11142,N_11825);
nor U13281 (N_13281,N_10815,N_11216);
xor U13282 (N_13282,N_11791,N_10413);
xor U13283 (N_13283,N_10772,N_11660);
xor U13284 (N_13284,N_10298,N_10537);
or U13285 (N_13285,N_10364,N_11175);
or U13286 (N_13286,N_10840,N_10653);
or U13287 (N_13287,N_11375,N_10170);
and U13288 (N_13288,N_11819,N_11772);
or U13289 (N_13289,N_10117,N_10745);
nand U13290 (N_13290,N_10448,N_10683);
and U13291 (N_13291,N_11244,N_10656);
xor U13292 (N_13292,N_11291,N_11683);
nor U13293 (N_13293,N_11996,N_10697);
nor U13294 (N_13294,N_11740,N_10546);
or U13295 (N_13295,N_10011,N_10005);
nor U13296 (N_13296,N_10550,N_11675);
or U13297 (N_13297,N_10084,N_11808);
or U13298 (N_13298,N_10542,N_10306);
xor U13299 (N_13299,N_10925,N_10689);
and U13300 (N_13300,N_11442,N_11331);
nor U13301 (N_13301,N_10714,N_10619);
nor U13302 (N_13302,N_11289,N_10437);
and U13303 (N_13303,N_11245,N_10131);
nor U13304 (N_13304,N_11618,N_10179);
nand U13305 (N_13305,N_10799,N_11632);
and U13306 (N_13306,N_10788,N_10338);
xor U13307 (N_13307,N_11790,N_10618);
nand U13308 (N_13308,N_11395,N_10304);
or U13309 (N_13309,N_11319,N_10240);
nand U13310 (N_13310,N_10027,N_11844);
xor U13311 (N_13311,N_10951,N_11277);
nor U13312 (N_13312,N_10563,N_11862);
nand U13313 (N_13313,N_11331,N_11108);
nand U13314 (N_13314,N_11899,N_10469);
xnor U13315 (N_13315,N_11489,N_11070);
nand U13316 (N_13316,N_10860,N_10548);
and U13317 (N_13317,N_11174,N_11308);
and U13318 (N_13318,N_11485,N_10513);
nor U13319 (N_13319,N_10917,N_10912);
nand U13320 (N_13320,N_10852,N_11791);
nor U13321 (N_13321,N_10553,N_11523);
or U13322 (N_13322,N_11370,N_11545);
or U13323 (N_13323,N_11428,N_10211);
or U13324 (N_13324,N_11194,N_10823);
and U13325 (N_13325,N_11509,N_10790);
or U13326 (N_13326,N_11941,N_11613);
xnor U13327 (N_13327,N_10326,N_10459);
or U13328 (N_13328,N_11420,N_10931);
and U13329 (N_13329,N_11947,N_10018);
xnor U13330 (N_13330,N_10253,N_10746);
nand U13331 (N_13331,N_10031,N_11732);
xor U13332 (N_13332,N_10229,N_10055);
nor U13333 (N_13333,N_10423,N_11196);
xnor U13334 (N_13334,N_10848,N_10715);
nor U13335 (N_13335,N_11644,N_10578);
xor U13336 (N_13336,N_11789,N_11787);
nor U13337 (N_13337,N_10129,N_10370);
and U13338 (N_13338,N_11766,N_10023);
nand U13339 (N_13339,N_11822,N_11377);
and U13340 (N_13340,N_11857,N_10323);
nor U13341 (N_13341,N_10482,N_10504);
xor U13342 (N_13342,N_11868,N_11983);
xnor U13343 (N_13343,N_10230,N_10322);
or U13344 (N_13344,N_11157,N_10671);
or U13345 (N_13345,N_11223,N_10713);
nor U13346 (N_13346,N_10800,N_11622);
nand U13347 (N_13347,N_11198,N_10708);
and U13348 (N_13348,N_10123,N_11189);
or U13349 (N_13349,N_11545,N_10527);
and U13350 (N_13350,N_11840,N_11123);
and U13351 (N_13351,N_10222,N_11210);
and U13352 (N_13352,N_11498,N_10457);
and U13353 (N_13353,N_11032,N_10543);
and U13354 (N_13354,N_11498,N_11666);
nand U13355 (N_13355,N_11508,N_10952);
xnor U13356 (N_13356,N_11159,N_10579);
nand U13357 (N_13357,N_10708,N_10796);
nor U13358 (N_13358,N_10808,N_11579);
nand U13359 (N_13359,N_11950,N_11369);
nand U13360 (N_13360,N_11189,N_11313);
nand U13361 (N_13361,N_10885,N_10097);
nor U13362 (N_13362,N_10902,N_11894);
and U13363 (N_13363,N_10973,N_10991);
nor U13364 (N_13364,N_11691,N_10799);
nor U13365 (N_13365,N_11851,N_11895);
and U13366 (N_13366,N_10078,N_11584);
xor U13367 (N_13367,N_11213,N_10080);
nor U13368 (N_13368,N_10526,N_11239);
or U13369 (N_13369,N_11950,N_11598);
and U13370 (N_13370,N_10108,N_10167);
xnor U13371 (N_13371,N_11735,N_11213);
and U13372 (N_13372,N_10714,N_10573);
nor U13373 (N_13373,N_10431,N_10698);
nor U13374 (N_13374,N_10760,N_10965);
xor U13375 (N_13375,N_10865,N_11147);
or U13376 (N_13376,N_11856,N_10021);
nor U13377 (N_13377,N_10893,N_10003);
nor U13378 (N_13378,N_10607,N_11792);
xnor U13379 (N_13379,N_11977,N_10906);
and U13380 (N_13380,N_10991,N_11433);
nor U13381 (N_13381,N_11874,N_11550);
nor U13382 (N_13382,N_10052,N_10188);
nor U13383 (N_13383,N_10856,N_10656);
or U13384 (N_13384,N_10675,N_10301);
and U13385 (N_13385,N_11244,N_11767);
and U13386 (N_13386,N_11929,N_11735);
xor U13387 (N_13387,N_11804,N_11200);
nand U13388 (N_13388,N_11047,N_10587);
nor U13389 (N_13389,N_10841,N_10880);
xnor U13390 (N_13390,N_11901,N_11116);
or U13391 (N_13391,N_11368,N_10622);
xor U13392 (N_13392,N_11375,N_11610);
or U13393 (N_13393,N_10726,N_10579);
nand U13394 (N_13394,N_11566,N_10115);
and U13395 (N_13395,N_10596,N_11522);
or U13396 (N_13396,N_11150,N_10212);
or U13397 (N_13397,N_11726,N_11426);
and U13398 (N_13398,N_10801,N_10920);
xnor U13399 (N_13399,N_10873,N_10166);
nand U13400 (N_13400,N_10783,N_10208);
and U13401 (N_13401,N_10380,N_11336);
nand U13402 (N_13402,N_11703,N_10983);
or U13403 (N_13403,N_10542,N_10966);
and U13404 (N_13404,N_10783,N_11910);
nor U13405 (N_13405,N_10764,N_11927);
nand U13406 (N_13406,N_10091,N_10087);
xor U13407 (N_13407,N_11190,N_10881);
nand U13408 (N_13408,N_10109,N_10589);
and U13409 (N_13409,N_10905,N_10816);
nand U13410 (N_13410,N_11589,N_10990);
nor U13411 (N_13411,N_10601,N_11629);
nand U13412 (N_13412,N_11096,N_11656);
and U13413 (N_13413,N_11076,N_10260);
nor U13414 (N_13414,N_10610,N_11869);
nor U13415 (N_13415,N_11128,N_10931);
and U13416 (N_13416,N_10439,N_10437);
and U13417 (N_13417,N_11558,N_11289);
xnor U13418 (N_13418,N_10772,N_10555);
xor U13419 (N_13419,N_11044,N_11794);
nor U13420 (N_13420,N_11485,N_10210);
or U13421 (N_13421,N_10941,N_11536);
xor U13422 (N_13422,N_10142,N_11896);
or U13423 (N_13423,N_11060,N_11848);
or U13424 (N_13424,N_10332,N_10409);
xor U13425 (N_13425,N_10236,N_10905);
and U13426 (N_13426,N_10939,N_11947);
or U13427 (N_13427,N_10313,N_11799);
xor U13428 (N_13428,N_11031,N_10722);
xnor U13429 (N_13429,N_10790,N_10478);
and U13430 (N_13430,N_10862,N_10544);
xor U13431 (N_13431,N_11994,N_11170);
xnor U13432 (N_13432,N_11777,N_10527);
and U13433 (N_13433,N_10987,N_11613);
nor U13434 (N_13434,N_11113,N_10246);
xor U13435 (N_13435,N_10333,N_11070);
xor U13436 (N_13436,N_10541,N_11820);
nand U13437 (N_13437,N_11849,N_10070);
nor U13438 (N_13438,N_11648,N_11000);
nor U13439 (N_13439,N_10396,N_10496);
and U13440 (N_13440,N_10095,N_10152);
and U13441 (N_13441,N_11969,N_10833);
nor U13442 (N_13442,N_10531,N_10507);
nand U13443 (N_13443,N_11405,N_10581);
or U13444 (N_13444,N_10144,N_11031);
xor U13445 (N_13445,N_10451,N_11135);
nand U13446 (N_13446,N_11100,N_10450);
xnor U13447 (N_13447,N_11227,N_11918);
and U13448 (N_13448,N_11268,N_11768);
or U13449 (N_13449,N_10068,N_10149);
nor U13450 (N_13450,N_11284,N_11507);
nand U13451 (N_13451,N_10908,N_10037);
or U13452 (N_13452,N_11263,N_11147);
or U13453 (N_13453,N_10401,N_11742);
and U13454 (N_13454,N_10260,N_10344);
xor U13455 (N_13455,N_11872,N_10488);
or U13456 (N_13456,N_11087,N_11421);
and U13457 (N_13457,N_10833,N_11450);
nor U13458 (N_13458,N_10457,N_11849);
and U13459 (N_13459,N_11968,N_10186);
nand U13460 (N_13460,N_11610,N_10095);
or U13461 (N_13461,N_10514,N_11238);
and U13462 (N_13462,N_10658,N_10439);
nand U13463 (N_13463,N_10236,N_11245);
nand U13464 (N_13464,N_10012,N_11700);
xnor U13465 (N_13465,N_11488,N_10208);
nor U13466 (N_13466,N_10307,N_10107);
or U13467 (N_13467,N_11883,N_10307);
nor U13468 (N_13468,N_10877,N_11179);
or U13469 (N_13469,N_10837,N_10578);
nor U13470 (N_13470,N_11321,N_11200);
xor U13471 (N_13471,N_10738,N_10997);
nor U13472 (N_13472,N_11593,N_10310);
nand U13473 (N_13473,N_10495,N_10698);
nand U13474 (N_13474,N_11841,N_10047);
nand U13475 (N_13475,N_11380,N_11598);
nor U13476 (N_13476,N_11271,N_11779);
nor U13477 (N_13477,N_10147,N_11975);
and U13478 (N_13478,N_10148,N_10163);
and U13479 (N_13479,N_10195,N_10404);
nor U13480 (N_13480,N_10392,N_10882);
nand U13481 (N_13481,N_11524,N_10562);
and U13482 (N_13482,N_11128,N_10664);
nand U13483 (N_13483,N_10827,N_11652);
or U13484 (N_13484,N_10140,N_10952);
nand U13485 (N_13485,N_11113,N_11962);
xnor U13486 (N_13486,N_11443,N_10679);
nand U13487 (N_13487,N_10837,N_10539);
nand U13488 (N_13488,N_11615,N_10453);
or U13489 (N_13489,N_11514,N_11035);
xor U13490 (N_13490,N_10015,N_10913);
nand U13491 (N_13491,N_11663,N_10763);
nor U13492 (N_13492,N_10916,N_10258);
and U13493 (N_13493,N_11954,N_11395);
nand U13494 (N_13494,N_10384,N_11400);
or U13495 (N_13495,N_11396,N_10529);
xnor U13496 (N_13496,N_11081,N_11815);
and U13497 (N_13497,N_11008,N_11642);
or U13498 (N_13498,N_11179,N_11261);
or U13499 (N_13499,N_10189,N_11545);
nand U13500 (N_13500,N_11651,N_11757);
and U13501 (N_13501,N_11939,N_10995);
nor U13502 (N_13502,N_11600,N_10736);
or U13503 (N_13503,N_10071,N_11525);
nor U13504 (N_13504,N_10796,N_11378);
or U13505 (N_13505,N_11172,N_11642);
and U13506 (N_13506,N_10622,N_11971);
or U13507 (N_13507,N_11782,N_11454);
nor U13508 (N_13508,N_10878,N_11253);
nor U13509 (N_13509,N_11860,N_10821);
nor U13510 (N_13510,N_11678,N_11764);
nor U13511 (N_13511,N_11973,N_10090);
nand U13512 (N_13512,N_10944,N_10945);
or U13513 (N_13513,N_11251,N_11908);
nor U13514 (N_13514,N_10396,N_10973);
xnor U13515 (N_13515,N_10390,N_11414);
and U13516 (N_13516,N_10252,N_10294);
xor U13517 (N_13517,N_11802,N_11968);
or U13518 (N_13518,N_11027,N_10810);
nand U13519 (N_13519,N_10501,N_10154);
nand U13520 (N_13520,N_11588,N_10105);
and U13521 (N_13521,N_11828,N_10249);
xnor U13522 (N_13522,N_10685,N_10648);
and U13523 (N_13523,N_11335,N_10147);
or U13524 (N_13524,N_11326,N_10551);
xnor U13525 (N_13525,N_10386,N_10198);
nand U13526 (N_13526,N_11877,N_10694);
or U13527 (N_13527,N_10437,N_10562);
or U13528 (N_13528,N_10997,N_10052);
nand U13529 (N_13529,N_10971,N_11579);
nor U13530 (N_13530,N_10964,N_11865);
xor U13531 (N_13531,N_10221,N_10432);
nor U13532 (N_13532,N_10884,N_10900);
and U13533 (N_13533,N_11328,N_11782);
nor U13534 (N_13534,N_11127,N_11326);
or U13535 (N_13535,N_11247,N_10894);
xor U13536 (N_13536,N_10768,N_11217);
nand U13537 (N_13537,N_10957,N_11353);
nor U13538 (N_13538,N_11736,N_11045);
nor U13539 (N_13539,N_11280,N_11134);
xnor U13540 (N_13540,N_11457,N_10014);
xor U13541 (N_13541,N_10155,N_10277);
xnor U13542 (N_13542,N_10436,N_11519);
nor U13543 (N_13543,N_10813,N_11384);
xnor U13544 (N_13544,N_11556,N_10570);
and U13545 (N_13545,N_10360,N_10366);
nand U13546 (N_13546,N_10435,N_11129);
and U13547 (N_13547,N_10265,N_11869);
nor U13548 (N_13548,N_10202,N_10798);
nor U13549 (N_13549,N_10253,N_10696);
nor U13550 (N_13550,N_10972,N_11478);
nor U13551 (N_13551,N_11801,N_11928);
nand U13552 (N_13552,N_10527,N_11396);
or U13553 (N_13553,N_10413,N_11355);
or U13554 (N_13554,N_11409,N_11553);
or U13555 (N_13555,N_11903,N_11522);
xor U13556 (N_13556,N_10338,N_11514);
nand U13557 (N_13557,N_10033,N_11338);
nor U13558 (N_13558,N_11356,N_10936);
and U13559 (N_13559,N_11773,N_10004);
or U13560 (N_13560,N_10859,N_10576);
or U13561 (N_13561,N_11702,N_10422);
and U13562 (N_13562,N_10693,N_11964);
xnor U13563 (N_13563,N_11519,N_11454);
nor U13564 (N_13564,N_11109,N_10246);
nand U13565 (N_13565,N_10053,N_10809);
and U13566 (N_13566,N_10359,N_11525);
nand U13567 (N_13567,N_11027,N_10425);
or U13568 (N_13568,N_11021,N_11594);
or U13569 (N_13569,N_11319,N_10242);
xor U13570 (N_13570,N_11650,N_10373);
xnor U13571 (N_13571,N_10928,N_11156);
and U13572 (N_13572,N_11095,N_11497);
nand U13573 (N_13573,N_11811,N_11117);
and U13574 (N_13574,N_11068,N_11429);
or U13575 (N_13575,N_11126,N_10251);
nand U13576 (N_13576,N_11458,N_10295);
or U13577 (N_13577,N_10214,N_11646);
and U13578 (N_13578,N_10377,N_10066);
and U13579 (N_13579,N_11279,N_10821);
and U13580 (N_13580,N_10528,N_11199);
xnor U13581 (N_13581,N_10425,N_11587);
nand U13582 (N_13582,N_11855,N_10416);
xnor U13583 (N_13583,N_11662,N_10504);
nor U13584 (N_13584,N_10423,N_11289);
or U13585 (N_13585,N_11859,N_11971);
or U13586 (N_13586,N_10784,N_10530);
xor U13587 (N_13587,N_10572,N_11121);
or U13588 (N_13588,N_10600,N_10155);
nand U13589 (N_13589,N_10395,N_11747);
nand U13590 (N_13590,N_11207,N_10102);
xnor U13591 (N_13591,N_10478,N_11845);
xor U13592 (N_13592,N_11903,N_11037);
nand U13593 (N_13593,N_11184,N_11296);
nand U13594 (N_13594,N_11222,N_10183);
or U13595 (N_13595,N_10213,N_10342);
and U13596 (N_13596,N_11326,N_10078);
nand U13597 (N_13597,N_11119,N_11414);
or U13598 (N_13598,N_10057,N_10480);
nor U13599 (N_13599,N_10299,N_11159);
nand U13600 (N_13600,N_10816,N_10220);
nand U13601 (N_13601,N_11569,N_11926);
and U13602 (N_13602,N_10072,N_11008);
xnor U13603 (N_13603,N_10671,N_11894);
and U13604 (N_13604,N_10872,N_11257);
nor U13605 (N_13605,N_10689,N_10439);
nor U13606 (N_13606,N_11641,N_10163);
xor U13607 (N_13607,N_10724,N_11498);
and U13608 (N_13608,N_11778,N_10112);
nor U13609 (N_13609,N_11264,N_10834);
xnor U13610 (N_13610,N_11624,N_10685);
xnor U13611 (N_13611,N_10718,N_11548);
or U13612 (N_13612,N_10851,N_11377);
xnor U13613 (N_13613,N_10332,N_11822);
and U13614 (N_13614,N_10405,N_10318);
nor U13615 (N_13615,N_11588,N_10485);
nand U13616 (N_13616,N_10744,N_11565);
xor U13617 (N_13617,N_11985,N_10494);
xor U13618 (N_13618,N_11935,N_11677);
nand U13619 (N_13619,N_11555,N_10462);
xnor U13620 (N_13620,N_10201,N_11393);
nor U13621 (N_13621,N_10434,N_11248);
and U13622 (N_13622,N_10900,N_11450);
nor U13623 (N_13623,N_11642,N_10741);
nand U13624 (N_13624,N_10055,N_11718);
and U13625 (N_13625,N_11989,N_10064);
or U13626 (N_13626,N_10958,N_11561);
xnor U13627 (N_13627,N_11216,N_10714);
nor U13628 (N_13628,N_10806,N_11797);
nor U13629 (N_13629,N_11975,N_11221);
nand U13630 (N_13630,N_11137,N_11800);
xor U13631 (N_13631,N_11258,N_10440);
or U13632 (N_13632,N_10422,N_11617);
nand U13633 (N_13633,N_10792,N_11582);
nand U13634 (N_13634,N_10776,N_11685);
xnor U13635 (N_13635,N_10447,N_11165);
xnor U13636 (N_13636,N_11581,N_11445);
and U13637 (N_13637,N_10880,N_10760);
or U13638 (N_13638,N_11808,N_11356);
nand U13639 (N_13639,N_10766,N_11550);
xnor U13640 (N_13640,N_10392,N_10496);
nand U13641 (N_13641,N_10992,N_11077);
or U13642 (N_13642,N_11281,N_10912);
xnor U13643 (N_13643,N_10479,N_11846);
and U13644 (N_13644,N_11434,N_10365);
and U13645 (N_13645,N_10071,N_11917);
and U13646 (N_13646,N_10475,N_10884);
and U13647 (N_13647,N_10269,N_11834);
or U13648 (N_13648,N_11697,N_11783);
or U13649 (N_13649,N_10273,N_11662);
xnor U13650 (N_13650,N_11771,N_10642);
nor U13651 (N_13651,N_11584,N_10585);
xnor U13652 (N_13652,N_11325,N_10854);
or U13653 (N_13653,N_11392,N_10981);
and U13654 (N_13654,N_11208,N_11461);
and U13655 (N_13655,N_11437,N_11182);
nor U13656 (N_13656,N_10789,N_11743);
xor U13657 (N_13657,N_10761,N_10139);
nor U13658 (N_13658,N_11884,N_11246);
nor U13659 (N_13659,N_11503,N_10340);
xor U13660 (N_13660,N_11660,N_10365);
or U13661 (N_13661,N_11263,N_10038);
or U13662 (N_13662,N_10338,N_11737);
xnor U13663 (N_13663,N_11583,N_10064);
or U13664 (N_13664,N_11750,N_11858);
nor U13665 (N_13665,N_11856,N_10799);
xor U13666 (N_13666,N_11437,N_11003);
and U13667 (N_13667,N_11004,N_11408);
and U13668 (N_13668,N_10730,N_10848);
nand U13669 (N_13669,N_10479,N_11963);
or U13670 (N_13670,N_11470,N_10341);
nor U13671 (N_13671,N_11174,N_11131);
nand U13672 (N_13672,N_11200,N_10019);
xnor U13673 (N_13673,N_11327,N_11138);
or U13674 (N_13674,N_10858,N_11450);
nor U13675 (N_13675,N_10394,N_11429);
and U13676 (N_13676,N_11371,N_11994);
or U13677 (N_13677,N_10380,N_11563);
or U13678 (N_13678,N_10171,N_11612);
or U13679 (N_13679,N_10887,N_10257);
or U13680 (N_13680,N_11517,N_10957);
or U13681 (N_13681,N_11803,N_11413);
xnor U13682 (N_13682,N_11819,N_10798);
and U13683 (N_13683,N_11359,N_11198);
xnor U13684 (N_13684,N_10247,N_10828);
nand U13685 (N_13685,N_11679,N_10415);
nand U13686 (N_13686,N_10355,N_11622);
or U13687 (N_13687,N_10014,N_10336);
nor U13688 (N_13688,N_11013,N_10168);
nor U13689 (N_13689,N_10025,N_10059);
and U13690 (N_13690,N_11795,N_11278);
or U13691 (N_13691,N_10980,N_11630);
and U13692 (N_13692,N_10741,N_10863);
nand U13693 (N_13693,N_10907,N_10599);
or U13694 (N_13694,N_10889,N_11613);
nand U13695 (N_13695,N_10793,N_10272);
xnor U13696 (N_13696,N_10340,N_11693);
or U13697 (N_13697,N_10826,N_11603);
and U13698 (N_13698,N_11062,N_10118);
nor U13699 (N_13699,N_10104,N_10871);
nor U13700 (N_13700,N_10517,N_11796);
xnor U13701 (N_13701,N_11350,N_11161);
xor U13702 (N_13702,N_11010,N_10165);
nand U13703 (N_13703,N_11513,N_10122);
xnor U13704 (N_13704,N_11879,N_11114);
nor U13705 (N_13705,N_10789,N_11224);
xnor U13706 (N_13706,N_10586,N_11697);
or U13707 (N_13707,N_11236,N_10633);
nor U13708 (N_13708,N_11002,N_10505);
nand U13709 (N_13709,N_11198,N_10287);
xor U13710 (N_13710,N_11231,N_10111);
nor U13711 (N_13711,N_11613,N_11057);
or U13712 (N_13712,N_11001,N_10921);
nand U13713 (N_13713,N_11048,N_11881);
nand U13714 (N_13714,N_10488,N_11650);
xor U13715 (N_13715,N_11861,N_11882);
nand U13716 (N_13716,N_11959,N_11949);
or U13717 (N_13717,N_10733,N_10541);
and U13718 (N_13718,N_11198,N_10712);
or U13719 (N_13719,N_11139,N_11551);
and U13720 (N_13720,N_11502,N_10520);
nand U13721 (N_13721,N_11212,N_10688);
nor U13722 (N_13722,N_10803,N_11167);
nand U13723 (N_13723,N_10226,N_10572);
and U13724 (N_13724,N_11576,N_11167);
and U13725 (N_13725,N_11326,N_11188);
nor U13726 (N_13726,N_10686,N_11455);
nor U13727 (N_13727,N_10990,N_11448);
xor U13728 (N_13728,N_11377,N_10464);
nor U13729 (N_13729,N_10761,N_11550);
or U13730 (N_13730,N_10095,N_10790);
nand U13731 (N_13731,N_11675,N_10974);
nor U13732 (N_13732,N_10734,N_11001);
nand U13733 (N_13733,N_10551,N_10083);
xor U13734 (N_13734,N_10811,N_10846);
or U13735 (N_13735,N_10551,N_11608);
nand U13736 (N_13736,N_10801,N_10063);
xnor U13737 (N_13737,N_11271,N_10002);
or U13738 (N_13738,N_10525,N_11795);
and U13739 (N_13739,N_11980,N_11190);
and U13740 (N_13740,N_10052,N_10989);
and U13741 (N_13741,N_11476,N_11977);
nand U13742 (N_13742,N_10238,N_11308);
or U13743 (N_13743,N_11888,N_11337);
xor U13744 (N_13744,N_11950,N_11065);
nor U13745 (N_13745,N_10346,N_11885);
or U13746 (N_13746,N_10299,N_11139);
nor U13747 (N_13747,N_10152,N_11192);
and U13748 (N_13748,N_11835,N_10829);
xnor U13749 (N_13749,N_11005,N_11094);
nand U13750 (N_13750,N_10348,N_10948);
and U13751 (N_13751,N_10309,N_11238);
or U13752 (N_13752,N_11542,N_11338);
or U13753 (N_13753,N_10066,N_11201);
nor U13754 (N_13754,N_11295,N_10955);
nor U13755 (N_13755,N_11095,N_10495);
or U13756 (N_13756,N_11019,N_10840);
nand U13757 (N_13757,N_10778,N_11794);
xnor U13758 (N_13758,N_10829,N_10217);
xor U13759 (N_13759,N_10361,N_10788);
or U13760 (N_13760,N_11687,N_11785);
and U13761 (N_13761,N_10686,N_10440);
nor U13762 (N_13762,N_10523,N_10558);
xor U13763 (N_13763,N_10282,N_10447);
and U13764 (N_13764,N_10222,N_11097);
and U13765 (N_13765,N_11289,N_11606);
and U13766 (N_13766,N_11337,N_11469);
nand U13767 (N_13767,N_10225,N_11910);
nor U13768 (N_13768,N_10521,N_10114);
or U13769 (N_13769,N_11532,N_11641);
or U13770 (N_13770,N_10685,N_10765);
xnor U13771 (N_13771,N_10889,N_11375);
nand U13772 (N_13772,N_11607,N_11687);
nand U13773 (N_13773,N_11246,N_10617);
nor U13774 (N_13774,N_11254,N_10623);
nor U13775 (N_13775,N_11087,N_10291);
nor U13776 (N_13776,N_11768,N_11589);
or U13777 (N_13777,N_10548,N_11234);
or U13778 (N_13778,N_11992,N_11739);
and U13779 (N_13779,N_10844,N_10057);
nand U13780 (N_13780,N_10196,N_10154);
xnor U13781 (N_13781,N_11625,N_10658);
or U13782 (N_13782,N_10499,N_10195);
or U13783 (N_13783,N_10047,N_10941);
nand U13784 (N_13784,N_10467,N_10749);
and U13785 (N_13785,N_11944,N_11279);
nand U13786 (N_13786,N_11276,N_10049);
xor U13787 (N_13787,N_11863,N_11874);
nor U13788 (N_13788,N_11581,N_11658);
xnor U13789 (N_13789,N_10914,N_11090);
nor U13790 (N_13790,N_10492,N_11049);
nand U13791 (N_13791,N_11831,N_11747);
nand U13792 (N_13792,N_10801,N_11736);
and U13793 (N_13793,N_10344,N_10298);
nand U13794 (N_13794,N_10942,N_11886);
nand U13795 (N_13795,N_11659,N_10409);
nand U13796 (N_13796,N_10057,N_10541);
or U13797 (N_13797,N_10616,N_11766);
and U13798 (N_13798,N_11019,N_11963);
and U13799 (N_13799,N_11685,N_10437);
and U13800 (N_13800,N_11917,N_11914);
nand U13801 (N_13801,N_10396,N_11663);
xnor U13802 (N_13802,N_11917,N_11033);
and U13803 (N_13803,N_11192,N_10852);
xnor U13804 (N_13804,N_10349,N_10029);
or U13805 (N_13805,N_11567,N_10323);
nor U13806 (N_13806,N_10701,N_11412);
xnor U13807 (N_13807,N_10288,N_11253);
or U13808 (N_13808,N_10556,N_11585);
nor U13809 (N_13809,N_10687,N_11244);
nor U13810 (N_13810,N_11624,N_11386);
nor U13811 (N_13811,N_11694,N_10524);
nand U13812 (N_13812,N_10454,N_11199);
and U13813 (N_13813,N_10927,N_11314);
nor U13814 (N_13814,N_10450,N_10318);
or U13815 (N_13815,N_10805,N_11588);
and U13816 (N_13816,N_10398,N_10432);
nand U13817 (N_13817,N_11184,N_10850);
nor U13818 (N_13818,N_10153,N_11483);
or U13819 (N_13819,N_11617,N_10134);
nand U13820 (N_13820,N_10912,N_10804);
or U13821 (N_13821,N_10402,N_10271);
nor U13822 (N_13822,N_11913,N_10809);
nand U13823 (N_13823,N_11828,N_11097);
nor U13824 (N_13824,N_10484,N_10258);
nor U13825 (N_13825,N_11180,N_10795);
nand U13826 (N_13826,N_10623,N_11788);
nor U13827 (N_13827,N_10187,N_11321);
xor U13828 (N_13828,N_10075,N_11150);
xor U13829 (N_13829,N_10068,N_10056);
xnor U13830 (N_13830,N_11204,N_11016);
or U13831 (N_13831,N_10471,N_10770);
and U13832 (N_13832,N_11848,N_10472);
or U13833 (N_13833,N_10037,N_11305);
nor U13834 (N_13834,N_10963,N_10329);
nor U13835 (N_13835,N_10412,N_10804);
or U13836 (N_13836,N_11183,N_10872);
and U13837 (N_13837,N_10399,N_11173);
nand U13838 (N_13838,N_10446,N_11890);
xor U13839 (N_13839,N_11952,N_11022);
xor U13840 (N_13840,N_10755,N_10499);
or U13841 (N_13841,N_10923,N_10041);
xor U13842 (N_13842,N_10421,N_11928);
xnor U13843 (N_13843,N_11401,N_11488);
or U13844 (N_13844,N_11717,N_11163);
nor U13845 (N_13845,N_11774,N_11514);
and U13846 (N_13846,N_11508,N_10581);
nand U13847 (N_13847,N_10492,N_11768);
xnor U13848 (N_13848,N_11424,N_11321);
or U13849 (N_13849,N_11691,N_11071);
nor U13850 (N_13850,N_11436,N_11968);
and U13851 (N_13851,N_10683,N_10710);
nand U13852 (N_13852,N_10680,N_10143);
and U13853 (N_13853,N_10920,N_11763);
or U13854 (N_13854,N_10034,N_11390);
or U13855 (N_13855,N_10215,N_11021);
or U13856 (N_13856,N_10254,N_10538);
or U13857 (N_13857,N_11388,N_10015);
nor U13858 (N_13858,N_10314,N_10797);
and U13859 (N_13859,N_10118,N_10629);
nand U13860 (N_13860,N_10879,N_11711);
nor U13861 (N_13861,N_11717,N_11822);
and U13862 (N_13862,N_10976,N_11471);
nor U13863 (N_13863,N_10987,N_10172);
nor U13864 (N_13864,N_10519,N_10169);
nor U13865 (N_13865,N_11999,N_11674);
or U13866 (N_13866,N_11756,N_11180);
xnor U13867 (N_13867,N_11993,N_11901);
nor U13868 (N_13868,N_10680,N_10907);
and U13869 (N_13869,N_10416,N_10955);
xor U13870 (N_13870,N_11877,N_11306);
and U13871 (N_13871,N_10660,N_11749);
nand U13872 (N_13872,N_11972,N_11672);
xor U13873 (N_13873,N_10962,N_10227);
nor U13874 (N_13874,N_10713,N_10872);
nand U13875 (N_13875,N_10984,N_11426);
and U13876 (N_13876,N_10225,N_11340);
or U13877 (N_13877,N_10005,N_11558);
xor U13878 (N_13878,N_11584,N_11853);
nand U13879 (N_13879,N_11850,N_10064);
or U13880 (N_13880,N_10553,N_10068);
xor U13881 (N_13881,N_11909,N_11424);
or U13882 (N_13882,N_10001,N_11222);
nor U13883 (N_13883,N_10556,N_10687);
nor U13884 (N_13884,N_10373,N_10128);
xor U13885 (N_13885,N_11363,N_10154);
xor U13886 (N_13886,N_10122,N_10176);
or U13887 (N_13887,N_10882,N_10345);
xor U13888 (N_13888,N_11380,N_11220);
or U13889 (N_13889,N_11294,N_10845);
nand U13890 (N_13890,N_11777,N_11910);
or U13891 (N_13891,N_10088,N_11480);
and U13892 (N_13892,N_10732,N_11424);
xor U13893 (N_13893,N_10787,N_11075);
or U13894 (N_13894,N_11589,N_10453);
nor U13895 (N_13895,N_10207,N_11422);
and U13896 (N_13896,N_10163,N_10468);
or U13897 (N_13897,N_10843,N_11967);
nor U13898 (N_13898,N_10084,N_11391);
xnor U13899 (N_13899,N_11484,N_11914);
or U13900 (N_13900,N_11534,N_10630);
xnor U13901 (N_13901,N_10592,N_10661);
xor U13902 (N_13902,N_11434,N_10079);
and U13903 (N_13903,N_11938,N_11520);
xor U13904 (N_13904,N_11633,N_10047);
nand U13905 (N_13905,N_11545,N_11309);
and U13906 (N_13906,N_10996,N_10599);
nor U13907 (N_13907,N_10002,N_11014);
xnor U13908 (N_13908,N_11582,N_11251);
xor U13909 (N_13909,N_11764,N_10452);
nand U13910 (N_13910,N_11452,N_11003);
or U13911 (N_13911,N_11080,N_10011);
and U13912 (N_13912,N_10942,N_11055);
or U13913 (N_13913,N_10288,N_10287);
and U13914 (N_13914,N_10981,N_11473);
nand U13915 (N_13915,N_11493,N_10199);
nor U13916 (N_13916,N_10910,N_11347);
xnor U13917 (N_13917,N_10578,N_11365);
nand U13918 (N_13918,N_11849,N_10617);
and U13919 (N_13919,N_10372,N_10894);
or U13920 (N_13920,N_10968,N_10656);
and U13921 (N_13921,N_11655,N_11041);
nand U13922 (N_13922,N_11964,N_11323);
or U13923 (N_13923,N_10144,N_11804);
and U13924 (N_13924,N_11626,N_11148);
and U13925 (N_13925,N_10187,N_11217);
nor U13926 (N_13926,N_10639,N_11306);
or U13927 (N_13927,N_11734,N_10181);
nand U13928 (N_13928,N_10761,N_11997);
or U13929 (N_13929,N_11048,N_10912);
and U13930 (N_13930,N_11575,N_11436);
nand U13931 (N_13931,N_10759,N_10818);
and U13932 (N_13932,N_11210,N_11742);
nand U13933 (N_13933,N_11601,N_10950);
xor U13934 (N_13934,N_10945,N_11992);
nand U13935 (N_13935,N_11362,N_10680);
and U13936 (N_13936,N_11968,N_10617);
nor U13937 (N_13937,N_11190,N_11058);
or U13938 (N_13938,N_11158,N_10859);
xor U13939 (N_13939,N_11577,N_10299);
xnor U13940 (N_13940,N_10026,N_10533);
xnor U13941 (N_13941,N_10493,N_10652);
nand U13942 (N_13942,N_10332,N_11664);
and U13943 (N_13943,N_10443,N_10832);
and U13944 (N_13944,N_11147,N_11868);
or U13945 (N_13945,N_11673,N_10108);
nand U13946 (N_13946,N_10611,N_10735);
or U13947 (N_13947,N_11129,N_10742);
and U13948 (N_13948,N_10078,N_10616);
or U13949 (N_13949,N_11659,N_10927);
or U13950 (N_13950,N_11900,N_10335);
or U13951 (N_13951,N_11416,N_10572);
xnor U13952 (N_13952,N_11401,N_10671);
and U13953 (N_13953,N_10986,N_10425);
nand U13954 (N_13954,N_10260,N_10421);
and U13955 (N_13955,N_10800,N_11291);
nand U13956 (N_13956,N_11914,N_10998);
nand U13957 (N_13957,N_11140,N_10797);
nand U13958 (N_13958,N_11321,N_10389);
or U13959 (N_13959,N_10376,N_11699);
and U13960 (N_13960,N_11519,N_10197);
or U13961 (N_13961,N_10685,N_11548);
nand U13962 (N_13962,N_11445,N_10351);
and U13963 (N_13963,N_10840,N_10172);
nor U13964 (N_13964,N_10724,N_11265);
and U13965 (N_13965,N_10702,N_11343);
xor U13966 (N_13966,N_11448,N_10292);
nor U13967 (N_13967,N_10561,N_10556);
and U13968 (N_13968,N_11122,N_10820);
xnor U13969 (N_13969,N_11338,N_10946);
or U13970 (N_13970,N_10040,N_10389);
and U13971 (N_13971,N_11953,N_10451);
xnor U13972 (N_13972,N_11889,N_11987);
nand U13973 (N_13973,N_11530,N_10761);
nor U13974 (N_13974,N_11705,N_10781);
nand U13975 (N_13975,N_10576,N_11149);
or U13976 (N_13976,N_11290,N_11474);
or U13977 (N_13977,N_11175,N_11453);
nand U13978 (N_13978,N_11517,N_10951);
and U13979 (N_13979,N_10010,N_10645);
or U13980 (N_13980,N_11672,N_10276);
nor U13981 (N_13981,N_11483,N_11902);
nand U13982 (N_13982,N_10521,N_10204);
xor U13983 (N_13983,N_10647,N_11569);
or U13984 (N_13984,N_11151,N_10928);
nor U13985 (N_13985,N_10023,N_10862);
or U13986 (N_13986,N_11810,N_11777);
and U13987 (N_13987,N_10439,N_11632);
or U13988 (N_13988,N_11189,N_11371);
nand U13989 (N_13989,N_11003,N_10432);
nand U13990 (N_13990,N_10430,N_11259);
xor U13991 (N_13991,N_11165,N_10478);
nand U13992 (N_13992,N_11686,N_10507);
nor U13993 (N_13993,N_11340,N_10404);
or U13994 (N_13994,N_10068,N_10173);
xnor U13995 (N_13995,N_11984,N_11299);
xnor U13996 (N_13996,N_10855,N_11190);
nand U13997 (N_13997,N_11016,N_11717);
and U13998 (N_13998,N_11515,N_10530);
and U13999 (N_13999,N_11271,N_10549);
xnor U14000 (N_14000,N_12979,N_12135);
nand U14001 (N_14001,N_13437,N_12369);
and U14002 (N_14002,N_12271,N_13443);
and U14003 (N_14003,N_12580,N_12280);
and U14004 (N_14004,N_13276,N_12416);
nand U14005 (N_14005,N_12449,N_13470);
nor U14006 (N_14006,N_13594,N_12187);
or U14007 (N_14007,N_13825,N_12037);
xor U14008 (N_14008,N_12503,N_12809);
and U14009 (N_14009,N_13273,N_12098);
or U14010 (N_14010,N_13182,N_13327);
or U14011 (N_14011,N_13923,N_12113);
xor U14012 (N_14012,N_13718,N_12013);
or U14013 (N_14013,N_12793,N_12070);
nor U14014 (N_14014,N_13572,N_13476);
and U14015 (N_14015,N_12907,N_12851);
nor U14016 (N_14016,N_13863,N_12519);
and U14017 (N_14017,N_13017,N_12870);
and U14018 (N_14018,N_12159,N_12983);
and U14019 (N_14019,N_13044,N_12530);
nor U14020 (N_14020,N_13577,N_13891);
xnor U14021 (N_14021,N_13786,N_13199);
nand U14022 (N_14022,N_13355,N_13085);
and U14023 (N_14023,N_13641,N_12458);
xor U14024 (N_14024,N_12996,N_12457);
nand U14025 (N_14025,N_13097,N_13219);
nand U14026 (N_14026,N_13388,N_12584);
xor U14027 (N_14027,N_13868,N_12840);
or U14028 (N_14028,N_13142,N_13463);
xnor U14029 (N_14029,N_12975,N_13560);
and U14030 (N_14030,N_13288,N_13481);
nand U14031 (N_14031,N_13191,N_12314);
xnor U14032 (N_14032,N_13499,N_13066);
nor U14033 (N_14033,N_12427,N_12299);
or U14034 (N_14034,N_13264,N_12150);
or U14035 (N_14035,N_12495,N_13284);
and U14036 (N_14036,N_13658,N_13965);
or U14037 (N_14037,N_12431,N_13311);
and U14038 (N_14038,N_12913,N_13974);
xor U14039 (N_14039,N_13550,N_12345);
nand U14040 (N_14040,N_13365,N_12992);
xnor U14041 (N_14041,N_13565,N_12838);
nand U14042 (N_14042,N_13862,N_12570);
and U14043 (N_14043,N_13096,N_13615);
nor U14044 (N_14044,N_13490,N_12977);
nand U14045 (N_14045,N_13796,N_13477);
xor U14046 (N_14046,N_12665,N_12388);
xor U14047 (N_14047,N_12354,N_12428);
or U14048 (N_14048,N_13023,N_13968);
and U14049 (N_14049,N_13702,N_13239);
or U14050 (N_14050,N_13911,N_13743);
or U14051 (N_14051,N_13075,N_12245);
nand U14052 (N_14052,N_12560,N_13788);
xor U14053 (N_14053,N_13526,N_13914);
or U14054 (N_14054,N_13186,N_13335);
nand U14055 (N_14055,N_12529,N_12933);
nand U14056 (N_14056,N_13492,N_12036);
nor U14057 (N_14057,N_13649,N_13026);
and U14058 (N_14058,N_13227,N_12836);
and U14059 (N_14059,N_13852,N_12286);
and U14060 (N_14060,N_12089,N_12585);
nand U14061 (N_14061,N_13394,N_12243);
or U14062 (N_14062,N_13736,N_13206);
and U14063 (N_14063,N_12408,N_13527);
nor U14064 (N_14064,N_13606,N_13875);
nand U14065 (N_14065,N_12643,N_13515);
and U14066 (N_14066,N_13580,N_12682);
nand U14067 (N_14067,N_13292,N_13928);
or U14068 (N_14068,N_12039,N_12334);
nor U14069 (N_14069,N_13558,N_13067);
nand U14070 (N_14070,N_13832,N_13287);
nand U14071 (N_14071,N_13626,N_12805);
nor U14072 (N_14072,N_12515,N_12256);
nand U14073 (N_14073,N_13694,N_13548);
nor U14074 (N_14074,N_13830,N_12956);
and U14075 (N_14075,N_12722,N_12831);
xor U14076 (N_14076,N_13433,N_13233);
nor U14077 (N_14077,N_13908,N_12974);
and U14078 (N_14078,N_12523,N_12787);
and U14079 (N_14079,N_13418,N_12466);
nand U14080 (N_14080,N_12075,N_12756);
nor U14081 (N_14081,N_12511,N_13586);
xor U14082 (N_14082,N_13715,N_12950);
nor U14083 (N_14083,N_13359,N_12220);
nand U14084 (N_14084,N_13346,N_13351);
and U14085 (N_14085,N_13913,N_12661);
xnor U14086 (N_14086,N_13814,N_12946);
and U14087 (N_14087,N_13556,N_12845);
xnor U14088 (N_14088,N_12074,N_12072);
and U14089 (N_14089,N_13552,N_12967);
and U14090 (N_14090,N_13881,N_13345);
and U14091 (N_14091,N_12798,N_12603);
xor U14092 (N_14092,N_13534,N_13740);
and U14093 (N_14093,N_13505,N_12729);
or U14094 (N_14094,N_12359,N_12197);
nor U14095 (N_14095,N_12060,N_12772);
xnor U14096 (N_14096,N_12500,N_13302);
xnor U14097 (N_14097,N_13555,N_13471);
nand U14098 (N_14098,N_13673,N_12569);
or U14099 (N_14099,N_12848,N_12090);
nor U14100 (N_14100,N_12049,N_12367);
nor U14101 (N_14101,N_12347,N_12274);
nand U14102 (N_14102,N_13757,N_13575);
and U14103 (N_14103,N_12909,N_13624);
nor U14104 (N_14104,N_13431,N_13289);
and U14105 (N_14105,N_12423,N_12216);
nor U14106 (N_14106,N_12281,N_13275);
and U14107 (N_14107,N_13245,N_12324);
nand U14108 (N_14108,N_13013,N_12658);
and U14109 (N_14109,N_12827,N_12490);
and U14110 (N_14110,N_12728,N_13945);
or U14111 (N_14111,N_12817,N_12673);
xor U14112 (N_14112,N_12011,N_12684);
xor U14113 (N_14113,N_13309,N_13818);
xor U14114 (N_14114,N_13135,N_12080);
nor U14115 (N_14115,N_13171,N_12409);
nand U14116 (N_14116,N_13978,N_13668);
nand U14117 (N_14117,N_12142,N_13268);
or U14118 (N_14118,N_13343,N_13189);
and U14119 (N_14119,N_12394,N_13425);
or U14120 (N_14120,N_12514,N_12140);
and U14121 (N_14121,N_12073,N_13544);
or U14122 (N_14122,N_13942,N_12877);
nor U14123 (N_14123,N_12137,N_13455);
nor U14124 (N_14124,N_13525,N_13600);
and U14125 (N_14125,N_12048,N_13432);
nor U14126 (N_14126,N_13799,N_12826);
and U14127 (N_14127,N_13277,N_13175);
or U14128 (N_14128,N_12126,N_12475);
xnor U14129 (N_14129,N_12768,N_12634);
xor U14130 (N_14130,N_13887,N_13733);
and U14131 (N_14131,N_12619,N_13041);
xor U14132 (N_14132,N_12723,N_12232);
nand U14133 (N_14133,N_13435,N_13701);
nand U14134 (N_14134,N_12066,N_13783);
and U14135 (N_14135,N_12835,N_13308);
or U14136 (N_14136,N_12578,N_13953);
nor U14137 (N_14137,N_12686,N_12970);
nand U14138 (N_14138,N_12943,N_12172);
nor U14139 (N_14139,N_12901,N_12596);
nand U14140 (N_14140,N_13250,N_13994);
nor U14141 (N_14141,N_13138,N_13174);
nor U14142 (N_14142,N_13159,N_13291);
or U14143 (N_14143,N_12714,N_12749);
nand U14144 (N_14144,N_13404,N_12564);
nor U14145 (N_14145,N_12815,N_12551);
nand U14146 (N_14146,N_12790,N_13062);
nand U14147 (N_14147,N_12154,N_12244);
xor U14148 (N_14148,N_12069,N_13720);
nor U14149 (N_14149,N_12356,N_12847);
and U14150 (N_14150,N_13108,N_12719);
xor U14151 (N_14151,N_12116,N_13927);
xor U14152 (N_14152,N_13734,N_13620);
nor U14153 (N_14153,N_13132,N_13926);
nand U14154 (N_14154,N_12857,N_12200);
and U14155 (N_14155,N_12591,N_12443);
and U14156 (N_14156,N_13350,N_12635);
nor U14157 (N_14157,N_12293,N_12944);
and U14158 (N_14158,N_12233,N_12513);
xnor U14159 (N_14159,N_12794,N_12807);
nand U14160 (N_14160,N_12770,N_12818);
xnor U14161 (N_14161,N_13936,N_12065);
xor U14162 (N_14162,N_12370,N_13050);
xnor U14163 (N_14163,N_13065,N_13194);
nand U14164 (N_14164,N_13693,N_13363);
nand U14165 (N_14165,N_13458,N_13969);
and U14166 (N_14166,N_12672,N_13161);
and U14167 (N_14167,N_13497,N_13155);
and U14168 (N_14168,N_12027,N_12867);
nand U14169 (N_14169,N_12023,N_12246);
nand U14170 (N_14170,N_12616,N_13508);
nand U14171 (N_14171,N_12181,N_12986);
xnor U14172 (N_14172,N_12812,N_12639);
nand U14173 (N_14173,N_12025,N_13637);
and U14174 (N_14174,N_13835,N_13376);
nor U14175 (N_14175,N_12823,N_12978);
or U14176 (N_14176,N_12516,N_13819);
nand U14177 (N_14177,N_13040,N_13670);
xnor U14178 (N_14178,N_13638,N_13681);
nand U14179 (N_14179,N_13697,N_12864);
and U14180 (N_14180,N_13741,N_13695);
and U14181 (N_14181,N_12067,N_13920);
nand U14182 (N_14182,N_12327,N_13551);
or U14183 (N_14183,N_12808,N_12429);
xnor U14184 (N_14184,N_12678,N_12020);
and U14185 (N_14185,N_12664,N_12572);
or U14186 (N_14186,N_13218,N_12064);
or U14187 (N_14187,N_13679,N_12078);
nand U14188 (N_14188,N_13398,N_12206);
nor U14189 (N_14189,N_12365,N_13313);
xor U14190 (N_14190,N_12786,N_13970);
nor U14191 (N_14191,N_13622,N_13721);
xor U14192 (N_14192,N_12600,N_13479);
nand U14193 (N_14193,N_12556,N_13669);
xor U14194 (N_14194,N_13775,N_13358);
nor U14195 (N_14195,N_12111,N_12712);
and U14196 (N_14196,N_13181,N_13434);
nor U14197 (N_14197,N_12637,N_12084);
and U14198 (N_14198,N_13102,N_12631);
xnor U14199 (N_14199,N_12526,N_13472);
nand U14200 (N_14200,N_12883,N_13342);
or U14201 (N_14201,N_12052,N_12758);
nand U14202 (N_14202,N_12254,N_13530);
nand U14203 (N_14203,N_13301,N_12653);
nor U14204 (N_14204,N_13440,N_12963);
and U14205 (N_14205,N_12353,N_13506);
or U14206 (N_14206,N_12364,N_13635);
nor U14207 (N_14207,N_12028,N_12437);
nand U14208 (N_14208,N_12467,N_12995);
nor U14209 (N_14209,N_12735,N_13267);
and U14210 (N_14210,N_12902,N_13707);
or U14211 (N_14211,N_12122,N_13977);
and U14212 (N_14212,N_12480,N_12830);
nor U14213 (N_14213,N_12498,N_13730);
or U14214 (N_14214,N_13991,N_12892);
and U14215 (N_14215,N_12479,N_12229);
or U14216 (N_14216,N_13823,N_12785);
nor U14217 (N_14217,N_13517,N_13086);
nand U14218 (N_14218,N_12333,N_13858);
xnor U14219 (N_14219,N_12789,N_12397);
nor U14220 (N_14220,N_13906,N_13957);
nand U14221 (N_14221,N_13598,N_13018);
nand U14222 (N_14222,N_13371,N_13400);
nor U14223 (N_14223,N_13469,N_13630);
and U14224 (N_14224,N_12488,N_13771);
and U14225 (N_14225,N_13032,N_13270);
nor U14226 (N_14226,N_12966,N_12985);
nand U14227 (N_14227,N_12783,N_12973);
nand U14228 (N_14228,N_13263,N_12932);
xnor U14229 (N_14229,N_13120,N_12934);
and U14230 (N_14230,N_13008,N_13068);
and U14231 (N_14231,N_13348,N_12435);
nor U14232 (N_14232,N_13223,N_12169);
or U14233 (N_14233,N_12898,N_13762);
nor U14234 (N_14234,N_12218,N_12453);
and U14235 (N_14235,N_12706,N_12125);
and U14236 (N_14236,N_12257,N_12760);
nor U14237 (N_14237,N_13100,N_13379);
nand U14238 (N_14238,N_13765,N_13905);
nor U14239 (N_14239,N_12800,N_12920);
xor U14240 (N_14240,N_12026,N_13979);
or U14241 (N_14241,N_12131,N_12338);
nand U14242 (N_14242,N_12699,N_12710);
and U14243 (N_14243,N_13072,N_12228);
nand U14244 (N_14244,N_13043,N_12589);
nor U14245 (N_14245,N_12108,N_12348);
xor U14246 (N_14246,N_13093,N_13930);
xor U14247 (N_14247,N_12965,N_13869);
and U14248 (N_14248,N_13468,N_12846);
or U14249 (N_14249,N_12313,N_12656);
and U14250 (N_14250,N_12262,N_12180);
nand U14251 (N_14251,N_13304,N_12510);
nand U14252 (N_14252,N_13004,N_12765);
and U14253 (N_14253,N_13048,N_12605);
xnor U14254 (N_14254,N_13639,N_13397);
xnor U14255 (N_14255,N_12024,N_13326);
xnor U14256 (N_14256,N_13893,N_12548);
xnor U14257 (N_14257,N_13522,N_12509);
nand U14258 (N_14258,N_12925,N_12700);
nand U14259 (N_14259,N_12235,N_13807);
or U14260 (N_14260,N_12693,N_12602);
xor U14261 (N_14261,N_13107,N_12102);
nor U14262 (N_14262,N_12717,N_13111);
xor U14263 (N_14263,N_13759,N_12378);
xnor U14264 (N_14264,N_13939,N_13449);
and U14265 (N_14265,N_12337,N_13029);
or U14266 (N_14266,N_13060,N_13320);
xor U14267 (N_14267,N_13648,N_13137);
nand U14268 (N_14268,N_13524,N_12414);
nand U14269 (N_14269,N_12696,N_12754);
xor U14270 (N_14270,N_13964,N_12019);
nand U14271 (N_14271,N_12307,N_13898);
nor U14272 (N_14272,N_13423,N_12814);
and U14273 (N_14273,N_13528,N_13752);
and U14274 (N_14274,N_12389,N_13420);
nor U14275 (N_14275,N_13878,N_13691);
xnor U14276 (N_14276,N_12780,N_13981);
nor U14277 (N_14277,N_12962,N_13871);
nand U14278 (N_14278,N_13021,N_13574);
xnor U14279 (N_14279,N_12954,N_12915);
xor U14280 (N_14280,N_13450,N_12788);
xnor U14281 (N_14281,N_13587,N_12162);
or U14282 (N_14282,N_12465,N_12834);
or U14283 (N_14283,N_12076,N_13012);
nor U14284 (N_14284,N_13564,N_13387);
nand U14285 (N_14285,N_12178,N_12566);
xnor U14286 (N_14286,N_13466,N_13801);
or U14287 (N_14287,N_12375,N_13375);
xnor U14288 (N_14288,N_13054,N_12816);
nor U14289 (N_14289,N_12177,N_13407);
and U14290 (N_14290,N_13602,N_13859);
nor U14291 (N_14291,N_12247,N_13607);
xnor U14292 (N_14292,N_12456,N_12042);
xnor U14293 (N_14293,N_13087,N_12911);
nand U14294 (N_14294,N_12419,N_12208);
xnor U14295 (N_14295,N_13772,N_13349);
nand U14296 (N_14296,N_12227,N_13485);
xor U14297 (N_14297,N_13610,N_12432);
xor U14298 (N_14298,N_12761,N_12340);
nand U14299 (N_14299,N_12879,N_13584);
xnor U14300 (N_14300,N_12179,N_12980);
nand U14301 (N_14301,N_13170,N_13570);
and U14302 (N_14302,N_12949,N_12007);
nor U14303 (N_14303,N_13993,N_12123);
or U14304 (N_14304,N_13849,N_12033);
and U14305 (N_14305,N_12399,N_12441);
nand U14306 (N_14306,N_13827,N_13665);
nand U14307 (N_14307,N_13051,N_13634);
xnor U14308 (N_14308,N_12046,N_12553);
or U14309 (N_14309,N_12527,N_13767);
nor U14310 (N_14310,N_13502,N_13361);
or U14311 (N_14311,N_13163,N_13180);
xor U14312 (N_14312,N_12797,N_12751);
xnor U14313 (N_14313,N_13019,N_12725);
nand U14314 (N_14314,N_12420,N_13674);
or U14315 (N_14315,N_12031,N_12576);
xor U14316 (N_14316,N_13971,N_13145);
and U14317 (N_14317,N_12802,N_12343);
nor U14318 (N_14318,N_13738,N_13999);
xor U14319 (N_14319,N_13549,N_12624);
and U14320 (N_14320,N_12905,N_13710);
nor U14321 (N_14321,N_13139,N_12595);
nor U14322 (N_14322,N_12483,N_12282);
nor U14323 (N_14323,N_12470,N_13184);
nor U14324 (N_14324,N_12310,N_13922);
and U14325 (N_14325,N_12391,N_13436);
and U14326 (N_14326,N_12899,N_13201);
nor U14327 (N_14327,N_12539,N_13136);
and U14328 (N_14328,N_12743,N_13333);
or U14329 (N_14329,N_12976,N_13243);
xnor U14330 (N_14330,N_12741,N_12190);
and U14331 (N_14331,N_13805,N_13446);
or U14332 (N_14332,N_12138,N_12234);
and U14333 (N_14333,N_13882,N_12828);
xnor U14334 (N_14334,N_12171,N_12574);
nand U14335 (N_14335,N_13536,N_12663);
or U14336 (N_14336,N_13148,N_13104);
or U14337 (N_14337,N_13412,N_12330);
xnor U14338 (N_14338,N_12371,N_13391);
nand U14339 (N_14339,N_13415,N_12189);
nand U14340 (N_14340,N_13076,N_13011);
xor U14341 (N_14341,N_12559,N_13937);
and U14342 (N_14342,N_13057,N_12862);
and U14343 (N_14343,N_12211,N_13990);
or U14344 (N_14344,N_13842,N_13402);
or U14345 (N_14345,N_13542,N_13405);
xor U14346 (N_14346,N_13178,N_13252);
nand U14347 (N_14347,N_13079,N_13232);
and U14348 (N_14348,N_12919,N_12960);
nand U14349 (N_14349,N_12844,N_13895);
and U14350 (N_14350,N_13056,N_13656);
nand U14351 (N_14351,N_12439,N_13885);
and U14352 (N_14352,N_13298,N_12690);
nand U14353 (N_14353,N_13103,N_13095);
and U14354 (N_14354,N_13495,N_13168);
or U14355 (N_14355,N_13151,N_13467);
nor U14356 (N_14356,N_12077,N_13246);
and U14357 (N_14357,N_12015,N_12926);
or U14358 (N_14358,N_13566,N_12999);
xor U14359 (N_14359,N_13010,N_13234);
and U14360 (N_14360,N_13633,N_13966);
and U14361 (N_14361,N_13897,N_12536);
nor U14362 (N_14362,N_12489,N_13909);
nand U14363 (N_14363,N_13677,N_12146);
nand U14364 (N_14364,N_12240,N_13323);
xor U14365 (N_14365,N_13078,N_12438);
or U14366 (N_14366,N_12452,N_12612);
and U14367 (N_14367,N_12604,N_13793);
or U14368 (N_14368,N_13535,N_12900);
and U14369 (N_14369,N_12914,N_12196);
and U14370 (N_14370,N_13664,N_13597);
nor U14371 (N_14371,N_13925,N_12198);
xnor U14372 (N_14372,N_12681,N_13657);
and U14373 (N_14373,N_13370,N_13384);
nand U14374 (N_14374,N_13187,N_13419);
xor U14375 (N_14375,N_13876,N_12744);
nand U14376 (N_14376,N_13112,N_12418);
nand U14377 (N_14377,N_12339,N_12504);
nand U14378 (N_14378,N_12223,N_13557);
xor U14379 (N_14379,N_12859,N_13442);
or U14380 (N_14380,N_13791,N_12941);
nor U14381 (N_14381,N_13153,N_13009);
or U14382 (N_14382,N_12331,N_12799);
or U14383 (N_14383,N_12878,N_13237);
nor U14384 (N_14384,N_13512,N_13873);
nand U14385 (N_14385,N_13372,N_12611);
nor U14386 (N_14386,N_12520,N_13997);
nand U14387 (N_14387,N_13452,N_13954);
nand U14388 (N_14388,N_12746,N_12547);
nor U14389 (N_14389,N_13778,N_12363);
nand U14390 (N_14390,N_13498,N_13623);
and U14391 (N_14391,N_13618,N_12732);
or U14392 (N_14392,N_12546,N_13478);
and U14393 (N_14393,N_13339,N_12091);
nand U14394 (N_14394,N_12022,N_12104);
nand U14395 (N_14395,N_12872,N_13133);
xnor U14396 (N_14396,N_13687,N_12182);
and U14397 (N_14397,N_12193,N_13840);
nand U14398 (N_14398,N_13728,N_13518);
or U14399 (N_14399,N_12170,N_13005);
and U14400 (N_14400,N_12156,N_12936);
and U14401 (N_14401,N_12477,N_12461);
nand U14402 (N_14402,N_12173,N_12352);
nor U14403 (N_14403,N_13373,N_13073);
and U14404 (N_14404,N_12929,N_12528);
and U14405 (N_14405,N_13509,N_12110);
nor U14406 (N_14406,N_12311,N_12044);
and U14407 (N_14407,N_12820,N_13049);
nor U14408 (N_14408,N_12618,N_12646);
nor U14409 (N_14409,N_13453,N_13763);
and U14410 (N_14410,N_12561,N_13430);
xor U14411 (N_14411,N_12998,N_12454);
or U14412 (N_14412,N_12669,N_13774);
and U14413 (N_14413,N_13935,N_12264);
and U14414 (N_14414,N_13683,N_12540);
nor U14415 (N_14415,N_13190,N_12448);
or U14416 (N_14416,N_13396,N_12627);
and U14417 (N_14417,N_13236,N_13255);
xor U14418 (N_14418,N_12373,N_12265);
or U14419 (N_14419,N_12521,N_13003);
xor U14420 (N_14420,N_12051,N_12697);
xnor U14421 (N_14421,N_13907,N_13228);
and U14422 (N_14422,N_13356,N_13114);
or U14423 (N_14423,N_12912,N_13027);
nand U14424 (N_14424,N_12395,N_13627);
and U14425 (N_14425,N_13000,N_12942);
nor U14426 (N_14426,N_12451,N_13883);
or U14427 (N_14427,N_13744,N_12811);
and U14428 (N_14428,N_13629,N_13824);
or U14429 (N_14429,N_13248,N_12004);
xnor U14430 (N_14430,N_12422,N_13105);
or U14431 (N_14431,N_12757,N_13924);
and U14432 (N_14432,N_12473,N_12647);
nor U14433 (N_14433,N_13797,N_13956);
and U14434 (N_14434,N_13675,N_13143);
xnor U14435 (N_14435,N_12632,N_13947);
xnor U14436 (N_14436,N_12779,N_13847);
and U14437 (N_14437,N_13521,N_13619);
or U14438 (N_14438,N_12279,N_12212);
xnor U14439 (N_14439,N_13428,N_13621);
or U14440 (N_14440,N_12318,N_12379);
xor U14441 (N_14441,N_13070,N_12813);
nand U14442 (N_14442,N_12215,N_13061);
xnor U14443 (N_14443,N_13089,N_13632);
nand U14444 (N_14444,N_12614,N_12219);
xnor U14445 (N_14445,N_12849,N_13754);
nand U14446 (N_14446,N_13154,N_13815);
xnor U14447 (N_14447,N_13781,N_13879);
nor U14448 (N_14448,N_12106,N_13663);
nor U14449 (N_14449,N_13147,N_13385);
or U14450 (N_14450,N_13886,N_13328);
nand U14451 (N_14451,N_12382,N_13739);
nor U14452 (N_14452,N_13982,N_13465);
and U14453 (N_14453,N_13015,N_13406);
xnor U14454 (N_14454,N_13213,N_12476);
and U14455 (N_14455,N_12225,N_13401);
xor U14456 (N_14456,N_12124,N_12620);
and U14457 (N_14457,N_13296,N_13306);
nor U14458 (N_14458,N_13812,N_12677);
nor U14459 (N_14459,N_13848,N_13667);
nand U14460 (N_14460,N_12917,N_13742);
xor U14461 (N_14461,N_12842,N_12869);
or U14462 (N_14462,N_13853,N_12598);
nor U14463 (N_14463,N_13902,N_12101);
or U14464 (N_14464,N_12119,N_12662);
nand U14465 (N_14465,N_12839,N_12298);
and U14466 (N_14466,N_13052,N_13192);
nand U14467 (N_14467,N_12541,N_12755);
or U14468 (N_14468,N_12103,N_13438);
nor U14469 (N_14469,N_12679,N_12384);
nor U14470 (N_14470,N_12916,N_12115);
xor U14471 (N_14471,N_13039,N_12550);
nor U14472 (N_14472,N_13366,N_12517);
nand U14473 (N_14473,N_12165,N_13210);
nor U14474 (N_14474,N_12532,N_12440);
and U14475 (N_14475,N_12209,N_12592);
xor U14476 (N_14476,N_13034,N_12594);
and U14477 (N_14477,N_13919,N_12093);
and U14478 (N_14478,N_13751,N_13045);
nor U14479 (N_14479,N_12342,N_12336);
and U14480 (N_14480,N_13803,N_12961);
nor U14481 (N_14481,N_12463,N_12638);
nor U14482 (N_14482,N_12775,N_12676);
or U14483 (N_14483,N_13682,N_12450);
and U14484 (N_14484,N_12716,N_12648);
and U14485 (N_14485,N_12698,N_12392);
or U14486 (N_14486,N_12300,N_12297);
nor U14487 (N_14487,N_13773,N_13631);
nand U14488 (N_14488,N_12733,N_12107);
and U14489 (N_14489,N_13688,N_13064);
and U14490 (N_14490,N_13386,N_12544);
nor U14491 (N_14491,N_12117,N_12577);
and U14492 (N_14492,N_12804,N_13447);
xnor U14493 (N_14493,N_12459,N_12401);
nand U14494 (N_14494,N_12701,N_13459);
nand U14495 (N_14495,N_12615,N_12058);
xor U14496 (N_14496,N_13377,N_13785);
nor U14497 (N_14497,N_13599,N_12579);
xor U14498 (N_14498,N_12175,N_13732);
and U14499 (N_14499,N_12573,N_12442);
xnor U14500 (N_14500,N_12341,N_13417);
xnor U14501 (N_14501,N_13834,N_12411);
xnor U14502 (N_14502,N_12922,N_12133);
nand U14503 (N_14503,N_12100,N_12485);
or U14504 (N_14504,N_13134,N_13307);
xor U14505 (N_14505,N_13424,N_13578);
nand U14506 (N_14506,N_12088,N_13963);
and U14507 (N_14507,N_13253,N_12155);
and U14508 (N_14508,N_13496,N_12613);
nand U14509 (N_14509,N_13124,N_12667);
nand U14510 (N_14510,N_12781,N_13725);
nand U14511 (N_14511,N_13338,N_12599);
nand U14512 (N_14512,N_12989,N_13880);
or U14513 (N_14513,N_12997,N_13241);
nand U14514 (N_14514,N_13934,N_13729);
or U14515 (N_14515,N_12259,N_13719);
or U14516 (N_14516,N_13059,N_12890);
nor U14517 (N_14517,N_12657,N_13197);
and U14518 (N_14518,N_13098,N_12085);
nor U14519 (N_14519,N_12132,N_12358);
xor U14520 (N_14520,N_12792,N_13900);
nor U14521 (N_14521,N_12904,N_12621);
or U14522 (N_14522,N_13272,N_12406);
xnor U14523 (N_14523,N_13949,N_13381);
nand U14524 (N_14524,N_12854,N_13101);
xor U14525 (N_14525,N_13884,N_12263);
or U14526 (N_14526,N_13461,N_12947);
xor U14527 (N_14527,N_12718,N_13212);
nand U14528 (N_14528,N_13160,N_12005);
xor U14529 (N_14529,N_12446,N_13860);
nor U14530 (N_14530,N_12763,N_13360);
nand U14531 (N_14531,N_13617,N_13951);
and U14532 (N_14532,N_13251,N_12272);
nand U14533 (N_14533,N_12567,N_12972);
and U14534 (N_14534,N_12875,N_13533);
nor U14535 (N_14535,N_13486,N_13156);
nor U14536 (N_14536,N_12689,N_13576);
or U14537 (N_14537,N_13144,N_13689);
nor U14538 (N_14538,N_13317,N_12054);
nor U14539 (N_14539,N_12778,N_13007);
nand U14540 (N_14540,N_13655,N_12708);
nor U14541 (N_14541,N_12994,N_13747);
or U14542 (N_14542,N_13297,N_12660);
or U14543 (N_14543,N_13053,N_13867);
and U14544 (N_14544,N_12032,N_12670);
nor U14545 (N_14545,N_12285,N_13146);
and U14546 (N_14546,N_13531,N_12893);
and U14547 (N_14547,N_12151,N_13699);
and U14548 (N_14548,N_13305,N_12305);
or U14549 (N_14549,N_12655,N_13917);
xnor U14550 (N_14550,N_13177,N_12161);
nand U14551 (N_14551,N_12468,N_13749);
nor U14552 (N_14552,N_12981,N_12201);
and U14553 (N_14553,N_13768,N_13014);
or U14554 (N_14554,N_12207,N_12897);
and U14555 (N_14555,N_13484,N_13608);
or U14556 (N_14556,N_13164,N_13713);
or U14557 (N_14557,N_13322,N_12711);
nand U14558 (N_14558,N_12871,N_12315);
xor U14559 (N_14559,N_12806,N_13271);
or U14560 (N_14560,N_12649,N_12887);
nor U14561 (N_14561,N_12505,N_12149);
nor U14562 (N_14562,N_12413,N_13193);
or U14563 (N_14563,N_12720,N_13454);
nor U14564 (N_14564,N_13659,N_13579);
xor U14565 (N_14565,N_13336,N_12043);
and U14566 (N_14566,N_13959,N_13929);
nand U14567 (N_14567,N_12764,N_13414);
xor U14568 (N_14568,N_12292,N_13393);
nor U14569 (N_14569,N_12948,N_13811);
or U14570 (N_14570,N_13779,N_13321);
nand U14571 (N_14571,N_13167,N_12127);
xor U14572 (N_14572,N_13047,N_13226);
and U14573 (N_14573,N_13962,N_12400);
and U14574 (N_14574,N_13382,N_12012);
xor U14575 (N_14575,N_13295,N_12852);
nand U14576 (N_14576,N_12056,N_12464);
nor U14577 (N_14577,N_13861,N_12222);
nand U14578 (N_14578,N_12837,N_13709);
xnor U14579 (N_14579,N_12704,N_13870);
nor U14580 (N_14580,N_13445,N_12555);
or U14581 (N_14581,N_13205,N_13987);
nor U14582 (N_14582,N_13033,N_12321);
nor U14583 (N_14583,N_13069,N_13955);
xnor U14584 (N_14584,N_12351,N_13547);
or U14585 (N_14585,N_13094,N_13782);
and U14586 (N_14586,N_13441,N_12885);
and U14587 (N_14587,N_12008,N_13127);
or U14588 (N_14588,N_13121,N_12059);
and U14589 (N_14589,N_12955,N_13353);
and U14590 (N_14590,N_13501,N_13614);
and U14591 (N_14591,N_12494,N_12147);
nor U14592 (N_14592,N_12194,N_13113);
nand U14593 (N_14593,N_13590,N_13158);
nor U14594 (N_14594,N_13750,N_13399);
or U14595 (N_14595,N_13383,N_13724);
xor U14596 (N_14596,N_12009,N_13642);
nand U14597 (N_14597,N_13242,N_13538);
and U14598 (N_14598,N_12554,N_13421);
nand U14599 (N_14599,N_13904,N_12583);
and U14600 (N_14600,N_13392,N_12128);
or U14601 (N_14601,N_13046,N_13532);
nor U14602 (N_14602,N_12276,N_13312);
and U14603 (N_14603,N_13474,N_13031);
and U14604 (N_14604,N_13211,N_13865);
nand U14605 (N_14605,N_12302,N_13507);
or U14606 (N_14606,N_13519,N_12114);
xor U14607 (N_14607,N_12773,N_12045);
nand U14608 (N_14608,N_12269,N_13464);
xor U14609 (N_14609,N_13706,N_12118);
xor U14610 (N_14610,N_12927,N_13554);
xor U14611 (N_14611,N_13462,N_13813);
xor U14612 (N_14612,N_12144,N_12289);
nand U14613 (N_14613,N_12882,N_13543);
xor U14614 (N_14614,N_13416,N_13916);
or U14615 (N_14615,N_12275,N_12081);
nor U14616 (N_14616,N_12957,N_12407);
or U14617 (N_14617,N_12810,N_12323);
xor U14618 (N_14618,N_12908,N_13931);
xor U14619 (N_14619,N_12425,N_13475);
and U14620 (N_14620,N_12303,N_12568);
and U14621 (N_14621,N_12668,N_12086);
or U14622 (N_14622,N_12562,N_12644);
nor U14623 (N_14623,N_12930,N_12843);
xor U14624 (N_14624,N_12478,N_13976);
nand U14625 (N_14625,N_13761,N_13992);
nor U14626 (N_14626,N_12750,N_13220);
and U14627 (N_14627,N_12447,N_13777);
nand U14628 (N_14628,N_13310,N_12237);
nor U14629 (N_14629,N_13357,N_12290);
or U14630 (N_14630,N_12841,N_13810);
or U14631 (N_14631,N_12436,N_13520);
nand U14632 (N_14632,N_13894,N_12164);
xor U14633 (N_14633,N_12287,N_13705);
nand U14634 (N_14634,N_13585,N_13081);
xor U14635 (N_14635,N_13808,N_13020);
and U14636 (N_14636,N_13244,N_12360);
and U14637 (N_14637,N_13690,N_13225);
xor U14638 (N_14638,N_13038,N_12691);
nor U14639 (N_14639,N_12833,N_13961);
and U14640 (N_14640,N_13082,N_12623);
and U14641 (N_14641,N_13787,N_12021);
or U14642 (N_14642,N_12876,N_12174);
and U14643 (N_14643,N_12694,N_13836);
or U14644 (N_14644,N_12214,N_12398);
nor U14645 (N_14645,N_12522,N_13367);
or U14646 (N_14646,N_12964,N_13006);
nand U14647 (N_14647,N_13755,N_12959);
and U14648 (N_14648,N_12923,N_13846);
nor U14649 (N_14649,N_12715,N_13247);
or U14650 (N_14650,N_12796,N_12747);
xnor U14651 (N_14651,N_12304,N_12990);
nand U14652 (N_14652,N_12312,N_12152);
xor U14653 (N_14653,N_12061,N_13983);
or U14654 (N_14654,N_13604,N_12168);
or U14655 (N_14655,N_12121,N_13214);
nor U14656 (N_14656,N_13195,N_13422);
or U14657 (N_14657,N_12380,N_13660);
xor U14658 (N_14658,N_13230,N_13503);
or U14659 (N_14659,N_12270,N_12226);
or U14660 (N_14660,N_12471,N_13126);
and U14661 (N_14661,N_13844,N_13457);
or U14662 (N_14662,N_13776,N_13354);
nand U14663 (N_14663,N_12112,N_13222);
and U14664 (N_14664,N_13410,N_13516);
or U14665 (N_14665,N_13989,N_13698);
or U14666 (N_14666,N_13426,N_13016);
or U14667 (N_14667,N_12737,N_13932);
and U14668 (N_14668,N_13571,N_12278);
nor U14669 (N_14669,N_12628,N_12727);
and U14670 (N_14670,N_12041,N_12350);
and U14671 (N_14671,N_13332,N_12782);
xor U14672 (N_14672,N_13973,N_12531);
xor U14673 (N_14673,N_12248,N_12491);
nand U14674 (N_14674,N_13269,N_13055);
nand U14675 (N_14675,N_13352,N_13745);
xor U14676 (N_14676,N_12460,N_13612);
xnor U14677 (N_14677,N_13409,N_12291);
nor U14678 (N_14678,N_13795,N_13240);
nor U14679 (N_14679,N_13165,N_13723);
or U14680 (N_14680,N_13259,N_13563);
nor U14681 (N_14681,N_12006,N_12549);
xnor U14682 (N_14682,N_12642,N_13504);
nor U14683 (N_14683,N_12266,N_13537);
and U14684 (N_14684,N_13002,N_13074);
nor U14685 (N_14685,N_12736,N_13480);
or U14686 (N_14686,N_13746,N_13123);
or U14687 (N_14687,N_12654,N_12745);
xor U14688 (N_14688,N_13611,N_13756);
nand U14689 (N_14689,N_13249,N_13510);
nand U14690 (N_14690,N_12167,N_12821);
or U14691 (N_14691,N_13001,N_12316);
and U14692 (N_14692,N_13910,N_12606);
xor U14693 (N_14693,N_13717,N_13331);
and U14694 (N_14694,N_12971,N_12707);
and U14695 (N_14695,N_13395,N_12376);
or U14696 (N_14696,N_13562,N_12575);
xor U14697 (N_14697,N_13603,N_12349);
or U14698 (N_14698,N_12249,N_13022);
nor U14699 (N_14699,N_13413,N_13802);
nor U14700 (N_14700,N_12134,N_12001);
nor U14701 (N_14701,N_13540,N_12410);
or U14702 (N_14702,N_13829,N_13573);
nand U14703 (N_14703,N_13283,N_13950);
and U14704 (N_14704,N_13588,N_13972);
nand U14705 (N_14705,N_12176,N_12224);
nand U14706 (N_14706,N_13661,N_12250);
xor U14707 (N_14707,N_12703,N_12709);
nor U14708 (N_14708,N_13216,N_13092);
or U14709 (N_14709,N_12771,N_13369);
nand U14710 (N_14710,N_13316,N_13899);
xnor U14711 (N_14711,N_13300,N_13493);
xnor U14712 (N_14712,N_12738,N_13903);
nor U14713 (N_14713,N_12850,N_12186);
nand U14714 (N_14714,N_12724,N_12185);
or U14715 (N_14715,N_13589,N_13857);
xnor U14716 (N_14716,N_12499,N_13559);
nor U14717 (N_14717,N_12597,N_12277);
nor U14718 (N_14718,N_13362,N_12784);
nor U14719 (N_14719,N_12481,N_13940);
nand U14720 (N_14720,N_13727,N_13198);
nor U14721 (N_14721,N_12545,N_13282);
and U14722 (N_14722,N_13714,N_13099);
or U14723 (N_14723,N_13948,N_12238);
xnor U14724 (N_14724,N_12769,N_12381);
and U14725 (N_14725,N_13601,N_12357);
xor U14726 (N_14726,N_12674,N_12099);
or U14727 (N_14727,N_13169,N_12740);
nand U14728 (N_14728,N_12387,N_12322);
or U14729 (N_14729,N_12748,N_12188);
and U14730 (N_14730,N_12063,N_13324);
and U14731 (N_14731,N_13279,N_12506);
xor U14732 (N_14732,N_12587,N_13806);
xnor U14733 (N_14733,N_12210,N_12630);
nand U14734 (N_14734,N_13877,N_13254);
nor U14735 (N_14735,N_12759,N_13591);
xor U14736 (N_14736,N_13686,N_12294);
or U14737 (N_14737,N_12969,N_12415);
or U14738 (N_14738,N_13314,N_12924);
xnor U14739 (N_14739,N_12486,N_13653);
nand U14740 (N_14740,N_12158,N_13337);
or U14741 (N_14741,N_13258,N_13613);
nand U14742 (N_14742,N_13200,N_12524);
xnor U14743 (N_14743,N_12306,N_13162);
and U14744 (N_14744,N_12991,N_12319);
and U14745 (N_14745,N_12038,N_12641);
nand U14746 (N_14746,N_13636,N_13188);
and U14747 (N_14747,N_13896,N_13794);
or U14748 (N_14748,N_13854,N_13605);
and U14749 (N_14749,N_13609,N_12332);
nor U14750 (N_14750,N_13511,N_12484);
nand U14751 (N_14751,N_13262,N_13488);
nand U14752 (N_14752,N_13278,N_13889);
xor U14753 (N_14753,N_12267,N_13647);
xor U14754 (N_14754,N_12884,N_13784);
xor U14755 (N_14755,N_13274,N_13592);
and U14756 (N_14756,N_12731,N_13645);
nand U14757 (N_14757,N_12405,N_12993);
nor U14758 (N_14758,N_13888,N_13822);
and U14759 (N_14759,N_12688,N_12910);
xor U14760 (N_14760,N_12296,N_12472);
nor U14761 (N_14761,N_12000,N_13915);
and U14762 (N_14762,N_13364,N_12958);
nor U14763 (N_14763,N_12940,N_12017);
xor U14764 (N_14764,N_12774,N_13790);
nand U14765 (N_14765,N_12687,N_13514);
and U14766 (N_14766,N_13838,N_12239);
or U14767 (N_14767,N_13960,N_13330);
or U14768 (N_14768,N_12087,N_13985);
nor U14769 (N_14769,N_12582,N_12894);
or U14770 (N_14770,N_12874,N_13831);
nand U14771 (N_14771,N_12258,N_12047);
xnor U14772 (N_14772,N_13260,N_12825);
nand U14773 (N_14773,N_13541,N_13988);
and U14774 (N_14774,N_13817,N_12863);
nand U14775 (N_14775,N_13851,N_13821);
and U14776 (N_14776,N_13281,N_13828);
and U14777 (N_14777,N_12866,N_13083);
xnor U14778 (N_14778,N_12096,N_12268);
xnor U14779 (N_14779,N_12903,N_13403);
nor U14780 (N_14780,N_12518,N_13341);
nand U14781 (N_14781,N_12721,N_12094);
nor U14782 (N_14782,N_13980,N_13770);
and U14783 (N_14783,N_13116,N_12801);
nand U14784 (N_14784,N_12230,N_12609);
xnor U14785 (N_14785,N_13553,N_12120);
or U14786 (N_14786,N_13294,N_12105);
or U14787 (N_14787,N_13892,N_12588);
nand U14788 (N_14788,N_12873,N_13118);
nand U14789 (N_14789,N_13117,N_12355);
nand U14790 (N_14790,N_12329,N_13700);
and U14791 (N_14791,N_12685,N_13952);
and U14792 (N_14792,N_12861,N_12284);
nand U14793 (N_14793,N_13037,N_13529);
and U14794 (N_14794,N_12068,N_13444);
nand U14795 (N_14795,N_12675,N_12622);
xnor U14796 (N_14796,N_12650,N_13077);
nand U14797 (N_14797,N_12493,N_13224);
and U14798 (N_14798,N_12434,N_12148);
xnor U14799 (N_14799,N_12931,N_12645);
and U14800 (N_14800,N_12029,N_12533);
nand U14801 (N_14801,N_13737,N_13943);
and U14802 (N_14802,N_12988,N_12362);
nor U14803 (N_14803,N_13666,N_13473);
xnor U14804 (N_14804,N_12542,N_12629);
xnor U14805 (N_14805,N_12881,N_13692);
xor U14806 (N_14806,N_12403,N_13800);
xnor U14807 (N_14807,N_12083,N_13091);
and U14808 (N_14808,N_12508,N_13685);
nand U14809 (N_14809,N_13716,N_13024);
and U14810 (N_14810,N_13106,N_13176);
or U14811 (N_14811,N_13115,N_12053);
or U14812 (N_14812,N_13712,N_12565);
nand U14813 (N_14813,N_12184,N_13640);
and U14814 (N_14814,N_12377,N_13643);
and U14815 (N_14815,N_13758,N_12636);
or U14816 (N_14816,N_12424,N_12683);
nand U14817 (N_14817,N_12203,N_13231);
nand U14818 (N_14818,N_13183,N_12617);
and U14819 (N_14819,N_12512,N_12143);
nand U14820 (N_14820,N_13439,N_12507);
and U14821 (N_14821,N_12626,N_13680);
or U14822 (N_14822,N_13769,N_12014);
and U14823 (N_14823,N_13837,N_13513);
nand U14824 (N_14824,N_13944,N_12593);
xnor U14825 (N_14825,N_13286,N_13798);
nor U14826 (N_14826,N_13229,N_13539);
and U14827 (N_14827,N_13489,N_12251);
and U14828 (N_14828,N_12141,N_13036);
xnor U14829 (N_14829,N_13764,N_13872);
nor U14830 (N_14830,N_12855,N_12659);
nand U14831 (N_14831,N_12308,N_13726);
or U14832 (N_14832,N_12695,N_12462);
nor U14833 (N_14833,N_12581,N_13140);
nand U14834 (N_14834,N_13080,N_12860);
nor U14835 (N_14835,N_13217,N_13650);
or U14836 (N_14836,N_13389,N_12195);
nor U14837 (N_14837,N_13545,N_13130);
or U14838 (N_14838,N_12153,N_13651);
or U14839 (N_14839,N_13596,N_12030);
nand U14840 (N_14840,N_12040,N_13933);
xor U14841 (N_14841,N_12938,N_12766);
xor U14842 (N_14842,N_13128,N_12776);
nor U14843 (N_14843,N_12320,N_13265);
nor U14844 (N_14844,N_13792,N_12803);
xnor U14845 (N_14845,N_13753,N_12543);
nand U14846 (N_14846,N_13678,N_12501);
and U14847 (N_14847,N_12928,N_12987);
nand U14848 (N_14848,N_13334,N_12010);
nor U14849 (N_14849,N_12433,N_13429);
or U14850 (N_14850,N_13122,N_12199);
nand U14851 (N_14851,N_12487,N_12537);
xnor U14852 (N_14852,N_12474,N_13561);
nor U14853 (N_14853,N_13207,N_13030);
nand U14854 (N_14854,N_13185,N_13157);
nand U14855 (N_14855,N_13221,N_12139);
or U14856 (N_14856,N_12557,N_12968);
xor U14857 (N_14857,N_13676,N_12145);
nor U14858 (N_14858,N_12444,N_13874);
and U14859 (N_14859,N_13833,N_12426);
or U14860 (N_14860,N_13975,N_12261);
nor U14861 (N_14861,N_13347,N_13644);
nand U14862 (N_14862,N_13119,N_13684);
xnor U14863 (N_14863,N_12002,N_12984);
nor U14864 (N_14864,N_12412,N_13662);
and U14865 (N_14865,N_13172,N_13938);
nand U14866 (N_14866,N_13129,N_13921);
and U14867 (N_14867,N_12309,N_13285);
or U14868 (N_14868,N_12607,N_12079);
nand U14869 (N_14869,N_13408,N_12982);
and U14870 (N_14870,N_13063,N_13652);
nor U14871 (N_14871,N_13315,N_12344);
nand U14872 (N_14872,N_12003,N_13748);
nand U14873 (N_14873,N_13238,N_12160);
and U14874 (N_14874,N_12326,N_12253);
or U14875 (N_14875,N_12283,N_12328);
nand U14876 (N_14876,N_12325,N_12260);
nand U14877 (N_14877,N_12651,N_13546);
xnor U14878 (N_14878,N_13084,N_12819);
nand U14879 (N_14879,N_12445,N_12390);
or U14880 (N_14880,N_12858,N_12082);
and U14881 (N_14881,N_12726,N_12136);
and U14882 (N_14882,N_13152,N_12895);
or U14883 (N_14883,N_13125,N_13173);
and U14884 (N_14884,N_12482,N_13378);
nand U14885 (N_14885,N_12889,N_13704);
or U14886 (N_14886,N_12610,N_12666);
or U14887 (N_14887,N_12288,N_12295);
and U14888 (N_14888,N_13941,N_12163);
xnor U14889 (N_14889,N_13890,N_13593);
or U14890 (N_14890,N_12374,N_12906);
nand U14891 (N_14891,N_13711,N_12166);
and U14892 (N_14892,N_13567,N_12832);
or U14893 (N_14893,N_13110,N_12213);
nor U14894 (N_14894,N_12095,N_13996);
xor U14895 (N_14895,N_12538,N_13582);
xor U14896 (N_14896,N_12455,N_12055);
xor U14897 (N_14897,N_13318,N_12034);
xor U14898 (N_14898,N_12018,N_13150);
or U14899 (N_14899,N_13280,N_12372);
and U14900 (N_14900,N_12204,N_13984);
nor U14901 (N_14901,N_13703,N_12937);
nor U14902 (N_14902,N_13864,N_12853);
xnor U14903 (N_14903,N_12205,N_12742);
nor U14904 (N_14904,N_13215,N_13202);
nand U14905 (N_14905,N_12502,N_13583);
nand U14906 (N_14906,N_12880,N_12951);
or U14907 (N_14907,N_12888,N_13487);
nand U14908 (N_14908,N_12590,N_12886);
or U14909 (N_14909,N_13625,N_13303);
or U14910 (N_14910,N_13196,N_13998);
nor U14911 (N_14911,N_12671,N_13261);
or U14912 (N_14912,N_12368,N_13995);
or U14913 (N_14913,N_13918,N_13843);
nor U14914 (N_14914,N_12335,N_13946);
or U14915 (N_14915,N_12393,N_12525);
or U14916 (N_14916,N_12935,N_13491);
and U14917 (N_14917,N_13325,N_13845);
nor U14918 (N_14918,N_13780,N_13986);
and U14919 (N_14919,N_12680,N_12713);
nor U14920 (N_14920,N_12856,N_13569);
or U14921 (N_14921,N_13646,N_12252);
nand U14922 (N_14922,N_13581,N_12945);
nand U14923 (N_14923,N_13482,N_12563);
nor U14924 (N_14924,N_12404,N_12273);
and U14925 (N_14925,N_12192,N_12016);
nand U14926 (N_14926,N_12497,N_12753);
xor U14927 (N_14927,N_12202,N_13299);
or U14928 (N_14928,N_12829,N_12777);
nor U14929 (N_14929,N_12221,N_13149);
xnor U14930 (N_14930,N_13290,N_13568);
or U14931 (N_14931,N_12217,N_13448);
or U14932 (N_14932,N_13257,N_12386);
xnor U14933 (N_14933,N_12752,N_13866);
or U14934 (N_14934,N_12402,N_12952);
nor U14935 (N_14935,N_12062,N_12346);
and U14936 (N_14936,N_13109,N_12097);
xnor U14937 (N_14937,N_12191,N_13967);
or U14938 (N_14938,N_12552,N_12918);
nand U14939 (N_14939,N_13766,N_13912);
or U14940 (N_14940,N_13735,N_12366);
nor U14941 (N_14941,N_13235,N_13380);
nor U14942 (N_14942,N_13839,N_12035);
nand U14943 (N_14943,N_12558,N_13319);
nor U14944 (N_14944,N_12601,N_13850);
xnor U14945 (N_14945,N_13722,N_12396);
nand U14946 (N_14946,N_12692,N_13809);
nand U14947 (N_14947,N_13028,N_13856);
nor U14948 (N_14948,N_13293,N_12231);
nand U14949 (N_14949,N_13789,N_13483);
and U14950 (N_14950,N_13025,N_13266);
xor U14951 (N_14951,N_12385,N_12953);
and U14952 (N_14952,N_12183,N_13411);
nor U14953 (N_14953,N_12496,N_13460);
xor U14954 (N_14954,N_13256,N_12767);
or U14955 (N_14955,N_12417,N_12157);
nand U14956 (N_14956,N_12361,N_13451);
xnor U14957 (N_14957,N_12050,N_12762);
nand U14958 (N_14958,N_13595,N_12071);
nor U14959 (N_14959,N_12608,N_12109);
nand U14960 (N_14960,N_13958,N_12891);
and U14961 (N_14961,N_13179,N_12865);
or U14962 (N_14962,N_13696,N_12469);
nand U14963 (N_14963,N_13340,N_13374);
nand U14964 (N_14964,N_13088,N_12640);
nand U14965 (N_14965,N_12492,N_13141);
nor U14966 (N_14966,N_12868,N_12822);
nor U14967 (N_14967,N_12241,N_13731);
nor U14968 (N_14968,N_13820,N_13035);
or U14969 (N_14969,N_13203,N_13901);
nand U14970 (N_14970,N_12534,N_13523);
xnor U14971 (N_14971,N_12130,N_13071);
nor U14972 (N_14972,N_12791,N_12255);
nand U14973 (N_14973,N_12633,N_13816);
and U14974 (N_14974,N_12092,N_13166);
nand U14975 (N_14975,N_13654,N_12242);
and U14976 (N_14976,N_13672,N_12571);
xor U14977 (N_14977,N_13760,N_13090);
and U14978 (N_14978,N_13671,N_13804);
xnor U14979 (N_14979,N_13204,N_13708);
nor U14980 (N_14980,N_12730,N_13494);
nand U14981 (N_14981,N_12795,N_12383);
or U14982 (N_14982,N_12129,N_13131);
nor U14983 (N_14983,N_13616,N_12625);
nor U14984 (N_14984,N_12921,N_13208);
and U14985 (N_14985,N_13329,N_12317);
or U14986 (N_14986,N_13390,N_12739);
and U14987 (N_14987,N_13058,N_13042);
or U14988 (N_14988,N_12652,N_12939);
or U14989 (N_14989,N_13855,N_12421);
xor U14990 (N_14990,N_12430,N_13427);
nor U14991 (N_14991,N_13209,N_12301);
nor U14992 (N_14992,N_12896,N_13500);
or U14993 (N_14993,N_12824,N_12057);
nand U14994 (N_14994,N_13344,N_12586);
or U14995 (N_14995,N_12535,N_12734);
xnor U14996 (N_14996,N_13368,N_12702);
or U14997 (N_14997,N_13456,N_13841);
xor U14998 (N_14998,N_12236,N_13628);
nor U14999 (N_14999,N_12705,N_13826);
and U15000 (N_15000,N_12344,N_12131);
xor U15001 (N_15001,N_12950,N_12521);
nand U15002 (N_15002,N_12602,N_13659);
nand U15003 (N_15003,N_12550,N_13765);
and U15004 (N_15004,N_12903,N_12796);
and U15005 (N_15005,N_12645,N_13302);
or U15006 (N_15006,N_12714,N_13086);
nor U15007 (N_15007,N_13191,N_13925);
or U15008 (N_15008,N_12363,N_12554);
xnor U15009 (N_15009,N_13427,N_12365);
and U15010 (N_15010,N_12440,N_13168);
nor U15011 (N_15011,N_12740,N_12210);
nand U15012 (N_15012,N_12078,N_12758);
xnor U15013 (N_15013,N_13412,N_13044);
nor U15014 (N_15014,N_13775,N_13132);
or U15015 (N_15015,N_12856,N_12435);
nor U15016 (N_15016,N_13489,N_13570);
or U15017 (N_15017,N_12702,N_12694);
or U15018 (N_15018,N_12573,N_12579);
xnor U15019 (N_15019,N_13777,N_13891);
nand U15020 (N_15020,N_13620,N_12422);
nand U15021 (N_15021,N_13431,N_13875);
and U15022 (N_15022,N_13126,N_13950);
xnor U15023 (N_15023,N_12856,N_12923);
and U15024 (N_15024,N_13966,N_13112);
and U15025 (N_15025,N_12559,N_13479);
xor U15026 (N_15026,N_12823,N_12549);
xor U15027 (N_15027,N_13204,N_12700);
and U15028 (N_15028,N_12695,N_13066);
and U15029 (N_15029,N_12201,N_13044);
nand U15030 (N_15030,N_13148,N_12197);
xnor U15031 (N_15031,N_13104,N_12622);
or U15032 (N_15032,N_12117,N_13589);
or U15033 (N_15033,N_13325,N_12314);
nand U15034 (N_15034,N_12289,N_13256);
nor U15035 (N_15035,N_13248,N_13183);
xor U15036 (N_15036,N_12134,N_12290);
and U15037 (N_15037,N_13741,N_13686);
and U15038 (N_15038,N_12502,N_12344);
and U15039 (N_15039,N_13251,N_13925);
xnor U15040 (N_15040,N_13865,N_13079);
nand U15041 (N_15041,N_13063,N_12061);
or U15042 (N_15042,N_12799,N_12657);
nand U15043 (N_15043,N_13201,N_13863);
or U15044 (N_15044,N_12445,N_13510);
xnor U15045 (N_15045,N_13984,N_12167);
and U15046 (N_15046,N_13223,N_12321);
nand U15047 (N_15047,N_13443,N_12122);
xor U15048 (N_15048,N_13088,N_12101);
nor U15049 (N_15049,N_12495,N_13313);
xor U15050 (N_15050,N_13811,N_12196);
nor U15051 (N_15051,N_13351,N_12297);
nor U15052 (N_15052,N_12403,N_12771);
xor U15053 (N_15053,N_13855,N_12246);
nor U15054 (N_15054,N_13336,N_13344);
nor U15055 (N_15055,N_12154,N_12015);
nor U15056 (N_15056,N_13615,N_13633);
nand U15057 (N_15057,N_13161,N_12130);
xnor U15058 (N_15058,N_12785,N_12900);
nor U15059 (N_15059,N_12636,N_13555);
or U15060 (N_15060,N_12448,N_13399);
and U15061 (N_15061,N_12723,N_12427);
and U15062 (N_15062,N_12432,N_12018);
nand U15063 (N_15063,N_12327,N_12472);
xor U15064 (N_15064,N_13986,N_12401);
and U15065 (N_15065,N_13934,N_13407);
nand U15066 (N_15066,N_13775,N_12136);
nor U15067 (N_15067,N_13449,N_12235);
xor U15068 (N_15068,N_13417,N_12676);
nand U15069 (N_15069,N_13952,N_12260);
nor U15070 (N_15070,N_13526,N_13489);
and U15071 (N_15071,N_12977,N_13647);
xor U15072 (N_15072,N_12799,N_12604);
nand U15073 (N_15073,N_13889,N_13985);
nand U15074 (N_15074,N_13650,N_13987);
nand U15075 (N_15075,N_12411,N_12216);
or U15076 (N_15076,N_12608,N_13110);
or U15077 (N_15077,N_13659,N_12773);
nand U15078 (N_15078,N_12564,N_12640);
and U15079 (N_15079,N_13684,N_13845);
xor U15080 (N_15080,N_12949,N_13764);
nor U15081 (N_15081,N_13288,N_12413);
nand U15082 (N_15082,N_12260,N_12661);
xor U15083 (N_15083,N_13771,N_13003);
or U15084 (N_15084,N_13032,N_12795);
xor U15085 (N_15085,N_13852,N_12195);
or U15086 (N_15086,N_13027,N_12197);
nand U15087 (N_15087,N_13193,N_13145);
xnor U15088 (N_15088,N_12576,N_12076);
xor U15089 (N_15089,N_13152,N_13917);
or U15090 (N_15090,N_13528,N_12517);
nor U15091 (N_15091,N_13966,N_13427);
nor U15092 (N_15092,N_13013,N_13667);
xor U15093 (N_15093,N_13545,N_12850);
xor U15094 (N_15094,N_13247,N_13354);
and U15095 (N_15095,N_13229,N_12558);
or U15096 (N_15096,N_13175,N_13090);
nand U15097 (N_15097,N_12431,N_13690);
and U15098 (N_15098,N_13987,N_13612);
or U15099 (N_15099,N_13392,N_13286);
nand U15100 (N_15100,N_12491,N_12676);
nand U15101 (N_15101,N_12146,N_13285);
or U15102 (N_15102,N_13993,N_12325);
nand U15103 (N_15103,N_12799,N_13320);
nand U15104 (N_15104,N_12867,N_12291);
nand U15105 (N_15105,N_13802,N_13061);
or U15106 (N_15106,N_12641,N_12834);
or U15107 (N_15107,N_13866,N_13781);
or U15108 (N_15108,N_13742,N_13741);
and U15109 (N_15109,N_13784,N_13052);
nor U15110 (N_15110,N_12515,N_13380);
and U15111 (N_15111,N_12839,N_13793);
and U15112 (N_15112,N_13969,N_13530);
nor U15113 (N_15113,N_13295,N_12096);
and U15114 (N_15114,N_13359,N_12720);
or U15115 (N_15115,N_13418,N_13604);
or U15116 (N_15116,N_13731,N_12619);
xnor U15117 (N_15117,N_13720,N_12161);
nand U15118 (N_15118,N_12294,N_12981);
nor U15119 (N_15119,N_12717,N_12952);
nand U15120 (N_15120,N_12391,N_12320);
nor U15121 (N_15121,N_13529,N_12741);
nand U15122 (N_15122,N_12228,N_12127);
and U15123 (N_15123,N_12134,N_13585);
nor U15124 (N_15124,N_12442,N_13547);
or U15125 (N_15125,N_12033,N_12107);
nand U15126 (N_15126,N_13897,N_13128);
or U15127 (N_15127,N_13012,N_13061);
or U15128 (N_15128,N_13935,N_13856);
or U15129 (N_15129,N_12234,N_12772);
or U15130 (N_15130,N_12820,N_13032);
nand U15131 (N_15131,N_12687,N_13074);
and U15132 (N_15132,N_12443,N_13662);
nor U15133 (N_15133,N_12778,N_13353);
xnor U15134 (N_15134,N_12515,N_12929);
and U15135 (N_15135,N_13224,N_12160);
and U15136 (N_15136,N_12081,N_12399);
nor U15137 (N_15137,N_12632,N_12178);
and U15138 (N_15138,N_12528,N_12690);
or U15139 (N_15139,N_12756,N_13352);
nand U15140 (N_15140,N_12827,N_13432);
or U15141 (N_15141,N_12777,N_13207);
and U15142 (N_15142,N_13121,N_12600);
and U15143 (N_15143,N_13977,N_12178);
or U15144 (N_15144,N_12970,N_13024);
or U15145 (N_15145,N_12140,N_13679);
xnor U15146 (N_15146,N_13065,N_13062);
and U15147 (N_15147,N_12187,N_13793);
and U15148 (N_15148,N_12212,N_13415);
nand U15149 (N_15149,N_13051,N_12095);
or U15150 (N_15150,N_12231,N_12852);
xor U15151 (N_15151,N_13953,N_13188);
and U15152 (N_15152,N_12796,N_12113);
and U15153 (N_15153,N_13344,N_13385);
nand U15154 (N_15154,N_13508,N_13790);
or U15155 (N_15155,N_13305,N_12979);
nor U15156 (N_15156,N_13799,N_12233);
nor U15157 (N_15157,N_12743,N_12286);
nor U15158 (N_15158,N_12118,N_12157);
nor U15159 (N_15159,N_12870,N_12592);
xor U15160 (N_15160,N_13228,N_12452);
or U15161 (N_15161,N_13162,N_13004);
nor U15162 (N_15162,N_13281,N_12507);
nand U15163 (N_15163,N_12352,N_13849);
and U15164 (N_15164,N_13531,N_13330);
and U15165 (N_15165,N_13844,N_12222);
or U15166 (N_15166,N_12382,N_12094);
nand U15167 (N_15167,N_13326,N_12670);
nor U15168 (N_15168,N_13805,N_12063);
nor U15169 (N_15169,N_12228,N_13147);
xor U15170 (N_15170,N_12203,N_13668);
nor U15171 (N_15171,N_12794,N_12229);
xnor U15172 (N_15172,N_13034,N_13696);
and U15173 (N_15173,N_12544,N_13811);
nand U15174 (N_15174,N_13503,N_13039);
xor U15175 (N_15175,N_12217,N_12560);
xnor U15176 (N_15176,N_12771,N_12564);
nand U15177 (N_15177,N_13193,N_13956);
nor U15178 (N_15178,N_12593,N_13861);
or U15179 (N_15179,N_13814,N_12456);
and U15180 (N_15180,N_12638,N_13744);
nor U15181 (N_15181,N_13937,N_12744);
and U15182 (N_15182,N_12900,N_13081);
or U15183 (N_15183,N_13305,N_12937);
nand U15184 (N_15184,N_13879,N_13023);
xor U15185 (N_15185,N_13330,N_13881);
xnor U15186 (N_15186,N_13874,N_13687);
or U15187 (N_15187,N_12563,N_13330);
and U15188 (N_15188,N_12772,N_12351);
and U15189 (N_15189,N_13804,N_13513);
nor U15190 (N_15190,N_12515,N_12381);
nand U15191 (N_15191,N_13570,N_13781);
xor U15192 (N_15192,N_13802,N_12897);
nor U15193 (N_15193,N_12765,N_13500);
nor U15194 (N_15194,N_13905,N_12031);
xor U15195 (N_15195,N_12095,N_12823);
or U15196 (N_15196,N_13506,N_12063);
nor U15197 (N_15197,N_13334,N_13719);
nor U15198 (N_15198,N_12459,N_12247);
nand U15199 (N_15199,N_12875,N_13995);
xor U15200 (N_15200,N_12140,N_13840);
or U15201 (N_15201,N_12169,N_12736);
xnor U15202 (N_15202,N_12308,N_13094);
or U15203 (N_15203,N_13656,N_12886);
nor U15204 (N_15204,N_13372,N_12543);
xnor U15205 (N_15205,N_12039,N_13271);
xor U15206 (N_15206,N_13708,N_12069);
nor U15207 (N_15207,N_13452,N_12382);
and U15208 (N_15208,N_12090,N_12539);
and U15209 (N_15209,N_12244,N_12141);
nand U15210 (N_15210,N_13316,N_12590);
xnor U15211 (N_15211,N_13640,N_12567);
and U15212 (N_15212,N_13594,N_13192);
nor U15213 (N_15213,N_12246,N_12966);
nor U15214 (N_15214,N_12280,N_13767);
nor U15215 (N_15215,N_12645,N_12563);
xor U15216 (N_15216,N_13007,N_13113);
nor U15217 (N_15217,N_13629,N_12119);
nand U15218 (N_15218,N_12218,N_12380);
and U15219 (N_15219,N_13137,N_13385);
xnor U15220 (N_15220,N_13349,N_12057);
and U15221 (N_15221,N_12889,N_13320);
nor U15222 (N_15222,N_12517,N_13989);
nand U15223 (N_15223,N_13021,N_13675);
or U15224 (N_15224,N_13904,N_13405);
and U15225 (N_15225,N_12026,N_13263);
nand U15226 (N_15226,N_12533,N_12316);
and U15227 (N_15227,N_13138,N_12581);
or U15228 (N_15228,N_12138,N_12001);
xor U15229 (N_15229,N_12715,N_12687);
nor U15230 (N_15230,N_12829,N_12946);
xor U15231 (N_15231,N_13310,N_13402);
nor U15232 (N_15232,N_12523,N_13909);
nor U15233 (N_15233,N_12448,N_12107);
or U15234 (N_15234,N_12312,N_13127);
or U15235 (N_15235,N_13443,N_13918);
nor U15236 (N_15236,N_12289,N_12688);
or U15237 (N_15237,N_13798,N_13919);
nand U15238 (N_15238,N_13908,N_12548);
or U15239 (N_15239,N_12661,N_12730);
xnor U15240 (N_15240,N_12884,N_12422);
and U15241 (N_15241,N_12878,N_12949);
nand U15242 (N_15242,N_12664,N_13741);
xnor U15243 (N_15243,N_13585,N_12623);
or U15244 (N_15244,N_12789,N_13302);
nand U15245 (N_15245,N_12674,N_13308);
nand U15246 (N_15246,N_12976,N_13559);
nand U15247 (N_15247,N_12300,N_12047);
and U15248 (N_15248,N_12421,N_13555);
or U15249 (N_15249,N_13742,N_13818);
nor U15250 (N_15250,N_13726,N_13085);
nor U15251 (N_15251,N_13145,N_12078);
xnor U15252 (N_15252,N_12354,N_12595);
nor U15253 (N_15253,N_12825,N_13426);
or U15254 (N_15254,N_13160,N_13832);
xor U15255 (N_15255,N_13023,N_12704);
nor U15256 (N_15256,N_12109,N_13606);
and U15257 (N_15257,N_13532,N_13084);
xnor U15258 (N_15258,N_12928,N_12657);
xnor U15259 (N_15259,N_12299,N_13835);
xnor U15260 (N_15260,N_12136,N_12922);
or U15261 (N_15261,N_12879,N_13786);
or U15262 (N_15262,N_13196,N_13100);
xor U15263 (N_15263,N_12998,N_12602);
nand U15264 (N_15264,N_13156,N_13514);
and U15265 (N_15265,N_12793,N_12289);
and U15266 (N_15266,N_13106,N_13687);
and U15267 (N_15267,N_13028,N_12931);
xor U15268 (N_15268,N_13195,N_12508);
nor U15269 (N_15269,N_13040,N_12040);
nand U15270 (N_15270,N_13650,N_13854);
nor U15271 (N_15271,N_12229,N_12207);
nand U15272 (N_15272,N_12353,N_12632);
nor U15273 (N_15273,N_12534,N_13018);
xor U15274 (N_15274,N_13454,N_12340);
nand U15275 (N_15275,N_12278,N_13952);
xor U15276 (N_15276,N_12901,N_13924);
or U15277 (N_15277,N_13789,N_12590);
nand U15278 (N_15278,N_12409,N_13366);
or U15279 (N_15279,N_13969,N_12034);
nor U15280 (N_15280,N_13883,N_13014);
nor U15281 (N_15281,N_13249,N_12643);
xnor U15282 (N_15282,N_12478,N_12023);
nand U15283 (N_15283,N_13492,N_13728);
nand U15284 (N_15284,N_13904,N_13518);
nand U15285 (N_15285,N_13067,N_12531);
or U15286 (N_15286,N_13776,N_13068);
or U15287 (N_15287,N_13826,N_12999);
nor U15288 (N_15288,N_12232,N_12722);
nor U15289 (N_15289,N_12395,N_12236);
nor U15290 (N_15290,N_13208,N_12454);
or U15291 (N_15291,N_12631,N_13847);
or U15292 (N_15292,N_13276,N_13649);
and U15293 (N_15293,N_13190,N_13766);
nor U15294 (N_15294,N_13278,N_12071);
or U15295 (N_15295,N_12138,N_12668);
nor U15296 (N_15296,N_13298,N_12884);
xor U15297 (N_15297,N_12933,N_12429);
nand U15298 (N_15298,N_12664,N_13538);
nand U15299 (N_15299,N_13365,N_12683);
and U15300 (N_15300,N_12179,N_13915);
xnor U15301 (N_15301,N_12053,N_12887);
xor U15302 (N_15302,N_12548,N_13808);
nand U15303 (N_15303,N_12087,N_13234);
nand U15304 (N_15304,N_13446,N_12933);
and U15305 (N_15305,N_12313,N_12282);
nor U15306 (N_15306,N_13288,N_12112);
xnor U15307 (N_15307,N_12468,N_12384);
xnor U15308 (N_15308,N_12388,N_13445);
nor U15309 (N_15309,N_13009,N_12453);
nor U15310 (N_15310,N_12321,N_13103);
nor U15311 (N_15311,N_13830,N_13652);
xnor U15312 (N_15312,N_12688,N_12057);
and U15313 (N_15313,N_12601,N_12717);
nand U15314 (N_15314,N_13063,N_12877);
and U15315 (N_15315,N_13376,N_12961);
nor U15316 (N_15316,N_13415,N_12171);
or U15317 (N_15317,N_12121,N_12005);
xnor U15318 (N_15318,N_13609,N_12569);
xnor U15319 (N_15319,N_12152,N_12804);
nor U15320 (N_15320,N_13837,N_12729);
nor U15321 (N_15321,N_13337,N_12682);
nand U15322 (N_15322,N_12812,N_13410);
and U15323 (N_15323,N_13075,N_12315);
or U15324 (N_15324,N_12884,N_12289);
or U15325 (N_15325,N_12103,N_13900);
or U15326 (N_15326,N_12289,N_13816);
nand U15327 (N_15327,N_13353,N_13379);
or U15328 (N_15328,N_12467,N_12183);
or U15329 (N_15329,N_13685,N_13338);
and U15330 (N_15330,N_13135,N_13455);
nand U15331 (N_15331,N_13255,N_12806);
nor U15332 (N_15332,N_13465,N_13166);
or U15333 (N_15333,N_13195,N_12793);
or U15334 (N_15334,N_12476,N_12791);
nand U15335 (N_15335,N_13756,N_12371);
xor U15336 (N_15336,N_12433,N_12107);
nor U15337 (N_15337,N_12235,N_12196);
nor U15338 (N_15338,N_12417,N_13370);
or U15339 (N_15339,N_13249,N_12595);
nor U15340 (N_15340,N_12257,N_13649);
or U15341 (N_15341,N_12386,N_12720);
and U15342 (N_15342,N_13275,N_13235);
or U15343 (N_15343,N_12566,N_12016);
xnor U15344 (N_15344,N_12936,N_12593);
xnor U15345 (N_15345,N_13939,N_12156);
or U15346 (N_15346,N_13217,N_13196);
and U15347 (N_15347,N_12524,N_12469);
nor U15348 (N_15348,N_12401,N_12076);
and U15349 (N_15349,N_13854,N_12005);
nor U15350 (N_15350,N_12713,N_12402);
or U15351 (N_15351,N_13320,N_12544);
nor U15352 (N_15352,N_12736,N_12267);
or U15353 (N_15353,N_12983,N_13139);
nand U15354 (N_15354,N_13619,N_12478);
and U15355 (N_15355,N_12013,N_12253);
or U15356 (N_15356,N_12127,N_12545);
nand U15357 (N_15357,N_12291,N_12553);
nand U15358 (N_15358,N_13764,N_12869);
or U15359 (N_15359,N_13550,N_12678);
nand U15360 (N_15360,N_13755,N_12067);
nand U15361 (N_15361,N_12766,N_12826);
or U15362 (N_15362,N_12828,N_12584);
or U15363 (N_15363,N_13623,N_12506);
nor U15364 (N_15364,N_13813,N_13359);
and U15365 (N_15365,N_13201,N_12980);
nor U15366 (N_15366,N_12445,N_12214);
or U15367 (N_15367,N_12933,N_13282);
or U15368 (N_15368,N_13927,N_13071);
xnor U15369 (N_15369,N_13474,N_13052);
and U15370 (N_15370,N_13384,N_12177);
and U15371 (N_15371,N_12094,N_13934);
and U15372 (N_15372,N_12527,N_13828);
or U15373 (N_15373,N_13882,N_13569);
nand U15374 (N_15374,N_12703,N_12415);
xor U15375 (N_15375,N_12433,N_13491);
and U15376 (N_15376,N_12754,N_12847);
and U15377 (N_15377,N_12173,N_13904);
nand U15378 (N_15378,N_12585,N_13452);
xor U15379 (N_15379,N_13202,N_12466);
nor U15380 (N_15380,N_13744,N_12276);
nor U15381 (N_15381,N_13566,N_12950);
xor U15382 (N_15382,N_12950,N_12270);
nand U15383 (N_15383,N_12068,N_12605);
or U15384 (N_15384,N_12732,N_12003);
or U15385 (N_15385,N_13978,N_12597);
xnor U15386 (N_15386,N_12613,N_13266);
or U15387 (N_15387,N_12822,N_13926);
and U15388 (N_15388,N_12117,N_12009);
nand U15389 (N_15389,N_12110,N_12849);
xnor U15390 (N_15390,N_12022,N_12569);
or U15391 (N_15391,N_13930,N_13084);
xor U15392 (N_15392,N_13780,N_13654);
nand U15393 (N_15393,N_13743,N_12587);
nand U15394 (N_15394,N_12085,N_12378);
and U15395 (N_15395,N_13254,N_13361);
nand U15396 (N_15396,N_12523,N_12065);
or U15397 (N_15397,N_13951,N_13993);
or U15398 (N_15398,N_13252,N_13798);
and U15399 (N_15399,N_12460,N_12754);
nand U15400 (N_15400,N_13577,N_13845);
nand U15401 (N_15401,N_13542,N_12554);
or U15402 (N_15402,N_13850,N_13503);
and U15403 (N_15403,N_12698,N_13773);
or U15404 (N_15404,N_13135,N_12720);
nor U15405 (N_15405,N_13329,N_13727);
and U15406 (N_15406,N_12964,N_13455);
nor U15407 (N_15407,N_12530,N_12221);
nor U15408 (N_15408,N_12508,N_12565);
nand U15409 (N_15409,N_12257,N_13640);
or U15410 (N_15410,N_12564,N_12509);
and U15411 (N_15411,N_12371,N_13306);
and U15412 (N_15412,N_13658,N_12685);
xor U15413 (N_15413,N_13875,N_13807);
xnor U15414 (N_15414,N_13811,N_13958);
xnor U15415 (N_15415,N_13029,N_13671);
and U15416 (N_15416,N_13521,N_12127);
xnor U15417 (N_15417,N_12475,N_13503);
or U15418 (N_15418,N_12200,N_12486);
xnor U15419 (N_15419,N_12106,N_13832);
and U15420 (N_15420,N_12916,N_12811);
nor U15421 (N_15421,N_12322,N_13902);
nor U15422 (N_15422,N_13317,N_13066);
xnor U15423 (N_15423,N_12981,N_13085);
or U15424 (N_15424,N_12543,N_13172);
xnor U15425 (N_15425,N_13125,N_12648);
xor U15426 (N_15426,N_13144,N_12124);
nor U15427 (N_15427,N_13078,N_12521);
nor U15428 (N_15428,N_13583,N_13902);
nand U15429 (N_15429,N_13231,N_12472);
and U15430 (N_15430,N_13532,N_13441);
nor U15431 (N_15431,N_13216,N_12178);
and U15432 (N_15432,N_12909,N_12244);
or U15433 (N_15433,N_13953,N_12340);
and U15434 (N_15434,N_12302,N_12287);
xnor U15435 (N_15435,N_13021,N_12148);
and U15436 (N_15436,N_12037,N_13947);
xnor U15437 (N_15437,N_12588,N_12482);
xnor U15438 (N_15438,N_13255,N_13872);
nor U15439 (N_15439,N_13796,N_13664);
and U15440 (N_15440,N_12972,N_12440);
nand U15441 (N_15441,N_13073,N_12780);
or U15442 (N_15442,N_12806,N_13159);
xor U15443 (N_15443,N_13615,N_13318);
xor U15444 (N_15444,N_12229,N_12886);
or U15445 (N_15445,N_12757,N_12489);
xnor U15446 (N_15446,N_12872,N_13114);
and U15447 (N_15447,N_12179,N_12491);
xnor U15448 (N_15448,N_12760,N_12679);
or U15449 (N_15449,N_12049,N_13524);
and U15450 (N_15450,N_13190,N_12342);
or U15451 (N_15451,N_13724,N_12646);
or U15452 (N_15452,N_12354,N_13873);
xor U15453 (N_15453,N_13983,N_13375);
nor U15454 (N_15454,N_13614,N_12802);
or U15455 (N_15455,N_12010,N_13965);
nor U15456 (N_15456,N_13158,N_13374);
and U15457 (N_15457,N_13834,N_13448);
and U15458 (N_15458,N_12474,N_12067);
and U15459 (N_15459,N_12762,N_12651);
nand U15460 (N_15460,N_12171,N_12411);
nor U15461 (N_15461,N_13824,N_13709);
nor U15462 (N_15462,N_13033,N_13967);
nand U15463 (N_15463,N_13054,N_12900);
nor U15464 (N_15464,N_13663,N_13719);
xor U15465 (N_15465,N_12234,N_13533);
nand U15466 (N_15466,N_13946,N_13709);
xor U15467 (N_15467,N_13643,N_12087);
and U15468 (N_15468,N_12019,N_12978);
nor U15469 (N_15469,N_12420,N_13162);
and U15470 (N_15470,N_13821,N_13651);
nand U15471 (N_15471,N_13131,N_13562);
nand U15472 (N_15472,N_13151,N_13508);
and U15473 (N_15473,N_13438,N_13133);
or U15474 (N_15474,N_12138,N_12650);
nand U15475 (N_15475,N_13413,N_12560);
and U15476 (N_15476,N_12164,N_13518);
xor U15477 (N_15477,N_12291,N_12102);
xor U15478 (N_15478,N_13688,N_12177);
or U15479 (N_15479,N_12219,N_12183);
or U15480 (N_15480,N_12280,N_13305);
nor U15481 (N_15481,N_12035,N_13608);
xor U15482 (N_15482,N_12758,N_13924);
xnor U15483 (N_15483,N_13595,N_12836);
nor U15484 (N_15484,N_12964,N_13747);
xor U15485 (N_15485,N_13276,N_13532);
nor U15486 (N_15486,N_13537,N_12513);
nand U15487 (N_15487,N_12232,N_12069);
and U15488 (N_15488,N_12627,N_12187);
nor U15489 (N_15489,N_13694,N_12799);
or U15490 (N_15490,N_13813,N_12375);
or U15491 (N_15491,N_12148,N_12527);
nand U15492 (N_15492,N_13154,N_12184);
nand U15493 (N_15493,N_13831,N_13290);
or U15494 (N_15494,N_12611,N_13573);
or U15495 (N_15495,N_12969,N_13555);
xnor U15496 (N_15496,N_12738,N_13053);
nand U15497 (N_15497,N_13469,N_13189);
nand U15498 (N_15498,N_13343,N_12669);
or U15499 (N_15499,N_13222,N_12869);
nor U15500 (N_15500,N_12874,N_12605);
xor U15501 (N_15501,N_12546,N_13283);
nand U15502 (N_15502,N_12170,N_12673);
nand U15503 (N_15503,N_12955,N_12919);
and U15504 (N_15504,N_12971,N_12555);
or U15505 (N_15505,N_12441,N_13039);
nor U15506 (N_15506,N_12456,N_12323);
xnor U15507 (N_15507,N_12631,N_12686);
and U15508 (N_15508,N_13013,N_13776);
nor U15509 (N_15509,N_12985,N_12673);
and U15510 (N_15510,N_13378,N_13131);
nand U15511 (N_15511,N_12848,N_13119);
nand U15512 (N_15512,N_13345,N_13870);
xor U15513 (N_15513,N_13471,N_12556);
nand U15514 (N_15514,N_12294,N_12639);
or U15515 (N_15515,N_12901,N_13005);
nor U15516 (N_15516,N_12596,N_12428);
and U15517 (N_15517,N_13158,N_13601);
xnor U15518 (N_15518,N_13872,N_13629);
and U15519 (N_15519,N_12298,N_13368);
nand U15520 (N_15520,N_13138,N_12440);
or U15521 (N_15521,N_12836,N_13954);
nand U15522 (N_15522,N_13380,N_12846);
and U15523 (N_15523,N_12917,N_12759);
and U15524 (N_15524,N_13914,N_13217);
xor U15525 (N_15525,N_12260,N_12000);
xor U15526 (N_15526,N_12656,N_13296);
xnor U15527 (N_15527,N_13459,N_13998);
and U15528 (N_15528,N_13886,N_12114);
nand U15529 (N_15529,N_12798,N_13845);
or U15530 (N_15530,N_13478,N_12538);
and U15531 (N_15531,N_12362,N_12048);
or U15532 (N_15532,N_12983,N_12173);
nor U15533 (N_15533,N_13301,N_13335);
or U15534 (N_15534,N_12099,N_12263);
nand U15535 (N_15535,N_13364,N_13377);
nor U15536 (N_15536,N_12942,N_13042);
nand U15537 (N_15537,N_12969,N_12963);
nor U15538 (N_15538,N_13112,N_13455);
nor U15539 (N_15539,N_13723,N_12530);
and U15540 (N_15540,N_13465,N_12664);
or U15541 (N_15541,N_13768,N_12643);
or U15542 (N_15542,N_13053,N_13504);
and U15543 (N_15543,N_12421,N_12383);
and U15544 (N_15544,N_13438,N_13679);
xor U15545 (N_15545,N_12649,N_13640);
nor U15546 (N_15546,N_12110,N_12403);
nor U15547 (N_15547,N_12459,N_12639);
nor U15548 (N_15548,N_13077,N_12338);
or U15549 (N_15549,N_12067,N_12459);
nand U15550 (N_15550,N_12122,N_12851);
nand U15551 (N_15551,N_12251,N_12806);
xnor U15552 (N_15552,N_12925,N_12349);
nor U15553 (N_15553,N_13315,N_12402);
and U15554 (N_15554,N_13323,N_13252);
and U15555 (N_15555,N_13004,N_13398);
nor U15556 (N_15556,N_13524,N_13890);
xnor U15557 (N_15557,N_12420,N_12335);
and U15558 (N_15558,N_12595,N_12997);
or U15559 (N_15559,N_12870,N_12403);
nor U15560 (N_15560,N_12677,N_12455);
or U15561 (N_15561,N_13386,N_12001);
or U15562 (N_15562,N_13368,N_12102);
nor U15563 (N_15563,N_12748,N_12468);
or U15564 (N_15564,N_13175,N_13837);
nor U15565 (N_15565,N_13046,N_12300);
nand U15566 (N_15566,N_13763,N_12906);
and U15567 (N_15567,N_13359,N_12440);
and U15568 (N_15568,N_13641,N_12732);
xnor U15569 (N_15569,N_12603,N_13792);
nor U15570 (N_15570,N_12079,N_13980);
xor U15571 (N_15571,N_12363,N_13750);
nand U15572 (N_15572,N_12590,N_12752);
or U15573 (N_15573,N_12036,N_13211);
nor U15574 (N_15574,N_12323,N_12160);
nand U15575 (N_15575,N_12575,N_12984);
xnor U15576 (N_15576,N_12605,N_12246);
nand U15577 (N_15577,N_12067,N_13325);
xnor U15578 (N_15578,N_13012,N_12567);
nand U15579 (N_15579,N_13872,N_13740);
nor U15580 (N_15580,N_13532,N_12310);
and U15581 (N_15581,N_12320,N_13932);
or U15582 (N_15582,N_13287,N_12697);
nand U15583 (N_15583,N_13490,N_13126);
xnor U15584 (N_15584,N_12973,N_12621);
nor U15585 (N_15585,N_12498,N_13699);
or U15586 (N_15586,N_13479,N_13017);
or U15587 (N_15587,N_12575,N_12541);
and U15588 (N_15588,N_12781,N_13589);
nand U15589 (N_15589,N_13055,N_12117);
xnor U15590 (N_15590,N_12164,N_12291);
and U15591 (N_15591,N_13400,N_13039);
xor U15592 (N_15592,N_13402,N_13064);
nor U15593 (N_15593,N_12808,N_13199);
xnor U15594 (N_15594,N_12157,N_13501);
nor U15595 (N_15595,N_13259,N_13472);
and U15596 (N_15596,N_12160,N_13891);
and U15597 (N_15597,N_12932,N_12826);
nand U15598 (N_15598,N_13355,N_13845);
nor U15599 (N_15599,N_13947,N_12973);
and U15600 (N_15600,N_13972,N_12558);
xnor U15601 (N_15601,N_12773,N_13257);
or U15602 (N_15602,N_12273,N_12762);
nor U15603 (N_15603,N_12066,N_12791);
nand U15604 (N_15604,N_13117,N_13215);
nor U15605 (N_15605,N_13736,N_13637);
or U15606 (N_15606,N_13460,N_12301);
nand U15607 (N_15607,N_13892,N_12761);
nor U15608 (N_15608,N_13048,N_13715);
and U15609 (N_15609,N_13153,N_12636);
xor U15610 (N_15610,N_13233,N_13420);
nor U15611 (N_15611,N_13126,N_12238);
and U15612 (N_15612,N_13496,N_13003);
nor U15613 (N_15613,N_13723,N_12966);
xnor U15614 (N_15614,N_13010,N_12606);
or U15615 (N_15615,N_13974,N_12573);
nand U15616 (N_15616,N_12587,N_12416);
nor U15617 (N_15617,N_13668,N_13876);
xor U15618 (N_15618,N_12807,N_12891);
nand U15619 (N_15619,N_13555,N_12054);
nand U15620 (N_15620,N_13228,N_12662);
and U15621 (N_15621,N_12223,N_13098);
nor U15622 (N_15622,N_13561,N_13824);
nor U15623 (N_15623,N_12619,N_12330);
nor U15624 (N_15624,N_13038,N_13791);
nor U15625 (N_15625,N_12721,N_13990);
or U15626 (N_15626,N_13853,N_12346);
xnor U15627 (N_15627,N_13130,N_13238);
xor U15628 (N_15628,N_12195,N_13083);
nand U15629 (N_15629,N_13811,N_13520);
and U15630 (N_15630,N_13851,N_13599);
and U15631 (N_15631,N_13584,N_12630);
nor U15632 (N_15632,N_13515,N_13637);
xor U15633 (N_15633,N_12577,N_13391);
and U15634 (N_15634,N_13341,N_12664);
nand U15635 (N_15635,N_13130,N_12275);
nand U15636 (N_15636,N_12433,N_13039);
nor U15637 (N_15637,N_12034,N_12206);
or U15638 (N_15638,N_13986,N_13989);
nand U15639 (N_15639,N_13085,N_12684);
or U15640 (N_15640,N_13307,N_12001);
nand U15641 (N_15641,N_13953,N_13586);
nor U15642 (N_15642,N_12874,N_13593);
xor U15643 (N_15643,N_13640,N_12572);
or U15644 (N_15644,N_12139,N_12128);
xnor U15645 (N_15645,N_12485,N_13810);
and U15646 (N_15646,N_13196,N_13195);
and U15647 (N_15647,N_13602,N_12635);
xnor U15648 (N_15648,N_12884,N_12007);
nor U15649 (N_15649,N_12667,N_13741);
and U15650 (N_15650,N_12277,N_13231);
and U15651 (N_15651,N_13528,N_12309);
nor U15652 (N_15652,N_13536,N_12029);
xor U15653 (N_15653,N_13647,N_13618);
nor U15654 (N_15654,N_12246,N_13624);
xnor U15655 (N_15655,N_12706,N_13215);
nor U15656 (N_15656,N_12662,N_13297);
and U15657 (N_15657,N_13654,N_12876);
nand U15658 (N_15658,N_12230,N_12378);
nor U15659 (N_15659,N_12936,N_13623);
xor U15660 (N_15660,N_12058,N_13900);
and U15661 (N_15661,N_13405,N_13775);
and U15662 (N_15662,N_12348,N_13840);
nor U15663 (N_15663,N_13383,N_12402);
or U15664 (N_15664,N_12373,N_12640);
xnor U15665 (N_15665,N_13572,N_12269);
or U15666 (N_15666,N_13774,N_13756);
or U15667 (N_15667,N_12370,N_12501);
nand U15668 (N_15668,N_12389,N_12515);
nand U15669 (N_15669,N_13544,N_12680);
or U15670 (N_15670,N_12925,N_12641);
nor U15671 (N_15671,N_13424,N_12821);
nand U15672 (N_15672,N_13788,N_13236);
and U15673 (N_15673,N_13615,N_13247);
or U15674 (N_15674,N_13885,N_13304);
or U15675 (N_15675,N_12199,N_13744);
nor U15676 (N_15676,N_13822,N_12791);
or U15677 (N_15677,N_12365,N_12603);
or U15678 (N_15678,N_12064,N_13106);
and U15679 (N_15679,N_12618,N_13893);
nand U15680 (N_15680,N_13533,N_13837);
and U15681 (N_15681,N_12061,N_13440);
and U15682 (N_15682,N_12273,N_13422);
nand U15683 (N_15683,N_13375,N_13197);
nand U15684 (N_15684,N_13236,N_12126);
xnor U15685 (N_15685,N_12488,N_12556);
xor U15686 (N_15686,N_13675,N_12540);
xnor U15687 (N_15687,N_13118,N_12011);
nand U15688 (N_15688,N_12712,N_13728);
nor U15689 (N_15689,N_13419,N_12027);
nand U15690 (N_15690,N_12632,N_12279);
and U15691 (N_15691,N_12644,N_12557);
nor U15692 (N_15692,N_12521,N_12265);
xnor U15693 (N_15693,N_12337,N_12749);
nand U15694 (N_15694,N_12701,N_12187);
nand U15695 (N_15695,N_13853,N_12664);
or U15696 (N_15696,N_13802,N_13306);
xor U15697 (N_15697,N_12963,N_13803);
xor U15698 (N_15698,N_12850,N_13376);
nor U15699 (N_15699,N_13046,N_13689);
nand U15700 (N_15700,N_12764,N_12265);
and U15701 (N_15701,N_13244,N_13726);
nor U15702 (N_15702,N_13744,N_12974);
nand U15703 (N_15703,N_13149,N_12889);
or U15704 (N_15704,N_13718,N_13282);
or U15705 (N_15705,N_12566,N_13864);
xor U15706 (N_15706,N_12257,N_12873);
nor U15707 (N_15707,N_13015,N_13631);
nor U15708 (N_15708,N_12401,N_12301);
xor U15709 (N_15709,N_13265,N_12820);
nand U15710 (N_15710,N_13470,N_12921);
and U15711 (N_15711,N_12251,N_12256);
and U15712 (N_15712,N_12982,N_13587);
nor U15713 (N_15713,N_12874,N_13685);
nor U15714 (N_15714,N_12866,N_12961);
xnor U15715 (N_15715,N_12827,N_13963);
xor U15716 (N_15716,N_13732,N_13939);
nor U15717 (N_15717,N_12196,N_12986);
xnor U15718 (N_15718,N_13483,N_13783);
xor U15719 (N_15719,N_13389,N_12927);
nor U15720 (N_15720,N_13563,N_12774);
or U15721 (N_15721,N_12997,N_12678);
xnor U15722 (N_15722,N_12869,N_12261);
nor U15723 (N_15723,N_13013,N_12146);
nor U15724 (N_15724,N_13006,N_12941);
or U15725 (N_15725,N_13439,N_13706);
xor U15726 (N_15726,N_12185,N_13634);
and U15727 (N_15727,N_12038,N_13747);
or U15728 (N_15728,N_13635,N_12502);
xnor U15729 (N_15729,N_12152,N_13363);
or U15730 (N_15730,N_13795,N_13189);
nand U15731 (N_15731,N_12089,N_12771);
nor U15732 (N_15732,N_13514,N_13726);
nand U15733 (N_15733,N_13111,N_12830);
xnor U15734 (N_15734,N_13180,N_12489);
xnor U15735 (N_15735,N_12737,N_12979);
xor U15736 (N_15736,N_13319,N_12827);
nand U15737 (N_15737,N_13397,N_12815);
or U15738 (N_15738,N_12026,N_13637);
nand U15739 (N_15739,N_12996,N_12668);
nor U15740 (N_15740,N_13347,N_12625);
or U15741 (N_15741,N_13322,N_12536);
nor U15742 (N_15742,N_12947,N_12976);
nor U15743 (N_15743,N_12900,N_13929);
xor U15744 (N_15744,N_13908,N_13505);
xor U15745 (N_15745,N_13813,N_13146);
nor U15746 (N_15746,N_12348,N_12002);
xnor U15747 (N_15747,N_12555,N_13623);
or U15748 (N_15748,N_12565,N_12389);
nand U15749 (N_15749,N_13281,N_13114);
and U15750 (N_15750,N_12491,N_13509);
nand U15751 (N_15751,N_13646,N_13988);
nand U15752 (N_15752,N_13270,N_12889);
and U15753 (N_15753,N_12023,N_12825);
xor U15754 (N_15754,N_13128,N_12668);
and U15755 (N_15755,N_12612,N_12144);
xor U15756 (N_15756,N_13626,N_12696);
xor U15757 (N_15757,N_12821,N_13510);
and U15758 (N_15758,N_13240,N_12098);
xnor U15759 (N_15759,N_12270,N_12679);
nor U15760 (N_15760,N_13135,N_13838);
and U15761 (N_15761,N_12625,N_12629);
nor U15762 (N_15762,N_12261,N_13582);
nand U15763 (N_15763,N_13365,N_13746);
nor U15764 (N_15764,N_13001,N_12189);
xor U15765 (N_15765,N_13743,N_13091);
nand U15766 (N_15766,N_12588,N_12726);
nand U15767 (N_15767,N_12686,N_13523);
or U15768 (N_15768,N_13199,N_13840);
and U15769 (N_15769,N_12575,N_13743);
and U15770 (N_15770,N_13615,N_12304);
nor U15771 (N_15771,N_13402,N_13725);
or U15772 (N_15772,N_12434,N_12023);
or U15773 (N_15773,N_13486,N_13002);
xor U15774 (N_15774,N_13365,N_12969);
or U15775 (N_15775,N_13620,N_12254);
nand U15776 (N_15776,N_13619,N_13913);
nor U15777 (N_15777,N_13234,N_13328);
nor U15778 (N_15778,N_12513,N_12403);
nor U15779 (N_15779,N_12983,N_13676);
nor U15780 (N_15780,N_12271,N_13812);
and U15781 (N_15781,N_13026,N_12335);
or U15782 (N_15782,N_13560,N_13791);
nor U15783 (N_15783,N_12421,N_13089);
or U15784 (N_15784,N_13615,N_13091);
nand U15785 (N_15785,N_12880,N_13346);
xnor U15786 (N_15786,N_13137,N_13761);
nor U15787 (N_15787,N_12111,N_12032);
nand U15788 (N_15788,N_12441,N_13648);
nor U15789 (N_15789,N_13438,N_12226);
or U15790 (N_15790,N_13387,N_13396);
nor U15791 (N_15791,N_12997,N_13406);
and U15792 (N_15792,N_12849,N_12988);
nor U15793 (N_15793,N_13293,N_13890);
or U15794 (N_15794,N_12992,N_13808);
and U15795 (N_15795,N_12547,N_13257);
or U15796 (N_15796,N_12801,N_12634);
nor U15797 (N_15797,N_13801,N_12336);
or U15798 (N_15798,N_13702,N_13376);
nand U15799 (N_15799,N_12912,N_13135);
or U15800 (N_15800,N_12174,N_12995);
nand U15801 (N_15801,N_12836,N_13053);
nor U15802 (N_15802,N_13487,N_13789);
nor U15803 (N_15803,N_12370,N_12913);
nand U15804 (N_15804,N_13058,N_12282);
and U15805 (N_15805,N_13277,N_12580);
and U15806 (N_15806,N_13608,N_13195);
or U15807 (N_15807,N_13658,N_13423);
and U15808 (N_15808,N_12413,N_13554);
or U15809 (N_15809,N_13767,N_13199);
nand U15810 (N_15810,N_13556,N_13637);
nor U15811 (N_15811,N_13812,N_13183);
xnor U15812 (N_15812,N_12651,N_13906);
and U15813 (N_15813,N_12510,N_13521);
nor U15814 (N_15814,N_13843,N_13750);
nand U15815 (N_15815,N_13859,N_13705);
xnor U15816 (N_15816,N_12202,N_13059);
nor U15817 (N_15817,N_13893,N_13409);
nor U15818 (N_15818,N_12724,N_13757);
and U15819 (N_15819,N_13516,N_12431);
or U15820 (N_15820,N_12989,N_13649);
nand U15821 (N_15821,N_12843,N_13934);
and U15822 (N_15822,N_13837,N_13189);
nand U15823 (N_15823,N_12185,N_12256);
nor U15824 (N_15824,N_13959,N_12308);
nor U15825 (N_15825,N_13894,N_13412);
and U15826 (N_15826,N_13602,N_12852);
xnor U15827 (N_15827,N_13804,N_13016);
and U15828 (N_15828,N_13487,N_13783);
or U15829 (N_15829,N_13707,N_13448);
nand U15830 (N_15830,N_12049,N_12983);
nand U15831 (N_15831,N_13539,N_12134);
or U15832 (N_15832,N_13828,N_12807);
nand U15833 (N_15833,N_13350,N_12070);
nor U15834 (N_15834,N_12003,N_12170);
nor U15835 (N_15835,N_12366,N_13232);
or U15836 (N_15836,N_13346,N_12521);
nand U15837 (N_15837,N_12718,N_12303);
or U15838 (N_15838,N_12529,N_12910);
and U15839 (N_15839,N_13982,N_13412);
nor U15840 (N_15840,N_12498,N_13743);
and U15841 (N_15841,N_13649,N_13645);
nor U15842 (N_15842,N_13212,N_12523);
nor U15843 (N_15843,N_13956,N_13027);
xnor U15844 (N_15844,N_12430,N_12471);
nor U15845 (N_15845,N_12130,N_13215);
nor U15846 (N_15846,N_12762,N_13170);
nand U15847 (N_15847,N_12516,N_12813);
or U15848 (N_15848,N_13549,N_13350);
or U15849 (N_15849,N_12708,N_13872);
xnor U15850 (N_15850,N_12816,N_12452);
or U15851 (N_15851,N_12683,N_12596);
or U15852 (N_15852,N_12330,N_12261);
xnor U15853 (N_15853,N_12833,N_12148);
nor U15854 (N_15854,N_13152,N_13690);
nor U15855 (N_15855,N_13833,N_12860);
and U15856 (N_15856,N_12070,N_13393);
or U15857 (N_15857,N_12248,N_13352);
xor U15858 (N_15858,N_13569,N_13762);
and U15859 (N_15859,N_13292,N_13231);
nand U15860 (N_15860,N_13987,N_13442);
and U15861 (N_15861,N_13418,N_12997);
and U15862 (N_15862,N_12781,N_13994);
or U15863 (N_15863,N_12871,N_13111);
or U15864 (N_15864,N_13233,N_12324);
xnor U15865 (N_15865,N_12774,N_13068);
or U15866 (N_15866,N_12008,N_13221);
or U15867 (N_15867,N_12594,N_12203);
nor U15868 (N_15868,N_12975,N_12920);
xnor U15869 (N_15869,N_13753,N_12225);
and U15870 (N_15870,N_13498,N_13823);
nor U15871 (N_15871,N_13226,N_13292);
or U15872 (N_15872,N_13631,N_12404);
nor U15873 (N_15873,N_12572,N_13016);
xnor U15874 (N_15874,N_12105,N_12183);
xnor U15875 (N_15875,N_13856,N_12048);
or U15876 (N_15876,N_13574,N_13846);
nor U15877 (N_15877,N_12716,N_13391);
or U15878 (N_15878,N_13023,N_13370);
and U15879 (N_15879,N_13928,N_13197);
nand U15880 (N_15880,N_12277,N_13382);
or U15881 (N_15881,N_13768,N_13703);
nand U15882 (N_15882,N_12272,N_12920);
and U15883 (N_15883,N_12305,N_13090);
or U15884 (N_15884,N_13213,N_13262);
and U15885 (N_15885,N_12778,N_12879);
xor U15886 (N_15886,N_13056,N_12056);
nor U15887 (N_15887,N_13290,N_13759);
xnor U15888 (N_15888,N_12133,N_12506);
or U15889 (N_15889,N_13690,N_12987);
nor U15890 (N_15890,N_12641,N_12740);
and U15891 (N_15891,N_12129,N_13729);
and U15892 (N_15892,N_13959,N_13190);
nand U15893 (N_15893,N_13002,N_13335);
nand U15894 (N_15894,N_12838,N_13992);
xor U15895 (N_15895,N_13381,N_12600);
xnor U15896 (N_15896,N_12306,N_12541);
nand U15897 (N_15897,N_13413,N_13152);
nor U15898 (N_15898,N_12736,N_12509);
nor U15899 (N_15899,N_13847,N_13103);
nand U15900 (N_15900,N_13203,N_13477);
and U15901 (N_15901,N_13185,N_12917);
or U15902 (N_15902,N_12515,N_12461);
and U15903 (N_15903,N_12571,N_13088);
nand U15904 (N_15904,N_12459,N_13953);
nand U15905 (N_15905,N_12095,N_12908);
and U15906 (N_15906,N_13900,N_12310);
and U15907 (N_15907,N_12670,N_12095);
xnor U15908 (N_15908,N_13995,N_12870);
or U15909 (N_15909,N_13152,N_13723);
and U15910 (N_15910,N_12656,N_13870);
and U15911 (N_15911,N_13098,N_12491);
nand U15912 (N_15912,N_12660,N_12217);
or U15913 (N_15913,N_12923,N_12626);
and U15914 (N_15914,N_13740,N_12463);
xnor U15915 (N_15915,N_13777,N_13459);
nand U15916 (N_15916,N_12769,N_12973);
or U15917 (N_15917,N_13267,N_13611);
nand U15918 (N_15918,N_13843,N_12798);
or U15919 (N_15919,N_13558,N_12534);
nand U15920 (N_15920,N_12673,N_12373);
nor U15921 (N_15921,N_13286,N_12765);
nor U15922 (N_15922,N_13207,N_13770);
xor U15923 (N_15923,N_13979,N_13177);
and U15924 (N_15924,N_12179,N_12884);
or U15925 (N_15925,N_13000,N_12016);
nor U15926 (N_15926,N_13895,N_12741);
or U15927 (N_15927,N_13454,N_12436);
or U15928 (N_15928,N_12000,N_12020);
nor U15929 (N_15929,N_13000,N_12495);
xnor U15930 (N_15930,N_12348,N_12571);
xnor U15931 (N_15931,N_12568,N_13440);
and U15932 (N_15932,N_12015,N_12748);
nand U15933 (N_15933,N_13835,N_13215);
or U15934 (N_15934,N_13733,N_13727);
and U15935 (N_15935,N_13386,N_12177);
xnor U15936 (N_15936,N_12614,N_12425);
or U15937 (N_15937,N_12630,N_13335);
or U15938 (N_15938,N_12076,N_13795);
xor U15939 (N_15939,N_13407,N_13309);
xnor U15940 (N_15940,N_13137,N_13209);
nor U15941 (N_15941,N_13909,N_13928);
and U15942 (N_15942,N_12257,N_13066);
or U15943 (N_15943,N_12995,N_12304);
and U15944 (N_15944,N_13780,N_13382);
and U15945 (N_15945,N_13448,N_12504);
nand U15946 (N_15946,N_12369,N_13683);
nor U15947 (N_15947,N_12030,N_13217);
or U15948 (N_15948,N_13405,N_13583);
nor U15949 (N_15949,N_12261,N_12640);
nor U15950 (N_15950,N_13663,N_13677);
xnor U15951 (N_15951,N_13455,N_13157);
and U15952 (N_15952,N_12196,N_13525);
nor U15953 (N_15953,N_13668,N_12006);
or U15954 (N_15954,N_12975,N_12310);
and U15955 (N_15955,N_12579,N_13409);
or U15956 (N_15956,N_13490,N_12352);
nor U15957 (N_15957,N_13726,N_12999);
xor U15958 (N_15958,N_13955,N_13780);
or U15959 (N_15959,N_13658,N_12672);
or U15960 (N_15960,N_13650,N_13645);
nor U15961 (N_15961,N_13812,N_12686);
nor U15962 (N_15962,N_12650,N_12809);
or U15963 (N_15963,N_12756,N_13878);
or U15964 (N_15964,N_13584,N_12624);
nor U15965 (N_15965,N_12985,N_13161);
nor U15966 (N_15966,N_13803,N_12269);
nor U15967 (N_15967,N_13682,N_12004);
xnor U15968 (N_15968,N_12793,N_12424);
or U15969 (N_15969,N_13912,N_13032);
nor U15970 (N_15970,N_13425,N_12599);
nor U15971 (N_15971,N_12718,N_13626);
xor U15972 (N_15972,N_12881,N_12137);
or U15973 (N_15973,N_12742,N_12855);
or U15974 (N_15974,N_12891,N_12597);
xnor U15975 (N_15975,N_12148,N_13122);
nand U15976 (N_15976,N_13810,N_13774);
or U15977 (N_15977,N_13779,N_13879);
and U15978 (N_15978,N_13423,N_13566);
nor U15979 (N_15979,N_12255,N_12362);
or U15980 (N_15980,N_13906,N_13642);
and U15981 (N_15981,N_13510,N_12191);
nor U15982 (N_15982,N_12524,N_13656);
nor U15983 (N_15983,N_13861,N_12697);
xnor U15984 (N_15984,N_13298,N_12854);
and U15985 (N_15985,N_12248,N_13118);
xnor U15986 (N_15986,N_12915,N_13436);
nand U15987 (N_15987,N_12415,N_12833);
and U15988 (N_15988,N_12176,N_12298);
or U15989 (N_15989,N_13899,N_12580);
nand U15990 (N_15990,N_12225,N_13714);
nor U15991 (N_15991,N_12685,N_13766);
nor U15992 (N_15992,N_13019,N_13971);
nor U15993 (N_15993,N_13876,N_13697);
nor U15994 (N_15994,N_12469,N_13299);
or U15995 (N_15995,N_13039,N_13546);
or U15996 (N_15996,N_12985,N_12110);
nor U15997 (N_15997,N_13340,N_12114);
nor U15998 (N_15998,N_13070,N_12283);
and U15999 (N_15999,N_12000,N_13659);
xor U16000 (N_16000,N_15252,N_14991);
or U16001 (N_16001,N_15361,N_15853);
and U16002 (N_16002,N_14888,N_14900);
xnor U16003 (N_16003,N_15593,N_15752);
nand U16004 (N_16004,N_14213,N_14621);
xor U16005 (N_16005,N_14580,N_14251);
nor U16006 (N_16006,N_15193,N_15538);
nand U16007 (N_16007,N_14185,N_15598);
and U16008 (N_16008,N_15787,N_15207);
and U16009 (N_16009,N_14723,N_15984);
nand U16010 (N_16010,N_15269,N_14980);
xnor U16011 (N_16011,N_15052,N_15778);
or U16012 (N_16012,N_15905,N_14081);
xor U16013 (N_16013,N_14042,N_15917);
or U16014 (N_16014,N_14082,N_15619);
xnor U16015 (N_16015,N_14786,N_15099);
and U16016 (N_16016,N_15213,N_15795);
or U16017 (N_16017,N_15459,N_14170);
or U16018 (N_16018,N_14003,N_15203);
or U16019 (N_16019,N_14499,N_15974);
or U16020 (N_16020,N_14222,N_14891);
xnor U16021 (N_16021,N_15492,N_14628);
nor U16022 (N_16022,N_15955,N_15500);
or U16023 (N_16023,N_14243,N_15676);
nor U16024 (N_16024,N_15146,N_14393);
xor U16025 (N_16025,N_14895,N_14138);
nand U16026 (N_16026,N_15864,N_15703);
nor U16027 (N_16027,N_15686,N_15507);
nor U16028 (N_16028,N_14121,N_15910);
xnor U16029 (N_16029,N_14157,N_15541);
nand U16030 (N_16030,N_15005,N_15401);
and U16031 (N_16031,N_14369,N_14007);
nor U16032 (N_16032,N_15161,N_14982);
nand U16033 (N_16033,N_15840,N_14406);
and U16034 (N_16034,N_15986,N_14261);
and U16035 (N_16035,N_14533,N_14549);
nor U16036 (N_16036,N_15334,N_15165);
or U16037 (N_16037,N_14716,N_15468);
or U16038 (N_16038,N_14504,N_14464);
nand U16039 (N_16039,N_14180,N_15596);
or U16040 (N_16040,N_14748,N_15384);
and U16041 (N_16041,N_15025,N_15808);
nor U16042 (N_16042,N_15960,N_14355);
nand U16043 (N_16043,N_15822,N_15738);
xor U16044 (N_16044,N_14939,N_15914);
nor U16045 (N_16045,N_15043,N_15101);
nand U16046 (N_16046,N_15994,N_14932);
or U16047 (N_16047,N_15510,N_15713);
and U16048 (N_16048,N_14266,N_15368);
xor U16049 (N_16049,N_14061,N_14139);
and U16050 (N_16050,N_14233,N_15728);
nor U16051 (N_16051,N_15545,N_14951);
or U16052 (N_16052,N_15457,N_14855);
or U16053 (N_16053,N_15897,N_15532);
nand U16054 (N_16054,N_14290,N_15751);
xnor U16055 (N_16055,N_15668,N_15402);
or U16056 (N_16056,N_14218,N_14709);
and U16057 (N_16057,N_14445,N_15606);
nand U16058 (N_16058,N_15559,N_14682);
nor U16059 (N_16059,N_14732,N_15259);
nand U16060 (N_16060,N_14777,N_14197);
xnor U16061 (N_16061,N_14426,N_14526);
and U16062 (N_16062,N_15879,N_15815);
or U16063 (N_16063,N_15341,N_14642);
or U16064 (N_16064,N_14427,N_14946);
nand U16065 (N_16065,N_14800,N_14944);
or U16066 (N_16066,N_14017,N_14196);
xor U16067 (N_16067,N_15968,N_15925);
or U16068 (N_16068,N_15178,N_15022);
nand U16069 (N_16069,N_15153,N_14662);
or U16070 (N_16070,N_15659,N_15015);
nor U16071 (N_16071,N_14490,N_14816);
nor U16072 (N_16072,N_14027,N_15944);
or U16073 (N_16073,N_15965,N_14713);
nand U16074 (N_16074,N_14351,N_15961);
nand U16075 (N_16075,N_15313,N_14189);
xor U16076 (N_16076,N_15154,N_15527);
xnor U16077 (N_16077,N_15571,N_14764);
nand U16078 (N_16078,N_15243,N_14433);
xor U16079 (N_16079,N_14485,N_14738);
or U16080 (N_16080,N_15087,N_14765);
xor U16081 (N_16081,N_14000,N_14563);
nand U16082 (N_16082,N_15376,N_14238);
nand U16083 (N_16083,N_15764,N_14740);
xor U16084 (N_16084,N_14179,N_14651);
or U16085 (N_16085,N_15958,N_14320);
xor U16086 (N_16086,N_15066,N_15589);
nand U16087 (N_16087,N_14616,N_14190);
nand U16088 (N_16088,N_15836,N_15031);
xor U16089 (N_16089,N_15236,N_15581);
xnor U16090 (N_16090,N_15997,N_14408);
nand U16091 (N_16091,N_15913,N_14497);
nand U16092 (N_16092,N_15705,N_14404);
or U16093 (N_16093,N_15851,N_14273);
nand U16094 (N_16094,N_14542,N_15938);
xor U16095 (N_16095,N_15192,N_15184);
nand U16096 (N_16096,N_14309,N_15274);
or U16097 (N_16097,N_15328,N_15518);
nand U16098 (N_16098,N_15338,N_14057);
and U16099 (N_16099,N_15565,N_14609);
nor U16100 (N_16100,N_14399,N_14114);
and U16101 (N_16101,N_14739,N_14931);
and U16102 (N_16102,N_15880,N_14669);
nand U16103 (N_16103,N_14085,N_14921);
nand U16104 (N_16104,N_14594,N_15075);
nand U16105 (N_16105,N_14817,N_14650);
or U16106 (N_16106,N_14286,N_14859);
or U16107 (N_16107,N_15803,N_14502);
nand U16108 (N_16108,N_14488,N_14354);
and U16109 (N_16109,N_15516,N_15360);
xor U16110 (N_16110,N_14249,N_14768);
or U16111 (N_16111,N_15786,N_15050);
or U16112 (N_16112,N_15824,N_14819);
xor U16113 (N_16113,N_15455,N_14152);
xor U16114 (N_16114,N_15172,N_15119);
and U16115 (N_16115,N_15284,N_15158);
xnor U16116 (N_16116,N_15688,N_15734);
and U16117 (N_16117,N_15973,N_14566);
nor U16118 (N_16118,N_14582,N_14903);
or U16119 (N_16119,N_15859,N_14592);
nor U16120 (N_16120,N_15117,N_15051);
or U16121 (N_16121,N_14443,N_14648);
nand U16122 (N_16122,N_15520,N_15749);
or U16123 (N_16123,N_14176,N_14687);
and U16124 (N_16124,N_15980,N_14323);
nand U16125 (N_16125,N_14788,N_15215);
or U16126 (N_16126,N_15448,N_14572);
nor U16127 (N_16127,N_15414,N_14094);
and U16128 (N_16128,N_15471,N_15077);
and U16129 (N_16129,N_15497,N_14407);
nand U16130 (N_16130,N_14242,N_14230);
nand U16131 (N_16131,N_15428,N_15354);
nor U16132 (N_16132,N_14269,N_14348);
or U16133 (N_16133,N_14008,N_14937);
nor U16134 (N_16134,N_15273,N_15489);
xnor U16135 (N_16135,N_14342,N_15018);
xnor U16136 (N_16136,N_14289,N_14071);
nor U16137 (N_16137,N_14904,N_14102);
nand U16138 (N_16138,N_15232,N_15693);
nand U16139 (N_16139,N_15970,N_14759);
xnor U16140 (N_16140,N_15297,N_15763);
nand U16141 (N_16141,N_14078,N_14164);
xnor U16142 (N_16142,N_15180,N_15941);
or U16143 (N_16143,N_15903,N_14851);
or U16144 (N_16144,N_14885,N_15060);
nor U16145 (N_16145,N_15307,N_15198);
or U16146 (N_16146,N_14599,N_15057);
and U16147 (N_16147,N_15138,N_15814);
or U16148 (N_16148,N_15181,N_15791);
and U16149 (N_16149,N_14097,N_14161);
nor U16150 (N_16150,N_15271,N_15927);
xor U16151 (N_16151,N_15512,N_15476);
and U16152 (N_16152,N_14292,N_14675);
or U16153 (N_16153,N_14935,N_14610);
or U16154 (N_16154,N_15535,N_14298);
nand U16155 (N_16155,N_15023,N_14147);
nor U16156 (N_16156,N_14612,N_15936);
or U16157 (N_16157,N_15280,N_15542);
nand U16158 (N_16158,N_15849,N_15242);
nand U16159 (N_16159,N_14052,N_14828);
or U16160 (N_16160,N_15648,N_15540);
nor U16161 (N_16161,N_15250,N_14201);
nand U16162 (N_16162,N_15238,N_14391);
and U16163 (N_16163,N_15921,N_15844);
nor U16164 (N_16164,N_14259,N_15386);
or U16165 (N_16165,N_14514,N_14084);
nand U16166 (N_16166,N_15951,N_15590);
or U16167 (N_16167,N_14573,N_15707);
or U16168 (N_16168,N_14608,N_15140);
or U16169 (N_16169,N_14395,N_14118);
nand U16170 (N_16170,N_15353,N_14952);
nand U16171 (N_16171,N_15754,N_14949);
xnor U16172 (N_16172,N_14225,N_15320);
or U16173 (N_16173,N_15079,N_15901);
xnor U16174 (N_16174,N_15987,N_14554);
or U16175 (N_16175,N_15549,N_15094);
or U16176 (N_16176,N_14380,N_15257);
and U16177 (N_16177,N_15682,N_14749);
or U16178 (N_16178,N_14840,N_15852);
nand U16179 (N_16179,N_14571,N_14969);
nor U16180 (N_16180,N_14970,N_14537);
and U16181 (N_16181,N_15244,N_14231);
xor U16182 (N_16182,N_15027,N_14543);
nor U16183 (N_16183,N_15097,N_15331);
nand U16184 (N_16184,N_15335,N_15522);
nand U16185 (N_16185,N_15890,N_14678);
xor U16186 (N_16186,N_14449,N_15318);
nand U16187 (N_16187,N_14334,N_15314);
nand U16188 (N_16188,N_14054,N_15253);
xnor U16189 (N_16189,N_14555,N_15841);
nor U16190 (N_16190,N_15595,N_15976);
and U16191 (N_16191,N_15826,N_15784);
nand U16192 (N_16192,N_15133,N_14950);
and U16193 (N_16193,N_15219,N_14145);
or U16194 (N_16194,N_14524,N_15503);
and U16195 (N_16195,N_14785,N_15644);
nor U16196 (N_16196,N_15486,N_14725);
and U16197 (N_16197,N_14093,N_14479);
nand U16198 (N_16198,N_14034,N_14194);
xor U16199 (N_16199,N_14862,N_14486);
nor U16200 (N_16200,N_15632,N_15744);
xnor U16201 (N_16201,N_15287,N_15209);
or U16202 (N_16202,N_15646,N_14523);
and U16203 (N_16203,N_15139,N_15715);
xor U16204 (N_16204,N_15305,N_14156);
and U16205 (N_16205,N_14367,N_14207);
and U16206 (N_16206,N_14839,N_15332);
or U16207 (N_16207,N_14452,N_14656);
and U16208 (N_16208,N_15775,N_14858);
nand U16209 (N_16209,N_14693,N_14271);
and U16210 (N_16210,N_14753,N_14352);
xnor U16211 (N_16211,N_14328,N_14585);
xor U16212 (N_16212,N_14370,N_14096);
xor U16213 (N_16213,N_15347,N_14297);
nor U16214 (N_16214,N_15689,N_14310);
nand U16215 (N_16215,N_15669,N_14113);
and U16216 (N_16216,N_15926,N_14477);
xnor U16217 (N_16217,N_15964,N_14849);
nor U16218 (N_16218,N_14807,N_14856);
nand U16219 (N_16219,N_14577,N_14235);
and U16220 (N_16220,N_15714,N_15816);
nor U16221 (N_16221,N_14830,N_15700);
nand U16222 (N_16222,N_15010,N_14559);
and U16223 (N_16223,N_15874,N_15316);
xnor U16224 (N_16224,N_15144,N_14468);
or U16225 (N_16225,N_14804,N_14615);
and U16226 (N_16226,N_14316,N_15883);
nand U16227 (N_16227,N_15102,N_14154);
nand U16228 (N_16228,N_14378,N_15760);
and U16229 (N_16229,N_14134,N_14876);
xor U16230 (N_16230,N_15429,N_15706);
xor U16231 (N_16231,N_14945,N_14265);
nor U16232 (N_16232,N_14948,N_15221);
nand U16233 (N_16233,N_14841,N_14624);
nor U16234 (N_16234,N_14232,N_15679);
nand U16235 (N_16235,N_15798,N_14066);
nand U16236 (N_16236,N_15909,N_14493);
and U16237 (N_16237,N_14847,N_15629);
or U16238 (N_16238,N_14663,N_14250);
nor U16239 (N_16239,N_15061,N_15963);
xor U16240 (N_16240,N_14371,N_14453);
nor U16241 (N_16241,N_15828,N_15275);
xnor U16242 (N_16242,N_14569,N_15690);
nor U16243 (N_16243,N_15095,N_14784);
nor U16244 (N_16244,N_15171,N_15090);
xor U16245 (N_16245,N_15548,N_14275);
nor U16246 (N_16246,N_14115,N_15260);
and U16247 (N_16247,N_15074,N_14644);
or U16248 (N_16248,N_14516,N_15317);
and U16249 (N_16249,N_14974,N_14806);
xor U16250 (N_16250,N_14029,N_14984);
xor U16251 (N_16251,N_15266,N_14210);
and U16252 (N_16252,N_14771,N_14133);
and U16253 (N_16253,N_14508,N_15922);
nand U16254 (N_16254,N_15762,N_15829);
xor U16255 (N_16255,N_15641,N_14364);
or U16256 (N_16256,N_15096,N_15400);
xor U16257 (N_16257,N_14155,N_15390);
xor U16258 (N_16258,N_15391,N_14747);
xor U16259 (N_16259,N_14968,N_14347);
xor U16260 (N_16260,N_14002,N_14295);
nand U16261 (N_16261,N_14183,N_14724);
xor U16262 (N_16262,N_14482,N_14023);
nand U16263 (N_16263,N_14270,N_15085);
nor U16264 (N_16264,N_15456,N_15820);
and U16265 (N_16265,N_15159,N_15996);
xor U16266 (N_16266,N_15251,N_14503);
and U16267 (N_16267,N_14229,N_14392);
xnor U16268 (N_16268,N_15191,N_14215);
nand U16269 (N_16269,N_14619,N_14832);
nor U16270 (N_16270,N_15654,N_15792);
or U16271 (N_16271,N_15939,N_15033);
nand U16272 (N_16272,N_14412,N_15506);
nor U16273 (N_16273,N_14424,N_14734);
nand U16274 (N_16274,N_15048,N_15053);
or U16275 (N_16275,N_15560,N_15666);
nor U16276 (N_16276,N_14241,N_15194);
and U16277 (N_16277,N_14032,N_15670);
and U16278 (N_16278,N_15365,N_15416);
or U16279 (N_16279,N_14611,N_14564);
and U16280 (N_16280,N_14127,N_15835);
xor U16281 (N_16281,N_14635,N_15933);
and U16282 (N_16282,N_15604,N_15067);
and U16283 (N_16283,N_15058,N_14613);
and U16284 (N_16284,N_15345,N_14976);
xor U16285 (N_16285,N_14671,N_15531);
nand U16286 (N_16286,N_14415,N_14505);
nand U16287 (N_16287,N_15461,N_15114);
or U16288 (N_16288,N_14198,N_14763);
xnor U16289 (N_16289,N_15674,N_15957);
nand U16290 (N_16290,N_15569,N_15585);
xnor U16291 (N_16291,N_15623,N_15753);
xor U16292 (N_16292,N_15759,N_15245);
or U16293 (N_16293,N_15349,N_15037);
nor U16294 (N_16294,N_14825,N_14743);
xor U16295 (N_16295,N_14660,N_14177);
xor U16296 (N_16296,N_15574,N_15108);
xnor U16297 (N_16297,N_14153,N_14659);
nand U16298 (N_16298,N_14040,N_15672);
nand U16299 (N_16299,N_14792,N_15279);
nor U16300 (N_16300,N_14059,N_15070);
nand U16301 (N_16301,N_14575,N_15126);
nand U16302 (N_16302,N_14532,N_15302);
and U16303 (N_16303,N_14556,N_15054);
xnor U16304 (N_16304,N_14487,N_14869);
nand U16305 (N_16305,N_14212,N_14496);
nand U16306 (N_16306,N_15573,N_14513);
and U16307 (N_16307,N_14691,N_14668);
or U16308 (N_16308,N_15536,N_15256);
xnor U16309 (N_16309,N_14518,N_14587);
nand U16310 (N_16310,N_14857,N_15240);
nand U16311 (N_16311,N_14353,N_15105);
or U16312 (N_16312,N_14398,N_14998);
nor U16313 (N_16313,N_14964,N_14755);
xnor U16314 (N_16314,N_14820,N_14252);
or U16315 (N_16315,N_14882,N_14603);
nor U16316 (N_16316,N_14489,N_14538);
xnor U16317 (N_16317,N_15602,N_14924);
or U16318 (N_16318,N_14462,N_15121);
nand U16319 (N_16319,N_14208,N_14861);
and U16320 (N_16320,N_15130,N_14247);
and U16321 (N_16321,N_15785,N_14962);
nor U16322 (N_16322,N_14814,N_14553);
and U16323 (N_16323,N_14751,N_15296);
nand U16324 (N_16324,N_14961,N_14907);
or U16325 (N_16325,N_14824,N_14448);
nand U16326 (N_16326,N_14137,N_15867);
or U16327 (N_16327,N_15807,N_15773);
nor U16328 (N_16328,N_15036,N_15479);
or U16329 (N_16329,N_14065,N_15721);
nor U16330 (N_16330,N_15469,N_15233);
nand U16331 (N_16331,N_15230,N_14704);
nand U16332 (N_16332,N_14602,N_15134);
xnor U16333 (N_16333,N_15582,N_14349);
xnor U16334 (N_16334,N_15026,N_15865);
or U16335 (N_16335,N_14385,N_14087);
and U16336 (N_16336,N_15306,N_15222);
nand U16337 (N_16337,N_14983,N_15182);
or U16338 (N_16338,N_15528,N_14776);
or U16339 (N_16339,N_15691,N_14868);
and U16340 (N_16340,N_14469,N_14637);
nand U16341 (N_16341,N_15562,N_14037);
nand U16342 (N_16342,N_14174,N_15356);
and U16343 (N_16343,N_15463,N_14216);
nand U16344 (N_16344,N_15768,N_15127);
or U16345 (N_16345,N_14810,N_15065);
xor U16346 (N_16346,N_15988,N_15854);
nor U16347 (N_16347,N_15810,N_14228);
and U16348 (N_16348,N_14780,N_15285);
or U16349 (N_16349,N_15049,N_15993);
nand U16350 (N_16350,N_15896,N_15626);
nor U16351 (N_16351,N_15726,N_15825);
xnor U16352 (N_16352,N_14793,N_14670);
or U16353 (N_16353,N_14451,N_14836);
and U16354 (N_16354,N_15908,N_14707);
nor U16355 (N_16355,N_15720,N_14267);
nor U16356 (N_16356,N_14975,N_15110);
nand U16357 (N_16357,N_14717,N_14001);
xor U16358 (N_16358,N_15972,N_14745);
or U16359 (N_16359,N_15199,N_15224);
nor U16360 (N_16360,N_14796,N_15592);
or U16361 (N_16361,N_15609,N_14943);
or U16362 (N_16362,N_14500,N_15080);
and U16363 (N_16363,N_14432,N_14035);
and U16364 (N_16364,N_15364,N_15343);
xor U16365 (N_16365,N_15832,N_14160);
xor U16366 (N_16366,N_14940,N_14507);
and U16367 (N_16367,N_14044,N_15782);
or U16368 (N_16368,N_15151,N_15515);
xor U16369 (N_16369,N_15868,N_14902);
or U16370 (N_16370,N_14425,N_15651);
and U16371 (N_16371,N_14004,N_14438);
and U16372 (N_16372,N_14812,N_15480);
nand U16373 (N_16373,N_14586,N_15678);
nor U16374 (N_16374,N_14927,N_15124);
and U16375 (N_16375,N_14301,N_15216);
xor U16376 (N_16376,N_14418,N_14992);
xnor U16377 (N_16377,N_15729,N_14892);
or U16378 (N_16378,N_14540,N_15580);
xnor U16379 (N_16379,N_14760,N_14111);
or U16380 (N_16380,N_14144,N_14973);
nor U16381 (N_16381,N_14423,N_15024);
xnor U16382 (N_16382,N_15451,N_14718);
or U16383 (N_16383,N_14698,N_14068);
nor U16384 (N_16384,N_15949,N_14018);
nor U16385 (N_16385,N_14531,N_14224);
nand U16386 (N_16386,N_15223,N_15697);
and U16387 (N_16387,N_14972,N_14722);
xnor U16388 (N_16388,N_14649,N_15157);
nand U16389 (N_16389,N_15856,N_14798);
and U16390 (N_16390,N_14996,N_14654);
nand U16391 (N_16391,N_14521,N_14421);
xnor U16392 (N_16392,N_14545,N_14712);
and U16393 (N_16393,N_14607,N_15104);
or U16394 (N_16394,N_15385,N_15603);
nand U16395 (N_16395,N_14633,N_14844);
nand U16396 (N_16396,N_14278,N_15501);
nor U16397 (N_16397,N_15757,N_14064);
or U16398 (N_16398,N_15911,N_15575);
nand U16399 (N_16399,N_15149,N_15712);
or U16400 (N_16400,N_14255,N_15442);
or U16401 (N_16401,N_15292,N_14695);
nor U16402 (N_16402,N_15664,N_15387);
nor U16403 (N_16403,N_15197,N_15467);
and U16404 (N_16404,N_14430,N_14597);
nor U16405 (N_16405,N_15612,N_14730);
xnor U16406 (N_16406,N_15931,N_15427);
xor U16407 (N_16407,N_15942,N_14396);
nand U16408 (N_16408,N_15152,N_15635);
and U16409 (N_16409,N_15089,N_15838);
and U16410 (N_16410,N_15444,N_14471);
nand U16411 (N_16411,N_14519,N_15267);
nor U16412 (N_16412,N_14770,N_14481);
nand U16413 (N_16413,N_15355,N_14509);
and U16414 (N_16414,N_15329,N_14359);
and U16415 (N_16415,N_15568,N_15711);
xor U16416 (N_16416,N_15310,N_15556);
nand U16417 (N_16417,N_15981,N_14282);
and U16418 (N_16418,N_15381,N_14262);
nand U16419 (N_16419,N_14645,N_14813);
nor U16420 (N_16420,N_14576,N_14886);
nor U16421 (N_16421,N_15561,N_14604);
xnor U16422 (N_16422,N_14994,N_15016);
xor U16423 (N_16423,N_14165,N_15484);
and U16424 (N_16424,N_15796,N_14986);
or U16425 (N_16425,N_15966,N_15150);
nand U16426 (N_16426,N_14304,N_14036);
and U16427 (N_16427,N_14120,N_15881);
and U16428 (N_16428,N_14220,N_15587);
xor U16429 (N_16429,N_14429,N_14492);
or U16430 (N_16430,N_14331,N_14256);
xor U16431 (N_16431,N_15876,N_15290);
nor U16432 (N_16432,N_15483,N_14458);
or U16433 (N_16433,N_14182,N_14963);
and U16434 (N_16434,N_15550,N_14205);
and U16435 (N_16435,N_15372,N_15702);
nand U16436 (N_16436,N_15817,N_15382);
or U16437 (N_16437,N_15742,N_15790);
or U16438 (N_16438,N_15336,N_15954);
or U16439 (N_16439,N_15107,N_15657);
or U16440 (N_16440,N_14570,N_15430);
and U16441 (N_16441,N_15009,N_14890);
nand U16442 (N_16442,N_15680,N_14667);
or U16443 (N_16443,N_14442,N_15147);
nor U16444 (N_16444,N_14827,N_15723);
and U16445 (N_16445,N_14305,N_14846);
and U16446 (N_16446,N_15142,N_14033);
nand U16447 (N_16447,N_15375,N_14794);
nand U16448 (N_16448,N_15247,N_15886);
and U16449 (N_16449,N_14384,N_14063);
and U16450 (N_16450,N_15842,N_14629);
nor U16451 (N_16451,N_15708,N_14799);
nand U16452 (N_16452,N_15268,N_14560);
nor U16453 (N_16453,N_15396,N_14618);
or U16454 (N_16454,N_15068,N_14641);
nor U16455 (N_16455,N_15615,N_14528);
and U16456 (N_16456,N_15201,N_15777);
xor U16457 (N_16457,N_14478,N_15464);
xor U16458 (N_16458,N_14089,N_15299);
and U16459 (N_16459,N_14236,N_14746);
nor U16460 (N_16460,N_15724,N_15611);
xor U16461 (N_16461,N_14646,N_14326);
and U16462 (N_16462,N_14226,N_15999);
nor U16463 (N_16463,N_14506,N_14417);
xor U16464 (N_16464,N_14906,N_15344);
and U16465 (N_16465,N_15630,N_15627);
and U16466 (N_16466,N_15474,N_14731);
xor U16467 (N_16467,N_15918,N_15406);
xor U16468 (N_16468,N_15866,N_15677);
nand U16469 (N_16469,N_15055,N_15979);
nor U16470 (N_16470,N_15028,N_15263);
or U16471 (N_16471,N_14515,N_14593);
and U16472 (N_16472,N_15358,N_15491);
xor U16473 (N_16473,N_14941,N_14446);
nor U16474 (N_16474,N_15405,N_15920);
nand U16475 (N_16475,N_15225,N_15799);
nor U16476 (N_16476,N_14596,N_14631);
nor U16477 (N_16477,N_14522,N_14450);
nand U16478 (N_16478,N_15413,N_14204);
and U16479 (N_16479,N_15935,N_15975);
xnor U16480 (N_16480,N_14439,N_14617);
and U16481 (N_16481,N_15698,N_14159);
nand U16482 (N_16482,N_14248,N_14726);
or U16483 (N_16483,N_15893,N_14080);
nand U16484 (N_16484,N_15505,N_14317);
xnor U16485 (N_16485,N_15877,N_14627);
xnor U16486 (N_16486,N_15719,N_15246);
and U16487 (N_16487,N_14132,N_15433);
and U16488 (N_16488,N_14480,N_14175);
nand U16489 (N_16489,N_14658,N_14172);
nand U16490 (N_16490,N_14108,N_14823);
nor U16491 (N_16491,N_15694,N_15586);
nand U16492 (N_16492,N_15887,N_15989);
nor U16493 (N_16493,N_15132,N_14254);
and U16494 (N_16494,N_15131,N_15465);
or U16495 (N_16495,N_14562,N_15286);
nand U16496 (N_16496,N_14041,N_14428);
and U16497 (N_16497,N_15063,N_15848);
nand U16498 (N_16498,N_14308,N_15684);
or U16499 (N_16499,N_14838,N_14595);
and U16500 (N_16500,N_14899,N_14472);
nand U16501 (N_16501,N_14447,N_15946);
xnor U16502 (N_16502,N_15032,N_15929);
nand U16503 (N_16503,N_14512,N_14729);
and U16504 (N_16504,N_14742,N_14960);
nor U16505 (N_16505,N_15044,N_15681);
xor U16506 (N_16506,N_14021,N_14547);
xnor U16507 (N_16507,N_15440,N_14039);
nand U16508 (N_16508,N_15438,N_15618);
or U16509 (N_16509,N_15017,N_15185);
or U16510 (N_16510,N_15534,N_14284);
nand U16511 (N_16511,N_14677,N_15326);
nor U16512 (N_16512,N_15188,N_14852);
xnor U16513 (N_16513,N_15969,N_15741);
xor U16514 (N_16514,N_15855,N_14676);
and U16515 (N_16515,N_15420,N_15991);
nor U16516 (N_16516,N_14291,N_14956);
nand U16517 (N_16517,N_14100,N_15187);
nor U16518 (N_16518,N_14126,N_14703);
xor U16519 (N_16519,N_14045,N_15733);
or U16520 (N_16520,N_15858,N_14583);
nor U16521 (N_16521,N_14436,N_14541);
nand U16522 (N_16522,N_15350,N_14579);
or U16523 (N_16523,N_14318,N_14337);
nand U16524 (N_16524,N_15953,N_15020);
xor U16525 (N_16525,N_14590,N_14455);
or U16526 (N_16526,N_15059,N_15303);
nor U16527 (N_16527,N_15640,N_14079);
or U16528 (N_16528,N_14083,N_14192);
and U16529 (N_16529,N_15092,N_15291);
nor U16530 (N_16530,N_14062,N_15607);
nand U16531 (N_16531,N_15731,N_14845);
nor U16532 (N_16532,N_14379,N_15437);
or U16533 (N_16533,N_15819,N_14501);
xnor U16534 (N_16534,N_15802,N_14019);
nand U16535 (N_16535,N_14591,N_15493);
xor U16536 (N_16536,N_15478,N_14701);
or U16537 (N_16537,N_14938,N_15870);
nor U16538 (N_16538,N_14377,N_15628);
nor U16539 (N_16539,N_14795,N_15412);
and U16540 (N_16540,N_15177,N_14589);
nand U16541 (N_16541,N_15511,N_14146);
nand U16542 (N_16542,N_14601,N_14614);
xor U16543 (N_16543,N_15488,N_14955);
or U16544 (N_16544,N_15793,N_14005);
nand U16545 (N_16545,N_15293,N_14200);
xor U16546 (N_16546,N_14735,N_15315);
xnor U16547 (N_16547,N_14733,N_15766);
xnor U16548 (N_16548,N_14958,N_14842);
nor U16549 (N_16549,N_15636,N_15649);
nand U16550 (N_16550,N_14680,N_15393);
nand U16551 (N_16551,N_15769,N_14274);
nand U16552 (N_16552,N_15912,N_15449);
xor U16553 (N_16553,N_15398,N_15671);
xor U16554 (N_16554,N_15205,N_15339);
and U16555 (N_16555,N_15620,N_14870);
xor U16556 (N_16556,N_14752,N_14878);
nand U16557 (N_16557,N_15818,N_14474);
or U16558 (N_16558,N_14965,N_14706);
and U16559 (N_16559,N_15823,N_14848);
xnor U16560 (N_16560,N_14652,N_14979);
or U16561 (N_16561,N_15779,N_15034);
xor U16562 (N_16562,N_15195,N_14315);
or U16563 (N_16563,N_14244,N_14894);
nor U16564 (N_16564,N_14544,N_15928);
nand U16565 (N_16565,N_14803,N_15530);
nor U16566 (N_16566,N_14914,N_15956);
and U16567 (N_16567,N_14598,N_15300);
nand U16568 (N_16568,N_15977,N_14674);
and U16569 (N_16569,N_14981,N_15289);
nor U16570 (N_16570,N_15496,N_14313);
xnor U16571 (N_16571,N_15552,N_15915);
nor U16572 (N_16572,N_14917,N_14168);
or U16573 (N_16573,N_15294,N_15389);
or U16574 (N_16574,N_14434,N_14319);
nand U16575 (N_16575,N_14867,N_14330);
or U16576 (N_16576,N_15660,N_15019);
xor U16577 (N_16577,N_15789,N_15116);
and U16578 (N_16578,N_14009,N_14936);
nor U16579 (N_16579,N_15261,N_15426);
and U16580 (N_16580,N_14258,N_15322);
or U16581 (N_16581,N_14413,N_15621);
nor U16582 (N_16582,N_14689,N_14123);
and U16583 (N_16583,N_14142,N_15175);
or U16584 (N_16584,N_14877,N_14774);
xor U16585 (N_16585,N_15091,N_15872);
nand U16586 (N_16586,N_15524,N_15164);
and U16587 (N_16587,N_14708,N_15419);
and U16588 (N_16588,N_14105,N_15517);
or U16589 (N_16589,N_14277,N_14990);
nor U16590 (N_16590,N_14060,N_15176);
nor U16591 (N_16591,N_15717,N_15447);
nor U16592 (N_16592,N_15924,N_15578);
xnor U16593 (N_16593,N_15882,N_15758);
xnor U16594 (N_16594,N_14498,N_15324);
or U16595 (N_16595,N_14779,N_15229);
or U16596 (N_16596,N_14634,N_15579);
xor U16597 (N_16597,N_14069,N_15967);
nand U16598 (N_16598,N_15128,N_15039);
or U16599 (N_16599,N_14107,N_14769);
nor U16600 (N_16600,N_15663,N_14095);
and U16601 (N_16601,N_14638,N_15342);
nand U16602 (N_16602,N_14790,N_15411);
and U16603 (N_16603,N_15502,N_14643);
nor U16604 (N_16604,N_14031,N_14772);
xnor U16605 (N_16605,N_14038,N_15136);
and U16606 (N_16606,N_14929,N_15226);
xnor U16607 (N_16607,N_15656,N_15394);
and U16608 (N_16608,N_14195,N_14829);
and U16609 (N_16609,N_14705,N_15605);
and U16610 (N_16610,N_14227,N_14808);
or U16611 (N_16611,N_15446,N_14557);
and U16612 (N_16612,N_14758,N_15639);
or U16613 (N_16613,N_15827,N_15008);
nand U16614 (N_16614,N_14880,N_15069);
and U16615 (N_16615,N_14345,N_15359);
and U16616 (N_16616,N_15084,N_14715);
or U16617 (N_16617,N_15482,N_15415);
or U16618 (N_16618,N_14112,N_15123);
or U16619 (N_16619,N_14362,N_14510);
and U16620 (N_16620,N_15937,N_14539);
nor U16621 (N_16621,N_15143,N_15083);
nand U16622 (N_16622,N_15900,N_15673);
xnor U16623 (N_16623,N_15539,N_15148);
nand U16624 (N_16624,N_14178,N_15608);
and U16625 (N_16625,N_15812,N_15166);
or U16626 (N_16626,N_15995,N_15473);
xnor U16627 (N_16627,N_15716,N_14293);
nand U16628 (N_16628,N_15687,N_14957);
and U16629 (N_16629,N_14672,N_15748);
nand U16630 (N_16630,N_14150,N_14837);
nor U16631 (N_16631,N_15042,N_15513);
and U16632 (N_16632,N_15323,N_15041);
xnor U16633 (N_16633,N_15950,N_15701);
nand U16634 (N_16634,N_15509,N_15231);
nand U16635 (N_16635,N_15035,N_15813);
xor U16636 (N_16636,N_14167,N_15417);
nor U16637 (N_16637,N_15523,N_14245);
nor U16638 (N_16638,N_14767,N_14299);
and U16639 (N_16639,N_14466,N_14454);
or U16640 (N_16640,N_15543,N_15454);
xor U16641 (N_16641,N_14025,N_14484);
nor U16642 (N_16642,N_14411,N_15470);
nor U16643 (N_16643,N_15658,N_14016);
nor U16644 (N_16644,N_15907,N_15990);
and U16645 (N_16645,N_15780,N_14387);
nand U16646 (N_16646,N_15735,N_15408);
xor U16647 (N_16647,N_14141,N_15410);
xor U16648 (N_16648,N_15650,N_14815);
and U16649 (N_16649,N_14014,N_14874);
xor U16650 (N_16650,N_15521,N_15647);
xnor U16651 (N_16651,N_14101,N_15845);
or U16652 (N_16652,N_14394,N_15869);
xor U16653 (N_16653,N_14140,N_14077);
nor U16654 (N_16654,N_15895,N_15743);
nand U16655 (N_16655,N_15434,N_15529);
and U16656 (N_16656,N_14605,N_15930);
or U16657 (N_16657,N_15030,N_15740);
and U16658 (N_16658,N_14206,N_14551);
xnor U16659 (N_16659,N_15371,N_14022);
nor U16660 (N_16660,N_15722,N_14476);
or U16661 (N_16661,N_15830,N_15241);
and U16662 (N_16662,N_15811,N_14459);
and U16663 (N_16663,N_15472,N_15264);
and U16664 (N_16664,N_14381,N_14344);
nor U16665 (N_16665,N_15173,N_15013);
or U16666 (N_16666,N_15462,N_14401);
nor U16667 (N_16667,N_14075,N_15439);
and U16668 (N_16668,N_15898,N_14221);
and U16669 (N_16669,N_15971,N_15227);
nand U16670 (N_16670,N_15453,N_14728);
nand U16671 (N_16671,N_14681,N_15373);
nor U16672 (N_16672,N_14333,N_15183);
nor U16673 (N_16673,N_14329,N_15378);
nor U16674 (N_16674,N_15774,N_14971);
nand U16675 (N_16675,N_15422,N_14881);
xnor U16676 (N_16676,N_15072,N_14360);
xor U16677 (N_16677,N_15747,N_15435);
or U16678 (N_16678,N_14199,N_15526);
and U16679 (N_16679,N_14757,N_14327);
nand U16680 (N_16680,N_15367,N_14711);
xnor U16681 (N_16681,N_15544,N_14073);
or U16682 (N_16682,N_15667,N_14926);
and U16683 (N_16683,N_15088,N_14376);
or U16684 (N_16684,N_14050,N_14091);
or U16685 (N_16685,N_15254,N_14420);
and U16686 (N_16686,N_15312,N_14416);
and U16687 (N_16687,N_15418,N_15235);
xor U16688 (N_16688,N_15801,N_15098);
nand U16689 (N_16689,N_15397,N_14581);
and U16690 (N_16690,N_15902,N_14440);
or U16691 (N_16691,N_14187,N_15584);
nor U16692 (N_16692,N_14721,N_14473);
xor U16693 (N_16693,N_15888,N_14090);
xnor U16694 (N_16694,N_14287,N_14397);
and U16695 (N_16695,N_15125,N_15661);
and U16696 (N_16696,N_14911,N_15208);
nand U16697 (N_16697,N_15002,N_15234);
and U16698 (N_16698,N_15045,N_15262);
and U16699 (N_16699,N_15380,N_14088);
xor U16700 (N_16700,N_14322,N_14997);
nor U16701 (N_16701,N_14801,N_14910);
xnor U16702 (N_16702,N_15767,N_14928);
and U16703 (N_16703,N_14302,N_14787);
nor U16704 (N_16704,N_15395,N_15519);
nor U16705 (N_16705,N_14632,N_15112);
or U16706 (N_16706,N_14437,N_14744);
nor U16707 (N_16707,N_14223,N_15567);
or U16708 (N_16708,N_15106,N_14527);
nand U16709 (N_16709,N_14809,N_15652);
nor U16710 (N_16710,N_15843,N_15730);
nor U16711 (N_16711,N_15514,N_14802);
xnor U16712 (N_16712,N_14104,N_15404);
nor U16713 (N_16713,N_14169,N_15959);
or U16714 (N_16714,N_14374,N_15466);
xnor U16715 (N_16715,N_14546,N_14389);
and U16716 (N_16716,N_14257,N_15952);
or U16717 (N_16717,N_15369,N_14372);
and U16718 (N_16718,N_15546,N_14296);
nor U16719 (N_16719,N_14163,N_15308);
nand U16720 (N_16720,N_14246,N_15076);
xnor U16721 (N_16721,N_14130,N_14568);
nor U16722 (N_16722,N_15992,N_14475);
nand U16723 (N_16723,N_15217,N_14756);
nor U16724 (N_16724,N_14873,N_14128);
or U16725 (N_16725,N_15062,N_15452);
nor U16726 (N_16726,N_14930,N_14918);
nor U16727 (N_16727,N_15327,N_14999);
and U16728 (N_16728,N_15081,N_14117);
nand U16729 (N_16729,N_14410,N_14116);
nand U16730 (N_16730,N_14696,N_15445);
nor U16731 (N_16731,N_15894,N_15270);
nor U16732 (N_16732,N_14626,N_14098);
nor U16733 (N_16733,N_14306,N_15288);
nand U16734 (N_16734,N_15357,N_14388);
and U16735 (N_16735,N_15304,N_14149);
and U16736 (N_16736,N_14076,N_14444);
nand U16737 (N_16737,N_14630,N_14805);
nor U16738 (N_16738,N_14151,N_14623);
nor U16739 (N_16739,N_14288,N_14915);
or U16740 (N_16740,N_14055,N_14240);
or U16741 (N_16741,N_15346,N_14171);
xnor U16742 (N_16742,N_15553,N_15932);
nand U16743 (N_16743,N_15948,N_14622);
and U16744 (N_16744,N_15739,N_14901);
and U16745 (N_16745,N_15196,N_15403);
nor U16746 (N_16746,N_14122,N_15040);
nor U16747 (N_16747,N_15631,N_15007);
nor U16748 (N_16748,N_15156,N_15837);
nand U16749 (N_16749,N_14993,N_14103);
nor U16750 (N_16750,N_14260,N_14219);
nand U16751 (N_16751,N_15978,N_14390);
nand U16752 (N_16752,N_15135,N_14661);
xor U16753 (N_16753,N_15770,N_14272);
and U16754 (N_16754,N_14209,N_14099);
nor U16755 (N_16755,N_15934,N_15370);
and U16756 (N_16756,N_14831,N_15809);
nor U16757 (N_16757,N_15301,N_14778);
xnor U16758 (N_16758,N_15504,N_15012);
and U16759 (N_16759,N_14191,N_14750);
nand U16760 (N_16760,N_14727,N_15407);
nand U16761 (N_16761,N_15210,N_14335);
and U16762 (N_16762,N_15399,N_15732);
or U16763 (N_16763,N_15564,N_14314);
nor U16764 (N_16764,N_15046,N_14386);
nand U16765 (N_16765,N_15388,N_14463);
nor U16766 (N_16766,N_15737,N_15597);
or U16767 (N_16767,N_14173,N_15736);
or U16768 (N_16768,N_14552,N_15554);
or U16769 (N_16769,N_15889,N_15846);
nand U16770 (N_16770,N_15162,N_14811);
nor U16771 (N_16771,N_14699,N_14865);
and U16772 (N_16772,N_14015,N_14866);
and U16773 (N_16773,N_15137,N_14821);
xor U16774 (N_16774,N_14822,N_14346);
nand U16775 (N_16775,N_15776,N_14129);
xor U16776 (N_16776,N_15599,N_14775);
nor U16777 (N_16777,N_15551,N_14214);
and U16778 (N_16778,N_14860,N_15211);
nand U16779 (N_16779,N_15014,N_14536);
or U16780 (N_16780,N_15064,N_15725);
or U16781 (N_16781,N_14766,N_14186);
xnor U16782 (N_16782,N_14053,N_15570);
or U16783 (N_16783,N_14188,N_15424);
nor U16784 (N_16784,N_15860,N_14056);
and U16785 (N_16785,N_14942,N_14640);
and U16786 (N_16786,N_15189,N_15662);
xor U16787 (N_16787,N_14409,N_14853);
nor U16788 (N_16788,N_14653,N_15475);
or U16789 (N_16789,N_15692,N_15755);
xor U16790 (N_16790,N_15155,N_15600);
xor U16791 (N_16791,N_14340,N_15533);
and U16792 (N_16792,N_15337,N_14339);
and U16793 (N_16793,N_14977,N_14897);
nand U16794 (N_16794,N_15850,N_14584);
nand U16795 (N_16795,N_14923,N_14988);
nand U16796 (N_16796,N_14441,N_15904);
nor U16797 (N_16797,N_14119,N_15141);
nor U16798 (N_16798,N_14686,N_14350);
or U16799 (N_16799,N_14158,N_15485);
and U16800 (N_16800,N_15011,N_15696);
nor U16801 (N_16801,N_15871,N_14465);
or U16802 (N_16802,N_15436,N_14402);
or U16803 (N_16803,N_15348,N_14535);
or U16804 (N_16804,N_14953,N_14781);
xnor U16805 (N_16805,N_15885,N_15572);
nor U16806 (N_16806,N_15122,N_15113);
and U16807 (N_16807,N_15642,N_14736);
or U16808 (N_16808,N_14303,N_14967);
nand U16809 (N_16809,N_14782,N_14363);
and U16810 (N_16810,N_14919,N_15555);
and U16811 (N_16811,N_15298,N_15458);
xnor U16812 (N_16812,N_15174,N_14636);
nand U16813 (N_16813,N_15940,N_14162);
and U16814 (N_16814,N_14072,N_15204);
nand U16815 (N_16815,N_14124,N_14720);
xor U16816 (N_16816,N_15272,N_15985);
and U16817 (N_16817,N_15118,N_14202);
nor U16818 (N_16818,N_15001,N_15321);
xor U16819 (N_16819,N_14639,N_14558);
and U16820 (N_16820,N_14048,N_15494);
nor U16821 (N_16821,N_15746,N_15431);
nor U16822 (N_16822,N_14673,N_14995);
nand U16823 (N_16823,N_15863,N_15258);
or U16824 (N_16824,N_15591,N_15167);
and U16825 (N_16825,N_14383,N_15443);
xor U16826 (N_16826,N_14143,N_14797);
and U16827 (N_16827,N_14606,N_15220);
xnor U16828 (N_16828,N_14234,N_14922);
nor U16829 (N_16829,N_15547,N_14684);
nor U16830 (N_16830,N_15004,N_15919);
or U16831 (N_16831,N_14135,N_15683);
and U16832 (N_16832,N_15800,N_14343);
and U16833 (N_16833,N_15249,N_14565);
xor U16834 (N_16834,N_15093,N_15029);
and U16835 (N_16835,N_14239,N_15129);
and U16836 (N_16836,N_15685,N_14491);
xnor U16837 (N_16837,N_15379,N_15655);
or U16838 (N_16838,N_14561,N_14700);
xnor U16839 (N_16839,N_14460,N_14959);
or U16840 (N_16840,N_14754,N_15771);
and U16841 (N_16841,N_14697,N_15982);
nor U16842 (N_16842,N_14365,N_14525);
or U16843 (N_16843,N_14664,N_14947);
nand U16844 (N_16844,N_14461,N_15794);
or U16845 (N_16845,N_15645,N_15566);
nand U16846 (N_16846,N_14702,N_15237);
xor U16847 (N_16847,N_14989,N_14620);
and U16848 (N_16848,N_14414,N_14431);
xnor U16849 (N_16849,N_14457,N_15255);
xnor U16850 (N_16850,N_14511,N_15745);
nand U16851 (N_16851,N_15425,N_14548);
or U16852 (N_16852,N_15638,N_15325);
nand U16853 (N_16853,N_15916,N_14312);
or U16854 (N_16854,N_14148,N_14400);
and U16855 (N_16855,N_15340,N_15583);
xnor U16856 (N_16856,N_14006,N_14181);
or U16857 (N_16857,N_15200,N_15278);
nor U16858 (N_16858,N_14013,N_15423);
or U16859 (N_16859,N_14762,N_15179);
or U16860 (N_16860,N_14761,N_15056);
nand U16861 (N_16861,N_15857,N_15111);
and U16862 (N_16862,N_14070,N_14074);
xnor U16863 (N_16863,N_14883,N_14916);
nand U16864 (N_16864,N_15862,N_14912);
nand U16865 (N_16865,N_14985,N_15038);
xnor U16866 (N_16866,N_14435,N_15202);
xor U16867 (N_16867,N_14714,N_15710);
and U16868 (N_16868,N_14184,N_14872);
or U16869 (N_16869,N_14456,N_15021);
nand U16870 (N_16870,N_15875,N_14683);
nand U16871 (N_16871,N_14276,N_15495);
and U16872 (N_16872,N_15481,N_14920);
xor U16873 (N_16873,N_15295,N_15821);
and U16874 (N_16874,N_15281,N_15884);
xor U16875 (N_16875,N_14737,N_14109);
and U16876 (N_16876,N_14356,N_14136);
nand U16877 (N_16877,N_14361,N_15490);
xnor U16878 (N_16878,N_14026,N_14854);
nand U16879 (N_16879,N_14338,N_15839);
nand U16880 (N_16880,N_14193,N_14366);
xor U16881 (N_16881,N_15082,N_15508);
nor U16882 (N_16882,N_15363,N_14325);
nand U16883 (N_16883,N_14368,N_15362);
nor U16884 (N_16884,N_14843,N_14049);
and U16885 (N_16885,N_15477,N_14574);
and U16886 (N_16886,N_15613,N_15617);
and U16887 (N_16887,N_14283,N_15878);
xnor U16888 (N_16888,N_14203,N_15078);
and U16889 (N_16889,N_14826,N_15761);
nand U16890 (N_16890,N_15103,N_15718);
and U16891 (N_16891,N_15168,N_14166);
xnor U16892 (N_16892,N_14382,N_15906);
and U16893 (N_16893,N_15576,N_14905);
xnor U16894 (N_16894,N_15577,N_14307);
nand U16895 (N_16895,N_14529,N_15073);
or U16896 (N_16896,N_15498,N_15333);
nand U16897 (N_16897,N_14818,N_14294);
or U16898 (N_16898,N_14909,N_14012);
or U16899 (N_16899,N_14332,N_14324);
or U16900 (N_16900,N_14600,N_15891);
nor U16901 (N_16901,N_15366,N_15892);
or U16902 (N_16902,N_15374,N_14470);
nor U16903 (N_16903,N_15633,N_15392);
nor U16904 (N_16904,N_14483,N_14237);
and U16905 (N_16905,N_14889,N_14517);
nor U16906 (N_16906,N_15947,N_15377);
nand U16907 (N_16907,N_15071,N_15006);
xnor U16908 (N_16908,N_15772,N_15806);
nand U16909 (N_16909,N_15351,N_14966);
nand U16910 (N_16910,N_14898,N_15675);
xor U16911 (N_16911,N_15537,N_15983);
or U16912 (N_16912,N_15861,N_14679);
and U16913 (N_16913,N_14131,N_15588);
or U16914 (N_16914,N_14879,N_15109);
and U16915 (N_16915,N_14887,N_14913);
xnor U16916 (N_16916,N_15160,N_15601);
nor U16917 (N_16917,N_14692,N_15499);
or U16918 (N_16918,N_14657,N_14211);
or U16919 (N_16919,N_15450,N_14110);
or U16920 (N_16920,N_14494,N_14467);
or U16921 (N_16921,N_14741,N_14925);
and U16922 (N_16922,N_14688,N_15000);
xnor U16923 (N_16923,N_15186,N_14020);
nand U16924 (N_16924,N_14217,N_14403);
nand U16925 (N_16925,N_15624,N_14665);
nand U16926 (N_16926,N_15783,N_15003);
nor U16927 (N_16927,N_14690,N_14263);
nand U16928 (N_16928,N_15563,N_14710);
nor U16929 (N_16929,N_14896,N_14685);
xor U16930 (N_16930,N_15643,N_14253);
xnor U16931 (N_16931,N_15923,N_15873);
or U16932 (N_16932,N_14373,N_15557);
nor U16933 (N_16933,N_15319,N_15804);
or U16934 (N_16934,N_14279,N_14280);
and U16935 (N_16935,N_15330,N_14047);
xnor U16936 (N_16936,N_14567,N_15190);
and U16937 (N_16937,N_15899,N_15206);
nand U16938 (N_16938,N_14086,N_14028);
nand U16939 (N_16939,N_15276,N_14791);
nand U16940 (N_16940,N_15265,N_15283);
nand U16941 (N_16941,N_14357,N_15163);
xor U16942 (N_16942,N_14281,N_14694);
xnor U16943 (N_16943,N_15047,N_14933);
xnor U16944 (N_16944,N_14871,N_15214);
xor U16945 (N_16945,N_15699,N_14835);
or U16946 (N_16946,N_14666,N_15170);
and U16947 (N_16947,N_15765,N_15120);
and U16948 (N_16948,N_15282,N_14010);
and U16949 (N_16949,N_14106,N_14834);
nor U16950 (N_16950,N_15797,N_14405);
xnor U16951 (N_16951,N_15409,N_15383);
xnor U16952 (N_16952,N_15704,N_15847);
nand U16953 (N_16953,N_15727,N_15637);
nand U16954 (N_16954,N_14893,N_14520);
nand U16955 (N_16955,N_15634,N_14268);
and U16956 (N_16956,N_15115,N_15695);
nor U16957 (N_16957,N_15998,N_14311);
or U16958 (N_16958,N_14011,N_14783);
nand U16959 (N_16959,N_15622,N_14534);
or U16960 (N_16960,N_15831,N_15709);
xnor U16961 (N_16961,N_15962,N_14850);
nor U16962 (N_16962,N_14495,N_14987);
or U16963 (N_16963,N_15277,N_14321);
and U16964 (N_16964,N_15421,N_15145);
nand U16965 (N_16965,N_14647,N_14024);
or U16966 (N_16966,N_14264,N_15625);
and U16967 (N_16967,N_14588,N_15653);
nor U16968 (N_16968,N_14934,N_14030);
and U16969 (N_16969,N_15616,N_15833);
nand U16970 (N_16970,N_14978,N_14863);
nor U16971 (N_16971,N_14067,N_15086);
nand U16972 (N_16972,N_15610,N_15441);
nor U16973 (N_16973,N_14875,N_15665);
nor U16974 (N_16974,N_15311,N_14864);
nor U16975 (N_16975,N_15558,N_14625);
xor U16976 (N_16976,N_15750,N_14578);
and U16977 (N_16977,N_15614,N_14092);
or U16978 (N_16978,N_15945,N_15309);
and U16979 (N_16979,N_14655,N_14908);
and U16980 (N_16980,N_14954,N_15943);
and U16981 (N_16981,N_15460,N_14051);
xor U16982 (N_16982,N_14046,N_14550);
xnor U16983 (N_16983,N_15788,N_15487);
and U16984 (N_16984,N_14341,N_15834);
nor U16985 (N_16985,N_15100,N_14336);
and U16986 (N_16986,N_15228,N_15218);
nor U16987 (N_16987,N_15756,N_14058);
and U16988 (N_16988,N_14833,N_14530);
nand U16989 (N_16989,N_15781,N_15594);
xor U16990 (N_16990,N_15352,N_14719);
nor U16991 (N_16991,N_15432,N_15239);
nand U16992 (N_16992,N_14789,N_14422);
and U16993 (N_16993,N_14884,N_14375);
xnor U16994 (N_16994,N_14125,N_15212);
nand U16995 (N_16995,N_15805,N_14285);
or U16996 (N_16996,N_15169,N_15525);
xor U16997 (N_16997,N_14358,N_14300);
or U16998 (N_16998,N_14043,N_14773);
nor U16999 (N_16999,N_14419,N_15248);
or U17000 (N_17000,N_15136,N_14963);
xnor U17001 (N_17001,N_15903,N_14238);
or U17002 (N_17002,N_15772,N_15521);
or U17003 (N_17003,N_15908,N_14531);
xor U17004 (N_17004,N_14512,N_15023);
or U17005 (N_17005,N_15463,N_15199);
or U17006 (N_17006,N_15554,N_15244);
xnor U17007 (N_17007,N_15384,N_15174);
nor U17008 (N_17008,N_14371,N_14341);
xor U17009 (N_17009,N_14250,N_14040);
xor U17010 (N_17010,N_14384,N_14521);
xor U17011 (N_17011,N_15113,N_15169);
nand U17012 (N_17012,N_15496,N_14314);
nand U17013 (N_17013,N_14548,N_15004);
nor U17014 (N_17014,N_15069,N_14442);
xor U17015 (N_17015,N_15502,N_14857);
nand U17016 (N_17016,N_15012,N_14561);
and U17017 (N_17017,N_14265,N_14888);
nand U17018 (N_17018,N_14703,N_15008);
xor U17019 (N_17019,N_14537,N_14879);
and U17020 (N_17020,N_14268,N_15998);
nor U17021 (N_17021,N_14846,N_15110);
nand U17022 (N_17022,N_14409,N_14063);
and U17023 (N_17023,N_14561,N_15806);
nand U17024 (N_17024,N_14409,N_15043);
xor U17025 (N_17025,N_14304,N_14869);
nand U17026 (N_17026,N_15154,N_15101);
nor U17027 (N_17027,N_15871,N_15755);
or U17028 (N_17028,N_14365,N_15699);
xor U17029 (N_17029,N_14973,N_14996);
or U17030 (N_17030,N_14232,N_14103);
xnor U17031 (N_17031,N_15754,N_14000);
and U17032 (N_17032,N_14203,N_14294);
or U17033 (N_17033,N_15513,N_15780);
xor U17034 (N_17034,N_14549,N_15832);
and U17035 (N_17035,N_15676,N_15152);
nand U17036 (N_17036,N_14468,N_15579);
xnor U17037 (N_17037,N_14492,N_15571);
or U17038 (N_17038,N_15789,N_15900);
xor U17039 (N_17039,N_14979,N_15551);
nor U17040 (N_17040,N_15178,N_15972);
xor U17041 (N_17041,N_14244,N_14575);
and U17042 (N_17042,N_14587,N_15740);
nor U17043 (N_17043,N_15315,N_15962);
nand U17044 (N_17044,N_14130,N_14184);
nor U17045 (N_17045,N_14474,N_15428);
and U17046 (N_17046,N_15877,N_14229);
or U17047 (N_17047,N_14531,N_15634);
xnor U17048 (N_17048,N_15695,N_14541);
or U17049 (N_17049,N_15543,N_15837);
nor U17050 (N_17050,N_14418,N_15775);
nand U17051 (N_17051,N_15622,N_15233);
nor U17052 (N_17052,N_14888,N_14561);
nand U17053 (N_17053,N_15549,N_14594);
xor U17054 (N_17054,N_14499,N_15600);
xnor U17055 (N_17055,N_14104,N_14445);
nand U17056 (N_17056,N_15779,N_15802);
nand U17057 (N_17057,N_14510,N_14078);
nor U17058 (N_17058,N_14012,N_15626);
xor U17059 (N_17059,N_14577,N_15476);
and U17060 (N_17060,N_15822,N_14167);
xnor U17061 (N_17061,N_14595,N_14755);
and U17062 (N_17062,N_15522,N_14100);
and U17063 (N_17063,N_15259,N_15174);
nand U17064 (N_17064,N_15858,N_15576);
nand U17065 (N_17065,N_14664,N_15568);
nor U17066 (N_17066,N_15941,N_15011);
or U17067 (N_17067,N_14548,N_14946);
xor U17068 (N_17068,N_15316,N_15357);
nand U17069 (N_17069,N_15471,N_15969);
or U17070 (N_17070,N_15565,N_15869);
xor U17071 (N_17071,N_15656,N_14094);
xor U17072 (N_17072,N_14165,N_14376);
nor U17073 (N_17073,N_15217,N_14847);
xnor U17074 (N_17074,N_15069,N_14426);
and U17075 (N_17075,N_15932,N_14749);
or U17076 (N_17076,N_15653,N_15873);
nor U17077 (N_17077,N_14969,N_15750);
xor U17078 (N_17078,N_14781,N_15168);
nor U17079 (N_17079,N_15776,N_14015);
or U17080 (N_17080,N_15444,N_15714);
and U17081 (N_17081,N_14575,N_14799);
nor U17082 (N_17082,N_14657,N_15856);
and U17083 (N_17083,N_15911,N_14090);
nand U17084 (N_17084,N_14793,N_15419);
nand U17085 (N_17085,N_15943,N_15018);
xnor U17086 (N_17086,N_15715,N_14927);
xnor U17087 (N_17087,N_14918,N_15064);
or U17088 (N_17088,N_15390,N_15757);
nand U17089 (N_17089,N_15704,N_15690);
or U17090 (N_17090,N_14211,N_14671);
or U17091 (N_17091,N_15622,N_14350);
and U17092 (N_17092,N_15056,N_15139);
nor U17093 (N_17093,N_14035,N_14659);
and U17094 (N_17094,N_14933,N_15576);
or U17095 (N_17095,N_14901,N_15403);
and U17096 (N_17096,N_14048,N_15879);
and U17097 (N_17097,N_15029,N_15521);
or U17098 (N_17098,N_14141,N_15659);
nand U17099 (N_17099,N_15370,N_15803);
or U17100 (N_17100,N_14723,N_14463);
xnor U17101 (N_17101,N_15857,N_15123);
xnor U17102 (N_17102,N_14647,N_14151);
or U17103 (N_17103,N_14902,N_14184);
and U17104 (N_17104,N_14153,N_15817);
or U17105 (N_17105,N_15383,N_14763);
or U17106 (N_17106,N_14441,N_14125);
and U17107 (N_17107,N_14260,N_15184);
or U17108 (N_17108,N_15250,N_15285);
nand U17109 (N_17109,N_15044,N_14061);
xnor U17110 (N_17110,N_14313,N_14493);
xnor U17111 (N_17111,N_14727,N_14859);
xnor U17112 (N_17112,N_14341,N_15891);
nor U17113 (N_17113,N_15829,N_15726);
or U17114 (N_17114,N_14499,N_15789);
nand U17115 (N_17115,N_14936,N_14639);
or U17116 (N_17116,N_14597,N_14339);
and U17117 (N_17117,N_14144,N_14637);
nand U17118 (N_17118,N_14438,N_15577);
or U17119 (N_17119,N_15803,N_14052);
xnor U17120 (N_17120,N_15211,N_15644);
nand U17121 (N_17121,N_15590,N_15023);
nand U17122 (N_17122,N_15634,N_14351);
nor U17123 (N_17123,N_15948,N_15120);
nor U17124 (N_17124,N_14326,N_14586);
and U17125 (N_17125,N_15159,N_14326);
xnor U17126 (N_17126,N_14936,N_14384);
or U17127 (N_17127,N_14583,N_15983);
nor U17128 (N_17128,N_14588,N_14942);
xnor U17129 (N_17129,N_15100,N_15866);
and U17130 (N_17130,N_14534,N_14539);
xor U17131 (N_17131,N_14705,N_15091);
nor U17132 (N_17132,N_15387,N_15656);
nand U17133 (N_17133,N_15330,N_14920);
xor U17134 (N_17134,N_14776,N_15655);
and U17135 (N_17135,N_14546,N_15264);
or U17136 (N_17136,N_14902,N_15281);
nand U17137 (N_17137,N_15154,N_15362);
or U17138 (N_17138,N_14035,N_14573);
nor U17139 (N_17139,N_14440,N_15828);
and U17140 (N_17140,N_15725,N_14476);
nor U17141 (N_17141,N_14547,N_14707);
nand U17142 (N_17142,N_15154,N_15848);
xor U17143 (N_17143,N_15260,N_14410);
nand U17144 (N_17144,N_14062,N_14212);
nand U17145 (N_17145,N_15686,N_14421);
nor U17146 (N_17146,N_14755,N_14032);
nor U17147 (N_17147,N_14322,N_15023);
nand U17148 (N_17148,N_15164,N_15506);
nand U17149 (N_17149,N_14582,N_15688);
nor U17150 (N_17150,N_14907,N_15869);
xnor U17151 (N_17151,N_15923,N_14223);
and U17152 (N_17152,N_14723,N_14318);
xnor U17153 (N_17153,N_14914,N_14693);
xor U17154 (N_17154,N_14407,N_14571);
nor U17155 (N_17155,N_15554,N_15310);
xor U17156 (N_17156,N_14123,N_14889);
xor U17157 (N_17157,N_15530,N_15654);
nor U17158 (N_17158,N_14083,N_14274);
and U17159 (N_17159,N_14791,N_14643);
nor U17160 (N_17160,N_14166,N_14684);
xnor U17161 (N_17161,N_14925,N_14060);
nor U17162 (N_17162,N_15685,N_14573);
and U17163 (N_17163,N_14741,N_14400);
xor U17164 (N_17164,N_14640,N_14753);
and U17165 (N_17165,N_15355,N_15638);
or U17166 (N_17166,N_14617,N_14630);
and U17167 (N_17167,N_14953,N_15404);
xnor U17168 (N_17168,N_14248,N_15837);
nor U17169 (N_17169,N_14786,N_15579);
xor U17170 (N_17170,N_15101,N_15487);
nand U17171 (N_17171,N_15044,N_15515);
and U17172 (N_17172,N_15582,N_14895);
nor U17173 (N_17173,N_15644,N_15635);
and U17174 (N_17174,N_14945,N_15564);
and U17175 (N_17175,N_15031,N_15386);
nand U17176 (N_17176,N_15526,N_14302);
and U17177 (N_17177,N_15102,N_15145);
xnor U17178 (N_17178,N_14685,N_15733);
nand U17179 (N_17179,N_15257,N_14754);
nand U17180 (N_17180,N_15158,N_14571);
nor U17181 (N_17181,N_14932,N_15303);
xor U17182 (N_17182,N_14958,N_14231);
and U17183 (N_17183,N_15952,N_14602);
nand U17184 (N_17184,N_14831,N_14933);
xnor U17185 (N_17185,N_15260,N_14857);
and U17186 (N_17186,N_14032,N_15875);
nand U17187 (N_17187,N_14003,N_15282);
nor U17188 (N_17188,N_15856,N_15655);
or U17189 (N_17189,N_14734,N_14210);
nand U17190 (N_17190,N_14085,N_15570);
nand U17191 (N_17191,N_15290,N_15357);
and U17192 (N_17192,N_14165,N_14606);
nand U17193 (N_17193,N_15850,N_15817);
xnor U17194 (N_17194,N_15860,N_15044);
and U17195 (N_17195,N_15107,N_14326);
nor U17196 (N_17196,N_15620,N_14957);
xnor U17197 (N_17197,N_14057,N_14766);
xnor U17198 (N_17198,N_15537,N_15372);
or U17199 (N_17199,N_15486,N_15350);
nor U17200 (N_17200,N_15742,N_15024);
nor U17201 (N_17201,N_15595,N_14331);
xnor U17202 (N_17202,N_14562,N_15973);
nand U17203 (N_17203,N_14964,N_14606);
nor U17204 (N_17204,N_15346,N_14539);
or U17205 (N_17205,N_14969,N_14721);
and U17206 (N_17206,N_14903,N_14642);
or U17207 (N_17207,N_14924,N_15489);
or U17208 (N_17208,N_14086,N_15747);
nor U17209 (N_17209,N_15052,N_14363);
xor U17210 (N_17210,N_14173,N_15489);
or U17211 (N_17211,N_14017,N_15543);
and U17212 (N_17212,N_14661,N_14200);
xnor U17213 (N_17213,N_15398,N_15707);
nand U17214 (N_17214,N_15623,N_14708);
nor U17215 (N_17215,N_15850,N_14856);
and U17216 (N_17216,N_14500,N_15850);
xnor U17217 (N_17217,N_15433,N_14391);
or U17218 (N_17218,N_14674,N_14730);
nor U17219 (N_17219,N_14471,N_14260);
or U17220 (N_17220,N_15262,N_15736);
and U17221 (N_17221,N_15198,N_14006);
and U17222 (N_17222,N_15755,N_14629);
or U17223 (N_17223,N_15165,N_15188);
xor U17224 (N_17224,N_15627,N_15361);
and U17225 (N_17225,N_14566,N_14642);
and U17226 (N_17226,N_15201,N_14181);
and U17227 (N_17227,N_14506,N_15903);
and U17228 (N_17228,N_15038,N_14363);
or U17229 (N_17229,N_15751,N_15966);
or U17230 (N_17230,N_14010,N_15379);
nor U17231 (N_17231,N_15148,N_15196);
nand U17232 (N_17232,N_15087,N_15697);
and U17233 (N_17233,N_15395,N_15401);
nand U17234 (N_17234,N_15949,N_15462);
or U17235 (N_17235,N_15712,N_14285);
or U17236 (N_17236,N_14073,N_15786);
nor U17237 (N_17237,N_15252,N_14819);
nand U17238 (N_17238,N_14443,N_14174);
or U17239 (N_17239,N_14185,N_15186);
or U17240 (N_17240,N_15897,N_15908);
nand U17241 (N_17241,N_15443,N_14830);
nor U17242 (N_17242,N_15170,N_15865);
or U17243 (N_17243,N_15261,N_15739);
and U17244 (N_17244,N_15285,N_14827);
and U17245 (N_17245,N_15730,N_15231);
or U17246 (N_17246,N_15693,N_15466);
or U17247 (N_17247,N_14105,N_14359);
nand U17248 (N_17248,N_15926,N_15634);
and U17249 (N_17249,N_14589,N_14301);
nand U17250 (N_17250,N_15500,N_15869);
nor U17251 (N_17251,N_15598,N_14363);
xnor U17252 (N_17252,N_14232,N_15468);
or U17253 (N_17253,N_14881,N_14266);
and U17254 (N_17254,N_15259,N_15273);
xnor U17255 (N_17255,N_14723,N_15186);
xor U17256 (N_17256,N_15051,N_15076);
or U17257 (N_17257,N_14181,N_14908);
or U17258 (N_17258,N_14496,N_15452);
or U17259 (N_17259,N_15224,N_15058);
or U17260 (N_17260,N_15250,N_14389);
nand U17261 (N_17261,N_14729,N_14778);
nand U17262 (N_17262,N_15153,N_15782);
or U17263 (N_17263,N_14488,N_14638);
or U17264 (N_17264,N_14638,N_14228);
or U17265 (N_17265,N_15742,N_15827);
and U17266 (N_17266,N_14134,N_14289);
or U17267 (N_17267,N_14128,N_14775);
and U17268 (N_17268,N_14625,N_15769);
nor U17269 (N_17269,N_15946,N_15241);
nor U17270 (N_17270,N_15902,N_14450);
nor U17271 (N_17271,N_14433,N_15630);
or U17272 (N_17272,N_15221,N_14325);
and U17273 (N_17273,N_14619,N_15905);
or U17274 (N_17274,N_15473,N_14908);
and U17275 (N_17275,N_14991,N_15074);
nor U17276 (N_17276,N_14094,N_14687);
nand U17277 (N_17277,N_14689,N_14775);
nor U17278 (N_17278,N_14309,N_14303);
nand U17279 (N_17279,N_14331,N_15494);
nor U17280 (N_17280,N_14359,N_14838);
nor U17281 (N_17281,N_15421,N_15375);
xor U17282 (N_17282,N_15108,N_14308);
and U17283 (N_17283,N_14833,N_15753);
nor U17284 (N_17284,N_14316,N_14044);
or U17285 (N_17285,N_14445,N_14717);
xor U17286 (N_17286,N_14034,N_14346);
xnor U17287 (N_17287,N_14265,N_15178);
or U17288 (N_17288,N_15684,N_14477);
or U17289 (N_17289,N_14565,N_15547);
nor U17290 (N_17290,N_14769,N_15429);
and U17291 (N_17291,N_15582,N_15280);
nand U17292 (N_17292,N_14762,N_15965);
or U17293 (N_17293,N_15175,N_15186);
and U17294 (N_17294,N_14156,N_15191);
or U17295 (N_17295,N_14783,N_14501);
xor U17296 (N_17296,N_14071,N_15647);
nor U17297 (N_17297,N_14672,N_14033);
and U17298 (N_17298,N_14964,N_14157);
xor U17299 (N_17299,N_14497,N_14938);
or U17300 (N_17300,N_15580,N_15490);
nand U17301 (N_17301,N_14632,N_14810);
xor U17302 (N_17302,N_14053,N_15018);
or U17303 (N_17303,N_15819,N_15732);
xnor U17304 (N_17304,N_14231,N_14608);
and U17305 (N_17305,N_15749,N_15654);
and U17306 (N_17306,N_14214,N_15649);
xnor U17307 (N_17307,N_15825,N_15012);
and U17308 (N_17308,N_14838,N_15451);
and U17309 (N_17309,N_15111,N_14681);
or U17310 (N_17310,N_14035,N_15152);
nand U17311 (N_17311,N_15013,N_14028);
xnor U17312 (N_17312,N_15931,N_15032);
nand U17313 (N_17313,N_15605,N_15644);
nor U17314 (N_17314,N_14448,N_15163);
xor U17315 (N_17315,N_14616,N_14357);
nand U17316 (N_17316,N_15320,N_15032);
nand U17317 (N_17317,N_15370,N_14881);
nor U17318 (N_17318,N_15792,N_15072);
nand U17319 (N_17319,N_15258,N_14778);
or U17320 (N_17320,N_15411,N_14372);
nand U17321 (N_17321,N_15860,N_14199);
and U17322 (N_17322,N_15111,N_15928);
nor U17323 (N_17323,N_14071,N_15732);
xor U17324 (N_17324,N_14220,N_15524);
nand U17325 (N_17325,N_15012,N_14068);
and U17326 (N_17326,N_14634,N_15681);
xor U17327 (N_17327,N_15518,N_14869);
or U17328 (N_17328,N_14519,N_15910);
nand U17329 (N_17329,N_15507,N_15100);
xnor U17330 (N_17330,N_14564,N_15039);
nand U17331 (N_17331,N_15146,N_15819);
or U17332 (N_17332,N_15739,N_15049);
xor U17333 (N_17333,N_14824,N_14328);
xor U17334 (N_17334,N_15998,N_14404);
xor U17335 (N_17335,N_15430,N_14363);
nor U17336 (N_17336,N_15465,N_14513);
or U17337 (N_17337,N_14677,N_15260);
nor U17338 (N_17338,N_15655,N_15695);
and U17339 (N_17339,N_15018,N_15738);
and U17340 (N_17340,N_15358,N_14660);
and U17341 (N_17341,N_15687,N_15930);
nand U17342 (N_17342,N_14767,N_15547);
nor U17343 (N_17343,N_15465,N_14581);
nand U17344 (N_17344,N_14949,N_14548);
or U17345 (N_17345,N_14763,N_15126);
or U17346 (N_17346,N_14861,N_14766);
nor U17347 (N_17347,N_15800,N_14407);
nor U17348 (N_17348,N_15056,N_14532);
xor U17349 (N_17349,N_14530,N_14353);
or U17350 (N_17350,N_14001,N_15646);
or U17351 (N_17351,N_14269,N_14898);
nand U17352 (N_17352,N_15631,N_15943);
xor U17353 (N_17353,N_14980,N_14153);
xnor U17354 (N_17354,N_15410,N_14540);
nor U17355 (N_17355,N_15591,N_14716);
or U17356 (N_17356,N_15048,N_14727);
or U17357 (N_17357,N_15685,N_15866);
xor U17358 (N_17358,N_15236,N_15336);
nand U17359 (N_17359,N_14799,N_15377);
or U17360 (N_17360,N_14452,N_15395);
nand U17361 (N_17361,N_15713,N_15148);
xor U17362 (N_17362,N_14060,N_14464);
nand U17363 (N_17363,N_14798,N_14485);
or U17364 (N_17364,N_14063,N_15832);
or U17365 (N_17365,N_14614,N_15555);
or U17366 (N_17366,N_14251,N_14246);
xor U17367 (N_17367,N_14201,N_14355);
xor U17368 (N_17368,N_14763,N_14411);
xor U17369 (N_17369,N_15286,N_15042);
nor U17370 (N_17370,N_15973,N_15884);
and U17371 (N_17371,N_15507,N_15647);
xnor U17372 (N_17372,N_14538,N_14003);
and U17373 (N_17373,N_14871,N_15593);
xor U17374 (N_17374,N_14778,N_15936);
nor U17375 (N_17375,N_14532,N_15850);
nand U17376 (N_17376,N_14523,N_15643);
xor U17377 (N_17377,N_15735,N_15625);
or U17378 (N_17378,N_14336,N_15833);
nor U17379 (N_17379,N_14587,N_15820);
and U17380 (N_17380,N_15596,N_14212);
nor U17381 (N_17381,N_14912,N_14962);
and U17382 (N_17382,N_15559,N_15271);
or U17383 (N_17383,N_15530,N_15531);
xnor U17384 (N_17384,N_15655,N_14464);
xor U17385 (N_17385,N_15597,N_15164);
nor U17386 (N_17386,N_15065,N_15465);
xor U17387 (N_17387,N_15681,N_15922);
or U17388 (N_17388,N_15450,N_14048);
and U17389 (N_17389,N_14824,N_15646);
and U17390 (N_17390,N_14035,N_14118);
or U17391 (N_17391,N_14850,N_14834);
or U17392 (N_17392,N_14668,N_15994);
nor U17393 (N_17393,N_14336,N_15857);
or U17394 (N_17394,N_15105,N_15119);
xor U17395 (N_17395,N_14173,N_14052);
or U17396 (N_17396,N_15264,N_15159);
nor U17397 (N_17397,N_14256,N_15420);
xnor U17398 (N_17398,N_14219,N_15450);
or U17399 (N_17399,N_15533,N_15624);
nand U17400 (N_17400,N_15314,N_15242);
xnor U17401 (N_17401,N_15844,N_15406);
and U17402 (N_17402,N_14580,N_15239);
and U17403 (N_17403,N_14770,N_15174);
or U17404 (N_17404,N_14283,N_14875);
and U17405 (N_17405,N_15699,N_14373);
nand U17406 (N_17406,N_15418,N_14110);
and U17407 (N_17407,N_14735,N_15169);
nand U17408 (N_17408,N_14048,N_15946);
nand U17409 (N_17409,N_15070,N_14763);
nor U17410 (N_17410,N_15948,N_15957);
xor U17411 (N_17411,N_14214,N_15459);
nor U17412 (N_17412,N_15470,N_15502);
or U17413 (N_17413,N_15117,N_15860);
and U17414 (N_17414,N_15056,N_14440);
xor U17415 (N_17415,N_15421,N_14832);
xor U17416 (N_17416,N_15123,N_14128);
nand U17417 (N_17417,N_14109,N_14019);
nand U17418 (N_17418,N_15728,N_14059);
or U17419 (N_17419,N_15027,N_15238);
and U17420 (N_17420,N_15069,N_15060);
nand U17421 (N_17421,N_15965,N_15634);
nand U17422 (N_17422,N_15255,N_14289);
and U17423 (N_17423,N_14635,N_15528);
and U17424 (N_17424,N_14317,N_14660);
or U17425 (N_17425,N_14053,N_14035);
or U17426 (N_17426,N_14000,N_14293);
xnor U17427 (N_17427,N_15952,N_15415);
nand U17428 (N_17428,N_14483,N_15284);
nor U17429 (N_17429,N_15189,N_14563);
nand U17430 (N_17430,N_15519,N_15359);
nand U17431 (N_17431,N_14787,N_15955);
nor U17432 (N_17432,N_14049,N_14741);
xor U17433 (N_17433,N_14675,N_15812);
or U17434 (N_17434,N_15800,N_15148);
or U17435 (N_17435,N_15422,N_14830);
or U17436 (N_17436,N_14519,N_15133);
nand U17437 (N_17437,N_14324,N_14667);
xnor U17438 (N_17438,N_14235,N_15228);
nand U17439 (N_17439,N_14609,N_14248);
and U17440 (N_17440,N_14696,N_15673);
nor U17441 (N_17441,N_14775,N_15253);
nor U17442 (N_17442,N_14024,N_14442);
nand U17443 (N_17443,N_15423,N_15201);
and U17444 (N_17444,N_15520,N_15005);
nand U17445 (N_17445,N_14112,N_14516);
or U17446 (N_17446,N_15408,N_14605);
xor U17447 (N_17447,N_14424,N_15004);
or U17448 (N_17448,N_14193,N_14246);
nand U17449 (N_17449,N_15644,N_15705);
nand U17450 (N_17450,N_14090,N_14481);
or U17451 (N_17451,N_14926,N_14227);
and U17452 (N_17452,N_14750,N_15744);
xor U17453 (N_17453,N_15974,N_15601);
and U17454 (N_17454,N_15819,N_14479);
xor U17455 (N_17455,N_15286,N_14219);
xor U17456 (N_17456,N_14453,N_15028);
xor U17457 (N_17457,N_15302,N_15696);
xnor U17458 (N_17458,N_14311,N_14640);
or U17459 (N_17459,N_14382,N_15214);
and U17460 (N_17460,N_15373,N_14170);
or U17461 (N_17461,N_15271,N_15768);
xnor U17462 (N_17462,N_15142,N_15856);
or U17463 (N_17463,N_15977,N_14128);
nor U17464 (N_17464,N_14050,N_14018);
xor U17465 (N_17465,N_15119,N_14665);
and U17466 (N_17466,N_15648,N_15038);
nor U17467 (N_17467,N_15244,N_15906);
xnor U17468 (N_17468,N_14829,N_14802);
or U17469 (N_17469,N_14380,N_14770);
nand U17470 (N_17470,N_14977,N_15488);
and U17471 (N_17471,N_14896,N_14479);
nand U17472 (N_17472,N_14437,N_15578);
and U17473 (N_17473,N_15057,N_15377);
xor U17474 (N_17474,N_14029,N_15350);
and U17475 (N_17475,N_15952,N_15032);
or U17476 (N_17476,N_14360,N_14868);
nand U17477 (N_17477,N_14220,N_15268);
nor U17478 (N_17478,N_14331,N_15760);
or U17479 (N_17479,N_15264,N_15145);
nand U17480 (N_17480,N_15975,N_14239);
nand U17481 (N_17481,N_14741,N_14574);
xor U17482 (N_17482,N_14230,N_15958);
and U17483 (N_17483,N_15866,N_15509);
xor U17484 (N_17484,N_15010,N_15926);
and U17485 (N_17485,N_14596,N_14851);
or U17486 (N_17486,N_15773,N_14498);
and U17487 (N_17487,N_15599,N_15682);
xor U17488 (N_17488,N_15600,N_14621);
and U17489 (N_17489,N_15640,N_14686);
or U17490 (N_17490,N_15213,N_14005);
or U17491 (N_17491,N_15838,N_14676);
or U17492 (N_17492,N_15559,N_14030);
xnor U17493 (N_17493,N_14149,N_14308);
or U17494 (N_17494,N_15253,N_15656);
or U17495 (N_17495,N_15780,N_15932);
and U17496 (N_17496,N_15901,N_14877);
nor U17497 (N_17497,N_15420,N_15029);
nand U17498 (N_17498,N_15291,N_14353);
or U17499 (N_17499,N_14751,N_15350);
nand U17500 (N_17500,N_15978,N_14873);
xnor U17501 (N_17501,N_14722,N_14779);
nor U17502 (N_17502,N_15847,N_14770);
nor U17503 (N_17503,N_15227,N_14568);
nand U17504 (N_17504,N_15446,N_15223);
nor U17505 (N_17505,N_15377,N_15646);
nand U17506 (N_17506,N_14276,N_14466);
nand U17507 (N_17507,N_14597,N_15816);
and U17508 (N_17508,N_15102,N_14140);
and U17509 (N_17509,N_14754,N_14383);
or U17510 (N_17510,N_15249,N_15831);
xnor U17511 (N_17511,N_14753,N_14379);
xor U17512 (N_17512,N_15073,N_15173);
nand U17513 (N_17513,N_14615,N_15563);
xnor U17514 (N_17514,N_14752,N_14059);
nor U17515 (N_17515,N_15223,N_14977);
nand U17516 (N_17516,N_15210,N_15142);
nor U17517 (N_17517,N_14838,N_14852);
nor U17518 (N_17518,N_14090,N_15329);
and U17519 (N_17519,N_14145,N_15586);
nor U17520 (N_17520,N_15838,N_15317);
and U17521 (N_17521,N_15088,N_14076);
nor U17522 (N_17522,N_15320,N_15901);
nor U17523 (N_17523,N_15579,N_14460);
or U17524 (N_17524,N_15479,N_15624);
nand U17525 (N_17525,N_14864,N_15447);
nor U17526 (N_17526,N_15246,N_14181);
and U17527 (N_17527,N_15796,N_14611);
and U17528 (N_17528,N_15003,N_14369);
or U17529 (N_17529,N_14617,N_15179);
xor U17530 (N_17530,N_15408,N_14713);
and U17531 (N_17531,N_14597,N_14546);
and U17532 (N_17532,N_14278,N_14741);
nand U17533 (N_17533,N_15061,N_14267);
xor U17534 (N_17534,N_14506,N_14327);
nor U17535 (N_17535,N_14655,N_14001);
xnor U17536 (N_17536,N_14570,N_15679);
xnor U17537 (N_17537,N_14579,N_15654);
nand U17538 (N_17538,N_15090,N_15403);
xor U17539 (N_17539,N_15263,N_14175);
or U17540 (N_17540,N_14243,N_15102);
nor U17541 (N_17541,N_14141,N_15753);
and U17542 (N_17542,N_14867,N_14073);
and U17543 (N_17543,N_15469,N_14201);
nor U17544 (N_17544,N_14896,N_14329);
nor U17545 (N_17545,N_14937,N_15693);
or U17546 (N_17546,N_14961,N_15156);
xor U17547 (N_17547,N_15500,N_14577);
nand U17548 (N_17548,N_14700,N_14063);
or U17549 (N_17549,N_14442,N_14603);
or U17550 (N_17550,N_14251,N_14363);
or U17551 (N_17551,N_15010,N_15642);
nor U17552 (N_17552,N_14495,N_14654);
nand U17553 (N_17553,N_15462,N_15375);
nor U17554 (N_17554,N_15228,N_14877);
or U17555 (N_17555,N_15709,N_15660);
and U17556 (N_17556,N_15247,N_15195);
nor U17557 (N_17557,N_15517,N_15016);
nor U17558 (N_17558,N_14532,N_14625);
xnor U17559 (N_17559,N_14191,N_15472);
nor U17560 (N_17560,N_15433,N_15961);
nor U17561 (N_17561,N_14626,N_15550);
nor U17562 (N_17562,N_14198,N_14248);
nand U17563 (N_17563,N_15916,N_14273);
nand U17564 (N_17564,N_14406,N_14348);
or U17565 (N_17565,N_15287,N_15850);
or U17566 (N_17566,N_14331,N_15876);
xnor U17567 (N_17567,N_15277,N_14458);
and U17568 (N_17568,N_14137,N_15816);
and U17569 (N_17569,N_14320,N_15351);
and U17570 (N_17570,N_15953,N_15317);
and U17571 (N_17571,N_15397,N_14834);
nand U17572 (N_17572,N_14676,N_14068);
nor U17573 (N_17573,N_15053,N_15696);
or U17574 (N_17574,N_14435,N_15149);
or U17575 (N_17575,N_15896,N_14230);
and U17576 (N_17576,N_15347,N_15174);
xor U17577 (N_17577,N_14487,N_14264);
xor U17578 (N_17578,N_14866,N_14394);
or U17579 (N_17579,N_14154,N_14562);
or U17580 (N_17580,N_14745,N_14924);
nor U17581 (N_17581,N_14633,N_15137);
xor U17582 (N_17582,N_14097,N_14413);
nor U17583 (N_17583,N_14046,N_14133);
and U17584 (N_17584,N_15935,N_14840);
and U17585 (N_17585,N_15576,N_14690);
nor U17586 (N_17586,N_14629,N_15878);
xnor U17587 (N_17587,N_15052,N_14694);
nor U17588 (N_17588,N_15602,N_15366);
xor U17589 (N_17589,N_14816,N_14699);
and U17590 (N_17590,N_15304,N_14573);
nand U17591 (N_17591,N_14668,N_14808);
and U17592 (N_17592,N_14383,N_15346);
or U17593 (N_17593,N_15880,N_15352);
xor U17594 (N_17594,N_14620,N_14091);
and U17595 (N_17595,N_15352,N_14912);
nand U17596 (N_17596,N_14321,N_14399);
xnor U17597 (N_17597,N_14698,N_15993);
nand U17598 (N_17598,N_15676,N_14802);
nand U17599 (N_17599,N_14349,N_15708);
nand U17600 (N_17600,N_15838,N_15230);
xor U17601 (N_17601,N_14300,N_14364);
xnor U17602 (N_17602,N_14581,N_15921);
and U17603 (N_17603,N_14254,N_15581);
nand U17604 (N_17604,N_15404,N_14847);
nor U17605 (N_17605,N_14046,N_15348);
nor U17606 (N_17606,N_14807,N_15106);
and U17607 (N_17607,N_14771,N_14160);
and U17608 (N_17608,N_15366,N_14957);
nand U17609 (N_17609,N_14193,N_14471);
nand U17610 (N_17610,N_15239,N_14687);
or U17611 (N_17611,N_15704,N_14968);
and U17612 (N_17612,N_15261,N_15444);
nand U17613 (N_17613,N_14181,N_15755);
or U17614 (N_17614,N_14052,N_15025);
nor U17615 (N_17615,N_15575,N_14919);
nand U17616 (N_17616,N_15557,N_15649);
nand U17617 (N_17617,N_14207,N_14755);
xnor U17618 (N_17618,N_14023,N_14819);
and U17619 (N_17619,N_14840,N_14011);
nand U17620 (N_17620,N_14926,N_15162);
or U17621 (N_17621,N_14825,N_14453);
xnor U17622 (N_17622,N_14543,N_15604);
and U17623 (N_17623,N_15668,N_15651);
nand U17624 (N_17624,N_15324,N_15425);
nand U17625 (N_17625,N_15022,N_14506);
xnor U17626 (N_17626,N_14447,N_15352);
and U17627 (N_17627,N_15870,N_15924);
nor U17628 (N_17628,N_14567,N_14779);
xor U17629 (N_17629,N_15058,N_15408);
nand U17630 (N_17630,N_15290,N_14541);
and U17631 (N_17631,N_14723,N_14738);
xnor U17632 (N_17632,N_14733,N_15520);
xnor U17633 (N_17633,N_15382,N_14541);
or U17634 (N_17634,N_14047,N_15638);
nand U17635 (N_17635,N_14491,N_15474);
nand U17636 (N_17636,N_14907,N_14984);
xnor U17637 (N_17637,N_15733,N_14259);
xor U17638 (N_17638,N_14098,N_14360);
nand U17639 (N_17639,N_15700,N_14381);
and U17640 (N_17640,N_15884,N_15738);
nor U17641 (N_17641,N_14883,N_15499);
nor U17642 (N_17642,N_14755,N_14120);
xor U17643 (N_17643,N_14585,N_15234);
xor U17644 (N_17644,N_15417,N_14574);
xor U17645 (N_17645,N_14952,N_14323);
nor U17646 (N_17646,N_14831,N_14758);
nor U17647 (N_17647,N_15793,N_14836);
xnor U17648 (N_17648,N_15762,N_14021);
nand U17649 (N_17649,N_14868,N_14476);
nor U17650 (N_17650,N_14843,N_15636);
or U17651 (N_17651,N_14100,N_14551);
nor U17652 (N_17652,N_14631,N_14193);
nor U17653 (N_17653,N_14782,N_15125);
nand U17654 (N_17654,N_14075,N_15904);
nor U17655 (N_17655,N_14506,N_15665);
or U17656 (N_17656,N_14338,N_15834);
nor U17657 (N_17657,N_15163,N_14483);
or U17658 (N_17658,N_15561,N_15488);
nand U17659 (N_17659,N_14231,N_15515);
nand U17660 (N_17660,N_14859,N_15990);
or U17661 (N_17661,N_15316,N_14394);
or U17662 (N_17662,N_14899,N_14836);
or U17663 (N_17663,N_14362,N_14120);
and U17664 (N_17664,N_15616,N_14179);
and U17665 (N_17665,N_15210,N_14522);
or U17666 (N_17666,N_15957,N_15550);
xnor U17667 (N_17667,N_14340,N_15399);
nand U17668 (N_17668,N_14635,N_14956);
or U17669 (N_17669,N_14657,N_14431);
or U17670 (N_17670,N_14170,N_14187);
nor U17671 (N_17671,N_14429,N_15932);
nor U17672 (N_17672,N_14906,N_15865);
nor U17673 (N_17673,N_14891,N_15589);
xnor U17674 (N_17674,N_14301,N_14501);
nand U17675 (N_17675,N_14036,N_14627);
nand U17676 (N_17676,N_14897,N_14078);
and U17677 (N_17677,N_14421,N_14789);
nand U17678 (N_17678,N_14234,N_14660);
nand U17679 (N_17679,N_15113,N_14538);
or U17680 (N_17680,N_15230,N_15766);
or U17681 (N_17681,N_14407,N_14608);
nand U17682 (N_17682,N_15608,N_14691);
nor U17683 (N_17683,N_14808,N_15356);
nand U17684 (N_17684,N_14881,N_14334);
and U17685 (N_17685,N_15443,N_15806);
and U17686 (N_17686,N_14476,N_14301);
xor U17687 (N_17687,N_15073,N_14420);
nor U17688 (N_17688,N_15698,N_14556);
and U17689 (N_17689,N_14069,N_14034);
and U17690 (N_17690,N_14728,N_14223);
nor U17691 (N_17691,N_15939,N_14361);
nand U17692 (N_17692,N_15183,N_14861);
nand U17693 (N_17693,N_15604,N_15531);
xnor U17694 (N_17694,N_15795,N_15874);
and U17695 (N_17695,N_15944,N_14454);
or U17696 (N_17696,N_15916,N_14498);
and U17697 (N_17697,N_15723,N_14888);
xor U17698 (N_17698,N_14034,N_15543);
xor U17699 (N_17699,N_15301,N_15231);
nand U17700 (N_17700,N_15196,N_14426);
nand U17701 (N_17701,N_14650,N_14452);
xor U17702 (N_17702,N_14992,N_15783);
nor U17703 (N_17703,N_14829,N_15842);
nand U17704 (N_17704,N_15167,N_15473);
or U17705 (N_17705,N_15971,N_15396);
or U17706 (N_17706,N_14123,N_15047);
nand U17707 (N_17707,N_15800,N_15124);
nor U17708 (N_17708,N_15535,N_15740);
or U17709 (N_17709,N_15668,N_15882);
or U17710 (N_17710,N_14544,N_14432);
nor U17711 (N_17711,N_14956,N_15016);
nor U17712 (N_17712,N_15782,N_15711);
or U17713 (N_17713,N_14924,N_14016);
or U17714 (N_17714,N_14155,N_15500);
nand U17715 (N_17715,N_14823,N_15748);
xnor U17716 (N_17716,N_14066,N_15740);
and U17717 (N_17717,N_14648,N_15004);
nand U17718 (N_17718,N_14436,N_14970);
nand U17719 (N_17719,N_15233,N_15195);
or U17720 (N_17720,N_15722,N_14878);
or U17721 (N_17721,N_14216,N_15307);
and U17722 (N_17722,N_15815,N_15701);
or U17723 (N_17723,N_14898,N_15431);
nor U17724 (N_17724,N_15190,N_14473);
xnor U17725 (N_17725,N_14353,N_15476);
xor U17726 (N_17726,N_15794,N_14100);
or U17727 (N_17727,N_15942,N_14730);
nor U17728 (N_17728,N_14132,N_15333);
or U17729 (N_17729,N_14998,N_15447);
nor U17730 (N_17730,N_15595,N_15287);
nor U17731 (N_17731,N_15782,N_14384);
nand U17732 (N_17732,N_15336,N_14435);
or U17733 (N_17733,N_14714,N_15317);
nor U17734 (N_17734,N_15131,N_14059);
xor U17735 (N_17735,N_15461,N_14142);
nand U17736 (N_17736,N_15041,N_15064);
nor U17737 (N_17737,N_14325,N_14523);
and U17738 (N_17738,N_14506,N_15921);
xor U17739 (N_17739,N_14514,N_15071);
and U17740 (N_17740,N_14299,N_14287);
and U17741 (N_17741,N_14453,N_14431);
and U17742 (N_17742,N_14455,N_14615);
nand U17743 (N_17743,N_15724,N_14480);
xnor U17744 (N_17744,N_15543,N_15178);
xor U17745 (N_17745,N_14011,N_14778);
and U17746 (N_17746,N_15109,N_15043);
nand U17747 (N_17747,N_14209,N_14512);
nor U17748 (N_17748,N_14611,N_15970);
nor U17749 (N_17749,N_14598,N_14084);
and U17750 (N_17750,N_14394,N_15601);
nand U17751 (N_17751,N_14156,N_14258);
nand U17752 (N_17752,N_14305,N_15165);
nand U17753 (N_17753,N_15125,N_14485);
xor U17754 (N_17754,N_14657,N_15172);
and U17755 (N_17755,N_15626,N_15706);
nand U17756 (N_17756,N_14644,N_15092);
nor U17757 (N_17757,N_15769,N_15505);
and U17758 (N_17758,N_15142,N_15681);
xor U17759 (N_17759,N_15373,N_15235);
nor U17760 (N_17760,N_14706,N_14108);
and U17761 (N_17761,N_14816,N_15251);
nand U17762 (N_17762,N_15764,N_14553);
xor U17763 (N_17763,N_14967,N_14537);
or U17764 (N_17764,N_15307,N_15084);
nand U17765 (N_17765,N_14396,N_15462);
nor U17766 (N_17766,N_14208,N_14175);
or U17767 (N_17767,N_15936,N_14162);
nand U17768 (N_17768,N_14772,N_15681);
or U17769 (N_17769,N_15274,N_14197);
xor U17770 (N_17770,N_14773,N_14754);
nand U17771 (N_17771,N_15801,N_15130);
nand U17772 (N_17772,N_15276,N_14953);
nand U17773 (N_17773,N_14203,N_14288);
nor U17774 (N_17774,N_14844,N_14150);
nor U17775 (N_17775,N_15949,N_14034);
and U17776 (N_17776,N_14721,N_14457);
nor U17777 (N_17777,N_15435,N_15740);
xnor U17778 (N_17778,N_14225,N_14047);
and U17779 (N_17779,N_14195,N_14675);
and U17780 (N_17780,N_14504,N_15227);
xor U17781 (N_17781,N_15151,N_14439);
nand U17782 (N_17782,N_15446,N_14383);
nor U17783 (N_17783,N_15904,N_14088);
xor U17784 (N_17784,N_15351,N_14136);
nor U17785 (N_17785,N_14045,N_14943);
nand U17786 (N_17786,N_15590,N_15598);
or U17787 (N_17787,N_15971,N_14781);
xor U17788 (N_17788,N_14055,N_15365);
and U17789 (N_17789,N_15582,N_14261);
and U17790 (N_17790,N_14365,N_14715);
nor U17791 (N_17791,N_15258,N_15686);
xnor U17792 (N_17792,N_15586,N_15788);
nor U17793 (N_17793,N_15378,N_15935);
or U17794 (N_17794,N_15168,N_15116);
xor U17795 (N_17795,N_15926,N_15560);
nand U17796 (N_17796,N_15765,N_15768);
and U17797 (N_17797,N_14526,N_15285);
nand U17798 (N_17798,N_14674,N_14061);
nor U17799 (N_17799,N_14251,N_15205);
and U17800 (N_17800,N_15046,N_15002);
or U17801 (N_17801,N_15373,N_14774);
and U17802 (N_17802,N_15260,N_15175);
nand U17803 (N_17803,N_15709,N_15073);
or U17804 (N_17804,N_14502,N_14571);
nor U17805 (N_17805,N_15077,N_15043);
xor U17806 (N_17806,N_14725,N_14793);
and U17807 (N_17807,N_15782,N_15713);
nand U17808 (N_17808,N_14652,N_15364);
nand U17809 (N_17809,N_15180,N_14428);
nand U17810 (N_17810,N_15304,N_14943);
and U17811 (N_17811,N_14836,N_15249);
xor U17812 (N_17812,N_14848,N_14769);
xor U17813 (N_17813,N_14937,N_14261);
or U17814 (N_17814,N_14386,N_14850);
or U17815 (N_17815,N_15671,N_14656);
nand U17816 (N_17816,N_15066,N_14615);
or U17817 (N_17817,N_15201,N_15571);
and U17818 (N_17818,N_15361,N_14274);
nor U17819 (N_17819,N_15995,N_15389);
or U17820 (N_17820,N_15766,N_14421);
xnor U17821 (N_17821,N_15510,N_15625);
or U17822 (N_17822,N_14878,N_14511);
and U17823 (N_17823,N_14778,N_14717);
and U17824 (N_17824,N_15845,N_15155);
nand U17825 (N_17825,N_15302,N_14782);
nor U17826 (N_17826,N_15562,N_14068);
or U17827 (N_17827,N_14390,N_14928);
nand U17828 (N_17828,N_15798,N_15751);
and U17829 (N_17829,N_14185,N_15506);
nor U17830 (N_17830,N_15030,N_14621);
nor U17831 (N_17831,N_15972,N_15031);
xor U17832 (N_17832,N_15316,N_14295);
nor U17833 (N_17833,N_14505,N_15879);
and U17834 (N_17834,N_14521,N_15863);
nor U17835 (N_17835,N_14289,N_14040);
or U17836 (N_17836,N_14070,N_14907);
or U17837 (N_17837,N_15213,N_14527);
xor U17838 (N_17838,N_14209,N_15530);
xnor U17839 (N_17839,N_14892,N_15023);
and U17840 (N_17840,N_15995,N_14928);
and U17841 (N_17841,N_14035,N_15334);
xnor U17842 (N_17842,N_15248,N_15407);
or U17843 (N_17843,N_15214,N_14591);
or U17844 (N_17844,N_14166,N_15550);
or U17845 (N_17845,N_15354,N_15474);
and U17846 (N_17846,N_14691,N_15868);
and U17847 (N_17847,N_14999,N_15062);
nand U17848 (N_17848,N_15478,N_15950);
or U17849 (N_17849,N_14544,N_15048);
nand U17850 (N_17850,N_14404,N_15528);
or U17851 (N_17851,N_14892,N_14616);
nand U17852 (N_17852,N_15539,N_15307);
nor U17853 (N_17853,N_14296,N_14245);
or U17854 (N_17854,N_14549,N_15854);
nor U17855 (N_17855,N_15288,N_14265);
and U17856 (N_17856,N_15129,N_15114);
and U17857 (N_17857,N_15757,N_14474);
and U17858 (N_17858,N_15717,N_14343);
and U17859 (N_17859,N_15870,N_15969);
xnor U17860 (N_17860,N_15080,N_15429);
and U17861 (N_17861,N_15144,N_14428);
xnor U17862 (N_17862,N_15402,N_14020);
nand U17863 (N_17863,N_15982,N_15411);
xor U17864 (N_17864,N_14163,N_14509);
and U17865 (N_17865,N_15883,N_15711);
and U17866 (N_17866,N_14305,N_15323);
nor U17867 (N_17867,N_14684,N_15822);
or U17868 (N_17868,N_15612,N_15607);
nand U17869 (N_17869,N_14753,N_15516);
nor U17870 (N_17870,N_14734,N_14101);
and U17871 (N_17871,N_15974,N_15908);
or U17872 (N_17872,N_14557,N_14666);
or U17873 (N_17873,N_15976,N_14679);
xor U17874 (N_17874,N_14508,N_14007);
nor U17875 (N_17875,N_14657,N_14442);
or U17876 (N_17876,N_14385,N_14282);
nor U17877 (N_17877,N_15291,N_15712);
or U17878 (N_17878,N_14425,N_15117);
nor U17879 (N_17879,N_15857,N_15178);
and U17880 (N_17880,N_15936,N_15511);
or U17881 (N_17881,N_14784,N_14206);
nor U17882 (N_17882,N_14347,N_14179);
xor U17883 (N_17883,N_14785,N_15501);
and U17884 (N_17884,N_14228,N_14829);
nor U17885 (N_17885,N_14272,N_15581);
nand U17886 (N_17886,N_14210,N_14979);
nand U17887 (N_17887,N_14649,N_15163);
or U17888 (N_17888,N_14363,N_15542);
xnor U17889 (N_17889,N_15727,N_14524);
nand U17890 (N_17890,N_15241,N_15598);
nand U17891 (N_17891,N_15253,N_14484);
and U17892 (N_17892,N_15493,N_15436);
nor U17893 (N_17893,N_15578,N_14838);
nand U17894 (N_17894,N_14346,N_15370);
and U17895 (N_17895,N_14692,N_15095);
xnor U17896 (N_17896,N_15909,N_14067);
or U17897 (N_17897,N_15165,N_14690);
xnor U17898 (N_17898,N_14842,N_14864);
or U17899 (N_17899,N_15803,N_15487);
xor U17900 (N_17900,N_15283,N_15972);
nor U17901 (N_17901,N_15229,N_15492);
xnor U17902 (N_17902,N_15927,N_15534);
or U17903 (N_17903,N_15894,N_14843);
or U17904 (N_17904,N_14173,N_15228);
nor U17905 (N_17905,N_14653,N_14928);
and U17906 (N_17906,N_14714,N_14589);
or U17907 (N_17907,N_15340,N_15829);
or U17908 (N_17908,N_15604,N_14611);
nand U17909 (N_17909,N_15048,N_15499);
or U17910 (N_17910,N_14143,N_15266);
and U17911 (N_17911,N_14790,N_15372);
nor U17912 (N_17912,N_15160,N_15738);
nor U17913 (N_17913,N_15499,N_14693);
nand U17914 (N_17914,N_14303,N_15446);
or U17915 (N_17915,N_14978,N_14671);
or U17916 (N_17916,N_14193,N_14604);
or U17917 (N_17917,N_14436,N_15993);
xnor U17918 (N_17918,N_15935,N_15629);
nand U17919 (N_17919,N_15479,N_15944);
and U17920 (N_17920,N_14120,N_15822);
xor U17921 (N_17921,N_15317,N_15927);
xor U17922 (N_17922,N_14429,N_14478);
and U17923 (N_17923,N_15266,N_15770);
or U17924 (N_17924,N_14847,N_15158);
or U17925 (N_17925,N_15854,N_15420);
xor U17926 (N_17926,N_14795,N_14220);
and U17927 (N_17927,N_15293,N_14490);
and U17928 (N_17928,N_15227,N_14870);
and U17929 (N_17929,N_15703,N_14552);
nand U17930 (N_17930,N_14695,N_15886);
nor U17931 (N_17931,N_14469,N_14697);
xor U17932 (N_17932,N_14148,N_15154);
or U17933 (N_17933,N_15233,N_14794);
and U17934 (N_17934,N_15865,N_14176);
and U17935 (N_17935,N_15156,N_15939);
and U17936 (N_17936,N_14962,N_15571);
xnor U17937 (N_17937,N_15643,N_14867);
or U17938 (N_17938,N_15245,N_15614);
and U17939 (N_17939,N_15487,N_15512);
and U17940 (N_17940,N_15892,N_15313);
xnor U17941 (N_17941,N_15694,N_15475);
nor U17942 (N_17942,N_14787,N_15227);
nand U17943 (N_17943,N_14543,N_14322);
nand U17944 (N_17944,N_15264,N_15338);
xnor U17945 (N_17945,N_14223,N_14506);
nand U17946 (N_17946,N_14586,N_15222);
nand U17947 (N_17947,N_15466,N_14318);
xor U17948 (N_17948,N_15311,N_15607);
or U17949 (N_17949,N_14420,N_14831);
nor U17950 (N_17950,N_15153,N_14275);
xnor U17951 (N_17951,N_14864,N_15944);
nand U17952 (N_17952,N_15206,N_14075);
nor U17953 (N_17953,N_14399,N_14552);
nand U17954 (N_17954,N_15031,N_14524);
nand U17955 (N_17955,N_15507,N_15549);
xor U17956 (N_17956,N_15840,N_14064);
and U17957 (N_17957,N_15606,N_15392);
nand U17958 (N_17958,N_15921,N_15205);
and U17959 (N_17959,N_15529,N_14551);
and U17960 (N_17960,N_14096,N_15823);
nor U17961 (N_17961,N_14951,N_14528);
xnor U17962 (N_17962,N_15402,N_15794);
xnor U17963 (N_17963,N_14631,N_15587);
xor U17964 (N_17964,N_14474,N_15759);
and U17965 (N_17965,N_14534,N_15388);
and U17966 (N_17966,N_14894,N_14720);
or U17967 (N_17967,N_14669,N_14303);
nand U17968 (N_17968,N_14389,N_14341);
and U17969 (N_17969,N_14125,N_15071);
nor U17970 (N_17970,N_14037,N_15492);
nor U17971 (N_17971,N_15446,N_15304);
xor U17972 (N_17972,N_14258,N_14516);
nor U17973 (N_17973,N_15624,N_14802);
and U17974 (N_17974,N_15597,N_14695);
xnor U17975 (N_17975,N_14645,N_15527);
or U17976 (N_17976,N_15590,N_14776);
nand U17977 (N_17977,N_14083,N_15743);
nor U17978 (N_17978,N_15328,N_14879);
nand U17979 (N_17979,N_15318,N_14791);
and U17980 (N_17980,N_15211,N_15582);
or U17981 (N_17981,N_15438,N_14797);
xnor U17982 (N_17982,N_15398,N_15200);
or U17983 (N_17983,N_15717,N_14437);
nor U17984 (N_17984,N_15098,N_15148);
nand U17985 (N_17985,N_14594,N_15543);
nor U17986 (N_17986,N_15624,N_14413);
nor U17987 (N_17987,N_14191,N_14667);
nand U17988 (N_17988,N_15606,N_15922);
nand U17989 (N_17989,N_15611,N_14046);
nand U17990 (N_17990,N_15630,N_15829);
nand U17991 (N_17991,N_15870,N_15115);
nor U17992 (N_17992,N_14622,N_14137);
and U17993 (N_17993,N_14051,N_15799);
xor U17994 (N_17994,N_15347,N_15456);
and U17995 (N_17995,N_15970,N_15760);
xnor U17996 (N_17996,N_15318,N_15239);
nand U17997 (N_17997,N_15375,N_14526);
nor U17998 (N_17998,N_15052,N_15960);
xnor U17999 (N_17999,N_15473,N_15469);
or U18000 (N_18000,N_16531,N_16157);
and U18001 (N_18001,N_16668,N_17402);
and U18002 (N_18002,N_16959,N_16426);
and U18003 (N_18003,N_16336,N_16038);
or U18004 (N_18004,N_17231,N_17528);
nand U18005 (N_18005,N_16395,N_17172);
or U18006 (N_18006,N_17039,N_16517);
or U18007 (N_18007,N_16958,N_16684);
nand U18008 (N_18008,N_17356,N_17941);
nand U18009 (N_18009,N_16881,N_16381);
or U18010 (N_18010,N_16377,N_17094);
or U18011 (N_18011,N_17724,N_16156);
xor U18012 (N_18012,N_16745,N_17992);
nor U18013 (N_18013,N_16616,N_17346);
xnor U18014 (N_18014,N_17970,N_17793);
and U18015 (N_18015,N_17519,N_17440);
or U18016 (N_18016,N_17608,N_17731);
nand U18017 (N_18017,N_16901,N_17108);
and U18018 (N_18018,N_16170,N_16705);
nor U18019 (N_18019,N_17980,N_17304);
xor U18020 (N_18020,N_17076,N_17553);
and U18021 (N_18021,N_17461,N_16895);
nor U18022 (N_18022,N_17091,N_17743);
and U18023 (N_18023,N_16573,N_17267);
or U18024 (N_18024,N_17698,N_17432);
or U18025 (N_18025,N_16441,N_17053);
xor U18026 (N_18026,N_17863,N_16561);
nand U18027 (N_18027,N_17224,N_17976);
xnor U18028 (N_18028,N_17423,N_17771);
xor U18029 (N_18029,N_17398,N_16743);
nand U18030 (N_18030,N_17012,N_17547);
xnor U18031 (N_18031,N_17119,N_16950);
xnor U18032 (N_18032,N_16342,N_17165);
nor U18033 (N_18033,N_17985,N_16594);
and U18034 (N_18034,N_17549,N_17657);
xnor U18035 (N_18035,N_16197,N_16001);
and U18036 (N_18036,N_17428,N_16279);
and U18037 (N_18037,N_16435,N_16368);
xor U18038 (N_18038,N_17275,N_17033);
nand U18039 (N_18039,N_16422,N_17691);
and U18040 (N_18040,N_16367,N_17372);
nor U18041 (N_18041,N_16434,N_17185);
and U18042 (N_18042,N_17931,N_16521);
xnor U18043 (N_18043,N_17288,N_16070);
or U18044 (N_18044,N_17125,N_16524);
nor U18045 (N_18045,N_17854,N_17090);
nor U18046 (N_18046,N_16412,N_17445);
and U18047 (N_18047,N_17601,N_16563);
and U18048 (N_18048,N_16662,N_16045);
nor U18049 (N_18049,N_17830,N_16604);
or U18050 (N_18050,N_16482,N_16960);
xnor U18051 (N_18051,N_16344,N_17485);
nand U18052 (N_18052,N_16077,N_16364);
nor U18053 (N_18053,N_17093,N_16299);
nand U18054 (N_18054,N_17487,N_16549);
nand U18055 (N_18055,N_17268,N_17826);
and U18056 (N_18056,N_17087,N_17531);
nor U18057 (N_18057,N_16719,N_16736);
or U18058 (N_18058,N_16453,N_17686);
xnor U18059 (N_18059,N_16935,N_16614);
or U18060 (N_18060,N_17236,N_17962);
xor U18061 (N_18061,N_17943,N_16980);
nor U18062 (N_18062,N_17321,N_16021);
and U18063 (N_18063,N_17891,N_16927);
xor U18064 (N_18064,N_17458,N_17124);
nand U18065 (N_18065,N_16809,N_17562);
or U18066 (N_18066,N_17895,N_16853);
and U18067 (N_18067,N_16108,N_17987);
or U18068 (N_18068,N_16158,N_16995);
or U18069 (N_18069,N_17331,N_16909);
nand U18070 (N_18070,N_16866,N_17928);
xnor U18071 (N_18071,N_16069,N_17182);
nand U18072 (N_18072,N_16824,N_17322);
nor U18073 (N_18073,N_17490,N_16635);
or U18074 (N_18074,N_17259,N_17038);
nand U18075 (N_18075,N_17750,N_17362);
nor U18076 (N_18076,N_16298,N_16555);
or U18077 (N_18077,N_16421,N_17235);
nor U18078 (N_18078,N_17251,N_16716);
nand U18079 (N_18079,N_16815,N_16078);
xor U18080 (N_18080,N_17955,N_16354);
nand U18081 (N_18081,N_16964,N_17779);
xnor U18082 (N_18082,N_16496,N_17064);
xor U18083 (N_18083,N_16418,N_17568);
nor U18084 (N_18084,N_17320,N_16707);
and U18085 (N_18085,N_17856,N_16807);
or U18086 (N_18086,N_17969,N_16908);
or U18087 (N_18087,N_16530,N_16945);
and U18088 (N_18088,N_17246,N_16844);
nor U18089 (N_18089,N_17438,N_17245);
and U18090 (N_18090,N_16355,N_17068);
and U18091 (N_18091,N_16763,N_17619);
nor U18092 (N_18092,N_16822,N_16951);
nand U18093 (N_18093,N_17984,N_16181);
and U18094 (N_18094,N_16526,N_17873);
and U18095 (N_18095,N_17279,N_16138);
xor U18096 (N_18096,N_16989,N_17489);
nand U18097 (N_18097,N_16969,N_17898);
and U18098 (N_18098,N_17991,N_16557);
and U18099 (N_18099,N_17617,N_16293);
nor U18100 (N_18100,N_17517,N_16952);
nor U18101 (N_18101,N_16024,N_16667);
nand U18102 (N_18102,N_17130,N_17846);
or U18103 (N_18103,N_17741,N_17369);
or U18104 (N_18104,N_16320,N_17887);
or U18105 (N_18105,N_17406,N_17083);
nor U18106 (N_18106,N_17579,N_16379);
or U18107 (N_18107,N_16494,N_16553);
and U18108 (N_18108,N_17735,N_17632);
xnor U18109 (N_18109,N_16456,N_16839);
nand U18110 (N_18110,N_16227,N_16750);
xnor U18111 (N_18111,N_17760,N_17794);
nor U18112 (N_18112,N_16501,N_17047);
xnor U18113 (N_18113,N_17483,N_16359);
nand U18114 (N_18114,N_17169,N_17569);
xor U18115 (N_18115,N_16440,N_16335);
xor U18116 (N_18116,N_17388,N_16663);
or U18117 (N_18117,N_17805,N_17052);
nand U18118 (N_18118,N_16455,N_16117);
and U18119 (N_18119,N_16328,N_17013);
and U18120 (N_18120,N_16163,N_17503);
xnor U18121 (N_18121,N_16887,N_16398);
xor U18122 (N_18122,N_17082,N_16762);
or U18123 (N_18123,N_16698,N_16308);
nor U18124 (N_18124,N_16796,N_17782);
nand U18125 (N_18125,N_17494,N_16782);
or U18126 (N_18126,N_17069,N_17103);
nor U18127 (N_18127,N_17383,N_16444);
and U18128 (N_18128,N_17370,N_17946);
nand U18129 (N_18129,N_16489,N_17202);
and U18130 (N_18130,N_16975,N_16845);
or U18131 (N_18131,N_17447,N_16110);
and U18132 (N_18132,N_16739,N_16244);
or U18133 (N_18133,N_16589,N_16066);
and U18134 (N_18134,N_16143,N_16934);
xnor U18135 (N_18135,N_17729,N_17152);
and U18136 (N_18136,N_17936,N_17371);
nand U18137 (N_18137,N_17436,N_16136);
xor U18138 (N_18138,N_16900,N_16431);
or U18139 (N_18139,N_16481,N_16650);
xnor U18140 (N_18140,N_17473,N_17335);
and U18141 (N_18141,N_17376,N_17089);
xor U18142 (N_18142,N_16546,N_17136);
or U18143 (N_18143,N_17211,N_17102);
nand U18144 (N_18144,N_17162,N_16034);
nand U18145 (N_18145,N_17692,N_17871);
nor U18146 (N_18146,N_16888,N_16100);
nand U18147 (N_18147,N_16926,N_16920);
nor U18148 (N_18148,N_17964,N_17084);
and U18149 (N_18149,N_16903,N_16597);
or U18150 (N_18150,N_17128,N_16384);
nor U18151 (N_18151,N_16838,N_17904);
or U18152 (N_18152,N_16089,N_17265);
xor U18153 (N_18153,N_17159,N_17277);
nand U18154 (N_18154,N_16661,N_17008);
nor U18155 (N_18155,N_16488,N_17109);
nor U18156 (N_18156,N_16651,N_16169);
xor U18157 (N_18157,N_16309,N_16943);
and U18158 (N_18158,N_17627,N_17394);
nor U18159 (N_18159,N_16141,N_17937);
nor U18160 (N_18160,N_16751,N_17700);
or U18161 (N_18161,N_17051,N_16288);
nand U18162 (N_18162,N_16334,N_17187);
xor U18163 (N_18163,N_17542,N_16697);
xor U18164 (N_18164,N_17551,N_16775);
or U18165 (N_18165,N_17550,N_17944);
nand U18166 (N_18166,N_17066,N_17806);
xnor U18167 (N_18167,N_17416,N_16011);
and U18168 (N_18168,N_16883,N_17032);
nand U18169 (N_18169,N_17430,N_16500);
or U18170 (N_18170,N_16723,N_17634);
xor U18171 (N_18171,N_17882,N_17845);
and U18172 (N_18172,N_16201,N_17683);
nand U18173 (N_18173,N_17009,N_16812);
or U18174 (N_18174,N_16889,N_17557);
or U18175 (N_18175,N_17253,N_17753);
xnor U18176 (N_18176,N_16990,N_17841);
xnor U18177 (N_18177,N_17527,N_17770);
or U18178 (N_18178,N_16856,N_17607);
and U18179 (N_18179,N_16267,N_17983);
or U18180 (N_18180,N_17546,N_17639);
xor U18181 (N_18181,N_17513,N_16596);
nand U18182 (N_18182,N_16074,N_16305);
nand U18183 (N_18183,N_16884,N_16930);
and U18184 (N_18184,N_17704,N_16852);
or U18185 (N_18185,N_17380,N_16084);
and U18186 (N_18186,N_16946,N_17583);
xnor U18187 (N_18187,N_17431,N_16353);
xor U18188 (N_18188,N_17533,N_17828);
nor U18189 (N_18189,N_17341,N_17474);
nand U18190 (N_18190,N_16673,N_16487);
nor U18191 (N_18191,N_17041,N_16544);
nand U18192 (N_18192,N_16522,N_17821);
xnor U18193 (N_18193,N_17726,N_16327);
nor U18194 (N_18194,N_16701,N_17932);
or U18195 (N_18195,N_16675,N_17139);
nor U18196 (N_18196,N_17464,N_17006);
xnor U18197 (N_18197,N_16362,N_16102);
nand U18198 (N_18198,N_17392,N_17777);
or U18199 (N_18199,N_16532,N_17342);
nand U18200 (N_18200,N_17712,N_17405);
and U18201 (N_18201,N_16027,N_16185);
or U18202 (N_18202,N_16874,N_16509);
xor U18203 (N_18203,N_17397,N_16459);
and U18204 (N_18204,N_16670,N_17104);
xnor U18205 (N_18205,N_17641,N_16741);
or U18206 (N_18206,N_16864,N_16240);
and U18207 (N_18207,N_16265,N_17669);
nor U18208 (N_18208,N_16712,N_16800);
and U18209 (N_18209,N_16880,N_16140);
nand U18210 (N_18210,N_16865,N_16725);
xor U18211 (N_18211,N_17243,N_17488);
and U18212 (N_18212,N_16198,N_17061);
nand U18213 (N_18213,N_16803,N_17186);
or U18214 (N_18214,N_16630,N_16634);
nor U18215 (N_18215,N_16237,N_16000);
xor U18216 (N_18216,N_16872,N_16049);
nor U18217 (N_18217,N_17018,N_16988);
xnor U18218 (N_18218,N_17306,N_16817);
nand U18219 (N_18219,N_17294,N_17667);
nor U18220 (N_18220,N_17674,N_17857);
or U18221 (N_18221,N_17633,N_16470);
and U18222 (N_18222,N_17822,N_16828);
and U18223 (N_18223,N_17905,N_16764);
or U18224 (N_18224,N_16813,N_16028);
nor U18225 (N_18225,N_16569,N_16176);
xor U18226 (N_18226,N_17520,N_16540);
xor U18227 (N_18227,N_16939,N_16598);
xnor U18228 (N_18228,N_17188,N_17518);
and U18229 (N_18229,N_17646,N_16525);
or U18230 (N_18230,N_17525,N_16632);
nor U18231 (N_18231,N_16985,N_17690);
and U18232 (N_18232,N_17734,N_16241);
nor U18233 (N_18233,N_16849,N_16829);
nand U18234 (N_18234,N_16080,N_16119);
xnor U18235 (N_18235,N_16399,N_17552);
xnor U18236 (N_18236,N_16221,N_16579);
and U18237 (N_18237,N_16996,N_17659);
nand U18238 (N_18238,N_16093,N_16647);
nand U18239 (N_18239,N_17373,N_16250);
and U18240 (N_18240,N_16644,N_17400);
or U18241 (N_18241,N_16213,N_17466);
or U18242 (N_18242,N_17647,N_17902);
and U18243 (N_18243,N_17271,N_16006);
nand U18244 (N_18244,N_17786,N_17914);
nand U18245 (N_18245,N_17001,N_16735);
and U18246 (N_18246,N_17209,N_16624);
nor U18247 (N_18247,N_17878,N_17880);
xnor U18248 (N_18248,N_16897,N_16311);
nand U18249 (N_18249,N_16107,N_17301);
and U18250 (N_18250,N_16154,N_16877);
nand U18251 (N_18251,N_16721,N_16660);
nor U18252 (N_18252,N_16404,N_16506);
xnor U18253 (N_18253,N_16203,N_17129);
or U18254 (N_18254,N_16846,N_17471);
xor U18255 (N_18255,N_17442,N_17570);
and U18256 (N_18256,N_17010,N_17628);
nand U18257 (N_18257,N_16599,N_16423);
xor U18258 (N_18258,N_17879,N_16373);
nor U18259 (N_18259,N_17592,N_16669);
nor U18260 (N_18260,N_16101,N_16122);
xor U18261 (N_18261,N_16297,N_17589);
xnor U18262 (N_18262,N_16977,N_17446);
nand U18263 (N_18263,N_16436,N_16276);
xnor U18264 (N_18264,N_17216,N_17935);
or U18265 (N_18265,N_16858,N_17584);
xor U18266 (N_18266,N_16340,N_17208);
xor U18267 (N_18267,N_16017,N_17972);
and U18268 (N_18268,N_16523,N_17204);
xnor U18269 (N_18269,N_17529,N_16683);
nand U18270 (N_18270,N_17756,N_17758);
xor U18271 (N_18271,N_17284,N_17606);
xnor U18272 (N_18272,N_16665,N_17459);
or U18273 (N_18273,N_17926,N_17078);
nor U18274 (N_18274,N_16711,N_16976);
nor U18275 (N_18275,N_17708,N_17142);
xor U18276 (N_18276,N_16015,N_16005);
xor U18277 (N_18277,N_16300,N_16729);
nor U18278 (N_18278,N_17853,N_17282);
nand U18279 (N_18279,N_16868,N_16837);
nor U18280 (N_18280,N_16035,N_16202);
nand U18281 (N_18281,N_16871,N_17834);
nor U18282 (N_18282,N_17333,N_16539);
nor U18283 (N_18283,N_16648,N_17610);
and U18284 (N_18284,N_17979,N_16007);
xor U18285 (N_18285,N_17965,N_17448);
xor U18286 (N_18286,N_17482,N_17860);
and U18287 (N_18287,N_17994,N_17024);
xor U18288 (N_18288,N_16036,N_16442);
xnor U18289 (N_18289,N_17126,N_16681);
and U18290 (N_18290,N_17577,N_17548);
and U18291 (N_18291,N_17989,N_16462);
nand U18292 (N_18292,N_17276,N_17100);
or U18293 (N_18293,N_17951,N_17117);
xor U18294 (N_18294,N_17063,N_17353);
xnor U18295 (N_18295,N_17347,N_17776);
xor U18296 (N_18296,N_16814,N_17167);
nor U18297 (N_18297,N_16702,N_16642);
and U18298 (N_18298,N_17950,N_17654);
or U18299 (N_18299,N_16755,N_17661);
xnor U18300 (N_18300,N_17868,N_16495);
or U18301 (N_18301,N_16406,N_17769);
nor U18302 (N_18302,N_17198,N_17191);
or U18303 (N_18303,N_16284,N_16571);
or U18304 (N_18304,N_17644,N_16037);
nor U18305 (N_18305,N_16533,N_17254);
nor U18306 (N_18306,N_17007,N_16730);
xnor U18307 (N_18307,N_17508,N_17449);
nand U18308 (N_18308,N_17214,N_17739);
or U18309 (N_18309,N_17832,N_17986);
and U18310 (N_18310,N_16551,N_16057);
nor U18311 (N_18311,N_16709,N_16728);
nor U18312 (N_18312,N_16123,N_16727);
or U18313 (N_18313,N_16899,N_17855);
xor U18314 (N_18314,N_16637,N_17164);
nand U18315 (N_18315,N_17435,N_17207);
xnor U18316 (N_18316,N_17960,N_16556);
nor U18317 (N_18317,N_17813,N_17916);
or U18318 (N_18318,N_17261,N_16583);
and U18319 (N_18319,N_17827,N_17355);
or U18320 (N_18320,N_17505,N_17509);
or U18321 (N_18321,N_17316,N_17391);
xor U18322 (N_18322,N_16165,N_17924);
and U18323 (N_18323,N_17496,N_17414);
and U18324 (N_18324,N_17472,N_17278);
or U18325 (N_18325,N_16870,N_17893);
or U18326 (N_18326,N_16629,N_17071);
nor U18327 (N_18327,N_17651,N_16348);
xor U18328 (N_18328,N_17266,N_16978);
nand U18329 (N_18329,N_17839,N_17219);
nand U18330 (N_18330,N_16262,N_17718);
and U18331 (N_18331,N_16235,N_16717);
or U18332 (N_18332,N_16582,N_16286);
and U18333 (N_18333,N_16720,N_17740);
nand U18334 (N_18334,N_16068,N_16692);
xnor U18335 (N_18335,N_16620,N_16780);
and U18336 (N_18336,N_17598,N_16061);
xnor U18337 (N_18337,N_16639,N_17377);
xor U18338 (N_18338,N_17819,N_16792);
or U18339 (N_18339,N_17798,N_16578);
and U18340 (N_18340,N_16438,N_17767);
nand U18341 (N_18341,N_17721,N_16403);
nor U18342 (N_18342,N_17810,N_16568);
or U18343 (N_18343,N_16010,N_16149);
and U18344 (N_18344,N_16636,N_17307);
nor U18345 (N_18345,N_16797,N_16854);
and U18346 (N_18346,N_16282,N_16454);
and U18347 (N_18347,N_17410,N_16559);
or U18348 (N_18348,N_17714,N_16216);
xor U18349 (N_18349,N_16111,N_16627);
xor U18350 (N_18350,N_16774,N_17982);
nand U18351 (N_18351,N_16703,N_17566);
and U18352 (N_18352,N_17910,N_17359);
or U18353 (N_18353,N_16484,N_16260);
or U18354 (N_18354,N_16894,N_17919);
and U18355 (N_18355,N_17002,N_17155);
xor U18356 (N_18356,N_17176,N_16891);
nand U18357 (N_18357,N_17016,N_17419);
or U18358 (N_18358,N_16558,N_16292);
and U18359 (N_18359,N_17157,N_16173);
or U18360 (N_18360,N_17707,N_16307);
nand U18361 (N_18361,N_17521,N_17652);
and U18362 (N_18362,N_17274,N_16974);
nor U18363 (N_18363,N_17604,N_16962);
nand U18364 (N_18364,N_17844,N_16137);
xor U18365 (N_18365,N_17801,N_17611);
nand U18366 (N_18366,N_16323,N_17722);
and U18367 (N_18367,N_16219,N_17427);
and U18368 (N_18368,N_17475,N_17825);
and U18369 (N_18369,N_17842,N_16679);
nor U18370 (N_18370,N_17947,N_17189);
or U18371 (N_18371,N_17404,N_17463);
and U18372 (N_18372,N_17417,N_17501);
nor U18373 (N_18373,N_16312,N_16082);
and U18374 (N_18374,N_16593,N_17334);
nor U18375 (N_18375,N_17178,N_17365);
or U18376 (N_18376,N_17889,N_16352);
or U18377 (N_18377,N_16911,N_16033);
or U18378 (N_18378,N_16249,N_16686);
xnor U18379 (N_18379,N_17133,N_17057);
xor U18380 (N_18380,N_16936,N_17468);
and U18381 (N_18381,N_17759,N_17328);
and U18382 (N_18382,N_16491,N_16331);
or U18383 (N_18383,N_17539,N_17800);
xor U18384 (N_18384,N_17649,N_17273);
nor U18385 (N_18385,N_16004,N_17096);
xnor U18386 (N_18386,N_16690,N_16124);
or U18387 (N_18387,N_17723,N_17263);
nor U18388 (N_18388,N_17077,N_17462);
and U18389 (N_18389,N_16464,N_17203);
nand U18390 (N_18390,N_16550,N_16139);
or U18391 (N_18391,N_17314,N_16788);
nand U18392 (N_18392,N_17455,N_16758);
nand U18393 (N_18393,N_17351,N_17673);
or U18394 (N_18394,N_16645,N_17578);
nand U18395 (N_18395,N_17545,N_17280);
nor U18396 (N_18396,N_16254,N_16724);
or U18397 (N_18397,N_16103,N_16982);
nor U18398 (N_18398,N_17114,N_16357);
nor U18399 (N_18399,N_16228,N_17218);
or U18400 (N_18400,N_16979,N_17030);
or U18401 (N_18401,N_16079,N_17981);
nor U18402 (N_18402,N_17797,N_16178);
nand U18403 (N_18403,N_16086,N_17787);
and U18404 (N_18404,N_16003,N_16699);
nand U18405 (N_18405,N_16904,N_17792);
nor U18406 (N_18406,N_17510,N_16230);
nand U18407 (N_18407,N_17507,N_17506);
or U18408 (N_18408,N_17134,N_16121);
xor U18409 (N_18409,N_16268,N_17581);
or U18410 (N_18410,N_16562,N_16840);
xnor U18411 (N_18411,N_16275,N_16700);
or U18412 (N_18412,N_16125,N_16825);
xor U18413 (N_18413,N_17939,N_17662);
nand U18414 (N_18414,N_17558,N_17424);
and U18415 (N_18415,N_17004,N_17381);
xnor U18416 (N_18416,N_16259,N_16789);
nor U18417 (N_18417,N_16882,N_17311);
nand U18418 (N_18418,N_16574,N_16674);
and U18419 (N_18419,N_17146,N_16430);
xnor U18420 (N_18420,N_17850,N_16941);
or U18421 (N_18421,N_16302,N_16694);
or U18422 (N_18422,N_17368,N_16126);
nand U18423 (N_18423,N_17618,N_17585);
and U18424 (N_18424,N_17948,N_17364);
nand U18425 (N_18425,N_16655,N_17180);
and U18426 (N_18426,N_17808,N_16973);
xnor U18427 (N_18427,N_17894,N_16025);
nand U18428 (N_18428,N_17961,N_16704);
nor U18429 (N_18429,N_16830,N_16785);
xnor U18430 (N_18430,N_17681,N_16051);
and U18431 (N_18431,N_17451,N_16180);
nand U18432 (N_18432,N_16835,N_17945);
xnor U18433 (N_18433,N_17345,N_16433);
or U18434 (N_18434,N_16691,N_17768);
xor U18435 (N_18435,N_17166,N_17684);
xor U18436 (N_18436,N_17666,N_16746);
or U18437 (N_18437,N_16022,N_16109);
or U18438 (N_18438,N_16097,N_16928);
or U18439 (N_18439,N_17378,N_16390);
xnor U18440 (N_18440,N_17861,N_16625);
or U18441 (N_18441,N_17678,N_16515);
and U18442 (N_18442,N_17403,N_17967);
xor U18443 (N_18443,N_16280,N_17859);
or U18444 (N_18444,N_17701,N_16878);
nand U18445 (N_18445,N_17453,N_17147);
and U18446 (N_18446,N_16113,N_17366);
xor U18447 (N_18447,N_16182,N_17014);
nor U18448 (N_18448,N_17422,N_16287);
xnor U18449 (N_18449,N_16347,N_17361);
and U18450 (N_18450,N_16850,N_16925);
nor U18451 (N_18451,N_16233,N_16791);
nor U18452 (N_18452,N_17222,N_16446);
or U18453 (N_18453,N_16492,N_17746);
nor U18454 (N_18454,N_16777,N_17221);
or U18455 (N_18455,N_16094,N_17865);
xor U18456 (N_18456,N_16688,N_17055);
xnor U18457 (N_18457,N_16095,N_16740);
nor U18458 (N_18458,N_16810,N_16548);
or U18459 (N_18459,N_17412,N_17564);
xor U18460 (N_18460,N_16917,N_16938);
and U18461 (N_18461,N_17387,N_17688);
nand U18462 (N_18462,N_16341,N_16190);
xor U18463 (N_18463,N_17903,N_17241);
and U18464 (N_18464,N_16961,N_16458);
nor U18465 (N_18465,N_16547,N_16767);
nor U18466 (N_18466,N_16383,N_17193);
or U18467 (N_18467,N_17795,N_16948);
nor U18468 (N_18468,N_16319,N_17054);
or U18469 (N_18469,N_17867,N_17154);
nor U18470 (N_18470,N_17151,N_17837);
or U18471 (N_18471,N_16304,N_16536);
nor U18472 (N_18472,N_17418,N_16765);
nand U18473 (N_18473,N_17663,N_16325);
nand U18474 (N_18474,N_17612,N_16296);
xnor U18475 (N_18475,N_17396,N_17137);
nand U18476 (N_18476,N_17095,N_16225);
or U18477 (N_18477,N_16088,N_17120);
and U18478 (N_18478,N_16414,N_17535);
nand U18479 (N_18479,N_17804,N_17113);
or U18480 (N_18480,N_16255,N_17660);
or U18481 (N_18481,N_16892,N_17493);
xnor U18482 (N_18482,N_17298,N_17325);
xor U18483 (N_18483,N_17065,N_17824);
nand U18484 (N_18484,N_17358,N_17622);
and U18485 (N_18485,N_16998,N_17693);
xor U18486 (N_18486,N_17866,N_17258);
xnor U18487 (N_18487,N_17917,N_16360);
or U18488 (N_18488,N_16640,N_16738);
and U18489 (N_18489,N_16223,N_16372);
and U18490 (N_18490,N_16214,N_17689);
nand U18491 (N_18491,N_17292,N_17732);
and U18492 (N_18492,N_16389,N_16339);
or U18493 (N_18493,N_16243,N_16040);
nor U18494 (N_18494,N_17122,N_16552);
xnor U18495 (N_18495,N_16447,N_17900);
xnor U18496 (N_18496,N_16607,N_17590);
or U18497 (N_18497,N_17600,N_16012);
and U18498 (N_18498,N_16685,N_16294);
nand U18499 (N_18499,N_16043,N_17374);
nor U18500 (N_18500,N_17597,N_17687);
and U18501 (N_18501,N_17599,N_17922);
nand U18502 (N_18502,N_16566,N_16916);
xnor U18503 (N_18503,N_16567,N_17602);
nand U18504 (N_18504,N_17144,N_16718);
nand U18505 (N_18505,N_17401,N_17021);
and U18506 (N_18506,N_16041,N_17349);
nand U18507 (N_18507,N_17615,N_16090);
and U18508 (N_18508,N_16167,N_16653);
or U18509 (N_18509,N_16753,N_16714);
xnor U18510 (N_18510,N_16622,N_16477);
and U18511 (N_18511,N_16303,N_16575);
or U18512 (N_18512,N_17680,N_16316);
xor U18513 (N_18513,N_16166,N_16261);
and U18514 (N_18514,N_16062,N_17029);
nor U18515 (N_18515,N_17603,N_16783);
nand U18516 (N_18516,N_17028,N_17309);
xnor U18517 (N_18517,N_17058,N_17042);
nor U18518 (N_18518,N_16873,N_16065);
nand U18519 (N_18519,N_17296,N_16405);
nor U18520 (N_18520,N_17831,N_17481);
xnor U18521 (N_18521,N_16425,N_17523);
or U18522 (N_18522,N_17959,N_17260);
nor U18523 (N_18523,N_16358,N_16248);
nor U18524 (N_18524,N_16385,N_16968);
and U18525 (N_18525,N_16680,N_16473);
nand U18526 (N_18526,N_16270,N_17337);
nand U18527 (N_18527,N_17469,N_16063);
xor U18528 (N_18528,N_16768,N_16333);
nand U18529 (N_18529,N_16171,N_17702);
and U18530 (N_18530,N_17747,N_17150);
nand U18531 (N_18531,N_16511,N_16184);
and U18532 (N_18532,N_16046,N_16565);
and U18533 (N_18533,N_16587,N_16475);
nand U18534 (N_18534,N_16991,N_17088);
or U18535 (N_18535,N_17421,N_17308);
xnor U18536 (N_18536,N_17588,N_16285);
and U18537 (N_18537,N_16733,N_16821);
or U18538 (N_18538,N_16196,N_16710);
xor U18539 (N_18539,N_17499,N_17215);
xor U18540 (N_18540,N_16378,N_16580);
and U18541 (N_18541,N_16072,N_16879);
or U18542 (N_18542,N_17354,N_17762);
nand U18543 (N_18543,N_16811,N_17876);
nand U18544 (N_18544,N_17799,N_16147);
and U18545 (N_18545,N_16924,N_17695);
nor U18546 (N_18546,N_17697,N_16451);
and U18547 (N_18547,N_16457,N_16773);
nand U18548 (N_18548,N_16461,N_16029);
nor U18549 (N_18549,N_17479,N_16204);
or U18550 (N_18550,N_17299,N_16120);
xor U18551 (N_18551,N_16055,N_16460);
nor U18552 (N_18552,N_17596,N_16696);
or U18553 (N_18553,N_16915,N_16400);
and U18554 (N_18554,N_17676,N_17317);
xor U18555 (N_18555,N_16605,N_17785);
nor U18556 (N_18556,N_17210,N_16490);
and U18557 (N_18557,N_16315,N_16150);
nor U18558 (N_18558,N_17067,N_17239);
nor U18559 (N_18559,N_17281,N_16401);
and U18560 (N_18560,N_16224,N_16999);
xor U18561 (N_18561,N_17037,N_16098);
nand U18562 (N_18562,N_16847,N_17930);
nand U18563 (N_18563,N_17194,N_16416);
and U18564 (N_18564,N_17820,N_17360);
nand U18565 (N_18565,N_17778,N_17899);
and U18566 (N_18566,N_16617,N_16600);
nor U18567 (N_18567,N_16199,N_17343);
or U18568 (N_18568,N_17060,N_17862);
and U18569 (N_18569,N_17290,N_16572);
xnor U18570 (N_18570,N_16476,N_17195);
nand U18571 (N_18571,N_17228,N_16295);
and U18572 (N_18572,N_16452,N_16393);
or U18573 (N_18573,N_17140,N_17285);
nand U18574 (N_18574,N_16937,N_16631);
or U18575 (N_18575,N_16754,N_16474);
nor U18576 (N_18576,N_17719,N_17538);
nor U18577 (N_18577,N_17237,N_17196);
nor U18578 (N_18578,N_16678,N_16693);
or U18579 (N_18579,N_16480,N_16291);
or U18580 (N_18580,N_16397,N_17720);
nand U18581 (N_18581,N_17877,N_16192);
nor U18582 (N_18582,N_16886,N_16450);
or U18583 (N_18583,N_16633,N_16621);
xnor U18584 (N_18584,N_17648,N_17460);
nand U18585 (N_18585,N_16483,N_17318);
nand U18586 (N_18586,N_17348,N_17725);
xnor U18587 (N_18587,N_16469,N_17847);
or U18588 (N_18588,N_16893,N_17363);
and U18589 (N_18589,N_17338,N_16966);
and U18590 (N_18590,N_16820,N_17534);
and U18591 (N_18591,N_16326,N_16263);
and U18592 (N_18592,N_16595,N_17815);
or U18593 (N_18593,N_16026,N_17123);
xnor U18594 (N_18594,N_17803,N_17796);
nand U18595 (N_18595,N_17477,N_17415);
nand U18596 (N_18596,N_16602,N_16843);
xnor U18597 (N_18597,N_16842,N_17918);
nand U18598 (N_18598,N_16402,N_17995);
or U18599 (N_18599,N_16609,N_17645);
and U18600 (N_18600,N_16689,N_17554);
xor U18601 (N_18601,N_17892,N_17225);
xor U18602 (N_18602,N_17624,N_17336);
xnor U18603 (N_18603,N_17870,N_17829);
nor U18604 (N_18604,N_16417,N_16770);
nor U18605 (N_18605,N_17145,N_16795);
and U18606 (N_18606,N_17174,N_16756);
xor U18607 (N_18607,N_16677,N_16424);
nand U18608 (N_18608,N_16584,N_16499);
or U18609 (N_18609,N_16955,N_17738);
nand U18610 (N_18610,N_16232,N_17044);
and U18611 (N_18611,N_17395,N_16902);
or U18612 (N_18612,N_16047,N_17197);
and U18613 (N_18613,N_17925,N_17480);
or U18614 (N_18614,N_17572,N_17375);
and U18615 (N_18615,N_17727,N_17300);
or U18616 (N_18616,N_16588,N_17699);
and U18617 (N_18617,N_17205,N_17213);
nand U18618 (N_18618,N_16330,N_16067);
nor U18619 (N_18619,N_16472,N_17685);
or U18620 (N_18620,N_17011,N_16972);
nand U18621 (N_18621,N_17514,N_17399);
xor U18622 (N_18622,N_17389,N_17694);
xnor U18623 (N_18623,N_16222,N_16050);
nor U18624 (N_18624,N_16869,N_16238);
and U18625 (N_18625,N_16671,N_17872);
and U18626 (N_18626,N_16044,N_17230);
and U18627 (N_18627,N_16392,N_17629);
or U18628 (N_18628,N_16212,N_17201);
nor U18629 (N_18629,N_16271,N_16349);
or U18630 (N_18630,N_17884,N_16855);
or U18631 (N_18631,N_17497,N_17256);
xnor U18632 (N_18632,N_17997,N_16570);
nand U18633 (N_18633,N_16752,N_17240);
nor U18634 (N_18634,N_16172,N_17035);
or U18635 (N_18635,N_17929,N_16345);
nand U18636 (N_18636,N_16859,N_17637);
nor U18637 (N_18637,N_17783,N_17444);
and U18638 (N_18638,N_16687,N_16921);
and U18639 (N_18639,N_16769,N_16970);
or U18640 (N_18640,N_16542,N_17788);
nand U18641 (N_18641,N_17357,N_17048);
or U18642 (N_18642,N_16274,N_17457);
xnor U18643 (N_18643,N_17470,N_17175);
nor U18644 (N_18644,N_16831,N_17106);
nor U18645 (N_18645,N_16808,N_17906);
xor U18646 (N_18646,N_17420,N_16396);
nor U18647 (N_18647,N_16971,N_17890);
nor U18648 (N_18648,N_16189,N_16415);
xnor U18649 (N_18649,N_17390,N_16258);
or U18650 (N_18650,N_17560,N_16498);
and U18651 (N_18651,N_16281,N_17183);
nand U18652 (N_18652,N_17217,N_16056);
xor U18653 (N_18653,N_16363,N_17319);
nand U18654 (N_18654,N_16505,N_17433);
xnor U18655 (N_18655,N_16177,N_17949);
xor U18656 (N_18656,N_17233,N_17764);
xnor U18657 (N_18657,N_16060,N_17110);
or U18658 (N_18658,N_16134,N_16014);
xor U18659 (N_18659,N_16042,N_17541);
or U18660 (N_18660,N_17498,N_17181);
and U18661 (N_18661,N_17658,N_17671);
xnor U18662 (N_18662,N_16804,N_17250);
nand U18663 (N_18663,N_17074,N_17326);
or U18664 (N_18664,N_17665,N_16471);
nand U18665 (N_18665,N_17034,N_16153);
and U18666 (N_18666,N_17023,N_17112);
nor U18667 (N_18667,N_16160,N_17567);
or U18668 (N_18668,N_16641,N_16913);
or U18669 (N_18669,N_17733,N_16207);
nor U18670 (N_18670,N_17963,N_16659);
nor U18671 (N_18671,N_16923,N_16146);
xnor U18672 (N_18672,N_17956,N_16407);
nand U18673 (N_18673,N_16467,N_16486);
xor U18674 (N_18674,N_17027,N_16048);
xor U18675 (N_18675,N_16115,N_17163);
and U18676 (N_18676,N_16514,N_17426);
or U18677 (N_18677,N_16283,N_17575);
nor U18678 (N_18678,N_16907,N_16351);
nor U18679 (N_18679,N_16766,N_16508);
xor U18680 (N_18680,N_17025,N_16052);
and U18681 (N_18681,N_16576,N_17848);
nand U18682 (N_18682,N_16619,N_17352);
xnor U18683 (N_18683,N_16242,N_16322);
or U18684 (N_18684,N_17156,N_17059);
xor U18685 (N_18685,N_16799,N_16654);
nand U18686 (N_18686,N_17177,N_16940);
and U18687 (N_18687,N_17875,N_17556);
xnor U18688 (N_18688,N_16220,N_17086);
nor U18689 (N_18689,N_16466,N_17511);
xnor U18690 (N_18690,N_16761,N_16929);
and U18691 (N_18691,N_16520,N_17050);
xor U18692 (N_18692,N_16130,N_16772);
or U18693 (N_18693,N_16085,N_16114);
nand U18694 (N_18694,N_17580,N_17838);
nor U18695 (N_18695,N_16419,N_16096);
xnor U18696 (N_18696,N_17226,N_17532);
nor U18697 (N_18697,N_17968,N_16152);
nand U18698 (N_18698,N_16919,N_16957);
or U18699 (N_18699,N_16666,N_17452);
xnor U18700 (N_18700,N_16510,N_16272);
and U18701 (N_18701,N_17500,N_17626);
nand U18702 (N_18702,N_17536,N_16581);
nand U18703 (N_18703,N_17851,N_17677);
xnor U18704 (N_18704,N_17297,N_17912);
and U18705 (N_18705,N_17653,N_17101);
or U18706 (N_18706,N_16497,N_16944);
or U18707 (N_18707,N_16099,N_17324);
nand U18708 (N_18708,N_17897,N_17291);
or U18709 (N_18709,N_17015,N_17555);
nor U18710 (N_18710,N_17242,N_16519);
xor U18711 (N_18711,N_17940,N_17537);
or U18712 (N_18712,N_16695,N_17141);
or U18713 (N_18713,N_16369,N_17814);
nand U18714 (N_18714,N_17135,N_17515);
and U18715 (N_18715,N_16375,N_17625);
nor U18716 (N_18716,N_17817,N_16314);
xnor U18717 (N_18717,N_16512,N_17679);
nand U18718 (N_18718,N_17737,N_16188);
and U18719 (N_18719,N_17411,N_16183);
and U18720 (N_18720,N_17710,N_17524);
and U18721 (N_18721,N_16318,N_16253);
nand U18722 (N_18722,N_17703,N_17954);
nor U18723 (N_18723,N_16427,N_16543);
or U18724 (N_18724,N_16246,N_16365);
nand U18725 (N_18725,N_17003,N_16914);
and U18726 (N_18726,N_16586,N_17313);
and U18727 (N_18727,N_17565,N_17302);
xnor U18728 (N_18728,N_17247,N_16116);
and U18729 (N_18729,N_17005,N_17227);
or U18730 (N_18730,N_17046,N_16252);
nor U18731 (N_18731,N_17312,N_17999);
nand U18732 (N_18732,N_16211,N_16608);
nand U18733 (N_18733,N_17332,N_16610);
and U18734 (N_18734,N_17773,N_17257);
xnor U18735 (N_18735,N_17544,N_16175);
xor U18736 (N_18736,N_16071,N_16672);
or U18737 (N_18737,N_17736,N_16906);
nand U18738 (N_18738,N_17874,N_17730);
or U18739 (N_18739,N_17031,N_16361);
or U18740 (N_18740,N_16781,N_17593);
or U18741 (N_18741,N_17017,N_16922);
or U18742 (N_18742,N_17642,N_16993);
or U18743 (N_18743,N_16144,N_17062);
nand U18744 (N_18744,N_16413,N_16208);
nand U18745 (N_18745,N_16805,N_17573);
xor U18746 (N_18746,N_16778,N_17909);
nor U18747 (N_18747,N_17942,N_16603);
nor U18748 (N_18748,N_17200,N_17766);
nand U18749 (N_18749,N_16087,N_16931);
nor U18750 (N_18750,N_17283,N_17056);
nand U18751 (N_18751,N_16905,N_17327);
nor U18752 (N_18752,N_17184,N_16161);
and U18753 (N_18753,N_16513,N_16819);
and U18754 (N_18754,N_17836,N_17881);
xnor U18755 (N_18755,N_16749,N_16310);
nor U18756 (N_18756,N_16649,N_17774);
xor U18757 (N_18757,N_16448,N_17675);
nor U18758 (N_18758,N_17467,N_17835);
and U18759 (N_18759,N_16118,N_17576);
xnor U18760 (N_18760,N_17437,N_17709);
or U18761 (N_18761,N_16554,N_17161);
nor U18762 (N_18762,N_16918,N_16485);
and U18763 (N_18763,N_17045,N_16806);
nand U18764 (N_18764,N_17127,N_17772);
nor U18765 (N_18765,N_17978,N_16757);
or U18766 (N_18766,N_16463,N_16428);
nor U18767 (N_18767,N_16890,N_17049);
nand U18768 (N_18768,N_16992,N_16128);
xnor U18769 (N_18769,N_17858,N_16657);
xnor U18770 (N_18770,N_16388,N_16439);
xnor U18771 (N_18771,N_17385,N_16942);
nand U18772 (N_18772,N_16612,N_17491);
or U18773 (N_18773,N_16997,N_16376);
and U18774 (N_18774,N_16896,N_17971);
and U18775 (N_18775,N_16953,N_16493);
xnor U18776 (N_18776,N_16981,N_16408);
or U18777 (N_18777,N_17907,N_16290);
nor U18778 (N_18778,N_17781,N_16545);
or U18779 (N_18779,N_16465,N_16321);
nand U18780 (N_18780,N_17742,N_17705);
nand U18781 (N_18781,N_16105,N_17131);
or U18782 (N_18782,N_16410,N_16737);
and U18783 (N_18783,N_17075,N_17670);
nand U18784 (N_18784,N_17486,N_16002);
nor U18785 (N_18785,N_16289,N_17249);
or U18786 (N_18786,N_16145,N_16541);
or U18787 (N_18787,N_17852,N_16256);
nor U18788 (N_18788,N_16818,N_16264);
or U18789 (N_18789,N_16611,N_16186);
xnor U18790 (N_18790,N_16502,N_17775);
xnor U18791 (N_18791,N_16932,N_17765);
nand U18792 (N_18792,N_16503,N_16643);
and U18793 (N_18793,N_17901,N_16277);
or U18794 (N_18794,N_17269,N_17160);
nand U18795 (N_18795,N_16016,N_16528);
xor U18796 (N_18796,N_17310,N_17636);
nor U18797 (N_18797,N_17640,N_16591);
or U18798 (N_18798,N_16032,N_17289);
nand U18799 (N_18799,N_16786,N_17339);
or U18800 (N_18800,N_16798,N_17933);
and U18801 (N_18801,N_16301,N_17315);
xnor U18802 (N_18802,N_16234,N_16019);
xor U18803 (N_18803,N_16251,N_17179);
or U18804 (N_18804,N_17595,N_17582);
nand U18805 (N_18805,N_16538,N_17158);
nand U18806 (N_18806,N_17913,N_17105);
xnor U18807 (N_18807,N_17305,N_17643);
or U18808 (N_18808,N_17809,N_16420);
nand U18809 (N_18809,N_16031,N_16577);
nand U18810 (N_18810,N_17439,N_16910);
nand U18811 (N_18811,N_17476,N_17526);
and U18812 (N_18812,N_17026,N_16432);
nor U18813 (N_18813,N_17220,N_17888);
and U18814 (N_18814,N_16239,N_16194);
and U18815 (N_18815,N_17244,N_17780);
and U18816 (N_18816,N_16857,N_16374);
nor U18817 (N_18817,N_17711,N_17303);
xnor U18818 (N_18818,N_16338,N_16209);
nand U18819 (N_18819,N_16064,N_16478);
or U18820 (N_18820,N_17036,N_16247);
nand U18821 (N_18821,N_17413,N_17330);
xnor U18822 (N_18822,N_16986,N_17631);
nand U18823 (N_18823,N_17264,N_16257);
nand U18824 (N_18824,N_16370,N_16059);
nor U18825 (N_18825,N_16860,N_17744);
or U18826 (N_18826,N_17092,N_17286);
or U18827 (N_18827,N_16437,N_16142);
nand U18828 (N_18828,N_16984,N_16449);
xor U18829 (N_18829,N_17072,N_17111);
or U18830 (N_18830,N_16106,N_16210);
or U18831 (N_18831,N_17192,N_17344);
nor U18832 (N_18832,N_16994,N_17070);
nand U18833 (N_18833,N_16537,N_17543);
and U18834 (N_18834,N_16479,N_17908);
and U18835 (N_18835,N_17173,N_16947);
nor U18836 (N_18836,N_16826,N_16626);
or U18837 (N_18837,N_16350,N_16229);
nand U18838 (N_18838,N_16638,N_17749);
nor U18839 (N_18839,N_16231,N_16226);
xnor U18840 (N_18840,N_17085,N_16956);
nor U18841 (N_18841,N_16371,N_17802);
nand U18842 (N_18842,N_16191,N_16535);
xnor U18843 (N_18843,N_17869,N_16076);
xnor U18844 (N_18844,N_16023,N_17255);
or U18845 (N_18845,N_17143,N_16861);
nand U18846 (N_18846,N_17382,N_16083);
nand U18847 (N_18847,N_17807,N_17998);
nor U18848 (N_18848,N_17456,N_17754);
or U18849 (N_18849,N_17586,N_17594);
and U18850 (N_18850,N_16790,N_16802);
nor U18851 (N_18851,N_17745,N_17616);
and U18852 (N_18852,N_17118,N_17952);
nor U18853 (N_18853,N_16613,N_17170);
nor U18854 (N_18854,N_16967,N_17522);
or U18855 (N_18855,N_16236,N_16159);
or U18856 (N_18856,N_17682,N_16784);
nand U18857 (N_18857,N_16356,N_16133);
nor U18858 (N_18858,N_17020,N_17886);
nand U18859 (N_18859,N_16590,N_17081);
xor U18860 (N_18860,N_16217,N_16104);
nor U18861 (N_18861,N_17811,N_17149);
or U18862 (N_18862,N_17099,N_17350);
xnor U18863 (N_18863,N_17443,N_16386);
or U18864 (N_18864,N_17728,N_16885);
nor U18865 (N_18865,N_17920,N_16715);
nor U18866 (N_18866,N_16726,N_16949);
nand U18867 (N_18867,N_17408,N_16875);
or U18868 (N_18868,N_16963,N_16615);
nor U18869 (N_18869,N_16269,N_16658);
and U18870 (N_18870,N_16516,N_16129);
nand U18871 (N_18871,N_17883,N_16073);
nand U18872 (N_18872,N_17591,N_16793);
or U18873 (N_18873,N_17784,N_17367);
xnor U18874 (N_18874,N_16215,N_16468);
nand U18875 (N_18875,N_17571,N_17295);
and U18876 (N_18876,N_17717,N_17993);
xnor U18877 (N_18877,N_16380,N_17621);
and U18878 (N_18878,N_17934,N_16833);
xor U18879 (N_18879,N_16747,N_16081);
or U18880 (N_18880,N_16564,N_16092);
or U18881 (N_18881,N_17696,N_16054);
nand U18882 (N_18882,N_17171,N_16346);
nand U18883 (N_18883,N_17040,N_17614);
or U18884 (N_18884,N_16278,N_17097);
or U18885 (N_18885,N_17272,N_17153);
nor U18886 (N_18886,N_17843,N_16205);
xor U18887 (N_18887,N_17715,N_16382);
nand U18888 (N_18888,N_16391,N_16771);
or U18889 (N_18889,N_16664,N_16013);
nor U18890 (N_18890,N_16794,N_17849);
and U18891 (N_18891,N_17229,N_17073);
nand U18892 (N_18892,N_17540,N_17664);
nor U18893 (N_18893,N_16008,N_16218);
nand U18894 (N_18894,N_17990,N_16507);
xnor U18895 (N_18895,N_16527,N_17609);
and U18896 (N_18896,N_16155,N_17502);
nand U18897 (N_18897,N_17516,N_17953);
nor U18898 (N_18898,N_16776,N_17262);
xnor U18899 (N_18899,N_17465,N_17495);
nand U18900 (N_18900,N_16039,N_17190);
nor U18901 (N_18901,N_17885,N_17977);
nand U18902 (N_18902,N_17079,N_17789);
nor U18903 (N_18903,N_16332,N_16834);
nand U18904 (N_18904,N_16127,N_16618);
and U18905 (N_18905,N_17752,N_16445);
and U18906 (N_18906,N_16343,N_16030);
nand U18907 (N_18907,N_16020,N_17896);
nand U18908 (N_18908,N_17716,N_16744);
and U18909 (N_18909,N_17973,N_16429);
or U18910 (N_18910,N_16317,N_17974);
or U18911 (N_18911,N_16759,N_17672);
or U18912 (N_18912,N_16411,N_17248);
nor U18913 (N_18913,N_17121,N_17620);
xor U18914 (N_18914,N_16053,N_17000);
xnor U18915 (N_18915,N_16135,N_17975);
and U18916 (N_18916,N_17098,N_17650);
or U18917 (N_18917,N_16164,N_16748);
and U18918 (N_18918,N_16706,N_16187);
nand U18919 (N_18919,N_16760,N_16851);
or U18920 (N_18920,N_16787,N_17441);
and U18921 (N_18921,N_16731,N_16734);
xor U18922 (N_18922,N_16018,N_16443);
nand U18923 (N_18923,N_16965,N_17713);
or U18924 (N_18924,N_17323,N_16266);
nand U18925 (N_18925,N_17923,N_17655);
and U18926 (N_18926,N_17988,N_17623);
and U18927 (N_18927,N_17790,N_17958);
xor U18928 (N_18928,N_17425,N_16623);
nor U18929 (N_18929,N_17238,N_16606);
nor U18930 (N_18930,N_16801,N_16245);
nand U18931 (N_18931,N_17833,N_17450);
nor U18932 (N_18932,N_17340,N_17454);
and U18933 (N_18933,N_16162,N_17434);
and U18934 (N_18934,N_17384,N_17429);
nand U18935 (N_18935,N_16009,N_16862);
and U18936 (N_18936,N_17638,N_17751);
nor U18937 (N_18937,N_17022,N_16148);
and U18938 (N_18938,N_17504,N_17812);
or U18939 (N_18939,N_16306,N_17252);
or U18940 (N_18940,N_17927,N_17605);
nor U18941 (N_18941,N_16848,N_16708);
nor U18942 (N_18942,N_16646,N_16876);
xor U18943 (N_18943,N_16676,N_17199);
nand U18944 (N_18944,N_16058,N_16816);
and U18945 (N_18945,N_17791,N_16983);
nor U18946 (N_18946,N_16652,N_17492);
xnor U18947 (N_18947,N_16324,N_16682);
nor U18948 (N_18948,N_17864,N_17656);
or U18949 (N_18949,N_17818,N_17635);
xnor U18950 (N_18950,N_17668,N_16206);
or U18951 (N_18951,N_17138,N_17212);
nand U18952 (N_18952,N_17206,N_16898);
or U18953 (N_18953,N_17386,N_17574);
xnor U18954 (N_18954,N_16628,N_16179);
nor U18955 (N_18955,N_16529,N_17116);
nand U18956 (N_18956,N_17921,N_16779);
and U18957 (N_18957,N_17911,N_16912);
nand U18958 (N_18958,N_16273,N_16827);
or U18959 (N_18959,N_17232,N_16394);
and U18960 (N_18960,N_16518,N_17478);
and U18961 (N_18961,N_16151,N_16933);
nor U18962 (N_18962,N_17757,N_17530);
xor U18963 (N_18963,N_16313,N_16732);
nand U18964 (N_18964,N_17561,N_17484);
and U18965 (N_18965,N_16601,N_17996);
nand U18966 (N_18966,N_16200,N_16329);
xor U18967 (N_18967,N_17043,N_16742);
xnor U18968 (N_18968,N_16387,N_17270);
nor U18969 (N_18969,N_17840,N_17966);
or U18970 (N_18970,N_16132,N_17512);
nor U18971 (N_18971,N_16409,N_16534);
nor U18972 (N_18972,N_17748,N_17407);
and U18973 (N_18973,N_17957,N_16131);
xnor U18974 (N_18974,N_16168,N_17223);
and U18975 (N_18975,N_17816,N_17329);
or U18976 (N_18976,N_16713,N_16722);
nor U18977 (N_18977,N_17287,N_17115);
nand U18978 (N_18978,N_16195,N_16836);
or U18979 (N_18979,N_17563,N_17019);
or U18980 (N_18980,N_17409,N_16987);
or U18981 (N_18981,N_17938,N_17706);
and U18982 (N_18982,N_17915,N_17763);
xnor U18983 (N_18983,N_16075,N_16863);
nor U18984 (N_18984,N_17132,N_17761);
nor U18985 (N_18985,N_17613,N_16112);
and U18986 (N_18986,N_17755,N_16656);
nand U18987 (N_18987,N_16091,N_16337);
nand U18988 (N_18988,N_17293,N_17234);
nor U18989 (N_18989,N_17107,N_16560);
and U18990 (N_18990,N_16585,N_17379);
nand U18991 (N_18991,N_16954,N_17587);
nand U18992 (N_18992,N_17080,N_16366);
xor U18993 (N_18993,N_17148,N_16592);
nor U18994 (N_18994,N_17559,N_17168);
nand U18995 (N_18995,N_16193,N_17630);
or U18996 (N_18996,N_16832,N_16867);
and U18997 (N_18997,N_17823,N_16823);
and U18998 (N_18998,N_16174,N_17393);
or U18999 (N_18999,N_16504,N_16841);
and U19000 (N_19000,N_17962,N_16666);
xnor U19001 (N_19001,N_16484,N_17896);
nand U19002 (N_19002,N_16206,N_16560);
nor U19003 (N_19003,N_17029,N_17537);
xnor U19004 (N_19004,N_17260,N_17777);
and U19005 (N_19005,N_17369,N_17353);
xnor U19006 (N_19006,N_16358,N_16756);
xnor U19007 (N_19007,N_17905,N_17254);
xor U19008 (N_19008,N_17660,N_17186);
or U19009 (N_19009,N_17749,N_17924);
nor U19010 (N_19010,N_17027,N_16752);
nand U19011 (N_19011,N_16082,N_17269);
and U19012 (N_19012,N_16485,N_17836);
nand U19013 (N_19013,N_17225,N_16565);
or U19014 (N_19014,N_17373,N_16693);
or U19015 (N_19015,N_16604,N_16091);
xor U19016 (N_19016,N_16581,N_17360);
and U19017 (N_19017,N_17318,N_17082);
or U19018 (N_19018,N_17038,N_17615);
nand U19019 (N_19019,N_16772,N_16902);
nand U19020 (N_19020,N_16699,N_17273);
nor U19021 (N_19021,N_16613,N_16595);
nand U19022 (N_19022,N_16962,N_17821);
and U19023 (N_19023,N_16798,N_17362);
or U19024 (N_19024,N_16038,N_16121);
xnor U19025 (N_19025,N_17596,N_16441);
or U19026 (N_19026,N_16741,N_17185);
nand U19027 (N_19027,N_17774,N_17749);
xor U19028 (N_19028,N_17495,N_17484);
nor U19029 (N_19029,N_16626,N_16674);
and U19030 (N_19030,N_17876,N_17225);
nor U19031 (N_19031,N_16245,N_16736);
nor U19032 (N_19032,N_16684,N_16224);
nand U19033 (N_19033,N_16882,N_17436);
nand U19034 (N_19034,N_16034,N_16587);
or U19035 (N_19035,N_16088,N_17293);
nand U19036 (N_19036,N_16127,N_16773);
xnor U19037 (N_19037,N_16597,N_17193);
xnor U19038 (N_19038,N_17905,N_16027);
nand U19039 (N_19039,N_17742,N_16954);
nand U19040 (N_19040,N_16033,N_16335);
and U19041 (N_19041,N_17344,N_17960);
nand U19042 (N_19042,N_17067,N_17406);
nor U19043 (N_19043,N_17564,N_16294);
xnor U19044 (N_19044,N_17239,N_17612);
nor U19045 (N_19045,N_17950,N_17991);
and U19046 (N_19046,N_16699,N_17659);
nor U19047 (N_19047,N_16828,N_16776);
xnor U19048 (N_19048,N_16124,N_17226);
and U19049 (N_19049,N_16760,N_17225);
xnor U19050 (N_19050,N_17442,N_17732);
nand U19051 (N_19051,N_16279,N_17920);
xor U19052 (N_19052,N_16707,N_17694);
or U19053 (N_19053,N_17130,N_17216);
nor U19054 (N_19054,N_17296,N_16107);
and U19055 (N_19055,N_16426,N_17525);
and U19056 (N_19056,N_17442,N_16727);
or U19057 (N_19057,N_17903,N_17648);
or U19058 (N_19058,N_17451,N_16526);
nand U19059 (N_19059,N_17679,N_16068);
nor U19060 (N_19060,N_17492,N_16493);
or U19061 (N_19061,N_17603,N_16657);
nand U19062 (N_19062,N_17816,N_17656);
xnor U19063 (N_19063,N_17937,N_16071);
or U19064 (N_19064,N_17910,N_16850);
and U19065 (N_19065,N_16989,N_17242);
xnor U19066 (N_19066,N_17243,N_17858);
and U19067 (N_19067,N_16383,N_16648);
nor U19068 (N_19068,N_17544,N_16828);
nand U19069 (N_19069,N_16051,N_16624);
xnor U19070 (N_19070,N_16351,N_17046);
nor U19071 (N_19071,N_17080,N_16901);
nor U19072 (N_19072,N_17527,N_17478);
nor U19073 (N_19073,N_17130,N_17126);
xnor U19074 (N_19074,N_17630,N_17378);
xnor U19075 (N_19075,N_16658,N_17253);
nand U19076 (N_19076,N_16355,N_17084);
nor U19077 (N_19077,N_16700,N_16290);
and U19078 (N_19078,N_17670,N_16679);
and U19079 (N_19079,N_17312,N_17757);
nand U19080 (N_19080,N_16177,N_16924);
and U19081 (N_19081,N_16952,N_16757);
nand U19082 (N_19082,N_17035,N_16769);
or U19083 (N_19083,N_17611,N_17898);
xnor U19084 (N_19084,N_17163,N_16388);
nand U19085 (N_19085,N_17624,N_16845);
nand U19086 (N_19086,N_16165,N_16243);
nor U19087 (N_19087,N_16262,N_17732);
and U19088 (N_19088,N_17457,N_17058);
nand U19089 (N_19089,N_17222,N_16315);
nor U19090 (N_19090,N_17912,N_16817);
xnor U19091 (N_19091,N_16813,N_16570);
or U19092 (N_19092,N_17927,N_16030);
nor U19093 (N_19093,N_16602,N_17244);
nor U19094 (N_19094,N_17630,N_16273);
nor U19095 (N_19095,N_16749,N_17810);
and U19096 (N_19096,N_17819,N_16480);
xor U19097 (N_19097,N_17183,N_16960);
xor U19098 (N_19098,N_17655,N_17323);
or U19099 (N_19099,N_16057,N_16060);
xor U19100 (N_19100,N_17093,N_17223);
nor U19101 (N_19101,N_17654,N_17403);
nor U19102 (N_19102,N_16902,N_17616);
or U19103 (N_19103,N_17015,N_17553);
and U19104 (N_19104,N_17339,N_16736);
nor U19105 (N_19105,N_17111,N_17789);
nand U19106 (N_19106,N_17329,N_17579);
and U19107 (N_19107,N_16524,N_17818);
xnor U19108 (N_19108,N_16727,N_16203);
xor U19109 (N_19109,N_17766,N_17013);
and U19110 (N_19110,N_16545,N_16723);
and U19111 (N_19111,N_16359,N_16149);
nand U19112 (N_19112,N_17820,N_16603);
xnor U19113 (N_19113,N_17540,N_16144);
nand U19114 (N_19114,N_16416,N_16892);
and U19115 (N_19115,N_17901,N_17753);
nor U19116 (N_19116,N_17764,N_16241);
xnor U19117 (N_19117,N_16182,N_17506);
nand U19118 (N_19118,N_17839,N_17557);
and U19119 (N_19119,N_16468,N_17726);
or U19120 (N_19120,N_17575,N_17077);
and U19121 (N_19121,N_17907,N_16583);
nand U19122 (N_19122,N_17083,N_16810);
xnor U19123 (N_19123,N_16126,N_16713);
xnor U19124 (N_19124,N_16272,N_16779);
xnor U19125 (N_19125,N_16855,N_17850);
or U19126 (N_19126,N_17285,N_16274);
nand U19127 (N_19127,N_16215,N_17288);
xnor U19128 (N_19128,N_17708,N_17743);
xor U19129 (N_19129,N_16101,N_16045);
nor U19130 (N_19130,N_17162,N_16730);
and U19131 (N_19131,N_17514,N_16512);
nand U19132 (N_19132,N_16136,N_16832);
nor U19133 (N_19133,N_16250,N_17362);
nand U19134 (N_19134,N_16737,N_17704);
or U19135 (N_19135,N_17800,N_17446);
xnor U19136 (N_19136,N_16984,N_17067);
nor U19137 (N_19137,N_16757,N_17658);
and U19138 (N_19138,N_16831,N_17668);
nand U19139 (N_19139,N_17915,N_16719);
nor U19140 (N_19140,N_17913,N_16366);
or U19141 (N_19141,N_17271,N_16193);
nor U19142 (N_19142,N_16571,N_17057);
or U19143 (N_19143,N_17503,N_16566);
and U19144 (N_19144,N_17052,N_17313);
or U19145 (N_19145,N_16505,N_17714);
or U19146 (N_19146,N_17984,N_17593);
nor U19147 (N_19147,N_17852,N_17619);
or U19148 (N_19148,N_16857,N_16916);
and U19149 (N_19149,N_16968,N_17627);
or U19150 (N_19150,N_17648,N_16924);
or U19151 (N_19151,N_16617,N_17838);
nand U19152 (N_19152,N_17518,N_17592);
xnor U19153 (N_19153,N_17243,N_16414);
and U19154 (N_19154,N_16861,N_17638);
nor U19155 (N_19155,N_17070,N_16843);
or U19156 (N_19156,N_17106,N_17935);
nor U19157 (N_19157,N_17036,N_17903);
and U19158 (N_19158,N_17652,N_17215);
or U19159 (N_19159,N_17597,N_16635);
xor U19160 (N_19160,N_17943,N_17276);
nor U19161 (N_19161,N_17348,N_16135);
or U19162 (N_19162,N_17591,N_16940);
and U19163 (N_19163,N_16504,N_17087);
nand U19164 (N_19164,N_16098,N_17756);
or U19165 (N_19165,N_16330,N_16417);
nor U19166 (N_19166,N_16961,N_17633);
or U19167 (N_19167,N_16409,N_17740);
xnor U19168 (N_19168,N_16923,N_16866);
nor U19169 (N_19169,N_17586,N_16774);
nand U19170 (N_19170,N_16961,N_16846);
nor U19171 (N_19171,N_16281,N_16901);
xnor U19172 (N_19172,N_17257,N_17658);
nand U19173 (N_19173,N_16731,N_17786);
xnor U19174 (N_19174,N_16529,N_17486);
or U19175 (N_19175,N_17778,N_16451);
or U19176 (N_19176,N_17751,N_16230);
xor U19177 (N_19177,N_16735,N_16579);
nor U19178 (N_19178,N_16710,N_17705);
and U19179 (N_19179,N_16057,N_17344);
xnor U19180 (N_19180,N_17579,N_16957);
nor U19181 (N_19181,N_16734,N_17834);
or U19182 (N_19182,N_16403,N_16327);
or U19183 (N_19183,N_16681,N_17630);
nand U19184 (N_19184,N_17285,N_16606);
nand U19185 (N_19185,N_16155,N_17657);
and U19186 (N_19186,N_16087,N_17315);
nand U19187 (N_19187,N_16522,N_16130);
nor U19188 (N_19188,N_16422,N_16328);
nor U19189 (N_19189,N_17652,N_16571);
or U19190 (N_19190,N_16713,N_17016);
nand U19191 (N_19191,N_16486,N_17150);
or U19192 (N_19192,N_16005,N_17077);
nand U19193 (N_19193,N_17892,N_17232);
nor U19194 (N_19194,N_16938,N_17130);
xor U19195 (N_19195,N_17758,N_17262);
and U19196 (N_19196,N_17643,N_16983);
xnor U19197 (N_19197,N_16812,N_17323);
and U19198 (N_19198,N_17524,N_16503);
nor U19199 (N_19199,N_17985,N_17238);
or U19200 (N_19200,N_16913,N_16121);
or U19201 (N_19201,N_16468,N_17056);
xor U19202 (N_19202,N_17099,N_16417);
nor U19203 (N_19203,N_17383,N_16891);
or U19204 (N_19204,N_17177,N_17884);
xnor U19205 (N_19205,N_16250,N_17416);
nand U19206 (N_19206,N_16325,N_17560);
nor U19207 (N_19207,N_16649,N_17746);
or U19208 (N_19208,N_16615,N_16419);
nand U19209 (N_19209,N_16741,N_16655);
nand U19210 (N_19210,N_16301,N_17495);
xor U19211 (N_19211,N_17726,N_16507);
or U19212 (N_19212,N_16444,N_17344);
nand U19213 (N_19213,N_16617,N_17262);
or U19214 (N_19214,N_17051,N_16950);
or U19215 (N_19215,N_17436,N_16877);
xnor U19216 (N_19216,N_17844,N_17692);
or U19217 (N_19217,N_16500,N_16595);
or U19218 (N_19218,N_16568,N_16335);
nor U19219 (N_19219,N_16660,N_16689);
nor U19220 (N_19220,N_17911,N_16911);
xor U19221 (N_19221,N_17496,N_16291);
xnor U19222 (N_19222,N_17016,N_17863);
nand U19223 (N_19223,N_17837,N_16278);
nand U19224 (N_19224,N_16246,N_17345);
nor U19225 (N_19225,N_17256,N_17424);
xor U19226 (N_19226,N_16968,N_17863);
nor U19227 (N_19227,N_17006,N_16032);
nand U19228 (N_19228,N_16135,N_16972);
and U19229 (N_19229,N_16717,N_16539);
or U19230 (N_19230,N_17920,N_16567);
xor U19231 (N_19231,N_16527,N_16283);
or U19232 (N_19232,N_17802,N_16863);
nor U19233 (N_19233,N_17703,N_17371);
or U19234 (N_19234,N_16602,N_16243);
xnor U19235 (N_19235,N_17571,N_16116);
nor U19236 (N_19236,N_17150,N_16595);
and U19237 (N_19237,N_17677,N_16131);
or U19238 (N_19238,N_17676,N_16594);
nand U19239 (N_19239,N_17501,N_17471);
nand U19240 (N_19240,N_16130,N_17747);
and U19241 (N_19241,N_16052,N_16214);
and U19242 (N_19242,N_17124,N_16394);
nand U19243 (N_19243,N_17607,N_16961);
or U19244 (N_19244,N_16258,N_16120);
nor U19245 (N_19245,N_16988,N_17998);
and U19246 (N_19246,N_16215,N_16418);
xnor U19247 (N_19247,N_17651,N_17262);
and U19248 (N_19248,N_16835,N_16381);
and U19249 (N_19249,N_17122,N_16168);
nor U19250 (N_19250,N_16591,N_16623);
and U19251 (N_19251,N_17393,N_17012);
or U19252 (N_19252,N_16730,N_16520);
nand U19253 (N_19253,N_16898,N_16529);
xnor U19254 (N_19254,N_17450,N_17704);
nand U19255 (N_19255,N_17174,N_17097);
nor U19256 (N_19256,N_17346,N_16295);
nor U19257 (N_19257,N_17543,N_16528);
nor U19258 (N_19258,N_16352,N_16800);
nor U19259 (N_19259,N_16815,N_17312);
or U19260 (N_19260,N_16346,N_16977);
or U19261 (N_19261,N_17606,N_16030);
nor U19262 (N_19262,N_17639,N_17477);
nand U19263 (N_19263,N_16005,N_17134);
or U19264 (N_19264,N_16636,N_16256);
xnor U19265 (N_19265,N_17088,N_16757);
nand U19266 (N_19266,N_17803,N_16414);
xnor U19267 (N_19267,N_16271,N_17979);
and U19268 (N_19268,N_16058,N_16617);
or U19269 (N_19269,N_17293,N_17763);
and U19270 (N_19270,N_16473,N_17013);
xor U19271 (N_19271,N_16087,N_17716);
or U19272 (N_19272,N_16113,N_17131);
nand U19273 (N_19273,N_17091,N_17731);
nor U19274 (N_19274,N_16923,N_16432);
or U19275 (N_19275,N_17244,N_17716);
or U19276 (N_19276,N_17340,N_17730);
xor U19277 (N_19277,N_17953,N_16578);
or U19278 (N_19278,N_17695,N_16717);
nor U19279 (N_19279,N_17475,N_16729);
nand U19280 (N_19280,N_16408,N_16062);
and U19281 (N_19281,N_16151,N_17016);
or U19282 (N_19282,N_16928,N_16134);
xor U19283 (N_19283,N_17401,N_16609);
nor U19284 (N_19284,N_17346,N_17962);
nand U19285 (N_19285,N_16450,N_16843);
nor U19286 (N_19286,N_16781,N_16307);
nor U19287 (N_19287,N_16381,N_16014);
and U19288 (N_19288,N_17749,N_16130);
nand U19289 (N_19289,N_17170,N_17847);
nand U19290 (N_19290,N_16157,N_16262);
or U19291 (N_19291,N_17469,N_17123);
and U19292 (N_19292,N_17487,N_17750);
nand U19293 (N_19293,N_17582,N_16079);
or U19294 (N_19294,N_17093,N_17065);
nand U19295 (N_19295,N_16399,N_16477);
xor U19296 (N_19296,N_17524,N_16929);
xor U19297 (N_19297,N_17490,N_17535);
nand U19298 (N_19298,N_16134,N_17826);
xnor U19299 (N_19299,N_17346,N_17979);
nand U19300 (N_19300,N_17593,N_17361);
and U19301 (N_19301,N_16168,N_17351);
or U19302 (N_19302,N_16304,N_17133);
nand U19303 (N_19303,N_17183,N_17292);
and U19304 (N_19304,N_16308,N_17811);
nor U19305 (N_19305,N_17345,N_17471);
and U19306 (N_19306,N_16028,N_16508);
and U19307 (N_19307,N_16817,N_17153);
nand U19308 (N_19308,N_16611,N_16671);
nor U19309 (N_19309,N_16108,N_16229);
or U19310 (N_19310,N_16638,N_17569);
or U19311 (N_19311,N_16126,N_16262);
nor U19312 (N_19312,N_16242,N_16529);
or U19313 (N_19313,N_17314,N_17899);
xnor U19314 (N_19314,N_17005,N_17877);
and U19315 (N_19315,N_16074,N_16488);
nor U19316 (N_19316,N_16529,N_17280);
or U19317 (N_19317,N_16920,N_17475);
nand U19318 (N_19318,N_16751,N_16822);
or U19319 (N_19319,N_16080,N_17581);
xor U19320 (N_19320,N_16003,N_17976);
and U19321 (N_19321,N_17102,N_16719);
or U19322 (N_19322,N_17714,N_16975);
or U19323 (N_19323,N_17033,N_16513);
nor U19324 (N_19324,N_17752,N_16058);
nor U19325 (N_19325,N_16044,N_16095);
nor U19326 (N_19326,N_17062,N_17735);
nor U19327 (N_19327,N_16047,N_16811);
xnor U19328 (N_19328,N_16156,N_17438);
nand U19329 (N_19329,N_16104,N_17296);
xnor U19330 (N_19330,N_16091,N_16879);
nor U19331 (N_19331,N_17868,N_16606);
nor U19332 (N_19332,N_16718,N_17519);
and U19333 (N_19333,N_17828,N_16857);
nand U19334 (N_19334,N_17134,N_16632);
or U19335 (N_19335,N_16235,N_17476);
and U19336 (N_19336,N_17801,N_16788);
and U19337 (N_19337,N_16984,N_16346);
xnor U19338 (N_19338,N_17587,N_17259);
nor U19339 (N_19339,N_17970,N_17362);
nand U19340 (N_19340,N_17556,N_17988);
xnor U19341 (N_19341,N_17882,N_16561);
or U19342 (N_19342,N_16228,N_16768);
nand U19343 (N_19343,N_17631,N_17493);
and U19344 (N_19344,N_17692,N_17069);
nand U19345 (N_19345,N_16424,N_17675);
nand U19346 (N_19346,N_17383,N_16211);
or U19347 (N_19347,N_17550,N_16140);
nor U19348 (N_19348,N_16847,N_17119);
xor U19349 (N_19349,N_17044,N_17004);
or U19350 (N_19350,N_16704,N_16781);
and U19351 (N_19351,N_16808,N_17406);
xnor U19352 (N_19352,N_17083,N_17130);
and U19353 (N_19353,N_16137,N_16294);
and U19354 (N_19354,N_17593,N_17119);
nand U19355 (N_19355,N_16742,N_16951);
or U19356 (N_19356,N_16757,N_17835);
and U19357 (N_19357,N_16807,N_17336);
or U19358 (N_19358,N_17802,N_17432);
nand U19359 (N_19359,N_16851,N_16622);
and U19360 (N_19360,N_17983,N_17761);
nand U19361 (N_19361,N_17646,N_16803);
and U19362 (N_19362,N_16061,N_17831);
and U19363 (N_19363,N_17093,N_17893);
nor U19364 (N_19364,N_16210,N_16861);
nor U19365 (N_19365,N_16026,N_16699);
and U19366 (N_19366,N_16281,N_16848);
or U19367 (N_19367,N_17227,N_16024);
nor U19368 (N_19368,N_17561,N_16755);
xnor U19369 (N_19369,N_17429,N_17300);
nand U19370 (N_19370,N_16240,N_17150);
nor U19371 (N_19371,N_16995,N_17057);
or U19372 (N_19372,N_17956,N_17920);
or U19373 (N_19373,N_17903,N_16390);
or U19374 (N_19374,N_17579,N_17897);
nand U19375 (N_19375,N_16155,N_17344);
and U19376 (N_19376,N_16536,N_16115);
or U19377 (N_19377,N_17742,N_16028);
nor U19378 (N_19378,N_16651,N_16548);
and U19379 (N_19379,N_16888,N_16168);
or U19380 (N_19380,N_16171,N_16871);
or U19381 (N_19381,N_16060,N_16510);
nor U19382 (N_19382,N_17410,N_16339);
or U19383 (N_19383,N_16817,N_17301);
nor U19384 (N_19384,N_16732,N_17837);
and U19385 (N_19385,N_17530,N_16942);
or U19386 (N_19386,N_16787,N_16539);
nor U19387 (N_19387,N_16075,N_16239);
and U19388 (N_19388,N_16010,N_16384);
nand U19389 (N_19389,N_16385,N_17369);
xnor U19390 (N_19390,N_16454,N_17384);
nor U19391 (N_19391,N_16927,N_16881);
nor U19392 (N_19392,N_16918,N_17849);
nand U19393 (N_19393,N_16242,N_16695);
and U19394 (N_19394,N_16574,N_17384);
nor U19395 (N_19395,N_17898,N_17025);
nor U19396 (N_19396,N_17186,N_16143);
or U19397 (N_19397,N_16290,N_17075);
xnor U19398 (N_19398,N_16934,N_16354);
xor U19399 (N_19399,N_16364,N_17950);
nand U19400 (N_19400,N_17095,N_17214);
nand U19401 (N_19401,N_17990,N_17827);
nor U19402 (N_19402,N_16217,N_17387);
xor U19403 (N_19403,N_16278,N_17747);
and U19404 (N_19404,N_17152,N_16226);
xor U19405 (N_19405,N_17855,N_17767);
nand U19406 (N_19406,N_17010,N_16693);
xnor U19407 (N_19407,N_16936,N_16329);
xor U19408 (N_19408,N_16842,N_16391);
or U19409 (N_19409,N_16480,N_16370);
nor U19410 (N_19410,N_17065,N_17236);
or U19411 (N_19411,N_16240,N_16225);
nand U19412 (N_19412,N_16990,N_16705);
nor U19413 (N_19413,N_17432,N_17024);
nand U19414 (N_19414,N_17893,N_17962);
nor U19415 (N_19415,N_16936,N_17103);
xor U19416 (N_19416,N_16477,N_17351);
nor U19417 (N_19417,N_17166,N_17836);
nand U19418 (N_19418,N_17419,N_17281);
and U19419 (N_19419,N_17670,N_16802);
nor U19420 (N_19420,N_16021,N_17554);
or U19421 (N_19421,N_17257,N_17742);
nand U19422 (N_19422,N_16718,N_17970);
nand U19423 (N_19423,N_17208,N_16042);
nand U19424 (N_19424,N_16856,N_16225);
and U19425 (N_19425,N_16475,N_16853);
or U19426 (N_19426,N_16148,N_16266);
and U19427 (N_19427,N_16938,N_17042);
xor U19428 (N_19428,N_17940,N_16343);
nand U19429 (N_19429,N_16102,N_17177);
and U19430 (N_19430,N_17323,N_16119);
xnor U19431 (N_19431,N_17872,N_17178);
xor U19432 (N_19432,N_16299,N_16283);
or U19433 (N_19433,N_16012,N_17304);
nand U19434 (N_19434,N_16354,N_16229);
xnor U19435 (N_19435,N_16463,N_16567);
xor U19436 (N_19436,N_16492,N_16604);
xor U19437 (N_19437,N_16523,N_17578);
nand U19438 (N_19438,N_17641,N_16159);
xnor U19439 (N_19439,N_16673,N_16932);
xnor U19440 (N_19440,N_17853,N_16092);
and U19441 (N_19441,N_17482,N_17532);
xnor U19442 (N_19442,N_17838,N_17073);
nand U19443 (N_19443,N_17016,N_17486);
or U19444 (N_19444,N_17620,N_17565);
nor U19445 (N_19445,N_16502,N_17962);
xnor U19446 (N_19446,N_17710,N_16084);
and U19447 (N_19447,N_16850,N_16293);
and U19448 (N_19448,N_17156,N_17130);
nor U19449 (N_19449,N_16389,N_16502);
and U19450 (N_19450,N_17821,N_16717);
xor U19451 (N_19451,N_17190,N_17506);
and U19452 (N_19452,N_17705,N_16549);
or U19453 (N_19453,N_17851,N_17651);
nor U19454 (N_19454,N_17651,N_16563);
nand U19455 (N_19455,N_16231,N_16328);
or U19456 (N_19456,N_16174,N_17237);
xnor U19457 (N_19457,N_16164,N_16872);
xor U19458 (N_19458,N_17778,N_16963);
nand U19459 (N_19459,N_17221,N_16871);
nand U19460 (N_19460,N_17460,N_16533);
and U19461 (N_19461,N_17188,N_17143);
and U19462 (N_19462,N_17521,N_16417);
and U19463 (N_19463,N_17117,N_17751);
or U19464 (N_19464,N_16293,N_17399);
xnor U19465 (N_19465,N_16726,N_17820);
nand U19466 (N_19466,N_17001,N_16824);
nand U19467 (N_19467,N_17111,N_17246);
nand U19468 (N_19468,N_16566,N_17938);
nor U19469 (N_19469,N_16170,N_17202);
nor U19470 (N_19470,N_16299,N_16712);
and U19471 (N_19471,N_17032,N_17049);
or U19472 (N_19472,N_16983,N_16434);
xnor U19473 (N_19473,N_16877,N_16819);
xor U19474 (N_19474,N_17176,N_17665);
and U19475 (N_19475,N_16039,N_17998);
and U19476 (N_19476,N_16229,N_16188);
xor U19477 (N_19477,N_17682,N_16439);
nor U19478 (N_19478,N_16063,N_17861);
and U19479 (N_19479,N_16294,N_17381);
nor U19480 (N_19480,N_17977,N_16539);
nor U19481 (N_19481,N_16048,N_16834);
or U19482 (N_19482,N_16723,N_16334);
nand U19483 (N_19483,N_16776,N_16866);
and U19484 (N_19484,N_16075,N_17037);
and U19485 (N_19485,N_17028,N_16832);
or U19486 (N_19486,N_16440,N_16505);
nand U19487 (N_19487,N_17838,N_16661);
nor U19488 (N_19488,N_17014,N_16014);
and U19489 (N_19489,N_16764,N_16589);
xnor U19490 (N_19490,N_17954,N_17642);
nor U19491 (N_19491,N_17153,N_16853);
nor U19492 (N_19492,N_16904,N_17161);
and U19493 (N_19493,N_17593,N_17229);
nor U19494 (N_19494,N_17676,N_17947);
xor U19495 (N_19495,N_16106,N_16150);
xnor U19496 (N_19496,N_17215,N_16001);
xnor U19497 (N_19497,N_17558,N_16743);
or U19498 (N_19498,N_17840,N_17894);
or U19499 (N_19499,N_16991,N_16046);
and U19500 (N_19500,N_16539,N_17495);
or U19501 (N_19501,N_16681,N_16176);
nor U19502 (N_19502,N_17100,N_16005);
nor U19503 (N_19503,N_17266,N_17980);
xor U19504 (N_19504,N_16774,N_17243);
xor U19505 (N_19505,N_16234,N_16439);
nor U19506 (N_19506,N_17688,N_16638);
and U19507 (N_19507,N_17921,N_16307);
nand U19508 (N_19508,N_16863,N_17761);
or U19509 (N_19509,N_16730,N_17403);
nand U19510 (N_19510,N_17689,N_17137);
and U19511 (N_19511,N_17563,N_16202);
nand U19512 (N_19512,N_16597,N_16717);
xnor U19513 (N_19513,N_17680,N_16505);
nand U19514 (N_19514,N_16707,N_17407);
nor U19515 (N_19515,N_17890,N_17614);
and U19516 (N_19516,N_17831,N_16247);
and U19517 (N_19517,N_16351,N_16812);
nand U19518 (N_19518,N_17870,N_17658);
nand U19519 (N_19519,N_17447,N_17987);
and U19520 (N_19520,N_17636,N_16223);
and U19521 (N_19521,N_16006,N_16635);
or U19522 (N_19522,N_17292,N_16900);
nor U19523 (N_19523,N_16641,N_17107);
nor U19524 (N_19524,N_16497,N_17020);
or U19525 (N_19525,N_16314,N_16679);
and U19526 (N_19526,N_16693,N_17744);
and U19527 (N_19527,N_17656,N_16436);
and U19528 (N_19528,N_17761,N_16664);
xor U19529 (N_19529,N_16341,N_17653);
or U19530 (N_19530,N_17997,N_17184);
xnor U19531 (N_19531,N_17397,N_17227);
or U19532 (N_19532,N_16828,N_17273);
nand U19533 (N_19533,N_16716,N_17742);
and U19534 (N_19534,N_17849,N_16096);
xor U19535 (N_19535,N_16669,N_17651);
and U19536 (N_19536,N_17386,N_16742);
or U19537 (N_19537,N_16848,N_17706);
and U19538 (N_19538,N_16934,N_17159);
and U19539 (N_19539,N_16508,N_16034);
or U19540 (N_19540,N_16316,N_16091);
nand U19541 (N_19541,N_17468,N_16024);
or U19542 (N_19542,N_17245,N_16065);
and U19543 (N_19543,N_16155,N_17092);
nor U19544 (N_19544,N_17792,N_16358);
or U19545 (N_19545,N_16346,N_16430);
nor U19546 (N_19546,N_16468,N_16145);
and U19547 (N_19547,N_16018,N_16279);
xnor U19548 (N_19548,N_17897,N_17665);
or U19549 (N_19549,N_16513,N_17111);
xnor U19550 (N_19550,N_17468,N_16026);
xnor U19551 (N_19551,N_16016,N_17933);
xor U19552 (N_19552,N_16747,N_16559);
nand U19553 (N_19553,N_17819,N_16302);
xor U19554 (N_19554,N_16297,N_16686);
xor U19555 (N_19555,N_16043,N_17344);
and U19556 (N_19556,N_16468,N_17944);
and U19557 (N_19557,N_17153,N_17642);
nor U19558 (N_19558,N_17179,N_16531);
xor U19559 (N_19559,N_17081,N_16335);
xnor U19560 (N_19560,N_17035,N_17822);
nor U19561 (N_19561,N_17066,N_17831);
nor U19562 (N_19562,N_16546,N_16484);
or U19563 (N_19563,N_17115,N_17624);
or U19564 (N_19564,N_16109,N_17934);
xnor U19565 (N_19565,N_17679,N_16080);
nand U19566 (N_19566,N_17860,N_17986);
nand U19567 (N_19567,N_16119,N_17223);
xnor U19568 (N_19568,N_17424,N_16598);
and U19569 (N_19569,N_16891,N_17805);
nand U19570 (N_19570,N_17515,N_16338);
xor U19571 (N_19571,N_16240,N_17798);
or U19572 (N_19572,N_16629,N_16019);
xnor U19573 (N_19573,N_16403,N_16471);
nor U19574 (N_19574,N_17233,N_16480);
and U19575 (N_19575,N_17698,N_16886);
and U19576 (N_19576,N_17439,N_16786);
and U19577 (N_19577,N_16098,N_17586);
or U19578 (N_19578,N_17587,N_16193);
xnor U19579 (N_19579,N_16285,N_16003);
nor U19580 (N_19580,N_16867,N_16583);
nand U19581 (N_19581,N_16071,N_17992);
xor U19582 (N_19582,N_17594,N_17993);
and U19583 (N_19583,N_16260,N_17782);
nor U19584 (N_19584,N_16219,N_17480);
nor U19585 (N_19585,N_16379,N_17800);
and U19586 (N_19586,N_16311,N_16367);
nand U19587 (N_19587,N_17390,N_16905);
xor U19588 (N_19588,N_17744,N_17021);
and U19589 (N_19589,N_17262,N_16334);
xor U19590 (N_19590,N_16602,N_17126);
and U19591 (N_19591,N_17357,N_17928);
nor U19592 (N_19592,N_16088,N_16768);
xnor U19593 (N_19593,N_17316,N_17196);
nor U19594 (N_19594,N_16986,N_17087);
xor U19595 (N_19595,N_17142,N_16814);
nand U19596 (N_19596,N_16145,N_17037);
and U19597 (N_19597,N_16115,N_17233);
nor U19598 (N_19598,N_17197,N_16802);
xnor U19599 (N_19599,N_17476,N_17617);
or U19600 (N_19600,N_17754,N_16444);
and U19601 (N_19601,N_16127,N_17828);
or U19602 (N_19602,N_16650,N_17174);
xor U19603 (N_19603,N_16106,N_16941);
nor U19604 (N_19604,N_16330,N_16226);
nor U19605 (N_19605,N_16690,N_16586);
and U19606 (N_19606,N_16413,N_17884);
nand U19607 (N_19607,N_17842,N_16808);
and U19608 (N_19608,N_17155,N_16577);
nor U19609 (N_19609,N_17715,N_16388);
nand U19610 (N_19610,N_17086,N_16298);
nand U19611 (N_19611,N_16581,N_17367);
nand U19612 (N_19612,N_17499,N_16684);
or U19613 (N_19613,N_17883,N_17510);
or U19614 (N_19614,N_16700,N_17454);
xor U19615 (N_19615,N_16414,N_17469);
or U19616 (N_19616,N_17545,N_16449);
and U19617 (N_19617,N_17871,N_17980);
nor U19618 (N_19618,N_17710,N_17556);
or U19619 (N_19619,N_17775,N_16561);
nor U19620 (N_19620,N_17903,N_17597);
nor U19621 (N_19621,N_17450,N_16045);
nand U19622 (N_19622,N_16798,N_16796);
and U19623 (N_19623,N_17115,N_16085);
or U19624 (N_19624,N_16352,N_17758);
or U19625 (N_19625,N_17054,N_17359);
nor U19626 (N_19626,N_17878,N_16824);
or U19627 (N_19627,N_16211,N_16655);
and U19628 (N_19628,N_17539,N_17295);
or U19629 (N_19629,N_17271,N_17114);
xor U19630 (N_19630,N_17735,N_17848);
nand U19631 (N_19631,N_17391,N_16196);
or U19632 (N_19632,N_16489,N_16783);
xor U19633 (N_19633,N_16571,N_16638);
and U19634 (N_19634,N_16081,N_17439);
nand U19635 (N_19635,N_17061,N_16347);
or U19636 (N_19636,N_17122,N_16590);
and U19637 (N_19637,N_16126,N_16933);
nor U19638 (N_19638,N_16708,N_17592);
nor U19639 (N_19639,N_16985,N_16289);
or U19640 (N_19640,N_17181,N_16166);
or U19641 (N_19641,N_17502,N_16799);
nand U19642 (N_19642,N_17526,N_17653);
nand U19643 (N_19643,N_16298,N_16162);
nand U19644 (N_19644,N_16945,N_16147);
and U19645 (N_19645,N_17751,N_16706);
and U19646 (N_19646,N_17254,N_17104);
xor U19647 (N_19647,N_17823,N_16093);
and U19648 (N_19648,N_17115,N_16847);
nor U19649 (N_19649,N_16854,N_16558);
nand U19650 (N_19650,N_16361,N_17354);
and U19651 (N_19651,N_17643,N_17961);
or U19652 (N_19652,N_17601,N_16244);
xor U19653 (N_19653,N_17163,N_16056);
xor U19654 (N_19654,N_16169,N_17422);
xnor U19655 (N_19655,N_17652,N_16537);
nor U19656 (N_19656,N_16462,N_16032);
xnor U19657 (N_19657,N_17354,N_16652);
nor U19658 (N_19658,N_17097,N_17821);
and U19659 (N_19659,N_16764,N_16117);
nand U19660 (N_19660,N_17369,N_16357);
nor U19661 (N_19661,N_17225,N_17475);
nand U19662 (N_19662,N_17761,N_17229);
nor U19663 (N_19663,N_16420,N_17179);
or U19664 (N_19664,N_17445,N_17605);
xor U19665 (N_19665,N_17651,N_17585);
or U19666 (N_19666,N_16207,N_16867);
and U19667 (N_19667,N_16431,N_16684);
xor U19668 (N_19668,N_16136,N_16208);
xnor U19669 (N_19669,N_17555,N_16176);
xor U19670 (N_19670,N_17547,N_16736);
and U19671 (N_19671,N_16241,N_17119);
xnor U19672 (N_19672,N_16422,N_17011);
nor U19673 (N_19673,N_17881,N_16449);
nand U19674 (N_19674,N_16891,N_17345);
or U19675 (N_19675,N_17869,N_17576);
nor U19676 (N_19676,N_17376,N_16129);
nand U19677 (N_19677,N_16740,N_17856);
or U19678 (N_19678,N_17607,N_17632);
and U19679 (N_19679,N_17153,N_17483);
nor U19680 (N_19680,N_16792,N_17088);
xnor U19681 (N_19681,N_16828,N_17515);
and U19682 (N_19682,N_16010,N_17257);
nor U19683 (N_19683,N_16295,N_16117);
and U19684 (N_19684,N_17006,N_17930);
or U19685 (N_19685,N_17484,N_16409);
and U19686 (N_19686,N_17900,N_16498);
nor U19687 (N_19687,N_16419,N_17821);
xor U19688 (N_19688,N_17430,N_16405);
xnor U19689 (N_19689,N_17650,N_16645);
and U19690 (N_19690,N_17675,N_16761);
and U19691 (N_19691,N_16434,N_16948);
nand U19692 (N_19692,N_17410,N_16560);
nand U19693 (N_19693,N_17683,N_16045);
xor U19694 (N_19694,N_17625,N_16390);
or U19695 (N_19695,N_16469,N_16143);
nor U19696 (N_19696,N_17162,N_17722);
nand U19697 (N_19697,N_16245,N_16617);
xnor U19698 (N_19698,N_17022,N_16407);
or U19699 (N_19699,N_16644,N_16345);
and U19700 (N_19700,N_16441,N_17872);
or U19701 (N_19701,N_17899,N_17686);
nand U19702 (N_19702,N_16673,N_17932);
or U19703 (N_19703,N_16325,N_16811);
nand U19704 (N_19704,N_17213,N_16139);
and U19705 (N_19705,N_17057,N_17625);
and U19706 (N_19706,N_17955,N_17663);
xnor U19707 (N_19707,N_16308,N_16686);
and U19708 (N_19708,N_17777,N_17395);
or U19709 (N_19709,N_16032,N_16563);
nand U19710 (N_19710,N_16489,N_16374);
or U19711 (N_19711,N_17068,N_17153);
or U19712 (N_19712,N_16088,N_17717);
or U19713 (N_19713,N_17766,N_16360);
and U19714 (N_19714,N_16636,N_17355);
xor U19715 (N_19715,N_16168,N_17978);
and U19716 (N_19716,N_16774,N_16464);
nand U19717 (N_19717,N_17797,N_17121);
and U19718 (N_19718,N_16069,N_16802);
xnor U19719 (N_19719,N_17975,N_17288);
or U19720 (N_19720,N_16478,N_17372);
nor U19721 (N_19721,N_16249,N_17649);
nand U19722 (N_19722,N_16896,N_16034);
and U19723 (N_19723,N_17631,N_16279);
xor U19724 (N_19724,N_16074,N_17285);
and U19725 (N_19725,N_17990,N_16048);
nor U19726 (N_19726,N_16923,N_16162);
nor U19727 (N_19727,N_17676,N_16209);
nand U19728 (N_19728,N_16730,N_17678);
xnor U19729 (N_19729,N_16342,N_17216);
xnor U19730 (N_19730,N_17707,N_16308);
xnor U19731 (N_19731,N_17566,N_16136);
or U19732 (N_19732,N_16586,N_17840);
xnor U19733 (N_19733,N_16209,N_16208);
and U19734 (N_19734,N_17960,N_16953);
xnor U19735 (N_19735,N_17911,N_16371);
nor U19736 (N_19736,N_17483,N_17437);
nand U19737 (N_19737,N_17891,N_16328);
or U19738 (N_19738,N_16271,N_16403);
and U19739 (N_19739,N_17902,N_17335);
and U19740 (N_19740,N_16685,N_17224);
nor U19741 (N_19741,N_16979,N_16744);
nor U19742 (N_19742,N_17105,N_16480);
nor U19743 (N_19743,N_16762,N_17384);
xor U19744 (N_19744,N_16797,N_16257);
nor U19745 (N_19745,N_16877,N_17941);
nor U19746 (N_19746,N_17346,N_16485);
or U19747 (N_19747,N_17261,N_16047);
and U19748 (N_19748,N_17941,N_17844);
xor U19749 (N_19749,N_17314,N_17016);
nand U19750 (N_19750,N_16985,N_17096);
nand U19751 (N_19751,N_17801,N_17918);
xor U19752 (N_19752,N_17646,N_17554);
xor U19753 (N_19753,N_17888,N_16054);
or U19754 (N_19754,N_16931,N_17822);
nor U19755 (N_19755,N_16331,N_16530);
nand U19756 (N_19756,N_17332,N_16043);
xor U19757 (N_19757,N_16094,N_17601);
or U19758 (N_19758,N_17570,N_16683);
nand U19759 (N_19759,N_17949,N_16844);
and U19760 (N_19760,N_17725,N_16782);
xor U19761 (N_19761,N_17113,N_16640);
xor U19762 (N_19762,N_17099,N_16380);
nor U19763 (N_19763,N_16871,N_17905);
or U19764 (N_19764,N_17078,N_16679);
nand U19765 (N_19765,N_17864,N_16698);
and U19766 (N_19766,N_16276,N_16885);
nand U19767 (N_19767,N_16167,N_17734);
xor U19768 (N_19768,N_17486,N_16230);
nor U19769 (N_19769,N_16123,N_16369);
or U19770 (N_19770,N_17796,N_16035);
xnor U19771 (N_19771,N_17603,N_17449);
and U19772 (N_19772,N_17355,N_17466);
xor U19773 (N_19773,N_17004,N_16515);
nor U19774 (N_19774,N_17808,N_16046);
xor U19775 (N_19775,N_16526,N_17268);
or U19776 (N_19776,N_16176,N_17254);
and U19777 (N_19777,N_16842,N_16323);
nand U19778 (N_19778,N_16252,N_17189);
nand U19779 (N_19779,N_17020,N_17807);
nand U19780 (N_19780,N_16520,N_17204);
nor U19781 (N_19781,N_16685,N_16927);
nor U19782 (N_19782,N_17213,N_17614);
nand U19783 (N_19783,N_17676,N_17481);
or U19784 (N_19784,N_16115,N_16153);
nor U19785 (N_19785,N_17157,N_16450);
or U19786 (N_19786,N_16964,N_16739);
xor U19787 (N_19787,N_16168,N_16926);
xor U19788 (N_19788,N_17151,N_16944);
and U19789 (N_19789,N_17025,N_16672);
xor U19790 (N_19790,N_16625,N_16980);
xnor U19791 (N_19791,N_16081,N_17659);
and U19792 (N_19792,N_17953,N_16488);
nor U19793 (N_19793,N_16055,N_16135);
xor U19794 (N_19794,N_16689,N_16597);
nor U19795 (N_19795,N_17521,N_17213);
xnor U19796 (N_19796,N_16927,N_16314);
and U19797 (N_19797,N_16904,N_16968);
nand U19798 (N_19798,N_16654,N_17128);
nand U19799 (N_19799,N_16224,N_17241);
xnor U19800 (N_19800,N_17537,N_17100);
nand U19801 (N_19801,N_17414,N_17450);
nand U19802 (N_19802,N_17676,N_17732);
xnor U19803 (N_19803,N_17459,N_17997);
or U19804 (N_19804,N_16019,N_17921);
or U19805 (N_19805,N_17222,N_16027);
and U19806 (N_19806,N_17830,N_17462);
xor U19807 (N_19807,N_16663,N_17034);
nor U19808 (N_19808,N_16055,N_17486);
or U19809 (N_19809,N_17148,N_17625);
nand U19810 (N_19810,N_17496,N_17309);
nand U19811 (N_19811,N_16764,N_17497);
xor U19812 (N_19812,N_17571,N_17512);
nand U19813 (N_19813,N_17889,N_17177);
xor U19814 (N_19814,N_16622,N_16561);
nor U19815 (N_19815,N_17112,N_16250);
xor U19816 (N_19816,N_16814,N_16149);
xor U19817 (N_19817,N_16701,N_17657);
nand U19818 (N_19818,N_16802,N_17980);
and U19819 (N_19819,N_16593,N_16807);
nand U19820 (N_19820,N_17262,N_16231);
nor U19821 (N_19821,N_17260,N_16694);
xnor U19822 (N_19822,N_17184,N_17620);
nor U19823 (N_19823,N_17450,N_16428);
nand U19824 (N_19824,N_16252,N_17035);
or U19825 (N_19825,N_16744,N_16279);
or U19826 (N_19826,N_17246,N_17605);
nand U19827 (N_19827,N_16913,N_16634);
nand U19828 (N_19828,N_16711,N_16772);
and U19829 (N_19829,N_17457,N_17268);
or U19830 (N_19830,N_17987,N_17497);
and U19831 (N_19831,N_17750,N_17491);
nor U19832 (N_19832,N_17176,N_17858);
nor U19833 (N_19833,N_17152,N_17290);
or U19834 (N_19834,N_16280,N_16144);
and U19835 (N_19835,N_16445,N_17148);
and U19836 (N_19836,N_17913,N_17137);
nor U19837 (N_19837,N_17212,N_16218);
nor U19838 (N_19838,N_17052,N_17053);
xnor U19839 (N_19839,N_17750,N_16838);
or U19840 (N_19840,N_17051,N_16611);
xnor U19841 (N_19841,N_17054,N_17013);
xor U19842 (N_19842,N_16011,N_16863);
and U19843 (N_19843,N_16354,N_17865);
nand U19844 (N_19844,N_17532,N_16992);
nor U19845 (N_19845,N_17070,N_17322);
xor U19846 (N_19846,N_16836,N_16849);
nor U19847 (N_19847,N_17058,N_16613);
nor U19848 (N_19848,N_16903,N_17186);
or U19849 (N_19849,N_16760,N_16940);
or U19850 (N_19850,N_16002,N_16567);
nand U19851 (N_19851,N_16762,N_17375);
nand U19852 (N_19852,N_16824,N_16358);
xor U19853 (N_19853,N_16146,N_16684);
xor U19854 (N_19854,N_16825,N_17571);
nor U19855 (N_19855,N_17688,N_16406);
nor U19856 (N_19856,N_17124,N_16111);
nor U19857 (N_19857,N_17884,N_16898);
and U19858 (N_19858,N_16696,N_17985);
and U19859 (N_19859,N_16973,N_17540);
xnor U19860 (N_19860,N_17510,N_16852);
or U19861 (N_19861,N_17357,N_17878);
or U19862 (N_19862,N_16918,N_17300);
and U19863 (N_19863,N_16655,N_16278);
nand U19864 (N_19864,N_16370,N_17157);
nand U19865 (N_19865,N_17341,N_17892);
and U19866 (N_19866,N_17166,N_17324);
and U19867 (N_19867,N_17910,N_17385);
xnor U19868 (N_19868,N_17688,N_16259);
or U19869 (N_19869,N_17555,N_16261);
nand U19870 (N_19870,N_16677,N_16361);
or U19871 (N_19871,N_16472,N_17752);
nand U19872 (N_19872,N_17984,N_17495);
xnor U19873 (N_19873,N_16203,N_16437);
and U19874 (N_19874,N_17332,N_17284);
or U19875 (N_19875,N_17591,N_16041);
and U19876 (N_19876,N_16319,N_16919);
nor U19877 (N_19877,N_16871,N_17257);
xor U19878 (N_19878,N_17615,N_17932);
xnor U19879 (N_19879,N_16079,N_17509);
nand U19880 (N_19880,N_16460,N_17585);
nand U19881 (N_19881,N_16385,N_17325);
and U19882 (N_19882,N_17064,N_17886);
xor U19883 (N_19883,N_16528,N_16014);
xor U19884 (N_19884,N_16180,N_17607);
or U19885 (N_19885,N_16266,N_17522);
or U19886 (N_19886,N_17897,N_16014);
or U19887 (N_19887,N_16827,N_16630);
nand U19888 (N_19888,N_16956,N_17377);
or U19889 (N_19889,N_17174,N_16184);
and U19890 (N_19890,N_17326,N_17068);
nand U19891 (N_19891,N_16821,N_17619);
nor U19892 (N_19892,N_17608,N_16627);
xor U19893 (N_19893,N_16003,N_17019);
xnor U19894 (N_19894,N_17672,N_17880);
nor U19895 (N_19895,N_16863,N_16918);
nor U19896 (N_19896,N_17083,N_17764);
xnor U19897 (N_19897,N_16353,N_17657);
nor U19898 (N_19898,N_17235,N_16546);
xor U19899 (N_19899,N_16813,N_16629);
nand U19900 (N_19900,N_16817,N_17082);
or U19901 (N_19901,N_16667,N_17968);
xor U19902 (N_19902,N_16571,N_17489);
and U19903 (N_19903,N_17866,N_17479);
and U19904 (N_19904,N_17106,N_17566);
and U19905 (N_19905,N_16262,N_16038);
xor U19906 (N_19906,N_16509,N_17933);
nand U19907 (N_19907,N_17837,N_17345);
nor U19908 (N_19908,N_16361,N_17792);
and U19909 (N_19909,N_16363,N_16511);
nand U19910 (N_19910,N_17532,N_17760);
and U19911 (N_19911,N_16758,N_16767);
and U19912 (N_19912,N_16236,N_16395);
nand U19913 (N_19913,N_17347,N_17842);
or U19914 (N_19914,N_17133,N_17585);
and U19915 (N_19915,N_17033,N_16700);
nand U19916 (N_19916,N_16119,N_16621);
and U19917 (N_19917,N_16497,N_17582);
or U19918 (N_19918,N_16664,N_17560);
nor U19919 (N_19919,N_16368,N_16307);
and U19920 (N_19920,N_17327,N_16610);
or U19921 (N_19921,N_17300,N_17506);
nor U19922 (N_19922,N_16997,N_16873);
and U19923 (N_19923,N_17001,N_17146);
or U19924 (N_19924,N_17665,N_17034);
or U19925 (N_19925,N_16953,N_16002);
and U19926 (N_19926,N_17997,N_17022);
or U19927 (N_19927,N_17841,N_17091);
xor U19928 (N_19928,N_16283,N_16094);
and U19929 (N_19929,N_16734,N_17111);
nor U19930 (N_19930,N_17747,N_16079);
nor U19931 (N_19931,N_16036,N_16446);
and U19932 (N_19932,N_16325,N_16525);
nand U19933 (N_19933,N_16940,N_16103);
xor U19934 (N_19934,N_16433,N_16761);
nor U19935 (N_19935,N_17521,N_16427);
or U19936 (N_19936,N_17503,N_16315);
xnor U19937 (N_19937,N_16649,N_17446);
and U19938 (N_19938,N_17410,N_17237);
nor U19939 (N_19939,N_16914,N_17452);
and U19940 (N_19940,N_16457,N_16614);
xor U19941 (N_19941,N_16884,N_17288);
and U19942 (N_19942,N_16124,N_16775);
and U19943 (N_19943,N_17829,N_16582);
or U19944 (N_19944,N_16473,N_16285);
nor U19945 (N_19945,N_16274,N_17434);
nor U19946 (N_19946,N_17542,N_16876);
nor U19947 (N_19947,N_16963,N_17430);
or U19948 (N_19948,N_17587,N_17001);
nor U19949 (N_19949,N_17308,N_16368);
xnor U19950 (N_19950,N_17210,N_17135);
nand U19951 (N_19951,N_16582,N_16502);
or U19952 (N_19952,N_16935,N_16598);
nor U19953 (N_19953,N_17858,N_17401);
nor U19954 (N_19954,N_16371,N_17964);
xor U19955 (N_19955,N_17362,N_16981);
xor U19956 (N_19956,N_16388,N_16409);
and U19957 (N_19957,N_17498,N_17215);
or U19958 (N_19958,N_17698,N_17595);
nand U19959 (N_19959,N_17501,N_16225);
nand U19960 (N_19960,N_17129,N_17509);
or U19961 (N_19961,N_16422,N_17927);
nor U19962 (N_19962,N_16955,N_17818);
nand U19963 (N_19963,N_16672,N_17524);
nand U19964 (N_19964,N_17153,N_16645);
nand U19965 (N_19965,N_16240,N_17474);
xnor U19966 (N_19966,N_16388,N_17370);
or U19967 (N_19967,N_17975,N_17168);
xor U19968 (N_19968,N_16519,N_16136);
nand U19969 (N_19969,N_16733,N_17228);
nand U19970 (N_19970,N_17092,N_16770);
and U19971 (N_19971,N_17187,N_16333);
nand U19972 (N_19972,N_17472,N_16044);
xor U19973 (N_19973,N_16485,N_17873);
or U19974 (N_19974,N_17832,N_16220);
and U19975 (N_19975,N_16360,N_16259);
nor U19976 (N_19976,N_17203,N_17492);
nand U19977 (N_19977,N_17631,N_17954);
and U19978 (N_19978,N_16691,N_17811);
xnor U19979 (N_19979,N_17245,N_17750);
nand U19980 (N_19980,N_16716,N_17067);
nor U19981 (N_19981,N_16900,N_16293);
nor U19982 (N_19982,N_17569,N_16729);
xor U19983 (N_19983,N_17727,N_17385);
and U19984 (N_19984,N_17257,N_16625);
nand U19985 (N_19985,N_17184,N_16382);
xor U19986 (N_19986,N_17795,N_16601);
xor U19987 (N_19987,N_17965,N_16342);
and U19988 (N_19988,N_16789,N_17654);
nor U19989 (N_19989,N_16339,N_16874);
xnor U19990 (N_19990,N_17491,N_17230);
nand U19991 (N_19991,N_16259,N_16108);
and U19992 (N_19992,N_16855,N_16975);
and U19993 (N_19993,N_17973,N_16791);
or U19994 (N_19994,N_16034,N_16519);
nand U19995 (N_19995,N_17010,N_16464);
nand U19996 (N_19996,N_16009,N_17145);
and U19997 (N_19997,N_16568,N_16768);
nor U19998 (N_19998,N_16674,N_17389);
or U19999 (N_19999,N_16808,N_16031);
or UO_0 (O_0,N_19877,N_18769);
nand UO_1 (O_1,N_19186,N_18926);
nor UO_2 (O_2,N_18617,N_18412);
nor UO_3 (O_3,N_18106,N_19347);
nor UO_4 (O_4,N_18380,N_18679);
xnor UO_5 (O_5,N_19904,N_19955);
nand UO_6 (O_6,N_19643,N_18952);
nor UO_7 (O_7,N_19695,N_18929);
or UO_8 (O_8,N_18967,N_18627);
nand UO_9 (O_9,N_18141,N_18041);
nand UO_10 (O_10,N_19379,N_18973);
and UO_11 (O_11,N_18860,N_19563);
nand UO_12 (O_12,N_18554,N_18757);
xnor UO_13 (O_13,N_19680,N_19638);
nor UO_14 (O_14,N_18726,N_19461);
and UO_15 (O_15,N_19051,N_19453);
xnor UO_16 (O_16,N_18390,N_19690);
xnor UO_17 (O_17,N_19896,N_18869);
or UO_18 (O_18,N_19891,N_18817);
xnor UO_19 (O_19,N_19516,N_18748);
and UO_20 (O_20,N_19893,N_18675);
or UO_21 (O_21,N_18121,N_19603);
xnor UO_22 (O_22,N_18942,N_19102);
and UO_23 (O_23,N_19411,N_18013);
and UO_24 (O_24,N_18725,N_18824);
nand UO_25 (O_25,N_18110,N_19369);
nand UO_26 (O_26,N_19730,N_18169);
xor UO_27 (O_27,N_19240,N_19823);
nor UO_28 (O_28,N_18666,N_18338);
and UO_29 (O_29,N_19149,N_19203);
and UO_30 (O_30,N_19530,N_19789);
xnor UO_31 (O_31,N_19807,N_18045);
nor UO_32 (O_32,N_18095,N_18242);
and UO_33 (O_33,N_19123,N_19555);
nand UO_34 (O_34,N_18904,N_18198);
and UO_35 (O_35,N_19572,N_18466);
and UO_36 (O_36,N_18670,N_18381);
or UO_37 (O_37,N_19947,N_19064);
and UO_38 (O_38,N_19329,N_18373);
nand UO_39 (O_39,N_19501,N_19734);
xor UO_40 (O_40,N_18645,N_18934);
xnor UO_41 (O_41,N_19182,N_19754);
nor UO_42 (O_42,N_18255,N_19377);
or UO_43 (O_43,N_18598,N_19951);
xor UO_44 (O_44,N_19491,N_18426);
or UO_45 (O_45,N_19076,N_18614);
or UO_46 (O_46,N_19707,N_19444);
and UO_47 (O_47,N_19245,N_19856);
nor UO_48 (O_48,N_18637,N_19156);
and UO_49 (O_49,N_19243,N_19884);
nor UO_50 (O_50,N_18009,N_18528);
and UO_51 (O_51,N_19021,N_18231);
and UO_52 (O_52,N_18264,N_19879);
or UO_53 (O_53,N_18406,N_18222);
nor UO_54 (O_54,N_19757,N_19894);
xnor UO_55 (O_55,N_18657,N_19079);
and UO_56 (O_56,N_19790,N_18691);
or UO_57 (O_57,N_18520,N_19756);
and UO_58 (O_58,N_19388,N_19748);
and UO_59 (O_59,N_18132,N_19799);
and UO_60 (O_60,N_18833,N_18310);
nand UO_61 (O_61,N_18035,N_18127);
nor UO_62 (O_62,N_18079,N_19348);
xor UO_63 (O_63,N_19435,N_19525);
or UO_64 (O_64,N_18167,N_18667);
and UO_65 (O_65,N_18366,N_19284);
xnor UO_66 (O_66,N_19066,N_18839);
and UO_67 (O_67,N_18492,N_19866);
nand UO_68 (O_68,N_19164,N_18287);
nand UO_69 (O_69,N_18540,N_18100);
xor UO_70 (O_70,N_18285,N_19306);
nor UO_71 (O_71,N_19508,N_19242);
xor UO_72 (O_72,N_18468,N_18341);
or UO_73 (O_73,N_18205,N_19709);
nand UO_74 (O_74,N_18410,N_19503);
nor UO_75 (O_75,N_18513,N_19036);
and UO_76 (O_76,N_19294,N_19957);
and UO_77 (O_77,N_18344,N_19241);
or UO_78 (O_78,N_18368,N_18823);
nand UO_79 (O_79,N_18245,N_19477);
and UO_80 (O_80,N_18162,N_19305);
nor UO_81 (O_81,N_19252,N_19861);
nor UO_82 (O_82,N_18574,N_19030);
xor UO_83 (O_83,N_19755,N_18714);
nor UO_84 (O_84,N_18759,N_19520);
and UO_85 (O_85,N_18053,N_18621);
nand UO_86 (O_86,N_19249,N_19539);
and UO_87 (O_87,N_19522,N_19095);
nand UO_88 (O_88,N_18490,N_19333);
and UO_89 (O_89,N_18123,N_18436);
xor UO_90 (O_90,N_19615,N_19026);
or UO_91 (O_91,N_18370,N_18154);
nor UO_92 (O_92,N_19677,N_19371);
or UO_93 (O_93,N_19853,N_19213);
and UO_94 (O_94,N_19703,N_18421);
nand UO_95 (O_95,N_18752,N_19644);
xnor UO_96 (O_96,N_18267,N_19865);
nor UO_97 (O_97,N_19074,N_18212);
nand UO_98 (O_98,N_19806,N_18047);
and UO_99 (O_99,N_19413,N_18797);
xnor UO_100 (O_100,N_19056,N_18186);
nand UO_101 (O_101,N_19147,N_19763);
nand UO_102 (O_102,N_19826,N_19636);
and UO_103 (O_103,N_19353,N_19082);
nor UO_104 (O_104,N_18082,N_19380);
nor UO_105 (O_105,N_19460,N_18136);
nor UO_106 (O_106,N_18303,N_19960);
nand UO_107 (O_107,N_19218,N_18073);
or UO_108 (O_108,N_18887,N_19208);
xor UO_109 (O_109,N_19798,N_19446);
or UO_110 (O_110,N_19005,N_18234);
nor UO_111 (O_111,N_18580,N_18304);
and UO_112 (O_112,N_18453,N_18750);
nor UO_113 (O_113,N_18743,N_19131);
nor UO_114 (O_114,N_18152,N_19109);
nor UO_115 (O_115,N_18126,N_18781);
xnor UO_116 (O_116,N_19899,N_19895);
and UO_117 (O_117,N_19682,N_19510);
nor UO_118 (O_118,N_19339,N_18225);
nand UO_119 (O_119,N_18005,N_19216);
xnor UO_120 (O_120,N_18051,N_18049);
and UO_121 (O_121,N_18316,N_19758);
or UO_122 (O_122,N_18098,N_19611);
or UO_123 (O_123,N_18995,N_18867);
and UO_124 (O_124,N_19828,N_19264);
nor UO_125 (O_125,N_18026,N_19604);
xnor UO_126 (O_126,N_19011,N_18764);
or UO_127 (O_127,N_18710,N_18064);
and UO_128 (O_128,N_18334,N_19934);
or UO_129 (O_129,N_19569,N_18912);
xor UO_130 (O_130,N_18852,N_19499);
or UO_131 (O_131,N_19013,N_18501);
or UO_132 (O_132,N_19831,N_19846);
and UO_133 (O_133,N_18564,N_18572);
nand UO_134 (O_134,N_19159,N_18427);
nand UO_135 (O_135,N_19788,N_18915);
nor UO_136 (O_136,N_19640,N_19336);
xor UO_137 (O_137,N_19923,N_19577);
xnor UO_138 (O_138,N_19321,N_19436);
nor UO_139 (O_139,N_19832,N_18806);
nor UO_140 (O_140,N_18720,N_18447);
or UO_141 (O_141,N_18607,N_18963);
and UO_142 (O_142,N_19098,N_18060);
xor UO_143 (O_143,N_19169,N_18038);
xor UO_144 (O_144,N_19833,N_18204);
nor UO_145 (O_145,N_19309,N_19500);
and UO_146 (O_146,N_19743,N_18146);
and UO_147 (O_147,N_19338,N_19268);
and UO_148 (O_148,N_19769,N_19399);
nor UO_149 (O_149,N_19044,N_19260);
or UO_150 (O_150,N_19590,N_19685);
nand UO_151 (O_151,N_19829,N_19087);
nand UO_152 (O_152,N_19981,N_18069);
and UO_153 (O_153,N_18756,N_19070);
and UO_154 (O_154,N_19854,N_18924);
nor UO_155 (O_155,N_19671,N_18903);
or UO_156 (O_156,N_18991,N_18317);
or UO_157 (O_157,N_18307,N_19850);
nand UO_158 (O_158,N_19583,N_18914);
nor UO_159 (O_159,N_19836,N_18494);
and UO_160 (O_160,N_18919,N_18092);
nand UO_161 (O_161,N_18512,N_19714);
or UO_162 (O_162,N_19608,N_18842);
nand UO_163 (O_163,N_19152,N_18104);
or UO_164 (O_164,N_18550,N_18293);
and UO_165 (O_165,N_19907,N_19495);
and UO_166 (O_166,N_18033,N_18858);
xnor UO_167 (O_167,N_19528,N_19858);
xnor UO_168 (O_168,N_19198,N_19713);
nand UO_169 (O_169,N_19429,N_18101);
xnor UO_170 (O_170,N_18199,N_18040);
and UO_171 (O_171,N_19716,N_18227);
and UO_172 (O_172,N_19418,N_19537);
nor UO_173 (O_173,N_18190,N_19927);
and UO_174 (O_174,N_19281,N_19591);
xnor UO_175 (O_175,N_18588,N_18031);
nor UO_176 (O_176,N_19916,N_18548);
nand UO_177 (O_177,N_19073,N_18791);
nand UO_178 (O_178,N_19937,N_18108);
and UO_179 (O_179,N_18827,N_18160);
xnor UO_180 (O_180,N_18702,N_19581);
and UO_181 (O_181,N_19445,N_18346);
and UO_182 (O_182,N_18599,N_18724);
nor UO_183 (O_183,N_19738,N_18601);
or UO_184 (O_184,N_18118,N_18522);
xor UO_185 (O_185,N_19296,N_19540);
or UO_186 (O_186,N_18589,N_19272);
or UO_187 (O_187,N_18099,N_18918);
nand UO_188 (O_188,N_18841,N_19745);
nand UO_189 (O_189,N_18811,N_18763);
nor UO_190 (O_190,N_18354,N_18506);
nand UO_191 (O_191,N_19433,N_19363);
nor UO_192 (O_192,N_18323,N_18059);
nor UO_193 (O_193,N_18571,N_18252);
and UO_194 (O_194,N_18185,N_18423);
xnor UO_195 (O_195,N_19120,N_19416);
nand UO_196 (O_196,N_18612,N_18340);
or UO_197 (O_197,N_18719,N_19787);
nor UO_198 (O_198,N_19982,N_19857);
nor UO_199 (O_199,N_19533,N_18418);
nor UO_200 (O_200,N_18297,N_19674);
nor UO_201 (O_201,N_18074,N_18042);
xor UO_202 (O_202,N_18362,N_19061);
xnor UO_203 (O_203,N_18523,N_19995);
nand UO_204 (O_204,N_19548,N_18678);
nor UO_205 (O_205,N_19809,N_19261);
or UO_206 (O_206,N_19843,N_19304);
xnor UO_207 (O_207,N_18565,N_18774);
xor UO_208 (O_208,N_19053,N_18885);
and UO_209 (O_209,N_19293,N_19941);
nor UO_210 (O_210,N_19514,N_18592);
xnor UO_211 (O_211,N_19223,N_18969);
xnor UO_212 (O_212,N_19570,N_19897);
or UO_213 (O_213,N_18907,N_18218);
nor UO_214 (O_214,N_19952,N_18651);
xor UO_215 (O_215,N_19080,N_19323);
nor UO_216 (O_216,N_18168,N_19055);
or UO_217 (O_217,N_18940,N_18706);
or UO_218 (O_218,N_19817,N_19386);
xnor UO_219 (O_219,N_19341,N_18276);
and UO_220 (O_220,N_18145,N_18158);
or UO_221 (O_221,N_19732,N_18676);
nor UO_222 (O_222,N_18257,N_18873);
and UO_223 (O_223,N_18740,N_18476);
or UO_224 (O_224,N_19085,N_19298);
nand UO_225 (O_225,N_19964,N_19473);
or UO_226 (O_226,N_19483,N_18911);
or UO_227 (O_227,N_18897,N_19116);
or UO_228 (O_228,N_18137,N_19419);
xor UO_229 (O_229,N_19326,N_19234);
xnor UO_230 (O_230,N_19915,N_18531);
nand UO_231 (O_231,N_18057,N_19667);
nand UO_232 (O_232,N_18001,N_19906);
or UO_233 (O_233,N_18209,N_19599);
and UO_234 (O_234,N_19471,N_18682);
and UO_235 (O_235,N_18483,N_18745);
or UO_236 (O_236,N_18125,N_19468);
xnor UO_237 (O_237,N_18845,N_18067);
or UO_238 (O_238,N_18796,N_18700);
nor UO_239 (O_239,N_18730,N_19779);
nand UO_240 (O_240,N_18133,N_19124);
nor UO_241 (O_241,N_18196,N_19687);
nor UO_242 (O_242,N_19630,N_18619);
or UO_243 (O_243,N_19840,N_19430);
nor UO_244 (O_244,N_18142,N_18420);
or UO_245 (O_245,N_18262,N_18244);
or UO_246 (O_246,N_19892,N_19513);
and UO_247 (O_247,N_18871,N_18088);
nand UO_248 (O_248,N_19967,N_19770);
xnor UO_249 (O_249,N_18349,N_19282);
xor UO_250 (O_250,N_19875,N_19199);
and UO_251 (O_251,N_19316,N_19228);
nand UO_252 (O_252,N_19361,N_19616);
or UO_253 (O_253,N_18343,N_19637);
or UO_254 (O_254,N_19178,N_18644);
or UO_255 (O_255,N_18039,N_19233);
nor UO_256 (O_256,N_18853,N_19696);
xor UO_257 (O_257,N_18219,N_19773);
or UO_258 (O_258,N_18615,N_18439);
or UO_259 (O_259,N_18080,N_19031);
xor UO_260 (O_260,N_19727,N_19586);
nor UO_261 (O_261,N_18913,N_19362);
nand UO_262 (O_262,N_19251,N_18772);
or UO_263 (O_263,N_18486,N_19506);
xor UO_264 (O_264,N_18718,N_18417);
and UO_265 (O_265,N_18898,N_19992);
and UO_266 (O_266,N_19197,N_19417);
nand UO_267 (O_267,N_18703,N_19489);
xor UO_268 (O_268,N_18835,N_18202);
xor UO_269 (O_269,N_18646,N_19848);
xor UO_270 (O_270,N_18128,N_18351);
and UO_271 (O_271,N_18360,N_18329);
nor UO_272 (O_272,N_18773,N_19062);
and UO_273 (O_273,N_19717,N_19277);
xor UO_274 (O_274,N_18046,N_19270);
and UO_275 (O_275,N_18987,N_18116);
nand UO_276 (O_276,N_19104,N_19626);
or UO_277 (O_277,N_18586,N_19175);
nand UO_278 (O_278,N_18544,N_19389);
xnor UO_279 (O_279,N_19883,N_19553);
or UO_280 (O_280,N_19645,N_18179);
and UO_281 (O_281,N_18878,N_19742);
or UO_282 (O_282,N_19800,N_19813);
and UO_283 (O_283,N_18030,N_19519);
nand UO_284 (O_284,N_18538,N_19824);
and UO_285 (O_285,N_19775,N_19354);
or UO_286 (O_286,N_18464,N_18090);
xor UO_287 (O_287,N_18533,N_18699);
and UO_288 (O_288,N_18305,N_18629);
xnor UO_289 (O_289,N_18177,N_18489);
or UO_290 (O_290,N_18477,N_19868);
or UO_291 (O_291,N_19834,N_19467);
xnor UO_292 (O_292,N_19794,N_18551);
and UO_293 (O_293,N_19037,N_18006);
nand UO_294 (O_294,N_19401,N_18197);
and UO_295 (O_295,N_19155,N_18570);
xor UO_296 (O_296,N_18378,N_19852);
xnor UO_297 (O_297,N_18470,N_19122);
nor UO_298 (O_298,N_19008,N_19457);
nor UO_299 (O_299,N_19334,N_19784);
nor UO_300 (O_300,N_18686,N_18587);
or UO_301 (O_301,N_18216,N_19912);
nor UO_302 (O_302,N_19774,N_18534);
or UO_303 (O_303,N_19239,N_19975);
nor UO_304 (O_304,N_18992,N_19057);
and UO_305 (O_305,N_19451,N_19238);
xnor UO_306 (O_306,N_18594,N_18156);
and UO_307 (O_307,N_19969,N_18084);
or UO_308 (O_308,N_19255,N_18089);
xor UO_309 (O_309,N_18290,N_18744);
xor UO_310 (O_310,N_18019,N_19518);
and UO_311 (O_311,N_19367,N_18778);
or UO_312 (O_312,N_19126,N_18313);
and UO_313 (O_313,N_19052,N_19527);
nor UO_314 (O_314,N_19613,N_19803);
and UO_315 (O_315,N_19003,N_19511);
or UO_316 (O_316,N_18171,N_19562);
or UO_317 (O_317,N_18445,N_19276);
xor UO_318 (O_318,N_18113,N_19931);
nand UO_319 (O_319,N_18386,N_19165);
xnor UO_320 (O_320,N_19872,N_19001);
xor UO_321 (O_321,N_18451,N_19837);
nor UO_322 (O_322,N_18561,N_19881);
or UO_323 (O_323,N_19322,N_18639);
and UO_324 (O_324,N_19237,N_18062);
xnor UO_325 (O_325,N_19134,N_19780);
xor UO_326 (O_326,N_19426,N_18736);
or UO_327 (O_327,N_18640,N_18318);
xor UO_328 (O_328,N_18888,N_18484);
nand UO_329 (O_329,N_18359,N_18389);
and UO_330 (O_330,N_19614,N_19302);
and UO_331 (O_331,N_18668,N_19766);
nor UO_332 (O_332,N_18892,N_19971);
xor UO_333 (O_333,N_18664,N_19753);
or UO_334 (O_334,N_18462,N_19097);
and UO_335 (O_335,N_19619,N_19622);
nor UO_336 (O_336,N_19248,N_19166);
or UO_337 (O_337,N_18365,N_19634);
or UO_338 (O_338,N_18737,N_19431);
nand UO_339 (O_339,N_19108,N_19595);
nand UO_340 (O_340,N_19855,N_18779);
and UO_341 (O_341,N_18192,N_19689);
nand UO_342 (O_342,N_19917,N_18505);
nand UO_343 (O_343,N_19768,N_19113);
nor UO_344 (O_344,N_19439,N_18847);
and UO_345 (O_345,N_19765,N_19232);
or UO_346 (O_346,N_19258,N_18107);
nor UO_347 (O_347,N_19356,N_19534);
or UO_348 (O_348,N_19115,N_19507);
nor UO_349 (O_349,N_18810,N_19878);
or UO_350 (O_350,N_19089,N_19236);
and UO_351 (O_351,N_18511,N_18294);
xor UO_352 (O_352,N_19521,N_18821);
or UO_353 (O_353,N_18465,N_18274);
nand UO_354 (O_354,N_19532,N_19024);
or UO_355 (O_355,N_18993,N_18825);
nand UO_356 (O_356,N_19358,N_18717);
xnor UO_357 (O_357,N_18696,N_19459);
xor UO_358 (O_358,N_19929,N_19818);
and UO_359 (O_359,N_19141,N_19978);
nor UO_360 (O_360,N_18923,N_19202);
and UO_361 (O_361,N_18944,N_19132);
and UO_362 (O_362,N_19462,N_18659);
and UO_363 (O_363,N_19215,N_19889);
or UO_364 (O_364,N_19139,N_19541);
xnor UO_365 (O_365,N_19176,N_19396);
nand UO_366 (O_366,N_18739,N_18948);
xnor UO_367 (O_367,N_18596,N_18058);
nor UO_368 (O_368,N_18224,N_18861);
xnor UO_369 (O_369,N_18709,N_18174);
nor UO_370 (O_370,N_19966,N_19607);
xnor UO_371 (O_371,N_18093,N_19188);
xnor UO_372 (O_372,N_19009,N_19876);
or UO_373 (O_373,N_19761,N_18097);
nor UO_374 (O_374,N_19403,N_19454);
and UO_375 (O_375,N_18901,N_19578);
nand UO_376 (O_376,N_18278,N_18474);
nand UO_377 (O_377,N_19317,N_18721);
nor UO_378 (O_378,N_18481,N_18655);
and UO_379 (O_379,N_19220,N_19962);
nand UO_380 (O_380,N_18665,N_18363);
and UO_381 (O_381,N_18358,N_19722);
nand UO_382 (O_382,N_19177,N_19554);
and UO_383 (O_383,N_18980,N_18306);
nor UO_384 (O_384,N_18652,N_18413);
nand UO_385 (O_385,N_18864,N_19183);
or UO_386 (O_386,N_19121,N_18976);
nor UO_387 (O_387,N_19623,N_19873);
nor UO_388 (O_388,N_18529,N_19455);
or UO_389 (O_389,N_19744,N_18176);
nor UO_390 (O_390,N_19557,N_18183);
nand UO_391 (O_391,N_19808,N_18630);
and UO_392 (O_392,N_19926,N_19256);
or UO_393 (O_393,N_19664,N_18254);
nor UO_394 (O_394,N_18749,N_19487);
nor UO_395 (O_395,N_19844,N_19448);
nand UO_396 (O_396,N_18933,N_19484);
nor UO_397 (O_397,N_18124,N_19589);
or UO_398 (O_398,N_19880,N_19476);
xor UO_399 (O_399,N_18960,N_18383);
and UO_400 (O_400,N_18454,N_18552);
xor UO_401 (O_401,N_18705,N_18459);
and UO_402 (O_402,N_18555,N_18238);
and UO_403 (O_403,N_19890,N_18279);
and UO_404 (O_404,N_18938,N_18734);
xor UO_405 (O_405,N_18003,N_18525);
nor UO_406 (O_406,N_18836,N_19665);
and UO_407 (O_407,N_19512,N_19691);
nor UO_408 (O_408,N_18765,N_18435);
xnor UO_409 (O_409,N_18844,N_19368);
and UO_410 (O_410,N_19253,N_18025);
nor UO_411 (O_411,N_18953,N_18526);
or UO_412 (O_412,N_18256,N_18775);
nor UO_413 (O_413,N_18229,N_19472);
or UO_414 (O_414,N_19804,N_18939);
xor UO_415 (O_415,N_19342,N_19535);
and UO_416 (O_416,N_18191,N_19908);
xnor UO_417 (O_417,N_19792,N_19588);
xor UO_418 (O_418,N_18648,N_18102);
xnor UO_419 (O_419,N_18021,N_18786);
and UO_420 (O_420,N_18813,N_19020);
xor UO_421 (O_421,N_18475,N_18391);
xor UO_422 (O_422,N_18377,N_19905);
nor UO_423 (O_423,N_18339,N_19729);
xor UO_424 (O_424,N_19559,N_18315);
and UO_425 (O_425,N_18086,N_19273);
or UO_426 (O_426,N_19310,N_18002);
nor UO_427 (O_427,N_19606,N_19762);
and UO_428 (O_428,N_19355,N_18761);
xor UO_429 (O_429,N_19432,N_19303);
and UO_430 (O_430,N_19230,N_18450);
xnor UO_431 (O_431,N_18994,N_18295);
nor UO_432 (O_432,N_19320,N_19920);
and UO_433 (O_433,N_18798,N_19415);
nand UO_434 (O_434,N_18249,N_18044);
nor UO_435 (O_435,N_19701,N_18809);
or UO_436 (O_436,N_19274,N_19949);
and UO_437 (O_437,N_18947,N_18760);
nor UO_438 (O_438,N_19479,N_18240);
xnor UO_439 (O_439,N_19968,N_18965);
nand UO_440 (O_440,N_18579,N_18954);
or UO_441 (O_441,N_19579,N_18232);
and UO_442 (O_442,N_18850,N_19058);
xnor UO_443 (O_443,N_18680,N_19071);
xor UO_444 (O_444,N_19505,N_19096);
nand UO_445 (O_445,N_19576,N_19924);
and UO_446 (O_446,N_18502,N_18336);
and UO_447 (O_447,N_18814,N_18028);
nor UO_448 (O_448,N_19724,N_18016);
nor UO_449 (O_449,N_19028,N_19404);
nand UO_450 (O_450,N_18054,N_19536);
nand UO_451 (O_451,N_18201,N_19933);
nor UO_452 (O_452,N_19378,N_18497);
or UO_453 (O_453,N_19287,N_18122);
xor UO_454 (O_454,N_18496,N_18189);
and UO_455 (O_455,N_19084,N_18071);
xor UO_456 (O_456,N_18065,N_19428);
or UO_457 (O_457,N_19391,N_18524);
and UO_458 (O_458,N_18573,N_18181);
nand UO_459 (O_459,N_18425,N_18217);
xnor UO_460 (O_460,N_18353,N_19214);
xnor UO_461 (O_461,N_19315,N_18870);
or UO_462 (O_462,N_18762,N_18747);
or UO_463 (O_463,N_18155,N_18382);
xnor UO_464 (O_464,N_18899,N_19075);
nor UO_465 (O_465,N_18673,N_18348);
xor UO_466 (O_466,N_19746,N_19170);
and UO_467 (O_467,N_18138,N_19523);
nand UO_468 (O_468,N_18401,N_18677);
nor UO_469 (O_469,N_18273,N_18165);
or UO_470 (O_470,N_19493,N_18480);
and UO_471 (O_471,N_19652,N_18446);
and UO_472 (O_472,N_19192,N_19434);
or UO_473 (O_473,N_19065,N_18076);
and UO_474 (O_474,N_18784,N_18787);
nor UO_475 (O_475,N_18325,N_18419);
xnor UO_476 (O_476,N_19299,N_18590);
and UO_477 (O_477,N_19819,N_18857);
nand UO_478 (O_478,N_19802,N_19767);
nor UO_479 (O_479,N_19375,N_18893);
nor UO_480 (O_480,N_18180,N_19751);
and UO_481 (O_481,N_18024,N_19681);
and UO_482 (O_482,N_18433,N_18547);
xor UO_483 (O_483,N_18795,N_19440);
and UO_484 (O_484,N_18854,N_19475);
xnor UO_485 (O_485,N_18392,N_19721);
nand UO_486 (O_486,N_19150,N_18442);
nor UO_487 (O_487,N_18029,N_19810);
and UO_488 (O_488,N_18335,N_18471);
xnor UO_489 (O_489,N_18558,N_18129);
nand UO_490 (O_490,N_19048,N_19946);
and UO_491 (O_491,N_18925,N_19550);
or UO_492 (O_492,N_18658,N_18488);
or UO_493 (O_493,N_18269,N_19189);
nor UO_494 (O_494,N_19014,N_18105);
xor UO_495 (O_495,N_19584,N_19033);
nor UO_496 (O_496,N_19795,N_18443);
or UO_497 (O_497,N_19250,N_18770);
nand UO_498 (O_498,N_19482,N_19335);
nor UO_499 (O_499,N_19827,N_18131);
nand UO_500 (O_500,N_19700,N_19262);
nand UO_501 (O_501,N_18921,N_19777);
and UO_502 (O_502,N_19602,N_18299);
nor UO_503 (O_503,N_18050,N_19863);
and UO_504 (O_504,N_19191,N_18920);
and UO_505 (O_505,N_18837,N_19269);
or UO_506 (O_506,N_19620,N_18188);
xor UO_507 (O_507,N_19699,N_18135);
and UO_508 (O_508,N_19373,N_18711);
nand UO_509 (O_509,N_19225,N_19088);
nor UO_510 (O_510,N_19295,N_19494);
xnor UO_511 (O_511,N_18260,N_19247);
nor UO_512 (O_512,N_19723,N_18210);
nand UO_513 (O_513,N_18751,N_19542);
nand UO_514 (O_514,N_19161,N_19345);
nand UO_515 (O_515,N_18220,N_18626);
xnor UO_516 (O_516,N_18566,N_19114);
and UO_517 (O_517,N_18239,N_18010);
xnor UO_518 (O_518,N_18620,N_19601);
nor UO_519 (O_519,N_18000,N_19936);
nand UO_520 (O_520,N_19911,N_19480);
nor UO_521 (O_521,N_18157,N_19672);
or UO_522 (O_522,N_18081,N_19785);
or UO_523 (O_523,N_19776,N_18330);
nand UO_524 (O_524,N_18251,N_19580);
nor UO_525 (O_525,N_18332,N_18958);
nor UO_526 (O_526,N_18072,N_19181);
nor UO_527 (O_527,N_18103,N_18656);
nor UO_528 (O_528,N_19662,N_18321);
nand UO_529 (O_529,N_19888,N_19330);
nor UO_530 (O_530,N_18403,N_18868);
and UO_531 (O_531,N_18519,N_19659);
nand UO_532 (O_532,N_19488,N_18402);
xnor UO_533 (O_533,N_18514,N_18746);
xnor UO_534 (O_534,N_19726,N_18077);
or UO_535 (O_535,N_19259,N_19886);
nor UO_536 (O_536,N_19953,N_18491);
nand UO_537 (O_537,N_19515,N_18014);
nand UO_538 (O_538,N_19688,N_19706);
nand UO_539 (O_539,N_19582,N_19366);
nor UO_540 (O_540,N_19212,N_19190);
xnor UO_541 (O_541,N_18593,N_19921);
and UO_542 (O_542,N_19509,N_18731);
nor UO_543 (O_543,N_18441,N_18504);
and UO_544 (O_544,N_19466,N_19497);
nand UO_545 (O_545,N_19424,N_18187);
or UO_546 (O_546,N_18802,N_18361);
or UO_547 (O_547,N_19381,N_18962);
nor UO_548 (O_548,N_19728,N_18374);
or UO_549 (O_549,N_19291,N_18984);
nand UO_550 (O_550,N_18968,N_18527);
xnor UO_551 (O_551,N_19452,N_19091);
nor UO_552 (O_552,N_18034,N_19991);
or UO_553 (O_553,N_19441,N_19712);
nand UO_554 (O_554,N_18576,N_18729);
and UO_555 (O_555,N_18326,N_19693);
and UO_556 (O_556,N_18581,N_18961);
or UO_557 (O_557,N_18559,N_19319);
or UO_558 (O_558,N_18568,N_18008);
and UO_559 (O_559,N_18616,N_18553);
xor UO_560 (O_560,N_19385,N_18879);
xor UO_561 (O_561,N_18261,N_18367);
nor UO_562 (O_562,N_18270,N_18910);
or UO_563 (O_563,N_19231,N_19168);
nand UO_564 (O_564,N_18203,N_19206);
nand UO_565 (O_565,N_18078,N_18007);
or UO_566 (O_566,N_18661,N_19594);
and UO_567 (O_567,N_19200,N_18440);
nand UO_568 (O_568,N_18755,N_19110);
nor UO_569 (O_569,N_18182,N_19384);
xnor UO_570 (O_570,N_18866,N_19449);
xor UO_571 (O_571,N_19913,N_18148);
or UO_572 (O_572,N_19597,N_18395);
or UO_573 (O_573,N_18820,N_19312);
nand UO_574 (O_574,N_19300,N_19195);
xnor UO_575 (O_575,N_19112,N_18634);
nand UO_576 (O_576,N_19592,N_18716);
or UO_577 (O_577,N_18543,N_19167);
or UO_578 (O_578,N_18472,N_19816);
nor UO_579 (O_579,N_19633,N_19474);
or UO_580 (O_580,N_19450,N_19129);
nor UO_581 (O_581,N_18022,N_19370);
nor UO_582 (O_582,N_19422,N_18130);
nand UO_583 (O_583,N_18253,N_18606);
xnor UO_584 (O_584,N_19812,N_19574);
and UO_585 (O_585,N_18517,N_18562);
or UO_586 (O_586,N_18094,N_18681);
xnor UO_587 (O_587,N_18012,N_19543);
or UO_588 (O_588,N_19327,N_19990);
nor UO_589 (O_589,N_19311,N_18688);
and UO_590 (O_590,N_19022,N_19568);
nor UO_591 (O_591,N_19196,N_18376);
nor UO_592 (O_592,N_18371,N_19351);
or UO_593 (O_593,N_19984,N_19617);
nand UO_594 (O_594,N_19292,N_18604);
nor UO_595 (O_595,N_19328,N_19337);
xnor UO_596 (O_596,N_18309,N_18863);
nand UO_597 (O_597,N_19420,N_19958);
xor UO_598 (O_598,N_18998,N_18056);
and UO_599 (O_599,N_19596,N_18438);
nor UO_600 (O_600,N_18916,N_19651);
nor UO_601 (O_601,N_18048,N_19103);
or UO_602 (O_602,N_19650,N_19267);
and UO_603 (O_603,N_19545,N_19194);
nor UO_604 (O_604,N_19697,N_18302);
xnor UO_605 (O_605,N_19882,N_18263);
and UO_606 (O_606,N_18884,N_19997);
nand UO_607 (O_607,N_18908,N_19010);
and UO_608 (O_608,N_18430,N_18859);
or UO_609 (O_609,N_19106,N_19346);
xor UO_610 (O_610,N_19408,N_19027);
or UO_611 (O_611,N_19077,N_18622);
and UO_612 (O_612,N_19711,N_19012);
nor UO_613 (O_613,N_18741,N_19571);
nor UO_614 (O_614,N_18387,N_19821);
xnor UO_615 (O_615,N_19344,N_18609);
xnor UO_616 (O_616,N_18613,N_19365);
xor UO_617 (O_617,N_18713,N_19526);
xor UO_618 (O_618,N_18521,N_18723);
or UO_619 (O_619,N_19624,N_19111);
nand UO_620 (O_620,N_18635,N_19653);
nand UO_621 (O_621,N_19410,N_19137);
or UO_622 (O_622,N_18355,N_18922);
xor UO_623 (O_623,N_19625,N_18405);
xor UO_624 (O_624,N_19314,N_19708);
xor UO_625 (O_625,N_18292,N_18134);
nor UO_626 (O_626,N_19771,N_18460);
or UO_627 (O_627,N_19222,N_18036);
or UO_628 (O_628,N_19669,N_19948);
nand UO_629 (O_629,N_19538,N_19961);
or UO_630 (O_630,N_18027,N_19490);
xor UO_631 (O_631,N_18337,N_18535);
and UO_632 (O_632,N_18793,N_19204);
and UO_633 (O_633,N_18456,N_18780);
or UO_634 (O_634,N_19107,N_18461);
and UO_635 (O_635,N_18715,N_18055);
xnor UO_636 (O_636,N_19552,N_18610);
xnor UO_637 (O_637,N_18017,N_18999);
nand UO_638 (O_638,N_18004,N_18672);
nor UO_639 (O_639,N_19332,N_19627);
xor UO_640 (O_640,N_18935,N_19845);
and UO_641 (O_641,N_19083,N_18815);
nor UO_642 (O_642,N_18416,N_18978);
or UO_643 (O_643,N_18411,N_19072);
or UO_644 (O_644,N_18541,N_19646);
and UO_645 (O_645,N_19063,N_19340);
nor UO_646 (O_646,N_19127,N_19786);
xnor UO_647 (O_647,N_19517,N_19173);
nor UO_648 (O_648,N_18241,N_18930);
nor UO_649 (O_649,N_19945,N_18653);
nand UO_650 (O_650,N_19556,N_19822);
nand UO_651 (O_651,N_18970,N_18674);
or UO_652 (O_652,N_18979,N_18347);
and UO_653 (O_653,N_19678,N_18794);
nand UO_654 (O_654,N_18328,N_19987);
xor UO_655 (O_655,N_19119,N_19360);
xnor UO_656 (O_656,N_19443,N_19725);
xor UO_657 (O_657,N_19985,N_18818);
and UO_658 (O_658,N_19567,N_18927);
or UO_659 (O_659,N_19397,N_18518);
nand UO_660 (O_660,N_18597,N_19862);
nor UO_661 (O_661,N_18037,N_18828);
and UO_662 (O_662,N_18856,N_18298);
or UO_663 (O_663,N_18111,N_18693);
nand UO_664 (O_664,N_18955,N_19737);
nand UO_665 (O_665,N_19049,N_18971);
xor UO_666 (O_666,N_18469,N_19227);
nand UO_667 (O_667,N_19163,N_18689);
and UO_668 (O_668,N_18883,N_19673);
nand UO_669 (O_669,N_19778,N_19395);
nor UO_670 (O_670,N_19244,N_19585);
xnor UO_671 (O_671,N_18018,N_19932);
nand UO_672 (O_672,N_18964,N_19041);
xor UO_673 (O_673,N_19412,N_18647);
nor UO_674 (O_674,N_18990,N_19898);
nor UO_675 (O_675,N_19221,N_18173);
nand UO_676 (O_676,N_18660,N_18301);
nand UO_677 (O_677,N_18300,N_18800);
or UO_678 (O_678,N_18642,N_18345);
nor UO_679 (O_679,N_19485,N_19902);
and UO_680 (O_680,N_18221,N_19160);
and UO_681 (O_681,N_18785,N_18463);
or UO_682 (O_682,N_18891,N_18877);
xor UO_683 (O_683,N_19201,N_18583);
nand UO_684 (O_684,N_19394,N_19492);
nor UO_685 (O_685,N_18331,N_19343);
nor UO_686 (O_686,N_18595,N_19942);
nand UO_687 (O_687,N_19587,N_19040);
nand UO_688 (O_688,N_19157,N_19018);
nand UO_689 (O_689,N_18989,N_18208);
nor UO_690 (O_690,N_19830,N_18928);
and UO_691 (O_691,N_19078,N_18889);
and UO_692 (O_692,N_19791,N_19654);
and UO_693 (O_693,N_18886,N_18246);
nor UO_694 (O_694,N_18479,N_19764);
or UO_695 (O_695,N_19702,N_19560);
nor UO_696 (O_696,N_18832,N_19859);
and UO_697 (O_697,N_19285,N_19747);
or UO_698 (O_698,N_18457,N_18259);
nor UO_699 (O_699,N_19976,N_19983);
xnor UO_700 (O_700,N_18388,N_19612);
or UO_701 (O_701,N_18385,N_18650);
and UO_702 (O_702,N_19144,N_19938);
xnor UO_703 (O_703,N_19609,N_19679);
and UO_704 (O_704,N_19447,N_18379);
nand UO_705 (O_705,N_18662,N_18758);
and UO_706 (O_706,N_18139,N_19263);
nor UO_707 (O_707,N_19382,N_19017);
nor UO_708 (O_708,N_19839,N_18375);
and UO_709 (O_709,N_18322,N_18214);
and UO_710 (O_710,N_19463,N_19950);
or UO_711 (O_711,N_18975,N_19099);
and UO_712 (O_712,N_18372,N_18546);
nor UO_713 (O_713,N_19387,N_18628);
or UO_714 (O_714,N_18766,N_18698);
nand UO_715 (O_715,N_18140,N_18286);
nor UO_716 (O_716,N_19067,N_18654);
and UO_717 (O_717,N_18478,N_18849);
and UO_718 (O_718,N_19086,N_18830);
and UO_719 (O_719,N_18803,N_18109);
or UO_720 (O_720,N_18692,N_19162);
nor UO_721 (O_721,N_18150,N_18738);
and UO_722 (O_722,N_18996,N_18603);
xnor UO_723 (O_723,N_19741,N_19524);
and UO_724 (O_724,N_19657,N_18364);
and UO_725 (O_725,N_19814,N_18697);
xnor UO_726 (O_726,N_19979,N_19631);
nor UO_727 (O_727,N_18807,N_18194);
nand UO_728 (O_728,N_19301,N_19647);
nand UO_729 (O_729,N_18950,N_19209);
nand UO_730 (O_730,N_18536,N_18175);
or UO_731 (O_731,N_18510,N_18327);
nand UO_732 (O_732,N_18671,N_18909);
or UO_733 (O_733,N_19034,N_18195);
and UO_734 (O_734,N_18384,N_18144);
and UO_735 (O_735,N_18683,N_18143);
or UO_736 (O_736,N_19558,N_18455);
and UO_737 (O_737,N_18695,N_19675);
and UO_738 (O_738,N_18789,N_19797);
nand UO_739 (O_739,N_19136,N_18556);
and UO_740 (O_740,N_18091,N_18396);
nor UO_741 (O_741,N_19733,N_19849);
and UO_742 (O_742,N_18211,N_18846);
nor UO_743 (O_743,N_18848,N_19297);
and UO_744 (O_744,N_19719,N_18567);
and UO_745 (O_745,N_19437,N_19133);
xnor UO_746 (O_746,N_18618,N_19090);
and UO_747 (O_747,N_18808,N_18397);
or UO_748 (O_748,N_18467,N_19698);
nor UO_749 (O_749,N_19069,N_18569);
xnor UO_750 (O_750,N_19464,N_19171);
nor UO_751 (O_751,N_19735,N_18632);
nor UO_752 (O_752,N_19414,N_18499);
nand UO_753 (O_753,N_18545,N_18070);
nor UO_754 (O_754,N_18582,N_19996);
and UO_755 (O_755,N_19235,N_18166);
xnor UO_756 (O_756,N_18237,N_19145);
and UO_757 (O_757,N_18272,N_19715);
nor UO_758 (O_758,N_18083,N_18409);
nand UO_759 (O_759,N_19400,N_19390);
and UO_760 (O_760,N_19944,N_18288);
or UO_761 (O_761,N_18782,N_19265);
nand UO_762 (O_762,N_19731,N_19740);
and UO_763 (O_763,N_18872,N_19928);
nand UO_764 (O_764,N_18495,N_19023);
or UO_765 (O_765,N_19308,N_19047);
nor UO_766 (O_766,N_18284,N_18282);
xor UO_767 (O_767,N_18838,N_19350);
or UO_768 (O_768,N_19456,N_19874);
nor UO_769 (O_769,N_18394,N_18408);
nor UO_770 (O_770,N_18875,N_19019);
or UO_771 (O_771,N_18352,N_18608);
nor UO_772 (O_772,N_18694,N_18431);
xor UO_773 (O_773,N_18085,N_19910);
nor UO_774 (O_774,N_18200,N_18314);
nor UO_775 (O_775,N_19184,N_18742);
nor UO_776 (O_776,N_18114,N_19393);
nand UO_777 (O_777,N_18342,N_18207);
nand UO_778 (O_778,N_19847,N_19092);
and UO_779 (O_779,N_19704,N_18015);
xnor UO_780 (O_780,N_19988,N_19546);
nor UO_781 (O_781,N_18161,N_18448);
and UO_782 (O_782,N_18268,N_19648);
nand UO_783 (O_783,N_19649,N_19864);
nand UO_784 (O_784,N_19993,N_19998);
nor UO_785 (O_785,N_18941,N_18398);
nor UO_786 (O_786,N_18937,N_18399);
or UO_787 (O_787,N_19943,N_18902);
xor UO_788 (O_788,N_19940,N_18633);
or UO_789 (O_789,N_19364,N_18247);
nand UO_790 (O_790,N_18277,N_19635);
or UO_791 (O_791,N_19486,N_19465);
and UO_792 (O_792,N_19035,N_19504);
or UO_793 (O_793,N_18946,N_18754);
nor UO_794 (O_794,N_19146,N_19405);
nand UO_795 (O_795,N_18066,N_19666);
nor UO_796 (O_796,N_18061,N_19739);
xnor UO_797 (O_797,N_19100,N_19684);
and UO_798 (O_798,N_18170,N_18788);
nor UO_799 (O_799,N_19286,N_19925);
or UO_800 (O_800,N_19039,N_19593);
or UO_801 (O_801,N_19901,N_19438);
nand UO_802 (O_802,N_18147,N_19496);
nand UO_803 (O_803,N_18117,N_19885);
or UO_804 (O_804,N_18226,N_19143);
and UO_805 (O_805,N_19801,N_19994);
xor UO_806 (O_806,N_19922,N_18685);
nor UO_807 (O_807,N_18452,N_19187);
and UO_808 (O_808,N_19974,N_19442);
or UO_809 (O_809,N_19458,N_18153);
nand UO_810 (O_810,N_18957,N_18516);
nand UO_811 (O_811,N_19398,N_18687);
or UO_812 (O_812,N_18549,N_19796);
nand UO_813 (O_813,N_18233,N_19006);
or UO_814 (O_814,N_18605,N_19125);
and UO_815 (O_815,N_18515,N_18193);
or UO_816 (O_816,N_19406,N_19138);
or UO_817 (O_817,N_18959,N_18115);
nor UO_818 (O_818,N_19349,N_18983);
and UO_819 (O_819,N_19470,N_18905);
nand UO_820 (O_820,N_18087,N_19081);
and UO_821 (O_821,N_18767,N_19618);
nand UO_822 (O_822,N_18407,N_19004);
and UO_823 (O_823,N_19825,N_19935);
nor UO_824 (O_824,N_18585,N_18974);
nand UO_825 (O_825,N_18643,N_18816);
nor UO_826 (O_826,N_19117,N_18735);
and UO_827 (O_827,N_19811,N_18690);
xnor UO_828 (O_828,N_18560,N_18493);
and UO_829 (O_829,N_19498,N_18151);
xnor UO_830 (O_830,N_18424,N_18822);
and UO_831 (O_831,N_19642,N_18728);
xor UO_832 (O_832,N_18498,N_18611);
nand UO_833 (O_833,N_18840,N_18172);
nand UO_834 (O_834,N_19564,N_18855);
nor UO_835 (O_835,N_19909,N_18434);
xor UO_836 (O_836,N_19842,N_18829);
and UO_837 (O_837,N_18280,N_19610);
xor UO_838 (O_838,N_18874,N_18400);
xnor UO_839 (O_839,N_18900,N_19963);
nand UO_840 (O_840,N_19676,N_19598);
xor UO_841 (O_841,N_19660,N_18163);
and UO_842 (O_842,N_19289,N_18149);
and UO_843 (O_843,N_19628,N_18895);
xnor UO_844 (O_844,N_19392,N_18768);
xor UO_845 (O_845,N_19060,N_19352);
xor UO_846 (O_846,N_18804,N_19205);
and UO_847 (O_847,N_19887,N_19663);
or UO_848 (O_848,N_19000,N_18178);
and UO_849 (O_849,N_18704,N_19007);
and UO_850 (O_850,N_18563,N_18432);
xor UO_851 (O_851,N_18790,N_19421);
or UO_852 (O_852,N_19871,N_18223);
xnor UO_853 (O_853,N_19283,N_19002);
nor UO_854 (O_854,N_19142,N_19211);
or UO_855 (O_855,N_19668,N_18966);
nand UO_856 (O_856,N_19750,N_19068);
nor UO_857 (O_857,N_18732,N_18350);
and UO_858 (O_858,N_19639,N_19692);
nor UO_859 (O_859,N_19565,N_18414);
nand UO_860 (O_860,N_18444,N_18068);
or UO_861 (O_861,N_18248,N_18311);
and UO_862 (O_862,N_19973,N_18638);
nor UO_863 (O_863,N_18043,N_18473);
nand UO_864 (O_864,N_19694,N_19153);
nand UO_865 (O_865,N_19870,N_19641);
xnor UO_866 (O_866,N_18602,N_18663);
xnor UO_867 (O_867,N_18575,N_18415);
xor UO_868 (O_868,N_18972,N_19783);
or UO_869 (O_869,N_19118,N_18733);
xnor UO_870 (O_870,N_18951,N_19015);
nor UO_871 (O_871,N_19930,N_19661);
and UO_872 (O_872,N_19835,N_18112);
and UO_873 (O_873,N_19860,N_18669);
nor UO_874 (O_874,N_18458,N_19032);
and UO_875 (O_875,N_18320,N_18422);
or UO_876 (O_876,N_18623,N_18487);
nand UO_877 (O_877,N_19547,N_19529);
nand UO_878 (O_878,N_18982,N_18507);
nor UO_879 (O_879,N_18851,N_19970);
nor UO_880 (O_880,N_19867,N_18437);
and UO_881 (O_881,N_19174,N_18776);
and UO_882 (O_882,N_18712,N_19600);
nand UO_883 (O_883,N_19025,N_19841);
and UO_884 (O_884,N_19629,N_19986);
nand UO_885 (O_885,N_18799,N_19357);
and UO_886 (O_886,N_18206,N_19423);
xor UO_887 (O_887,N_18120,N_18428);
or UO_888 (O_888,N_18075,N_19900);
and UO_889 (O_889,N_18296,N_18258);
xnor UO_890 (O_890,N_18753,N_19566);
or UO_891 (O_891,N_19093,N_18291);
xnor UO_892 (O_892,N_18631,N_19760);
xnor UO_893 (O_893,N_18876,N_18880);
nor UO_894 (O_894,N_19531,N_19782);
and UO_895 (O_895,N_19266,N_18449);
or UO_896 (O_896,N_18539,N_18584);
nor UO_897 (O_897,N_18023,N_19254);
and UO_898 (O_898,N_18862,N_19059);
nand UO_899 (O_899,N_18369,N_19658);
nand UO_900 (O_900,N_18243,N_18932);
or UO_901 (O_901,N_18393,N_18020);
and UO_902 (O_902,N_18805,N_18801);
and UO_903 (O_903,N_18591,N_18826);
and UO_904 (O_904,N_18917,N_18052);
nand UO_905 (O_905,N_18708,N_19151);
or UO_906 (O_906,N_19977,N_18281);
xnor UO_907 (O_907,N_18357,N_19999);
or UO_908 (O_908,N_19217,N_18275);
nand UO_909 (O_909,N_19409,N_18271);
and UO_910 (O_910,N_19290,N_18324);
nor UO_911 (O_911,N_19179,N_18956);
nor UO_912 (O_912,N_19838,N_19154);
and UO_913 (O_913,N_18557,N_19101);
and UO_914 (O_914,N_19425,N_19180);
and UO_915 (O_915,N_18945,N_19359);
nand UO_916 (O_916,N_19105,N_18250);
and UO_917 (O_917,N_19805,N_19655);
nand UO_918 (O_918,N_19128,N_19210);
xnor UO_919 (O_919,N_19279,N_18997);
xor UO_920 (O_920,N_18986,N_19621);
or UO_921 (O_921,N_19325,N_19207);
xnor UO_922 (O_922,N_19324,N_19130);
and UO_923 (O_923,N_18159,N_19980);
xor UO_924 (O_924,N_19551,N_19632);
or UO_925 (O_925,N_18894,N_19972);
xor UO_926 (O_926,N_19224,N_18213);
xnor UO_927 (O_927,N_18164,N_18119);
nor UO_928 (O_928,N_18482,N_18096);
nand UO_929 (O_929,N_18312,N_19939);
xnor UO_930 (O_930,N_18865,N_18319);
or UO_931 (O_931,N_18265,N_19954);
nand UO_932 (O_932,N_19759,N_19372);
nor UO_933 (O_933,N_18577,N_18429);
nand UO_934 (O_934,N_18230,N_18508);
and UO_935 (O_935,N_19736,N_18641);
and UO_936 (O_936,N_18356,N_19172);
nand UO_937 (O_937,N_18896,N_18936);
nor UO_938 (O_938,N_19042,N_18988);
nand UO_939 (O_939,N_19914,N_19965);
xnor UO_940 (O_940,N_19148,N_18985);
nand UO_941 (O_941,N_18636,N_18981);
nor UO_942 (O_942,N_19318,N_18308);
nand UO_943 (O_943,N_19313,N_18532);
nand UO_944 (O_944,N_19478,N_19374);
nand UO_945 (O_945,N_19851,N_19331);
nand UO_946 (O_946,N_19561,N_19918);
xnor UO_947 (O_947,N_18943,N_19656);
nor UO_948 (O_948,N_19956,N_18777);
xnor UO_949 (O_949,N_19502,N_18404);
and UO_950 (O_950,N_18684,N_19407);
or UO_951 (O_951,N_18783,N_18228);
xor UO_952 (O_952,N_18215,N_18235);
or UO_953 (O_953,N_18949,N_19903);
nor UO_954 (O_954,N_18063,N_18843);
nor UO_955 (O_955,N_18509,N_18624);
nor UO_956 (O_956,N_19016,N_19054);
and UO_957 (O_957,N_19275,N_19193);
nand UO_958 (O_958,N_19229,N_19670);
nand UO_959 (O_959,N_19271,N_19815);
and UO_960 (O_960,N_19246,N_18727);
nand UO_961 (O_961,N_19544,N_19226);
nor UO_962 (O_962,N_19686,N_19718);
nor UO_963 (O_963,N_19140,N_18578);
or UO_964 (O_964,N_18707,N_18819);
and UO_965 (O_965,N_18011,N_19045);
and UO_966 (O_966,N_19781,N_19683);
xor UO_967 (O_967,N_19094,N_19710);
or UO_968 (O_968,N_18834,N_19705);
xnor UO_969 (O_969,N_19402,N_18906);
nor UO_970 (O_970,N_18283,N_19959);
nand UO_971 (O_971,N_18701,N_18530);
and UO_972 (O_972,N_19720,N_19752);
nor UO_973 (O_973,N_18503,N_18333);
nand UO_974 (O_974,N_18792,N_18722);
nor UO_975 (O_975,N_19050,N_19869);
or UO_976 (O_976,N_19280,N_19820);
nor UO_977 (O_977,N_18032,N_18931);
nor UO_978 (O_978,N_18542,N_19029);
nand UO_979 (O_979,N_19575,N_19278);
nor UO_980 (O_980,N_19573,N_18485);
nor UO_981 (O_981,N_19772,N_19919);
or UO_982 (O_982,N_19135,N_18881);
and UO_983 (O_983,N_19307,N_19749);
xor UO_984 (O_984,N_18890,N_18600);
xnor UO_985 (O_985,N_19257,N_18500);
xor UO_986 (O_986,N_18812,N_19605);
and UO_987 (O_987,N_19989,N_19158);
and UO_988 (O_988,N_19793,N_18537);
or UO_989 (O_989,N_18882,N_18977);
or UO_990 (O_990,N_18625,N_19481);
nor UO_991 (O_991,N_19549,N_19469);
nor UO_992 (O_992,N_19288,N_19219);
nand UO_993 (O_993,N_19046,N_19185);
xnor UO_994 (O_994,N_18289,N_19038);
nand UO_995 (O_995,N_18831,N_18649);
nor UO_996 (O_996,N_18236,N_18266);
and UO_997 (O_997,N_18771,N_19383);
nor UO_998 (O_998,N_19427,N_19376);
nor UO_999 (O_999,N_18184,N_19043);
nor UO_1000 (O_1000,N_19274,N_19544);
or UO_1001 (O_1001,N_19665,N_18882);
nor UO_1002 (O_1002,N_19672,N_19830);
xnor UO_1003 (O_1003,N_19875,N_18047);
and UO_1004 (O_1004,N_19598,N_18827);
and UO_1005 (O_1005,N_18809,N_18827);
and UO_1006 (O_1006,N_18579,N_19921);
and UO_1007 (O_1007,N_19006,N_18850);
nand UO_1008 (O_1008,N_19931,N_18890);
xor UO_1009 (O_1009,N_18088,N_18638);
nand UO_1010 (O_1010,N_18344,N_18110);
nor UO_1011 (O_1011,N_19656,N_19247);
nand UO_1012 (O_1012,N_19280,N_18611);
and UO_1013 (O_1013,N_18037,N_19262);
nand UO_1014 (O_1014,N_18142,N_18512);
nand UO_1015 (O_1015,N_18078,N_18350);
and UO_1016 (O_1016,N_19805,N_18492);
and UO_1017 (O_1017,N_18921,N_18328);
or UO_1018 (O_1018,N_19683,N_18312);
nand UO_1019 (O_1019,N_19882,N_18438);
or UO_1020 (O_1020,N_18967,N_18974);
xnor UO_1021 (O_1021,N_19363,N_18269);
and UO_1022 (O_1022,N_18790,N_18702);
xor UO_1023 (O_1023,N_18102,N_19060);
or UO_1024 (O_1024,N_18225,N_19584);
or UO_1025 (O_1025,N_18792,N_19450);
or UO_1026 (O_1026,N_19405,N_18008);
or UO_1027 (O_1027,N_19602,N_19256);
xnor UO_1028 (O_1028,N_18659,N_19296);
and UO_1029 (O_1029,N_18112,N_19364);
nand UO_1030 (O_1030,N_18858,N_18048);
nor UO_1031 (O_1031,N_18076,N_18328);
xor UO_1032 (O_1032,N_18664,N_19101);
nor UO_1033 (O_1033,N_19828,N_19107);
and UO_1034 (O_1034,N_19163,N_19506);
xnor UO_1035 (O_1035,N_18927,N_18501);
or UO_1036 (O_1036,N_19057,N_19554);
nand UO_1037 (O_1037,N_19730,N_18763);
nand UO_1038 (O_1038,N_18003,N_19171);
xnor UO_1039 (O_1039,N_19325,N_19162);
or UO_1040 (O_1040,N_19823,N_19877);
nor UO_1041 (O_1041,N_19614,N_18453);
xor UO_1042 (O_1042,N_19222,N_18006);
or UO_1043 (O_1043,N_18668,N_19837);
nand UO_1044 (O_1044,N_19588,N_18446);
xor UO_1045 (O_1045,N_18828,N_19056);
nor UO_1046 (O_1046,N_18804,N_18081);
nand UO_1047 (O_1047,N_19414,N_18912);
or UO_1048 (O_1048,N_19945,N_19641);
nand UO_1049 (O_1049,N_19123,N_19532);
xnor UO_1050 (O_1050,N_18810,N_19736);
or UO_1051 (O_1051,N_18569,N_19856);
xnor UO_1052 (O_1052,N_19463,N_18666);
nand UO_1053 (O_1053,N_18993,N_19758);
and UO_1054 (O_1054,N_18394,N_18113);
nand UO_1055 (O_1055,N_18747,N_19059);
nor UO_1056 (O_1056,N_19912,N_18567);
xor UO_1057 (O_1057,N_18803,N_18502);
nand UO_1058 (O_1058,N_18914,N_18233);
and UO_1059 (O_1059,N_18662,N_18180);
nand UO_1060 (O_1060,N_18882,N_18327);
xnor UO_1061 (O_1061,N_18934,N_19291);
xor UO_1062 (O_1062,N_19254,N_19222);
xnor UO_1063 (O_1063,N_18309,N_19409);
nand UO_1064 (O_1064,N_18817,N_18325);
and UO_1065 (O_1065,N_19283,N_18161);
nand UO_1066 (O_1066,N_19405,N_19418);
nand UO_1067 (O_1067,N_18698,N_19733);
or UO_1068 (O_1068,N_19538,N_18257);
nand UO_1069 (O_1069,N_18275,N_19685);
nor UO_1070 (O_1070,N_18369,N_19820);
or UO_1071 (O_1071,N_19120,N_18838);
xnor UO_1072 (O_1072,N_18485,N_19354);
and UO_1073 (O_1073,N_19362,N_18382);
or UO_1074 (O_1074,N_18548,N_19830);
and UO_1075 (O_1075,N_19560,N_18024);
nor UO_1076 (O_1076,N_19132,N_19196);
and UO_1077 (O_1077,N_19517,N_18596);
and UO_1078 (O_1078,N_18439,N_18014);
xnor UO_1079 (O_1079,N_19619,N_18733);
and UO_1080 (O_1080,N_19435,N_18760);
xnor UO_1081 (O_1081,N_19743,N_19134);
or UO_1082 (O_1082,N_18743,N_19862);
and UO_1083 (O_1083,N_18774,N_19276);
and UO_1084 (O_1084,N_19739,N_19392);
or UO_1085 (O_1085,N_19981,N_18907);
xor UO_1086 (O_1086,N_19152,N_19740);
xor UO_1087 (O_1087,N_19701,N_18412);
nand UO_1088 (O_1088,N_18619,N_19455);
xor UO_1089 (O_1089,N_19096,N_18775);
nand UO_1090 (O_1090,N_18725,N_19533);
nor UO_1091 (O_1091,N_18497,N_19567);
nor UO_1092 (O_1092,N_19551,N_18015);
and UO_1093 (O_1093,N_19403,N_19813);
nand UO_1094 (O_1094,N_18490,N_19740);
or UO_1095 (O_1095,N_19392,N_19462);
nand UO_1096 (O_1096,N_19373,N_18965);
and UO_1097 (O_1097,N_19322,N_18004);
nor UO_1098 (O_1098,N_18994,N_18762);
nor UO_1099 (O_1099,N_18560,N_19067);
nand UO_1100 (O_1100,N_19771,N_19809);
or UO_1101 (O_1101,N_18160,N_19676);
nand UO_1102 (O_1102,N_19572,N_18451);
or UO_1103 (O_1103,N_19625,N_19629);
or UO_1104 (O_1104,N_19550,N_18317);
nor UO_1105 (O_1105,N_18904,N_18445);
nor UO_1106 (O_1106,N_19293,N_18982);
nand UO_1107 (O_1107,N_18758,N_19305);
and UO_1108 (O_1108,N_18924,N_18144);
and UO_1109 (O_1109,N_18744,N_19798);
nand UO_1110 (O_1110,N_18440,N_18088);
xnor UO_1111 (O_1111,N_18026,N_19694);
nand UO_1112 (O_1112,N_19402,N_18896);
nor UO_1113 (O_1113,N_18416,N_18937);
and UO_1114 (O_1114,N_19928,N_18509);
and UO_1115 (O_1115,N_18949,N_19636);
or UO_1116 (O_1116,N_19852,N_19197);
or UO_1117 (O_1117,N_18215,N_18814);
xnor UO_1118 (O_1118,N_19425,N_19067);
nand UO_1119 (O_1119,N_19024,N_18290);
xor UO_1120 (O_1120,N_19871,N_18605);
xnor UO_1121 (O_1121,N_18876,N_19007);
xnor UO_1122 (O_1122,N_18662,N_18982);
or UO_1123 (O_1123,N_18508,N_18709);
or UO_1124 (O_1124,N_19985,N_18464);
nor UO_1125 (O_1125,N_19579,N_18551);
nor UO_1126 (O_1126,N_19521,N_19622);
nor UO_1127 (O_1127,N_18329,N_18659);
nand UO_1128 (O_1128,N_18179,N_19654);
and UO_1129 (O_1129,N_18186,N_19700);
or UO_1130 (O_1130,N_19806,N_18175);
xnor UO_1131 (O_1131,N_19598,N_19645);
nand UO_1132 (O_1132,N_19168,N_19549);
nand UO_1133 (O_1133,N_18911,N_18803);
nand UO_1134 (O_1134,N_19454,N_19139);
or UO_1135 (O_1135,N_19854,N_18047);
or UO_1136 (O_1136,N_19650,N_19004);
xor UO_1137 (O_1137,N_18372,N_19854);
xnor UO_1138 (O_1138,N_19710,N_19651);
or UO_1139 (O_1139,N_18217,N_18069);
xnor UO_1140 (O_1140,N_19126,N_19241);
or UO_1141 (O_1141,N_18944,N_19967);
and UO_1142 (O_1142,N_19304,N_18404);
and UO_1143 (O_1143,N_18002,N_19689);
and UO_1144 (O_1144,N_18425,N_19052);
or UO_1145 (O_1145,N_19929,N_18626);
nand UO_1146 (O_1146,N_18969,N_18980);
xnor UO_1147 (O_1147,N_18108,N_19177);
xor UO_1148 (O_1148,N_19664,N_18257);
xor UO_1149 (O_1149,N_19603,N_18537);
or UO_1150 (O_1150,N_19749,N_18942);
or UO_1151 (O_1151,N_18137,N_19142);
or UO_1152 (O_1152,N_18461,N_19587);
nor UO_1153 (O_1153,N_19013,N_19873);
nor UO_1154 (O_1154,N_18743,N_19040);
nand UO_1155 (O_1155,N_18455,N_18196);
or UO_1156 (O_1156,N_19905,N_18957);
nand UO_1157 (O_1157,N_18858,N_18916);
nand UO_1158 (O_1158,N_18352,N_18330);
and UO_1159 (O_1159,N_18703,N_19914);
xor UO_1160 (O_1160,N_18773,N_18657);
and UO_1161 (O_1161,N_18342,N_18897);
or UO_1162 (O_1162,N_19714,N_19759);
nand UO_1163 (O_1163,N_18050,N_18623);
or UO_1164 (O_1164,N_19409,N_18746);
nand UO_1165 (O_1165,N_18233,N_19493);
nor UO_1166 (O_1166,N_19350,N_18716);
nor UO_1167 (O_1167,N_19256,N_19693);
and UO_1168 (O_1168,N_19254,N_18929);
and UO_1169 (O_1169,N_19386,N_18814);
or UO_1170 (O_1170,N_18805,N_18804);
xnor UO_1171 (O_1171,N_19123,N_18420);
and UO_1172 (O_1172,N_19937,N_19038);
nor UO_1173 (O_1173,N_19765,N_19276);
and UO_1174 (O_1174,N_19021,N_18227);
nor UO_1175 (O_1175,N_18419,N_19586);
nand UO_1176 (O_1176,N_19900,N_19351);
nand UO_1177 (O_1177,N_18629,N_19722);
or UO_1178 (O_1178,N_19025,N_19071);
or UO_1179 (O_1179,N_18173,N_19942);
nor UO_1180 (O_1180,N_19452,N_19949);
and UO_1181 (O_1181,N_18339,N_18107);
xor UO_1182 (O_1182,N_18354,N_19012);
nand UO_1183 (O_1183,N_18559,N_18350);
nand UO_1184 (O_1184,N_18632,N_18320);
nand UO_1185 (O_1185,N_19706,N_18141);
or UO_1186 (O_1186,N_19440,N_18334);
and UO_1187 (O_1187,N_18471,N_19964);
xnor UO_1188 (O_1188,N_19656,N_18962);
or UO_1189 (O_1189,N_19671,N_18897);
nor UO_1190 (O_1190,N_19957,N_19879);
and UO_1191 (O_1191,N_19879,N_18812);
nand UO_1192 (O_1192,N_19385,N_18591);
xor UO_1193 (O_1193,N_18453,N_18144);
nor UO_1194 (O_1194,N_19565,N_18197);
nand UO_1195 (O_1195,N_18283,N_18109);
nor UO_1196 (O_1196,N_19475,N_19406);
or UO_1197 (O_1197,N_19381,N_19698);
and UO_1198 (O_1198,N_18295,N_18464);
nor UO_1199 (O_1199,N_18292,N_19076);
or UO_1200 (O_1200,N_19175,N_19302);
nor UO_1201 (O_1201,N_18522,N_18871);
nand UO_1202 (O_1202,N_19641,N_19093);
and UO_1203 (O_1203,N_18327,N_18724);
and UO_1204 (O_1204,N_19831,N_18970);
and UO_1205 (O_1205,N_19738,N_19990);
and UO_1206 (O_1206,N_19410,N_19841);
xnor UO_1207 (O_1207,N_19268,N_18372);
and UO_1208 (O_1208,N_18600,N_19727);
xnor UO_1209 (O_1209,N_19650,N_18758);
nand UO_1210 (O_1210,N_18589,N_19032);
and UO_1211 (O_1211,N_19599,N_18890);
nand UO_1212 (O_1212,N_18620,N_19937);
or UO_1213 (O_1213,N_19902,N_18788);
or UO_1214 (O_1214,N_18608,N_18795);
or UO_1215 (O_1215,N_18453,N_18143);
and UO_1216 (O_1216,N_18371,N_18149);
or UO_1217 (O_1217,N_19879,N_19934);
and UO_1218 (O_1218,N_18334,N_18639);
nor UO_1219 (O_1219,N_19688,N_18890);
nand UO_1220 (O_1220,N_19577,N_19703);
nand UO_1221 (O_1221,N_18560,N_18686);
or UO_1222 (O_1222,N_18452,N_18871);
xor UO_1223 (O_1223,N_18869,N_19771);
and UO_1224 (O_1224,N_19617,N_19977);
xor UO_1225 (O_1225,N_19960,N_18931);
xor UO_1226 (O_1226,N_18036,N_18242);
and UO_1227 (O_1227,N_19627,N_19888);
nor UO_1228 (O_1228,N_19634,N_19683);
and UO_1229 (O_1229,N_18666,N_18656);
xnor UO_1230 (O_1230,N_18986,N_18943);
and UO_1231 (O_1231,N_19500,N_18572);
xor UO_1232 (O_1232,N_19233,N_18307);
nand UO_1233 (O_1233,N_18052,N_19703);
nor UO_1234 (O_1234,N_19524,N_19175);
nor UO_1235 (O_1235,N_18657,N_18377);
or UO_1236 (O_1236,N_19937,N_19300);
or UO_1237 (O_1237,N_18876,N_19824);
xor UO_1238 (O_1238,N_18537,N_18290);
nor UO_1239 (O_1239,N_18839,N_19147);
xor UO_1240 (O_1240,N_18740,N_19166);
nand UO_1241 (O_1241,N_18522,N_18086);
nand UO_1242 (O_1242,N_18046,N_18343);
xnor UO_1243 (O_1243,N_18196,N_19619);
or UO_1244 (O_1244,N_19546,N_18168);
xor UO_1245 (O_1245,N_18972,N_19470);
and UO_1246 (O_1246,N_19288,N_19852);
and UO_1247 (O_1247,N_19377,N_19691);
xor UO_1248 (O_1248,N_19682,N_19327);
nand UO_1249 (O_1249,N_18448,N_19076);
nand UO_1250 (O_1250,N_18257,N_19587);
and UO_1251 (O_1251,N_18175,N_18111);
and UO_1252 (O_1252,N_18407,N_18725);
nand UO_1253 (O_1253,N_18036,N_19016);
xnor UO_1254 (O_1254,N_19838,N_18754);
xor UO_1255 (O_1255,N_19429,N_19645);
nor UO_1256 (O_1256,N_18826,N_18329);
nor UO_1257 (O_1257,N_18068,N_19022);
xnor UO_1258 (O_1258,N_19919,N_19900);
nor UO_1259 (O_1259,N_18460,N_19173);
nor UO_1260 (O_1260,N_19632,N_18045);
or UO_1261 (O_1261,N_19912,N_19102);
xor UO_1262 (O_1262,N_19256,N_18017);
or UO_1263 (O_1263,N_19637,N_18777);
nor UO_1264 (O_1264,N_18175,N_19670);
xor UO_1265 (O_1265,N_19402,N_18793);
xor UO_1266 (O_1266,N_18741,N_18264);
nor UO_1267 (O_1267,N_18465,N_18059);
and UO_1268 (O_1268,N_18169,N_19386);
nand UO_1269 (O_1269,N_19733,N_18381);
or UO_1270 (O_1270,N_19622,N_18085);
or UO_1271 (O_1271,N_19949,N_19797);
nand UO_1272 (O_1272,N_19664,N_18854);
nand UO_1273 (O_1273,N_18782,N_18632);
xnor UO_1274 (O_1274,N_19328,N_18022);
nand UO_1275 (O_1275,N_19342,N_18742);
nor UO_1276 (O_1276,N_18309,N_19430);
and UO_1277 (O_1277,N_19759,N_19529);
or UO_1278 (O_1278,N_19432,N_19073);
or UO_1279 (O_1279,N_19980,N_18235);
nand UO_1280 (O_1280,N_19608,N_18385);
nand UO_1281 (O_1281,N_18648,N_19411);
and UO_1282 (O_1282,N_19165,N_19835);
nand UO_1283 (O_1283,N_19015,N_19904);
or UO_1284 (O_1284,N_19183,N_19533);
or UO_1285 (O_1285,N_18353,N_18990);
xnor UO_1286 (O_1286,N_19766,N_18040);
or UO_1287 (O_1287,N_19568,N_19642);
and UO_1288 (O_1288,N_18723,N_18597);
nor UO_1289 (O_1289,N_18993,N_19755);
xor UO_1290 (O_1290,N_19599,N_19472);
xor UO_1291 (O_1291,N_19199,N_19092);
xnor UO_1292 (O_1292,N_19109,N_19110);
xor UO_1293 (O_1293,N_18463,N_18855);
and UO_1294 (O_1294,N_18477,N_19103);
or UO_1295 (O_1295,N_18794,N_19259);
nand UO_1296 (O_1296,N_19910,N_19762);
nand UO_1297 (O_1297,N_19141,N_19965);
or UO_1298 (O_1298,N_18011,N_19344);
nand UO_1299 (O_1299,N_19789,N_19568);
and UO_1300 (O_1300,N_18407,N_19581);
and UO_1301 (O_1301,N_19481,N_18468);
or UO_1302 (O_1302,N_18975,N_19127);
nand UO_1303 (O_1303,N_19411,N_19271);
and UO_1304 (O_1304,N_19435,N_18629);
nor UO_1305 (O_1305,N_18895,N_18683);
and UO_1306 (O_1306,N_18537,N_18797);
or UO_1307 (O_1307,N_19502,N_18301);
nor UO_1308 (O_1308,N_19757,N_19023);
nor UO_1309 (O_1309,N_19024,N_19242);
xnor UO_1310 (O_1310,N_19909,N_19904);
and UO_1311 (O_1311,N_19674,N_18045);
nand UO_1312 (O_1312,N_19246,N_18591);
nor UO_1313 (O_1313,N_19670,N_18875);
xor UO_1314 (O_1314,N_18119,N_18305);
and UO_1315 (O_1315,N_18224,N_18698);
xor UO_1316 (O_1316,N_19220,N_19267);
and UO_1317 (O_1317,N_18864,N_19276);
nand UO_1318 (O_1318,N_18783,N_19562);
and UO_1319 (O_1319,N_19015,N_19854);
xor UO_1320 (O_1320,N_19119,N_19384);
or UO_1321 (O_1321,N_18238,N_19961);
and UO_1322 (O_1322,N_19400,N_18028);
or UO_1323 (O_1323,N_19945,N_19381);
xor UO_1324 (O_1324,N_19365,N_18645);
nand UO_1325 (O_1325,N_18128,N_19176);
nand UO_1326 (O_1326,N_18174,N_18814);
and UO_1327 (O_1327,N_18669,N_18048);
or UO_1328 (O_1328,N_18088,N_19750);
xnor UO_1329 (O_1329,N_18276,N_19152);
nand UO_1330 (O_1330,N_18423,N_18347);
xnor UO_1331 (O_1331,N_19686,N_18198);
nor UO_1332 (O_1332,N_19901,N_18261);
xnor UO_1333 (O_1333,N_18824,N_18988);
nand UO_1334 (O_1334,N_18394,N_18820);
and UO_1335 (O_1335,N_19776,N_19958);
xnor UO_1336 (O_1336,N_19355,N_19409);
nor UO_1337 (O_1337,N_18937,N_18614);
nor UO_1338 (O_1338,N_18967,N_19434);
nor UO_1339 (O_1339,N_19455,N_19978);
or UO_1340 (O_1340,N_19172,N_19622);
xnor UO_1341 (O_1341,N_18069,N_18369);
nor UO_1342 (O_1342,N_18553,N_18242);
nor UO_1343 (O_1343,N_19394,N_18150);
nand UO_1344 (O_1344,N_18888,N_18708);
nand UO_1345 (O_1345,N_18253,N_19238);
or UO_1346 (O_1346,N_18730,N_18676);
nor UO_1347 (O_1347,N_19265,N_19310);
xnor UO_1348 (O_1348,N_19918,N_18514);
nand UO_1349 (O_1349,N_19606,N_18139);
or UO_1350 (O_1350,N_18099,N_19376);
nand UO_1351 (O_1351,N_18132,N_18140);
or UO_1352 (O_1352,N_18494,N_19698);
or UO_1353 (O_1353,N_18469,N_18729);
nor UO_1354 (O_1354,N_19783,N_19334);
or UO_1355 (O_1355,N_19324,N_19212);
nor UO_1356 (O_1356,N_19610,N_18898);
or UO_1357 (O_1357,N_18404,N_18980);
and UO_1358 (O_1358,N_19807,N_18741);
nand UO_1359 (O_1359,N_19227,N_19665);
and UO_1360 (O_1360,N_18717,N_18410);
nor UO_1361 (O_1361,N_19469,N_19315);
nor UO_1362 (O_1362,N_18665,N_18437);
or UO_1363 (O_1363,N_19415,N_19485);
or UO_1364 (O_1364,N_19993,N_19312);
xnor UO_1365 (O_1365,N_19150,N_19894);
nor UO_1366 (O_1366,N_19838,N_18889);
nor UO_1367 (O_1367,N_18009,N_19505);
or UO_1368 (O_1368,N_19046,N_19421);
nor UO_1369 (O_1369,N_19075,N_19355);
or UO_1370 (O_1370,N_19939,N_19593);
nand UO_1371 (O_1371,N_19613,N_18817);
or UO_1372 (O_1372,N_19167,N_18113);
nand UO_1373 (O_1373,N_19060,N_18361);
or UO_1374 (O_1374,N_18692,N_18245);
xor UO_1375 (O_1375,N_18644,N_19468);
nor UO_1376 (O_1376,N_18314,N_18620);
nand UO_1377 (O_1377,N_19929,N_19353);
or UO_1378 (O_1378,N_18137,N_18801);
nor UO_1379 (O_1379,N_19811,N_19745);
nor UO_1380 (O_1380,N_19128,N_18273);
nand UO_1381 (O_1381,N_19524,N_18341);
nor UO_1382 (O_1382,N_18270,N_19996);
nor UO_1383 (O_1383,N_18353,N_18221);
nor UO_1384 (O_1384,N_18555,N_19834);
nor UO_1385 (O_1385,N_18666,N_18454);
nand UO_1386 (O_1386,N_18962,N_19633);
or UO_1387 (O_1387,N_19055,N_19872);
nor UO_1388 (O_1388,N_19114,N_19885);
and UO_1389 (O_1389,N_19094,N_19636);
or UO_1390 (O_1390,N_19703,N_18290);
xor UO_1391 (O_1391,N_18797,N_18380);
or UO_1392 (O_1392,N_19039,N_18673);
xnor UO_1393 (O_1393,N_19732,N_19573);
or UO_1394 (O_1394,N_18103,N_18247);
and UO_1395 (O_1395,N_19830,N_19154);
xnor UO_1396 (O_1396,N_19065,N_19326);
xnor UO_1397 (O_1397,N_19026,N_19656);
or UO_1398 (O_1398,N_18704,N_18309);
nor UO_1399 (O_1399,N_18647,N_18150);
nand UO_1400 (O_1400,N_18529,N_18493);
nand UO_1401 (O_1401,N_19793,N_19817);
and UO_1402 (O_1402,N_19740,N_18828);
xnor UO_1403 (O_1403,N_18946,N_19694);
xnor UO_1404 (O_1404,N_19377,N_19580);
and UO_1405 (O_1405,N_18082,N_19657);
xnor UO_1406 (O_1406,N_18399,N_18392);
and UO_1407 (O_1407,N_19586,N_19811);
nor UO_1408 (O_1408,N_18088,N_18862);
nand UO_1409 (O_1409,N_18814,N_18671);
xnor UO_1410 (O_1410,N_19278,N_19588);
and UO_1411 (O_1411,N_19381,N_19494);
or UO_1412 (O_1412,N_18653,N_18044);
and UO_1413 (O_1413,N_19920,N_19986);
nand UO_1414 (O_1414,N_18562,N_19293);
or UO_1415 (O_1415,N_19456,N_18935);
nand UO_1416 (O_1416,N_18429,N_18304);
and UO_1417 (O_1417,N_18089,N_19141);
nor UO_1418 (O_1418,N_18498,N_19425);
nand UO_1419 (O_1419,N_19444,N_19183);
nand UO_1420 (O_1420,N_19556,N_19323);
and UO_1421 (O_1421,N_19215,N_19298);
nand UO_1422 (O_1422,N_19717,N_18768);
or UO_1423 (O_1423,N_18059,N_18582);
nand UO_1424 (O_1424,N_18092,N_19649);
or UO_1425 (O_1425,N_18499,N_18957);
nor UO_1426 (O_1426,N_18635,N_19579);
and UO_1427 (O_1427,N_19316,N_19207);
nor UO_1428 (O_1428,N_18855,N_18393);
or UO_1429 (O_1429,N_19807,N_18540);
nand UO_1430 (O_1430,N_19793,N_19346);
xnor UO_1431 (O_1431,N_18309,N_18483);
nor UO_1432 (O_1432,N_19134,N_19897);
or UO_1433 (O_1433,N_18108,N_18114);
nand UO_1434 (O_1434,N_18920,N_18577);
and UO_1435 (O_1435,N_18865,N_18355);
nor UO_1436 (O_1436,N_18195,N_19235);
and UO_1437 (O_1437,N_18980,N_18565);
and UO_1438 (O_1438,N_19384,N_18593);
nand UO_1439 (O_1439,N_19589,N_19266);
nand UO_1440 (O_1440,N_18854,N_18810);
nor UO_1441 (O_1441,N_19832,N_19540);
or UO_1442 (O_1442,N_18867,N_19669);
xor UO_1443 (O_1443,N_19372,N_19922);
or UO_1444 (O_1444,N_18541,N_19717);
xnor UO_1445 (O_1445,N_19608,N_18907);
xnor UO_1446 (O_1446,N_18634,N_18578);
nor UO_1447 (O_1447,N_18819,N_19224);
and UO_1448 (O_1448,N_18787,N_18254);
xor UO_1449 (O_1449,N_18678,N_19787);
and UO_1450 (O_1450,N_19596,N_19328);
nor UO_1451 (O_1451,N_19833,N_19449);
and UO_1452 (O_1452,N_19854,N_19208);
nor UO_1453 (O_1453,N_18843,N_18971);
nand UO_1454 (O_1454,N_18261,N_18590);
xor UO_1455 (O_1455,N_19870,N_18554);
and UO_1456 (O_1456,N_18217,N_19706);
nor UO_1457 (O_1457,N_19578,N_18013);
or UO_1458 (O_1458,N_19592,N_19968);
and UO_1459 (O_1459,N_18450,N_18636);
nand UO_1460 (O_1460,N_18205,N_18715);
and UO_1461 (O_1461,N_19899,N_18130);
or UO_1462 (O_1462,N_19280,N_19769);
and UO_1463 (O_1463,N_18598,N_18205);
and UO_1464 (O_1464,N_19262,N_18375);
or UO_1465 (O_1465,N_19217,N_19805);
and UO_1466 (O_1466,N_19022,N_19966);
or UO_1467 (O_1467,N_19030,N_19359);
xor UO_1468 (O_1468,N_19609,N_19290);
and UO_1469 (O_1469,N_19519,N_19687);
nand UO_1470 (O_1470,N_18365,N_19207);
xnor UO_1471 (O_1471,N_19877,N_18987);
nor UO_1472 (O_1472,N_18850,N_19377);
or UO_1473 (O_1473,N_18088,N_19939);
and UO_1474 (O_1474,N_19504,N_19433);
or UO_1475 (O_1475,N_19159,N_18019);
nor UO_1476 (O_1476,N_19824,N_18358);
nor UO_1477 (O_1477,N_19209,N_19698);
nand UO_1478 (O_1478,N_19432,N_18952);
xor UO_1479 (O_1479,N_19593,N_19401);
nor UO_1480 (O_1480,N_19927,N_19069);
and UO_1481 (O_1481,N_19102,N_19446);
nor UO_1482 (O_1482,N_18708,N_18921);
and UO_1483 (O_1483,N_18114,N_18869);
nor UO_1484 (O_1484,N_19758,N_18267);
nand UO_1485 (O_1485,N_19572,N_18743);
or UO_1486 (O_1486,N_18231,N_19216);
and UO_1487 (O_1487,N_18544,N_19999);
or UO_1488 (O_1488,N_19307,N_19353);
nor UO_1489 (O_1489,N_18650,N_18623);
or UO_1490 (O_1490,N_18557,N_19069);
and UO_1491 (O_1491,N_18739,N_18066);
and UO_1492 (O_1492,N_19462,N_18990);
nor UO_1493 (O_1493,N_19360,N_19132);
nor UO_1494 (O_1494,N_18175,N_18072);
or UO_1495 (O_1495,N_18754,N_19719);
or UO_1496 (O_1496,N_19479,N_18069);
nor UO_1497 (O_1497,N_19829,N_19328);
or UO_1498 (O_1498,N_19766,N_18353);
nor UO_1499 (O_1499,N_19874,N_19659);
nand UO_1500 (O_1500,N_18824,N_18808);
nand UO_1501 (O_1501,N_19717,N_19720);
nand UO_1502 (O_1502,N_19565,N_18291);
and UO_1503 (O_1503,N_18806,N_18953);
nor UO_1504 (O_1504,N_19508,N_18556);
and UO_1505 (O_1505,N_19064,N_19524);
nor UO_1506 (O_1506,N_19912,N_18830);
nor UO_1507 (O_1507,N_18721,N_19419);
and UO_1508 (O_1508,N_18029,N_19006);
and UO_1509 (O_1509,N_19192,N_19410);
nand UO_1510 (O_1510,N_19634,N_18872);
and UO_1511 (O_1511,N_18489,N_19301);
or UO_1512 (O_1512,N_19395,N_19812);
or UO_1513 (O_1513,N_19900,N_18258);
nand UO_1514 (O_1514,N_18319,N_19056);
xor UO_1515 (O_1515,N_19547,N_18524);
xor UO_1516 (O_1516,N_18605,N_19975);
xnor UO_1517 (O_1517,N_18749,N_19813);
nor UO_1518 (O_1518,N_18561,N_18990);
nor UO_1519 (O_1519,N_19495,N_19655);
nor UO_1520 (O_1520,N_19188,N_18599);
or UO_1521 (O_1521,N_18774,N_18511);
xnor UO_1522 (O_1522,N_19470,N_19066);
and UO_1523 (O_1523,N_18584,N_19751);
nand UO_1524 (O_1524,N_19160,N_19584);
nor UO_1525 (O_1525,N_18451,N_18755);
or UO_1526 (O_1526,N_18817,N_19471);
xnor UO_1527 (O_1527,N_18470,N_19674);
nor UO_1528 (O_1528,N_18698,N_19013);
nor UO_1529 (O_1529,N_18601,N_19635);
xnor UO_1530 (O_1530,N_18531,N_18471);
nor UO_1531 (O_1531,N_19122,N_19644);
nor UO_1532 (O_1532,N_18273,N_19029);
xor UO_1533 (O_1533,N_19993,N_18216);
and UO_1534 (O_1534,N_18323,N_18460);
nor UO_1535 (O_1535,N_19190,N_19865);
nand UO_1536 (O_1536,N_19878,N_19695);
nor UO_1537 (O_1537,N_19339,N_19485);
or UO_1538 (O_1538,N_19924,N_18487);
or UO_1539 (O_1539,N_18443,N_19418);
or UO_1540 (O_1540,N_18569,N_19157);
or UO_1541 (O_1541,N_18911,N_18734);
and UO_1542 (O_1542,N_18071,N_19359);
xnor UO_1543 (O_1543,N_18514,N_18856);
and UO_1544 (O_1544,N_18714,N_19192);
or UO_1545 (O_1545,N_18637,N_19315);
or UO_1546 (O_1546,N_19026,N_19216);
or UO_1547 (O_1547,N_18311,N_18424);
xor UO_1548 (O_1548,N_19212,N_18659);
and UO_1549 (O_1549,N_19076,N_18078);
nor UO_1550 (O_1550,N_18400,N_19813);
xor UO_1551 (O_1551,N_19788,N_18232);
xor UO_1552 (O_1552,N_19445,N_18930);
xnor UO_1553 (O_1553,N_18260,N_19724);
nor UO_1554 (O_1554,N_19896,N_18414);
nor UO_1555 (O_1555,N_18172,N_18592);
nor UO_1556 (O_1556,N_19765,N_18104);
or UO_1557 (O_1557,N_19583,N_18676);
nor UO_1558 (O_1558,N_19389,N_19065);
nand UO_1559 (O_1559,N_19659,N_18568);
and UO_1560 (O_1560,N_19989,N_19872);
nand UO_1561 (O_1561,N_18846,N_19908);
nand UO_1562 (O_1562,N_19764,N_18481);
xnor UO_1563 (O_1563,N_18724,N_19158);
nand UO_1564 (O_1564,N_19093,N_18830);
xor UO_1565 (O_1565,N_19353,N_19101);
nor UO_1566 (O_1566,N_18560,N_19821);
xor UO_1567 (O_1567,N_18410,N_18002);
or UO_1568 (O_1568,N_19846,N_18882);
and UO_1569 (O_1569,N_18877,N_18309);
or UO_1570 (O_1570,N_19758,N_19776);
xnor UO_1571 (O_1571,N_19628,N_19963);
or UO_1572 (O_1572,N_18466,N_18850);
or UO_1573 (O_1573,N_19263,N_19605);
xor UO_1574 (O_1574,N_19820,N_18877);
nand UO_1575 (O_1575,N_19114,N_18921);
nor UO_1576 (O_1576,N_18828,N_18478);
nand UO_1577 (O_1577,N_19995,N_18375);
nor UO_1578 (O_1578,N_18719,N_19595);
nand UO_1579 (O_1579,N_19630,N_19117);
and UO_1580 (O_1580,N_18000,N_18029);
and UO_1581 (O_1581,N_19904,N_19405);
nand UO_1582 (O_1582,N_19497,N_18178);
and UO_1583 (O_1583,N_19110,N_19454);
or UO_1584 (O_1584,N_18699,N_18650);
or UO_1585 (O_1585,N_19024,N_18089);
nand UO_1586 (O_1586,N_19721,N_19539);
xnor UO_1587 (O_1587,N_18471,N_19199);
nand UO_1588 (O_1588,N_19091,N_18691);
nand UO_1589 (O_1589,N_19893,N_18434);
nand UO_1590 (O_1590,N_18406,N_18046);
and UO_1591 (O_1591,N_18900,N_19571);
and UO_1592 (O_1592,N_18771,N_19860);
or UO_1593 (O_1593,N_19124,N_18704);
or UO_1594 (O_1594,N_19196,N_18623);
xnor UO_1595 (O_1595,N_18513,N_19048);
xor UO_1596 (O_1596,N_19812,N_18948);
and UO_1597 (O_1597,N_18536,N_19667);
or UO_1598 (O_1598,N_18238,N_19344);
nor UO_1599 (O_1599,N_18075,N_18793);
xor UO_1600 (O_1600,N_19335,N_19255);
nor UO_1601 (O_1601,N_18731,N_18392);
or UO_1602 (O_1602,N_19805,N_18665);
and UO_1603 (O_1603,N_19553,N_19921);
and UO_1604 (O_1604,N_19008,N_18813);
nand UO_1605 (O_1605,N_19643,N_19936);
xor UO_1606 (O_1606,N_19399,N_19654);
nor UO_1607 (O_1607,N_18109,N_19012);
and UO_1608 (O_1608,N_19586,N_18991);
xnor UO_1609 (O_1609,N_19817,N_19814);
xnor UO_1610 (O_1610,N_18942,N_19617);
or UO_1611 (O_1611,N_19245,N_18721);
or UO_1612 (O_1612,N_18092,N_18603);
nor UO_1613 (O_1613,N_19195,N_19440);
or UO_1614 (O_1614,N_18463,N_19636);
or UO_1615 (O_1615,N_18771,N_18227);
nand UO_1616 (O_1616,N_18842,N_19865);
and UO_1617 (O_1617,N_19437,N_18293);
or UO_1618 (O_1618,N_19373,N_18829);
nor UO_1619 (O_1619,N_19096,N_18472);
nor UO_1620 (O_1620,N_18746,N_19023);
xor UO_1621 (O_1621,N_19512,N_19162);
or UO_1622 (O_1622,N_18540,N_18782);
nand UO_1623 (O_1623,N_19370,N_19223);
xnor UO_1624 (O_1624,N_19664,N_18139);
or UO_1625 (O_1625,N_18429,N_18513);
or UO_1626 (O_1626,N_19423,N_19062);
nand UO_1627 (O_1627,N_19544,N_19023);
xor UO_1628 (O_1628,N_18180,N_18271);
nand UO_1629 (O_1629,N_19442,N_19524);
nand UO_1630 (O_1630,N_19751,N_19306);
or UO_1631 (O_1631,N_18649,N_18128);
nand UO_1632 (O_1632,N_19119,N_19239);
nor UO_1633 (O_1633,N_19822,N_19424);
nor UO_1634 (O_1634,N_19836,N_18767);
nand UO_1635 (O_1635,N_19039,N_18987);
and UO_1636 (O_1636,N_18925,N_19159);
xnor UO_1637 (O_1637,N_18321,N_19890);
nor UO_1638 (O_1638,N_19063,N_18815);
or UO_1639 (O_1639,N_19339,N_19177);
nand UO_1640 (O_1640,N_19581,N_18221);
nor UO_1641 (O_1641,N_19582,N_18361);
xnor UO_1642 (O_1642,N_19218,N_19361);
nor UO_1643 (O_1643,N_19304,N_18313);
and UO_1644 (O_1644,N_18865,N_19525);
and UO_1645 (O_1645,N_18553,N_18916);
or UO_1646 (O_1646,N_19135,N_19995);
or UO_1647 (O_1647,N_18646,N_19122);
nor UO_1648 (O_1648,N_19280,N_18517);
nand UO_1649 (O_1649,N_19931,N_18692);
xnor UO_1650 (O_1650,N_18657,N_18694);
xnor UO_1651 (O_1651,N_18593,N_19138);
nor UO_1652 (O_1652,N_19551,N_19778);
nand UO_1653 (O_1653,N_18905,N_19185);
nand UO_1654 (O_1654,N_19619,N_18940);
nor UO_1655 (O_1655,N_19911,N_18844);
nand UO_1656 (O_1656,N_18790,N_19059);
and UO_1657 (O_1657,N_19338,N_18672);
xor UO_1658 (O_1658,N_18988,N_19858);
and UO_1659 (O_1659,N_19401,N_18468);
and UO_1660 (O_1660,N_19387,N_18653);
nor UO_1661 (O_1661,N_19176,N_19802);
xnor UO_1662 (O_1662,N_18030,N_19141);
xor UO_1663 (O_1663,N_19862,N_19857);
nand UO_1664 (O_1664,N_18401,N_18042);
and UO_1665 (O_1665,N_19691,N_18776);
nand UO_1666 (O_1666,N_19032,N_19657);
or UO_1667 (O_1667,N_18703,N_18617);
nor UO_1668 (O_1668,N_19246,N_19387);
and UO_1669 (O_1669,N_19748,N_18783);
or UO_1670 (O_1670,N_18388,N_18099);
nand UO_1671 (O_1671,N_19334,N_19632);
and UO_1672 (O_1672,N_19093,N_18021);
nor UO_1673 (O_1673,N_19991,N_19310);
and UO_1674 (O_1674,N_18372,N_19664);
nand UO_1675 (O_1675,N_18077,N_18508);
nor UO_1676 (O_1676,N_18602,N_19795);
nand UO_1677 (O_1677,N_18848,N_18275);
xor UO_1678 (O_1678,N_18366,N_19969);
xnor UO_1679 (O_1679,N_18856,N_19271);
xor UO_1680 (O_1680,N_18979,N_18931);
nand UO_1681 (O_1681,N_19498,N_18361);
nor UO_1682 (O_1682,N_18780,N_18582);
and UO_1683 (O_1683,N_19154,N_18319);
or UO_1684 (O_1684,N_19115,N_18331);
xnor UO_1685 (O_1685,N_18064,N_18892);
xnor UO_1686 (O_1686,N_19670,N_18765);
nand UO_1687 (O_1687,N_19927,N_18709);
xor UO_1688 (O_1688,N_19073,N_19908);
xor UO_1689 (O_1689,N_19457,N_18592);
and UO_1690 (O_1690,N_19092,N_18003);
or UO_1691 (O_1691,N_19305,N_18207);
or UO_1692 (O_1692,N_19880,N_19199);
nor UO_1693 (O_1693,N_18622,N_18818);
or UO_1694 (O_1694,N_19665,N_18068);
or UO_1695 (O_1695,N_18854,N_19785);
and UO_1696 (O_1696,N_18125,N_19636);
and UO_1697 (O_1697,N_19894,N_18948);
and UO_1698 (O_1698,N_19373,N_19686);
nand UO_1699 (O_1699,N_18700,N_18579);
nand UO_1700 (O_1700,N_19855,N_18358);
nor UO_1701 (O_1701,N_19899,N_19491);
or UO_1702 (O_1702,N_19463,N_18496);
nor UO_1703 (O_1703,N_18146,N_18958);
nand UO_1704 (O_1704,N_18905,N_19832);
xor UO_1705 (O_1705,N_18447,N_19407);
nand UO_1706 (O_1706,N_19243,N_18670);
xnor UO_1707 (O_1707,N_19287,N_18963);
nand UO_1708 (O_1708,N_18749,N_19670);
or UO_1709 (O_1709,N_19588,N_19451);
and UO_1710 (O_1710,N_19980,N_18457);
nand UO_1711 (O_1711,N_19003,N_18534);
or UO_1712 (O_1712,N_18531,N_19305);
or UO_1713 (O_1713,N_18581,N_18191);
and UO_1714 (O_1714,N_19050,N_19333);
xnor UO_1715 (O_1715,N_18926,N_18927);
nor UO_1716 (O_1716,N_19671,N_19335);
xnor UO_1717 (O_1717,N_18286,N_18626);
or UO_1718 (O_1718,N_19485,N_19021);
or UO_1719 (O_1719,N_18174,N_18505);
xnor UO_1720 (O_1720,N_19363,N_18127);
nor UO_1721 (O_1721,N_18465,N_18927);
nor UO_1722 (O_1722,N_19974,N_19043);
or UO_1723 (O_1723,N_19567,N_19790);
or UO_1724 (O_1724,N_19101,N_18207);
xor UO_1725 (O_1725,N_19879,N_19688);
xor UO_1726 (O_1726,N_19799,N_18143);
and UO_1727 (O_1727,N_18081,N_18470);
or UO_1728 (O_1728,N_18373,N_19665);
nor UO_1729 (O_1729,N_19438,N_19041);
nand UO_1730 (O_1730,N_18627,N_19576);
nand UO_1731 (O_1731,N_18065,N_19129);
xnor UO_1732 (O_1732,N_19346,N_19808);
nand UO_1733 (O_1733,N_19937,N_19130);
or UO_1734 (O_1734,N_18240,N_18937);
or UO_1735 (O_1735,N_19319,N_19571);
nand UO_1736 (O_1736,N_19220,N_19559);
or UO_1737 (O_1737,N_18177,N_18839);
or UO_1738 (O_1738,N_19409,N_18425);
nor UO_1739 (O_1739,N_18118,N_18318);
or UO_1740 (O_1740,N_19948,N_19260);
nand UO_1741 (O_1741,N_19904,N_18148);
xor UO_1742 (O_1742,N_19972,N_18712);
nand UO_1743 (O_1743,N_19910,N_19824);
or UO_1744 (O_1744,N_19617,N_19126);
or UO_1745 (O_1745,N_19854,N_19458);
nor UO_1746 (O_1746,N_18652,N_18077);
xor UO_1747 (O_1747,N_18130,N_19856);
nor UO_1748 (O_1748,N_19006,N_19797);
nor UO_1749 (O_1749,N_19571,N_19954);
or UO_1750 (O_1750,N_19883,N_19478);
or UO_1751 (O_1751,N_18995,N_18438);
nor UO_1752 (O_1752,N_19708,N_18203);
or UO_1753 (O_1753,N_19695,N_18429);
and UO_1754 (O_1754,N_19467,N_19424);
nand UO_1755 (O_1755,N_19318,N_19794);
nor UO_1756 (O_1756,N_19088,N_18240);
nor UO_1757 (O_1757,N_18557,N_18030);
nor UO_1758 (O_1758,N_19734,N_19119);
xnor UO_1759 (O_1759,N_18448,N_18943);
nand UO_1760 (O_1760,N_19642,N_18915);
or UO_1761 (O_1761,N_18530,N_18862);
nand UO_1762 (O_1762,N_19942,N_19820);
nor UO_1763 (O_1763,N_18574,N_18486);
nor UO_1764 (O_1764,N_18059,N_19996);
nand UO_1765 (O_1765,N_18252,N_19325);
nand UO_1766 (O_1766,N_18626,N_18874);
nor UO_1767 (O_1767,N_19768,N_19892);
nor UO_1768 (O_1768,N_19982,N_19308);
nand UO_1769 (O_1769,N_19505,N_18765);
nand UO_1770 (O_1770,N_19643,N_18215);
nand UO_1771 (O_1771,N_18123,N_18667);
or UO_1772 (O_1772,N_18847,N_19693);
or UO_1773 (O_1773,N_18310,N_18316);
or UO_1774 (O_1774,N_19459,N_19733);
and UO_1775 (O_1775,N_19428,N_19486);
and UO_1776 (O_1776,N_19787,N_19534);
and UO_1777 (O_1777,N_19159,N_19605);
nor UO_1778 (O_1778,N_19186,N_19294);
nand UO_1779 (O_1779,N_18732,N_19153);
xor UO_1780 (O_1780,N_19366,N_19986);
or UO_1781 (O_1781,N_18723,N_18163);
or UO_1782 (O_1782,N_19903,N_18536);
nand UO_1783 (O_1783,N_18599,N_18693);
nand UO_1784 (O_1784,N_19295,N_19923);
xnor UO_1785 (O_1785,N_19235,N_18985);
nor UO_1786 (O_1786,N_18815,N_18255);
or UO_1787 (O_1787,N_18692,N_19164);
and UO_1788 (O_1788,N_19342,N_19405);
nor UO_1789 (O_1789,N_18033,N_18690);
xnor UO_1790 (O_1790,N_18359,N_18675);
or UO_1791 (O_1791,N_18969,N_18132);
and UO_1792 (O_1792,N_18758,N_19311);
nor UO_1793 (O_1793,N_18342,N_19436);
nor UO_1794 (O_1794,N_18130,N_19133);
nor UO_1795 (O_1795,N_19400,N_18831);
nor UO_1796 (O_1796,N_19450,N_18946);
xor UO_1797 (O_1797,N_18606,N_19755);
xnor UO_1798 (O_1798,N_19376,N_18763);
and UO_1799 (O_1799,N_19362,N_19292);
xnor UO_1800 (O_1800,N_19267,N_19167);
or UO_1801 (O_1801,N_19194,N_18142);
nand UO_1802 (O_1802,N_18567,N_19749);
nor UO_1803 (O_1803,N_18707,N_19992);
and UO_1804 (O_1804,N_19404,N_18490);
and UO_1805 (O_1805,N_19632,N_19788);
or UO_1806 (O_1806,N_18675,N_19612);
nand UO_1807 (O_1807,N_19375,N_18840);
xnor UO_1808 (O_1808,N_19145,N_19403);
nor UO_1809 (O_1809,N_18822,N_18664);
and UO_1810 (O_1810,N_18668,N_18710);
or UO_1811 (O_1811,N_18064,N_19287);
nor UO_1812 (O_1812,N_19795,N_18065);
and UO_1813 (O_1813,N_18029,N_18597);
and UO_1814 (O_1814,N_19134,N_19077);
nor UO_1815 (O_1815,N_19415,N_19649);
and UO_1816 (O_1816,N_18978,N_18857);
or UO_1817 (O_1817,N_19660,N_18356);
or UO_1818 (O_1818,N_18605,N_19817);
nand UO_1819 (O_1819,N_19768,N_19812);
and UO_1820 (O_1820,N_19103,N_19525);
and UO_1821 (O_1821,N_19944,N_19690);
nand UO_1822 (O_1822,N_18867,N_19766);
or UO_1823 (O_1823,N_19630,N_19326);
nor UO_1824 (O_1824,N_19889,N_18638);
or UO_1825 (O_1825,N_18899,N_19276);
nand UO_1826 (O_1826,N_18126,N_18053);
or UO_1827 (O_1827,N_19831,N_19094);
or UO_1828 (O_1828,N_18461,N_18304);
or UO_1829 (O_1829,N_19955,N_19930);
nand UO_1830 (O_1830,N_18423,N_18691);
nand UO_1831 (O_1831,N_19423,N_18542);
nor UO_1832 (O_1832,N_18798,N_18215);
xor UO_1833 (O_1833,N_19076,N_18335);
nand UO_1834 (O_1834,N_19663,N_18536);
xor UO_1835 (O_1835,N_18933,N_19071);
and UO_1836 (O_1836,N_18158,N_19906);
nor UO_1837 (O_1837,N_18436,N_19279);
and UO_1838 (O_1838,N_18965,N_19446);
nand UO_1839 (O_1839,N_18940,N_18985);
and UO_1840 (O_1840,N_18664,N_18295);
and UO_1841 (O_1841,N_18828,N_18432);
nor UO_1842 (O_1842,N_19775,N_19037);
or UO_1843 (O_1843,N_19220,N_18765);
nand UO_1844 (O_1844,N_19725,N_18914);
and UO_1845 (O_1845,N_18992,N_19887);
xor UO_1846 (O_1846,N_19794,N_18885);
and UO_1847 (O_1847,N_19272,N_18795);
nor UO_1848 (O_1848,N_18142,N_18772);
xor UO_1849 (O_1849,N_18051,N_19418);
nand UO_1850 (O_1850,N_18540,N_18553);
or UO_1851 (O_1851,N_18511,N_19655);
nand UO_1852 (O_1852,N_18470,N_18208);
or UO_1853 (O_1853,N_19059,N_19701);
nand UO_1854 (O_1854,N_18099,N_19310);
xor UO_1855 (O_1855,N_19589,N_18314);
nand UO_1856 (O_1856,N_19727,N_18342);
nand UO_1857 (O_1857,N_19707,N_19408);
nor UO_1858 (O_1858,N_19604,N_18284);
or UO_1859 (O_1859,N_19044,N_18341);
and UO_1860 (O_1860,N_18740,N_19249);
xor UO_1861 (O_1861,N_19143,N_18144);
nand UO_1862 (O_1862,N_18501,N_19534);
and UO_1863 (O_1863,N_19851,N_18448);
nand UO_1864 (O_1864,N_18424,N_19884);
xnor UO_1865 (O_1865,N_18811,N_18923);
or UO_1866 (O_1866,N_19624,N_18711);
or UO_1867 (O_1867,N_18355,N_19770);
nor UO_1868 (O_1868,N_18837,N_18694);
nand UO_1869 (O_1869,N_18395,N_19471);
nand UO_1870 (O_1870,N_18771,N_18902);
xor UO_1871 (O_1871,N_19885,N_18369);
and UO_1872 (O_1872,N_19522,N_18501);
xor UO_1873 (O_1873,N_19576,N_18815);
and UO_1874 (O_1874,N_18842,N_18368);
xor UO_1875 (O_1875,N_18464,N_18890);
nand UO_1876 (O_1876,N_19928,N_18274);
xnor UO_1877 (O_1877,N_18069,N_18965);
xor UO_1878 (O_1878,N_18802,N_18501);
xor UO_1879 (O_1879,N_19597,N_18692);
or UO_1880 (O_1880,N_18264,N_18483);
and UO_1881 (O_1881,N_19103,N_18311);
xnor UO_1882 (O_1882,N_19344,N_18423);
and UO_1883 (O_1883,N_18416,N_18902);
xor UO_1884 (O_1884,N_18116,N_18331);
nand UO_1885 (O_1885,N_19855,N_19929);
xnor UO_1886 (O_1886,N_18758,N_18944);
nand UO_1887 (O_1887,N_19280,N_18374);
nand UO_1888 (O_1888,N_19766,N_18266);
and UO_1889 (O_1889,N_19237,N_19599);
nand UO_1890 (O_1890,N_18847,N_18497);
xnor UO_1891 (O_1891,N_18839,N_19287);
nand UO_1892 (O_1892,N_18928,N_19282);
nor UO_1893 (O_1893,N_19494,N_19780);
nand UO_1894 (O_1894,N_19009,N_18515);
or UO_1895 (O_1895,N_19372,N_18826);
nor UO_1896 (O_1896,N_18439,N_19381);
xnor UO_1897 (O_1897,N_18219,N_18633);
or UO_1898 (O_1898,N_18377,N_18111);
nor UO_1899 (O_1899,N_18935,N_18892);
or UO_1900 (O_1900,N_18174,N_19076);
nand UO_1901 (O_1901,N_18609,N_18785);
xnor UO_1902 (O_1902,N_18958,N_19673);
and UO_1903 (O_1903,N_19508,N_19541);
nor UO_1904 (O_1904,N_19929,N_18852);
xor UO_1905 (O_1905,N_19532,N_18657);
or UO_1906 (O_1906,N_19579,N_18460);
nor UO_1907 (O_1907,N_19764,N_19384);
nand UO_1908 (O_1908,N_18026,N_18726);
nand UO_1909 (O_1909,N_19084,N_18602);
or UO_1910 (O_1910,N_18465,N_19795);
nand UO_1911 (O_1911,N_18896,N_18670);
and UO_1912 (O_1912,N_18120,N_18353);
or UO_1913 (O_1913,N_19119,N_19958);
nor UO_1914 (O_1914,N_19747,N_18623);
nand UO_1915 (O_1915,N_18635,N_18685);
and UO_1916 (O_1916,N_18494,N_19947);
nand UO_1917 (O_1917,N_19737,N_19684);
or UO_1918 (O_1918,N_18354,N_18719);
nor UO_1919 (O_1919,N_19705,N_19735);
nand UO_1920 (O_1920,N_18008,N_18930);
and UO_1921 (O_1921,N_19843,N_18915);
xor UO_1922 (O_1922,N_19518,N_19002);
nand UO_1923 (O_1923,N_19306,N_18448);
or UO_1924 (O_1924,N_19727,N_18223);
nor UO_1925 (O_1925,N_18692,N_19998);
nand UO_1926 (O_1926,N_19254,N_18601);
nor UO_1927 (O_1927,N_18286,N_18345);
and UO_1928 (O_1928,N_18229,N_18702);
nand UO_1929 (O_1929,N_18120,N_18249);
xnor UO_1930 (O_1930,N_18766,N_19987);
nand UO_1931 (O_1931,N_19158,N_18221);
and UO_1932 (O_1932,N_18378,N_18375);
or UO_1933 (O_1933,N_18858,N_18054);
or UO_1934 (O_1934,N_19128,N_19932);
nor UO_1935 (O_1935,N_19471,N_18242);
or UO_1936 (O_1936,N_18944,N_18038);
or UO_1937 (O_1937,N_18966,N_18958);
or UO_1938 (O_1938,N_19431,N_18716);
and UO_1939 (O_1939,N_19800,N_19382);
xor UO_1940 (O_1940,N_19642,N_18415);
xnor UO_1941 (O_1941,N_18877,N_19184);
nor UO_1942 (O_1942,N_18407,N_19490);
nand UO_1943 (O_1943,N_18479,N_19547);
nor UO_1944 (O_1944,N_19267,N_19593);
nor UO_1945 (O_1945,N_19014,N_19703);
nor UO_1946 (O_1946,N_18923,N_18703);
or UO_1947 (O_1947,N_18568,N_18792);
xnor UO_1948 (O_1948,N_19764,N_18597);
nor UO_1949 (O_1949,N_19925,N_19093);
xor UO_1950 (O_1950,N_19647,N_18237);
nor UO_1951 (O_1951,N_18825,N_19286);
nand UO_1952 (O_1952,N_18228,N_19627);
xor UO_1953 (O_1953,N_18837,N_18898);
xnor UO_1954 (O_1954,N_18813,N_19239);
nand UO_1955 (O_1955,N_19207,N_18409);
and UO_1956 (O_1956,N_18143,N_19073);
nand UO_1957 (O_1957,N_19294,N_19644);
and UO_1958 (O_1958,N_19376,N_19227);
or UO_1959 (O_1959,N_19367,N_18109);
and UO_1960 (O_1960,N_18003,N_18186);
nand UO_1961 (O_1961,N_19369,N_19590);
nor UO_1962 (O_1962,N_19254,N_19265);
or UO_1963 (O_1963,N_19670,N_19701);
nand UO_1964 (O_1964,N_18124,N_19108);
or UO_1965 (O_1965,N_19666,N_19967);
nand UO_1966 (O_1966,N_19470,N_19563);
nand UO_1967 (O_1967,N_19490,N_19687);
nand UO_1968 (O_1968,N_18584,N_19674);
xor UO_1969 (O_1969,N_18507,N_18550);
or UO_1970 (O_1970,N_18621,N_19499);
nor UO_1971 (O_1971,N_18780,N_19592);
nor UO_1972 (O_1972,N_18725,N_19754);
nor UO_1973 (O_1973,N_19448,N_19325);
nor UO_1974 (O_1974,N_18457,N_18020);
nor UO_1975 (O_1975,N_19457,N_18711);
and UO_1976 (O_1976,N_18968,N_18276);
xnor UO_1977 (O_1977,N_19127,N_19969);
nand UO_1978 (O_1978,N_19733,N_18903);
or UO_1979 (O_1979,N_18859,N_19888);
or UO_1980 (O_1980,N_18775,N_19120);
and UO_1981 (O_1981,N_19469,N_19896);
or UO_1982 (O_1982,N_18294,N_19946);
or UO_1983 (O_1983,N_18075,N_19159);
xnor UO_1984 (O_1984,N_19231,N_19541);
nor UO_1985 (O_1985,N_18617,N_18686);
or UO_1986 (O_1986,N_19521,N_19740);
or UO_1987 (O_1987,N_18171,N_18391);
xnor UO_1988 (O_1988,N_18552,N_18510);
xor UO_1989 (O_1989,N_18077,N_18442);
or UO_1990 (O_1990,N_19589,N_18400);
nor UO_1991 (O_1991,N_19336,N_18907);
and UO_1992 (O_1992,N_19517,N_18850);
and UO_1993 (O_1993,N_19975,N_19356);
nand UO_1994 (O_1994,N_18588,N_18073);
and UO_1995 (O_1995,N_19770,N_18629);
nor UO_1996 (O_1996,N_18711,N_19515);
xnor UO_1997 (O_1997,N_18187,N_18680);
and UO_1998 (O_1998,N_19667,N_19518);
nor UO_1999 (O_1999,N_18356,N_18752);
nor UO_2000 (O_2000,N_18728,N_18417);
or UO_2001 (O_2001,N_19861,N_18301);
xnor UO_2002 (O_2002,N_18832,N_18703);
xnor UO_2003 (O_2003,N_19033,N_18661);
xor UO_2004 (O_2004,N_19765,N_18058);
nand UO_2005 (O_2005,N_18534,N_19394);
nand UO_2006 (O_2006,N_19046,N_18224);
nor UO_2007 (O_2007,N_18357,N_18754);
nand UO_2008 (O_2008,N_18811,N_19358);
or UO_2009 (O_2009,N_18122,N_18026);
nand UO_2010 (O_2010,N_18166,N_19955);
nand UO_2011 (O_2011,N_19341,N_18272);
xnor UO_2012 (O_2012,N_18974,N_18862);
or UO_2013 (O_2013,N_18823,N_18070);
xor UO_2014 (O_2014,N_18289,N_19009);
xor UO_2015 (O_2015,N_19357,N_18562);
or UO_2016 (O_2016,N_18452,N_19928);
xnor UO_2017 (O_2017,N_18040,N_18843);
nand UO_2018 (O_2018,N_19738,N_18513);
xor UO_2019 (O_2019,N_18532,N_19021);
and UO_2020 (O_2020,N_19946,N_19633);
and UO_2021 (O_2021,N_18469,N_18522);
nor UO_2022 (O_2022,N_18543,N_18328);
and UO_2023 (O_2023,N_18289,N_18017);
xor UO_2024 (O_2024,N_19742,N_18530);
and UO_2025 (O_2025,N_18134,N_18353);
or UO_2026 (O_2026,N_19154,N_18757);
or UO_2027 (O_2027,N_19199,N_19566);
nand UO_2028 (O_2028,N_19059,N_19750);
nand UO_2029 (O_2029,N_18258,N_18981);
nand UO_2030 (O_2030,N_18646,N_18246);
and UO_2031 (O_2031,N_19708,N_19018);
nor UO_2032 (O_2032,N_19706,N_19798);
nor UO_2033 (O_2033,N_19783,N_18763);
nand UO_2034 (O_2034,N_19364,N_19200);
nand UO_2035 (O_2035,N_19520,N_18818);
xor UO_2036 (O_2036,N_18861,N_19677);
or UO_2037 (O_2037,N_18954,N_19706);
nor UO_2038 (O_2038,N_18436,N_18491);
and UO_2039 (O_2039,N_18855,N_18287);
or UO_2040 (O_2040,N_18908,N_19471);
and UO_2041 (O_2041,N_18479,N_19899);
nand UO_2042 (O_2042,N_18988,N_19479);
nand UO_2043 (O_2043,N_18156,N_19829);
nor UO_2044 (O_2044,N_18397,N_18667);
and UO_2045 (O_2045,N_18112,N_19491);
xor UO_2046 (O_2046,N_18495,N_18830);
or UO_2047 (O_2047,N_19924,N_18218);
and UO_2048 (O_2048,N_19980,N_19905);
nor UO_2049 (O_2049,N_18721,N_18879);
nor UO_2050 (O_2050,N_18042,N_19249);
nor UO_2051 (O_2051,N_18112,N_18199);
nor UO_2052 (O_2052,N_18653,N_19663);
and UO_2053 (O_2053,N_19835,N_19387);
nor UO_2054 (O_2054,N_18634,N_19296);
or UO_2055 (O_2055,N_18462,N_19738);
xor UO_2056 (O_2056,N_19897,N_18057);
xor UO_2057 (O_2057,N_19221,N_18339);
xor UO_2058 (O_2058,N_19343,N_19097);
nor UO_2059 (O_2059,N_19497,N_18657);
and UO_2060 (O_2060,N_19299,N_19501);
nand UO_2061 (O_2061,N_19086,N_18162);
xor UO_2062 (O_2062,N_19868,N_18259);
and UO_2063 (O_2063,N_19784,N_18983);
and UO_2064 (O_2064,N_18241,N_18774);
or UO_2065 (O_2065,N_18328,N_18332);
xor UO_2066 (O_2066,N_19258,N_19545);
xnor UO_2067 (O_2067,N_19415,N_19664);
nand UO_2068 (O_2068,N_19145,N_19727);
nand UO_2069 (O_2069,N_19703,N_18905);
nand UO_2070 (O_2070,N_19656,N_18417);
and UO_2071 (O_2071,N_19989,N_18866);
nor UO_2072 (O_2072,N_19020,N_19664);
xor UO_2073 (O_2073,N_19578,N_19501);
and UO_2074 (O_2074,N_18595,N_18076);
xnor UO_2075 (O_2075,N_19880,N_18561);
xnor UO_2076 (O_2076,N_19942,N_18702);
xnor UO_2077 (O_2077,N_19946,N_18844);
or UO_2078 (O_2078,N_18126,N_19946);
xor UO_2079 (O_2079,N_19165,N_19592);
nor UO_2080 (O_2080,N_19226,N_18284);
or UO_2081 (O_2081,N_18400,N_18577);
and UO_2082 (O_2082,N_18496,N_19359);
and UO_2083 (O_2083,N_18122,N_18142);
or UO_2084 (O_2084,N_18221,N_18591);
nand UO_2085 (O_2085,N_18618,N_19851);
or UO_2086 (O_2086,N_18335,N_19270);
or UO_2087 (O_2087,N_19339,N_19429);
nor UO_2088 (O_2088,N_19676,N_18332);
nand UO_2089 (O_2089,N_18013,N_18468);
or UO_2090 (O_2090,N_18845,N_18648);
and UO_2091 (O_2091,N_19617,N_19993);
xor UO_2092 (O_2092,N_18110,N_18569);
xor UO_2093 (O_2093,N_19243,N_19332);
xor UO_2094 (O_2094,N_19848,N_19998);
and UO_2095 (O_2095,N_18262,N_19120);
and UO_2096 (O_2096,N_19964,N_19723);
or UO_2097 (O_2097,N_18271,N_19747);
nor UO_2098 (O_2098,N_18944,N_18747);
or UO_2099 (O_2099,N_19996,N_19640);
nand UO_2100 (O_2100,N_19797,N_18447);
nand UO_2101 (O_2101,N_19398,N_19280);
xnor UO_2102 (O_2102,N_18728,N_18213);
nor UO_2103 (O_2103,N_19069,N_18411);
or UO_2104 (O_2104,N_19372,N_19506);
and UO_2105 (O_2105,N_19518,N_18461);
nor UO_2106 (O_2106,N_19760,N_18059);
xor UO_2107 (O_2107,N_19957,N_19175);
or UO_2108 (O_2108,N_19060,N_19377);
or UO_2109 (O_2109,N_18786,N_18855);
xnor UO_2110 (O_2110,N_18380,N_19211);
nor UO_2111 (O_2111,N_19585,N_18360);
nand UO_2112 (O_2112,N_19832,N_18935);
or UO_2113 (O_2113,N_18551,N_18703);
xnor UO_2114 (O_2114,N_19638,N_18631);
xor UO_2115 (O_2115,N_19787,N_19652);
nand UO_2116 (O_2116,N_19521,N_19273);
and UO_2117 (O_2117,N_18661,N_19524);
nor UO_2118 (O_2118,N_19138,N_18849);
nand UO_2119 (O_2119,N_18502,N_19775);
xnor UO_2120 (O_2120,N_19099,N_18771);
and UO_2121 (O_2121,N_19740,N_18352);
and UO_2122 (O_2122,N_18956,N_18430);
xnor UO_2123 (O_2123,N_19928,N_19579);
or UO_2124 (O_2124,N_18131,N_19182);
or UO_2125 (O_2125,N_19933,N_19910);
xor UO_2126 (O_2126,N_19975,N_18937);
or UO_2127 (O_2127,N_19435,N_18278);
xor UO_2128 (O_2128,N_19489,N_19303);
xnor UO_2129 (O_2129,N_19532,N_18295);
or UO_2130 (O_2130,N_18773,N_19765);
xnor UO_2131 (O_2131,N_18291,N_19752);
xnor UO_2132 (O_2132,N_19077,N_18029);
xor UO_2133 (O_2133,N_19984,N_19436);
or UO_2134 (O_2134,N_19662,N_18129);
or UO_2135 (O_2135,N_18026,N_18737);
or UO_2136 (O_2136,N_19439,N_19196);
or UO_2137 (O_2137,N_19323,N_19342);
and UO_2138 (O_2138,N_18764,N_19860);
nor UO_2139 (O_2139,N_19907,N_18431);
nor UO_2140 (O_2140,N_18295,N_18556);
nor UO_2141 (O_2141,N_18245,N_18080);
nand UO_2142 (O_2142,N_19785,N_19493);
and UO_2143 (O_2143,N_18736,N_18709);
nor UO_2144 (O_2144,N_19247,N_19063);
nor UO_2145 (O_2145,N_18346,N_19331);
or UO_2146 (O_2146,N_18073,N_19547);
or UO_2147 (O_2147,N_19756,N_18612);
xor UO_2148 (O_2148,N_19244,N_18601);
nor UO_2149 (O_2149,N_19245,N_19502);
and UO_2150 (O_2150,N_18518,N_19299);
nor UO_2151 (O_2151,N_19027,N_19900);
and UO_2152 (O_2152,N_18845,N_19033);
xor UO_2153 (O_2153,N_18399,N_19810);
nand UO_2154 (O_2154,N_18072,N_19453);
and UO_2155 (O_2155,N_18188,N_18454);
xnor UO_2156 (O_2156,N_18974,N_18210);
and UO_2157 (O_2157,N_19067,N_19763);
nor UO_2158 (O_2158,N_18818,N_18925);
or UO_2159 (O_2159,N_19327,N_18627);
nor UO_2160 (O_2160,N_19963,N_19588);
and UO_2161 (O_2161,N_19824,N_19607);
xnor UO_2162 (O_2162,N_19233,N_18372);
nor UO_2163 (O_2163,N_18442,N_18520);
or UO_2164 (O_2164,N_19622,N_18690);
xnor UO_2165 (O_2165,N_19526,N_18597);
nor UO_2166 (O_2166,N_18236,N_18530);
nand UO_2167 (O_2167,N_19078,N_18441);
or UO_2168 (O_2168,N_18986,N_18273);
nor UO_2169 (O_2169,N_19820,N_19946);
xor UO_2170 (O_2170,N_18065,N_19611);
nand UO_2171 (O_2171,N_18957,N_19429);
nand UO_2172 (O_2172,N_18707,N_19079);
nand UO_2173 (O_2173,N_18145,N_18407);
xor UO_2174 (O_2174,N_19742,N_19345);
nand UO_2175 (O_2175,N_19565,N_19717);
and UO_2176 (O_2176,N_18724,N_19799);
nand UO_2177 (O_2177,N_18436,N_18753);
nand UO_2178 (O_2178,N_19880,N_18662);
nand UO_2179 (O_2179,N_19358,N_18442);
or UO_2180 (O_2180,N_18407,N_18413);
and UO_2181 (O_2181,N_18765,N_19261);
or UO_2182 (O_2182,N_19952,N_19353);
xor UO_2183 (O_2183,N_18600,N_18215);
nand UO_2184 (O_2184,N_18586,N_19196);
nor UO_2185 (O_2185,N_18762,N_18211);
or UO_2186 (O_2186,N_18258,N_18900);
and UO_2187 (O_2187,N_18762,N_18822);
and UO_2188 (O_2188,N_19347,N_18992);
xor UO_2189 (O_2189,N_19486,N_18946);
nor UO_2190 (O_2190,N_19815,N_19852);
xor UO_2191 (O_2191,N_19772,N_18806);
or UO_2192 (O_2192,N_19682,N_19114);
nor UO_2193 (O_2193,N_19953,N_19747);
nor UO_2194 (O_2194,N_19818,N_19217);
or UO_2195 (O_2195,N_19217,N_18854);
and UO_2196 (O_2196,N_19414,N_18546);
xnor UO_2197 (O_2197,N_18656,N_18654);
nand UO_2198 (O_2198,N_19635,N_19814);
nand UO_2199 (O_2199,N_19574,N_18793);
or UO_2200 (O_2200,N_19938,N_18166);
nor UO_2201 (O_2201,N_18860,N_18341);
nand UO_2202 (O_2202,N_19860,N_19545);
xor UO_2203 (O_2203,N_18006,N_18444);
nand UO_2204 (O_2204,N_18270,N_19918);
nand UO_2205 (O_2205,N_18774,N_18721);
nand UO_2206 (O_2206,N_18371,N_19897);
nand UO_2207 (O_2207,N_18254,N_18746);
xnor UO_2208 (O_2208,N_18542,N_19389);
nand UO_2209 (O_2209,N_19106,N_19388);
nand UO_2210 (O_2210,N_19973,N_18383);
xnor UO_2211 (O_2211,N_19757,N_18989);
nor UO_2212 (O_2212,N_19783,N_19787);
nand UO_2213 (O_2213,N_19821,N_18236);
and UO_2214 (O_2214,N_18273,N_18486);
nand UO_2215 (O_2215,N_18030,N_19074);
xor UO_2216 (O_2216,N_19064,N_19896);
or UO_2217 (O_2217,N_18768,N_18813);
and UO_2218 (O_2218,N_19252,N_18418);
xnor UO_2219 (O_2219,N_19477,N_19211);
or UO_2220 (O_2220,N_19770,N_18165);
or UO_2221 (O_2221,N_19516,N_19021);
nor UO_2222 (O_2222,N_18865,N_18154);
xnor UO_2223 (O_2223,N_19172,N_19672);
xor UO_2224 (O_2224,N_18497,N_18239);
xnor UO_2225 (O_2225,N_19589,N_19748);
nand UO_2226 (O_2226,N_18686,N_18938);
and UO_2227 (O_2227,N_18001,N_18395);
and UO_2228 (O_2228,N_19393,N_18606);
nor UO_2229 (O_2229,N_19831,N_19660);
xnor UO_2230 (O_2230,N_18484,N_19573);
nand UO_2231 (O_2231,N_19214,N_18878);
nor UO_2232 (O_2232,N_18170,N_18964);
nand UO_2233 (O_2233,N_18194,N_19102);
xnor UO_2234 (O_2234,N_19537,N_19146);
nor UO_2235 (O_2235,N_18964,N_18019);
and UO_2236 (O_2236,N_19657,N_19624);
and UO_2237 (O_2237,N_18292,N_18520);
and UO_2238 (O_2238,N_18884,N_19199);
and UO_2239 (O_2239,N_19241,N_18657);
nor UO_2240 (O_2240,N_18988,N_19897);
xor UO_2241 (O_2241,N_18907,N_19177);
nor UO_2242 (O_2242,N_18941,N_18571);
nor UO_2243 (O_2243,N_19587,N_18548);
or UO_2244 (O_2244,N_19047,N_18760);
and UO_2245 (O_2245,N_18000,N_18500);
xor UO_2246 (O_2246,N_18226,N_18523);
or UO_2247 (O_2247,N_18368,N_18616);
nor UO_2248 (O_2248,N_19257,N_19084);
xnor UO_2249 (O_2249,N_19528,N_18728);
nor UO_2250 (O_2250,N_19936,N_18510);
nand UO_2251 (O_2251,N_18956,N_19630);
or UO_2252 (O_2252,N_18024,N_18585);
xor UO_2253 (O_2253,N_19133,N_19974);
nand UO_2254 (O_2254,N_19309,N_19708);
xor UO_2255 (O_2255,N_19503,N_19258);
nor UO_2256 (O_2256,N_18344,N_19151);
and UO_2257 (O_2257,N_19488,N_19940);
nand UO_2258 (O_2258,N_18435,N_19998);
or UO_2259 (O_2259,N_18079,N_19626);
nor UO_2260 (O_2260,N_18916,N_19706);
or UO_2261 (O_2261,N_19555,N_18215);
nor UO_2262 (O_2262,N_18142,N_19922);
or UO_2263 (O_2263,N_18806,N_19296);
nand UO_2264 (O_2264,N_18530,N_18910);
nand UO_2265 (O_2265,N_19603,N_18675);
nand UO_2266 (O_2266,N_19653,N_18038);
or UO_2267 (O_2267,N_18684,N_19666);
nand UO_2268 (O_2268,N_19766,N_19432);
or UO_2269 (O_2269,N_19892,N_18802);
or UO_2270 (O_2270,N_18285,N_18511);
and UO_2271 (O_2271,N_19537,N_19549);
and UO_2272 (O_2272,N_19937,N_19354);
or UO_2273 (O_2273,N_18022,N_19699);
and UO_2274 (O_2274,N_19462,N_19798);
nor UO_2275 (O_2275,N_18913,N_18135);
xnor UO_2276 (O_2276,N_19486,N_19566);
nand UO_2277 (O_2277,N_19007,N_18484);
and UO_2278 (O_2278,N_18206,N_18032);
and UO_2279 (O_2279,N_19433,N_19415);
nand UO_2280 (O_2280,N_19730,N_18376);
nor UO_2281 (O_2281,N_18865,N_19113);
nor UO_2282 (O_2282,N_19696,N_19411);
xor UO_2283 (O_2283,N_19339,N_18264);
nand UO_2284 (O_2284,N_19733,N_19344);
nand UO_2285 (O_2285,N_19044,N_18297);
or UO_2286 (O_2286,N_18987,N_18924);
nor UO_2287 (O_2287,N_19132,N_19432);
xnor UO_2288 (O_2288,N_18223,N_19526);
nand UO_2289 (O_2289,N_19356,N_18133);
nand UO_2290 (O_2290,N_18474,N_19448);
or UO_2291 (O_2291,N_18936,N_18853);
and UO_2292 (O_2292,N_19618,N_19356);
nand UO_2293 (O_2293,N_19148,N_18665);
nor UO_2294 (O_2294,N_19047,N_19315);
and UO_2295 (O_2295,N_19484,N_19446);
or UO_2296 (O_2296,N_19630,N_19034);
or UO_2297 (O_2297,N_18274,N_19343);
nor UO_2298 (O_2298,N_19374,N_19090);
xnor UO_2299 (O_2299,N_19632,N_18314);
and UO_2300 (O_2300,N_18881,N_19067);
nand UO_2301 (O_2301,N_18955,N_18470);
nor UO_2302 (O_2302,N_19158,N_18272);
xor UO_2303 (O_2303,N_19779,N_18360);
or UO_2304 (O_2304,N_18333,N_18431);
or UO_2305 (O_2305,N_18115,N_19858);
nand UO_2306 (O_2306,N_19428,N_18440);
or UO_2307 (O_2307,N_19115,N_19898);
nand UO_2308 (O_2308,N_18148,N_18334);
and UO_2309 (O_2309,N_19194,N_19292);
nor UO_2310 (O_2310,N_18028,N_19892);
nor UO_2311 (O_2311,N_19285,N_18352);
xor UO_2312 (O_2312,N_18921,N_18200);
or UO_2313 (O_2313,N_18973,N_18053);
xor UO_2314 (O_2314,N_18448,N_18217);
xnor UO_2315 (O_2315,N_18492,N_18465);
xor UO_2316 (O_2316,N_19605,N_18397);
xnor UO_2317 (O_2317,N_19884,N_19359);
nor UO_2318 (O_2318,N_18634,N_18829);
nor UO_2319 (O_2319,N_19670,N_18362);
xnor UO_2320 (O_2320,N_18206,N_18763);
or UO_2321 (O_2321,N_18953,N_19066);
nand UO_2322 (O_2322,N_18641,N_18272);
and UO_2323 (O_2323,N_18350,N_18603);
and UO_2324 (O_2324,N_18961,N_19200);
nor UO_2325 (O_2325,N_18072,N_19211);
xnor UO_2326 (O_2326,N_19779,N_19079);
or UO_2327 (O_2327,N_19536,N_18637);
or UO_2328 (O_2328,N_19801,N_19137);
nor UO_2329 (O_2329,N_19637,N_19403);
nand UO_2330 (O_2330,N_18065,N_18749);
nand UO_2331 (O_2331,N_18617,N_19980);
or UO_2332 (O_2332,N_18919,N_19763);
and UO_2333 (O_2333,N_18669,N_18056);
and UO_2334 (O_2334,N_18307,N_19954);
xnor UO_2335 (O_2335,N_19375,N_18416);
and UO_2336 (O_2336,N_19217,N_18663);
xnor UO_2337 (O_2337,N_19437,N_18063);
xor UO_2338 (O_2338,N_18235,N_18941);
nand UO_2339 (O_2339,N_18350,N_19492);
xnor UO_2340 (O_2340,N_19283,N_19070);
nor UO_2341 (O_2341,N_18734,N_19144);
nor UO_2342 (O_2342,N_18438,N_18853);
nor UO_2343 (O_2343,N_18437,N_18538);
and UO_2344 (O_2344,N_18955,N_18221);
nor UO_2345 (O_2345,N_18830,N_18537);
nand UO_2346 (O_2346,N_18600,N_18959);
nor UO_2347 (O_2347,N_19373,N_18096);
or UO_2348 (O_2348,N_19186,N_18512);
or UO_2349 (O_2349,N_18726,N_18982);
and UO_2350 (O_2350,N_19561,N_19983);
nor UO_2351 (O_2351,N_18931,N_18858);
nand UO_2352 (O_2352,N_19208,N_19108);
nor UO_2353 (O_2353,N_19691,N_19584);
or UO_2354 (O_2354,N_19060,N_18569);
or UO_2355 (O_2355,N_19964,N_18302);
or UO_2356 (O_2356,N_18947,N_18957);
xnor UO_2357 (O_2357,N_18521,N_18715);
nor UO_2358 (O_2358,N_18278,N_18354);
nor UO_2359 (O_2359,N_19789,N_18803);
or UO_2360 (O_2360,N_19233,N_18127);
nand UO_2361 (O_2361,N_18957,N_18756);
nand UO_2362 (O_2362,N_18124,N_18384);
nand UO_2363 (O_2363,N_18938,N_18918);
and UO_2364 (O_2364,N_19694,N_18779);
and UO_2365 (O_2365,N_18942,N_19702);
nor UO_2366 (O_2366,N_19860,N_19020);
or UO_2367 (O_2367,N_19727,N_18017);
or UO_2368 (O_2368,N_19985,N_19044);
xor UO_2369 (O_2369,N_19888,N_18078);
nand UO_2370 (O_2370,N_19196,N_19139);
or UO_2371 (O_2371,N_19192,N_19091);
nand UO_2372 (O_2372,N_18125,N_19518);
xor UO_2373 (O_2373,N_19992,N_18758);
nand UO_2374 (O_2374,N_18423,N_19921);
nand UO_2375 (O_2375,N_18749,N_19659);
and UO_2376 (O_2376,N_19298,N_19019);
xor UO_2377 (O_2377,N_18740,N_19630);
xor UO_2378 (O_2378,N_19181,N_19236);
and UO_2379 (O_2379,N_18003,N_19321);
xnor UO_2380 (O_2380,N_18909,N_18195);
nor UO_2381 (O_2381,N_18580,N_19017);
xnor UO_2382 (O_2382,N_19412,N_18924);
nor UO_2383 (O_2383,N_19808,N_18122);
and UO_2384 (O_2384,N_18029,N_19061);
nor UO_2385 (O_2385,N_19985,N_18861);
xnor UO_2386 (O_2386,N_19370,N_19021);
or UO_2387 (O_2387,N_18139,N_18607);
and UO_2388 (O_2388,N_19042,N_18413);
nand UO_2389 (O_2389,N_18257,N_19184);
xor UO_2390 (O_2390,N_18425,N_19146);
and UO_2391 (O_2391,N_18421,N_19388);
nor UO_2392 (O_2392,N_19321,N_19167);
xnor UO_2393 (O_2393,N_19501,N_18733);
and UO_2394 (O_2394,N_19873,N_19296);
nor UO_2395 (O_2395,N_18575,N_18185);
nor UO_2396 (O_2396,N_19291,N_18372);
xor UO_2397 (O_2397,N_19193,N_18504);
xnor UO_2398 (O_2398,N_18846,N_19233);
xor UO_2399 (O_2399,N_18611,N_18014);
xnor UO_2400 (O_2400,N_18692,N_19634);
nor UO_2401 (O_2401,N_19592,N_19816);
xnor UO_2402 (O_2402,N_19222,N_19022);
nor UO_2403 (O_2403,N_18206,N_18402);
and UO_2404 (O_2404,N_19542,N_18344);
nor UO_2405 (O_2405,N_18880,N_19190);
nand UO_2406 (O_2406,N_18799,N_19306);
and UO_2407 (O_2407,N_19404,N_19862);
nor UO_2408 (O_2408,N_19000,N_18131);
and UO_2409 (O_2409,N_19523,N_18454);
xnor UO_2410 (O_2410,N_18902,N_18085);
xnor UO_2411 (O_2411,N_18109,N_19311);
nand UO_2412 (O_2412,N_18232,N_19344);
or UO_2413 (O_2413,N_19826,N_18036);
xnor UO_2414 (O_2414,N_18015,N_19399);
and UO_2415 (O_2415,N_19253,N_18112);
and UO_2416 (O_2416,N_18571,N_19365);
xnor UO_2417 (O_2417,N_18127,N_18490);
xor UO_2418 (O_2418,N_18117,N_19938);
nand UO_2419 (O_2419,N_18988,N_19873);
xor UO_2420 (O_2420,N_19234,N_19925);
or UO_2421 (O_2421,N_18043,N_19959);
nand UO_2422 (O_2422,N_18409,N_18534);
or UO_2423 (O_2423,N_19194,N_19057);
xor UO_2424 (O_2424,N_18776,N_18361);
nor UO_2425 (O_2425,N_18195,N_18827);
xnor UO_2426 (O_2426,N_19006,N_19553);
nor UO_2427 (O_2427,N_19116,N_19619);
or UO_2428 (O_2428,N_18906,N_18545);
xor UO_2429 (O_2429,N_18566,N_18391);
nor UO_2430 (O_2430,N_18028,N_19160);
or UO_2431 (O_2431,N_18655,N_18702);
or UO_2432 (O_2432,N_18696,N_18879);
nor UO_2433 (O_2433,N_19021,N_18671);
xnor UO_2434 (O_2434,N_19114,N_19742);
and UO_2435 (O_2435,N_19158,N_19071);
and UO_2436 (O_2436,N_19856,N_19004);
nor UO_2437 (O_2437,N_19012,N_19291);
nor UO_2438 (O_2438,N_19599,N_18969);
or UO_2439 (O_2439,N_19924,N_18484);
or UO_2440 (O_2440,N_19260,N_18473);
nand UO_2441 (O_2441,N_18628,N_18638);
nor UO_2442 (O_2442,N_18437,N_19557);
or UO_2443 (O_2443,N_19244,N_18623);
and UO_2444 (O_2444,N_18895,N_18023);
and UO_2445 (O_2445,N_19582,N_18275);
xnor UO_2446 (O_2446,N_19086,N_19514);
xnor UO_2447 (O_2447,N_18424,N_19595);
nand UO_2448 (O_2448,N_18428,N_18146);
xnor UO_2449 (O_2449,N_18662,N_18644);
nand UO_2450 (O_2450,N_19859,N_19784);
and UO_2451 (O_2451,N_18117,N_18907);
nand UO_2452 (O_2452,N_19694,N_19702);
xor UO_2453 (O_2453,N_19689,N_18007);
nor UO_2454 (O_2454,N_18123,N_18336);
or UO_2455 (O_2455,N_19390,N_18624);
and UO_2456 (O_2456,N_19308,N_19310);
nor UO_2457 (O_2457,N_18762,N_18011);
nor UO_2458 (O_2458,N_19536,N_18408);
and UO_2459 (O_2459,N_18808,N_18750);
or UO_2460 (O_2460,N_18820,N_19415);
nand UO_2461 (O_2461,N_18376,N_19896);
xor UO_2462 (O_2462,N_18609,N_19773);
nor UO_2463 (O_2463,N_19048,N_18390);
and UO_2464 (O_2464,N_18784,N_18227);
xnor UO_2465 (O_2465,N_19984,N_19452);
nor UO_2466 (O_2466,N_19235,N_19191);
xor UO_2467 (O_2467,N_19435,N_18848);
and UO_2468 (O_2468,N_18196,N_19913);
nand UO_2469 (O_2469,N_19334,N_18556);
and UO_2470 (O_2470,N_19847,N_18246);
or UO_2471 (O_2471,N_18407,N_18356);
or UO_2472 (O_2472,N_19677,N_18488);
xor UO_2473 (O_2473,N_18649,N_18669);
and UO_2474 (O_2474,N_18070,N_18454);
xnor UO_2475 (O_2475,N_19611,N_18443);
or UO_2476 (O_2476,N_19127,N_19699);
or UO_2477 (O_2477,N_18141,N_18515);
nor UO_2478 (O_2478,N_18021,N_18337);
nand UO_2479 (O_2479,N_18243,N_19160);
or UO_2480 (O_2480,N_19565,N_18184);
nand UO_2481 (O_2481,N_18863,N_18475);
xor UO_2482 (O_2482,N_18289,N_19163);
xnor UO_2483 (O_2483,N_19360,N_18383);
and UO_2484 (O_2484,N_19890,N_19918);
nand UO_2485 (O_2485,N_18824,N_19344);
xor UO_2486 (O_2486,N_19870,N_19875);
and UO_2487 (O_2487,N_18560,N_18163);
nor UO_2488 (O_2488,N_19875,N_18658);
nor UO_2489 (O_2489,N_19200,N_19411);
nor UO_2490 (O_2490,N_18009,N_18462);
or UO_2491 (O_2491,N_19414,N_18630);
nor UO_2492 (O_2492,N_19738,N_19314);
nand UO_2493 (O_2493,N_18903,N_18700);
xor UO_2494 (O_2494,N_19382,N_18323);
or UO_2495 (O_2495,N_19595,N_18269);
or UO_2496 (O_2496,N_19399,N_18366);
and UO_2497 (O_2497,N_19077,N_19959);
or UO_2498 (O_2498,N_19848,N_18808);
nor UO_2499 (O_2499,N_18628,N_18974);
endmodule