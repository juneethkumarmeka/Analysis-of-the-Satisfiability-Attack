module basic_3000_30000_3500_10_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_614,In_1413);
or U1 (N_1,In_2605,In_2535);
or U2 (N_2,In_1036,In_106);
nand U3 (N_3,In_498,In_475);
nand U4 (N_4,In_943,In_1772);
nand U5 (N_5,In_1118,In_505);
nor U6 (N_6,In_784,In_797);
or U7 (N_7,In_1606,In_2524);
and U8 (N_8,In_1326,In_892);
and U9 (N_9,In_834,In_802);
or U10 (N_10,In_1378,In_2270);
and U11 (N_11,In_180,In_664);
nor U12 (N_12,In_2982,In_2445);
and U13 (N_13,In_2267,In_2264);
or U14 (N_14,In_2861,In_405);
or U15 (N_15,In_1720,In_2858);
nand U16 (N_16,In_2285,In_1385);
nor U17 (N_17,In_953,In_1092);
xnor U18 (N_18,In_912,In_2555);
nand U19 (N_19,In_1062,In_358);
nand U20 (N_20,In_267,In_379);
nand U21 (N_21,In_2490,In_2308);
and U22 (N_22,In_1512,In_2795);
nand U23 (N_23,In_2780,In_2303);
nor U24 (N_24,In_1745,In_1623);
xnor U25 (N_25,In_1996,In_1047);
nand U26 (N_26,In_1121,In_2055);
and U27 (N_27,In_36,In_2251);
or U28 (N_28,In_1415,In_1132);
and U29 (N_29,In_924,In_1247);
xnor U30 (N_30,In_2794,In_2167);
and U31 (N_31,In_1104,In_454);
or U32 (N_32,In_1881,In_559);
and U33 (N_33,In_1513,In_2822);
and U34 (N_34,In_537,In_1811);
nor U35 (N_35,In_2968,In_1451);
nand U36 (N_36,In_2975,In_2126);
nor U37 (N_37,In_1009,In_277);
nand U38 (N_38,In_856,In_1454);
or U39 (N_39,In_2897,In_1787);
and U40 (N_40,In_826,In_112);
nor U41 (N_41,In_920,In_2621);
nand U42 (N_42,In_1626,In_2883);
xor U43 (N_43,In_1674,In_2284);
nor U44 (N_44,In_932,In_299);
nand U45 (N_45,In_1568,In_1327);
and U46 (N_46,In_890,In_2204);
and U47 (N_47,In_1497,In_2375);
nand U48 (N_48,In_2581,In_350);
nand U49 (N_49,In_796,In_2446);
nand U50 (N_50,In_2349,In_122);
xor U51 (N_51,In_2112,In_538);
or U52 (N_52,In_251,In_775);
and U53 (N_53,In_2325,In_1686);
nand U54 (N_54,In_2109,In_2095);
and U55 (N_55,In_1145,In_1109);
nand U56 (N_56,In_1916,In_396);
nor U57 (N_57,In_624,In_2225);
or U58 (N_58,In_2986,In_562);
or U59 (N_59,In_1929,In_148);
nor U60 (N_60,In_973,In_991);
nand U61 (N_61,In_957,In_2350);
nor U62 (N_62,In_1622,In_2715);
or U63 (N_63,In_1046,In_34);
nor U64 (N_64,In_962,In_1562);
nor U65 (N_65,In_2012,In_2667);
or U66 (N_66,In_2076,In_2448);
nand U67 (N_67,In_1695,In_1802);
nand U68 (N_68,In_2923,In_2471);
and U69 (N_69,In_1320,In_1670);
nand U70 (N_70,In_2031,In_2518);
or U71 (N_71,In_2027,In_1723);
nor U72 (N_72,In_2165,In_160);
and U73 (N_73,In_1691,In_476);
and U74 (N_74,In_1767,In_730);
nor U75 (N_75,In_52,In_770);
nor U76 (N_76,In_2341,In_1039);
nor U77 (N_77,In_104,In_1575);
nand U78 (N_78,In_404,In_1131);
nor U79 (N_79,In_2769,In_906);
nand U80 (N_80,In_2280,In_2599);
and U81 (N_81,In_780,In_1263);
nand U82 (N_82,In_1958,In_2281);
nor U83 (N_83,In_172,In_1441);
nor U84 (N_84,In_1532,In_1099);
and U85 (N_85,In_2036,In_1147);
or U86 (N_86,In_2944,In_368);
nand U87 (N_87,In_818,In_930);
nor U88 (N_88,In_2347,In_2082);
nand U89 (N_89,In_1064,In_196);
and U90 (N_90,In_1872,In_315);
nand U91 (N_91,In_2185,In_72);
xor U92 (N_92,In_1294,In_1467);
nor U93 (N_93,In_2260,In_841);
nand U94 (N_94,In_254,In_2606);
nand U95 (N_95,In_80,In_2531);
nor U96 (N_96,In_309,In_258);
and U97 (N_97,In_1564,In_1439);
nand U98 (N_98,In_1422,In_2917);
or U99 (N_99,In_2866,In_748);
or U100 (N_100,In_2345,In_846);
and U101 (N_101,In_2406,In_895);
xor U102 (N_102,In_313,In_1915);
nor U103 (N_103,In_734,In_400);
or U104 (N_104,In_2133,In_39);
and U105 (N_105,In_1485,In_1480);
and U106 (N_106,In_2101,In_185);
and U107 (N_107,In_206,In_1344);
nand U108 (N_108,In_1502,In_89);
nand U109 (N_109,In_2910,In_903);
or U110 (N_110,In_675,In_2005);
xor U111 (N_111,In_591,In_1017);
nand U112 (N_112,In_293,In_183);
nor U113 (N_113,In_433,In_2206);
nor U114 (N_114,In_2263,In_670);
xor U115 (N_115,In_1057,In_2559);
or U116 (N_116,In_1144,In_1035);
and U117 (N_117,In_356,In_577);
xor U118 (N_118,In_153,In_1424);
nand U119 (N_119,In_2111,In_2142);
nor U120 (N_120,In_1637,In_2679);
nand U121 (N_121,In_29,In_2814);
nor U122 (N_122,In_2368,In_1126);
and U123 (N_123,In_945,In_332);
nor U124 (N_124,In_2132,In_213);
nor U125 (N_125,In_1117,In_1844);
nand U126 (N_126,In_465,In_338);
nand U127 (N_127,In_2389,In_124);
and U128 (N_128,In_2416,In_955);
nand U129 (N_129,In_609,In_742);
nor U130 (N_130,In_417,In_1604);
xor U131 (N_131,In_2556,In_2949);
and U132 (N_132,In_1572,In_1177);
xor U133 (N_133,In_1919,In_919);
nor U134 (N_134,In_1506,In_2728);
or U135 (N_135,In_1054,In_2907);
nor U136 (N_136,In_1668,In_2993);
xor U137 (N_137,In_1137,In_851);
nor U138 (N_138,In_462,In_540);
nand U139 (N_139,In_193,In_515);
or U140 (N_140,In_640,In_2707);
xnor U141 (N_141,In_386,In_2618);
or U142 (N_142,In_888,In_2331);
and U143 (N_143,In_1114,In_1164);
and U144 (N_144,In_1168,In_1854);
and U145 (N_145,In_2105,In_992);
and U146 (N_146,In_922,In_779);
and U147 (N_147,In_1152,In_2598);
nor U148 (N_148,In_1636,In_2739);
or U149 (N_149,In_2764,In_2746);
nand U150 (N_150,In_1585,In_114);
nor U151 (N_151,In_178,In_123);
or U152 (N_152,In_1329,In_2181);
nor U153 (N_153,In_2979,In_2878);
and U154 (N_154,In_1793,In_416);
xor U155 (N_155,In_2772,In_1207);
nand U156 (N_156,In_1722,In_2753);
nand U157 (N_157,In_286,In_2880);
nor U158 (N_158,In_1433,In_1423);
nand U159 (N_159,In_2336,In_2919);
and U160 (N_160,In_1859,In_2918);
nor U161 (N_161,In_1914,In_990);
and U162 (N_162,In_2073,In_2030);
or U163 (N_163,In_1944,In_1019);
nor U164 (N_164,In_255,In_494);
and U165 (N_165,In_1673,In_294);
nand U166 (N_166,In_894,In_1222);
nand U167 (N_167,In_1616,In_1307);
and U168 (N_168,In_1510,In_2934);
and U169 (N_169,In_64,In_2674);
nand U170 (N_170,In_2966,In_1101);
nand U171 (N_171,In_628,In_2213);
nor U172 (N_172,In_1221,In_135);
xor U173 (N_173,In_672,In_536);
nand U174 (N_174,In_1427,In_2094);
nand U175 (N_175,In_2190,In_2681);
xor U176 (N_176,In_1095,In_1728);
nor U177 (N_177,In_1250,In_2083);
or U178 (N_178,In_1217,In_1216);
nand U179 (N_179,In_1111,In_816);
nand U180 (N_180,In_17,In_247);
and U181 (N_181,In_1477,In_630);
or U182 (N_182,In_2961,In_944);
or U183 (N_183,In_899,In_2318);
nor U184 (N_184,In_715,In_1407);
nor U185 (N_185,In_2408,In_411);
and U186 (N_186,In_1633,In_1602);
nand U187 (N_187,In_1873,In_551);
or U188 (N_188,In_2623,In_268);
or U189 (N_189,In_2098,In_590);
and U190 (N_190,In_840,In_2965);
and U191 (N_191,In_2401,In_175);
and U192 (N_192,In_233,In_1912);
nand U193 (N_193,In_2649,In_980);
or U194 (N_194,In_1753,In_626);
nand U195 (N_195,In_1957,In_2150);
and U196 (N_196,In_394,In_2064);
and U197 (N_197,In_1841,In_271);
nor U198 (N_198,In_682,In_1831);
nand U199 (N_199,In_1078,In_882);
and U200 (N_200,In_317,In_1066);
and U201 (N_201,In_2841,In_1139);
and U202 (N_202,In_1848,In_2884);
or U203 (N_203,In_1534,In_1650);
xnor U204 (N_204,In_946,In_2259);
nand U205 (N_205,In_2542,In_1702);
nand U206 (N_206,In_2564,In_503);
xor U207 (N_207,In_2343,In_71);
xor U208 (N_208,In_1336,In_738);
nand U209 (N_209,In_1368,In_852);
xnor U210 (N_210,In_1192,In_2845);
nor U211 (N_211,In_1970,In_1815);
nor U212 (N_212,In_1648,In_2376);
and U213 (N_213,In_308,In_2943);
nand U214 (N_214,In_2796,In_663);
or U215 (N_215,In_1706,In_2740);
or U216 (N_216,In_1437,In_2977);
and U217 (N_217,In_897,In_1664);
nand U218 (N_218,In_1964,In_698);
nand U219 (N_219,In_2255,In_2237);
or U220 (N_220,In_137,In_1976);
nand U221 (N_221,In_401,In_2207);
and U222 (N_222,In_2220,In_259);
and U223 (N_223,In_2244,In_2592);
and U224 (N_224,In_374,In_704);
nand U225 (N_225,In_2671,In_1335);
nor U226 (N_226,In_2990,In_701);
or U227 (N_227,In_304,In_2775);
or U228 (N_228,In_63,In_32);
xnor U229 (N_229,In_2304,In_1136);
nand U230 (N_230,In_2664,In_1857);
nand U231 (N_231,In_2320,In_489);
or U232 (N_232,In_2449,In_212);
or U233 (N_233,In_599,In_1060);
nand U234 (N_234,In_20,In_312);
nand U235 (N_235,In_2026,In_1625);
nor U236 (N_236,In_1656,In_2676);
nor U237 (N_237,In_1138,In_688);
and U238 (N_238,In_69,In_2151);
or U239 (N_239,In_1624,In_813);
and U240 (N_240,In_342,In_2548);
or U241 (N_241,In_125,In_1516);
or U242 (N_242,In_1421,In_377);
or U243 (N_243,In_1820,In_1797);
xor U244 (N_244,In_865,In_200);
or U245 (N_245,In_2289,In_514);
and U246 (N_246,In_1484,In_1779);
and U247 (N_247,In_1600,In_2830);
and U248 (N_248,In_1399,In_1918);
nor U249 (N_249,In_2758,In_220);
or U250 (N_250,In_291,In_2940);
nor U251 (N_251,In_2125,In_2838);
or U252 (N_252,In_1795,In_1004);
or U253 (N_253,In_353,In_1088);
nor U254 (N_254,In_2591,In_1911);
and U255 (N_255,In_2896,In_2779);
nand U256 (N_256,In_2122,In_2154);
or U257 (N_257,In_2624,In_2103);
nand U258 (N_258,In_1402,In_1116);
and U259 (N_259,In_307,In_1876);
nor U260 (N_260,In_2087,In_2737);
nand U261 (N_261,In_2729,In_2374);
or U262 (N_262,In_1462,In_1994);
or U263 (N_263,In_2912,In_1094);
or U264 (N_264,In_219,In_1001);
nand U265 (N_265,In_2503,In_1498);
nor U266 (N_266,In_2079,In_654);
nand U267 (N_267,In_1612,In_2786);
nor U268 (N_268,In_2439,In_695);
nand U269 (N_269,In_1590,In_1328);
xor U270 (N_270,In_50,In_1734);
xnor U271 (N_271,In_1869,In_1159);
or U272 (N_272,In_2299,In_366);
nor U273 (N_273,In_250,In_2001);
nand U274 (N_274,In_2774,In_691);
nand U275 (N_275,In_480,In_781);
nor U276 (N_276,In_1704,In_2228);
xnor U277 (N_277,In_276,In_348);
xor U278 (N_278,In_2069,In_914);
nand U279 (N_279,In_1874,In_720);
and U280 (N_280,In_2987,In_1459);
nor U281 (N_281,In_869,In_1483);
and U282 (N_282,In_875,In_2392);
nand U283 (N_283,In_1031,In_157);
and U284 (N_284,In_483,In_2799);
nand U285 (N_285,In_1167,In_2359);
and U286 (N_286,In_2235,In_1660);
nor U287 (N_287,In_2424,In_2149);
and U288 (N_288,In_319,In_1866);
xor U289 (N_289,In_1629,In_812);
or U290 (N_290,In_2006,In_1188);
or U291 (N_291,In_1142,In_216);
nand U292 (N_292,In_2791,In_2309);
xor U293 (N_293,In_2295,In_188);
nand U294 (N_294,In_2283,In_466);
nand U295 (N_295,In_2600,In_1885);
and U296 (N_296,In_1791,In_2898);
and U297 (N_297,In_1941,In_1952);
nand U298 (N_298,In_603,In_633);
xor U299 (N_299,In_1890,In_2136);
nor U300 (N_300,In_2099,In_1191);
and U301 (N_301,In_2741,In_145);
and U302 (N_302,In_1229,In_2790);
or U303 (N_303,In_1341,In_978);
nand U304 (N_304,In_765,In_1269);
and U305 (N_305,In_597,In_2045);
nor U306 (N_306,In_1827,In_2981);
and U307 (N_307,In_1347,In_448);
nor U308 (N_308,In_300,In_2223);
and U309 (N_309,In_2538,In_1746);
and U310 (N_310,In_803,In_248);
nand U311 (N_311,In_1416,In_1428);
and U312 (N_312,In_2820,In_2022);
nand U313 (N_313,In_1264,In_646);
and U314 (N_314,In_2469,In_1375);
nor U315 (N_315,In_2817,In_1053);
nand U316 (N_316,In_1120,In_997);
nand U317 (N_317,In_2373,In_1900);
and U318 (N_318,In_2508,In_544);
or U319 (N_319,In_1014,In_227);
or U320 (N_320,In_1256,In_2666);
xnor U321 (N_321,In_1710,In_1331);
nor U322 (N_322,In_1124,In_2135);
nor U323 (N_323,In_371,In_388);
and U324 (N_324,In_2313,In_1531);
nor U325 (N_325,In_1141,In_2889);
xnor U326 (N_326,In_984,In_1835);
nand U327 (N_327,In_2199,In_1551);
xor U328 (N_328,In_2249,In_1097);
nor U329 (N_329,In_1640,In_2434);
or U330 (N_330,In_2307,In_182);
xor U331 (N_331,In_2049,In_390);
or U332 (N_332,In_381,In_1005);
and U333 (N_333,In_948,In_2500);
nor U334 (N_334,In_1830,In_1669);
nor U335 (N_335,In_635,In_1729);
or U336 (N_336,In_162,In_2689);
or U337 (N_337,In_1853,In_1404);
nor U338 (N_338,In_1582,In_256);
nand U339 (N_339,In_1350,In_2938);
nand U340 (N_340,In_1517,In_1230);
nand U341 (N_341,In_2396,In_2387);
xnor U342 (N_342,In_1226,In_2018);
or U343 (N_343,In_232,In_569);
and U344 (N_344,In_2275,In_2380);
and U345 (N_345,In_26,In_2491);
and U346 (N_346,In_2367,In_2330);
xor U347 (N_347,In_2608,In_1487);
and U348 (N_348,In_1405,In_1419);
or U349 (N_349,In_1103,In_526);
or U350 (N_350,In_1266,In_2166);
or U351 (N_351,In_1884,In_1533);
nor U352 (N_352,In_1609,In_863);
nand U353 (N_353,In_2025,In_1491);
or U354 (N_354,In_1822,In_1751);
and U355 (N_355,In_1816,In_2808);
and U356 (N_356,In_833,In_1832);
nand U357 (N_357,In_2075,In_2121);
nor U358 (N_358,In_2900,In_75);
nand U359 (N_359,In_1494,In_155);
and U360 (N_360,In_1236,In_518);
and U361 (N_361,In_2699,In_1865);
and U362 (N_362,In_558,In_421);
nand U363 (N_363,In_699,In_1284);
nand U364 (N_364,In_2333,In_1173);
or U365 (N_365,In_1542,In_2915);
and U366 (N_366,In_363,In_2381);
nor U367 (N_367,In_1356,In_2653);
and U368 (N_368,In_2855,In_2415);
nor U369 (N_369,In_2250,In_2390);
nor U370 (N_370,In_1917,In_59);
xnor U371 (N_371,In_1735,In_1134);
xor U372 (N_372,In_1429,In_941);
nand U373 (N_373,In_521,In_324);
nand U374 (N_374,In_2118,In_611);
xnor U375 (N_375,In_1050,In_999);
and U376 (N_376,In_393,In_2716);
nand U377 (N_377,In_1677,In_1218);
nand U378 (N_378,In_2593,In_1995);
xnor U379 (N_379,In_2634,In_1544);
or U380 (N_380,In_961,In_1698);
or U381 (N_381,In_836,In_913);
nor U382 (N_382,In_2474,In_44);
nor U383 (N_383,In_435,In_1093);
nor U384 (N_384,In_77,In_1271);
or U385 (N_385,In_1283,In_2847);
xor U386 (N_386,In_1212,In_2995);
and U387 (N_387,In_1408,In_2763);
and U388 (N_388,In_491,In_896);
or U389 (N_389,In_707,In_623);
nand U390 (N_390,In_685,In_2705);
nand U391 (N_391,In_2812,In_1690);
nand U392 (N_392,In_874,In_951);
nand U393 (N_393,In_1583,In_1200);
nand U394 (N_394,In_351,In_1863);
and U395 (N_395,In_1085,In_601);
nor U396 (N_396,In_195,In_2056);
xor U397 (N_397,In_1945,In_242);
nor U398 (N_398,In_1807,In_2827);
or U399 (N_399,In_408,In_2742);
and U400 (N_400,In_1856,In_419);
and U401 (N_401,In_1228,In_2143);
nand U402 (N_402,In_2933,In_214);
xor U403 (N_403,In_2361,In_79);
and U404 (N_404,In_1146,In_2159);
nand U405 (N_405,In_1987,In_1041);
or U406 (N_406,In_1395,In_1022);
nor U407 (N_407,In_340,In_620);
or U408 (N_408,In_103,In_2221);
and U409 (N_409,In_1071,In_1804);
or U410 (N_410,In_2115,In_12);
nor U411 (N_411,In_1715,In_2554);
and U412 (N_412,In_848,In_2463);
nand U413 (N_413,In_998,In_2130);
or U414 (N_414,In_1978,In_2454);
and U415 (N_415,In_1086,In_1537);
nor U416 (N_416,In_2733,In_2736);
nand U417 (N_417,In_2090,In_2301);
or U418 (N_418,In_2525,In_1798);
and U419 (N_419,In_1426,In_2410);
xor U420 (N_420,In_1638,In_573);
and U421 (N_421,In_1708,In_2534);
xnor U422 (N_422,In_759,In_2431);
and U423 (N_423,In_2048,In_1058);
nand U424 (N_424,In_48,In_2407);
nor U425 (N_425,In_1259,In_1748);
nand U426 (N_426,In_2175,In_832);
or U427 (N_427,In_1205,In_2787);
nand U428 (N_428,In_1090,In_1076);
nand U429 (N_429,In_345,In_2754);
xnor U430 (N_430,In_1267,In_1449);
or U431 (N_431,In_1956,In_636);
nor U432 (N_432,In_2247,In_1688);
nor U433 (N_433,In_2498,In_1045);
nand U434 (N_434,In_1496,In_502);
or U435 (N_435,In_2887,In_2825);
nor U436 (N_436,In_412,In_2706);
nand U437 (N_437,In_2583,In_60);
nand U438 (N_438,In_144,In_1842);
xor U439 (N_439,In_1089,In_2248);
nand U440 (N_440,In_2034,In_1755);
nand U441 (N_441,In_2395,In_1538);
nor U442 (N_442,In_2433,In_2520);
nand U443 (N_443,In_2496,In_901);
nor U444 (N_444,In_645,In_1409);
nor U445 (N_445,In_352,In_2063);
nor U446 (N_446,In_334,In_728);
and U447 (N_447,In_2364,In_1215);
and U448 (N_448,In_2033,In_1758);
or U449 (N_449,In_804,In_1002);
nor U450 (N_450,In_2879,In_1904);
or U451 (N_451,In_303,In_2515);
nand U452 (N_452,In_2971,In_975);
or U453 (N_453,In_746,In_782);
and U454 (N_454,In_2502,In_2890);
xnor U455 (N_455,In_1067,In_2924);
nand U456 (N_456,In_131,In_1418);
or U457 (N_457,In_1764,In_2651);
or U458 (N_458,In_985,In_85);
nand U459 (N_459,In_807,In_976);
nor U460 (N_460,In_2412,In_1683);
or U461 (N_461,In_2945,In_1174);
nor U462 (N_462,In_265,In_954);
nor U463 (N_463,In_1,In_1889);
nor U464 (N_464,In_2413,In_1410);
nor U465 (N_465,In_2584,In_471);
xor U466 (N_466,In_1971,In_1472);
nor U467 (N_467,In_380,In_2596);
xnor U468 (N_468,In_777,In_1369);
or U469 (N_469,In_58,In_1171);
and U470 (N_470,In_1028,In_1342);
or U471 (N_471,In_1059,In_1770);
or U472 (N_472,In_1270,In_38);
and U473 (N_473,In_809,In_638);
xnor U474 (N_474,In_2409,In_1343);
xor U475 (N_475,In_2656,In_343);
or U476 (N_476,In_1394,In_111);
and U477 (N_477,In_296,In_1705);
and U478 (N_478,In_2501,In_1460);
or U479 (N_479,In_1258,In_2062);
xnor U480 (N_480,In_2252,In_1011);
or U481 (N_481,In_2696,In_1296);
xnor U482 (N_482,In_1579,In_1322);
nand U483 (N_483,In_1340,In_2314);
and U484 (N_484,In_2639,In_1008);
nor U485 (N_485,In_1557,In_1950);
nand U486 (N_486,In_1659,In_621);
xnor U487 (N_487,In_2660,In_786);
and U488 (N_488,In_598,In_1849);
or U489 (N_489,In_373,In_904);
nand U490 (N_490,In_1543,In_531);
nor U491 (N_491,In_2635,In_1225);
and U492 (N_492,In_679,In_266);
or U493 (N_493,In_2494,In_2317);
xnor U494 (N_494,In_1774,In_305);
or U495 (N_495,In_1346,In_1027);
xnor U496 (N_496,In_2459,In_2579);
nand U497 (N_497,In_1913,In_2437);
and U498 (N_498,In_1727,In_2602);
nor U499 (N_499,In_1232,In_731);
nand U500 (N_500,In_1555,In_1522);
and U501 (N_501,In_1412,In_1069);
or U502 (N_502,In_2245,In_129);
and U503 (N_503,In_2750,In_1476);
nor U504 (N_504,In_330,In_1597);
or U505 (N_505,In_1578,In_721);
and U506 (N_506,In_2678,In_1376);
nor U507 (N_507,In_898,In_487);
nand U508 (N_508,In_2286,In_2371);
nand U509 (N_509,In_203,In_223);
nor U510 (N_510,In_2974,In_2455);
or U511 (N_511,In_2164,In_1707);
and U512 (N_512,In_2690,In_263);
and U513 (N_513,In_1280,In_886);
or U514 (N_514,In_861,In_2680);
nor U515 (N_515,In_2328,In_2310);
and U516 (N_516,In_2342,In_2436);
xor U517 (N_517,In_1909,In_121);
nor U518 (N_518,In_459,In_2119);
or U519 (N_519,In_490,In_986);
nand U520 (N_520,In_706,In_2954);
and U521 (N_521,In_1025,In_1389);
and U522 (N_522,In_1360,In_2980);
nor U523 (N_523,In_2507,In_768);
xnor U524 (N_524,In_78,In_1888);
and U525 (N_525,In_115,In_2174);
nand U526 (N_526,In_543,In_2505);
and U527 (N_527,In_2872,In_314);
nand U528 (N_528,In_1509,In_1275);
and U529 (N_529,In_2183,In_425);
or U530 (N_530,In_2572,In_284);
or U531 (N_531,In_602,In_1851);
or U532 (N_532,In_1072,In_2964);
or U533 (N_533,In_1665,In_2441);
nand U534 (N_534,In_2486,In_2573);
xnor U535 (N_535,In_2192,In_1684);
nor U536 (N_536,In_1962,In_1490);
nand U537 (N_537,In_2269,In_880);
and U538 (N_538,In_2102,In_8);
and U539 (N_539,In_2404,In_2776);
xor U540 (N_540,In_1096,In_1968);
nand U541 (N_541,In_500,In_292);
nand U542 (N_542,In_1006,In_105);
nand U543 (N_543,In_369,In_2901);
nor U544 (N_544,In_61,In_507);
and U545 (N_545,In_1773,In_1662);
or U546 (N_546,In_2802,In_2068);
and U547 (N_547,In_2687,In_2461);
or U548 (N_548,In_2234,In_87);
or U549 (N_549,In_2873,In_1763);
nand U550 (N_550,In_2526,In_2955);
and U551 (N_551,In_737,In_887);
xor U552 (N_552,In_1242,In_2080);
or U553 (N_553,In_152,In_1864);
nor U554 (N_554,In_1605,In_2178);
or U555 (N_555,In_237,In_1577);
and U556 (N_556,In_1826,In_2642);
and U557 (N_557,In_42,In_1529);
nor U558 (N_558,In_2570,In_2096);
and U559 (N_559,In_1618,In_497);
nor U560 (N_560,In_556,In_2517);
xor U561 (N_561,In_2337,In_449);
nand U562 (N_562,In_1313,In_1373);
and U563 (N_563,In_2784,In_923);
and U564 (N_564,In_1836,In_2391);
or U565 (N_565,In_2160,In_2636);
nor U566 (N_566,In_785,In_810);
or U567 (N_567,In_102,In_1023);
and U568 (N_568,In_2886,In_349);
nor U569 (N_569,In_150,In_1630);
and U570 (N_570,In_1430,In_2229);
nand U571 (N_571,In_668,In_967);
xor U572 (N_572,In_1391,In_2043);
or U573 (N_573,In_1949,In_647);
or U574 (N_574,In_492,In_1179);
nand U575 (N_575,In_1026,In_1922);
and U576 (N_576,In_1042,In_387);
or U577 (N_577,In_921,In_2107);
nor U578 (N_578,In_167,In_1634);
and U579 (N_579,In_2017,In_684);
nor U580 (N_580,In_1966,In_1048);
nor U581 (N_581,In_1233,In_2717);
and U582 (N_582,In_479,In_2279);
or U583 (N_583,In_928,In_2700);
and U584 (N_584,In_1495,In_644);
or U585 (N_585,In_81,In_1527);
nor U586 (N_586,In_2176,In_871);
nand U587 (N_587,In_727,In_2863);
or U588 (N_588,In_2616,In_1020);
nor U589 (N_589,In_2695,In_1573);
and U590 (N_590,In_1661,In_2853);
nand U591 (N_591,In_2116,In_1440);
or U592 (N_592,In_709,In_589);
nor U593 (N_593,In_1393,In_1289);
nor U594 (N_594,In_161,In_1312);
or U595 (N_595,In_2902,In_1223);
nor U596 (N_596,In_508,In_958);
nand U597 (N_597,In_2744,In_1074);
nor U598 (N_598,In_1515,In_92);
nand U599 (N_599,In_1211,In_627);
and U600 (N_600,In_680,In_1110);
or U601 (N_601,In_1486,In_1334);
nand U602 (N_602,In_1034,In_2932);
xnor U603 (N_603,In_1972,In_2629);
nor U604 (N_604,In_541,In_625);
xor U605 (N_605,In_1276,In_2806);
and U606 (N_606,In_1339,In_1300);
or U607 (N_607,In_1716,In_2258);
nor U608 (N_608,In_1306,In_1757);
and U609 (N_609,In_2540,In_2645);
and U610 (N_610,In_2460,In_2911);
and U611 (N_611,In_443,In_339);
nand U612 (N_612,In_1442,In_819);
nand U613 (N_613,In_1457,In_2173);
nand U614 (N_614,In_68,In_2261);
xor U615 (N_615,In_1033,In_482);
nor U616 (N_616,In_2013,In_2360);
and U617 (N_617,In_1828,In_253);
and U618 (N_618,In_2557,In_2113);
nor U619 (N_619,In_1241,In_1697);
xor U620 (N_620,In_1586,In_2868);
and U621 (N_621,In_608,In_101);
nor U622 (N_622,In_2541,In_2617);
nand U623 (N_623,In_2358,In_147);
or U624 (N_624,In_1161,In_306);
or U625 (N_625,In_2051,In_511);
and U626 (N_626,In_1100,In_966);
nand U627 (N_627,In_596,In_146);
nand U628 (N_628,In_2504,In_1295);
nand U629 (N_629,In_2292,In_1718);
nand U630 (N_630,In_1933,In_815);
nor U631 (N_631,In_552,In_236);
nand U632 (N_632,In_2628,In_2184);
nand U633 (N_633,In_1672,In_288);
or U634 (N_634,In_2108,In_2257);
or U635 (N_635,In_2803,In_2749);
or U636 (N_636,In_519,In_2837);
or U637 (N_637,In_2821,In_2089);
nand U638 (N_638,In_2353,In_2718);
nor U639 (N_639,In_1696,In_1601);
or U640 (N_640,In_876,In_1406);
xor U641 (N_641,In_422,In_1443);
and U642 (N_642,In_889,In_1977);
nand U643 (N_643,In_1926,In_2562);
xnor U644 (N_644,In_2801,In_1530);
and U645 (N_645,In_2231,In_2177);
and U646 (N_646,In_1989,In_2665);
nand U647 (N_647,In_1140,In_1362);
and U648 (N_648,In_260,In_311);
nor U649 (N_649,In_2348,In_2952);
or U650 (N_650,In_881,In_2646);
nand U651 (N_651,In_1740,In_1401);
and U652 (N_652,In_2464,In_2611);
and U653 (N_653,In_2423,In_629);
and U654 (N_654,In_2351,In_581);
and U655 (N_655,In_2654,In_915);
or U656 (N_656,In_134,In_2106);
xnor U657 (N_657,In_1536,In_2904);
and U658 (N_658,In_2430,In_1935);
and U659 (N_659,In_754,In_2042);
nor U660 (N_660,In_2382,In_2482);
nand U661 (N_661,In_142,In_2519);
and U662 (N_662,In_1272,In_1453);
nand U663 (N_663,In_1713,In_16);
nor U664 (N_664,In_1308,In_1540);
nor U665 (N_665,In_2195,In_2179);
and U666 (N_666,In_2465,In_2941);
nand U667 (N_667,In_2256,In_464);
or U668 (N_668,In_977,In_750);
nand U669 (N_669,In_2129,In_481);
nor U670 (N_670,In_2532,In_40);
or U671 (N_671,In_2338,In_1244);
or U672 (N_672,In_2053,In_1182);
or U673 (N_673,In_1645,In_2759);
and U674 (N_674,In_151,In_2035);
nor U675 (N_675,In_2274,In_1181);
or U676 (N_676,In_752,In_208);
and U677 (N_677,In_965,In_1281);
or U678 (N_678,In_426,In_2597);
and U679 (N_679,In_2205,In_7);
nand U680 (N_680,In_94,In_1252);
nand U681 (N_681,In_2340,In_1469);
or U682 (N_682,In_2484,In_811);
or U683 (N_683,In_467,In_606);
xnor U684 (N_684,In_2708,In_2589);
xnor U685 (N_685,In_1658,In_2893);
or U686 (N_686,In_2188,In_2726);
and U687 (N_687,In_868,In_181);
nor U688 (N_688,In_2804,In_2547);
xor U689 (N_689,In_1279,In_1372);
xor U690 (N_690,In_2957,In_2110);
and U691 (N_691,In_159,In_517);
or U692 (N_692,In_1463,In_1860);
nand U693 (N_693,In_964,In_329);
or U694 (N_694,In_2305,In_1273);
nor U695 (N_695,In_2641,In_2242);
and U696 (N_696,In_2146,In_655);
and U697 (N_697,In_1984,In_837);
nand U698 (N_698,In_911,In_2613);
xnor U699 (N_699,In_1325,In_2626);
or U700 (N_700,In_346,In_857);
and U701 (N_701,In_409,In_1203);
nand U702 (N_702,In_2644,In_2773);
nor U703 (N_703,In_2850,In_687);
xnor U704 (N_704,In_403,In_766);
nor U705 (N_705,In_2354,In_582);
nor U706 (N_706,In_822,In_1975);
nor U707 (N_707,In_2693,In_6);
and U708 (N_708,In_384,In_760);
nand U709 (N_709,In_2278,In_1492);
nand U710 (N_710,In_469,In_295);
and U711 (N_711,In_179,In_2161);
and U712 (N_712,In_84,In_2731);
or U713 (N_713,In_1932,In_2552);
nor U714 (N_714,In_1183,In_2948);
nor U715 (N_715,In_2521,In_1614);
nand U716 (N_716,In_2655,In_979);
nor U717 (N_717,In_1130,In_1447);
or U718 (N_718,In_713,In_273);
or U719 (N_719,In_858,In_918);
nand U720 (N_720,In_926,In_450);
and U721 (N_721,In_2240,In_2522);
nor U722 (N_722,In_54,In_35);
and U723 (N_723,In_2686,In_1445);
or U724 (N_724,In_827,In_745);
nor U725 (N_725,In_548,In_1545);
or U726 (N_726,In_2489,In_1761);
and U727 (N_727,In_2568,In_1709);
xnor U728 (N_728,In_2029,In_1920);
and U729 (N_729,In_1620,In_1352);
or U730 (N_730,In_1243,In_174);
nor U731 (N_731,In_1743,In_1044);
or U732 (N_732,In_1717,In_1384);
and U733 (N_733,In_864,In_283);
or U734 (N_734,In_2959,In_2397);
nor U735 (N_735,In_1817,In_468);
nor U736 (N_736,In_2162,In_1303);
or U737 (N_737,In_1077,In_2860);
or U738 (N_738,In_488,In_1210);
nand U739 (N_739,In_2647,In_824);
nor U740 (N_740,In_2456,In_2157);
nand U741 (N_741,In_1671,In_2086);
nand U742 (N_742,In_878,In_1871);
nand U743 (N_743,In_583,In_585);
nor U744 (N_744,In_66,In_808);
xnor U745 (N_745,In_287,In_1628);
and U746 (N_746,In_2834,In_74);
or U747 (N_747,In_2587,In_2362);
and U748 (N_748,In_429,In_347);
nand U749 (N_749,In_1029,In_189);
or U750 (N_750,In_673,In_2950);
nand U751 (N_751,In_397,In_1380);
xnor U752 (N_752,In_86,In_1750);
and U753 (N_753,In_568,In_1417);
and U754 (N_754,In_2277,In_1000);
xnor U755 (N_755,In_1018,In_1160);
xor U756 (N_756,In_2466,In_528);
nand U757 (N_757,In_1703,In_2607);
or U758 (N_758,In_477,In_674);
or U759 (N_759,In_2824,In_1896);
xnor U760 (N_760,In_995,In_2440);
nor U761 (N_761,In_2398,In_5);
or U762 (N_762,In_1112,In_1613);
nor U763 (N_763,In_2356,In_592);
and U764 (N_764,In_634,In_1654);
nand U765 (N_765,In_1148,In_1468);
nand U766 (N_766,In_2117,In_1310);
and U767 (N_767,In_641,In_829);
nor U768 (N_768,In_1581,In_436);
nand U769 (N_769,In_1015,In_842);
nor U770 (N_770,In_1268,In_1631);
nor U771 (N_771,In_2287,In_755);
and U772 (N_772,In_2612,In_1499);
or U773 (N_773,In_2156,In_2369);
nor U774 (N_774,In_726,In_2867);
or U775 (N_775,In_994,In_2882);
or U776 (N_776,In_2211,In_2846);
and U777 (N_777,In_1595,In_1759);
nand U778 (N_778,In_2230,In_1719);
nor U779 (N_779,In_2714,In_719);
xnor U780 (N_780,In_1425,In_723);
or U781 (N_781,In_1108,In_22);
nor U782 (N_782,In_2631,In_509);
nand U783 (N_783,In_2743,In_2435);
nand U784 (N_784,In_2402,In_2302);
or U785 (N_785,In_2124,In_138);
or U786 (N_786,In_364,In_1030);
xor U787 (N_787,In_2059,In_2481);
nand U788 (N_788,In_2983,In_947);
and U789 (N_789,In_2625,In_2357);
and U790 (N_790,In_1304,In_2047);
and U791 (N_791,In_1778,In_278);
nand U792 (N_792,In_712,In_1370);
and U793 (N_793,In_1901,In_2661);
nor U794 (N_794,In_1396,In_2958);
and U795 (N_795,In_270,In_1434);
xnor U796 (N_796,In_725,In_2996);
nand U797 (N_797,In_1366,In_1646);
or U798 (N_798,In_662,In_866);
or U799 (N_799,In_925,In_1599);
or U800 (N_800,In_365,In_733);
and U801 (N_801,In_2271,In_1435);
and U802 (N_802,In_2478,In_2202);
nor U803 (N_803,In_1998,In_2497);
nor U804 (N_804,In_744,In_2710);
nor U805 (N_805,In_184,In_1809);
and U806 (N_806,In_798,In_2123);
nand U807 (N_807,In_2411,In_1939);
nor U808 (N_808,In_2138,In_2929);
and U809 (N_809,In_1196,In_210);
nand U810 (N_810,In_141,In_2586);
or U811 (N_811,In_931,In_2272);
and U812 (N_812,In_605,In_136);
xnor U813 (N_813,In_1598,In_2595);
nand U814 (N_814,In_872,In_1318);
nand U815 (N_815,In_751,In_2088);
or U816 (N_816,In_2854,In_575);
xor U817 (N_817,In_2216,In_226);
nand U818 (N_818,In_1361,In_1891);
or U819 (N_819,In_439,In_2352);
nand U820 (N_820,In_814,In_2324);
and U821 (N_821,In_1566,In_1194);
or U822 (N_822,In_1286,In_2662);
nor U823 (N_823,In_2865,In_2899);
xnor U824 (N_824,In_2296,In_1037);
nand U825 (N_825,In_2298,In_243);
nand U826 (N_826,In_1556,In_1615);
xor U827 (N_827,In_2914,In_2007);
and U828 (N_828,In_2168,In_11);
or U829 (N_829,In_2008,In_2097);
nor U830 (N_830,In_1676,In_1726);
or U831 (N_831,In_2002,In_154);
nand U832 (N_832,In_2615,In_2319);
or U833 (N_833,In_830,In_2663);
or U834 (N_834,In_1986,In_2334);
xnor U835 (N_835,In_2857,In_686);
and U836 (N_836,In_2335,In_110);
or U837 (N_837,In_1013,In_2604);
nor U838 (N_838,In_2443,In_297);
xor U839 (N_839,In_862,In_1760);
and U840 (N_840,In_1187,In_1043);
nor U841 (N_841,In_2851,In_119);
and U842 (N_842,In_2322,In_1290);
nand U843 (N_843,In_2070,In_1554);
nand U844 (N_844,In_2692,In_1528);
nand U845 (N_845,In_823,In_1010);
xor U846 (N_846,In_2189,In_1169);
nand U847 (N_847,In_120,In_2523);
or U848 (N_848,In_2580,In_849);
and U849 (N_849,In_793,In_1621);
or U850 (N_850,In_1301,In_2363);
nor U851 (N_851,In_486,In_1507);
nor U852 (N_852,In_651,In_1087);
and U853 (N_853,In_2239,In_1559);
nor U854 (N_854,In_1052,In_2719);
or U855 (N_855,In_2290,In_289);
and U856 (N_856,In_1800,In_2724);
nand U857 (N_857,In_2227,In_2426);
or U858 (N_858,In_1927,In_788);
nor U859 (N_859,In_2963,In_91);
or U860 (N_860,In_143,In_2594);
xor U861 (N_861,In_1371,In_1098);
nand U862 (N_862,In_2876,In_1737);
nor U863 (N_863,In_831,In_2315);
xor U864 (N_864,In_1024,In_2432);
and U865 (N_865,In_376,In_1679);
nor U866 (N_866,In_2762,In_30);
or U867 (N_867,In_711,In_1570);
nor U868 (N_868,In_1282,In_413);
nand U869 (N_869,In_275,In_2293);
nor U870 (N_870,In_2777,In_2134);
nor U871 (N_871,In_2066,In_736);
nor U872 (N_872,In_2180,In_1765);
nand U873 (N_873,In_855,In_571);
and U874 (N_874,In_539,In_0);
or U875 (N_875,In_643,In_149);
nand U876 (N_876,In_2870,In_1297);
and U877 (N_877,In_1954,In_1667);
nor U878 (N_878,In_420,In_534);
or U879 (N_879,In_884,In_545);
nand U880 (N_880,In_2200,In_1730);
and U881 (N_881,In_2186,In_2669);
and U882 (N_882,In_2273,In_669);
nand U883 (N_883,In_1176,In_2632);
xnor U884 (N_884,In_1255,In_2386);
nor U885 (N_885,In_24,In_2691);
or U886 (N_886,In_1738,In_1080);
nor U887 (N_887,In_2316,In_2442);
nand U888 (N_888,In_1790,In_1923);
or U889 (N_889,In_697,In_1178);
nor U890 (N_890,In_410,In_2);
xnor U891 (N_891,In_2947,In_1999);
nor U892 (N_892,In_230,In_406);
xor U893 (N_893,In_934,In_1951);
nand U894 (N_894,In_1185,In_2028);
nand U895 (N_895,In_2462,In_43);
or U896 (N_896,In_2253,In_209);
nor U897 (N_897,In_2512,In_2539);
xor U898 (N_898,In_156,In_2148);
or U899 (N_899,In_2956,In_1063);
nand U900 (N_900,In_2372,In_1714);
xor U901 (N_901,In_1905,In_1821);
nand U902 (N_902,In_1068,In_2781);
nand U903 (N_903,In_2060,In_2832);
nand U904 (N_904,In_909,In_2745);
and U905 (N_905,In_128,In_1471);
and U906 (N_906,In_2236,In_1348);
and U907 (N_907,In_2480,In_215);
xor U908 (N_908,In_2771,In_658);
or U909 (N_909,In_693,In_414);
xnor U910 (N_910,In_2588,In_1184);
nor U911 (N_911,In_555,In_1675);
and U912 (N_912,In_1204,In_118);
nor U913 (N_913,In_2262,In_1903);
xor U914 (N_914,In_281,In_1032);
nand U915 (N_915,In_2985,In_2233);
and U916 (N_916,In_1783,In_1589);
nand U917 (N_917,In_1127,In_729);
nand U918 (N_918,In_2894,In_2311);
nor U919 (N_919,In_201,In_772);
nand U920 (N_920,In_1314,In_1458);
and U921 (N_921,In_2765,In_2930);
nor U922 (N_922,In_3,In_2294);
or U923 (N_923,In_1607,In_1450);
or U924 (N_924,In_2321,In_427);
nor U925 (N_925,In_1153,In_2670);
and U926 (N_926,In_616,In_1924);
nand U927 (N_927,In_2927,In_1814);
nor U928 (N_928,In_642,In_1363);
nor U929 (N_929,In_1643,In_1752);
and U930 (N_930,In_2421,In_395);
nand U931 (N_931,In_2020,In_235);
nor U932 (N_932,In_1254,In_1337);
nand U933 (N_933,In_1175,In_792);
nand U934 (N_934,In_1151,In_2152);
and U935 (N_935,In_565,In_1392);
xnor U936 (N_936,In_1711,In_1154);
nand U937 (N_937,In_2614,In_1237);
nor U938 (N_938,In_2761,In_211);
nand U939 (N_939,In_2037,In_1390);
or U940 (N_940,In_194,In_49);
nand U941 (N_941,In_996,In_2078);
or U942 (N_942,In_1379,In_1261);
nand U943 (N_943,In_2962,In_741);
nor U944 (N_944,In_1993,In_165);
xnor U945 (N_945,In_461,In_838);
or U946 (N_946,In_191,In_1603);
nand U947 (N_947,In_650,In_2536);
and U948 (N_948,In_2810,In_764);
nor U949 (N_949,In_1488,In_2420);
or U950 (N_950,In_850,In_902);
and U951 (N_951,In_2909,In_1948);
nor U952 (N_952,In_359,In_1887);
nand U953 (N_953,In_2475,In_108);
or U954 (N_954,In_2417,In_2575);
nand U955 (N_955,In_530,In_783);
nor U956 (N_956,In_2339,In_1481);
and U957 (N_957,In_1539,In_2429);
and U958 (N_958,In_1055,In_2477);
nand U959 (N_959,In_310,In_485);
nand U960 (N_960,In_2668,In_229);
nand U961 (N_961,In_1868,In_1635);
xnor U962 (N_962,In_2582,In_391);
and U963 (N_963,In_2770,In_1733);
or U964 (N_964,In_2450,In_1382);
or U965 (N_965,In_1158,In_57);
and U966 (N_966,In_1305,In_1567);
nor U967 (N_967,In_238,In_1357);
nand U968 (N_968,In_1594,In_51);
nand U969 (N_969,In_2513,In_1324);
or U970 (N_970,In_692,In_252);
and U971 (N_971,In_96,In_2738);
and U972 (N_972,In_891,In_2493);
nor U973 (N_973,In_2610,In_2329);
nor U974 (N_974,In_218,In_1201);
xnor U975 (N_975,In_1021,In_2537);
nand U976 (N_976,In_1619,In_27);
or U977 (N_977,In_192,In_2378);
nor U978 (N_978,In_2297,In_2683);
xnor U979 (N_979,In_438,In_1550);
nand U980 (N_980,In_520,In_1239);
nand U981 (N_981,In_938,In_2768);
and U982 (N_982,In_484,In_279);
xor U983 (N_983,In_1694,In_800);
xor U984 (N_984,In_968,In_2238);
or U985 (N_985,In_1647,In_331);
or U986 (N_986,In_1278,In_1682);
xor U987 (N_987,In_735,In_506);
or U988 (N_988,In_2447,In_910);
or U989 (N_989,In_2550,In_839);
or U990 (N_990,In_2400,In_65);
and U991 (N_991,In_463,In_1240);
or U992 (N_992,In_546,In_55);
nand U993 (N_993,In_1157,In_1470);
and U994 (N_994,In_2131,In_2638);
nand U995 (N_995,In_1747,In_1355);
xnor U996 (N_996,In_2384,In_198);
and U997 (N_997,In_2153,In_53);
xor U998 (N_998,In_761,In_2100);
nor U999 (N_999,In_474,In_1593);
and U1000 (N_1000,In_1330,In_1823);
and U1001 (N_1001,In_2725,In_2648);
nor U1002 (N_1002,In_2052,In_513);
nor U1003 (N_1003,In_2483,In_717);
and U1004 (N_1004,In_1930,In_2829);
nand U1005 (N_1005,In_1786,In_444);
nand U1006 (N_1006,In_496,In_989);
and U1007 (N_1007,In_1186,In_929);
nand U1008 (N_1008,In_1180,In_1782);
nor U1009 (N_1009,In_2171,In_2675);
nor U1010 (N_1010,In_2973,In_1910);
or U1011 (N_1011,In_1547,In_2479);
or U1012 (N_1012,In_845,In_917);
nor U1013 (N_1013,In_1893,In_1455);
or U1014 (N_1014,In_441,In_95);
and U1015 (N_1015,In_2241,In_847);
and U1016 (N_1016,In_2574,In_1776);
nor U1017 (N_1017,In_2811,In_2727);
and U1018 (N_1018,In_2355,In_499);
and U1019 (N_1019,In_2050,In_580);
or U1020 (N_1020,In_2903,In_817);
or U1021 (N_1021,In_2065,In_1248);
or U1022 (N_1022,In_1500,In_1374);
nand U1023 (N_1023,In_877,In_2545);
and U1024 (N_1024,In_1397,In_2137);
or U1025 (N_1025,In_522,In_67);
nand U1026 (N_1026,In_656,In_222);
or U1027 (N_1027,In_769,In_355);
nand U1028 (N_1028,In_1012,In_1238);
nor U1029 (N_1029,In_2024,In_2222);
nor U1030 (N_1030,In_453,In_1769);
nand U1031 (N_1031,In_1049,In_1155);
or U1032 (N_1032,In_1514,In_2473);
xor U1033 (N_1033,In_470,In_584);
nand U1034 (N_1034,In_2458,In_1411);
or U1035 (N_1035,In_2040,In_1899);
xnor U1036 (N_1036,In_290,In_791);
nand U1037 (N_1037,In_2032,In_2084);
or U1038 (N_1038,In_1260,In_1115);
or U1039 (N_1039,In_1475,In_501);
nor U1040 (N_1040,In_2561,In_578);
and U1041 (N_1041,In_2807,In_749);
and U1042 (N_1042,In_1766,In_1364);
nor U1043 (N_1043,In_2881,In_2704);
nand U1044 (N_1044,In_1003,In_743);
nor U1045 (N_1045,In_1333,In_1988);
nand U1046 (N_1046,In_257,In_1265);
or U1047 (N_1047,In_1701,In_127);
or U1048 (N_1048,In_354,In_402);
nand U1049 (N_1049,In_1359,In_1414);
nand U1050 (N_1050,In_2566,In_2839);
and U1051 (N_1051,In_939,In_383);
or U1052 (N_1052,In_2967,In_2326);
nor U1053 (N_1053,In_1805,In_33);
nand U1054 (N_1054,In_885,In_1293);
nand U1055 (N_1055,In_718,In_269);
or U1056 (N_1056,In_1843,In_1473);
nand U1057 (N_1057,In_437,In_2011);
and U1058 (N_1058,In_600,In_1523);
and U1059 (N_1059,In_2194,In_1961);
nor U1060 (N_1060,In_1546,In_1504);
and U1061 (N_1061,In_859,In_168);
xnor U1062 (N_1062,In_1808,In_2994);
and U1063 (N_1063,In_1122,In_274);
nand U1064 (N_1064,In_1801,In_1511);
or U1065 (N_1065,In_139,In_2016);
nand U1066 (N_1066,In_805,In_1653);
nor U1067 (N_1067,In_173,In_702);
and U1068 (N_1068,In_2677,In_703);
and U1069 (N_1069,In_1189,In_460);
xnor U1070 (N_1070,In_1736,In_1133);
nor U1071 (N_1071,In_677,In_1358);
or U1072 (N_1072,In_1553,In_2081);
and U1073 (N_1073,In_1209,In_1870);
or U1074 (N_1074,In_2767,In_323);
or U1075 (N_1075,In_2960,In_1792);
nand U1076 (N_1076,In_661,In_169);
or U1077 (N_1077,In_2509,In_2735);
nor U1078 (N_1078,In_1991,In_1775);
and U1079 (N_1079,In_2553,In_447);
and U1080 (N_1080,In_2071,In_301);
nand U1081 (N_1081,In_1655,In_1150);
nand U1082 (N_1082,In_1436,In_787);
or U1083 (N_1083,In_1125,In_2951);
nand U1084 (N_1084,In_2711,In_2969);
and U1085 (N_1085,In_2551,In_328);
or U1086 (N_1086,In_2394,In_619);
xor U1087 (N_1087,In_690,In_1466);
and U1088 (N_1088,In_2852,In_1377);
nor U1089 (N_1089,In_280,In_907);
or U1090 (N_1090,In_2877,In_1834);
nand U1091 (N_1091,In_1845,In_1724);
nand U1092 (N_1092,In_1897,In_1657);
nand U1093 (N_1093,In_1274,In_1689);
or U1094 (N_1094,In_988,In_1699);
or U1095 (N_1095,In_525,In_2922);
nor U1096 (N_1096,In_2529,In_2127);
nand U1097 (N_1097,In_949,In_1584);
nor U1098 (N_1098,In_1852,In_249);
or U1099 (N_1099,In_974,In_2658);
nor U1100 (N_1100,In_1091,In_171);
and U1101 (N_1101,In_2864,In_524);
and U1102 (N_1102,In_2182,In_221);
nor U1103 (N_1103,In_398,In_2453);
or U1104 (N_1104,In_2104,In_1611);
and U1105 (N_1105,In_2757,In_1886);
or U1106 (N_1106,In_905,In_2300);
or U1107 (N_1107,In_2003,In_1678);
xor U1108 (N_1108,In_963,In_2452);
or U1109 (N_1109,In_93,In_2577);
or U1110 (N_1110,In_1383,In_533);
nor U1111 (N_1111,In_2991,In_676);
nand U1112 (N_1112,In_1298,In_2976);
xnor U1113 (N_1113,In_431,In_586);
nor U1114 (N_1114,In_2457,In_333);
or U1115 (N_1115,In_870,In_1007);
or U1116 (N_1116,In_1894,In_2419);
and U1117 (N_1117,In_1680,In_2633);
nand U1118 (N_1118,In_570,In_4);
nor U1119 (N_1119,In_535,In_681);
nor U1120 (N_1120,In_2826,In_1855);
nor U1121 (N_1121,In_2495,In_1596);
nand U1122 (N_1122,In_2004,In_2578);
or U1123 (N_1123,In_2209,In_1493);
and U1124 (N_1124,In_1824,In_25);
and U1125 (N_1125,In_972,In_434);
nand U1126 (N_1126,In_1199,In_2530);
and U1127 (N_1127,In_2703,In_1285);
nand U1128 (N_1128,In_2291,In_2214);
and U1129 (N_1129,In_694,In_2630);
nand U1130 (N_1130,In_2609,In_576);
and U1131 (N_1131,In_2800,In_1796);
nand U1132 (N_1132,In_2210,In_2997);
nand U1133 (N_1133,In_2558,In_942);
and U1134 (N_1134,In_190,In_2158);
nor U1135 (N_1135,In_776,In_1651);
nor U1136 (N_1136,In_1902,In_825);
nor U1137 (N_1137,In_1317,In_1524);
or U1138 (N_1138,In_2590,In_854);
nor U1139 (N_1139,In_799,In_2366);
xor U1140 (N_1140,In_1803,In_1840);
nor U1141 (N_1141,In_1525,In_2418);
xnor U1142 (N_1142,In_1644,In_657);
xor U1143 (N_1143,In_2567,In_2622);
xor U1144 (N_1144,In_1875,In_2470);
nand U1145 (N_1145,In_19,In_2778);
and U1146 (N_1146,In_2438,In_2425);
xor U1147 (N_1147,In_1825,In_202);
nand U1148 (N_1148,In_637,In_1979);
nand U1149 (N_1149,In_418,In_2196);
nor U1150 (N_1150,In_2323,In_399);
xor U1151 (N_1151,In_2569,In_1789);
nand U1152 (N_1152,In_1985,In_1799);
or U1153 (N_1153,In_1565,In_2875);
nand U1154 (N_1154,In_2992,In_318);
and U1155 (N_1155,In_207,In_1535);
nor U1156 (N_1156,In_828,In_613);
nor U1157 (N_1157,In_2266,In_282);
xnor U1158 (N_1158,In_747,In_362);
xor U1159 (N_1159,In_458,In_2942);
nor U1160 (N_1160,In_572,In_2815);
nand U1161 (N_1161,In_2385,In_773);
nor U1162 (N_1162,In_1937,In_2685);
nor U1163 (N_1163,In_549,In_916);
nand U1164 (N_1164,In_604,In_1262);
and U1165 (N_1165,In_1420,In_264);
or U1166 (N_1166,In_456,In_2797);
nor U1167 (N_1167,In_2516,In_2155);
or U1168 (N_1168,In_1627,In_739);
xor U1169 (N_1169,In_1388,In_1982);
nor U1170 (N_1170,In_683,In_1367);
nand U1171 (N_1171,In_15,In_1921);
or U1172 (N_1172,In_341,In_2840);
nor U1173 (N_1173,In_2576,In_1806);
or U1174 (N_1174,In_2282,In_2874);
or U1175 (N_1175,In_1867,In_262);
or U1176 (N_1176,In_2215,In_563);
nor U1177 (N_1177,In_631,In_2563);
or U1178 (N_1178,In_806,In_2916);
nor U1179 (N_1179,In_1947,In_2198);
nand U1180 (N_1180,In_166,In_2925);
xor U1181 (N_1181,In_109,In_933);
and U1182 (N_1182,In_1739,In_1862);
xnor U1183 (N_1183,In_1084,In_2895);
or U1184 (N_1184,In_99,In_2147);
nand U1185 (N_1185,In_2939,In_547);
or U1186 (N_1186,In_671,In_2793);
and U1187 (N_1187,In_1591,In_163);
nor U1188 (N_1188,In_554,In_696);
or U1189 (N_1189,In_2972,In_1195);
or U1190 (N_1190,In_130,In_1432);
and U1191 (N_1191,In_2365,In_2888);
nor U1192 (N_1192,In_893,In_272);
nand U1193 (N_1193,In_2682,In_937);
and U1194 (N_1194,In_1742,In_10);
or U1195 (N_1195,In_2620,In_2114);
or U1196 (N_1196,In_2694,In_652);
or U1197 (N_1197,In_1810,In_2849);
or U1198 (N_1198,In_587,In_2405);
nor U1199 (N_1199,In_1291,In_1934);
xor U1200 (N_1200,In_2619,In_1083);
nand U1201 (N_1201,In_1666,In_1288);
and U1202 (N_1202,In_716,In_285);
and U1203 (N_1203,In_1231,In_361);
or U1204 (N_1204,In_705,In_204);
or U1205 (N_1205,In_771,In_1172);
and U1206 (N_1206,In_1925,In_473);
and U1207 (N_1207,In_821,In_88);
or U1208 (N_1208,In_2698,In_2701);
nand U1209 (N_1209,In_1503,In_1768);
nand U1210 (N_1210,In_2721,In_2288);
and U1211 (N_1211,In_1505,In_1992);
or U1212 (N_1212,In_1754,In_2760);
nor U1213 (N_1213,In_778,In_1166);
xor U1214 (N_1214,In_1474,In_1813);
or U1215 (N_1215,In_337,In_790);
or U1216 (N_1216,In_550,In_1878);
and U1217 (N_1217,In_1908,In_2970);
and U1218 (N_1218,In_2169,In_516);
xor U1219 (N_1219,In_445,In_2074);
nor U1220 (N_1220,In_1541,In_1906);
nand U1221 (N_1221,In_1943,In_2487);
and U1222 (N_1222,In_186,In_2046);
or U1223 (N_1223,In_2720,In_795);
nor U1224 (N_1224,In_1107,In_442);
or U1225 (N_1225,In_2869,In_1642);
nor U1226 (N_1226,In_574,In_1983);
and U1227 (N_1227,In_2327,In_2544);
or U1228 (N_1228,In_1219,In_1143);
nor U1229 (N_1229,In_2528,In_2543);
nand U1230 (N_1230,In_2788,In_2560);
and U1231 (N_1231,In_326,In_2010);
nand U1232 (N_1232,In_132,In_231);
and U1233 (N_1233,In_1663,In_430);
nor U1234 (N_1234,In_107,In_1877);
xor U1235 (N_1235,In_2414,In_1882);
nand U1236 (N_1236,In_2782,In_542);
nand U1237 (N_1237,In_2468,In_1837);
nor U1238 (N_1238,In_595,In_2998);
nand U1239 (N_1239,In_1351,In_2913);
or U1240 (N_1240,In_653,In_1936);
nor U1241 (N_1241,In_2208,In_2212);
nor U1242 (N_1242,In_2201,In_336);
or U1243 (N_1243,In_2747,In_2067);
or U1244 (N_1244,In_1354,In_2472);
and U1245 (N_1245,In_2862,In_2928);
nor U1246 (N_1246,In_2816,In_2510);
nor U1247 (N_1247,In_844,In_1785);
or U1248 (N_1248,In_1234,In_428);
and U1249 (N_1249,In_2844,In_177);
and U1250 (N_1250,In_455,In_2835);
xnor U1251 (N_1251,In_2885,In_2988);
or U1252 (N_1252,In_527,In_860);
nand U1253 (N_1253,In_415,In_710);
and U1254 (N_1254,In_1608,In_1721);
and U1255 (N_1255,In_648,In_2684);
xor U1256 (N_1256,In_1079,In_523);
xnor U1257 (N_1257,In_245,In_2243);
and U1258 (N_1258,In_1257,In_82);
nand U1259 (N_1259,In_2187,In_97);
nand U1260 (N_1260,In_1398,In_56);
nor U1261 (N_1261,In_504,In_667);
nand U1262 (N_1262,In_987,In_1938);
nand U1263 (N_1263,In_70,In_2798);
or U1264 (N_1264,In_1128,In_2488);
and U1265 (N_1265,In_618,In_2014);
or U1266 (N_1266,In_100,In_2828);
nor U1267 (N_1267,In_1287,In_2306);
nand U1268 (N_1268,In_1592,In_2549);
xor U1269 (N_1269,In_2836,In_2755);
and U1270 (N_1270,In_224,In_1712);
nor U1271 (N_1271,In_2571,In_1681);
and U1272 (N_1272,In_2709,In_1780);
nor U1273 (N_1273,In_722,In_1464);
and U1274 (N_1274,In_1400,In_1135);
and U1275 (N_1275,In_407,In_1381);
nor U1276 (N_1276,In_689,In_1073);
and U1277 (N_1277,In_495,In_2092);
nor U1278 (N_1278,In_1198,In_2688);
and U1279 (N_1279,In_588,In_98);
and U1280 (N_1280,In_1639,In_1741);
and U1281 (N_1281,In_767,In_1781);
nand U1282 (N_1282,In_2444,In_2041);
nand U1283 (N_1283,In_1253,In_76);
nand U1284 (N_1284,In_2637,In_2673);
or U1285 (N_1285,In_472,In_2792);
nor U1286 (N_1286,In_1311,In_2783);
or U1287 (N_1287,In_2921,In_820);
and U1288 (N_1288,In_2805,In_13);
or U1289 (N_1289,In_372,In_1149);
nor U1290 (N_1290,In_2009,In_2906);
nand U1291 (N_1291,In_2197,In_1129);
nand U1292 (N_1292,In_1907,In_1794);
or U1293 (N_1293,In_2054,In_843);
nor U1294 (N_1294,In_2224,In_1040);
nand U1295 (N_1295,In_37,In_1386);
nand U1296 (N_1296,In_2021,In_639);
or U1297 (N_1297,In_853,In_1227);
or U1298 (N_1298,In_234,In_2585);
and U1299 (N_1299,In_2265,In_1561);
or U1300 (N_1300,In_1960,In_1588);
or U1301 (N_1301,In_1549,In_1214);
and U1302 (N_1302,In_225,In_197);
xor U1303 (N_1303,In_1731,In_302);
nand U1304 (N_1304,In_2061,In_2751);
nor U1305 (N_1305,In_1251,In_322);
and U1306 (N_1306,In_2191,In_1065);
nor U1307 (N_1307,In_1465,In_678);
and U1308 (N_1308,In_1649,In_205);
and U1309 (N_1309,In_1056,In_2485);
or U1310 (N_1310,In_239,In_451);
xnor U1311 (N_1311,In_2085,In_512);
nor U1312 (N_1312,In_2946,In_940);
or U1313 (N_1313,In_935,In_529);
nand U1314 (N_1314,In_23,In_2226);
or U1315 (N_1315,In_2953,In_241);
and U1316 (N_1316,In_2422,In_983);
nand U1317 (N_1317,In_2657,In_1302);
nor U1318 (N_1318,In_1315,In_1967);
or U1319 (N_1319,In_2848,In_424);
nand U1320 (N_1320,In_1812,In_617);
nand U1321 (N_1321,In_47,In_2144);
nor U1322 (N_1322,In_493,In_1444);
nand U1323 (N_1323,In_561,In_1756);
nand U1324 (N_1324,In_1879,In_164);
or U1325 (N_1325,In_1580,In_612);
or U1326 (N_1326,In_2072,In_1725);
xnor U1327 (N_1327,In_2920,In_659);
nor U1328 (N_1328,In_2989,In_757);
nand U1329 (N_1329,In_579,In_649);
nor U1330 (N_1330,In_2672,In_1576);
or U1331 (N_1331,In_1928,In_1316);
nor U1332 (N_1332,In_1744,In_2120);
nor U1333 (N_1333,In_594,In_1452);
and U1334 (N_1334,In_566,In_756);
and U1335 (N_1335,In_1520,In_2403);
nor U1336 (N_1336,In_1162,In_1563);
and U1337 (N_1337,In_2659,In_28);
nand U1338 (N_1338,In_2818,In_2023);
nand U1339 (N_1339,In_2193,In_2276);
nand U1340 (N_1340,In_1461,In_2268);
nor U1341 (N_1341,In_660,In_2601);
nand U1342 (N_1342,In_2871,In_1700);
or U1343 (N_1343,In_320,In_1403);
or U1344 (N_1344,In_557,In_2730);
xnor U1345 (N_1345,In_2734,In_316);
xnor U1346 (N_1346,In_1518,In_1685);
and U1347 (N_1347,In_116,In_1245);
nand U1348 (N_1348,In_170,In_2019);
nand U1349 (N_1349,In_187,In_982);
nor U1350 (N_1350,In_2467,In_1387);
and U1351 (N_1351,In_2141,In_2044);
xor U1352 (N_1352,In_1208,In_1277);
nand U1353 (N_1353,In_1973,In_1165);
and U1354 (N_1354,In_1959,In_774);
or U1355 (N_1355,In_1501,In_2785);
nand U1356 (N_1356,In_2039,In_1955);
and U1357 (N_1357,In_14,In_1861);
nor U1358 (N_1358,In_952,In_2527);
nand U1359 (N_1359,In_2712,In_2217);
nor U1360 (N_1360,In_927,In_2937);
nand U1361 (N_1361,In_1081,In_1521);
nor U1362 (N_1362,In_665,In_1997);
nor U1363 (N_1363,In_1931,In_567);
nand U1364 (N_1364,In_140,In_385);
and U1365 (N_1365,In_2506,In_2451);
nor U1366 (N_1366,In_1456,In_873);
and U1367 (N_1367,In_158,In_392);
nor U1368 (N_1368,In_2399,In_2346);
and U1369 (N_1369,In_2377,In_908);
xor U1370 (N_1370,In_1353,In_90);
or U1371 (N_1371,In_2128,In_1846);
nor U1372 (N_1372,In_1519,In_1571);
nand U1373 (N_1373,In_1156,In_1788);
xor U1374 (N_1374,In_389,In_452);
nor U1375 (N_1375,In_936,In_375);
and U1376 (N_1376,In_2091,In_113);
nand U1377 (N_1377,In_2752,In_2643);
or U1378 (N_1378,In_1038,In_607);
or U1379 (N_1379,In_367,In_1478);
or U1380 (N_1380,In_1819,In_2722);
xnor U1381 (N_1381,In_700,In_1249);
xnor U1382 (N_1382,In_41,In_1235);
or U1383 (N_1383,In_1940,In_970);
nand U1384 (N_1384,In_2476,In_553);
nor U1385 (N_1385,In_2809,In_610);
or U1386 (N_1386,In_1202,In_133);
or U1387 (N_1387,In_1082,In_1980);
nand U1388 (N_1388,In_956,In_1113);
or U1389 (N_1389,In_2203,In_1119);
nand U1390 (N_1390,In_1777,In_228);
nand U1391 (N_1391,In_1075,In_1847);
or U1392 (N_1392,In_2170,In_1106);
and U1393 (N_1393,In_2984,In_217);
or U1394 (N_1394,In_1574,In_2842);
or U1395 (N_1395,In_1898,In_1338);
nor U1396 (N_1396,In_261,In_2232);
nor U1397 (N_1397,In_440,In_1784);
and U1398 (N_1398,In_879,In_1479);
nand U1399 (N_1399,In_21,In_2511);
or U1400 (N_1400,In_1981,In_2813);
and U1401 (N_1401,In_1438,In_1617);
nand U1402 (N_1402,In_2140,In_1693);
nor U1403 (N_1403,In_960,In_1632);
or U1404 (N_1404,In_666,In_1349);
nor U1405 (N_1405,In_1652,In_1732);
and U1406 (N_1406,In_2905,In_2246);
or U1407 (N_1407,In_1552,In_900);
nand U1408 (N_1408,In_2428,In_708);
nor U1409 (N_1409,In_240,In_1190);
nor U1410 (N_1410,In_1687,In_1365);
nor U1411 (N_1411,In_1224,In_2057);
or U1412 (N_1412,In_1548,In_446);
nor U1413 (N_1413,In_2499,In_83);
nand U1414 (N_1414,In_714,In_1170);
and U1415 (N_1415,In_2931,In_2533);
nor U1416 (N_1416,In_1858,In_622);
nand U1417 (N_1417,In_2766,In_1323);
nand U1418 (N_1418,In_758,In_2819);
xnor U1419 (N_1419,In_1762,In_969);
or U1420 (N_1420,In_423,In_2859);
xnor U1421 (N_1421,In_1895,In_789);
nand U1422 (N_1422,In_2218,In_2383);
nand U1423 (N_1423,In_2702,In_1123);
or U1424 (N_1424,In_2891,In_327);
nand U1425 (N_1425,In_1838,In_762);
and U1426 (N_1426,In_794,In_2492);
nand U1427 (N_1427,In_2139,In_2831);
xnor U1428 (N_1428,In_2370,In_1051);
and U1429 (N_1429,In_126,In_2603);
and U1430 (N_1430,In_1321,In_2254);
nor U1431 (N_1431,In_2427,In_740);
or U1432 (N_1432,In_1197,In_1446);
and U1433 (N_1433,In_1102,In_2038);
nand U1434 (N_1434,In_1560,In_1482);
and U1435 (N_1435,In_959,In_2388);
nand U1436 (N_1436,In_2713,In_2926);
or U1437 (N_1437,In_835,In_335);
nor U1438 (N_1438,In_2823,In_1771);
or U1439 (N_1439,In_801,In_117);
nand U1440 (N_1440,In_325,In_2789);
xor U1441 (N_1441,In_1508,In_2093);
or U1442 (N_1442,In_2172,In_357);
nand U1443 (N_1443,In_321,In_1641);
and U1444 (N_1444,In_1990,In_1569);
nor U1445 (N_1445,In_732,In_883);
nor U1446 (N_1446,In_2697,In_763);
nor U1447 (N_1447,In_1818,In_1833);
nor U1448 (N_1448,In_1299,In_2077);
and U1449 (N_1449,In_2379,In_62);
or U1450 (N_1450,In_2344,In_615);
nand U1451 (N_1451,In_2833,In_478);
or U1452 (N_1452,In_2546,In_1974);
or U1453 (N_1453,In_1880,In_344);
nand U1454 (N_1454,In_2723,In_1558);
and U1455 (N_1455,In_1193,In_2748);
or U1456 (N_1456,In_2908,In_1963);
or U1457 (N_1457,In_73,In_2978);
nor U1458 (N_1458,In_2219,In_1309);
or U1459 (N_1459,In_31,In_370);
nand U1460 (N_1460,In_382,In_2565);
nor U1461 (N_1461,In_2163,In_2843);
nand U1462 (N_1462,In_593,In_360);
nand U1463 (N_1463,In_2892,In_298);
nor U1464 (N_1464,In_2935,In_199);
xor U1465 (N_1465,In_1692,In_981);
and U1466 (N_1466,In_1070,In_18);
nor U1467 (N_1467,In_1292,In_244);
and U1468 (N_1468,In_2640,In_2652);
nor U1469 (N_1469,In_2145,In_457);
and U1470 (N_1470,In_46,In_1332);
nand U1471 (N_1471,In_2393,In_432);
and U1472 (N_1472,In_2000,In_1489);
nand U1473 (N_1473,In_45,In_1220);
and U1474 (N_1474,In_1105,In_2999);
nand U1475 (N_1475,In_724,In_753);
xnor U1476 (N_1476,In_1163,In_1883);
nor U1477 (N_1477,In_1345,In_9);
nor U1478 (N_1478,In_1213,In_2936);
and U1479 (N_1479,In_1749,In_564);
and U1480 (N_1480,In_1965,In_1206);
or U1481 (N_1481,In_1246,In_246);
nand U1482 (N_1482,In_2312,In_1061);
xnor U1483 (N_1483,In_2732,In_2514);
and U1484 (N_1484,In_1016,In_1526);
nor U1485 (N_1485,In_1448,In_176);
and U1486 (N_1486,In_2015,In_2756);
or U1487 (N_1487,In_1431,In_2058);
and U1488 (N_1488,In_1946,In_1587);
nand U1489 (N_1489,In_1953,In_1610);
nand U1490 (N_1490,In_950,In_2332);
nor U1491 (N_1491,In_1850,In_1892);
xor U1492 (N_1492,In_1942,In_378);
nand U1493 (N_1493,In_510,In_2650);
and U1494 (N_1494,In_1829,In_1969);
nor U1495 (N_1495,In_971,In_993);
or U1496 (N_1496,In_632,In_2856);
and U1497 (N_1497,In_1319,In_532);
nor U1498 (N_1498,In_867,In_2627);
or U1499 (N_1499,In_1839,In_560);
and U1500 (N_1500,In_759,In_2673);
nor U1501 (N_1501,In_2476,In_2185);
and U1502 (N_1502,In_720,In_1875);
xnor U1503 (N_1503,In_947,In_2356);
nor U1504 (N_1504,In_2045,In_2834);
and U1505 (N_1505,In_2562,In_213);
and U1506 (N_1506,In_2110,In_2473);
or U1507 (N_1507,In_891,In_1642);
nor U1508 (N_1508,In_2748,In_2524);
nand U1509 (N_1509,In_2531,In_640);
nand U1510 (N_1510,In_870,In_2865);
nand U1511 (N_1511,In_1392,In_916);
and U1512 (N_1512,In_1152,In_1899);
nand U1513 (N_1513,In_2901,In_1197);
nand U1514 (N_1514,In_2389,In_210);
or U1515 (N_1515,In_1489,In_2713);
or U1516 (N_1516,In_2740,In_1133);
nand U1517 (N_1517,In_1638,In_2569);
and U1518 (N_1518,In_749,In_942);
and U1519 (N_1519,In_2956,In_2260);
xor U1520 (N_1520,In_1946,In_2875);
and U1521 (N_1521,In_2093,In_824);
xor U1522 (N_1522,In_2197,In_220);
xnor U1523 (N_1523,In_114,In_1150);
and U1524 (N_1524,In_10,In_2602);
or U1525 (N_1525,In_2046,In_472);
nand U1526 (N_1526,In_1038,In_2457);
and U1527 (N_1527,In_609,In_2930);
nor U1528 (N_1528,In_1552,In_2655);
nor U1529 (N_1529,In_2127,In_2573);
and U1530 (N_1530,In_883,In_2563);
nand U1531 (N_1531,In_2611,In_1102);
or U1532 (N_1532,In_1065,In_1989);
and U1533 (N_1533,In_434,In_2572);
and U1534 (N_1534,In_1118,In_1670);
or U1535 (N_1535,In_1096,In_792);
nor U1536 (N_1536,In_2856,In_1355);
nand U1537 (N_1537,In_244,In_2199);
nor U1538 (N_1538,In_1354,In_198);
or U1539 (N_1539,In_2898,In_1488);
nor U1540 (N_1540,In_1979,In_1259);
xnor U1541 (N_1541,In_1877,In_1314);
or U1542 (N_1542,In_1885,In_2441);
nor U1543 (N_1543,In_2135,In_2895);
and U1544 (N_1544,In_570,In_970);
nor U1545 (N_1545,In_2593,In_1725);
xor U1546 (N_1546,In_2911,In_2344);
nor U1547 (N_1547,In_2948,In_370);
nand U1548 (N_1548,In_355,In_1290);
xnor U1549 (N_1549,In_2385,In_1485);
and U1550 (N_1550,In_2476,In_48);
nand U1551 (N_1551,In_2824,In_1102);
nor U1552 (N_1552,In_2270,In_1188);
nor U1553 (N_1553,In_2530,In_1230);
and U1554 (N_1554,In_575,In_1773);
xor U1555 (N_1555,In_1040,In_241);
nand U1556 (N_1556,In_1577,In_2788);
and U1557 (N_1557,In_2105,In_2009);
or U1558 (N_1558,In_2546,In_1221);
or U1559 (N_1559,In_255,In_671);
nor U1560 (N_1560,In_1804,In_2976);
nand U1561 (N_1561,In_2801,In_1452);
or U1562 (N_1562,In_2659,In_808);
or U1563 (N_1563,In_1097,In_1791);
xnor U1564 (N_1564,In_983,In_1419);
nand U1565 (N_1565,In_1194,In_2280);
xnor U1566 (N_1566,In_209,In_2127);
nor U1567 (N_1567,In_2933,In_1277);
xnor U1568 (N_1568,In_2538,In_379);
and U1569 (N_1569,In_141,In_1848);
and U1570 (N_1570,In_2492,In_2822);
and U1571 (N_1571,In_2819,In_2653);
xor U1572 (N_1572,In_1661,In_1138);
or U1573 (N_1573,In_2876,In_173);
xnor U1574 (N_1574,In_86,In_1384);
or U1575 (N_1575,In_1939,In_362);
or U1576 (N_1576,In_1911,In_2179);
or U1577 (N_1577,In_2045,In_850);
and U1578 (N_1578,In_1740,In_1288);
or U1579 (N_1579,In_1399,In_2102);
nor U1580 (N_1580,In_2202,In_1019);
or U1581 (N_1581,In_525,In_1036);
nand U1582 (N_1582,In_1560,In_235);
nor U1583 (N_1583,In_2836,In_1793);
xnor U1584 (N_1584,In_2335,In_496);
xor U1585 (N_1585,In_879,In_2783);
nand U1586 (N_1586,In_289,In_1431);
and U1587 (N_1587,In_1471,In_2355);
xnor U1588 (N_1588,In_2990,In_2016);
and U1589 (N_1589,In_1106,In_1048);
and U1590 (N_1590,In_2758,In_629);
nand U1591 (N_1591,In_2830,In_2147);
nor U1592 (N_1592,In_2864,In_1558);
nor U1593 (N_1593,In_1018,In_146);
and U1594 (N_1594,In_2033,In_1320);
nor U1595 (N_1595,In_885,In_1299);
or U1596 (N_1596,In_2393,In_2731);
nor U1597 (N_1597,In_1648,In_2536);
and U1598 (N_1598,In_9,In_1423);
and U1599 (N_1599,In_2156,In_2524);
or U1600 (N_1600,In_627,In_2776);
nor U1601 (N_1601,In_972,In_1164);
nand U1602 (N_1602,In_2691,In_2055);
nor U1603 (N_1603,In_1642,In_2921);
and U1604 (N_1604,In_403,In_2591);
or U1605 (N_1605,In_1816,In_1531);
nor U1606 (N_1606,In_227,In_2022);
nor U1607 (N_1607,In_2409,In_2250);
nand U1608 (N_1608,In_994,In_1703);
nor U1609 (N_1609,In_2710,In_1327);
nor U1610 (N_1610,In_598,In_1612);
nor U1611 (N_1611,In_1231,In_1844);
or U1612 (N_1612,In_2257,In_2035);
and U1613 (N_1613,In_2934,In_2049);
and U1614 (N_1614,In_316,In_2593);
xor U1615 (N_1615,In_59,In_1993);
nand U1616 (N_1616,In_1212,In_124);
xor U1617 (N_1617,In_404,In_1624);
nand U1618 (N_1618,In_1959,In_855);
or U1619 (N_1619,In_2464,In_1033);
nor U1620 (N_1620,In_2400,In_893);
nor U1621 (N_1621,In_2615,In_438);
xor U1622 (N_1622,In_14,In_2828);
nand U1623 (N_1623,In_487,In_159);
nor U1624 (N_1624,In_361,In_2149);
nor U1625 (N_1625,In_2958,In_969);
and U1626 (N_1626,In_989,In_1723);
and U1627 (N_1627,In_1527,In_1588);
nand U1628 (N_1628,In_991,In_1495);
or U1629 (N_1629,In_1050,In_2369);
or U1630 (N_1630,In_1987,In_2436);
or U1631 (N_1631,In_2202,In_426);
nand U1632 (N_1632,In_878,In_2878);
nand U1633 (N_1633,In_842,In_284);
and U1634 (N_1634,In_700,In_888);
nor U1635 (N_1635,In_2004,In_860);
or U1636 (N_1636,In_1867,In_2476);
or U1637 (N_1637,In_1790,In_1741);
and U1638 (N_1638,In_1263,In_2554);
xnor U1639 (N_1639,In_1382,In_1176);
nand U1640 (N_1640,In_1693,In_2930);
nor U1641 (N_1641,In_2014,In_1958);
nand U1642 (N_1642,In_866,In_1026);
or U1643 (N_1643,In_2628,In_2120);
nor U1644 (N_1644,In_63,In_121);
nor U1645 (N_1645,In_721,In_2941);
xnor U1646 (N_1646,In_1092,In_1912);
xnor U1647 (N_1647,In_2720,In_2330);
and U1648 (N_1648,In_219,In_1768);
and U1649 (N_1649,In_35,In_1213);
or U1650 (N_1650,In_299,In_1958);
nor U1651 (N_1651,In_2790,In_265);
nor U1652 (N_1652,In_848,In_248);
nor U1653 (N_1653,In_657,In_2492);
and U1654 (N_1654,In_476,In_1022);
or U1655 (N_1655,In_2228,In_455);
and U1656 (N_1656,In_138,In_1051);
and U1657 (N_1657,In_2589,In_2970);
or U1658 (N_1658,In_1344,In_2231);
nand U1659 (N_1659,In_2891,In_1882);
or U1660 (N_1660,In_962,In_1718);
or U1661 (N_1661,In_2680,In_2018);
and U1662 (N_1662,In_1133,In_79);
nand U1663 (N_1663,In_2415,In_2770);
or U1664 (N_1664,In_1175,In_2038);
xnor U1665 (N_1665,In_2435,In_2404);
nand U1666 (N_1666,In_1950,In_893);
nor U1667 (N_1667,In_216,In_1725);
nand U1668 (N_1668,In_798,In_2230);
and U1669 (N_1669,In_313,In_2958);
nand U1670 (N_1670,In_1771,In_2883);
xor U1671 (N_1671,In_1501,In_1403);
nor U1672 (N_1672,In_630,In_1458);
nand U1673 (N_1673,In_1836,In_2540);
or U1674 (N_1674,In_1233,In_1390);
nand U1675 (N_1675,In_1533,In_1661);
nor U1676 (N_1676,In_446,In_228);
or U1677 (N_1677,In_2512,In_725);
nor U1678 (N_1678,In_2304,In_1896);
xnor U1679 (N_1679,In_2054,In_2974);
nand U1680 (N_1680,In_1715,In_480);
and U1681 (N_1681,In_908,In_2718);
nor U1682 (N_1682,In_1410,In_447);
xor U1683 (N_1683,In_163,In_2309);
or U1684 (N_1684,In_11,In_257);
nor U1685 (N_1685,In_42,In_179);
or U1686 (N_1686,In_2745,In_2369);
and U1687 (N_1687,In_2733,In_2289);
nor U1688 (N_1688,In_2226,In_155);
and U1689 (N_1689,In_611,In_2136);
and U1690 (N_1690,In_1178,In_1900);
nor U1691 (N_1691,In_1179,In_269);
nor U1692 (N_1692,In_2095,In_122);
and U1693 (N_1693,In_909,In_952);
nand U1694 (N_1694,In_2918,In_127);
nor U1695 (N_1695,In_1903,In_2544);
and U1696 (N_1696,In_1332,In_2429);
and U1697 (N_1697,In_2455,In_1614);
nand U1698 (N_1698,In_1050,In_294);
and U1699 (N_1699,In_64,In_888);
and U1700 (N_1700,In_466,In_619);
or U1701 (N_1701,In_2329,In_1098);
or U1702 (N_1702,In_2305,In_811);
nor U1703 (N_1703,In_1263,In_2830);
nand U1704 (N_1704,In_2256,In_967);
and U1705 (N_1705,In_2320,In_1872);
or U1706 (N_1706,In_2404,In_1729);
nand U1707 (N_1707,In_2459,In_869);
or U1708 (N_1708,In_1081,In_805);
and U1709 (N_1709,In_1714,In_2047);
or U1710 (N_1710,In_489,In_512);
nor U1711 (N_1711,In_2608,In_2128);
or U1712 (N_1712,In_2429,In_964);
nor U1713 (N_1713,In_1966,In_2497);
nor U1714 (N_1714,In_2952,In_1578);
xor U1715 (N_1715,In_2308,In_245);
nor U1716 (N_1716,In_2970,In_2646);
or U1717 (N_1717,In_2324,In_202);
and U1718 (N_1718,In_335,In_541);
or U1719 (N_1719,In_710,In_286);
nand U1720 (N_1720,In_1911,In_1725);
and U1721 (N_1721,In_2006,In_537);
nand U1722 (N_1722,In_1108,In_848);
and U1723 (N_1723,In_1361,In_1535);
or U1724 (N_1724,In_574,In_2964);
or U1725 (N_1725,In_2352,In_91);
or U1726 (N_1726,In_51,In_2196);
nand U1727 (N_1727,In_1713,In_750);
nand U1728 (N_1728,In_785,In_1157);
nand U1729 (N_1729,In_2861,In_1185);
nor U1730 (N_1730,In_1740,In_1886);
and U1731 (N_1731,In_739,In_2143);
and U1732 (N_1732,In_72,In_2644);
nand U1733 (N_1733,In_780,In_312);
xor U1734 (N_1734,In_2159,In_1460);
or U1735 (N_1735,In_920,In_680);
and U1736 (N_1736,In_1057,In_2034);
xnor U1737 (N_1737,In_2834,In_2701);
nand U1738 (N_1738,In_144,In_2384);
xor U1739 (N_1739,In_2589,In_1332);
nor U1740 (N_1740,In_2801,In_691);
nand U1741 (N_1741,In_151,In_1618);
and U1742 (N_1742,In_1461,In_834);
and U1743 (N_1743,In_529,In_2192);
nand U1744 (N_1744,In_2862,In_1158);
or U1745 (N_1745,In_1448,In_2967);
or U1746 (N_1746,In_2580,In_1806);
or U1747 (N_1747,In_2122,In_2861);
nand U1748 (N_1748,In_345,In_1052);
and U1749 (N_1749,In_2195,In_2639);
nand U1750 (N_1750,In_2903,In_327);
nand U1751 (N_1751,In_2681,In_1397);
and U1752 (N_1752,In_1587,In_1287);
nor U1753 (N_1753,In_1790,In_1670);
and U1754 (N_1754,In_1705,In_2251);
nand U1755 (N_1755,In_1668,In_661);
nor U1756 (N_1756,In_6,In_2643);
xnor U1757 (N_1757,In_1844,In_2781);
or U1758 (N_1758,In_995,In_1104);
nor U1759 (N_1759,In_2858,In_1716);
and U1760 (N_1760,In_1142,In_1990);
nor U1761 (N_1761,In_460,In_2302);
nor U1762 (N_1762,In_1723,In_2266);
or U1763 (N_1763,In_2382,In_2644);
nor U1764 (N_1764,In_1477,In_1013);
or U1765 (N_1765,In_696,In_1442);
nand U1766 (N_1766,In_2489,In_2966);
nand U1767 (N_1767,In_2800,In_684);
and U1768 (N_1768,In_1131,In_1801);
and U1769 (N_1769,In_74,In_1123);
nand U1770 (N_1770,In_258,In_936);
nand U1771 (N_1771,In_2776,In_1805);
nand U1772 (N_1772,In_715,In_2576);
and U1773 (N_1773,In_2893,In_1446);
and U1774 (N_1774,In_1870,In_346);
nand U1775 (N_1775,In_2540,In_1701);
nor U1776 (N_1776,In_2129,In_23);
nor U1777 (N_1777,In_2255,In_648);
nor U1778 (N_1778,In_1694,In_2406);
nor U1779 (N_1779,In_377,In_533);
nand U1780 (N_1780,In_2173,In_206);
nand U1781 (N_1781,In_1010,In_1642);
and U1782 (N_1782,In_2547,In_1166);
nor U1783 (N_1783,In_1680,In_841);
and U1784 (N_1784,In_1061,In_2689);
nand U1785 (N_1785,In_366,In_389);
and U1786 (N_1786,In_638,In_1518);
nor U1787 (N_1787,In_1669,In_1781);
nor U1788 (N_1788,In_1693,In_1827);
xor U1789 (N_1789,In_333,In_2795);
nor U1790 (N_1790,In_29,In_2260);
or U1791 (N_1791,In_1350,In_101);
or U1792 (N_1792,In_866,In_2770);
or U1793 (N_1793,In_509,In_793);
and U1794 (N_1794,In_2430,In_1910);
xnor U1795 (N_1795,In_9,In_2732);
nor U1796 (N_1796,In_1854,In_145);
and U1797 (N_1797,In_1095,In_812);
nor U1798 (N_1798,In_1237,In_518);
or U1799 (N_1799,In_1397,In_1736);
nand U1800 (N_1800,In_2157,In_677);
and U1801 (N_1801,In_2931,In_1176);
or U1802 (N_1802,In_271,In_2055);
nor U1803 (N_1803,In_909,In_1794);
nand U1804 (N_1804,In_2003,In_2909);
nor U1805 (N_1805,In_2987,In_638);
and U1806 (N_1806,In_2047,In_1213);
and U1807 (N_1807,In_1771,In_754);
nand U1808 (N_1808,In_255,In_1393);
nor U1809 (N_1809,In_2570,In_1142);
nor U1810 (N_1810,In_362,In_2511);
xnor U1811 (N_1811,In_2742,In_2154);
nor U1812 (N_1812,In_1653,In_1142);
nand U1813 (N_1813,In_724,In_1634);
nor U1814 (N_1814,In_67,In_119);
and U1815 (N_1815,In_2029,In_1096);
and U1816 (N_1816,In_1100,In_1175);
nand U1817 (N_1817,In_342,In_2292);
nand U1818 (N_1818,In_545,In_279);
and U1819 (N_1819,In_315,In_2964);
nor U1820 (N_1820,In_2767,In_1161);
or U1821 (N_1821,In_1917,In_389);
or U1822 (N_1822,In_1127,In_796);
nand U1823 (N_1823,In_863,In_2341);
nand U1824 (N_1824,In_1263,In_1724);
nand U1825 (N_1825,In_588,In_2956);
or U1826 (N_1826,In_939,In_1141);
nand U1827 (N_1827,In_2972,In_493);
nor U1828 (N_1828,In_2051,In_1876);
or U1829 (N_1829,In_2652,In_486);
and U1830 (N_1830,In_799,In_1323);
or U1831 (N_1831,In_486,In_1544);
and U1832 (N_1832,In_213,In_2513);
and U1833 (N_1833,In_2747,In_2241);
or U1834 (N_1834,In_1578,In_2213);
nor U1835 (N_1835,In_2112,In_2390);
and U1836 (N_1836,In_19,In_2991);
nand U1837 (N_1837,In_2487,In_2214);
and U1838 (N_1838,In_1492,In_1204);
or U1839 (N_1839,In_1367,In_1265);
and U1840 (N_1840,In_1096,In_1666);
or U1841 (N_1841,In_108,In_2535);
and U1842 (N_1842,In_1679,In_1906);
nand U1843 (N_1843,In_669,In_1522);
or U1844 (N_1844,In_1921,In_834);
nand U1845 (N_1845,In_1225,In_1629);
nor U1846 (N_1846,In_1234,In_1323);
nor U1847 (N_1847,In_2087,In_231);
nor U1848 (N_1848,In_1897,In_1874);
nor U1849 (N_1849,In_765,In_2684);
nand U1850 (N_1850,In_2402,In_360);
or U1851 (N_1851,In_1970,In_638);
nand U1852 (N_1852,In_803,In_1674);
nand U1853 (N_1853,In_184,In_384);
and U1854 (N_1854,In_1506,In_681);
xor U1855 (N_1855,In_624,In_271);
or U1856 (N_1856,In_2225,In_1148);
nor U1857 (N_1857,In_564,In_1769);
or U1858 (N_1858,In_1219,In_2082);
and U1859 (N_1859,In_2973,In_2308);
xnor U1860 (N_1860,In_2672,In_126);
nand U1861 (N_1861,In_1062,In_2512);
nor U1862 (N_1862,In_2425,In_2513);
nor U1863 (N_1863,In_1174,In_1304);
nor U1864 (N_1864,In_1294,In_1739);
nand U1865 (N_1865,In_2212,In_2699);
or U1866 (N_1866,In_2251,In_243);
or U1867 (N_1867,In_1931,In_800);
nor U1868 (N_1868,In_2336,In_1184);
or U1869 (N_1869,In_1031,In_1920);
nor U1870 (N_1870,In_551,In_2040);
and U1871 (N_1871,In_2752,In_2592);
nand U1872 (N_1872,In_937,In_1617);
or U1873 (N_1873,In_1853,In_1697);
or U1874 (N_1874,In_2608,In_2704);
nand U1875 (N_1875,In_1914,In_1388);
xnor U1876 (N_1876,In_1457,In_2517);
nor U1877 (N_1877,In_1796,In_1490);
or U1878 (N_1878,In_2247,In_2878);
and U1879 (N_1879,In_733,In_1101);
nand U1880 (N_1880,In_2292,In_2451);
and U1881 (N_1881,In_865,In_1223);
or U1882 (N_1882,In_775,In_1558);
or U1883 (N_1883,In_930,In_1694);
nor U1884 (N_1884,In_810,In_635);
nand U1885 (N_1885,In_1477,In_855);
and U1886 (N_1886,In_382,In_1303);
and U1887 (N_1887,In_1825,In_1652);
nand U1888 (N_1888,In_1012,In_2651);
nand U1889 (N_1889,In_2323,In_1160);
nor U1890 (N_1890,In_2950,In_760);
nand U1891 (N_1891,In_1417,In_767);
or U1892 (N_1892,In_1792,In_373);
or U1893 (N_1893,In_1507,In_2274);
nand U1894 (N_1894,In_418,In_2719);
nor U1895 (N_1895,In_695,In_1418);
and U1896 (N_1896,In_397,In_1142);
nand U1897 (N_1897,In_250,In_841);
nor U1898 (N_1898,In_2589,In_496);
and U1899 (N_1899,In_435,In_1631);
and U1900 (N_1900,In_2008,In_1111);
nand U1901 (N_1901,In_836,In_437);
and U1902 (N_1902,In_696,In_526);
nand U1903 (N_1903,In_2201,In_1817);
and U1904 (N_1904,In_628,In_1753);
nor U1905 (N_1905,In_2460,In_1297);
nand U1906 (N_1906,In_1236,In_1992);
or U1907 (N_1907,In_1112,In_2955);
and U1908 (N_1908,In_1500,In_3);
or U1909 (N_1909,In_1291,In_1617);
nand U1910 (N_1910,In_834,In_2227);
nand U1911 (N_1911,In_1278,In_2906);
nand U1912 (N_1912,In_1705,In_676);
nand U1913 (N_1913,In_2105,In_2138);
and U1914 (N_1914,In_2575,In_2477);
or U1915 (N_1915,In_710,In_2696);
or U1916 (N_1916,In_2794,In_55);
nand U1917 (N_1917,In_1235,In_1983);
nor U1918 (N_1918,In_1536,In_1487);
or U1919 (N_1919,In_2851,In_1254);
or U1920 (N_1920,In_2214,In_2187);
nor U1921 (N_1921,In_2050,In_1076);
nand U1922 (N_1922,In_2742,In_1938);
nand U1923 (N_1923,In_434,In_1753);
nor U1924 (N_1924,In_479,In_1750);
xnor U1925 (N_1925,In_273,In_1302);
nor U1926 (N_1926,In_283,In_853);
nand U1927 (N_1927,In_807,In_642);
nor U1928 (N_1928,In_2430,In_1258);
nor U1929 (N_1929,In_2729,In_1905);
nand U1930 (N_1930,In_2373,In_592);
nand U1931 (N_1931,In_2520,In_1548);
nor U1932 (N_1932,In_764,In_1784);
nor U1933 (N_1933,In_473,In_382);
or U1934 (N_1934,In_1590,In_2600);
or U1935 (N_1935,In_1365,In_435);
nor U1936 (N_1936,In_566,In_1929);
and U1937 (N_1937,In_1240,In_43);
and U1938 (N_1938,In_2305,In_1577);
nand U1939 (N_1939,In_751,In_2390);
nand U1940 (N_1940,In_912,In_315);
and U1941 (N_1941,In_2927,In_2594);
and U1942 (N_1942,In_2494,In_2265);
or U1943 (N_1943,In_825,In_71);
nand U1944 (N_1944,In_1210,In_2672);
nand U1945 (N_1945,In_1888,In_932);
and U1946 (N_1946,In_2132,In_519);
nor U1947 (N_1947,In_1127,In_1814);
nand U1948 (N_1948,In_2540,In_1530);
and U1949 (N_1949,In_2766,In_1113);
or U1950 (N_1950,In_929,In_366);
and U1951 (N_1951,In_182,In_1014);
and U1952 (N_1952,In_639,In_2937);
or U1953 (N_1953,In_2256,In_1507);
and U1954 (N_1954,In_2452,In_882);
nand U1955 (N_1955,In_2158,In_1617);
nand U1956 (N_1956,In_1783,In_549);
xnor U1957 (N_1957,In_2578,In_1892);
and U1958 (N_1958,In_122,In_2159);
and U1959 (N_1959,In_835,In_666);
and U1960 (N_1960,In_677,In_1337);
nand U1961 (N_1961,In_1631,In_612);
and U1962 (N_1962,In_2656,In_199);
or U1963 (N_1963,In_709,In_2008);
or U1964 (N_1964,In_1692,In_2733);
or U1965 (N_1965,In_227,In_189);
or U1966 (N_1966,In_797,In_329);
nand U1967 (N_1967,In_176,In_2477);
nor U1968 (N_1968,In_1979,In_2473);
and U1969 (N_1969,In_259,In_2669);
and U1970 (N_1970,In_1200,In_223);
and U1971 (N_1971,In_730,In_389);
and U1972 (N_1972,In_768,In_1610);
xor U1973 (N_1973,In_316,In_2458);
or U1974 (N_1974,In_1991,In_274);
or U1975 (N_1975,In_2146,In_1470);
nand U1976 (N_1976,In_1510,In_1015);
xor U1977 (N_1977,In_2580,In_2302);
nand U1978 (N_1978,In_2380,In_2684);
nor U1979 (N_1979,In_2466,In_872);
nand U1980 (N_1980,In_1391,In_772);
xnor U1981 (N_1981,In_1098,In_1046);
and U1982 (N_1982,In_1495,In_413);
or U1983 (N_1983,In_679,In_1063);
or U1984 (N_1984,In_1068,In_2867);
or U1985 (N_1985,In_342,In_325);
xnor U1986 (N_1986,In_1676,In_276);
and U1987 (N_1987,In_457,In_243);
xnor U1988 (N_1988,In_2690,In_677);
or U1989 (N_1989,In_2637,In_1493);
nand U1990 (N_1990,In_1664,In_178);
xnor U1991 (N_1991,In_2101,In_1776);
and U1992 (N_1992,In_892,In_2502);
and U1993 (N_1993,In_1593,In_1197);
nand U1994 (N_1994,In_503,In_2848);
nand U1995 (N_1995,In_2684,In_2113);
nand U1996 (N_1996,In_59,In_511);
nand U1997 (N_1997,In_1621,In_1570);
and U1998 (N_1998,In_2211,In_2231);
xnor U1999 (N_1999,In_455,In_1258);
nor U2000 (N_2000,In_25,In_2336);
and U2001 (N_2001,In_788,In_522);
and U2002 (N_2002,In_2792,In_985);
nor U2003 (N_2003,In_1630,In_346);
and U2004 (N_2004,In_2134,In_1177);
and U2005 (N_2005,In_1064,In_1630);
nand U2006 (N_2006,In_2445,In_903);
nor U2007 (N_2007,In_2914,In_362);
nand U2008 (N_2008,In_1543,In_1223);
nor U2009 (N_2009,In_2646,In_2889);
or U2010 (N_2010,In_2644,In_1474);
or U2011 (N_2011,In_2815,In_1622);
xor U2012 (N_2012,In_2033,In_718);
nor U2013 (N_2013,In_2423,In_224);
and U2014 (N_2014,In_1527,In_1494);
nand U2015 (N_2015,In_1356,In_855);
or U2016 (N_2016,In_1196,In_1530);
and U2017 (N_2017,In_1060,In_1294);
nor U2018 (N_2018,In_141,In_1289);
nand U2019 (N_2019,In_563,In_1070);
and U2020 (N_2020,In_468,In_247);
nor U2021 (N_2021,In_2378,In_1301);
and U2022 (N_2022,In_2494,In_1403);
and U2023 (N_2023,In_1856,In_1630);
nand U2024 (N_2024,In_349,In_1461);
nand U2025 (N_2025,In_2334,In_1610);
or U2026 (N_2026,In_1477,In_2554);
and U2027 (N_2027,In_2646,In_2787);
nor U2028 (N_2028,In_1541,In_1475);
nor U2029 (N_2029,In_1595,In_2493);
and U2030 (N_2030,In_1137,In_1366);
nor U2031 (N_2031,In_2538,In_1877);
nor U2032 (N_2032,In_2863,In_667);
or U2033 (N_2033,In_73,In_2604);
nand U2034 (N_2034,In_2681,In_1434);
nor U2035 (N_2035,In_2978,In_2384);
nor U2036 (N_2036,In_1669,In_360);
nand U2037 (N_2037,In_1674,In_1639);
nand U2038 (N_2038,In_2446,In_1018);
or U2039 (N_2039,In_2043,In_1808);
or U2040 (N_2040,In_2362,In_797);
nor U2041 (N_2041,In_1076,In_2668);
and U2042 (N_2042,In_243,In_2362);
and U2043 (N_2043,In_1217,In_2768);
and U2044 (N_2044,In_1064,In_2046);
and U2045 (N_2045,In_517,In_1874);
nand U2046 (N_2046,In_2834,In_1548);
nand U2047 (N_2047,In_2349,In_484);
xnor U2048 (N_2048,In_1458,In_211);
nor U2049 (N_2049,In_2849,In_345);
and U2050 (N_2050,In_1668,In_1380);
nor U2051 (N_2051,In_1755,In_464);
or U2052 (N_2052,In_845,In_1871);
nor U2053 (N_2053,In_453,In_1893);
nor U2054 (N_2054,In_464,In_456);
xor U2055 (N_2055,In_198,In_1748);
nor U2056 (N_2056,In_1391,In_124);
nor U2057 (N_2057,In_467,In_1379);
and U2058 (N_2058,In_375,In_80);
or U2059 (N_2059,In_1528,In_2093);
nor U2060 (N_2060,In_2770,In_2672);
xor U2061 (N_2061,In_1133,In_1554);
nor U2062 (N_2062,In_655,In_1500);
xnor U2063 (N_2063,In_1872,In_1004);
and U2064 (N_2064,In_2673,In_68);
nand U2065 (N_2065,In_1273,In_1078);
xor U2066 (N_2066,In_1893,In_327);
and U2067 (N_2067,In_1716,In_570);
nand U2068 (N_2068,In_2532,In_1890);
nor U2069 (N_2069,In_2728,In_1708);
nor U2070 (N_2070,In_1899,In_604);
nand U2071 (N_2071,In_2131,In_319);
and U2072 (N_2072,In_436,In_55);
nand U2073 (N_2073,In_511,In_620);
xnor U2074 (N_2074,In_1897,In_2662);
xnor U2075 (N_2075,In_1733,In_2559);
and U2076 (N_2076,In_2363,In_1935);
nor U2077 (N_2077,In_1096,In_360);
nand U2078 (N_2078,In_2780,In_1167);
nand U2079 (N_2079,In_902,In_2509);
nand U2080 (N_2080,In_254,In_2450);
nand U2081 (N_2081,In_826,In_432);
xor U2082 (N_2082,In_642,In_54);
or U2083 (N_2083,In_2679,In_2567);
nor U2084 (N_2084,In_793,In_2969);
and U2085 (N_2085,In_1486,In_2174);
nor U2086 (N_2086,In_165,In_890);
or U2087 (N_2087,In_501,In_358);
and U2088 (N_2088,In_2173,In_2830);
or U2089 (N_2089,In_1430,In_2111);
nor U2090 (N_2090,In_490,In_740);
or U2091 (N_2091,In_577,In_603);
nor U2092 (N_2092,In_1712,In_1980);
xor U2093 (N_2093,In_305,In_2729);
nor U2094 (N_2094,In_2892,In_368);
nand U2095 (N_2095,In_2611,In_1188);
or U2096 (N_2096,In_1450,In_880);
and U2097 (N_2097,In_2111,In_2461);
nor U2098 (N_2098,In_1062,In_990);
or U2099 (N_2099,In_829,In_1652);
nor U2100 (N_2100,In_498,In_2167);
or U2101 (N_2101,In_1987,In_1315);
xor U2102 (N_2102,In_2254,In_1697);
nand U2103 (N_2103,In_1511,In_825);
nand U2104 (N_2104,In_843,In_2765);
nor U2105 (N_2105,In_1851,In_177);
nor U2106 (N_2106,In_691,In_200);
or U2107 (N_2107,In_2189,In_1687);
nor U2108 (N_2108,In_2026,In_1447);
or U2109 (N_2109,In_2502,In_1437);
nand U2110 (N_2110,In_1950,In_2646);
and U2111 (N_2111,In_2340,In_1398);
nor U2112 (N_2112,In_2800,In_2144);
or U2113 (N_2113,In_2858,In_953);
nor U2114 (N_2114,In_1599,In_2587);
and U2115 (N_2115,In_797,In_283);
and U2116 (N_2116,In_2824,In_2437);
and U2117 (N_2117,In_98,In_1839);
or U2118 (N_2118,In_2705,In_760);
or U2119 (N_2119,In_2633,In_224);
and U2120 (N_2120,In_932,In_1396);
nand U2121 (N_2121,In_1449,In_2582);
nand U2122 (N_2122,In_1415,In_1682);
and U2123 (N_2123,In_2237,In_2495);
nor U2124 (N_2124,In_872,In_1203);
and U2125 (N_2125,In_2296,In_2873);
or U2126 (N_2126,In_657,In_1363);
nand U2127 (N_2127,In_487,In_1495);
xor U2128 (N_2128,In_651,In_1202);
nor U2129 (N_2129,In_1763,In_1842);
nand U2130 (N_2130,In_1796,In_433);
nand U2131 (N_2131,In_2696,In_663);
and U2132 (N_2132,In_221,In_2845);
nand U2133 (N_2133,In_2949,In_858);
and U2134 (N_2134,In_942,In_435);
and U2135 (N_2135,In_1544,In_2353);
nor U2136 (N_2136,In_2737,In_488);
nor U2137 (N_2137,In_2349,In_405);
xnor U2138 (N_2138,In_2827,In_2256);
nor U2139 (N_2139,In_934,In_2331);
nor U2140 (N_2140,In_2167,In_1825);
and U2141 (N_2141,In_1701,In_1790);
nor U2142 (N_2142,In_2615,In_922);
or U2143 (N_2143,In_2114,In_1485);
nor U2144 (N_2144,In_2248,In_1539);
or U2145 (N_2145,In_445,In_1961);
nor U2146 (N_2146,In_1791,In_379);
or U2147 (N_2147,In_2367,In_543);
xnor U2148 (N_2148,In_557,In_1556);
nand U2149 (N_2149,In_2004,In_1468);
nand U2150 (N_2150,In_349,In_1757);
and U2151 (N_2151,In_1691,In_209);
nand U2152 (N_2152,In_2530,In_868);
or U2153 (N_2153,In_1111,In_479);
nand U2154 (N_2154,In_2273,In_1326);
nand U2155 (N_2155,In_2813,In_1308);
nand U2156 (N_2156,In_1613,In_904);
or U2157 (N_2157,In_2017,In_2113);
and U2158 (N_2158,In_1060,In_2908);
and U2159 (N_2159,In_2435,In_2675);
nand U2160 (N_2160,In_2960,In_1750);
nand U2161 (N_2161,In_809,In_1960);
nor U2162 (N_2162,In_650,In_157);
nor U2163 (N_2163,In_451,In_250);
xor U2164 (N_2164,In_1513,In_2514);
nor U2165 (N_2165,In_2438,In_2504);
xor U2166 (N_2166,In_2992,In_548);
nor U2167 (N_2167,In_1150,In_2694);
nand U2168 (N_2168,In_1341,In_1519);
nor U2169 (N_2169,In_1038,In_2914);
nor U2170 (N_2170,In_1655,In_1909);
nor U2171 (N_2171,In_1347,In_2245);
nand U2172 (N_2172,In_2618,In_193);
nor U2173 (N_2173,In_1850,In_1100);
and U2174 (N_2174,In_414,In_1636);
and U2175 (N_2175,In_989,In_2705);
xor U2176 (N_2176,In_307,In_245);
and U2177 (N_2177,In_2212,In_132);
and U2178 (N_2178,In_2680,In_1216);
and U2179 (N_2179,In_2826,In_2302);
and U2180 (N_2180,In_1049,In_1690);
nand U2181 (N_2181,In_700,In_1846);
nor U2182 (N_2182,In_2250,In_1935);
or U2183 (N_2183,In_1726,In_1311);
nand U2184 (N_2184,In_2995,In_60);
nor U2185 (N_2185,In_2763,In_425);
nand U2186 (N_2186,In_1008,In_696);
nand U2187 (N_2187,In_2476,In_1850);
nor U2188 (N_2188,In_911,In_2742);
and U2189 (N_2189,In_2826,In_2406);
nand U2190 (N_2190,In_1850,In_829);
or U2191 (N_2191,In_1390,In_2546);
xnor U2192 (N_2192,In_348,In_1155);
nand U2193 (N_2193,In_44,In_2299);
nand U2194 (N_2194,In_2220,In_2333);
and U2195 (N_2195,In_2974,In_1108);
and U2196 (N_2196,In_61,In_2857);
nand U2197 (N_2197,In_1161,In_2907);
or U2198 (N_2198,In_2455,In_2896);
or U2199 (N_2199,In_2621,In_27);
or U2200 (N_2200,In_1879,In_1844);
nor U2201 (N_2201,In_37,In_932);
nand U2202 (N_2202,In_2711,In_1659);
or U2203 (N_2203,In_1225,In_1549);
and U2204 (N_2204,In_1223,In_670);
and U2205 (N_2205,In_317,In_1541);
and U2206 (N_2206,In_519,In_2292);
or U2207 (N_2207,In_84,In_1402);
nand U2208 (N_2208,In_1069,In_291);
nand U2209 (N_2209,In_838,In_302);
xor U2210 (N_2210,In_2842,In_1783);
xnor U2211 (N_2211,In_2578,In_1247);
nand U2212 (N_2212,In_1528,In_2329);
or U2213 (N_2213,In_225,In_180);
and U2214 (N_2214,In_2013,In_957);
nor U2215 (N_2215,In_919,In_1243);
and U2216 (N_2216,In_2203,In_774);
and U2217 (N_2217,In_2439,In_2701);
nand U2218 (N_2218,In_2325,In_2342);
or U2219 (N_2219,In_1284,In_2558);
and U2220 (N_2220,In_126,In_810);
nor U2221 (N_2221,In_391,In_174);
nor U2222 (N_2222,In_1349,In_2074);
or U2223 (N_2223,In_2895,In_1666);
nand U2224 (N_2224,In_2017,In_2373);
nand U2225 (N_2225,In_576,In_839);
xnor U2226 (N_2226,In_768,In_1876);
nand U2227 (N_2227,In_2695,In_882);
and U2228 (N_2228,In_2321,In_1039);
nand U2229 (N_2229,In_2382,In_290);
nand U2230 (N_2230,In_332,In_1802);
or U2231 (N_2231,In_2130,In_839);
nor U2232 (N_2232,In_2772,In_549);
nor U2233 (N_2233,In_1105,In_2856);
or U2234 (N_2234,In_2883,In_290);
nand U2235 (N_2235,In_1168,In_1606);
or U2236 (N_2236,In_2409,In_715);
nor U2237 (N_2237,In_627,In_1800);
nor U2238 (N_2238,In_1461,In_1152);
nor U2239 (N_2239,In_2552,In_694);
nor U2240 (N_2240,In_2527,In_685);
nor U2241 (N_2241,In_1059,In_735);
nand U2242 (N_2242,In_1630,In_645);
and U2243 (N_2243,In_996,In_2346);
and U2244 (N_2244,In_2125,In_2062);
nand U2245 (N_2245,In_813,In_1699);
or U2246 (N_2246,In_1874,In_1448);
or U2247 (N_2247,In_1719,In_26);
nor U2248 (N_2248,In_2761,In_173);
or U2249 (N_2249,In_2308,In_2677);
nand U2250 (N_2250,In_1710,In_931);
or U2251 (N_2251,In_349,In_2795);
and U2252 (N_2252,In_2809,In_193);
nor U2253 (N_2253,In_1088,In_2731);
nor U2254 (N_2254,In_2729,In_1383);
nand U2255 (N_2255,In_2358,In_2561);
nand U2256 (N_2256,In_946,In_2047);
or U2257 (N_2257,In_1017,In_1614);
nand U2258 (N_2258,In_2310,In_2065);
or U2259 (N_2259,In_338,In_585);
nand U2260 (N_2260,In_1493,In_2689);
nand U2261 (N_2261,In_398,In_2527);
and U2262 (N_2262,In_207,In_2543);
nor U2263 (N_2263,In_2938,In_2905);
nand U2264 (N_2264,In_457,In_2125);
or U2265 (N_2265,In_2850,In_1639);
xor U2266 (N_2266,In_322,In_1057);
nor U2267 (N_2267,In_125,In_1594);
or U2268 (N_2268,In_1557,In_1920);
or U2269 (N_2269,In_1944,In_1458);
or U2270 (N_2270,In_2716,In_281);
and U2271 (N_2271,In_668,In_1137);
xor U2272 (N_2272,In_937,In_1014);
nand U2273 (N_2273,In_653,In_1686);
or U2274 (N_2274,In_2475,In_2236);
nand U2275 (N_2275,In_484,In_836);
and U2276 (N_2276,In_1760,In_113);
and U2277 (N_2277,In_1114,In_1716);
nand U2278 (N_2278,In_1675,In_964);
or U2279 (N_2279,In_454,In_1244);
nand U2280 (N_2280,In_2749,In_1558);
nor U2281 (N_2281,In_2234,In_1591);
or U2282 (N_2282,In_1158,In_1770);
and U2283 (N_2283,In_2531,In_918);
and U2284 (N_2284,In_815,In_967);
and U2285 (N_2285,In_1208,In_1125);
or U2286 (N_2286,In_1345,In_2349);
nand U2287 (N_2287,In_519,In_2328);
and U2288 (N_2288,In_1568,In_735);
nand U2289 (N_2289,In_1621,In_1919);
xor U2290 (N_2290,In_328,In_1932);
and U2291 (N_2291,In_2962,In_1152);
or U2292 (N_2292,In_2273,In_294);
and U2293 (N_2293,In_2942,In_1507);
xor U2294 (N_2294,In_2666,In_2957);
nor U2295 (N_2295,In_2324,In_137);
and U2296 (N_2296,In_1566,In_2510);
nor U2297 (N_2297,In_639,In_2821);
nand U2298 (N_2298,In_313,In_847);
nand U2299 (N_2299,In_2176,In_2256);
nand U2300 (N_2300,In_2199,In_1173);
xor U2301 (N_2301,In_1683,In_2015);
nor U2302 (N_2302,In_1000,In_2947);
nor U2303 (N_2303,In_580,In_631);
nor U2304 (N_2304,In_1140,In_948);
and U2305 (N_2305,In_1163,In_2714);
and U2306 (N_2306,In_2505,In_430);
or U2307 (N_2307,In_2364,In_432);
nor U2308 (N_2308,In_2779,In_1880);
and U2309 (N_2309,In_2981,In_1650);
xnor U2310 (N_2310,In_1843,In_2028);
or U2311 (N_2311,In_1783,In_1212);
or U2312 (N_2312,In_16,In_2140);
or U2313 (N_2313,In_827,In_46);
nor U2314 (N_2314,In_2237,In_541);
nand U2315 (N_2315,In_452,In_1269);
nor U2316 (N_2316,In_2279,In_2126);
and U2317 (N_2317,In_187,In_1537);
nor U2318 (N_2318,In_2356,In_2290);
or U2319 (N_2319,In_1438,In_2690);
and U2320 (N_2320,In_2319,In_2063);
and U2321 (N_2321,In_1189,In_1998);
nor U2322 (N_2322,In_1442,In_1828);
nand U2323 (N_2323,In_2419,In_2775);
and U2324 (N_2324,In_2518,In_29);
and U2325 (N_2325,In_2108,In_280);
nor U2326 (N_2326,In_2692,In_2850);
and U2327 (N_2327,In_872,In_2365);
nand U2328 (N_2328,In_2836,In_697);
nand U2329 (N_2329,In_1947,In_227);
xnor U2330 (N_2330,In_966,In_1394);
and U2331 (N_2331,In_1559,In_298);
and U2332 (N_2332,In_522,In_2101);
nor U2333 (N_2333,In_2335,In_2765);
nor U2334 (N_2334,In_2016,In_1807);
or U2335 (N_2335,In_1690,In_339);
nand U2336 (N_2336,In_1708,In_2105);
nor U2337 (N_2337,In_145,In_285);
or U2338 (N_2338,In_759,In_1234);
or U2339 (N_2339,In_445,In_783);
and U2340 (N_2340,In_1259,In_1857);
nor U2341 (N_2341,In_1289,In_382);
and U2342 (N_2342,In_1956,In_1752);
nor U2343 (N_2343,In_2548,In_1916);
xor U2344 (N_2344,In_1070,In_1151);
and U2345 (N_2345,In_1539,In_452);
nor U2346 (N_2346,In_321,In_2991);
and U2347 (N_2347,In_835,In_519);
and U2348 (N_2348,In_1306,In_1256);
nor U2349 (N_2349,In_1879,In_2681);
nand U2350 (N_2350,In_308,In_1815);
and U2351 (N_2351,In_2061,In_1237);
and U2352 (N_2352,In_2398,In_1664);
nor U2353 (N_2353,In_123,In_2389);
nand U2354 (N_2354,In_2980,In_309);
nand U2355 (N_2355,In_2970,In_1819);
nor U2356 (N_2356,In_603,In_2070);
and U2357 (N_2357,In_2195,In_2894);
and U2358 (N_2358,In_2117,In_2628);
or U2359 (N_2359,In_1205,In_2055);
and U2360 (N_2360,In_390,In_669);
nor U2361 (N_2361,In_796,In_451);
xor U2362 (N_2362,In_379,In_1772);
and U2363 (N_2363,In_762,In_2650);
nand U2364 (N_2364,In_2694,In_1673);
nand U2365 (N_2365,In_902,In_1287);
nor U2366 (N_2366,In_1879,In_330);
and U2367 (N_2367,In_2494,In_1029);
nand U2368 (N_2368,In_2611,In_1251);
nor U2369 (N_2369,In_2174,In_1090);
and U2370 (N_2370,In_1517,In_2571);
or U2371 (N_2371,In_2635,In_1914);
xnor U2372 (N_2372,In_604,In_1926);
and U2373 (N_2373,In_582,In_68);
nand U2374 (N_2374,In_953,In_1163);
nand U2375 (N_2375,In_43,In_1125);
or U2376 (N_2376,In_976,In_2546);
or U2377 (N_2377,In_64,In_1917);
or U2378 (N_2378,In_2914,In_1536);
or U2379 (N_2379,In_2067,In_311);
nand U2380 (N_2380,In_2640,In_1760);
nand U2381 (N_2381,In_2082,In_1257);
or U2382 (N_2382,In_2730,In_348);
nor U2383 (N_2383,In_78,In_2647);
or U2384 (N_2384,In_2907,In_2717);
nor U2385 (N_2385,In_851,In_952);
xnor U2386 (N_2386,In_357,In_1574);
or U2387 (N_2387,In_741,In_1484);
or U2388 (N_2388,In_2860,In_2066);
nor U2389 (N_2389,In_94,In_2504);
nor U2390 (N_2390,In_119,In_2760);
nand U2391 (N_2391,In_118,In_1988);
nand U2392 (N_2392,In_483,In_3);
nor U2393 (N_2393,In_480,In_2794);
nand U2394 (N_2394,In_1707,In_492);
nand U2395 (N_2395,In_2597,In_2552);
nor U2396 (N_2396,In_857,In_1380);
nor U2397 (N_2397,In_2999,In_216);
or U2398 (N_2398,In_2102,In_2942);
or U2399 (N_2399,In_2244,In_2604);
and U2400 (N_2400,In_2941,In_65);
or U2401 (N_2401,In_491,In_1939);
nand U2402 (N_2402,In_2984,In_2977);
xnor U2403 (N_2403,In_1447,In_1991);
nand U2404 (N_2404,In_146,In_340);
or U2405 (N_2405,In_2994,In_2212);
or U2406 (N_2406,In_2003,In_1978);
nor U2407 (N_2407,In_794,In_1783);
nor U2408 (N_2408,In_2730,In_2576);
and U2409 (N_2409,In_56,In_2985);
and U2410 (N_2410,In_957,In_2064);
or U2411 (N_2411,In_85,In_847);
nor U2412 (N_2412,In_1436,In_2518);
and U2413 (N_2413,In_2313,In_2019);
nand U2414 (N_2414,In_618,In_1121);
and U2415 (N_2415,In_2846,In_1982);
nand U2416 (N_2416,In_889,In_380);
and U2417 (N_2417,In_514,In_853);
nand U2418 (N_2418,In_2376,In_1533);
and U2419 (N_2419,In_1636,In_1148);
nand U2420 (N_2420,In_535,In_1387);
and U2421 (N_2421,In_2451,In_2148);
and U2422 (N_2422,In_1281,In_2612);
xnor U2423 (N_2423,In_2557,In_1080);
nand U2424 (N_2424,In_705,In_1035);
nand U2425 (N_2425,In_1759,In_685);
nor U2426 (N_2426,In_2702,In_1903);
or U2427 (N_2427,In_2098,In_2164);
or U2428 (N_2428,In_86,In_38);
and U2429 (N_2429,In_2862,In_1446);
xor U2430 (N_2430,In_2243,In_2909);
nand U2431 (N_2431,In_2910,In_88);
nand U2432 (N_2432,In_1066,In_121);
or U2433 (N_2433,In_2294,In_1758);
and U2434 (N_2434,In_801,In_1389);
and U2435 (N_2435,In_1685,In_826);
nor U2436 (N_2436,In_1447,In_506);
xnor U2437 (N_2437,In_1011,In_2488);
nor U2438 (N_2438,In_1717,In_498);
or U2439 (N_2439,In_2729,In_199);
and U2440 (N_2440,In_2909,In_1353);
and U2441 (N_2441,In_868,In_792);
nor U2442 (N_2442,In_139,In_2362);
and U2443 (N_2443,In_2792,In_2788);
and U2444 (N_2444,In_1172,In_2190);
nand U2445 (N_2445,In_1007,In_609);
nand U2446 (N_2446,In_556,In_1260);
and U2447 (N_2447,In_755,In_2802);
nor U2448 (N_2448,In_2280,In_2233);
nand U2449 (N_2449,In_2137,In_1153);
xor U2450 (N_2450,In_332,In_2667);
nand U2451 (N_2451,In_2179,In_805);
or U2452 (N_2452,In_1801,In_2858);
or U2453 (N_2453,In_545,In_2646);
and U2454 (N_2454,In_758,In_655);
and U2455 (N_2455,In_501,In_2058);
xor U2456 (N_2456,In_303,In_672);
xor U2457 (N_2457,In_2282,In_980);
xor U2458 (N_2458,In_208,In_1818);
and U2459 (N_2459,In_1431,In_1012);
and U2460 (N_2460,In_1056,In_2938);
nand U2461 (N_2461,In_2333,In_726);
nor U2462 (N_2462,In_2593,In_1827);
nand U2463 (N_2463,In_1556,In_1853);
nor U2464 (N_2464,In_63,In_2862);
or U2465 (N_2465,In_699,In_1384);
xor U2466 (N_2466,In_917,In_2995);
and U2467 (N_2467,In_2072,In_1541);
or U2468 (N_2468,In_690,In_1178);
xnor U2469 (N_2469,In_2103,In_1408);
nor U2470 (N_2470,In_1679,In_253);
nor U2471 (N_2471,In_2202,In_2253);
or U2472 (N_2472,In_240,In_1558);
nor U2473 (N_2473,In_542,In_2133);
nand U2474 (N_2474,In_2268,In_509);
and U2475 (N_2475,In_475,In_183);
nand U2476 (N_2476,In_1549,In_1271);
xor U2477 (N_2477,In_1574,In_1403);
nor U2478 (N_2478,In_2255,In_923);
nand U2479 (N_2479,In_2110,In_1238);
nor U2480 (N_2480,In_2305,In_1208);
nand U2481 (N_2481,In_2383,In_2333);
and U2482 (N_2482,In_1126,In_2502);
nand U2483 (N_2483,In_1064,In_847);
nor U2484 (N_2484,In_2046,In_2751);
nand U2485 (N_2485,In_39,In_1584);
xnor U2486 (N_2486,In_2368,In_1883);
nand U2487 (N_2487,In_2795,In_2940);
and U2488 (N_2488,In_301,In_466);
nand U2489 (N_2489,In_2479,In_1240);
nand U2490 (N_2490,In_508,In_969);
nand U2491 (N_2491,In_1638,In_1345);
xor U2492 (N_2492,In_1220,In_1069);
nor U2493 (N_2493,In_1769,In_2754);
or U2494 (N_2494,In_2703,In_1460);
or U2495 (N_2495,In_1372,In_1518);
or U2496 (N_2496,In_2916,In_1567);
nor U2497 (N_2497,In_2349,In_191);
and U2498 (N_2498,In_842,In_2425);
or U2499 (N_2499,In_2823,In_2003);
and U2500 (N_2500,In_2317,In_1548);
xor U2501 (N_2501,In_2162,In_109);
nor U2502 (N_2502,In_2132,In_1458);
and U2503 (N_2503,In_1427,In_1771);
nor U2504 (N_2504,In_1807,In_2969);
or U2505 (N_2505,In_2973,In_207);
or U2506 (N_2506,In_1538,In_1502);
nand U2507 (N_2507,In_1282,In_1909);
or U2508 (N_2508,In_692,In_1209);
nor U2509 (N_2509,In_526,In_1984);
or U2510 (N_2510,In_2007,In_2763);
nor U2511 (N_2511,In_2680,In_1895);
nor U2512 (N_2512,In_917,In_1242);
nand U2513 (N_2513,In_2898,In_1073);
xnor U2514 (N_2514,In_2908,In_2612);
nand U2515 (N_2515,In_2520,In_1397);
nand U2516 (N_2516,In_1342,In_2535);
nand U2517 (N_2517,In_2038,In_706);
nor U2518 (N_2518,In_2281,In_2431);
or U2519 (N_2519,In_2583,In_916);
xor U2520 (N_2520,In_2490,In_1667);
nand U2521 (N_2521,In_2250,In_284);
or U2522 (N_2522,In_736,In_746);
xor U2523 (N_2523,In_798,In_2513);
or U2524 (N_2524,In_570,In_2195);
nor U2525 (N_2525,In_1452,In_116);
and U2526 (N_2526,In_2396,In_2093);
and U2527 (N_2527,In_1607,In_1349);
or U2528 (N_2528,In_627,In_1133);
or U2529 (N_2529,In_326,In_96);
nor U2530 (N_2530,In_227,In_372);
nand U2531 (N_2531,In_2020,In_7);
nand U2532 (N_2532,In_2550,In_1963);
nand U2533 (N_2533,In_832,In_2134);
and U2534 (N_2534,In_2020,In_270);
nand U2535 (N_2535,In_2321,In_2989);
nor U2536 (N_2536,In_988,In_1746);
and U2537 (N_2537,In_191,In_1175);
nand U2538 (N_2538,In_1742,In_683);
and U2539 (N_2539,In_236,In_2973);
nor U2540 (N_2540,In_360,In_405);
xnor U2541 (N_2541,In_2176,In_2293);
nor U2542 (N_2542,In_140,In_2734);
or U2543 (N_2543,In_2256,In_1837);
nor U2544 (N_2544,In_1020,In_2734);
and U2545 (N_2545,In_2742,In_725);
or U2546 (N_2546,In_954,In_759);
nand U2547 (N_2547,In_1784,In_2110);
xnor U2548 (N_2548,In_1665,In_1453);
or U2549 (N_2549,In_312,In_897);
or U2550 (N_2550,In_1058,In_930);
nand U2551 (N_2551,In_2050,In_2449);
or U2552 (N_2552,In_1125,In_702);
nand U2553 (N_2553,In_1177,In_936);
and U2554 (N_2554,In_2541,In_1719);
nor U2555 (N_2555,In_1137,In_775);
nand U2556 (N_2556,In_1088,In_2310);
nand U2557 (N_2557,In_600,In_2641);
or U2558 (N_2558,In_1338,In_2109);
or U2559 (N_2559,In_1792,In_1191);
or U2560 (N_2560,In_2172,In_2754);
and U2561 (N_2561,In_1235,In_2833);
nand U2562 (N_2562,In_2029,In_1192);
or U2563 (N_2563,In_2312,In_2245);
or U2564 (N_2564,In_1506,In_1930);
or U2565 (N_2565,In_2189,In_112);
xnor U2566 (N_2566,In_42,In_2798);
xnor U2567 (N_2567,In_1543,In_667);
and U2568 (N_2568,In_24,In_784);
nand U2569 (N_2569,In_94,In_2310);
xor U2570 (N_2570,In_67,In_1242);
nand U2571 (N_2571,In_1139,In_2506);
nor U2572 (N_2572,In_1002,In_2651);
nor U2573 (N_2573,In_1818,In_2195);
nor U2574 (N_2574,In_1376,In_988);
xnor U2575 (N_2575,In_1175,In_703);
and U2576 (N_2576,In_1201,In_831);
nand U2577 (N_2577,In_2823,In_1798);
xnor U2578 (N_2578,In_2735,In_2974);
or U2579 (N_2579,In_1587,In_1215);
or U2580 (N_2580,In_2962,In_1632);
or U2581 (N_2581,In_267,In_1742);
nand U2582 (N_2582,In_515,In_2954);
and U2583 (N_2583,In_1952,In_4);
nor U2584 (N_2584,In_1612,In_1900);
nor U2585 (N_2585,In_254,In_2500);
xnor U2586 (N_2586,In_2864,In_319);
and U2587 (N_2587,In_1666,In_2810);
nor U2588 (N_2588,In_2980,In_872);
nor U2589 (N_2589,In_2519,In_1681);
nand U2590 (N_2590,In_1279,In_2080);
nand U2591 (N_2591,In_1241,In_761);
nand U2592 (N_2592,In_1988,In_2870);
nor U2593 (N_2593,In_48,In_886);
nor U2594 (N_2594,In_1367,In_1556);
and U2595 (N_2595,In_1474,In_2123);
and U2596 (N_2596,In_173,In_2442);
nor U2597 (N_2597,In_1742,In_1780);
nand U2598 (N_2598,In_1085,In_460);
nor U2599 (N_2599,In_1080,In_2853);
and U2600 (N_2600,In_418,In_1469);
nor U2601 (N_2601,In_1446,In_939);
nand U2602 (N_2602,In_2302,In_2349);
nor U2603 (N_2603,In_738,In_1950);
or U2604 (N_2604,In_950,In_2915);
nand U2605 (N_2605,In_1767,In_1210);
and U2606 (N_2606,In_1425,In_2466);
nand U2607 (N_2607,In_1175,In_1408);
nor U2608 (N_2608,In_1659,In_352);
nor U2609 (N_2609,In_1222,In_1085);
nand U2610 (N_2610,In_466,In_580);
nor U2611 (N_2611,In_1620,In_2485);
nor U2612 (N_2612,In_1214,In_2798);
and U2613 (N_2613,In_2012,In_1150);
nand U2614 (N_2614,In_597,In_968);
xor U2615 (N_2615,In_2492,In_1197);
nor U2616 (N_2616,In_2278,In_323);
or U2617 (N_2617,In_1796,In_2254);
xnor U2618 (N_2618,In_1557,In_2830);
or U2619 (N_2619,In_2078,In_2565);
nor U2620 (N_2620,In_2175,In_2702);
nor U2621 (N_2621,In_1224,In_1847);
or U2622 (N_2622,In_1814,In_128);
nor U2623 (N_2623,In_1932,In_1623);
and U2624 (N_2624,In_1236,In_1321);
or U2625 (N_2625,In_2672,In_214);
nand U2626 (N_2626,In_2881,In_759);
or U2627 (N_2627,In_2277,In_681);
and U2628 (N_2628,In_1372,In_2980);
or U2629 (N_2629,In_364,In_22);
or U2630 (N_2630,In_2180,In_2853);
and U2631 (N_2631,In_1727,In_2750);
nor U2632 (N_2632,In_1771,In_2796);
nor U2633 (N_2633,In_2489,In_2403);
and U2634 (N_2634,In_2147,In_2611);
nand U2635 (N_2635,In_1498,In_2230);
or U2636 (N_2636,In_17,In_2298);
nor U2637 (N_2637,In_1273,In_2795);
nand U2638 (N_2638,In_2566,In_360);
nor U2639 (N_2639,In_2681,In_1565);
xor U2640 (N_2640,In_2109,In_1373);
and U2641 (N_2641,In_1848,In_2183);
and U2642 (N_2642,In_916,In_463);
xor U2643 (N_2643,In_888,In_2886);
and U2644 (N_2644,In_2665,In_522);
xnor U2645 (N_2645,In_649,In_1003);
nor U2646 (N_2646,In_1737,In_1045);
and U2647 (N_2647,In_981,In_2422);
nor U2648 (N_2648,In_1995,In_2816);
nor U2649 (N_2649,In_2165,In_821);
nand U2650 (N_2650,In_1478,In_2781);
and U2651 (N_2651,In_1425,In_638);
nand U2652 (N_2652,In_629,In_560);
and U2653 (N_2653,In_815,In_1858);
nor U2654 (N_2654,In_2938,In_1260);
nor U2655 (N_2655,In_38,In_2661);
or U2656 (N_2656,In_457,In_426);
nand U2657 (N_2657,In_2143,In_2542);
xnor U2658 (N_2658,In_1830,In_108);
nand U2659 (N_2659,In_378,In_830);
or U2660 (N_2660,In_468,In_2071);
xor U2661 (N_2661,In_1681,In_94);
and U2662 (N_2662,In_1451,In_1619);
and U2663 (N_2663,In_918,In_2558);
and U2664 (N_2664,In_825,In_2495);
nand U2665 (N_2665,In_1421,In_2357);
nor U2666 (N_2666,In_281,In_426);
and U2667 (N_2667,In_470,In_1021);
nor U2668 (N_2668,In_254,In_1699);
or U2669 (N_2669,In_2756,In_295);
and U2670 (N_2670,In_2417,In_884);
and U2671 (N_2671,In_647,In_2240);
nor U2672 (N_2672,In_935,In_586);
and U2673 (N_2673,In_2248,In_2339);
nor U2674 (N_2674,In_981,In_454);
nor U2675 (N_2675,In_760,In_1262);
nand U2676 (N_2676,In_2915,In_867);
nor U2677 (N_2677,In_1935,In_1539);
nand U2678 (N_2678,In_94,In_1015);
and U2679 (N_2679,In_2228,In_110);
nand U2680 (N_2680,In_2600,In_2024);
nand U2681 (N_2681,In_345,In_1159);
nand U2682 (N_2682,In_947,In_560);
or U2683 (N_2683,In_45,In_920);
or U2684 (N_2684,In_907,In_2432);
or U2685 (N_2685,In_2809,In_811);
xor U2686 (N_2686,In_161,In_247);
nor U2687 (N_2687,In_437,In_1489);
nor U2688 (N_2688,In_2737,In_1918);
xnor U2689 (N_2689,In_2074,In_890);
nor U2690 (N_2690,In_2457,In_151);
xnor U2691 (N_2691,In_1222,In_2910);
nor U2692 (N_2692,In_232,In_1337);
xor U2693 (N_2693,In_60,In_1985);
nor U2694 (N_2694,In_2486,In_1423);
nor U2695 (N_2695,In_1208,In_1799);
nor U2696 (N_2696,In_1916,In_2526);
or U2697 (N_2697,In_587,In_1236);
nor U2698 (N_2698,In_1324,In_1244);
nor U2699 (N_2699,In_2222,In_17);
nand U2700 (N_2700,In_934,In_1109);
nand U2701 (N_2701,In_1622,In_1326);
nor U2702 (N_2702,In_1543,In_1202);
nand U2703 (N_2703,In_2496,In_1186);
nand U2704 (N_2704,In_2031,In_2125);
nand U2705 (N_2705,In_2009,In_1663);
xnor U2706 (N_2706,In_1962,In_698);
nor U2707 (N_2707,In_1552,In_261);
nor U2708 (N_2708,In_792,In_2952);
nand U2709 (N_2709,In_998,In_2586);
nor U2710 (N_2710,In_2259,In_1586);
and U2711 (N_2711,In_91,In_1332);
nand U2712 (N_2712,In_368,In_1023);
or U2713 (N_2713,In_630,In_1229);
xnor U2714 (N_2714,In_2953,In_1408);
or U2715 (N_2715,In_1138,In_2224);
nor U2716 (N_2716,In_2605,In_1778);
nor U2717 (N_2717,In_2272,In_1002);
xor U2718 (N_2718,In_2929,In_2237);
nor U2719 (N_2719,In_2370,In_603);
nand U2720 (N_2720,In_2366,In_1525);
or U2721 (N_2721,In_158,In_2689);
nand U2722 (N_2722,In_1524,In_2477);
nor U2723 (N_2723,In_2828,In_1961);
and U2724 (N_2724,In_2961,In_1702);
or U2725 (N_2725,In_2541,In_52);
nor U2726 (N_2726,In_1733,In_1551);
or U2727 (N_2727,In_741,In_2648);
nor U2728 (N_2728,In_863,In_1841);
nor U2729 (N_2729,In_2401,In_2180);
nand U2730 (N_2730,In_1833,In_2859);
nor U2731 (N_2731,In_1155,In_2147);
and U2732 (N_2732,In_1834,In_2317);
xor U2733 (N_2733,In_2065,In_978);
nor U2734 (N_2734,In_187,In_2128);
and U2735 (N_2735,In_1611,In_893);
nor U2736 (N_2736,In_988,In_2144);
and U2737 (N_2737,In_2839,In_1518);
or U2738 (N_2738,In_2302,In_2052);
nor U2739 (N_2739,In_534,In_784);
or U2740 (N_2740,In_956,In_2843);
nor U2741 (N_2741,In_454,In_2715);
and U2742 (N_2742,In_2787,In_2171);
xor U2743 (N_2743,In_2469,In_150);
or U2744 (N_2744,In_1626,In_211);
or U2745 (N_2745,In_2123,In_1418);
and U2746 (N_2746,In_1381,In_1639);
or U2747 (N_2747,In_2329,In_673);
or U2748 (N_2748,In_406,In_1392);
xnor U2749 (N_2749,In_287,In_707);
xnor U2750 (N_2750,In_2538,In_1756);
and U2751 (N_2751,In_2881,In_187);
and U2752 (N_2752,In_174,In_2835);
nand U2753 (N_2753,In_2657,In_1031);
or U2754 (N_2754,In_2946,In_1004);
or U2755 (N_2755,In_2328,In_1383);
and U2756 (N_2756,In_1063,In_2564);
nand U2757 (N_2757,In_1089,In_998);
nor U2758 (N_2758,In_627,In_783);
and U2759 (N_2759,In_86,In_2335);
nor U2760 (N_2760,In_673,In_1109);
nor U2761 (N_2761,In_65,In_324);
nand U2762 (N_2762,In_913,In_2621);
or U2763 (N_2763,In_271,In_2005);
nor U2764 (N_2764,In_2996,In_230);
xor U2765 (N_2765,In_1004,In_1369);
nor U2766 (N_2766,In_1158,In_2262);
xor U2767 (N_2767,In_1513,In_2030);
and U2768 (N_2768,In_31,In_2975);
nand U2769 (N_2769,In_2958,In_1790);
or U2770 (N_2770,In_605,In_2891);
and U2771 (N_2771,In_696,In_1648);
nor U2772 (N_2772,In_1102,In_1159);
and U2773 (N_2773,In_2040,In_985);
or U2774 (N_2774,In_196,In_185);
nor U2775 (N_2775,In_848,In_331);
nand U2776 (N_2776,In_2966,In_1266);
nor U2777 (N_2777,In_1402,In_1614);
nand U2778 (N_2778,In_944,In_2145);
nor U2779 (N_2779,In_2004,In_962);
or U2780 (N_2780,In_241,In_247);
or U2781 (N_2781,In_1045,In_1249);
xor U2782 (N_2782,In_426,In_2348);
nand U2783 (N_2783,In_2276,In_1011);
or U2784 (N_2784,In_938,In_2730);
and U2785 (N_2785,In_1686,In_2819);
and U2786 (N_2786,In_1255,In_32);
nor U2787 (N_2787,In_2467,In_2301);
xor U2788 (N_2788,In_2435,In_2147);
nand U2789 (N_2789,In_1321,In_2281);
nand U2790 (N_2790,In_1772,In_744);
or U2791 (N_2791,In_2538,In_1016);
nor U2792 (N_2792,In_607,In_1834);
and U2793 (N_2793,In_1251,In_1244);
nand U2794 (N_2794,In_852,In_1814);
or U2795 (N_2795,In_2553,In_1289);
nand U2796 (N_2796,In_1857,In_2606);
or U2797 (N_2797,In_1461,In_1574);
and U2798 (N_2798,In_923,In_2114);
nand U2799 (N_2799,In_2463,In_648);
and U2800 (N_2800,In_2115,In_625);
and U2801 (N_2801,In_1980,In_1251);
nand U2802 (N_2802,In_530,In_1802);
and U2803 (N_2803,In_2786,In_1392);
or U2804 (N_2804,In_2159,In_2742);
or U2805 (N_2805,In_2330,In_2961);
xnor U2806 (N_2806,In_429,In_2534);
and U2807 (N_2807,In_849,In_1574);
or U2808 (N_2808,In_196,In_718);
nand U2809 (N_2809,In_2473,In_175);
and U2810 (N_2810,In_2922,In_2994);
or U2811 (N_2811,In_620,In_378);
xnor U2812 (N_2812,In_403,In_826);
and U2813 (N_2813,In_1398,In_2183);
nand U2814 (N_2814,In_2600,In_2233);
nor U2815 (N_2815,In_1102,In_2010);
or U2816 (N_2816,In_858,In_1);
and U2817 (N_2817,In_1791,In_2750);
or U2818 (N_2818,In_1072,In_719);
and U2819 (N_2819,In_2312,In_2112);
nor U2820 (N_2820,In_1839,In_621);
and U2821 (N_2821,In_2254,In_1493);
xnor U2822 (N_2822,In_2668,In_2431);
or U2823 (N_2823,In_1719,In_1544);
and U2824 (N_2824,In_2649,In_1274);
and U2825 (N_2825,In_2527,In_1588);
or U2826 (N_2826,In_1019,In_1178);
nand U2827 (N_2827,In_13,In_1986);
or U2828 (N_2828,In_829,In_2516);
xor U2829 (N_2829,In_1536,In_505);
and U2830 (N_2830,In_1603,In_1340);
nand U2831 (N_2831,In_2782,In_707);
and U2832 (N_2832,In_294,In_1729);
and U2833 (N_2833,In_2884,In_1777);
nor U2834 (N_2834,In_1038,In_458);
and U2835 (N_2835,In_620,In_18);
and U2836 (N_2836,In_2981,In_2767);
or U2837 (N_2837,In_2182,In_971);
or U2838 (N_2838,In_369,In_151);
and U2839 (N_2839,In_63,In_1514);
xnor U2840 (N_2840,In_2104,In_483);
nand U2841 (N_2841,In_833,In_1136);
and U2842 (N_2842,In_2225,In_2348);
nor U2843 (N_2843,In_1091,In_1520);
or U2844 (N_2844,In_2903,In_585);
and U2845 (N_2845,In_771,In_2938);
and U2846 (N_2846,In_1467,In_2847);
or U2847 (N_2847,In_2290,In_1423);
or U2848 (N_2848,In_2563,In_55);
nor U2849 (N_2849,In_1027,In_1170);
nor U2850 (N_2850,In_283,In_2647);
and U2851 (N_2851,In_1248,In_279);
nand U2852 (N_2852,In_9,In_1502);
nand U2853 (N_2853,In_567,In_1009);
and U2854 (N_2854,In_2662,In_1657);
nand U2855 (N_2855,In_1189,In_1205);
or U2856 (N_2856,In_371,In_2995);
xor U2857 (N_2857,In_1636,In_1846);
and U2858 (N_2858,In_2300,In_970);
nand U2859 (N_2859,In_718,In_879);
nand U2860 (N_2860,In_2311,In_1531);
nand U2861 (N_2861,In_678,In_8);
or U2862 (N_2862,In_1482,In_1157);
nor U2863 (N_2863,In_364,In_1221);
or U2864 (N_2864,In_435,In_1186);
nand U2865 (N_2865,In_1507,In_476);
and U2866 (N_2866,In_1246,In_1003);
nor U2867 (N_2867,In_402,In_504);
xor U2868 (N_2868,In_1531,In_82);
or U2869 (N_2869,In_2157,In_1081);
or U2870 (N_2870,In_2169,In_2012);
and U2871 (N_2871,In_2892,In_1433);
nand U2872 (N_2872,In_1636,In_49);
or U2873 (N_2873,In_2822,In_2646);
nand U2874 (N_2874,In_2445,In_660);
nor U2875 (N_2875,In_375,In_1491);
nand U2876 (N_2876,In_197,In_675);
nor U2877 (N_2877,In_74,In_1515);
and U2878 (N_2878,In_1761,In_1084);
and U2879 (N_2879,In_2440,In_2459);
xor U2880 (N_2880,In_506,In_558);
and U2881 (N_2881,In_2831,In_263);
and U2882 (N_2882,In_2933,In_2703);
or U2883 (N_2883,In_305,In_477);
nor U2884 (N_2884,In_2076,In_209);
nor U2885 (N_2885,In_2572,In_158);
or U2886 (N_2886,In_2171,In_875);
or U2887 (N_2887,In_1551,In_2240);
and U2888 (N_2888,In_230,In_1301);
or U2889 (N_2889,In_1197,In_34);
xor U2890 (N_2890,In_1662,In_612);
nand U2891 (N_2891,In_1746,In_2429);
or U2892 (N_2892,In_2453,In_2620);
nand U2893 (N_2893,In_1231,In_1442);
and U2894 (N_2894,In_2949,In_2766);
or U2895 (N_2895,In_2500,In_954);
and U2896 (N_2896,In_1696,In_1156);
nor U2897 (N_2897,In_1545,In_2632);
nand U2898 (N_2898,In_2824,In_2178);
and U2899 (N_2899,In_2398,In_2724);
or U2900 (N_2900,In_1831,In_1042);
or U2901 (N_2901,In_1999,In_2161);
nand U2902 (N_2902,In_162,In_951);
or U2903 (N_2903,In_2444,In_1288);
and U2904 (N_2904,In_682,In_1041);
and U2905 (N_2905,In_1243,In_120);
nand U2906 (N_2906,In_1629,In_1268);
or U2907 (N_2907,In_1938,In_2066);
and U2908 (N_2908,In_1124,In_702);
nand U2909 (N_2909,In_1506,In_2395);
or U2910 (N_2910,In_2609,In_1937);
or U2911 (N_2911,In_2950,In_2045);
nand U2912 (N_2912,In_2942,In_2339);
nand U2913 (N_2913,In_2778,In_436);
or U2914 (N_2914,In_2856,In_118);
and U2915 (N_2915,In_235,In_1072);
xor U2916 (N_2916,In_1759,In_2120);
nand U2917 (N_2917,In_1313,In_2788);
nor U2918 (N_2918,In_1833,In_1840);
xnor U2919 (N_2919,In_1799,In_1624);
xor U2920 (N_2920,In_692,In_1037);
and U2921 (N_2921,In_2188,In_751);
or U2922 (N_2922,In_2816,In_2358);
and U2923 (N_2923,In_1289,In_2105);
and U2924 (N_2924,In_224,In_951);
nor U2925 (N_2925,In_2385,In_2634);
or U2926 (N_2926,In_1701,In_511);
nand U2927 (N_2927,In_2192,In_204);
or U2928 (N_2928,In_2259,In_1827);
and U2929 (N_2929,In_1521,In_2437);
nand U2930 (N_2930,In_1762,In_2498);
nor U2931 (N_2931,In_1616,In_1874);
nand U2932 (N_2932,In_1077,In_1700);
nor U2933 (N_2933,In_1801,In_2862);
and U2934 (N_2934,In_1693,In_1462);
xor U2935 (N_2935,In_1625,In_1930);
or U2936 (N_2936,In_991,In_247);
nor U2937 (N_2937,In_1284,In_1437);
xor U2938 (N_2938,In_2319,In_1179);
nand U2939 (N_2939,In_848,In_2829);
xor U2940 (N_2940,In_1631,In_337);
nand U2941 (N_2941,In_2785,In_1317);
or U2942 (N_2942,In_49,In_1361);
or U2943 (N_2943,In_2383,In_2830);
nor U2944 (N_2944,In_899,In_395);
nor U2945 (N_2945,In_2921,In_1290);
nor U2946 (N_2946,In_1630,In_1982);
or U2947 (N_2947,In_2761,In_1223);
nor U2948 (N_2948,In_1565,In_2629);
nand U2949 (N_2949,In_292,In_1101);
or U2950 (N_2950,In_1206,In_559);
nor U2951 (N_2951,In_1551,In_163);
nor U2952 (N_2952,In_2438,In_2930);
and U2953 (N_2953,In_2820,In_1605);
or U2954 (N_2954,In_329,In_2168);
or U2955 (N_2955,In_2259,In_676);
nor U2956 (N_2956,In_1961,In_2693);
or U2957 (N_2957,In_586,In_205);
nor U2958 (N_2958,In_1117,In_2920);
nand U2959 (N_2959,In_1302,In_2363);
xnor U2960 (N_2960,In_1401,In_119);
or U2961 (N_2961,In_2266,In_854);
nor U2962 (N_2962,In_2539,In_2947);
nand U2963 (N_2963,In_816,In_1816);
or U2964 (N_2964,In_630,In_1037);
xor U2965 (N_2965,In_1409,In_1226);
nand U2966 (N_2966,In_2080,In_998);
or U2967 (N_2967,In_2098,In_1616);
or U2968 (N_2968,In_1301,In_1295);
or U2969 (N_2969,In_1873,In_17);
and U2970 (N_2970,In_1264,In_2715);
and U2971 (N_2971,In_514,In_2706);
xnor U2972 (N_2972,In_721,In_1452);
and U2973 (N_2973,In_1098,In_197);
or U2974 (N_2974,In_1049,In_1299);
nand U2975 (N_2975,In_86,In_2969);
nand U2976 (N_2976,In_604,In_2367);
nor U2977 (N_2977,In_200,In_998);
nor U2978 (N_2978,In_340,In_2195);
or U2979 (N_2979,In_1047,In_2528);
and U2980 (N_2980,In_2978,In_2429);
nor U2981 (N_2981,In_1203,In_2992);
nand U2982 (N_2982,In_2509,In_1485);
xnor U2983 (N_2983,In_2504,In_1081);
or U2984 (N_2984,In_2652,In_176);
nor U2985 (N_2985,In_1257,In_1224);
nand U2986 (N_2986,In_1522,In_2770);
xnor U2987 (N_2987,In_1362,In_416);
nor U2988 (N_2988,In_757,In_1);
nand U2989 (N_2989,In_2542,In_1481);
and U2990 (N_2990,In_198,In_2134);
nand U2991 (N_2991,In_207,In_1);
nand U2992 (N_2992,In_764,In_1264);
nand U2993 (N_2993,In_2774,In_2676);
nand U2994 (N_2994,In_268,In_676);
nand U2995 (N_2995,In_2741,In_2402);
and U2996 (N_2996,In_1435,In_2305);
and U2997 (N_2997,In_1532,In_2256);
and U2998 (N_2998,In_1320,In_2849);
nor U2999 (N_2999,In_1153,In_1455);
and U3000 (N_3000,N_1424,N_1307);
xor U3001 (N_3001,N_2253,N_174);
or U3002 (N_3002,N_436,N_87);
or U3003 (N_3003,N_2462,N_2020);
and U3004 (N_3004,N_1443,N_543);
nor U3005 (N_3005,N_2074,N_2841);
xnor U3006 (N_3006,N_2983,N_1556);
and U3007 (N_3007,N_2380,N_1516);
nand U3008 (N_3008,N_253,N_729);
nor U3009 (N_3009,N_1731,N_1056);
and U3010 (N_3010,N_2732,N_1266);
or U3011 (N_3011,N_434,N_2252);
nor U3012 (N_3012,N_2338,N_566);
nor U3013 (N_3013,N_760,N_476);
nand U3014 (N_3014,N_1471,N_1198);
nand U3015 (N_3015,N_377,N_275);
or U3016 (N_3016,N_1296,N_1798);
or U3017 (N_3017,N_2586,N_722);
nand U3018 (N_3018,N_900,N_1292);
xor U3019 (N_3019,N_1553,N_1338);
and U3020 (N_3020,N_256,N_955);
or U3021 (N_3021,N_331,N_1495);
xor U3022 (N_3022,N_2613,N_2755);
nand U3023 (N_3023,N_2765,N_1470);
and U3024 (N_3024,N_1789,N_1919);
xnor U3025 (N_3025,N_2153,N_540);
nor U3026 (N_3026,N_724,N_1813);
nand U3027 (N_3027,N_136,N_2690);
and U3028 (N_3028,N_1468,N_2349);
nor U3029 (N_3029,N_134,N_2161);
nand U3030 (N_3030,N_672,N_107);
or U3031 (N_3031,N_718,N_2618);
and U3032 (N_3032,N_1230,N_804);
and U3033 (N_3033,N_1535,N_1854);
xnor U3034 (N_3034,N_2577,N_2470);
nand U3035 (N_3035,N_319,N_2762);
or U3036 (N_3036,N_2857,N_499);
nand U3037 (N_3037,N_2775,N_2715);
nand U3038 (N_3038,N_2193,N_1106);
or U3039 (N_3039,N_647,N_2474);
nor U3040 (N_3040,N_2124,N_1765);
nand U3041 (N_3041,N_465,N_1833);
or U3042 (N_3042,N_2482,N_439);
nand U3043 (N_3043,N_2754,N_2967);
nor U3044 (N_3044,N_2977,N_1145);
nor U3045 (N_3045,N_1025,N_770);
nand U3046 (N_3046,N_2522,N_1687);
nor U3047 (N_3047,N_757,N_2900);
or U3048 (N_3048,N_2845,N_2603);
and U3049 (N_3049,N_755,N_385);
nor U3050 (N_3050,N_2230,N_1152);
nor U3051 (N_3051,N_1206,N_297);
xor U3052 (N_3052,N_1707,N_1805);
or U3053 (N_3053,N_1140,N_1771);
and U3054 (N_3054,N_2363,N_2733);
nand U3055 (N_3055,N_151,N_1825);
nand U3056 (N_3056,N_621,N_1628);
and U3057 (N_3057,N_2808,N_2739);
nor U3058 (N_3058,N_2557,N_2449);
and U3059 (N_3059,N_1204,N_2578);
xnor U3060 (N_3060,N_656,N_166);
or U3061 (N_3061,N_2146,N_1255);
xnor U3062 (N_3062,N_667,N_2759);
and U3063 (N_3063,N_1908,N_1399);
xor U3064 (N_3064,N_2095,N_2552);
nand U3065 (N_3065,N_1984,N_2781);
or U3066 (N_3066,N_2719,N_1112);
nand U3067 (N_3067,N_740,N_2285);
nand U3068 (N_3068,N_1316,N_603);
nand U3069 (N_3069,N_1555,N_913);
nand U3070 (N_3070,N_2394,N_492);
and U3071 (N_3071,N_2378,N_1077);
nand U3072 (N_3072,N_576,N_2937);
nor U3073 (N_3073,N_141,N_1856);
or U3074 (N_3074,N_850,N_2620);
or U3075 (N_3075,N_1490,N_1462);
xnor U3076 (N_3076,N_514,N_2897);
nor U3077 (N_3077,N_1937,N_2676);
and U3078 (N_3078,N_1018,N_2495);
or U3079 (N_3079,N_985,N_184);
nand U3080 (N_3080,N_1498,N_649);
nor U3081 (N_3081,N_2393,N_1530);
nor U3082 (N_3082,N_2602,N_623);
and U3083 (N_3083,N_628,N_948);
xor U3084 (N_3084,N_869,N_2617);
and U3085 (N_3085,N_1743,N_1549);
and U3086 (N_3086,N_2023,N_1181);
xor U3087 (N_3087,N_1836,N_693);
nand U3088 (N_3088,N_844,N_2869);
xnor U3089 (N_3089,N_2718,N_1171);
nor U3090 (N_3090,N_1218,N_2880);
nand U3091 (N_3091,N_1941,N_2274);
nand U3092 (N_3092,N_1285,N_1269);
or U3093 (N_3093,N_2292,N_2228);
nand U3094 (N_3094,N_705,N_1815);
xor U3095 (N_3095,N_1527,N_2695);
or U3096 (N_3096,N_202,N_455);
and U3097 (N_3097,N_2863,N_2913);
nand U3098 (N_3098,N_1958,N_1184);
and U3099 (N_3099,N_2984,N_2317);
nor U3100 (N_3100,N_2486,N_1943);
or U3101 (N_3101,N_2717,N_83);
or U3102 (N_3102,N_1007,N_1410);
and U3103 (N_3103,N_1922,N_76);
and U3104 (N_3104,N_165,N_1475);
nand U3105 (N_3105,N_1416,N_2300);
nor U3106 (N_3106,N_1273,N_1890);
nor U3107 (N_3107,N_680,N_2288);
nor U3108 (N_3108,N_375,N_1483);
nand U3109 (N_3109,N_1863,N_735);
nor U3110 (N_3110,N_2390,N_824);
and U3111 (N_3111,N_673,N_2737);
or U3112 (N_3112,N_283,N_925);
and U3113 (N_3113,N_192,N_951);
nand U3114 (N_3114,N_2981,N_1658);
nand U3115 (N_3115,N_2409,N_1760);
nand U3116 (N_3116,N_2017,N_50);
xnor U3117 (N_3117,N_2953,N_1810);
or U3118 (N_3118,N_2121,N_1622);
nor U3119 (N_3119,N_1178,N_1644);
nand U3120 (N_3120,N_1076,N_753);
nor U3121 (N_3121,N_2885,N_1721);
or U3122 (N_3122,N_1071,N_2669);
nor U3123 (N_3123,N_2314,N_677);
nand U3124 (N_3124,N_2558,N_2091);
or U3125 (N_3125,N_82,N_2960);
nand U3126 (N_3126,N_922,N_641);
or U3127 (N_3127,N_205,N_2145);
nor U3128 (N_3128,N_1221,N_2432);
and U3129 (N_3129,N_1795,N_289);
nor U3130 (N_3130,N_1068,N_1092);
nor U3131 (N_3131,N_128,N_1869);
xor U3132 (N_3132,N_1915,N_935);
nand U3133 (N_3133,N_2233,N_1405);
or U3134 (N_3134,N_2174,N_62);
and U3135 (N_3135,N_1615,N_703);
nand U3136 (N_3136,N_1818,N_1010);
nor U3137 (N_3137,N_1695,N_1380);
nand U3138 (N_3138,N_2851,N_1492);
or U3139 (N_3139,N_734,N_339);
nor U3140 (N_3140,N_2659,N_1754);
nor U3141 (N_3141,N_1261,N_388);
and U3142 (N_3142,N_1084,N_247);
xor U3143 (N_3143,N_405,N_2853);
nor U3144 (N_3144,N_1747,N_191);
or U3145 (N_3145,N_1662,N_1752);
nor U3146 (N_3146,N_322,N_1790);
and U3147 (N_3147,N_2211,N_1169);
nand U3148 (N_3148,N_20,N_1602);
or U3149 (N_3149,N_2912,N_343);
and U3150 (N_3150,N_1668,N_961);
and U3151 (N_3151,N_493,N_1050);
nand U3152 (N_3152,N_1618,N_1323);
nand U3153 (N_3153,N_2219,N_2120);
and U3154 (N_3154,N_2569,N_1461);
nor U3155 (N_3155,N_80,N_1716);
or U3156 (N_3156,N_684,N_789);
and U3157 (N_3157,N_2537,N_430);
and U3158 (N_3158,N_944,N_1729);
or U3159 (N_3159,N_1609,N_2525);
or U3160 (N_3160,N_2599,N_2660);
xnor U3161 (N_3161,N_1271,N_611);
nor U3162 (N_3162,N_497,N_538);
xnor U3163 (N_3163,N_2591,N_84);
nor U3164 (N_3164,N_369,N_125);
nand U3165 (N_3165,N_148,N_2753);
nor U3166 (N_3166,N_2673,N_409);
nor U3167 (N_3167,N_2177,N_367);
nor U3168 (N_3168,N_2867,N_1256);
nand U3169 (N_3169,N_237,N_1481);
nor U3170 (N_3170,N_1087,N_1038);
nand U3171 (N_3171,N_2128,N_433);
and U3172 (N_3172,N_494,N_2928);
nand U3173 (N_3173,N_691,N_217);
and U3174 (N_3174,N_17,N_220);
nand U3175 (N_3175,N_173,N_2055);
nand U3176 (N_3176,N_2479,N_1375);
or U3177 (N_3177,N_2582,N_1748);
nor U3178 (N_3178,N_144,N_2011);
or U3179 (N_3179,N_2802,N_408);
and U3180 (N_3180,N_2090,N_1196);
and U3181 (N_3181,N_2117,N_301);
nand U3182 (N_3182,N_481,N_2284);
xor U3183 (N_3183,N_2678,N_1792);
nand U3184 (N_3184,N_2903,N_1965);
nor U3185 (N_3185,N_2226,N_241);
nor U3186 (N_3186,N_2901,N_2614);
nand U3187 (N_3187,N_1186,N_1193);
nand U3188 (N_3188,N_599,N_1816);
or U3189 (N_3189,N_1796,N_459);
or U3190 (N_3190,N_2748,N_2439);
nor U3191 (N_3191,N_1175,N_2447);
nand U3192 (N_3192,N_1939,N_391);
or U3193 (N_3193,N_2675,N_1598);
or U3194 (N_3194,N_1572,N_1121);
nor U3195 (N_3195,N_2823,N_577);
nor U3196 (N_3196,N_2371,N_1217);
and U3197 (N_3197,N_2631,N_1001);
and U3198 (N_3198,N_1868,N_2076);
or U3199 (N_3199,N_867,N_912);
nor U3200 (N_3200,N_618,N_1688);
nand U3201 (N_3201,N_1243,N_1069);
xnor U3202 (N_3202,N_1964,N_2255);
nor U3203 (N_3203,N_1968,N_969);
nand U3204 (N_3204,N_402,N_2952);
nor U3205 (N_3205,N_2195,N_2429);
or U3206 (N_3206,N_1061,N_1903);
xor U3207 (N_3207,N_1433,N_1096);
or U3208 (N_3208,N_257,N_2339);
nor U3209 (N_3209,N_2012,N_1111);
or U3210 (N_3210,N_449,N_742);
nor U3211 (N_3211,N_198,N_114);
nor U3212 (N_3212,N_1860,N_609);
nand U3213 (N_3213,N_2248,N_209);
nor U3214 (N_3214,N_314,N_346);
nand U3215 (N_3215,N_1673,N_194);
and U3216 (N_3216,N_490,N_2163);
nand U3217 (N_3217,N_2059,N_1710);
nand U3218 (N_3218,N_918,N_336);
or U3219 (N_3219,N_1918,N_2081);
nand U3220 (N_3220,N_966,N_1788);
nand U3221 (N_3221,N_2794,N_613);
nand U3222 (N_3222,N_2351,N_467);
and U3223 (N_3223,N_1513,N_57);
nand U3224 (N_3224,N_751,N_2914);
nand U3225 (N_3225,N_1130,N_1322);
xor U3226 (N_3226,N_61,N_2037);
nand U3227 (N_3227,N_1843,N_1222);
or U3228 (N_3228,N_120,N_1613);
nand U3229 (N_3229,N_1737,N_2107);
or U3230 (N_3230,N_2819,N_2511);
nand U3231 (N_3231,N_262,N_2746);
or U3232 (N_3232,N_1547,N_2624);
or U3233 (N_3233,N_1913,N_2144);
nor U3234 (N_3234,N_2742,N_1460);
or U3235 (N_3235,N_2308,N_728);
or U3236 (N_3236,N_2548,N_2041);
xnor U3237 (N_3237,N_2457,N_2600);
nor U3238 (N_3238,N_2353,N_999);
nand U3239 (N_3239,N_1957,N_1544);
nand U3240 (N_3240,N_2365,N_2000);
nand U3241 (N_3241,N_715,N_967);
and U3242 (N_3242,N_2609,N_1328);
and U3243 (N_3243,N_118,N_2435);
or U3244 (N_3244,N_2467,N_323);
nor U3245 (N_3245,N_1717,N_517);
or U3246 (N_3246,N_658,N_332);
nor U3247 (N_3247,N_2088,N_2372);
or U3248 (N_3248,N_326,N_2042);
xor U3249 (N_3249,N_1144,N_477);
xnor U3250 (N_3250,N_2369,N_934);
nand U3251 (N_3251,N_2889,N_2553);
or U3252 (N_3252,N_636,N_2818);
or U3253 (N_3253,N_2420,N_102);
and U3254 (N_3254,N_203,N_115);
and U3255 (N_3255,N_2347,N_1037);
and U3256 (N_3256,N_1146,N_424);
and U3257 (N_3257,N_1054,N_731);
or U3258 (N_3258,N_78,N_1368);
and U3259 (N_3259,N_2151,N_2422);
nand U3260 (N_3260,N_2519,N_2157);
and U3261 (N_3261,N_460,N_56);
nand U3262 (N_3262,N_2661,N_2871);
nand U3263 (N_3263,N_1436,N_1304);
nand U3264 (N_3264,N_2979,N_721);
or U3265 (N_3265,N_1298,N_1259);
or U3266 (N_3266,N_2374,N_2260);
nand U3267 (N_3267,N_2738,N_897);
nor U3268 (N_3268,N_612,N_1015);
and U3269 (N_3269,N_792,N_2813);
xnor U3270 (N_3270,N_608,N_2384);
or U3271 (N_3271,N_1314,N_726);
nor U3272 (N_3272,N_1905,N_905);
xor U3273 (N_3273,N_504,N_233);
or U3274 (N_3274,N_1596,N_988);
or U3275 (N_3275,N_2969,N_875);
and U3276 (N_3276,N_2777,N_2433);
nor U3277 (N_3277,N_1697,N_315);
nor U3278 (N_3278,N_525,N_2298);
nor U3279 (N_3279,N_2635,N_2683);
or U3280 (N_3280,N_1987,N_1227);
or U3281 (N_3281,N_2924,N_1728);
or U3282 (N_3282,N_547,N_1923);
and U3283 (N_3283,N_2080,N_2412);
xor U3284 (N_3284,N_2509,N_2968);
nor U3285 (N_3285,N_1751,N_1078);
xnor U3286 (N_3286,N_710,N_2050);
nand U3287 (N_3287,N_55,N_2139);
or U3288 (N_3288,N_2749,N_1998);
nand U3289 (N_3289,N_363,N_2580);
or U3290 (N_3290,N_555,N_2879);
and U3291 (N_3291,N_1701,N_1866);
or U3292 (N_3292,N_725,N_129);
nand U3293 (N_3293,N_978,N_1280);
nor U3294 (N_3294,N_1637,N_2465);
nor U3295 (N_3295,N_437,N_630);
and U3296 (N_3296,N_2442,N_2698);
and U3297 (N_3297,N_1875,N_2408);
or U3298 (N_3298,N_1525,N_463);
and U3299 (N_3299,N_1125,N_238);
xnor U3300 (N_3300,N_1288,N_99);
or U3301 (N_3301,N_2576,N_235);
or U3302 (N_3302,N_1422,N_1778);
xor U3303 (N_3303,N_2103,N_2450);
or U3304 (N_3304,N_2865,N_561);
and U3305 (N_3305,N_2181,N_1999);
nand U3306 (N_3306,N_907,N_643);
or U3307 (N_3307,N_806,N_2971);
and U3308 (N_3308,N_1826,N_327);
and U3309 (N_3309,N_2844,N_1299);
nor U3310 (N_3310,N_534,N_505);
and U3311 (N_3311,N_2957,N_733);
nand U3312 (N_3312,N_2533,N_1774);
and U3313 (N_3313,N_1254,N_840);
nand U3314 (N_3314,N_968,N_832);
or U3315 (N_3315,N_1270,N_1333);
or U3316 (N_3316,N_1750,N_2658);
and U3317 (N_3317,N_1772,N_1168);
nor U3318 (N_3318,N_2123,N_963);
xor U3319 (N_3319,N_898,N_2373);
nand U3320 (N_3320,N_2268,N_1372);
or U3321 (N_3321,N_139,N_1783);
and U3322 (N_3322,N_226,N_2206);
nor U3323 (N_3323,N_939,N_269);
nand U3324 (N_3324,N_373,N_744);
nor U3325 (N_3325,N_2136,N_172);
nand U3326 (N_3326,N_154,N_8);
nor U3327 (N_3327,N_364,N_2598);
or U3328 (N_3328,N_2478,N_1253);
nor U3329 (N_3329,N_2152,N_1847);
xor U3330 (N_3330,N_2313,N_271);
nand U3331 (N_3331,N_51,N_777);
xnor U3332 (N_3332,N_2119,N_2352);
xnor U3333 (N_3333,N_2856,N_97);
xnor U3334 (N_3334,N_2705,N_96);
and U3335 (N_3335,N_140,N_2238);
nand U3336 (N_3336,N_952,N_2938);
or U3337 (N_3337,N_2187,N_417);
nor U3338 (N_3338,N_1429,N_2007);
nand U3339 (N_3339,N_193,N_1088);
xor U3340 (N_3340,N_2305,N_2054);
nand U3341 (N_3341,N_1441,N_916);
nand U3342 (N_3342,N_2263,N_1862);
nor U3343 (N_3343,N_1009,N_1369);
nor U3344 (N_3344,N_1411,N_1502);
nor U3345 (N_3345,N_531,N_1766);
or U3346 (N_3346,N_1289,N_1741);
nand U3347 (N_3347,N_1265,N_654);
nor U3348 (N_3348,N_2048,N_2480);
or U3349 (N_3349,N_2484,N_941);
nor U3350 (N_3350,N_2512,N_1839);
nor U3351 (N_3351,N_2492,N_2743);
nand U3352 (N_3352,N_1714,N_2350);
xnor U3353 (N_3353,N_1366,N_1013);
xor U3354 (N_3354,N_1419,N_2677);
nand U3355 (N_3355,N_774,N_2340);
nand U3356 (N_3356,N_594,N_2791);
nand U3357 (N_3357,N_1402,N_484);
and U3358 (N_3358,N_60,N_1887);
nand U3359 (N_3359,N_1925,N_182);
and U3360 (N_3360,N_622,N_568);
xnor U3361 (N_3361,N_1491,N_2406);
or U3362 (N_3362,N_42,N_2655);
and U3363 (N_3363,N_1955,N_1749);
nor U3364 (N_3364,N_1725,N_2415);
nand U3365 (N_3365,N_2544,N_2584);
nand U3366 (N_3366,N_1075,N_2710);
and U3367 (N_3367,N_590,N_579);
nand U3368 (N_3368,N_1867,N_1157);
nand U3369 (N_3369,N_2684,N_591);
and U3370 (N_3370,N_2212,N_360);
nand U3371 (N_3371,N_1129,N_2421);
or U3372 (N_3372,N_983,N_1344);
nor U3373 (N_3373,N_1480,N_227);
xor U3374 (N_3374,N_1699,N_1006);
nor U3375 (N_3375,N_1359,N_1019);
nor U3376 (N_3376,N_666,N_2555);
xnor U3377 (N_3377,N_23,N_1407);
xnor U3378 (N_3378,N_2196,N_1542);
and U3379 (N_3379,N_2418,N_2273);
or U3380 (N_3380,N_1983,N_454);
nand U3381 (N_3381,N_18,N_1324);
nand U3382 (N_3382,N_117,N_2197);
nand U3383 (N_3383,N_2639,N_1016);
nor U3384 (N_3384,N_2280,N_697);
or U3385 (N_3385,N_1336,N_2164);
or U3386 (N_3386,N_2108,N_817);
nand U3387 (N_3387,N_2809,N_1028);
nand U3388 (N_3388,N_1924,N_1967);
or U3389 (N_3389,N_746,N_583);
xor U3390 (N_3390,N_2590,N_2815);
xor U3391 (N_3391,N_2905,N_2361);
nor U3392 (N_3392,N_2930,N_2670);
nand U3393 (N_3393,N_426,N_2391);
nand U3394 (N_3394,N_1235,N_244);
and U3395 (N_3395,N_1512,N_1817);
nand U3396 (N_3396,N_2927,N_1293);
nand U3397 (N_3397,N_2239,N_1108);
nor U3398 (N_3398,N_2225,N_975);
or U3399 (N_3399,N_2060,N_2083);
or U3400 (N_3400,N_48,N_808);
and U3401 (N_3401,N_485,N_1200);
and U3402 (N_3402,N_1312,N_340);
nor U3403 (N_3403,N_1430,N_2860);
or U3404 (N_3404,N_2534,N_2650);
and U3405 (N_3405,N_876,N_1962);
and U3406 (N_3406,N_2199,N_2807);
xnor U3407 (N_3407,N_27,N_535);
nor U3408 (N_3408,N_15,N_1489);
nand U3409 (N_3409,N_2965,N_1666);
and U3410 (N_3410,N_111,N_1985);
or U3411 (N_3411,N_2499,N_536);
and U3412 (N_3412,N_1238,N_2862);
xnor U3413 (N_3413,N_903,N_1570);
and U3414 (N_3414,N_2277,N_1397);
nor U3415 (N_3415,N_36,N_1199);
or U3416 (N_3416,N_2043,N_2475);
nand U3417 (N_3417,N_234,N_372);
and U3418 (N_3418,N_2357,N_355);
or U3419 (N_3419,N_1275,N_601);
and U3420 (N_3420,N_2382,N_44);
and U3421 (N_3421,N_2730,N_1494);
nor U3422 (N_3422,N_1352,N_163);
or U3423 (N_3423,N_468,N_736);
and U3424 (N_3424,N_1676,N_1248);
and U3425 (N_3425,N_2049,N_2720);
or U3426 (N_3426,N_981,N_2162);
nand U3427 (N_3427,N_769,N_940);
and U3428 (N_3428,N_1724,N_2192);
nor U3429 (N_3429,N_826,N_629);
or U3430 (N_3430,N_210,N_1386);
xor U3431 (N_3431,N_1354,N_2874);
nand U3432 (N_3432,N_1486,N_1537);
xnor U3433 (N_3433,N_2521,N_1095);
nor U3434 (N_3434,N_2140,N_785);
nand U3435 (N_3435,N_116,N_2220);
or U3436 (N_3436,N_807,N_2915);
nand U3437 (N_3437,N_610,N_32);
nand U3438 (N_3438,N_2191,N_1382);
and U3439 (N_3439,N_358,N_486);
and U3440 (N_3440,N_2697,N_1305);
nand U3441 (N_3441,N_1807,N_2771);
and U3442 (N_3442,N_1963,N_1723);
nand U3443 (N_3443,N_2626,N_906);
and U3444 (N_3444,N_187,N_278);
and U3445 (N_3445,N_52,N_2888);
and U3446 (N_3446,N_1727,N_2198);
nand U3447 (N_3447,N_124,N_1864);
or U3448 (N_3448,N_2535,N_2311);
nand U3449 (N_3449,N_1584,N_2579);
and U3450 (N_3450,N_1361,N_425);
and U3451 (N_3451,N_545,N_881);
or U3452 (N_3452,N_598,N_1024);
and U3453 (N_3453,N_990,N_526);
xor U3454 (N_3454,N_394,N_2891);
and U3455 (N_3455,N_2032,N_2894);
xnor U3456 (N_3456,N_2346,N_1646);
xnor U3457 (N_3457,N_2837,N_2096);
and U3458 (N_3458,N_2256,N_674);
or U3459 (N_3459,N_1309,N_1708);
and U3460 (N_3460,N_2118,N_1538);
or U3461 (N_3461,N_67,N_665);
and U3462 (N_3462,N_904,N_1091);
xor U3463 (N_3463,N_280,N_1260);
or U3464 (N_3464,N_1745,N_313);
and U3465 (N_3465,N_1995,N_14);
xor U3466 (N_3466,N_644,N_970);
or U3467 (N_3467,N_100,N_2185);
and U3468 (N_3468,N_1651,N_469);
xor U3469 (N_3469,N_720,N_2736);
nor U3470 (N_3470,N_783,N_2234);
nand U3471 (N_3471,N_2240,N_1906);
nor U3472 (N_3472,N_2179,N_1842);
and U3473 (N_3473,N_2942,N_1225);
nor U3474 (N_3474,N_1877,N_1563);
and U3475 (N_3475,N_2817,N_1661);
nand U3476 (N_3476,N_788,N_1488);
and U3477 (N_3477,N_2471,N_201);
and U3478 (N_3478,N_130,N_650);
nor U3479 (N_3479,N_683,N_1000);
and U3480 (N_3480,N_2079,N_2321);
nor U3481 (N_3481,N_1902,N_65);
nor U3482 (N_3482,N_2377,N_2150);
and U3483 (N_3483,N_1326,N_716);
and U3484 (N_3484,N_871,N_2821);
and U3485 (N_3485,N_2345,N_2038);
or U3486 (N_3486,N_2072,N_2434);
and U3487 (N_3487,N_2805,N_2806);
xnor U3488 (N_3488,N_518,N_94);
and U3489 (N_3489,N_635,N_1632);
or U3490 (N_3490,N_2703,N_2488);
or U3491 (N_3491,N_634,N_1051);
or U3492 (N_3492,N_2975,N_1073);
nand U3493 (N_3493,N_2543,N_150);
nor U3494 (N_3494,N_40,N_606);
nand U3495 (N_3495,N_1365,N_1374);
nand U3496 (N_3496,N_800,N_895);
or U3497 (N_3497,N_1927,N_1767);
or U3498 (N_3498,N_2637,N_1210);
nand U3499 (N_3499,N_2419,N_521);
and U3500 (N_3500,N_466,N_1466);
and U3501 (N_3501,N_213,N_1994);
nor U3502 (N_3502,N_564,N_2796);
nor U3503 (N_3503,N_2445,N_1319);
nand U3504 (N_3504,N_528,N_2583);
nand U3505 (N_3505,N_1916,N_2241);
or U3506 (N_3506,N_2254,N_1440);
nand U3507 (N_3507,N_2142,N_2362);
and U3508 (N_3508,N_2662,N_1231);
nor U3509 (N_3509,N_79,N_333);
and U3510 (N_3510,N_37,N_393);
or U3511 (N_3511,N_550,N_1347);
nor U3512 (N_3512,N_822,N_1601);
and U3513 (N_3513,N_1396,N_2295);
nor U3514 (N_3514,N_664,N_2704);
xnor U3515 (N_3515,N_1041,N_2638);
and U3516 (N_3516,N_2396,N_1127);
nor U3517 (N_3517,N_361,N_197);
nand U3518 (N_3518,N_1464,N_669);
nand U3519 (N_3519,N_1712,N_2461);
nor U3520 (N_3520,N_95,N_2058);
or U3521 (N_3521,N_567,N_1606);
nand U3522 (N_3522,N_614,N_1684);
nand U3523 (N_3523,N_767,N_563);
or U3524 (N_3524,N_2788,N_1715);
nor U3525 (N_3525,N_1294,N_414);
and U3526 (N_3526,N_1039,N_1938);
and U3527 (N_3527,N_1138,N_295);
xnor U3528 (N_3528,N_1616,N_1510);
nor U3529 (N_3529,N_1047,N_132);
nand U3530 (N_3530,N_1590,N_1340);
xnor U3531 (N_3531,N_272,N_1586);
nand U3532 (N_3532,N_229,N_2031);
xnor U3533 (N_3533,N_1428,N_1446);
or U3534 (N_3534,N_2368,N_380);
and U3535 (N_3535,N_1501,N_763);
nand U3536 (N_3536,N_1873,N_575);
nand U3537 (N_3537,N_997,N_2632);
nor U3538 (N_3538,N_453,N_1652);
xnor U3539 (N_3539,N_239,N_2100);
and U3540 (N_3540,N_2708,N_2886);
nand U3541 (N_3541,N_2798,N_1636);
nand U3542 (N_3542,N_1020,N_1614);
nand U3543 (N_3543,N_2324,N_321);
nor U3544 (N_3544,N_1733,N_159);
nor U3545 (N_3545,N_2604,N_2834);
and U3546 (N_3546,N_1786,N_1315);
or U3547 (N_3547,N_1581,N_2998);
and U3548 (N_3548,N_2711,N_882);
and U3549 (N_3549,N_1976,N_1508);
and U3550 (N_3550,N_70,N_1678);
nor U3551 (N_3551,N_2158,N_556);
nor U3552 (N_3552,N_2878,N_2870);
and U3553 (N_3553,N_1978,N_998);
xor U3554 (N_3554,N_548,N_2890);
xnor U3555 (N_3555,N_1002,N_937);
and U3556 (N_3556,N_2811,N_2294);
and U3557 (N_3557,N_2320,N_286);
nand U3558 (N_3558,N_2884,N_2858);
nand U3559 (N_3559,N_345,N_1300);
nand U3560 (N_3560,N_2940,N_1165);
xnor U3561 (N_3561,N_709,N_1625);
or U3562 (N_3562,N_1511,N_831);
xnor U3563 (N_3563,N_1233,N_2877);
xnor U3564 (N_3564,N_1763,N_1577);
nor U3565 (N_3565,N_1702,N_640);
nand U3566 (N_3566,N_480,N_862);
and U3567 (N_3567,N_977,N_330);
nand U3568 (N_3568,N_1355,N_2908);
nand U3569 (N_3569,N_2015,N_2652);
or U3570 (N_3570,N_1879,N_2898);
nand U3571 (N_3571,N_2987,N_1297);
or U3572 (N_3572,N_2504,N_415);
xor U3573 (N_3573,N_2948,N_2820);
or U3574 (N_3574,N_863,N_1610);
and U3575 (N_3575,N_2751,N_1162);
and U3576 (N_3576,N_1485,N_2355);
nand U3577 (N_3577,N_1690,N_1031);
and U3578 (N_3578,N_701,N_2116);
nor U3579 (N_3579,N_1286,N_2171);
or U3580 (N_3580,N_1738,N_1450);
and U3581 (N_3581,N_342,N_2105);
or U3582 (N_3582,N_341,N_741);
nand U3583 (N_3583,N_1996,N_1705);
nor U3584 (N_3584,N_368,N_2190);
and U3585 (N_3585,N_1263,N_1560);
xnor U3586 (N_3586,N_1654,N_1022);
nand U3587 (N_3587,N_1981,N_829);
nor U3588 (N_3588,N_2246,N_676);
nor U3589 (N_3589,N_153,N_1418);
and U3590 (N_3590,N_2358,N_799);
or U3591 (N_3591,N_929,N_383);
and U3592 (N_3592,N_2089,N_2651);
or U3593 (N_3593,N_1412,N_255);
nor U3594 (N_3594,N_2726,N_791);
xnor U3595 (N_3595,N_809,N_1401);
nand U3596 (N_3596,N_1043,N_761);
nor U3597 (N_3597,N_2148,N_1620);
or U3598 (N_3598,N_1952,N_2082);
xor U3599 (N_3599,N_2131,N_1809);
or U3600 (N_3600,N_2530,N_651);
nor U3601 (N_3601,N_2170,N_1770);
and U3602 (N_3602,N_1629,N_508);
and U3603 (N_3603,N_2341,N_1706);
nor U3604 (N_3604,N_58,N_81);
nor U3605 (N_3605,N_795,N_2178);
or U3606 (N_3606,N_1384,N_53);
nand U3607 (N_3607,N_243,N_2776);
nand U3608 (N_3608,N_2656,N_932);
nand U3609 (N_3609,N_2264,N_856);
and U3610 (N_3610,N_2567,N_1624);
and U3611 (N_3611,N_1546,N_1947);
nand U3612 (N_3612,N_1914,N_2056);
and U3613 (N_3613,N_1518,N_1313);
or U3614 (N_3614,N_747,N_2956);
nand U3615 (N_3615,N_1852,N_1268);
and U3616 (N_3616,N_1400,N_113);
or U3617 (N_3617,N_207,N_146);
and U3618 (N_3618,N_2682,N_407);
xor U3619 (N_3619,N_989,N_1819);
and U3620 (N_3620,N_230,N_2400);
nand U3621 (N_3621,N_7,N_902);
xnor U3622 (N_3622,N_2165,N_2114);
and U3623 (N_3623,N_382,N_980);
nor U3624 (N_3624,N_179,N_570);
nor U3625 (N_3625,N_2612,N_1659);
nand U3626 (N_3626,N_2934,N_936);
nor U3627 (N_3627,N_2279,N_2184);
nor U3628 (N_3628,N_1592,N_2619);
and U3629 (N_3629,N_9,N_1150);
nand U3630 (N_3630,N_274,N_1761);
and U3631 (N_3631,N_2030,N_2539);
nand U3632 (N_3632,N_1214,N_1302);
nand U3633 (N_3633,N_261,N_1437);
or U3634 (N_3634,N_631,N_745);
nor U3635 (N_3635,N_2014,N_1497);
or U3636 (N_3636,N_1250,N_1281);
nor U3637 (N_3637,N_2574,N_1665);
or U3638 (N_3638,N_2565,N_743);
nand U3639 (N_3639,N_2920,N_551);
nor U3640 (N_3640,N_211,N_2291);
or U3641 (N_3641,N_2303,N_1189);
and U3642 (N_3642,N_2787,N_2018);
xor U3643 (N_3643,N_1830,N_1387);
nand U3644 (N_3644,N_571,N_1979);
nand U3645 (N_3645,N_1246,N_2126);
nand U3646 (N_3646,N_1201,N_927);
nor U3647 (N_3647,N_2500,N_2770);
xor U3648 (N_3648,N_1378,N_2232);
or U3649 (N_3649,N_2127,N_2563);
xor U3650 (N_3650,N_1454,N_507);
nand U3651 (N_3651,N_1824,N_1893);
nor U3652 (N_3652,N_711,N_752);
nand U3653 (N_3653,N_2344,N_2911);
and U3654 (N_3654,N_189,N_1226);
or U3655 (N_3655,N_2297,N_419);
xor U3656 (N_3656,N_1070,N_1655);
and U3657 (N_3657,N_1109,N_1917);
nand U3658 (N_3658,N_2271,N_1931);
or U3659 (N_3659,N_2910,N_1012);
nand U3660 (N_3660,N_2554,N_2974);
nor U3661 (N_3661,N_830,N_2648);
or U3662 (N_3662,N_1427,N_356);
and U3663 (N_3663,N_164,N_2287);
nand U3664 (N_3664,N_445,N_63);
and U3665 (N_3665,N_1859,N_85);
and U3666 (N_3666,N_797,N_1083);
and U3667 (N_3667,N_1883,N_1920);
xnor U3668 (N_3668,N_818,N_2073);
and U3669 (N_3669,N_1604,N_304);
and U3670 (N_3670,N_1519,N_422);
nor U3671 (N_3671,N_1154,N_1827);
and U3672 (N_3672,N_2936,N_1696);
nor U3673 (N_3673,N_1787,N_1029);
nand U3674 (N_3674,N_250,N_749);
xnor U3675 (N_3675,N_2803,N_2404);
nor U3676 (N_3676,N_2485,N_1487);
nor U3677 (N_3677,N_2101,N_921);
or U3678 (N_3678,N_1040,N_1899);
nor U3679 (N_3679,N_1638,N_2494);
or U3680 (N_3680,N_2473,N_2545);
nand U3681 (N_3681,N_1974,N_1972);
nand U3682 (N_3682,N_2970,N_600);
or U3683 (N_3683,N_2343,N_885);
or U3684 (N_3684,N_1835,N_2712);
xnor U3685 (N_3685,N_479,N_585);
and U3686 (N_3686,N_2951,N_1257);
nor U3687 (N_3687,N_1909,N_645);
and U3688 (N_3688,N_2949,N_2647);
nand U3689 (N_3689,N_1635,N_1949);
nor U3690 (N_3690,N_1258,N_920);
and U3691 (N_3691,N_1871,N_737);
or U3692 (N_3692,N_2713,N_1228);
or U3693 (N_3693,N_5,N_1482);
and U3694 (N_3694,N_376,N_487);
or U3695 (N_3695,N_2585,N_2700);
nor U3696 (N_3696,N_2601,N_167);
or U3697 (N_3697,N_1432,N_138);
nor U3698 (N_3698,N_2706,N_823);
and U3699 (N_3699,N_738,N_1383);
and U3700 (N_3700,N_780,N_1858);
or U3701 (N_3701,N_1279,N_2999);
or U3702 (N_3702,N_162,N_334);
nor U3703 (N_3703,N_2680,N_1391);
or U3704 (N_3704,N_1642,N_1929);
or U3705 (N_3705,N_1532,N_2825);
or U3706 (N_3706,N_679,N_1837);
and U3707 (N_3707,N_2463,N_2416);
nor U3708 (N_3708,N_2078,N_1828);
and U3709 (N_3709,N_2201,N_2247);
nand U3710 (N_3710,N_589,N_2731);
nand U3711 (N_3711,N_1911,N_2166);
or U3712 (N_3712,N_1643,N_1209);
or U3713 (N_3713,N_1423,N_2481);
or U3714 (N_3714,N_2929,N_604);
nand U3715 (N_3715,N_2431,N_1241);
xor U3716 (N_3716,N_2194,N_1683);
nor U3717 (N_3717,N_1117,N_2026);
or U3718 (N_3718,N_2464,N_837);
xnor U3719 (N_3719,N_59,N_1469);
and U3720 (N_3720,N_2547,N_2945);
or U3721 (N_3721,N_1310,N_2933);
nand U3722 (N_3722,N_2964,N_2559);
xnor U3723 (N_3723,N_1892,N_2002);
nor U3724 (N_3724,N_1398,N_2290);
nand U3725 (N_3725,N_13,N_2180);
and U3726 (N_3726,N_2110,N_593);
and U3727 (N_3727,N_2094,N_1713);
nor U3728 (N_3728,N_2289,N_1948);
nor U3729 (N_3729,N_2070,N_1472);
and U3730 (N_3730,N_412,N_2923);
or U3731 (N_3731,N_958,N_1926);
nor U3732 (N_3732,N_2067,N_2596);
nor U3733 (N_3733,N_2636,N_88);
or U3734 (N_3734,N_2646,N_2996);
nand U3735 (N_3735,N_2995,N_1064);
nand U3736 (N_3736,N_626,N_652);
and U3737 (N_3737,N_387,N_552);
or U3738 (N_3738,N_859,N_2257);
or U3739 (N_3739,N_2672,N_1197);
and U3740 (N_3740,N_686,N_2398);
nand U3741 (N_3741,N_1568,N_1517);
and U3742 (N_3742,N_411,N_1252);
nand U3743 (N_3743,N_1005,N_2909);
xor U3744 (N_3744,N_2438,N_1846);
or U3745 (N_3745,N_1829,N_1139);
and U3746 (N_3746,N_2392,N_282);
or U3747 (N_3747,N_188,N_2780);
or U3748 (N_3748,N_1403,N_1634);
and U3749 (N_3749,N_771,N_303);
and U3750 (N_3750,N_511,N_473);
and U3751 (N_3751,N_798,N_2685);
nand U3752 (N_3752,N_1149,N_878);
nand U3753 (N_3753,N_2542,N_1709);
nand U3754 (N_3754,N_168,N_2946);
or U3755 (N_3755,N_2955,N_1335);
or U3756 (N_3756,N_717,N_103);
and U3757 (N_3757,N_1861,N_1928);
or U3758 (N_3758,N_2593,N_2608);
or U3759 (N_3759,N_1526,N_1036);
and U3760 (N_3760,N_1229,N_2004);
and U3761 (N_3761,N_317,N_979);
and U3762 (N_3762,N_773,N_397);
nor U3763 (N_3763,N_1190,N_1213);
or U3764 (N_3764,N_827,N_2972);
xnor U3765 (N_3765,N_2895,N_1605);
or U3766 (N_3766,N_764,N_1657);
nor U3767 (N_3767,N_1775,N_2573);
nor U3768 (N_3768,N_1574,N_1205);
nand U3769 (N_3769,N_1820,N_1768);
or U3770 (N_3770,N_183,N_973);
nand U3771 (N_3771,N_2529,N_685);
nand U3772 (N_3772,N_2528,N_2309);
and U3773 (N_3773,N_2021,N_143);
xor U3774 (N_3774,N_2506,N_2556);
nand U3775 (N_3775,N_1506,N_2827);
and U3776 (N_3776,N_1496,N_1782);
or U3777 (N_3777,N_778,N_2227);
or U3778 (N_3778,N_1362,N_584);
or U3779 (N_3779,N_1841,N_1379);
and U3780 (N_3780,N_2275,N_305);
or U3781 (N_3781,N_2657,N_588);
or U3782 (N_3782,N_1562,N_803);
nor U3783 (N_3783,N_500,N_11);
nor U3784 (N_3784,N_73,N_1389);
nor U3785 (N_3785,N_2138,N_1026);
nor U3786 (N_3786,N_835,N_1881);
nand U3787 (N_3787,N_2316,N_2978);
or U3788 (N_3788,N_1647,N_2587);
or U3789 (N_3789,N_131,N_1557);
or U3790 (N_3790,N_478,N_2507);
and U3791 (N_3791,N_1934,N_2019);
nand U3792 (N_3792,N_1034,N_510);
and U3793 (N_3793,N_232,N_646);
nor U3794 (N_3794,N_1576,N_2564);
and U3795 (N_3795,N_2186,N_1442);
nand U3796 (N_3796,N_2778,N_1524);
or U3797 (N_3797,N_759,N_438);
or U3798 (N_3798,N_1814,N_627);
nand U3799 (N_3799,N_2962,N_2203);
and U3800 (N_3800,N_231,N_2204);
nor U3801 (N_3801,N_1120,N_2760);
and U3802 (N_3802,N_2850,N_26);
or U3803 (N_3803,N_1477,N_1660);
xnor U3804 (N_3804,N_475,N_2792);
nand U3805 (N_3805,N_199,N_1617);
or U3806 (N_3806,N_527,N_1447);
xnor U3807 (N_3807,N_2882,N_2493);
nor U3808 (N_3808,N_765,N_350);
nor U3809 (N_3809,N_617,N_1182);
xnor U3810 (N_3810,N_1746,N_2109);
and U3811 (N_3811,N_6,N_949);
and U3812 (N_3812,N_30,N_105);
nor U3813 (N_3813,N_2084,N_2052);
nor U3814 (N_3814,N_1325,N_98);
xor U3815 (N_3815,N_1991,N_1891);
and U3816 (N_3816,N_401,N_1528);
or U3817 (N_3817,N_549,N_2622);
and U3818 (N_3818,N_1035,N_1128);
nor U3819 (N_3819,N_1133,N_1803);
and U3820 (N_3820,N_171,N_888);
nand U3821 (N_3821,N_976,N_1504);
and U3822 (N_3822,N_1693,N_756);
nand U3823 (N_3823,N_200,N_2642);
and U3824 (N_3824,N_2976,N_1573);
nor U3825 (N_3825,N_2231,N_1793);
nand U3826 (N_3826,N_1143,N_77);
nor U3827 (N_3827,N_2013,N_1773);
or U3828 (N_3828,N_1066,N_2514);
nand U3829 (N_3829,N_2840,N_1063);
nor U3830 (N_3830,N_2047,N_495);
and U3831 (N_3831,N_2502,N_41);
or U3832 (N_3832,N_865,N_2069);
nand U3833 (N_3833,N_554,N_348);
nand U3834 (N_3834,N_619,N_1329);
nor U3835 (N_3835,N_2643,N_21);
and U3836 (N_3836,N_1160,N_615);
or U3837 (N_3837,N_2606,N_1776);
nor U3838 (N_3838,N_1249,N_596);
or U3839 (N_3839,N_25,N_2010);
nand U3840 (N_3840,N_452,N_2768);
and U3841 (N_3841,N_2904,N_328);
nor U3842 (N_3842,N_2986,N_2896);
and U3843 (N_3843,N_2699,N_883);
nand U3844 (N_3844,N_857,N_1758);
nand U3845 (N_3845,N_2784,N_928);
or U3846 (N_3846,N_2403,N_1435);
nand U3847 (N_3847,N_1669,N_2812);
and U3848 (N_3848,N_24,N_2259);
or U3849 (N_3849,N_1639,N_1583);
or U3850 (N_3850,N_2561,N_2302);
or U3851 (N_3851,N_28,N_2188);
and U3852 (N_3852,N_1912,N_2779);
and U3853 (N_3853,N_638,N_1291);
nand U3854 (N_3854,N_2399,N_1626);
nor U3855 (N_3855,N_775,N_2312);
xor U3856 (N_3856,N_1377,N_1685);
nand U3857 (N_3857,N_1982,N_273);
and U3858 (N_3858,N_2572,N_45);
xor U3859 (N_3859,N_236,N_1534);
nor U3860 (N_3860,N_2527,N_1113);
nand U3861 (N_3861,N_175,N_2892);
or U3862 (N_3862,N_2902,N_894);
or U3863 (N_3863,N_2381,N_1371);
nand U3864 (N_3864,N_2202,N_1671);
nor U3865 (N_3865,N_982,N_2425);
nor U3866 (N_3866,N_251,N_1463);
and U3867 (N_3867,N_249,N_2458);
nand U3868 (N_3868,N_687,N_2941);
nand U3869 (N_3869,N_252,N_784);
nor U3870 (N_3870,N_890,N_1191);
or U3871 (N_3871,N_706,N_1588);
or U3872 (N_3872,N_2918,N_1882);
or U3873 (N_3873,N_1332,N_714);
nand U3874 (N_3874,N_34,N_648);
nand U3875 (N_3875,N_2668,N_964);
nor U3876 (N_3876,N_845,N_1008);
or U3877 (N_3877,N_413,N_2917);
or U3878 (N_3878,N_942,N_1003);
and U3879 (N_3879,N_899,N_2722);
or U3880 (N_3880,N_2707,N_1457);
nor U3881 (N_3881,N_421,N_768);
nand U3882 (N_3882,N_1207,N_2405);
and U3883 (N_3883,N_954,N_2440);
nand U3884 (N_3884,N_260,N_1575);
nor U3885 (N_3885,N_1621,N_2155);
nor U3886 (N_3886,N_2154,N_349);
nand U3887 (N_3887,N_2566,N_1267);
nor U3888 (N_3888,N_2315,N_1308);
or U3889 (N_3889,N_945,N_2286);
nor U3890 (N_3890,N_872,N_1413);
or U3891 (N_3891,N_1719,N_2469);
xnor U3892 (N_3892,N_2866,N_2129);
and U3893 (N_3893,N_1102,N_1910);
nand U3894 (N_3894,N_1124,N_625);
nor U3895 (N_3895,N_75,N_520);
or U3896 (N_3896,N_392,N_2693);
nor U3897 (N_3897,N_2001,N_224);
nand U3898 (N_3898,N_347,N_483);
or U3899 (N_3899,N_698,N_843);
nor U3900 (N_3900,N_2766,N_2854);
nor U3901 (N_3901,N_2848,N_2167);
xor U3902 (N_3902,N_1649,N_2980);
nor U3903 (N_3903,N_1156,N_877);
and U3904 (N_3904,N_678,N_2728);
nand U3905 (N_3905,N_101,N_398);
and U3906 (N_3906,N_359,N_2674);
nand U3907 (N_3907,N_1161,N_879);
nand U3908 (N_3908,N_1529,N_2411);
or U3909 (N_3909,N_2068,N_974);
nand U3910 (N_3910,N_135,N_222);
and U3911 (N_3911,N_2761,N_1283);
nor U3912 (N_3912,N_1571,N_2027);
and U3913 (N_3913,N_1845,N_1342);
or U3914 (N_3914,N_2276,N_2594);
nand U3915 (N_3915,N_1831,N_2795);
nand U3916 (N_3916,N_1969,N_2687);
or U3917 (N_3917,N_2159,N_1282);
nor U3918 (N_3918,N_842,N_2183);
nor U3919 (N_3919,N_713,N_157);
nor U3920 (N_3920,N_71,N_2546);
and U3921 (N_3921,N_2801,N_2466);
or U3922 (N_3922,N_1030,N_1640);
nor U3923 (N_3923,N_1033,N_1244);
or U3924 (N_3924,N_1935,N_1682);
nand U3925 (N_3925,N_1720,N_1045);
xnor U3926 (N_3926,N_1360,N_2443);
xnor U3927 (N_3927,N_316,N_816);
or U3928 (N_3928,N_655,N_69);
or U3929 (N_3929,N_482,N_1449);
nand U3930 (N_3930,N_2064,N_506);
nor U3931 (N_3931,N_218,N_2075);
and U3932 (N_3932,N_558,N_2065);
or U3933 (N_3933,N_2610,N_2063);
or U3934 (N_3934,N_2097,N_2062);
or U3935 (N_3935,N_995,N_312);
or U3936 (N_3936,N_671,N_2407);
and U3937 (N_3937,N_2057,N_186);
or U3938 (N_3938,N_0,N_2388);
or U3939 (N_3939,N_1287,N_1251);
and U3940 (N_3940,N_2843,N_1172);
nand U3941 (N_3941,N_2523,N_2611);
and U3942 (N_3942,N_2763,N_1415);
nor U3943 (N_3943,N_1505,N_108);
nand U3944 (N_3944,N_812,N_2686);
nor U3945 (N_3945,N_472,N_2106);
and U3946 (N_3946,N_1330,N_1394);
nand U3947 (N_3947,N_1880,N_2520);
nand U3948 (N_3948,N_1173,N_2797);
or U3949 (N_3949,N_1896,N_2483);
nand U3950 (N_3950,N_1907,N_1545);
nand U3951 (N_3951,N_284,N_2436);
or U3952 (N_3952,N_1677,N_155);
nor U3953 (N_3953,N_1971,N_1317);
nor U3954 (N_3954,N_836,N_2098);
or U3955 (N_3955,N_2786,N_440);
nor U3956 (N_3956,N_2654,N_2329);
or U3957 (N_3957,N_1742,N_1247);
and U3958 (N_3958,N_1290,N_1794);
or U3959 (N_3959,N_1195,N_1381);
nor U3960 (N_3960,N_1103,N_839);
nor U3961 (N_3961,N_1853,N_2040);
nor U3962 (N_3962,N_2490,N_1579);
nand U3963 (N_3963,N_137,N_1704);
xnor U3964 (N_3964,N_1090,N_2221);
or U3965 (N_3965,N_574,N_104);
and U3966 (N_3966,N_1812,N_820);
nand U3967 (N_3967,N_732,N_2033);
xor U3968 (N_3968,N_265,N_1757);
nor U3969 (N_3969,N_2132,N_2337);
and U3970 (N_3970,N_2376,N_2633);
or U3971 (N_3971,N_38,N_92);
nor U3972 (N_3972,N_2944,N_802);
nand U3973 (N_3973,N_1785,N_2387);
nand U3974 (N_3974,N_1101,N_2696);
nand U3975 (N_3975,N_1900,N_378);
xnor U3976 (N_3976,N_370,N_1067);
or U3977 (N_3977,N_1395,N_1448);
nand U3978 (N_3978,N_2838,N_47);
and U3979 (N_3979,N_503,N_1276);
nor U3980 (N_3980,N_1089,N_2282);
and U3981 (N_3981,N_2790,N_2267);
xnor U3982 (N_3982,N_2189,N_2774);
and U3983 (N_3983,N_2741,N_2235);
and U3984 (N_3984,N_1753,N_1167);
or U3985 (N_3985,N_2694,N_1566);
and U3986 (N_3986,N_123,N_381);
xor U3987 (N_3987,N_196,N_225);
nor U3988 (N_3988,N_464,N_1237);
and U3989 (N_3989,N_488,N_1587);
xor U3990 (N_3990,N_1653,N_1118);
or U3991 (N_3991,N_1211,N_2086);
nand U3992 (N_3992,N_1990,N_1274);
nor U3993 (N_3993,N_553,N_2503);
xor U3994 (N_3994,N_801,N_2143);
nor U3995 (N_3995,N_2322,N_1220);
nand U3996 (N_3996,N_2455,N_950);
nor U3997 (N_3997,N_2932,N_324);
or U3998 (N_3998,N_2649,N_708);
nand U3999 (N_3999,N_1303,N_2510);
and U4000 (N_4000,N_2961,N_668);
nand U4001 (N_4001,N_1081,N_1339);
or U4002 (N_4002,N_1453,N_74);
xnor U4003 (N_4003,N_2767,N_181);
nand U4004 (N_4004,N_572,N_335);
or U4005 (N_4005,N_2681,N_180);
nand U4006 (N_4006,N_2209,N_1295);
nand U4007 (N_4007,N_1500,N_1597);
nor U4008 (N_4008,N_1550,N_2518);
and U4009 (N_4009,N_1055,N_2982);
nor U4010 (N_4010,N_1956,N_268);
and U4011 (N_4011,N_2906,N_1694);
and U4012 (N_4012,N_2993,N_410);
nor U4013 (N_4013,N_559,N_2283);
nor U4014 (N_4014,N_423,N_1301);
and U4015 (N_4015,N_946,N_2859);
nand U4016 (N_4016,N_522,N_2441);
nand U4017 (N_4017,N_1507,N_2835);
xor U4018 (N_4018,N_616,N_2764);
and U4019 (N_4019,N_119,N_1135);
and U4020 (N_4020,N_2278,N_501);
and U4021 (N_4021,N_498,N_2477);
xnor U4022 (N_4022,N_573,N_810);
and U4023 (N_4023,N_1735,N_690);
nor U4024 (N_4024,N_2549,N_221);
or U4025 (N_4025,N_1367,N_2723);
nor U4026 (N_4026,N_2207,N_787);
or U4027 (N_4027,N_1779,N_1451);
nor U4028 (N_4028,N_1520,N_917);
nand U4029 (N_4029,N_523,N_1740);
or U4030 (N_4030,N_1960,N_2581);
or U4031 (N_4031,N_2628,N_1901);
nand U4032 (N_4032,N_1593,N_2281);
nand U4033 (N_4033,N_1060,N_2336);
or U4034 (N_4034,N_933,N_2333);
or U4035 (N_4035,N_748,N_2168);
xor U4036 (N_4036,N_2135,N_1953);
and U4037 (N_4037,N_2562,N_2688);
and U4038 (N_4038,N_1004,N_2423);
or U4039 (N_4039,N_1080,N_2692);
nor U4040 (N_4040,N_1177,N_281);
or U4041 (N_4041,N_2210,N_2531);
nand U4042 (N_4042,N_2799,N_310);
xnor U4043 (N_4043,N_1552,N_352);
and U4044 (N_4044,N_2417,N_1548);
nor U4045 (N_4045,N_1163,N_214);
nor U4046 (N_4046,N_2653,N_2757);
or U4047 (N_4047,N_1674,N_93);
nand U4048 (N_4048,N_1114,N_519);
nand U4049 (N_4049,N_2745,N_354);
or U4050 (N_4050,N_580,N_502);
and U4051 (N_4051,N_2985,N_1434);
nand U4052 (N_4052,N_156,N_441);
nand U4053 (N_4053,N_1153,N_1134);
or U4054 (N_4054,N_926,N_2725);
xor U4055 (N_4055,N_1058,N_2424);
and U4056 (N_4056,N_2645,N_639);
and U4057 (N_4057,N_1540,N_2370);
nand U4058 (N_4058,N_2085,N_1898);
and U4059 (N_4059,N_1234,N_1700);
or U4060 (N_4060,N_841,N_1633);
nor U4061 (N_4061,N_2701,N_2427);
nand U4062 (N_4062,N_1821,N_2729);
nor U4063 (N_4063,N_474,N_1886);
nor U4064 (N_4064,N_2800,N_1992);
xnor U4065 (N_4065,N_1185,N_1358);
nor U4066 (N_4066,N_1072,N_2663);
nand U4067 (N_4067,N_1736,N_2524);
or U4068 (N_4068,N_586,N_2839);
nand U4069 (N_4069,N_2921,N_2243);
and U4070 (N_4070,N_404,N_2111);
xnor U4071 (N_4071,N_1989,N_813);
or U4072 (N_4072,N_1474,N_854);
and U4073 (N_4073,N_524,N_110);
nand U4074 (N_4074,N_1414,N_821);
nand U4075 (N_4075,N_848,N_2716);
and U4076 (N_4076,N_2223,N_2141);
or U4077 (N_4077,N_1954,N_2133);
nand U4078 (N_4078,N_1122,N_1467);
or U4079 (N_4079,N_2325,N_442);
nor U4080 (N_4080,N_2926,N_1603);
nand U4081 (N_4081,N_2625,N_2829);
nand U4082 (N_4082,N_1048,N_353);
nor U4083 (N_4083,N_1692,N_2304);
and U4084 (N_4084,N_242,N_357);
nand U4085 (N_4085,N_2627,N_68);
nand U4086 (N_4086,N_259,N_1650);
nand U4087 (N_4087,N_1921,N_582);
and U4088 (N_4088,N_366,N_1607);
and U4089 (N_4089,N_833,N_2307);
or U4090 (N_4090,N_1426,N_739);
and U4091 (N_4091,N_1762,N_420);
nand U4092 (N_4092,N_2875,N_1142);
nand U4093 (N_4093,N_2112,N_2175);
and U4094 (N_4094,N_1800,N_1357);
or U4095 (N_4095,N_2272,N_294);
xor U4096 (N_4096,N_972,N_1388);
or U4097 (N_4097,N_2958,N_1834);
and U4098 (N_4098,N_886,N_1769);
and U4099 (N_4099,N_384,N_1933);
nand U4100 (N_4100,N_2452,N_2061);
or U4101 (N_4101,N_2451,N_931);
nand U4102 (N_4102,N_786,N_1648);
nand U4103 (N_4103,N_1582,N_2634);
or U4104 (N_4104,N_2306,N_1595);
xor U4105 (N_4105,N_1889,N_22);
nand U4106 (N_4106,N_2244,N_2515);
and U4107 (N_4107,N_2513,N_2756);
or U4108 (N_4108,N_1811,N_661);
nor U4109 (N_4109,N_1802,N_2025);
or U4110 (N_4110,N_1691,N_868);
and U4111 (N_4111,N_1804,N_796);
nand U4112 (N_4112,N_1331,N_1973);
nor U4113 (N_4113,N_2887,N_960);
and U4114 (N_4114,N_1017,N_2258);
and U4115 (N_4115,N_642,N_216);
nand U4116 (N_4116,N_1239,N_126);
and U4117 (N_4117,N_2009,N_2149);
nor U4118 (N_4118,N_1756,N_516);
nor U4119 (N_4119,N_855,N_1844);
nand U4120 (N_4120,N_1533,N_1689);
and U4121 (N_4121,N_2102,N_470);
and U4122 (N_4122,N_2691,N_1993);
and U4123 (N_4123,N_386,N_1567);
xnor U4124 (N_4124,N_947,N_1350);
nor U4125 (N_4125,N_418,N_779);
nor U4126 (N_4126,N_965,N_1318);
nor U4127 (N_4127,N_790,N_287);
and U4128 (N_4128,N_1726,N_443);
or U4129 (N_4129,N_719,N_2640);
or U4130 (N_4130,N_1348,N_258);
nand U4131 (N_4131,N_2629,N_245);
and U4132 (N_4132,N_2229,N_2005);
and U4133 (N_4133,N_2323,N_178);
or U4134 (N_4134,N_699,N_1730);
and U4135 (N_4135,N_754,N_1522);
xnor U4136 (N_4136,N_1722,N_860);
or U4137 (N_4137,N_185,N_959);
or U4138 (N_4138,N_858,N_240);
nor U4139 (N_4139,N_602,N_987);
or U4140 (N_4140,N_1363,N_2873);
nor U4141 (N_4141,N_308,N_696);
nor U4142 (N_4142,N_1663,N_1459);
or U4143 (N_4143,N_2208,N_112);
nor U4144 (N_4144,N_429,N_1098);
nor U4145 (N_4145,N_914,N_2036);
and U4146 (N_4146,N_529,N_1986);
nand U4147 (N_4147,N_2296,N_29);
nor U4148 (N_4148,N_2750,N_1611);
nand U4149 (N_4149,N_1670,N_938);
or U4150 (N_4150,N_2615,N_416);
and U4151 (N_4151,N_1493,N_1569);
nand U4152 (N_4152,N_1888,N_451);
nand U4153 (N_4153,N_1711,N_31);
and U4154 (N_4154,N_1176,N_814);
or U4155 (N_4155,N_2588,N_458);
and U4156 (N_4156,N_688,N_1997);
nand U4157 (N_4157,N_991,N_2607);
nand U4158 (N_4158,N_1732,N_2872);
and U4159 (N_4159,N_447,N_2724);
and U4160 (N_4160,N_279,N_1278);
nand U4161 (N_4161,N_2540,N_1936);
and U4162 (N_4162,N_2734,N_2832);
nand U4163 (N_4163,N_2496,N_1438);
nor U4164 (N_4164,N_2989,N_208);
nand U4165 (N_4165,N_811,N_2516);
or U4166 (N_4166,N_2319,N_266);
nand U4167 (N_4167,N_2831,N_446);
or U4168 (N_4168,N_2679,N_435);
or U4169 (N_4169,N_1021,N_1223);
or U4170 (N_4170,N_537,N_1599);
and U4171 (N_4171,N_1777,N_956);
nor U4172 (N_4172,N_1097,N_329);
or U4173 (N_4173,N_2213,N_2589);
nor U4174 (N_4174,N_2053,N_512);
xnor U4175 (N_4175,N_834,N_1123);
and U4176 (N_4176,N_2789,N_1046);
and U4177 (N_4177,N_338,N_190);
nor U4178 (N_4178,N_1105,N_1445);
nand U4179 (N_4179,N_986,N_1686);
nor U4180 (N_4180,N_2664,N_1183);
nor U4181 (N_4181,N_1849,N_1531);
nor U4182 (N_4182,N_2301,N_637);
or U4183 (N_4183,N_1349,N_2459);
and U4184 (N_4184,N_1561,N_2071);
xor U4185 (N_4185,N_1645,N_379);
nor U4186 (N_4186,N_870,N_2667);
or U4187 (N_4187,N_1840,N_1808);
nand U4188 (N_4188,N_2334,N_2402);
nand U4189 (N_4189,N_1656,N_142);
nor U4190 (N_4190,N_365,N_254);
xor U4191 (N_4191,N_1180,N_1703);
nand U4192 (N_4192,N_849,N_873);
nor U4193 (N_4193,N_318,N_2437);
or U4194 (N_4194,N_2342,N_578);
and U4195 (N_4195,N_1420,N_2099);
nor U4196 (N_4196,N_1672,N_2172);
or U4197 (N_4197,N_2487,N_122);
nand U4198 (N_4198,N_309,N_1431);
or U4199 (N_4199,N_403,N_1744);
nor U4200 (N_4200,N_2115,N_659);
xnor U4201 (N_4201,N_962,N_1216);
or U4202 (N_4202,N_2842,N_1082);
nor U4203 (N_4203,N_930,N_2769);
nand U4204 (N_4204,N_2430,N_1539);
and U4205 (N_4205,N_546,N_461);
nor U4206 (N_4206,N_2824,N_2401);
or U4207 (N_4207,N_2836,N_1942);
nand U4208 (N_4208,N_2216,N_228);
and U4209 (N_4209,N_2266,N_1589);
or U4210 (N_4210,N_782,N_219);
or U4211 (N_4211,N_246,N_1930);
and U4212 (N_4212,N_2446,N_1147);
nor U4213 (N_4213,N_712,N_1343);
and U4214 (N_4214,N_1417,N_19);
nand U4215 (N_4215,N_2428,N_2551);
nand U4216 (N_4216,N_2855,N_2044);
xor U4217 (N_4217,N_943,N_1631);
nor U4218 (N_4218,N_1155,N_2249);
nor U4219 (N_4219,N_351,N_288);
nor U4220 (N_4220,N_1409,N_2532);
or U4221 (N_4221,N_2935,N_1439);
nand U4222 (N_4222,N_1499,N_1393);
nand U4223 (N_4223,N_587,N_682);
or U4224 (N_4224,N_450,N_2709);
nand U4225 (N_4225,N_2250,N_66);
nand U4226 (N_4226,N_2200,N_2182);
and U4227 (N_4227,N_1215,N_293);
and U4228 (N_4228,N_2773,N_2822);
and U4229 (N_4229,N_1321,N_2575);
nor U4230 (N_4230,N_121,N_291);
nor U4231 (N_4231,N_1212,N_223);
or U4232 (N_4232,N_2666,N_2785);
nand U4233 (N_4233,N_1623,N_532);
nand U4234 (N_4234,N_539,N_1099);
or U4235 (N_4235,N_2134,N_1675);
or U4236 (N_4236,N_248,N_1897);
or U4237 (N_4237,N_1851,N_1473);
xnor U4238 (N_4238,N_2505,N_874);
nor U4239 (N_4239,N_2205,N_1946);
or U4240 (N_4240,N_2595,N_496);
and U4241 (N_4241,N_2497,N_1245);
nand U4242 (N_4242,N_2214,N_1057);
nand U4243 (N_4243,N_2242,N_2568);
nor U4244 (N_4244,N_681,N_64);
and U4245 (N_4245,N_2814,N_2868);
nor U4246 (N_4246,N_462,N_2104);
nand U4247 (N_4247,N_2147,N_2468);
nor U4248 (N_4248,N_1680,N_1627);
and U4249 (N_4249,N_1850,N_707);
nor U4250 (N_4250,N_2328,N_992);
and U4251 (N_4251,N_2735,N_689);
nand U4252 (N_4252,N_793,N_1373);
or U4253 (N_4253,N_1074,N_1110);
nor U4254 (N_4254,N_1541,N_971);
nor U4255 (N_4255,N_2087,N_595);
nor U4256 (N_4256,N_1327,N_1559);
and U4257 (N_4257,N_1014,N_2671);
and U4258 (N_4258,N_1052,N_892);
xor U4259 (N_4259,N_395,N_1042);
nor U4260 (N_4260,N_2997,N_2414);
or U4261 (N_4261,N_1136,N_1174);
or U4262 (N_4262,N_1232,N_758);
nand U4263 (N_4263,N_1764,N_1797);
nor U4264 (N_4264,N_2386,N_2024);
xnor U4265 (N_4265,N_1119,N_2541);
nor U4266 (N_4266,N_805,N_2160);
xor U4267 (N_4267,N_2570,N_1578);
nor U4268 (N_4268,N_2793,N_861);
and U4269 (N_4269,N_300,N_864);
nand U4270 (N_4270,N_2331,N_1799);
or U4271 (N_4271,N_2454,N_838);
nor U4272 (N_4272,N_1822,N_1192);
nand U4273 (N_4273,N_160,N_653);
and U4274 (N_4274,N_1641,N_39);
nor U4275 (N_4275,N_565,N_1100);
nand U4276 (N_4276,N_1959,N_2939);
and U4277 (N_4277,N_362,N_2130);
nand U4278 (N_4278,N_1944,N_1264);
or U4279 (N_4279,N_924,N_889);
nor U4280 (N_4280,N_2326,N_161);
and U4281 (N_4281,N_2721,N_1536);
nor U4282 (N_4282,N_772,N_212);
and U4283 (N_4283,N_2,N_1027);
nor U4284 (N_4284,N_86,N_344);
nand U4285 (N_4285,N_1564,N_557);
nor U4286 (N_4286,N_620,N_727);
xnor U4287 (N_4287,N_1855,N_2950);
and U4288 (N_4288,N_597,N_2772);
or U4289 (N_4289,N_1838,N_2318);
and U4290 (N_4290,N_106,N_2782);
xnor U4291 (N_4291,N_2426,N_264);
and U4292 (N_4292,N_1580,N_2954);
nand U4293 (N_4293,N_2375,N_127);
or U4294 (N_4294,N_2327,N_670);
nand U4295 (N_4295,N_1023,N_1585);
or U4296 (N_4296,N_1509,N_2389);
nand U4297 (N_4297,N_1681,N_195);
or U4298 (N_4298,N_2224,N_2045);
xnor U4299 (N_4299,N_2804,N_306);
xor U4300 (N_4300,N_2472,N_1219);
and U4301 (N_4301,N_2093,N_1202);
or U4302 (N_4302,N_1970,N_2237);
or U4303 (N_4303,N_2907,N_298);
nand U4304 (N_4304,N_457,N_147);
nor U4305 (N_4305,N_145,N_285);
or U4306 (N_4306,N_901,N_1132);
or U4307 (N_4307,N_2990,N_1608);
or U4308 (N_4308,N_1158,N_1698);
nor U4309 (N_4309,N_1179,N_2623);
nand U4310 (N_4310,N_581,N_1421);
xor U4311 (N_4311,N_2536,N_1049);
nand U4312 (N_4312,N_675,N_2861);
xnor U4313 (N_4313,N_1878,N_2876);
and U4314 (N_4314,N_828,N_406);
nor U4315 (N_4315,N_2354,N_1739);
xor U4316 (N_4316,N_730,N_1044);
nor U4317 (N_4317,N_993,N_1452);
or U4318 (N_4318,N_1356,N_1224);
and U4319 (N_4319,N_2367,N_2293);
nand U4320 (N_4320,N_2752,N_2991);
and U4321 (N_4321,N_1874,N_694);
nor U4322 (N_4322,N_605,N_1940);
nand U4323 (N_4323,N_887,N_1458);
nand U4324 (N_4324,N_923,N_2744);
nand U4325 (N_4325,N_2963,N_1801);
nor U4326 (N_4326,N_2456,N_2299);
or U4327 (N_4327,N_1865,N_1);
nand U4328 (N_4328,N_400,N_2262);
nor U4329 (N_4329,N_819,N_1306);
and U4330 (N_4330,N_1187,N_2173);
or U4331 (N_4331,N_2893,N_530);
nor U4332 (N_4332,N_2265,N_2833);
and U4333 (N_4333,N_2740,N_1619);
or U4334 (N_4334,N_1390,N_2830);
nand U4335 (N_4335,N_448,N_2034);
and U4336 (N_4336,N_1115,N_1630);
or U4337 (N_4337,N_1141,N_374);
nor U4338 (N_4338,N_1521,N_428);
or U4339 (N_4339,N_2702,N_542);
nor U4340 (N_4340,N_1364,N_16);
nor U4341 (N_4341,N_432,N_2489);
nor U4342 (N_4342,N_1284,N_2251);
and U4343 (N_4343,N_2931,N_633);
nand U4344 (N_4344,N_1406,N_1718);
nand U4345 (N_4345,N_176,N_866);
nand U4346 (N_4346,N_2864,N_1523);
nand U4347 (N_4347,N_204,N_2689);
or U4348 (N_4348,N_2051,N_2006);
nand U4349 (N_4349,N_371,N_2028);
and U4350 (N_4350,N_2783,N_1456);
nand U4351 (N_4351,N_1885,N_1554);
and U4352 (N_4352,N_607,N_90);
or U4353 (N_4353,N_1376,N_1781);
or U4354 (N_4354,N_2881,N_1977);
nand U4355 (N_4355,N_2476,N_2665);
or U4356 (N_4356,N_915,N_91);
nor U4357 (N_4357,N_431,N_2460);
or U4358 (N_4358,N_2560,N_276);
nor U4359 (N_4359,N_1484,N_2410);
nor U4360 (N_4360,N_337,N_2501);
nand U4361 (N_4361,N_1870,N_2137);
nor U4362 (N_4362,N_1277,N_953);
nand U4363 (N_4363,N_847,N_1159);
xnor U4364 (N_4364,N_723,N_49);
and U4365 (N_4365,N_2245,N_206);
or U4366 (N_4366,N_1337,N_2169);
xor U4367 (N_4367,N_2269,N_2444);
nand U4368 (N_4368,N_1667,N_311);
or U4369 (N_4369,N_169,N_515);
or U4370 (N_4370,N_2310,N_2359);
nand U4371 (N_4371,N_896,N_766);
or U4372 (N_4372,N_1784,N_957);
and U4373 (N_4373,N_1126,N_996);
nor U4374 (N_4374,N_2270,N_880);
nand U4375 (N_4375,N_2491,N_277);
nor U4376 (N_4376,N_1385,N_2008);
or U4377 (N_4377,N_702,N_2395);
nand U4378 (N_4378,N_1503,N_700);
and U4379 (N_4379,N_2959,N_33);
xnor U4380 (N_4380,N_1932,N_1455);
xnor U4381 (N_4381,N_307,N_1059);
nor U4382 (N_4382,N_1904,N_1966);
nor U4383 (N_4383,N_846,N_1262);
xnor U4384 (N_4384,N_299,N_1137);
nand U4385 (N_4385,N_267,N_884);
nand U4386 (N_4386,N_491,N_2379);
and U4387 (N_4387,N_1884,N_292);
or U4388 (N_4388,N_1558,N_1094);
nand U4389 (N_4389,N_2383,N_290);
nand U4390 (N_4390,N_35,N_456);
nor U4391 (N_4391,N_2758,N_1032);
nor U4392 (N_4392,N_270,N_1950);
nand U4393 (N_4393,N_1872,N_1062);
nand U4394 (N_4394,N_325,N_2916);
xor U4395 (N_4395,N_909,N_1170);
and U4396 (N_4396,N_2092,N_54);
or U4397 (N_4397,N_692,N_1408);
and U4398 (N_4398,N_2988,N_489);
nor U4399 (N_4399,N_1514,N_704);
and U4400 (N_4400,N_2077,N_1988);
nand U4401 (N_4401,N_852,N_1065);
and U4402 (N_4402,N_2222,N_1876);
nor U4403 (N_4403,N_1370,N_10);
and U4404 (N_4404,N_1832,N_509);
xor U4405 (N_4405,N_1240,N_2066);
xor U4406 (N_4406,N_1945,N_1465);
xnor U4407 (N_4407,N_2947,N_1551);
nand U4408 (N_4408,N_2641,N_2022);
nand U4409 (N_4409,N_109,N_3);
nor U4410 (N_4410,N_1345,N_1404);
xor U4411 (N_4411,N_1107,N_1208);
nand U4412 (N_4412,N_2046,N_1272);
and U4413 (N_4413,N_2335,N_1600);
xnor U4414 (N_4414,N_1476,N_320);
and U4415 (N_4415,N_2125,N_1311);
or U4416 (N_4416,N_560,N_1543);
nor U4417 (N_4417,N_1848,N_1164);
or U4418 (N_4418,N_1478,N_2003);
or U4419 (N_4419,N_427,N_908);
and U4420 (N_4420,N_2016,N_657);
nor U4421 (N_4421,N_2605,N_302);
nand U4422 (N_4422,N_794,N_1734);
or U4423 (N_4423,N_1780,N_2644);
and U4424 (N_4424,N_1116,N_1011);
or U4425 (N_4425,N_1188,N_2852);
nor U4426 (N_4426,N_695,N_1823);
and U4427 (N_4427,N_911,N_533);
nor U4428 (N_4428,N_541,N_994);
nor U4429 (N_4429,N_893,N_1975);
or U4430 (N_4430,N_851,N_2727);
nand U4431 (N_4431,N_2621,N_2517);
nand U4432 (N_4432,N_2332,N_2413);
and U4433 (N_4433,N_663,N_444);
or U4434 (N_4434,N_781,N_1334);
xor U4435 (N_4435,N_2592,N_2714);
nand U4436 (N_4436,N_43,N_2215);
or U4437 (N_4437,N_72,N_1594);
or U4438 (N_4438,N_149,N_1131);
nor U4439 (N_4439,N_891,N_2217);
nand U4440 (N_4440,N_1085,N_2826);
and U4441 (N_4441,N_2919,N_1148);
nor U4442 (N_4442,N_1151,N_158);
or U4443 (N_4443,N_1515,N_177);
or U4444 (N_4444,N_263,N_1053);
and U4445 (N_4445,N_2156,N_46);
and U4446 (N_4446,N_2847,N_984);
nand U4447 (N_4447,N_1346,N_152);
or U4448 (N_4448,N_2364,N_2925);
or U4449 (N_4449,N_2747,N_2498);
xnor U4450 (N_4450,N_1242,N_569);
nor U4451 (N_4451,N_215,N_1093);
and U4452 (N_4452,N_592,N_750);
or U4453 (N_4453,N_1351,N_389);
nor U4454 (N_4454,N_170,N_2846);
or U4455 (N_4455,N_1565,N_399);
nand U4456 (N_4456,N_2966,N_2883);
or U4457 (N_4457,N_2828,N_2348);
nand U4458 (N_4458,N_762,N_2538);
or U4459 (N_4459,N_2550,N_1612);
and U4460 (N_4460,N_624,N_825);
and U4461 (N_4461,N_544,N_2899);
nor U4462 (N_4462,N_513,N_2122);
nor U4463 (N_4463,N_2397,N_2508);
and U4464 (N_4464,N_1894,N_1341);
and U4465 (N_4465,N_1961,N_632);
nor U4466 (N_4466,N_2849,N_1895);
nor U4467 (N_4467,N_2992,N_390);
or U4468 (N_4468,N_1104,N_1203);
nor U4469 (N_4469,N_2360,N_1479);
or U4470 (N_4470,N_2630,N_2218);
and U4471 (N_4471,N_1791,N_2356);
xor U4472 (N_4472,N_1664,N_815);
nand U4473 (N_4473,N_2616,N_296);
or U4474 (N_4474,N_1236,N_89);
and U4475 (N_4475,N_1951,N_1194);
xnor U4476 (N_4476,N_1759,N_662);
xnor U4477 (N_4477,N_2453,N_660);
and U4478 (N_4478,N_2385,N_853);
nand U4479 (N_4479,N_2526,N_910);
nand U4480 (N_4480,N_2176,N_2973);
nor U4481 (N_4481,N_1679,N_396);
nand U4482 (N_4482,N_1857,N_471);
and U4483 (N_4483,N_2113,N_1353);
nor U4484 (N_4484,N_1980,N_2261);
nor U4485 (N_4485,N_12,N_1166);
nor U4486 (N_4486,N_776,N_2236);
and U4487 (N_4487,N_2330,N_2994);
and U4488 (N_4488,N_2571,N_1806);
or U4489 (N_4489,N_1755,N_2816);
and U4490 (N_4490,N_2448,N_562);
nor U4491 (N_4491,N_1444,N_133);
xor U4492 (N_4492,N_1591,N_2943);
nor U4493 (N_4493,N_1320,N_1392);
nor U4494 (N_4494,N_1425,N_2035);
nor U4495 (N_4495,N_1086,N_2922);
or U4496 (N_4496,N_2029,N_2366);
or U4497 (N_4497,N_2810,N_1079);
nor U4498 (N_4498,N_4,N_919);
and U4499 (N_4499,N_2039,N_2597);
or U4500 (N_4500,N_2973,N_954);
or U4501 (N_4501,N_2337,N_2143);
nand U4502 (N_4502,N_409,N_119);
nor U4503 (N_4503,N_2429,N_2334);
and U4504 (N_4504,N_478,N_2628);
nand U4505 (N_4505,N_833,N_189);
or U4506 (N_4506,N_1366,N_2774);
nor U4507 (N_4507,N_1319,N_6);
nor U4508 (N_4508,N_1706,N_2012);
nand U4509 (N_4509,N_1527,N_234);
xor U4510 (N_4510,N_2329,N_692);
nand U4511 (N_4511,N_2878,N_1399);
nor U4512 (N_4512,N_2232,N_2913);
and U4513 (N_4513,N_1843,N_1622);
nand U4514 (N_4514,N_377,N_292);
xnor U4515 (N_4515,N_1807,N_1136);
or U4516 (N_4516,N_1455,N_440);
xor U4517 (N_4517,N_1520,N_1951);
nor U4518 (N_4518,N_1426,N_2624);
nand U4519 (N_4519,N_752,N_842);
or U4520 (N_4520,N_99,N_626);
nand U4521 (N_4521,N_1823,N_1316);
and U4522 (N_4522,N_174,N_445);
or U4523 (N_4523,N_2786,N_2686);
nand U4524 (N_4524,N_2817,N_2144);
or U4525 (N_4525,N_2959,N_304);
and U4526 (N_4526,N_765,N_1729);
nand U4527 (N_4527,N_2206,N_1040);
nor U4528 (N_4528,N_2777,N_2094);
nor U4529 (N_4529,N_838,N_672);
nor U4530 (N_4530,N_2849,N_157);
nor U4531 (N_4531,N_596,N_2600);
nand U4532 (N_4532,N_259,N_886);
or U4533 (N_4533,N_2776,N_2426);
and U4534 (N_4534,N_2623,N_220);
or U4535 (N_4535,N_82,N_2164);
nand U4536 (N_4536,N_2266,N_1755);
and U4537 (N_4537,N_2673,N_2557);
and U4538 (N_4538,N_1132,N_699);
or U4539 (N_4539,N_2093,N_2477);
and U4540 (N_4540,N_2534,N_430);
and U4541 (N_4541,N_2063,N_1489);
nor U4542 (N_4542,N_101,N_2241);
nand U4543 (N_4543,N_2258,N_2391);
nor U4544 (N_4544,N_1111,N_320);
or U4545 (N_4545,N_1088,N_2223);
and U4546 (N_4546,N_532,N_2238);
or U4547 (N_4547,N_598,N_2797);
nand U4548 (N_4548,N_2756,N_1055);
nor U4549 (N_4549,N_1222,N_2419);
or U4550 (N_4550,N_250,N_283);
nor U4551 (N_4551,N_1986,N_2952);
nor U4552 (N_4552,N_1577,N_117);
nor U4553 (N_4553,N_420,N_2266);
and U4554 (N_4554,N_74,N_1552);
or U4555 (N_4555,N_663,N_37);
or U4556 (N_4556,N_2846,N_2315);
or U4557 (N_4557,N_1672,N_1859);
and U4558 (N_4558,N_2710,N_552);
xnor U4559 (N_4559,N_1032,N_2901);
and U4560 (N_4560,N_2866,N_1282);
nand U4561 (N_4561,N_5,N_2435);
nor U4562 (N_4562,N_2736,N_848);
or U4563 (N_4563,N_197,N_550);
nor U4564 (N_4564,N_2425,N_1886);
and U4565 (N_4565,N_170,N_2176);
and U4566 (N_4566,N_2962,N_2716);
nor U4567 (N_4567,N_2728,N_89);
and U4568 (N_4568,N_982,N_2410);
and U4569 (N_4569,N_1921,N_2041);
or U4570 (N_4570,N_432,N_361);
nor U4571 (N_4571,N_417,N_2116);
nor U4572 (N_4572,N_1050,N_1461);
or U4573 (N_4573,N_782,N_1932);
nor U4574 (N_4574,N_65,N_1717);
nor U4575 (N_4575,N_56,N_1106);
and U4576 (N_4576,N_368,N_285);
or U4577 (N_4577,N_2075,N_950);
or U4578 (N_4578,N_2785,N_1190);
nor U4579 (N_4579,N_183,N_2179);
nor U4580 (N_4580,N_2304,N_1432);
nor U4581 (N_4581,N_1140,N_2125);
nand U4582 (N_4582,N_2137,N_247);
and U4583 (N_4583,N_1290,N_1723);
nor U4584 (N_4584,N_2454,N_481);
nand U4585 (N_4585,N_1570,N_774);
nand U4586 (N_4586,N_1840,N_736);
or U4587 (N_4587,N_711,N_1693);
or U4588 (N_4588,N_524,N_394);
nor U4589 (N_4589,N_765,N_1327);
or U4590 (N_4590,N_1332,N_1508);
and U4591 (N_4591,N_393,N_1656);
nor U4592 (N_4592,N_916,N_2918);
and U4593 (N_4593,N_1735,N_123);
or U4594 (N_4594,N_600,N_1883);
and U4595 (N_4595,N_2568,N_964);
nand U4596 (N_4596,N_1760,N_1327);
xor U4597 (N_4597,N_61,N_945);
xnor U4598 (N_4598,N_1479,N_2661);
xor U4599 (N_4599,N_2943,N_1145);
nor U4600 (N_4600,N_2728,N_2048);
or U4601 (N_4601,N_1103,N_34);
xnor U4602 (N_4602,N_1825,N_1580);
and U4603 (N_4603,N_857,N_149);
nand U4604 (N_4604,N_2438,N_984);
and U4605 (N_4605,N_170,N_271);
nor U4606 (N_4606,N_1785,N_467);
and U4607 (N_4607,N_158,N_2162);
nand U4608 (N_4608,N_1032,N_1459);
and U4609 (N_4609,N_1372,N_471);
and U4610 (N_4610,N_2819,N_852);
or U4611 (N_4611,N_1310,N_438);
nor U4612 (N_4612,N_669,N_745);
and U4613 (N_4613,N_1326,N_563);
nand U4614 (N_4614,N_1603,N_2944);
and U4615 (N_4615,N_690,N_2394);
xnor U4616 (N_4616,N_923,N_1418);
or U4617 (N_4617,N_2222,N_1095);
and U4618 (N_4618,N_2744,N_2240);
nand U4619 (N_4619,N_2544,N_197);
nand U4620 (N_4620,N_64,N_2245);
xnor U4621 (N_4621,N_1698,N_2333);
xor U4622 (N_4622,N_576,N_2432);
nor U4623 (N_4623,N_1692,N_1926);
xnor U4624 (N_4624,N_2355,N_1135);
and U4625 (N_4625,N_1687,N_1894);
or U4626 (N_4626,N_1292,N_2624);
nand U4627 (N_4627,N_2127,N_627);
nor U4628 (N_4628,N_406,N_2491);
nor U4629 (N_4629,N_742,N_2431);
or U4630 (N_4630,N_2326,N_2156);
and U4631 (N_4631,N_343,N_474);
or U4632 (N_4632,N_1066,N_2804);
or U4633 (N_4633,N_439,N_785);
nor U4634 (N_4634,N_2965,N_928);
and U4635 (N_4635,N_1334,N_1307);
or U4636 (N_4636,N_1013,N_2885);
nor U4637 (N_4637,N_1000,N_469);
nand U4638 (N_4638,N_2877,N_1943);
or U4639 (N_4639,N_487,N_472);
and U4640 (N_4640,N_179,N_2580);
nor U4641 (N_4641,N_2859,N_1611);
and U4642 (N_4642,N_2066,N_1042);
and U4643 (N_4643,N_528,N_2458);
nor U4644 (N_4644,N_2928,N_107);
nor U4645 (N_4645,N_744,N_562);
and U4646 (N_4646,N_1477,N_1670);
nor U4647 (N_4647,N_1476,N_2136);
nand U4648 (N_4648,N_1532,N_2525);
and U4649 (N_4649,N_1063,N_682);
nor U4650 (N_4650,N_1624,N_810);
or U4651 (N_4651,N_382,N_588);
nor U4652 (N_4652,N_1233,N_2928);
and U4653 (N_4653,N_493,N_2803);
xnor U4654 (N_4654,N_1678,N_1912);
or U4655 (N_4655,N_385,N_1517);
or U4656 (N_4656,N_1418,N_428);
or U4657 (N_4657,N_1632,N_459);
nand U4658 (N_4658,N_1071,N_968);
nand U4659 (N_4659,N_690,N_1270);
or U4660 (N_4660,N_2125,N_1694);
and U4661 (N_4661,N_2915,N_1684);
and U4662 (N_4662,N_1872,N_2657);
or U4663 (N_4663,N_1128,N_1762);
xnor U4664 (N_4664,N_274,N_2139);
nand U4665 (N_4665,N_1820,N_514);
nand U4666 (N_4666,N_407,N_1398);
nand U4667 (N_4667,N_836,N_896);
nand U4668 (N_4668,N_638,N_21);
nor U4669 (N_4669,N_851,N_903);
and U4670 (N_4670,N_847,N_516);
or U4671 (N_4671,N_327,N_451);
and U4672 (N_4672,N_1880,N_1811);
and U4673 (N_4673,N_420,N_2487);
and U4674 (N_4674,N_469,N_2655);
nand U4675 (N_4675,N_1363,N_2266);
and U4676 (N_4676,N_944,N_1031);
nor U4677 (N_4677,N_2782,N_2380);
nand U4678 (N_4678,N_222,N_505);
nor U4679 (N_4679,N_186,N_2587);
and U4680 (N_4680,N_2248,N_429);
nor U4681 (N_4681,N_2787,N_774);
or U4682 (N_4682,N_608,N_428);
and U4683 (N_4683,N_74,N_1275);
nor U4684 (N_4684,N_138,N_403);
and U4685 (N_4685,N_1798,N_1563);
nor U4686 (N_4686,N_2469,N_1730);
or U4687 (N_4687,N_213,N_672);
nor U4688 (N_4688,N_2744,N_1444);
and U4689 (N_4689,N_2068,N_1451);
xnor U4690 (N_4690,N_1583,N_750);
and U4691 (N_4691,N_2692,N_2872);
or U4692 (N_4692,N_2125,N_2085);
nor U4693 (N_4693,N_1968,N_1379);
or U4694 (N_4694,N_1166,N_1387);
or U4695 (N_4695,N_2297,N_2179);
or U4696 (N_4696,N_2521,N_1525);
nor U4697 (N_4697,N_2596,N_425);
and U4698 (N_4698,N_1808,N_2214);
nor U4699 (N_4699,N_104,N_1714);
nor U4700 (N_4700,N_694,N_194);
nand U4701 (N_4701,N_728,N_2121);
nor U4702 (N_4702,N_1273,N_221);
nor U4703 (N_4703,N_293,N_1756);
nor U4704 (N_4704,N_412,N_566);
and U4705 (N_4705,N_2187,N_2151);
nand U4706 (N_4706,N_2941,N_545);
nand U4707 (N_4707,N_1788,N_1969);
and U4708 (N_4708,N_1929,N_2486);
nor U4709 (N_4709,N_1734,N_2657);
and U4710 (N_4710,N_2525,N_1837);
nor U4711 (N_4711,N_2390,N_1889);
or U4712 (N_4712,N_1595,N_1448);
or U4713 (N_4713,N_2830,N_979);
nand U4714 (N_4714,N_2371,N_1218);
nand U4715 (N_4715,N_830,N_664);
nor U4716 (N_4716,N_1878,N_1333);
nor U4717 (N_4717,N_2321,N_2930);
nand U4718 (N_4718,N_2724,N_1544);
or U4719 (N_4719,N_1668,N_1324);
nor U4720 (N_4720,N_1643,N_2924);
and U4721 (N_4721,N_505,N_1082);
nand U4722 (N_4722,N_594,N_599);
xor U4723 (N_4723,N_817,N_2500);
or U4724 (N_4724,N_1679,N_1977);
nand U4725 (N_4725,N_1659,N_1355);
or U4726 (N_4726,N_442,N_517);
nand U4727 (N_4727,N_1998,N_791);
nand U4728 (N_4728,N_2211,N_1619);
xor U4729 (N_4729,N_624,N_764);
nand U4730 (N_4730,N_1556,N_842);
xnor U4731 (N_4731,N_2172,N_447);
nor U4732 (N_4732,N_793,N_2458);
or U4733 (N_4733,N_727,N_1846);
nand U4734 (N_4734,N_2863,N_2697);
and U4735 (N_4735,N_2377,N_1417);
and U4736 (N_4736,N_375,N_1969);
or U4737 (N_4737,N_418,N_992);
xnor U4738 (N_4738,N_788,N_1691);
nor U4739 (N_4739,N_2021,N_808);
nor U4740 (N_4740,N_2579,N_478);
and U4741 (N_4741,N_1382,N_494);
or U4742 (N_4742,N_2994,N_1945);
nand U4743 (N_4743,N_2258,N_323);
or U4744 (N_4744,N_167,N_1612);
or U4745 (N_4745,N_264,N_2629);
or U4746 (N_4746,N_198,N_2848);
or U4747 (N_4747,N_1501,N_2603);
nand U4748 (N_4748,N_2284,N_1876);
or U4749 (N_4749,N_1911,N_1884);
nor U4750 (N_4750,N_1583,N_375);
and U4751 (N_4751,N_1785,N_2707);
or U4752 (N_4752,N_1011,N_2191);
nand U4753 (N_4753,N_2597,N_1282);
nor U4754 (N_4754,N_2560,N_100);
nand U4755 (N_4755,N_1136,N_2962);
nor U4756 (N_4756,N_1212,N_1578);
or U4757 (N_4757,N_2172,N_342);
and U4758 (N_4758,N_1715,N_2562);
xor U4759 (N_4759,N_687,N_310);
or U4760 (N_4760,N_2815,N_1847);
nor U4761 (N_4761,N_2534,N_606);
nand U4762 (N_4762,N_800,N_115);
and U4763 (N_4763,N_303,N_1342);
nand U4764 (N_4764,N_2050,N_1536);
xnor U4765 (N_4765,N_2699,N_1255);
xnor U4766 (N_4766,N_198,N_1384);
or U4767 (N_4767,N_1458,N_2647);
xnor U4768 (N_4768,N_1474,N_1964);
and U4769 (N_4769,N_2074,N_171);
or U4770 (N_4770,N_803,N_505);
nor U4771 (N_4771,N_1856,N_1610);
and U4772 (N_4772,N_728,N_407);
and U4773 (N_4773,N_972,N_2632);
and U4774 (N_4774,N_2615,N_1010);
nor U4775 (N_4775,N_399,N_2961);
xor U4776 (N_4776,N_2351,N_154);
nand U4777 (N_4777,N_673,N_2521);
nor U4778 (N_4778,N_2061,N_2391);
nor U4779 (N_4779,N_2353,N_2526);
nor U4780 (N_4780,N_1100,N_1009);
nor U4781 (N_4781,N_1173,N_1973);
nand U4782 (N_4782,N_1902,N_544);
and U4783 (N_4783,N_780,N_2291);
nand U4784 (N_4784,N_2647,N_1028);
nand U4785 (N_4785,N_328,N_1171);
and U4786 (N_4786,N_1070,N_1229);
nor U4787 (N_4787,N_1669,N_1739);
nor U4788 (N_4788,N_1127,N_1564);
nand U4789 (N_4789,N_2707,N_1044);
and U4790 (N_4790,N_819,N_101);
nand U4791 (N_4791,N_460,N_1806);
or U4792 (N_4792,N_2224,N_636);
nor U4793 (N_4793,N_1751,N_1456);
nor U4794 (N_4794,N_597,N_1411);
and U4795 (N_4795,N_1626,N_2048);
nand U4796 (N_4796,N_2557,N_24);
nand U4797 (N_4797,N_2008,N_2898);
and U4798 (N_4798,N_2230,N_2614);
xnor U4799 (N_4799,N_2891,N_1225);
and U4800 (N_4800,N_781,N_1165);
nand U4801 (N_4801,N_1604,N_957);
and U4802 (N_4802,N_1252,N_2128);
nand U4803 (N_4803,N_896,N_2355);
and U4804 (N_4804,N_1237,N_2747);
nor U4805 (N_4805,N_636,N_2931);
xnor U4806 (N_4806,N_1761,N_2806);
and U4807 (N_4807,N_302,N_225);
nand U4808 (N_4808,N_628,N_233);
and U4809 (N_4809,N_1981,N_1439);
or U4810 (N_4810,N_2062,N_1544);
nand U4811 (N_4811,N_2318,N_1721);
nand U4812 (N_4812,N_54,N_624);
nor U4813 (N_4813,N_1136,N_2939);
or U4814 (N_4814,N_634,N_896);
nand U4815 (N_4815,N_2305,N_1510);
or U4816 (N_4816,N_1504,N_244);
nand U4817 (N_4817,N_460,N_1570);
nor U4818 (N_4818,N_1641,N_2088);
or U4819 (N_4819,N_2773,N_56);
xor U4820 (N_4820,N_855,N_750);
and U4821 (N_4821,N_1665,N_2377);
nand U4822 (N_4822,N_94,N_843);
nor U4823 (N_4823,N_2184,N_2479);
nand U4824 (N_4824,N_2530,N_1121);
and U4825 (N_4825,N_2456,N_747);
and U4826 (N_4826,N_22,N_2362);
nor U4827 (N_4827,N_2788,N_1072);
or U4828 (N_4828,N_2502,N_1975);
and U4829 (N_4829,N_2698,N_1014);
nand U4830 (N_4830,N_2543,N_1698);
xor U4831 (N_4831,N_2194,N_1257);
nand U4832 (N_4832,N_2950,N_2552);
nand U4833 (N_4833,N_672,N_2076);
nand U4834 (N_4834,N_2913,N_499);
and U4835 (N_4835,N_2338,N_1082);
nor U4836 (N_4836,N_365,N_258);
nor U4837 (N_4837,N_379,N_422);
nand U4838 (N_4838,N_925,N_569);
nand U4839 (N_4839,N_2462,N_1433);
or U4840 (N_4840,N_2171,N_1829);
nand U4841 (N_4841,N_1425,N_23);
nand U4842 (N_4842,N_2394,N_1023);
nand U4843 (N_4843,N_1432,N_1228);
nor U4844 (N_4844,N_540,N_1428);
nand U4845 (N_4845,N_1170,N_2854);
and U4846 (N_4846,N_2961,N_1753);
xnor U4847 (N_4847,N_1599,N_1723);
nand U4848 (N_4848,N_1240,N_223);
nand U4849 (N_4849,N_699,N_2519);
and U4850 (N_4850,N_1397,N_962);
nor U4851 (N_4851,N_795,N_527);
nor U4852 (N_4852,N_844,N_731);
nor U4853 (N_4853,N_2529,N_2652);
and U4854 (N_4854,N_2157,N_1295);
nand U4855 (N_4855,N_986,N_828);
and U4856 (N_4856,N_1260,N_2793);
and U4857 (N_4857,N_354,N_1532);
or U4858 (N_4858,N_492,N_1562);
or U4859 (N_4859,N_2883,N_851);
and U4860 (N_4860,N_2415,N_1021);
and U4861 (N_4861,N_943,N_369);
nor U4862 (N_4862,N_252,N_160);
nand U4863 (N_4863,N_2138,N_1714);
nand U4864 (N_4864,N_385,N_402);
nor U4865 (N_4865,N_1908,N_1872);
nor U4866 (N_4866,N_1085,N_234);
nor U4867 (N_4867,N_1108,N_2062);
nor U4868 (N_4868,N_616,N_2666);
and U4869 (N_4869,N_2854,N_2108);
nand U4870 (N_4870,N_1614,N_415);
nor U4871 (N_4871,N_1111,N_2035);
and U4872 (N_4872,N_2518,N_289);
nand U4873 (N_4873,N_152,N_2200);
nor U4874 (N_4874,N_2441,N_4);
and U4875 (N_4875,N_1561,N_2228);
and U4876 (N_4876,N_2714,N_766);
nand U4877 (N_4877,N_866,N_1769);
and U4878 (N_4878,N_671,N_325);
or U4879 (N_4879,N_2495,N_2993);
and U4880 (N_4880,N_934,N_902);
nor U4881 (N_4881,N_372,N_351);
nor U4882 (N_4882,N_1009,N_2022);
nor U4883 (N_4883,N_1181,N_774);
nand U4884 (N_4884,N_355,N_653);
nand U4885 (N_4885,N_927,N_955);
or U4886 (N_4886,N_2364,N_2354);
nor U4887 (N_4887,N_767,N_2479);
nor U4888 (N_4888,N_74,N_1326);
nor U4889 (N_4889,N_2479,N_1021);
nor U4890 (N_4890,N_1580,N_2300);
nor U4891 (N_4891,N_2321,N_1953);
or U4892 (N_4892,N_824,N_2950);
nand U4893 (N_4893,N_2414,N_2248);
nor U4894 (N_4894,N_48,N_1470);
and U4895 (N_4895,N_910,N_878);
nor U4896 (N_4896,N_2173,N_390);
xor U4897 (N_4897,N_1214,N_2921);
or U4898 (N_4898,N_715,N_2241);
and U4899 (N_4899,N_1715,N_504);
and U4900 (N_4900,N_2741,N_517);
or U4901 (N_4901,N_1722,N_808);
xor U4902 (N_4902,N_1855,N_2045);
nand U4903 (N_4903,N_2470,N_30);
and U4904 (N_4904,N_2612,N_275);
nand U4905 (N_4905,N_2751,N_441);
nand U4906 (N_4906,N_2502,N_1581);
and U4907 (N_4907,N_2516,N_2695);
nand U4908 (N_4908,N_643,N_2151);
nand U4909 (N_4909,N_1459,N_2733);
and U4910 (N_4910,N_2690,N_2472);
nor U4911 (N_4911,N_2323,N_1495);
and U4912 (N_4912,N_514,N_1322);
nand U4913 (N_4913,N_1930,N_2065);
nor U4914 (N_4914,N_2586,N_697);
nor U4915 (N_4915,N_1975,N_62);
or U4916 (N_4916,N_1701,N_2310);
and U4917 (N_4917,N_778,N_1550);
or U4918 (N_4918,N_1803,N_2613);
or U4919 (N_4919,N_697,N_1467);
nand U4920 (N_4920,N_458,N_2110);
nor U4921 (N_4921,N_1361,N_753);
nor U4922 (N_4922,N_1721,N_2606);
nand U4923 (N_4923,N_656,N_1745);
and U4924 (N_4924,N_2097,N_1666);
nor U4925 (N_4925,N_84,N_26);
or U4926 (N_4926,N_2444,N_858);
and U4927 (N_4927,N_1368,N_310);
and U4928 (N_4928,N_1021,N_232);
nor U4929 (N_4929,N_158,N_1501);
or U4930 (N_4930,N_384,N_2048);
nand U4931 (N_4931,N_2629,N_2581);
and U4932 (N_4932,N_2597,N_1618);
or U4933 (N_4933,N_2652,N_2840);
or U4934 (N_4934,N_984,N_702);
and U4935 (N_4935,N_2851,N_2758);
and U4936 (N_4936,N_1179,N_1299);
nand U4937 (N_4937,N_311,N_1442);
and U4938 (N_4938,N_2486,N_1920);
or U4939 (N_4939,N_2719,N_2353);
or U4940 (N_4940,N_705,N_849);
or U4941 (N_4941,N_1103,N_2109);
and U4942 (N_4942,N_1134,N_2471);
nand U4943 (N_4943,N_692,N_890);
or U4944 (N_4944,N_2930,N_300);
or U4945 (N_4945,N_48,N_503);
and U4946 (N_4946,N_1507,N_2724);
nor U4947 (N_4947,N_286,N_2427);
or U4948 (N_4948,N_2928,N_744);
nor U4949 (N_4949,N_200,N_799);
nand U4950 (N_4950,N_2739,N_895);
and U4951 (N_4951,N_2070,N_593);
nand U4952 (N_4952,N_2508,N_2471);
or U4953 (N_4953,N_108,N_1146);
nor U4954 (N_4954,N_1905,N_2564);
xor U4955 (N_4955,N_2136,N_980);
and U4956 (N_4956,N_1333,N_302);
nand U4957 (N_4957,N_2402,N_2328);
nand U4958 (N_4958,N_1306,N_295);
nand U4959 (N_4959,N_336,N_2845);
and U4960 (N_4960,N_371,N_2073);
or U4961 (N_4961,N_1115,N_756);
nor U4962 (N_4962,N_1958,N_1557);
xnor U4963 (N_4963,N_1924,N_112);
and U4964 (N_4964,N_2875,N_1614);
nand U4965 (N_4965,N_2001,N_2042);
and U4966 (N_4966,N_692,N_770);
xor U4967 (N_4967,N_891,N_448);
and U4968 (N_4968,N_814,N_999);
xnor U4969 (N_4969,N_618,N_2242);
or U4970 (N_4970,N_2021,N_2505);
and U4971 (N_4971,N_1330,N_2061);
and U4972 (N_4972,N_1744,N_212);
nor U4973 (N_4973,N_1198,N_440);
or U4974 (N_4974,N_928,N_853);
xor U4975 (N_4975,N_1374,N_1790);
nand U4976 (N_4976,N_2125,N_1263);
xor U4977 (N_4977,N_1926,N_1816);
xor U4978 (N_4978,N_1152,N_1798);
and U4979 (N_4979,N_2221,N_1089);
xnor U4980 (N_4980,N_2060,N_2955);
nand U4981 (N_4981,N_2973,N_1497);
or U4982 (N_4982,N_359,N_601);
or U4983 (N_4983,N_2113,N_1660);
and U4984 (N_4984,N_71,N_1917);
nand U4985 (N_4985,N_2915,N_1085);
nor U4986 (N_4986,N_756,N_1821);
or U4987 (N_4987,N_328,N_2742);
nor U4988 (N_4988,N_2906,N_1813);
or U4989 (N_4989,N_505,N_1077);
nand U4990 (N_4990,N_2508,N_1882);
or U4991 (N_4991,N_898,N_1558);
nor U4992 (N_4992,N_1463,N_2182);
nor U4993 (N_4993,N_937,N_2796);
nor U4994 (N_4994,N_1861,N_1332);
or U4995 (N_4995,N_1876,N_1715);
nand U4996 (N_4996,N_302,N_1314);
or U4997 (N_4997,N_1711,N_1859);
nor U4998 (N_4998,N_2929,N_557);
and U4999 (N_4999,N_2007,N_2098);
nor U5000 (N_5000,N_852,N_1747);
xnor U5001 (N_5001,N_1583,N_1822);
nor U5002 (N_5002,N_2868,N_424);
nor U5003 (N_5003,N_2729,N_2072);
nand U5004 (N_5004,N_1280,N_832);
or U5005 (N_5005,N_317,N_2647);
nand U5006 (N_5006,N_132,N_2858);
xor U5007 (N_5007,N_2080,N_2150);
nand U5008 (N_5008,N_2127,N_1965);
nor U5009 (N_5009,N_1330,N_726);
nand U5010 (N_5010,N_1170,N_249);
or U5011 (N_5011,N_2873,N_1012);
and U5012 (N_5012,N_179,N_2046);
and U5013 (N_5013,N_1960,N_100);
nor U5014 (N_5014,N_2359,N_2058);
or U5015 (N_5015,N_863,N_464);
nand U5016 (N_5016,N_2142,N_1628);
nand U5017 (N_5017,N_1067,N_2534);
nand U5018 (N_5018,N_461,N_2717);
or U5019 (N_5019,N_1024,N_2109);
nand U5020 (N_5020,N_2604,N_1439);
nand U5021 (N_5021,N_1342,N_2218);
and U5022 (N_5022,N_964,N_2279);
or U5023 (N_5023,N_880,N_2326);
and U5024 (N_5024,N_2248,N_2095);
or U5025 (N_5025,N_649,N_1746);
nand U5026 (N_5026,N_690,N_1613);
nor U5027 (N_5027,N_1047,N_2422);
or U5028 (N_5028,N_2166,N_639);
xor U5029 (N_5029,N_2911,N_1776);
xnor U5030 (N_5030,N_2775,N_732);
nor U5031 (N_5031,N_2550,N_2353);
xor U5032 (N_5032,N_103,N_2469);
nand U5033 (N_5033,N_2960,N_2822);
or U5034 (N_5034,N_670,N_584);
or U5035 (N_5035,N_390,N_31);
or U5036 (N_5036,N_1175,N_2589);
xnor U5037 (N_5037,N_2714,N_342);
nand U5038 (N_5038,N_444,N_1394);
xnor U5039 (N_5039,N_2772,N_2046);
nand U5040 (N_5040,N_2767,N_1285);
and U5041 (N_5041,N_2934,N_1188);
nand U5042 (N_5042,N_876,N_2506);
xnor U5043 (N_5043,N_1863,N_96);
and U5044 (N_5044,N_1214,N_787);
and U5045 (N_5045,N_1723,N_2144);
nand U5046 (N_5046,N_724,N_2906);
nor U5047 (N_5047,N_2103,N_2571);
and U5048 (N_5048,N_1756,N_1766);
and U5049 (N_5049,N_1541,N_2792);
and U5050 (N_5050,N_948,N_608);
and U5051 (N_5051,N_1349,N_2832);
or U5052 (N_5052,N_2225,N_1016);
nand U5053 (N_5053,N_1357,N_1607);
or U5054 (N_5054,N_1775,N_1046);
and U5055 (N_5055,N_1941,N_2180);
and U5056 (N_5056,N_2935,N_2416);
or U5057 (N_5057,N_101,N_1495);
nand U5058 (N_5058,N_2342,N_953);
or U5059 (N_5059,N_2459,N_1690);
and U5060 (N_5060,N_2882,N_307);
or U5061 (N_5061,N_2217,N_1375);
and U5062 (N_5062,N_708,N_2787);
and U5063 (N_5063,N_648,N_622);
and U5064 (N_5064,N_1468,N_2016);
nor U5065 (N_5065,N_171,N_139);
and U5066 (N_5066,N_961,N_1633);
and U5067 (N_5067,N_1060,N_2708);
nor U5068 (N_5068,N_2120,N_954);
and U5069 (N_5069,N_1149,N_188);
and U5070 (N_5070,N_275,N_482);
nand U5071 (N_5071,N_2940,N_1217);
nor U5072 (N_5072,N_2325,N_1204);
nand U5073 (N_5073,N_1501,N_1441);
and U5074 (N_5074,N_371,N_356);
nor U5075 (N_5075,N_869,N_1584);
xor U5076 (N_5076,N_804,N_1564);
nor U5077 (N_5077,N_2178,N_79);
or U5078 (N_5078,N_2275,N_2350);
or U5079 (N_5079,N_1991,N_2219);
nand U5080 (N_5080,N_591,N_1284);
or U5081 (N_5081,N_458,N_2035);
or U5082 (N_5082,N_2,N_2796);
xnor U5083 (N_5083,N_2507,N_2418);
or U5084 (N_5084,N_1249,N_969);
nor U5085 (N_5085,N_2789,N_2347);
or U5086 (N_5086,N_1675,N_2824);
or U5087 (N_5087,N_704,N_1404);
nand U5088 (N_5088,N_575,N_2826);
xnor U5089 (N_5089,N_1822,N_1036);
nor U5090 (N_5090,N_764,N_2456);
nand U5091 (N_5091,N_867,N_800);
or U5092 (N_5092,N_1924,N_1858);
nor U5093 (N_5093,N_1667,N_2381);
or U5094 (N_5094,N_16,N_1688);
and U5095 (N_5095,N_262,N_1098);
nor U5096 (N_5096,N_2706,N_8);
or U5097 (N_5097,N_2748,N_2662);
and U5098 (N_5098,N_668,N_254);
nor U5099 (N_5099,N_2747,N_1818);
nor U5100 (N_5100,N_2991,N_1162);
nor U5101 (N_5101,N_2725,N_305);
nand U5102 (N_5102,N_2002,N_1756);
and U5103 (N_5103,N_2805,N_1293);
nor U5104 (N_5104,N_1982,N_1110);
or U5105 (N_5105,N_1995,N_472);
nand U5106 (N_5106,N_2561,N_804);
nand U5107 (N_5107,N_1004,N_66);
nand U5108 (N_5108,N_1010,N_371);
or U5109 (N_5109,N_2928,N_1994);
xnor U5110 (N_5110,N_923,N_1722);
nor U5111 (N_5111,N_854,N_136);
nor U5112 (N_5112,N_1062,N_2143);
or U5113 (N_5113,N_1509,N_2898);
or U5114 (N_5114,N_2302,N_2538);
nand U5115 (N_5115,N_1568,N_2529);
nor U5116 (N_5116,N_378,N_1536);
or U5117 (N_5117,N_708,N_2105);
xor U5118 (N_5118,N_278,N_1117);
or U5119 (N_5119,N_2344,N_765);
nand U5120 (N_5120,N_1294,N_2742);
xor U5121 (N_5121,N_2250,N_134);
and U5122 (N_5122,N_2636,N_2090);
or U5123 (N_5123,N_1813,N_2056);
nand U5124 (N_5124,N_1961,N_1253);
or U5125 (N_5125,N_2,N_319);
or U5126 (N_5126,N_2741,N_925);
nand U5127 (N_5127,N_1674,N_1107);
xor U5128 (N_5128,N_2216,N_2098);
nor U5129 (N_5129,N_1364,N_560);
xor U5130 (N_5130,N_2097,N_1395);
xor U5131 (N_5131,N_1715,N_1606);
nand U5132 (N_5132,N_77,N_1831);
nor U5133 (N_5133,N_1448,N_2934);
or U5134 (N_5134,N_2140,N_770);
xnor U5135 (N_5135,N_2531,N_1841);
nor U5136 (N_5136,N_2522,N_2739);
or U5137 (N_5137,N_477,N_42);
or U5138 (N_5138,N_377,N_2440);
xor U5139 (N_5139,N_1671,N_1906);
and U5140 (N_5140,N_2594,N_2772);
or U5141 (N_5141,N_1536,N_60);
and U5142 (N_5142,N_2352,N_209);
or U5143 (N_5143,N_1121,N_642);
nor U5144 (N_5144,N_1203,N_2401);
nand U5145 (N_5145,N_705,N_1289);
and U5146 (N_5146,N_2930,N_1065);
nor U5147 (N_5147,N_1380,N_1491);
or U5148 (N_5148,N_1112,N_1594);
and U5149 (N_5149,N_609,N_2197);
or U5150 (N_5150,N_2108,N_2179);
nor U5151 (N_5151,N_393,N_944);
nor U5152 (N_5152,N_706,N_31);
and U5153 (N_5153,N_2319,N_1823);
nand U5154 (N_5154,N_935,N_2808);
nand U5155 (N_5155,N_2428,N_402);
nand U5156 (N_5156,N_1091,N_392);
and U5157 (N_5157,N_1767,N_642);
xnor U5158 (N_5158,N_1492,N_2555);
nor U5159 (N_5159,N_2286,N_712);
nor U5160 (N_5160,N_81,N_2908);
nand U5161 (N_5161,N_831,N_1765);
nor U5162 (N_5162,N_2381,N_2021);
nand U5163 (N_5163,N_105,N_2163);
or U5164 (N_5164,N_1912,N_165);
nor U5165 (N_5165,N_2121,N_1585);
nor U5166 (N_5166,N_44,N_494);
and U5167 (N_5167,N_1680,N_2113);
or U5168 (N_5168,N_2955,N_1195);
nor U5169 (N_5169,N_1578,N_217);
and U5170 (N_5170,N_2936,N_791);
or U5171 (N_5171,N_1048,N_1757);
nor U5172 (N_5172,N_1534,N_986);
and U5173 (N_5173,N_2968,N_499);
or U5174 (N_5174,N_692,N_1983);
nor U5175 (N_5175,N_1744,N_1172);
xnor U5176 (N_5176,N_706,N_2397);
or U5177 (N_5177,N_1422,N_1339);
and U5178 (N_5178,N_2269,N_1046);
or U5179 (N_5179,N_2273,N_515);
or U5180 (N_5180,N_2266,N_629);
or U5181 (N_5181,N_1460,N_137);
nor U5182 (N_5182,N_1429,N_576);
nor U5183 (N_5183,N_621,N_165);
and U5184 (N_5184,N_2244,N_84);
or U5185 (N_5185,N_2654,N_2076);
nor U5186 (N_5186,N_2731,N_2901);
or U5187 (N_5187,N_697,N_2414);
nand U5188 (N_5188,N_2945,N_1608);
or U5189 (N_5189,N_561,N_1422);
nor U5190 (N_5190,N_2645,N_2943);
xor U5191 (N_5191,N_570,N_1915);
xor U5192 (N_5192,N_965,N_1853);
and U5193 (N_5193,N_2020,N_1538);
or U5194 (N_5194,N_2513,N_2391);
nor U5195 (N_5195,N_1028,N_1460);
nand U5196 (N_5196,N_87,N_1104);
xor U5197 (N_5197,N_2925,N_2988);
nand U5198 (N_5198,N_979,N_1331);
and U5199 (N_5199,N_1519,N_854);
nand U5200 (N_5200,N_2727,N_364);
or U5201 (N_5201,N_2544,N_295);
and U5202 (N_5202,N_35,N_758);
or U5203 (N_5203,N_1238,N_2905);
or U5204 (N_5204,N_1319,N_940);
or U5205 (N_5205,N_2175,N_256);
and U5206 (N_5206,N_2941,N_1487);
or U5207 (N_5207,N_837,N_2747);
nor U5208 (N_5208,N_2824,N_1378);
nand U5209 (N_5209,N_2940,N_1188);
nor U5210 (N_5210,N_172,N_2907);
and U5211 (N_5211,N_261,N_443);
or U5212 (N_5212,N_151,N_1514);
nand U5213 (N_5213,N_315,N_2498);
or U5214 (N_5214,N_2052,N_1868);
or U5215 (N_5215,N_2504,N_1037);
nand U5216 (N_5216,N_1664,N_2948);
xor U5217 (N_5217,N_601,N_542);
nor U5218 (N_5218,N_213,N_388);
nand U5219 (N_5219,N_2617,N_2492);
nor U5220 (N_5220,N_2280,N_2489);
nor U5221 (N_5221,N_53,N_247);
or U5222 (N_5222,N_2516,N_693);
nand U5223 (N_5223,N_1009,N_2290);
and U5224 (N_5224,N_329,N_694);
or U5225 (N_5225,N_840,N_590);
nor U5226 (N_5226,N_1559,N_2135);
nand U5227 (N_5227,N_811,N_1615);
nor U5228 (N_5228,N_1533,N_1827);
nor U5229 (N_5229,N_2824,N_2306);
nor U5230 (N_5230,N_2971,N_2060);
nor U5231 (N_5231,N_2856,N_2851);
nor U5232 (N_5232,N_2267,N_767);
or U5233 (N_5233,N_2095,N_2540);
nand U5234 (N_5234,N_1166,N_1091);
xor U5235 (N_5235,N_1183,N_2787);
nand U5236 (N_5236,N_2806,N_314);
nor U5237 (N_5237,N_2100,N_1612);
or U5238 (N_5238,N_2418,N_1227);
nor U5239 (N_5239,N_380,N_1784);
xor U5240 (N_5240,N_187,N_415);
nor U5241 (N_5241,N_2728,N_1562);
nor U5242 (N_5242,N_1704,N_2769);
and U5243 (N_5243,N_2920,N_2286);
and U5244 (N_5244,N_1773,N_2513);
nor U5245 (N_5245,N_1682,N_759);
or U5246 (N_5246,N_1431,N_1653);
nor U5247 (N_5247,N_346,N_2874);
and U5248 (N_5248,N_2682,N_1924);
nor U5249 (N_5249,N_2428,N_2271);
nand U5250 (N_5250,N_1640,N_32);
nand U5251 (N_5251,N_291,N_2784);
nor U5252 (N_5252,N_345,N_1003);
and U5253 (N_5253,N_2247,N_383);
and U5254 (N_5254,N_2398,N_1734);
or U5255 (N_5255,N_2732,N_1100);
nand U5256 (N_5256,N_3,N_2793);
and U5257 (N_5257,N_2695,N_2606);
xor U5258 (N_5258,N_2663,N_2850);
nor U5259 (N_5259,N_26,N_772);
nor U5260 (N_5260,N_949,N_440);
nor U5261 (N_5261,N_48,N_1123);
nor U5262 (N_5262,N_1539,N_461);
nand U5263 (N_5263,N_1308,N_1473);
and U5264 (N_5264,N_309,N_1933);
nor U5265 (N_5265,N_1178,N_2083);
or U5266 (N_5266,N_2863,N_2076);
or U5267 (N_5267,N_2508,N_2509);
nand U5268 (N_5268,N_765,N_1086);
xnor U5269 (N_5269,N_2604,N_1405);
nor U5270 (N_5270,N_1219,N_752);
nor U5271 (N_5271,N_22,N_2738);
nand U5272 (N_5272,N_2753,N_1501);
or U5273 (N_5273,N_1393,N_525);
nand U5274 (N_5274,N_2077,N_2469);
or U5275 (N_5275,N_1124,N_2871);
and U5276 (N_5276,N_500,N_531);
and U5277 (N_5277,N_1171,N_2651);
xnor U5278 (N_5278,N_856,N_2146);
or U5279 (N_5279,N_1493,N_1124);
nor U5280 (N_5280,N_1832,N_1718);
and U5281 (N_5281,N_1804,N_2822);
nor U5282 (N_5282,N_32,N_327);
nor U5283 (N_5283,N_2523,N_316);
or U5284 (N_5284,N_2742,N_820);
nand U5285 (N_5285,N_896,N_793);
or U5286 (N_5286,N_1544,N_2669);
nand U5287 (N_5287,N_1689,N_2590);
nor U5288 (N_5288,N_1802,N_123);
xor U5289 (N_5289,N_2223,N_776);
and U5290 (N_5290,N_1782,N_2638);
and U5291 (N_5291,N_1152,N_2139);
or U5292 (N_5292,N_1250,N_1234);
or U5293 (N_5293,N_2811,N_510);
nor U5294 (N_5294,N_2976,N_1064);
and U5295 (N_5295,N_2164,N_2263);
nor U5296 (N_5296,N_487,N_2128);
or U5297 (N_5297,N_1938,N_546);
nor U5298 (N_5298,N_2937,N_2863);
nor U5299 (N_5299,N_1723,N_1220);
nand U5300 (N_5300,N_74,N_2472);
nand U5301 (N_5301,N_53,N_246);
and U5302 (N_5302,N_2914,N_4);
and U5303 (N_5303,N_371,N_1918);
and U5304 (N_5304,N_2532,N_2371);
or U5305 (N_5305,N_1209,N_2973);
nand U5306 (N_5306,N_2887,N_1827);
nor U5307 (N_5307,N_2532,N_2971);
or U5308 (N_5308,N_429,N_1582);
and U5309 (N_5309,N_1111,N_878);
xnor U5310 (N_5310,N_484,N_1720);
nor U5311 (N_5311,N_617,N_2705);
and U5312 (N_5312,N_2125,N_717);
nor U5313 (N_5313,N_2605,N_2896);
nor U5314 (N_5314,N_1779,N_1973);
or U5315 (N_5315,N_1811,N_908);
or U5316 (N_5316,N_365,N_911);
or U5317 (N_5317,N_2231,N_473);
nor U5318 (N_5318,N_2598,N_2746);
nor U5319 (N_5319,N_1240,N_897);
or U5320 (N_5320,N_1824,N_2539);
or U5321 (N_5321,N_1057,N_2912);
nor U5322 (N_5322,N_951,N_141);
xnor U5323 (N_5323,N_2391,N_743);
xnor U5324 (N_5324,N_2225,N_2147);
and U5325 (N_5325,N_2825,N_268);
xnor U5326 (N_5326,N_2122,N_296);
nand U5327 (N_5327,N_541,N_0);
and U5328 (N_5328,N_655,N_407);
nand U5329 (N_5329,N_2042,N_1581);
nand U5330 (N_5330,N_2673,N_938);
xnor U5331 (N_5331,N_1920,N_2155);
or U5332 (N_5332,N_1204,N_2151);
nand U5333 (N_5333,N_858,N_2370);
and U5334 (N_5334,N_670,N_2029);
and U5335 (N_5335,N_2364,N_2179);
and U5336 (N_5336,N_727,N_1498);
and U5337 (N_5337,N_2079,N_970);
nand U5338 (N_5338,N_2520,N_1449);
and U5339 (N_5339,N_617,N_1848);
nand U5340 (N_5340,N_2955,N_317);
or U5341 (N_5341,N_442,N_104);
xnor U5342 (N_5342,N_1913,N_1094);
nor U5343 (N_5343,N_2692,N_1448);
nand U5344 (N_5344,N_15,N_926);
and U5345 (N_5345,N_2310,N_1507);
and U5346 (N_5346,N_1755,N_1427);
nand U5347 (N_5347,N_1351,N_2473);
or U5348 (N_5348,N_1744,N_1312);
or U5349 (N_5349,N_1637,N_1966);
nand U5350 (N_5350,N_369,N_1949);
and U5351 (N_5351,N_2118,N_2524);
nand U5352 (N_5352,N_2279,N_663);
or U5353 (N_5353,N_772,N_1736);
or U5354 (N_5354,N_2537,N_1678);
xor U5355 (N_5355,N_2349,N_2727);
or U5356 (N_5356,N_251,N_151);
or U5357 (N_5357,N_1903,N_1447);
and U5358 (N_5358,N_2829,N_1210);
nand U5359 (N_5359,N_1659,N_1526);
and U5360 (N_5360,N_589,N_2280);
nor U5361 (N_5361,N_334,N_1288);
nor U5362 (N_5362,N_1231,N_1669);
nand U5363 (N_5363,N_2376,N_2265);
or U5364 (N_5364,N_2123,N_362);
and U5365 (N_5365,N_605,N_1194);
nand U5366 (N_5366,N_1357,N_935);
xor U5367 (N_5367,N_2611,N_2131);
and U5368 (N_5368,N_625,N_1136);
nand U5369 (N_5369,N_2819,N_2706);
and U5370 (N_5370,N_847,N_2189);
nor U5371 (N_5371,N_2836,N_2994);
nor U5372 (N_5372,N_478,N_957);
nand U5373 (N_5373,N_1697,N_666);
or U5374 (N_5374,N_808,N_960);
and U5375 (N_5375,N_1756,N_1312);
and U5376 (N_5376,N_1022,N_1920);
or U5377 (N_5377,N_2859,N_2855);
or U5378 (N_5378,N_2221,N_2130);
nand U5379 (N_5379,N_2945,N_1755);
nand U5380 (N_5380,N_1475,N_207);
or U5381 (N_5381,N_1208,N_950);
nor U5382 (N_5382,N_2086,N_1707);
nor U5383 (N_5383,N_1084,N_1843);
nand U5384 (N_5384,N_784,N_2553);
nor U5385 (N_5385,N_2258,N_475);
xnor U5386 (N_5386,N_652,N_2214);
xor U5387 (N_5387,N_500,N_203);
or U5388 (N_5388,N_1618,N_858);
xnor U5389 (N_5389,N_2116,N_1307);
xor U5390 (N_5390,N_1891,N_1988);
and U5391 (N_5391,N_2202,N_819);
xnor U5392 (N_5392,N_2808,N_562);
nor U5393 (N_5393,N_520,N_607);
nor U5394 (N_5394,N_1517,N_118);
or U5395 (N_5395,N_1949,N_1177);
xnor U5396 (N_5396,N_1150,N_2086);
nor U5397 (N_5397,N_2121,N_906);
and U5398 (N_5398,N_463,N_1916);
and U5399 (N_5399,N_2382,N_1853);
or U5400 (N_5400,N_2052,N_2151);
nand U5401 (N_5401,N_1106,N_2379);
nand U5402 (N_5402,N_2357,N_2636);
and U5403 (N_5403,N_1171,N_1667);
and U5404 (N_5404,N_2329,N_1396);
nor U5405 (N_5405,N_2763,N_660);
and U5406 (N_5406,N_1692,N_745);
nand U5407 (N_5407,N_2467,N_93);
or U5408 (N_5408,N_263,N_1377);
or U5409 (N_5409,N_2124,N_1338);
or U5410 (N_5410,N_865,N_2144);
and U5411 (N_5411,N_512,N_2663);
and U5412 (N_5412,N_937,N_849);
xnor U5413 (N_5413,N_1107,N_2000);
or U5414 (N_5414,N_2914,N_1967);
and U5415 (N_5415,N_828,N_2098);
nor U5416 (N_5416,N_1997,N_1728);
and U5417 (N_5417,N_2890,N_1235);
or U5418 (N_5418,N_189,N_2533);
nand U5419 (N_5419,N_1181,N_1067);
nand U5420 (N_5420,N_28,N_2163);
xnor U5421 (N_5421,N_212,N_786);
nand U5422 (N_5422,N_1621,N_1791);
nand U5423 (N_5423,N_2135,N_1533);
or U5424 (N_5424,N_780,N_587);
nand U5425 (N_5425,N_1002,N_891);
and U5426 (N_5426,N_2550,N_2689);
nand U5427 (N_5427,N_1289,N_2917);
and U5428 (N_5428,N_1071,N_406);
nand U5429 (N_5429,N_814,N_304);
nor U5430 (N_5430,N_18,N_2635);
nand U5431 (N_5431,N_600,N_1889);
and U5432 (N_5432,N_591,N_667);
and U5433 (N_5433,N_950,N_2745);
and U5434 (N_5434,N_1456,N_2319);
and U5435 (N_5435,N_2715,N_197);
and U5436 (N_5436,N_1537,N_319);
xnor U5437 (N_5437,N_1222,N_905);
or U5438 (N_5438,N_656,N_1831);
nor U5439 (N_5439,N_1354,N_623);
nand U5440 (N_5440,N_1765,N_2997);
and U5441 (N_5441,N_1210,N_2803);
and U5442 (N_5442,N_2721,N_1631);
nor U5443 (N_5443,N_734,N_1661);
nor U5444 (N_5444,N_2677,N_2225);
nor U5445 (N_5445,N_1503,N_2732);
nor U5446 (N_5446,N_2712,N_1964);
or U5447 (N_5447,N_1404,N_2607);
xor U5448 (N_5448,N_541,N_1053);
nor U5449 (N_5449,N_2776,N_2015);
nand U5450 (N_5450,N_1368,N_17);
nor U5451 (N_5451,N_2334,N_2933);
nor U5452 (N_5452,N_1429,N_2823);
nor U5453 (N_5453,N_321,N_2676);
nor U5454 (N_5454,N_730,N_896);
nor U5455 (N_5455,N_2975,N_1333);
nor U5456 (N_5456,N_1052,N_805);
nand U5457 (N_5457,N_911,N_1021);
and U5458 (N_5458,N_625,N_2635);
and U5459 (N_5459,N_929,N_2670);
and U5460 (N_5460,N_1346,N_2235);
nand U5461 (N_5461,N_2946,N_829);
and U5462 (N_5462,N_273,N_478);
or U5463 (N_5463,N_1049,N_2739);
nor U5464 (N_5464,N_687,N_2813);
and U5465 (N_5465,N_1761,N_1850);
or U5466 (N_5466,N_1530,N_2099);
and U5467 (N_5467,N_418,N_2402);
or U5468 (N_5468,N_1512,N_431);
and U5469 (N_5469,N_1869,N_322);
and U5470 (N_5470,N_1618,N_2917);
or U5471 (N_5471,N_1286,N_1514);
nand U5472 (N_5472,N_610,N_1689);
or U5473 (N_5473,N_1565,N_2345);
and U5474 (N_5474,N_418,N_2630);
nand U5475 (N_5475,N_1088,N_1647);
or U5476 (N_5476,N_2245,N_166);
nor U5477 (N_5477,N_2922,N_798);
or U5478 (N_5478,N_2372,N_735);
nand U5479 (N_5479,N_1343,N_1689);
nor U5480 (N_5480,N_676,N_1319);
and U5481 (N_5481,N_1087,N_1934);
nor U5482 (N_5482,N_819,N_1179);
and U5483 (N_5483,N_2327,N_2440);
nand U5484 (N_5484,N_2820,N_2039);
and U5485 (N_5485,N_2386,N_1548);
nor U5486 (N_5486,N_1362,N_2362);
or U5487 (N_5487,N_90,N_395);
nor U5488 (N_5488,N_370,N_2791);
and U5489 (N_5489,N_212,N_1750);
nand U5490 (N_5490,N_130,N_2923);
nor U5491 (N_5491,N_1004,N_886);
nand U5492 (N_5492,N_2311,N_166);
nor U5493 (N_5493,N_1566,N_2063);
and U5494 (N_5494,N_245,N_401);
and U5495 (N_5495,N_1977,N_1571);
and U5496 (N_5496,N_933,N_1620);
or U5497 (N_5497,N_1809,N_1623);
or U5498 (N_5498,N_405,N_1989);
and U5499 (N_5499,N_1554,N_1304);
and U5500 (N_5500,N_1720,N_798);
nor U5501 (N_5501,N_684,N_2700);
nand U5502 (N_5502,N_1003,N_60);
nor U5503 (N_5503,N_613,N_729);
nand U5504 (N_5504,N_932,N_1945);
nor U5505 (N_5505,N_43,N_1323);
or U5506 (N_5506,N_240,N_2584);
xnor U5507 (N_5507,N_379,N_610);
and U5508 (N_5508,N_1730,N_453);
nand U5509 (N_5509,N_924,N_2335);
or U5510 (N_5510,N_2560,N_2062);
or U5511 (N_5511,N_2607,N_2352);
nand U5512 (N_5512,N_1940,N_1243);
or U5513 (N_5513,N_1649,N_1106);
or U5514 (N_5514,N_688,N_727);
and U5515 (N_5515,N_674,N_1192);
nand U5516 (N_5516,N_1434,N_2465);
or U5517 (N_5517,N_2293,N_1518);
nor U5518 (N_5518,N_2161,N_1665);
nor U5519 (N_5519,N_1872,N_935);
nor U5520 (N_5520,N_1328,N_1382);
nand U5521 (N_5521,N_322,N_2548);
nand U5522 (N_5522,N_599,N_1488);
xnor U5523 (N_5523,N_448,N_378);
nand U5524 (N_5524,N_1827,N_941);
and U5525 (N_5525,N_105,N_440);
or U5526 (N_5526,N_727,N_969);
xnor U5527 (N_5527,N_1717,N_2015);
xnor U5528 (N_5528,N_2141,N_1620);
or U5529 (N_5529,N_791,N_1655);
xnor U5530 (N_5530,N_2552,N_2943);
or U5531 (N_5531,N_637,N_2236);
xnor U5532 (N_5532,N_1535,N_1351);
or U5533 (N_5533,N_928,N_840);
nand U5534 (N_5534,N_116,N_2655);
and U5535 (N_5535,N_2609,N_744);
xor U5536 (N_5536,N_849,N_2179);
nand U5537 (N_5537,N_1970,N_2817);
nand U5538 (N_5538,N_1497,N_62);
and U5539 (N_5539,N_2759,N_2594);
nand U5540 (N_5540,N_466,N_1834);
and U5541 (N_5541,N_385,N_2976);
and U5542 (N_5542,N_2504,N_2321);
and U5543 (N_5543,N_78,N_1914);
or U5544 (N_5544,N_2647,N_1147);
or U5545 (N_5545,N_926,N_1369);
and U5546 (N_5546,N_125,N_607);
nand U5547 (N_5547,N_2781,N_724);
and U5548 (N_5548,N_2709,N_1539);
nor U5549 (N_5549,N_343,N_2227);
or U5550 (N_5550,N_45,N_1555);
and U5551 (N_5551,N_675,N_1223);
or U5552 (N_5552,N_2309,N_650);
and U5553 (N_5553,N_1193,N_2796);
or U5554 (N_5554,N_1291,N_1547);
nand U5555 (N_5555,N_1347,N_2964);
nor U5556 (N_5556,N_936,N_2811);
and U5557 (N_5557,N_640,N_2775);
nor U5558 (N_5558,N_204,N_1773);
xnor U5559 (N_5559,N_1480,N_1840);
or U5560 (N_5560,N_2262,N_1739);
or U5561 (N_5561,N_1073,N_2915);
nand U5562 (N_5562,N_2856,N_584);
or U5563 (N_5563,N_2630,N_136);
and U5564 (N_5564,N_273,N_420);
or U5565 (N_5565,N_757,N_2502);
nand U5566 (N_5566,N_2436,N_2529);
and U5567 (N_5567,N_2915,N_2628);
nor U5568 (N_5568,N_1886,N_480);
nor U5569 (N_5569,N_2415,N_1732);
and U5570 (N_5570,N_1550,N_74);
xor U5571 (N_5571,N_1531,N_1996);
nand U5572 (N_5572,N_2652,N_1273);
nor U5573 (N_5573,N_933,N_321);
and U5574 (N_5574,N_2230,N_2815);
nor U5575 (N_5575,N_1107,N_1408);
or U5576 (N_5576,N_2230,N_2431);
and U5577 (N_5577,N_1254,N_2291);
nand U5578 (N_5578,N_1863,N_2895);
and U5579 (N_5579,N_2831,N_2485);
nor U5580 (N_5580,N_38,N_986);
nor U5581 (N_5581,N_2091,N_2846);
or U5582 (N_5582,N_105,N_2612);
nand U5583 (N_5583,N_2692,N_2975);
nand U5584 (N_5584,N_420,N_646);
xnor U5585 (N_5585,N_1856,N_2964);
nand U5586 (N_5586,N_37,N_1582);
or U5587 (N_5587,N_2313,N_804);
or U5588 (N_5588,N_104,N_555);
nand U5589 (N_5589,N_1104,N_1278);
xnor U5590 (N_5590,N_2538,N_726);
nor U5591 (N_5591,N_2326,N_2643);
nor U5592 (N_5592,N_2907,N_364);
nor U5593 (N_5593,N_1863,N_2554);
nand U5594 (N_5594,N_603,N_1187);
nand U5595 (N_5595,N_982,N_2415);
or U5596 (N_5596,N_809,N_2918);
nand U5597 (N_5597,N_1312,N_2077);
nand U5598 (N_5598,N_431,N_2876);
nor U5599 (N_5599,N_1835,N_831);
nand U5600 (N_5600,N_1715,N_2145);
nand U5601 (N_5601,N_1833,N_825);
nand U5602 (N_5602,N_1055,N_2728);
nand U5603 (N_5603,N_663,N_2207);
and U5604 (N_5604,N_45,N_931);
or U5605 (N_5605,N_461,N_2598);
nor U5606 (N_5606,N_1139,N_558);
and U5607 (N_5607,N_665,N_2430);
or U5608 (N_5608,N_894,N_971);
nor U5609 (N_5609,N_1408,N_1855);
or U5610 (N_5610,N_1308,N_258);
and U5611 (N_5611,N_676,N_1180);
and U5612 (N_5612,N_2231,N_2209);
xnor U5613 (N_5613,N_405,N_1896);
nor U5614 (N_5614,N_2174,N_370);
nand U5615 (N_5615,N_1832,N_2125);
and U5616 (N_5616,N_284,N_577);
and U5617 (N_5617,N_2236,N_2065);
nand U5618 (N_5618,N_1946,N_2816);
nor U5619 (N_5619,N_2808,N_2305);
nor U5620 (N_5620,N_173,N_1223);
nand U5621 (N_5621,N_2153,N_1461);
nand U5622 (N_5622,N_1894,N_1744);
and U5623 (N_5623,N_1501,N_1984);
and U5624 (N_5624,N_387,N_2024);
or U5625 (N_5625,N_216,N_1886);
or U5626 (N_5626,N_938,N_2705);
nor U5627 (N_5627,N_2749,N_2878);
nor U5628 (N_5628,N_106,N_753);
and U5629 (N_5629,N_2586,N_33);
or U5630 (N_5630,N_396,N_906);
nor U5631 (N_5631,N_898,N_2517);
nor U5632 (N_5632,N_2600,N_1291);
xor U5633 (N_5633,N_950,N_2826);
or U5634 (N_5634,N_121,N_1782);
nand U5635 (N_5635,N_714,N_626);
and U5636 (N_5636,N_1182,N_2347);
nand U5637 (N_5637,N_1824,N_2471);
and U5638 (N_5638,N_2203,N_2689);
nand U5639 (N_5639,N_2073,N_2498);
xor U5640 (N_5640,N_2376,N_1270);
nor U5641 (N_5641,N_1625,N_1615);
and U5642 (N_5642,N_2645,N_1575);
nand U5643 (N_5643,N_2137,N_2208);
or U5644 (N_5644,N_1064,N_507);
nand U5645 (N_5645,N_60,N_2917);
nand U5646 (N_5646,N_2377,N_2605);
or U5647 (N_5647,N_2439,N_1378);
nor U5648 (N_5648,N_498,N_1169);
nand U5649 (N_5649,N_1342,N_1222);
or U5650 (N_5650,N_555,N_1152);
nor U5651 (N_5651,N_2654,N_2692);
nor U5652 (N_5652,N_2406,N_2687);
nand U5653 (N_5653,N_181,N_307);
and U5654 (N_5654,N_2314,N_2994);
and U5655 (N_5655,N_1463,N_1083);
and U5656 (N_5656,N_263,N_1972);
nor U5657 (N_5657,N_2166,N_717);
nor U5658 (N_5658,N_2913,N_441);
nor U5659 (N_5659,N_2657,N_1094);
nor U5660 (N_5660,N_736,N_2224);
or U5661 (N_5661,N_2318,N_693);
xor U5662 (N_5662,N_232,N_747);
xnor U5663 (N_5663,N_179,N_2583);
nor U5664 (N_5664,N_520,N_2595);
nor U5665 (N_5665,N_1826,N_206);
or U5666 (N_5666,N_1031,N_2497);
nand U5667 (N_5667,N_625,N_6);
and U5668 (N_5668,N_1182,N_186);
nor U5669 (N_5669,N_731,N_1496);
nor U5670 (N_5670,N_445,N_2351);
or U5671 (N_5671,N_1520,N_1312);
nand U5672 (N_5672,N_1127,N_2679);
nand U5673 (N_5673,N_2256,N_544);
nor U5674 (N_5674,N_1968,N_2721);
nand U5675 (N_5675,N_1076,N_2864);
nor U5676 (N_5676,N_526,N_275);
and U5677 (N_5677,N_148,N_760);
or U5678 (N_5678,N_2239,N_905);
or U5679 (N_5679,N_45,N_400);
or U5680 (N_5680,N_875,N_1989);
or U5681 (N_5681,N_2296,N_1982);
xnor U5682 (N_5682,N_479,N_2330);
or U5683 (N_5683,N_2339,N_992);
nor U5684 (N_5684,N_447,N_1476);
nor U5685 (N_5685,N_2886,N_899);
nand U5686 (N_5686,N_405,N_2115);
or U5687 (N_5687,N_2499,N_1336);
and U5688 (N_5688,N_630,N_186);
nor U5689 (N_5689,N_2694,N_684);
or U5690 (N_5690,N_1019,N_743);
or U5691 (N_5691,N_1202,N_2192);
and U5692 (N_5692,N_2407,N_2266);
nand U5693 (N_5693,N_925,N_177);
nand U5694 (N_5694,N_2142,N_2375);
or U5695 (N_5695,N_1780,N_304);
or U5696 (N_5696,N_1724,N_460);
or U5697 (N_5697,N_2028,N_765);
nor U5698 (N_5698,N_680,N_2907);
nor U5699 (N_5699,N_1662,N_10);
and U5700 (N_5700,N_2716,N_1512);
and U5701 (N_5701,N_370,N_1889);
xnor U5702 (N_5702,N_2785,N_882);
xor U5703 (N_5703,N_2362,N_1567);
and U5704 (N_5704,N_1691,N_1370);
xor U5705 (N_5705,N_1887,N_2478);
nand U5706 (N_5706,N_370,N_1906);
nand U5707 (N_5707,N_1607,N_273);
nand U5708 (N_5708,N_2992,N_2291);
nor U5709 (N_5709,N_130,N_1800);
and U5710 (N_5710,N_2211,N_2661);
and U5711 (N_5711,N_1813,N_2000);
xor U5712 (N_5712,N_1054,N_2260);
or U5713 (N_5713,N_426,N_8);
and U5714 (N_5714,N_2366,N_121);
or U5715 (N_5715,N_2307,N_215);
nand U5716 (N_5716,N_2570,N_1509);
nor U5717 (N_5717,N_201,N_1261);
and U5718 (N_5718,N_2616,N_1210);
nand U5719 (N_5719,N_2871,N_1776);
or U5720 (N_5720,N_1188,N_246);
nand U5721 (N_5721,N_1008,N_2806);
nor U5722 (N_5722,N_2481,N_396);
nand U5723 (N_5723,N_1099,N_1064);
nor U5724 (N_5724,N_1398,N_1482);
nor U5725 (N_5725,N_2723,N_2659);
and U5726 (N_5726,N_1640,N_1864);
nor U5727 (N_5727,N_1107,N_2291);
xor U5728 (N_5728,N_2348,N_537);
nand U5729 (N_5729,N_343,N_2680);
nor U5730 (N_5730,N_2608,N_888);
nor U5731 (N_5731,N_1199,N_1032);
nand U5732 (N_5732,N_2120,N_2242);
xor U5733 (N_5733,N_546,N_1651);
nand U5734 (N_5734,N_1237,N_54);
xnor U5735 (N_5735,N_2637,N_605);
nor U5736 (N_5736,N_467,N_766);
and U5737 (N_5737,N_2760,N_2045);
and U5738 (N_5738,N_376,N_1842);
nand U5739 (N_5739,N_2651,N_1325);
nor U5740 (N_5740,N_2120,N_743);
nand U5741 (N_5741,N_1485,N_1109);
nor U5742 (N_5742,N_962,N_1376);
or U5743 (N_5743,N_1560,N_146);
and U5744 (N_5744,N_907,N_2081);
nand U5745 (N_5745,N_984,N_2242);
or U5746 (N_5746,N_2111,N_1094);
xor U5747 (N_5747,N_2182,N_1887);
nand U5748 (N_5748,N_324,N_124);
nor U5749 (N_5749,N_2562,N_1339);
or U5750 (N_5750,N_300,N_1088);
nand U5751 (N_5751,N_619,N_2591);
and U5752 (N_5752,N_2646,N_1694);
xor U5753 (N_5753,N_1675,N_47);
or U5754 (N_5754,N_1853,N_1807);
xnor U5755 (N_5755,N_748,N_923);
nor U5756 (N_5756,N_2055,N_388);
xor U5757 (N_5757,N_1958,N_582);
nand U5758 (N_5758,N_2156,N_2428);
and U5759 (N_5759,N_2438,N_2919);
nor U5760 (N_5760,N_1147,N_2696);
and U5761 (N_5761,N_564,N_336);
nor U5762 (N_5762,N_1396,N_2356);
nand U5763 (N_5763,N_2742,N_601);
and U5764 (N_5764,N_1681,N_655);
and U5765 (N_5765,N_2444,N_870);
nor U5766 (N_5766,N_2471,N_913);
and U5767 (N_5767,N_1095,N_619);
nor U5768 (N_5768,N_1137,N_484);
nor U5769 (N_5769,N_683,N_2132);
and U5770 (N_5770,N_2138,N_1540);
or U5771 (N_5771,N_1434,N_1471);
and U5772 (N_5772,N_148,N_2943);
and U5773 (N_5773,N_629,N_1759);
nor U5774 (N_5774,N_1427,N_703);
or U5775 (N_5775,N_1510,N_1465);
nor U5776 (N_5776,N_2999,N_2204);
nand U5777 (N_5777,N_1933,N_911);
or U5778 (N_5778,N_2502,N_2374);
or U5779 (N_5779,N_1089,N_2927);
xor U5780 (N_5780,N_2638,N_1905);
nand U5781 (N_5781,N_2192,N_779);
xor U5782 (N_5782,N_2700,N_1501);
and U5783 (N_5783,N_474,N_2700);
and U5784 (N_5784,N_2595,N_2417);
xnor U5785 (N_5785,N_1993,N_2472);
nor U5786 (N_5786,N_172,N_2820);
nand U5787 (N_5787,N_2212,N_1899);
nand U5788 (N_5788,N_2287,N_1545);
and U5789 (N_5789,N_2062,N_2081);
nor U5790 (N_5790,N_1663,N_1057);
nor U5791 (N_5791,N_2644,N_1592);
nand U5792 (N_5792,N_4,N_1820);
nand U5793 (N_5793,N_731,N_2681);
and U5794 (N_5794,N_1070,N_1782);
and U5795 (N_5795,N_2336,N_693);
xnor U5796 (N_5796,N_2077,N_2466);
nand U5797 (N_5797,N_2679,N_2111);
nor U5798 (N_5798,N_676,N_977);
and U5799 (N_5799,N_1557,N_2853);
or U5800 (N_5800,N_437,N_556);
xor U5801 (N_5801,N_1932,N_182);
nor U5802 (N_5802,N_1845,N_1340);
nand U5803 (N_5803,N_2813,N_2142);
xor U5804 (N_5804,N_512,N_2256);
or U5805 (N_5805,N_1825,N_2646);
nand U5806 (N_5806,N_2909,N_1476);
or U5807 (N_5807,N_2480,N_1033);
or U5808 (N_5808,N_2358,N_861);
and U5809 (N_5809,N_1792,N_1707);
nand U5810 (N_5810,N_103,N_1705);
nand U5811 (N_5811,N_2972,N_1473);
or U5812 (N_5812,N_174,N_731);
or U5813 (N_5813,N_1632,N_1375);
and U5814 (N_5814,N_2593,N_390);
xor U5815 (N_5815,N_2323,N_155);
nand U5816 (N_5816,N_1137,N_2859);
nor U5817 (N_5817,N_684,N_2002);
nor U5818 (N_5818,N_2469,N_2903);
or U5819 (N_5819,N_2609,N_2513);
and U5820 (N_5820,N_632,N_1134);
or U5821 (N_5821,N_530,N_1134);
and U5822 (N_5822,N_231,N_2692);
nand U5823 (N_5823,N_176,N_1174);
xor U5824 (N_5824,N_2392,N_913);
and U5825 (N_5825,N_660,N_2733);
nand U5826 (N_5826,N_1677,N_2663);
or U5827 (N_5827,N_900,N_2045);
nor U5828 (N_5828,N_907,N_629);
nor U5829 (N_5829,N_1274,N_1442);
and U5830 (N_5830,N_2109,N_41);
nor U5831 (N_5831,N_715,N_2614);
nand U5832 (N_5832,N_855,N_1664);
nor U5833 (N_5833,N_2682,N_1546);
nand U5834 (N_5834,N_2278,N_778);
nand U5835 (N_5835,N_1193,N_2247);
or U5836 (N_5836,N_143,N_2338);
nor U5837 (N_5837,N_2483,N_2717);
nor U5838 (N_5838,N_984,N_1291);
nand U5839 (N_5839,N_1800,N_1696);
xor U5840 (N_5840,N_746,N_1514);
and U5841 (N_5841,N_2838,N_1845);
nand U5842 (N_5842,N_608,N_1416);
and U5843 (N_5843,N_648,N_413);
nor U5844 (N_5844,N_2516,N_1392);
or U5845 (N_5845,N_2466,N_2759);
or U5846 (N_5846,N_2253,N_1324);
or U5847 (N_5847,N_826,N_1579);
nand U5848 (N_5848,N_1534,N_467);
nand U5849 (N_5849,N_2374,N_908);
nand U5850 (N_5850,N_503,N_685);
or U5851 (N_5851,N_2392,N_2728);
or U5852 (N_5852,N_2880,N_2561);
nand U5853 (N_5853,N_1672,N_1006);
and U5854 (N_5854,N_2328,N_49);
and U5855 (N_5855,N_635,N_2014);
or U5856 (N_5856,N_1101,N_2323);
or U5857 (N_5857,N_1661,N_1597);
and U5858 (N_5858,N_2648,N_99);
nor U5859 (N_5859,N_2368,N_231);
and U5860 (N_5860,N_2236,N_765);
nand U5861 (N_5861,N_2476,N_2006);
nor U5862 (N_5862,N_1502,N_54);
or U5863 (N_5863,N_2634,N_259);
and U5864 (N_5864,N_553,N_1103);
nor U5865 (N_5865,N_567,N_2497);
nor U5866 (N_5866,N_2199,N_897);
nor U5867 (N_5867,N_1754,N_2555);
or U5868 (N_5868,N_216,N_577);
xnor U5869 (N_5869,N_1922,N_946);
or U5870 (N_5870,N_1653,N_830);
xor U5871 (N_5871,N_2103,N_2714);
nor U5872 (N_5872,N_2832,N_1929);
nand U5873 (N_5873,N_512,N_2283);
and U5874 (N_5874,N_237,N_1429);
nor U5875 (N_5875,N_2458,N_666);
nand U5876 (N_5876,N_524,N_2694);
xor U5877 (N_5877,N_386,N_243);
and U5878 (N_5878,N_677,N_255);
nor U5879 (N_5879,N_234,N_2805);
nand U5880 (N_5880,N_2251,N_1249);
nand U5881 (N_5881,N_1651,N_2033);
or U5882 (N_5882,N_1721,N_1237);
nor U5883 (N_5883,N_1893,N_2890);
or U5884 (N_5884,N_1943,N_2035);
or U5885 (N_5885,N_2853,N_1678);
or U5886 (N_5886,N_516,N_2439);
nor U5887 (N_5887,N_1607,N_2519);
and U5888 (N_5888,N_2949,N_606);
xor U5889 (N_5889,N_1435,N_292);
and U5890 (N_5890,N_2357,N_2074);
or U5891 (N_5891,N_855,N_489);
nand U5892 (N_5892,N_2646,N_2382);
nand U5893 (N_5893,N_2360,N_415);
nor U5894 (N_5894,N_805,N_2039);
nor U5895 (N_5895,N_1860,N_419);
nor U5896 (N_5896,N_959,N_869);
and U5897 (N_5897,N_2805,N_374);
nand U5898 (N_5898,N_2874,N_2928);
nand U5899 (N_5899,N_1397,N_1433);
nor U5900 (N_5900,N_1709,N_2376);
and U5901 (N_5901,N_1192,N_1696);
and U5902 (N_5902,N_1993,N_2652);
nor U5903 (N_5903,N_1424,N_593);
nand U5904 (N_5904,N_2912,N_740);
nor U5905 (N_5905,N_580,N_1629);
and U5906 (N_5906,N_1557,N_346);
nand U5907 (N_5907,N_2052,N_2576);
and U5908 (N_5908,N_241,N_2999);
and U5909 (N_5909,N_2620,N_725);
or U5910 (N_5910,N_1567,N_1928);
nand U5911 (N_5911,N_1052,N_554);
nor U5912 (N_5912,N_2321,N_2127);
nor U5913 (N_5913,N_602,N_1862);
nand U5914 (N_5914,N_877,N_1782);
nor U5915 (N_5915,N_1932,N_1955);
nand U5916 (N_5916,N_2821,N_944);
nor U5917 (N_5917,N_1226,N_987);
nand U5918 (N_5918,N_2609,N_1055);
nand U5919 (N_5919,N_509,N_1653);
and U5920 (N_5920,N_426,N_889);
nor U5921 (N_5921,N_2532,N_1120);
xnor U5922 (N_5922,N_2127,N_1815);
or U5923 (N_5923,N_2764,N_2428);
and U5924 (N_5924,N_721,N_127);
and U5925 (N_5925,N_511,N_1869);
or U5926 (N_5926,N_1514,N_1353);
nor U5927 (N_5927,N_511,N_1988);
or U5928 (N_5928,N_2801,N_2113);
nand U5929 (N_5929,N_1011,N_1263);
nor U5930 (N_5930,N_2469,N_393);
nand U5931 (N_5931,N_2749,N_816);
nor U5932 (N_5932,N_626,N_1709);
nand U5933 (N_5933,N_2998,N_2946);
nand U5934 (N_5934,N_2306,N_2366);
and U5935 (N_5935,N_35,N_1167);
nand U5936 (N_5936,N_867,N_1453);
xor U5937 (N_5937,N_1546,N_781);
nor U5938 (N_5938,N_693,N_2745);
or U5939 (N_5939,N_1935,N_2469);
or U5940 (N_5940,N_2856,N_1542);
nor U5941 (N_5941,N_2609,N_635);
and U5942 (N_5942,N_1570,N_605);
nor U5943 (N_5943,N_1781,N_2373);
or U5944 (N_5944,N_2501,N_1293);
nor U5945 (N_5945,N_696,N_568);
and U5946 (N_5946,N_2140,N_1460);
xor U5947 (N_5947,N_2492,N_1530);
nand U5948 (N_5948,N_1737,N_1541);
nor U5949 (N_5949,N_118,N_2171);
or U5950 (N_5950,N_2185,N_2060);
and U5951 (N_5951,N_2873,N_2233);
nand U5952 (N_5952,N_1099,N_746);
and U5953 (N_5953,N_2876,N_2338);
xnor U5954 (N_5954,N_2784,N_1398);
nor U5955 (N_5955,N_2827,N_2639);
or U5956 (N_5956,N_1181,N_2375);
nor U5957 (N_5957,N_2147,N_1664);
and U5958 (N_5958,N_613,N_267);
and U5959 (N_5959,N_1521,N_1787);
and U5960 (N_5960,N_2571,N_906);
nor U5961 (N_5961,N_303,N_2402);
xor U5962 (N_5962,N_1005,N_468);
or U5963 (N_5963,N_2711,N_780);
nor U5964 (N_5964,N_1365,N_1195);
nand U5965 (N_5965,N_2909,N_1620);
or U5966 (N_5966,N_2502,N_1400);
nand U5967 (N_5967,N_1422,N_2762);
or U5968 (N_5968,N_1383,N_1111);
nand U5969 (N_5969,N_1168,N_2812);
nor U5970 (N_5970,N_1131,N_1854);
and U5971 (N_5971,N_2119,N_2253);
xor U5972 (N_5972,N_1683,N_1887);
and U5973 (N_5973,N_2152,N_1355);
xor U5974 (N_5974,N_1364,N_2005);
nand U5975 (N_5975,N_2262,N_1309);
or U5976 (N_5976,N_2430,N_207);
nor U5977 (N_5977,N_750,N_1301);
nor U5978 (N_5978,N_1363,N_828);
xnor U5979 (N_5979,N_632,N_1949);
nor U5980 (N_5980,N_715,N_485);
nor U5981 (N_5981,N_190,N_119);
nor U5982 (N_5982,N_2670,N_1206);
nand U5983 (N_5983,N_2689,N_1058);
nor U5984 (N_5984,N_2022,N_1281);
and U5985 (N_5985,N_379,N_2373);
or U5986 (N_5986,N_1573,N_1709);
nor U5987 (N_5987,N_259,N_1974);
nor U5988 (N_5988,N_1666,N_108);
nor U5989 (N_5989,N_671,N_2087);
nor U5990 (N_5990,N_2206,N_289);
or U5991 (N_5991,N_28,N_2889);
and U5992 (N_5992,N_2662,N_418);
or U5993 (N_5993,N_2942,N_1915);
and U5994 (N_5994,N_1081,N_1549);
nor U5995 (N_5995,N_1933,N_2776);
nor U5996 (N_5996,N_681,N_656);
and U5997 (N_5997,N_1905,N_105);
or U5998 (N_5998,N_1521,N_2847);
or U5999 (N_5999,N_1838,N_2602);
and U6000 (N_6000,N_4421,N_5731);
nand U6001 (N_6001,N_5079,N_5535);
or U6002 (N_6002,N_4195,N_5235);
and U6003 (N_6003,N_5716,N_5825);
or U6004 (N_6004,N_4773,N_5915);
and U6005 (N_6005,N_3158,N_5369);
nor U6006 (N_6006,N_5984,N_4014);
xor U6007 (N_6007,N_5578,N_3670);
nand U6008 (N_6008,N_5151,N_5831);
and U6009 (N_6009,N_4279,N_4066);
nor U6010 (N_6010,N_4091,N_4904);
and U6011 (N_6011,N_3741,N_3606);
or U6012 (N_6012,N_3721,N_3645);
nand U6013 (N_6013,N_4393,N_5862);
nand U6014 (N_6014,N_3067,N_3246);
nor U6015 (N_6015,N_4707,N_3903);
and U6016 (N_6016,N_5962,N_5429);
nand U6017 (N_6017,N_4519,N_3001);
xnor U6018 (N_6018,N_5683,N_5750);
and U6019 (N_6019,N_3322,N_5426);
xor U6020 (N_6020,N_4876,N_4198);
xnor U6021 (N_6021,N_5153,N_3215);
nand U6022 (N_6022,N_4511,N_5131);
nor U6023 (N_6023,N_5680,N_3996);
or U6024 (N_6024,N_3119,N_4355);
and U6025 (N_6025,N_4555,N_4938);
xnor U6026 (N_6026,N_5207,N_5204);
and U6027 (N_6027,N_5262,N_3451);
or U6028 (N_6028,N_5619,N_3602);
and U6029 (N_6029,N_5743,N_3787);
nand U6030 (N_6030,N_4167,N_3271);
nand U6031 (N_6031,N_5434,N_5279);
or U6032 (N_6032,N_4108,N_3256);
or U6033 (N_6033,N_3648,N_5157);
nand U6034 (N_6034,N_5075,N_4064);
and U6035 (N_6035,N_3753,N_5183);
nor U6036 (N_6036,N_3751,N_5577);
nor U6037 (N_6037,N_3264,N_5382);
or U6038 (N_6038,N_4364,N_3534);
nor U6039 (N_6039,N_3675,N_4808);
nor U6040 (N_6040,N_5088,N_5686);
or U6041 (N_6041,N_3110,N_4281);
nand U6042 (N_6042,N_3413,N_4150);
nand U6043 (N_6043,N_5410,N_3330);
xor U6044 (N_6044,N_4331,N_3177);
xnor U6045 (N_6045,N_5900,N_3131);
nand U6046 (N_6046,N_4831,N_3209);
nand U6047 (N_6047,N_3354,N_5257);
and U6048 (N_6048,N_3399,N_5375);
and U6049 (N_6049,N_3937,N_4036);
xnor U6050 (N_6050,N_4851,N_3894);
nor U6051 (N_6051,N_4833,N_3196);
nor U6052 (N_6052,N_5753,N_5758);
and U6053 (N_6053,N_4688,N_3044);
and U6054 (N_6054,N_5352,N_3462);
and U6055 (N_6055,N_5569,N_4439);
and U6056 (N_6056,N_4772,N_4875);
or U6057 (N_6057,N_5013,N_5105);
nor U6058 (N_6058,N_5863,N_3369);
and U6059 (N_6059,N_5191,N_3156);
and U6060 (N_6060,N_3694,N_5781);
nor U6061 (N_6061,N_4411,N_3139);
or U6062 (N_6062,N_3512,N_5960);
and U6063 (N_6063,N_5361,N_5198);
xnor U6064 (N_6064,N_5790,N_5642);
nand U6065 (N_6065,N_4535,N_3896);
and U6066 (N_6066,N_3312,N_3036);
xnor U6067 (N_6067,N_5253,N_5584);
or U6068 (N_6068,N_4911,N_5208);
xnor U6069 (N_6069,N_5789,N_5154);
or U6070 (N_6070,N_4021,N_5745);
and U6071 (N_6071,N_4941,N_3338);
nand U6072 (N_6072,N_5993,N_3535);
and U6073 (N_6073,N_4897,N_3951);
xor U6074 (N_6074,N_4492,N_4129);
and U6075 (N_6075,N_5893,N_3207);
or U6076 (N_6076,N_3270,N_5195);
or U6077 (N_6077,N_5256,N_3785);
nor U6078 (N_6078,N_4209,N_4401);
xor U6079 (N_6079,N_5412,N_4780);
and U6080 (N_6080,N_4803,N_4319);
and U6081 (N_6081,N_3977,N_5231);
or U6082 (N_6082,N_3183,N_3251);
and U6083 (N_6083,N_5615,N_5327);
or U6084 (N_6084,N_4955,N_5189);
xnor U6085 (N_6085,N_4354,N_4922);
nor U6086 (N_6086,N_4667,N_5944);
or U6087 (N_6087,N_4450,N_4549);
or U6088 (N_6088,N_3565,N_3340);
xnor U6089 (N_6089,N_4696,N_4508);
or U6090 (N_6090,N_4154,N_4842);
nand U6091 (N_6091,N_4741,N_4750);
nand U6092 (N_6092,N_5925,N_3607);
nor U6093 (N_6093,N_4774,N_3892);
or U6094 (N_6094,N_3571,N_4845);
nand U6095 (N_6095,N_4087,N_5887);
nand U6096 (N_6096,N_5548,N_5769);
nand U6097 (N_6097,N_5518,N_3736);
nor U6098 (N_6098,N_3058,N_5665);
nand U6099 (N_6099,N_5715,N_5212);
nand U6100 (N_6100,N_4133,N_4823);
and U6101 (N_6101,N_4863,N_5138);
nor U6102 (N_6102,N_5744,N_4657);
nand U6103 (N_6103,N_5069,N_5842);
xor U6104 (N_6104,N_5200,N_3763);
nand U6105 (N_6105,N_5529,N_5346);
and U6106 (N_6106,N_5585,N_3883);
and U6107 (N_6107,N_5726,N_5551);
nand U6108 (N_6108,N_4380,N_4587);
nor U6109 (N_6109,N_3530,N_4998);
nor U6110 (N_6110,N_3150,N_3008);
nand U6111 (N_6111,N_3840,N_4383);
nand U6112 (N_6112,N_4692,N_4796);
nor U6113 (N_6113,N_3623,N_4344);
or U6114 (N_6114,N_4113,N_4822);
nor U6115 (N_6115,N_5123,N_3477);
or U6116 (N_6116,N_3831,N_3541);
nor U6117 (N_6117,N_5067,N_3885);
nor U6118 (N_6118,N_4274,N_4184);
or U6119 (N_6119,N_3710,N_3761);
nand U6120 (N_6120,N_5659,N_5975);
xnor U6121 (N_6121,N_4423,N_3418);
and U6122 (N_6122,N_4400,N_3819);
or U6123 (N_6123,N_3910,N_4948);
and U6124 (N_6124,N_3812,N_5306);
nor U6125 (N_6125,N_4871,N_4857);
nand U6126 (N_6126,N_3428,N_5017);
nand U6127 (N_6127,N_4560,N_3358);
nor U6128 (N_6128,N_3536,N_3460);
or U6129 (N_6129,N_5633,N_4665);
or U6130 (N_6130,N_5763,N_3279);
xor U6131 (N_6131,N_3070,N_3668);
and U6132 (N_6132,N_4708,N_5794);
xor U6133 (N_6133,N_3442,N_3574);
and U6134 (N_6134,N_3936,N_3441);
or U6135 (N_6135,N_5823,N_4470);
nand U6136 (N_6136,N_4789,N_3144);
nand U6137 (N_6137,N_5821,N_4105);
nand U6138 (N_6138,N_5439,N_5152);
nor U6139 (N_6139,N_5994,N_3682);
nor U6140 (N_6140,N_5421,N_4020);
nor U6141 (N_6141,N_4314,N_5610);
nand U6142 (N_6142,N_3076,N_4614);
nor U6143 (N_6143,N_4542,N_3174);
xnor U6144 (N_6144,N_4957,N_4077);
or U6145 (N_6145,N_4507,N_5675);
or U6146 (N_6146,N_3305,N_4194);
or U6147 (N_6147,N_4451,N_4047);
nor U6148 (N_6148,N_4709,N_3148);
nand U6149 (N_6149,N_3643,N_3778);
nand U6150 (N_6150,N_4583,N_5180);
nor U6151 (N_6151,N_5221,N_4616);
nor U6152 (N_6152,N_3096,N_4111);
nand U6153 (N_6153,N_5612,N_5621);
and U6154 (N_6154,N_4865,N_4747);
or U6155 (N_6155,N_5210,N_3514);
nor U6156 (N_6156,N_4680,N_4196);
and U6157 (N_6157,N_5567,N_4266);
xnor U6158 (N_6158,N_5654,N_4921);
xor U6159 (N_6159,N_5689,N_4001);
nor U6160 (N_6160,N_5700,N_5423);
and U6161 (N_6161,N_4043,N_3866);
and U6162 (N_6162,N_5016,N_3856);
xor U6163 (N_6163,N_4454,N_4443);
nor U6164 (N_6164,N_5852,N_4104);
nor U6165 (N_6165,N_4982,N_4365);
nand U6166 (N_6166,N_5135,N_4388);
nand U6167 (N_6167,N_5799,N_3781);
nand U6168 (N_6168,N_4147,N_3810);
and U6169 (N_6169,N_5630,N_4699);
nand U6170 (N_6170,N_4112,N_3968);
xnor U6171 (N_6171,N_3306,N_3527);
or U6172 (N_6172,N_3962,N_3265);
xor U6173 (N_6173,N_4270,N_5844);
nor U6174 (N_6174,N_4448,N_4757);
and U6175 (N_6175,N_5358,N_3170);
and U6176 (N_6176,N_4582,N_5566);
nand U6177 (N_6177,N_3956,N_3238);
nand U6178 (N_6178,N_3884,N_4821);
or U6179 (N_6179,N_5169,N_3543);
and U6180 (N_6180,N_5943,N_5812);
nor U6181 (N_6181,N_3045,N_3234);
and U6182 (N_6182,N_5658,N_3093);
nand U6183 (N_6183,N_5310,N_4034);
nand U6184 (N_6184,N_3876,N_5953);
or U6185 (N_6185,N_5575,N_4053);
and U6186 (N_6186,N_5809,N_5912);
nor U6187 (N_6187,N_5864,N_5225);
nand U6188 (N_6188,N_5004,N_4513);
nor U6189 (N_6189,N_5942,N_3415);
nand U6190 (N_6190,N_5990,N_5236);
nor U6191 (N_6191,N_5534,N_3194);
or U6192 (N_6192,N_4491,N_3783);
and U6193 (N_6193,N_5752,N_4217);
or U6194 (N_6194,N_4381,N_4810);
or U6195 (N_6195,N_3872,N_4601);
xor U6196 (N_6196,N_5587,N_4025);
or U6197 (N_6197,N_4418,N_4755);
and U6198 (N_6198,N_4520,N_3376);
nand U6199 (N_6199,N_5599,N_4533);
or U6200 (N_6200,N_4640,N_5111);
nand U6201 (N_6201,N_4452,N_4990);
nor U6202 (N_6202,N_4927,N_5401);
nor U6203 (N_6203,N_5285,N_4122);
xor U6204 (N_6204,N_5528,N_4946);
nor U6205 (N_6205,N_4449,N_5093);
or U6206 (N_6206,N_4063,N_5568);
nor U6207 (N_6207,N_5589,N_4242);
and U6208 (N_6208,N_4647,N_5552);
xor U6209 (N_6209,N_4799,N_3315);
xnor U6210 (N_6210,N_3718,N_5931);
or U6211 (N_6211,N_3311,N_5907);
nand U6212 (N_6212,N_4148,N_3284);
nor U6213 (N_6213,N_4838,N_4844);
or U6214 (N_6214,N_4888,N_5701);
xnor U6215 (N_6215,N_5638,N_4445);
or U6216 (N_6216,N_4989,N_5342);
or U6217 (N_6217,N_4033,N_5362);
nor U6218 (N_6218,N_5649,N_3104);
nor U6219 (N_6219,N_3538,N_5114);
xor U6220 (N_6220,N_3383,N_4310);
or U6221 (N_6221,N_5238,N_5655);
and U6222 (N_6222,N_5274,N_5388);
or U6223 (N_6223,N_3920,N_3957);
or U6224 (N_6224,N_3438,N_3537);
nor U6225 (N_6225,N_3362,N_5640);
and U6226 (N_6226,N_5590,N_3683);
or U6227 (N_6227,N_3554,N_4284);
nand U6228 (N_6228,N_3899,N_5699);
nor U6229 (N_6229,N_5291,N_5264);
or U6230 (N_6230,N_5333,N_4356);
and U6231 (N_6231,N_3134,N_4642);
or U6232 (N_6232,N_5930,N_4347);
and U6233 (N_6233,N_5168,N_5433);
xnor U6234 (N_6234,N_5515,N_4644);
nor U6235 (N_6235,N_4246,N_4556);
or U6236 (N_6236,N_4885,N_4362);
nor U6237 (N_6237,N_5720,N_4992);
nor U6238 (N_6238,N_3969,N_4480);
xnor U6239 (N_6239,N_4444,N_5541);
and U6240 (N_6240,N_5116,N_4545);
or U6241 (N_6241,N_4239,N_5300);
nor U6242 (N_6242,N_3000,N_3933);
nand U6243 (N_6243,N_3587,N_5422);
nand U6244 (N_6244,N_5160,N_5603);
xnor U6245 (N_6245,N_3600,N_3770);
and U6246 (N_6246,N_5586,N_3949);
nor U6247 (N_6247,N_5787,N_4585);
and U6248 (N_6248,N_5970,N_5187);
and U6249 (N_6249,N_4767,N_4031);
and U6250 (N_6250,N_3553,N_4602);
nor U6251 (N_6251,N_4711,N_3175);
or U6252 (N_6252,N_4051,N_4220);
nor U6253 (N_6253,N_3931,N_3808);
nor U6254 (N_6254,N_5450,N_5058);
or U6255 (N_6255,N_3344,N_4930);
nand U6256 (N_6256,N_4429,N_5365);
nand U6257 (N_6257,N_3649,N_3463);
and U6258 (N_6258,N_5676,N_4224);
or U6259 (N_6259,N_5695,N_3510);
nor U6260 (N_6260,N_5202,N_3408);
nor U6261 (N_6261,N_3749,N_3955);
or U6262 (N_6262,N_5739,N_5501);
or U6263 (N_6263,N_5836,N_5428);
nand U6264 (N_6264,N_3267,N_3755);
nor U6265 (N_6265,N_4233,N_5020);
and U6266 (N_6266,N_5512,N_3118);
nand U6267 (N_6267,N_3459,N_4517);
and U6268 (N_6268,N_3976,N_3739);
or U6269 (N_6269,N_5038,N_5560);
nor U6270 (N_6270,N_3456,N_4328);
nand U6271 (N_6271,N_4038,N_4461);
xor U6272 (N_6272,N_5628,N_4285);
nand U6273 (N_6273,N_5527,N_4742);
or U6274 (N_6274,N_5980,N_5413);
nand U6275 (N_6275,N_5951,N_5513);
xor U6276 (N_6276,N_3203,N_3720);
nand U6277 (N_6277,N_5060,N_5049);
and U6278 (N_6278,N_5351,N_3266);
nor U6279 (N_6279,N_3403,N_3125);
and U6280 (N_6280,N_5670,N_3392);
and U6281 (N_6281,N_5708,N_4849);
and U6282 (N_6282,N_4761,N_3359);
nand U6283 (N_6283,N_3690,N_3128);
nor U6284 (N_6284,N_3659,N_3786);
or U6285 (N_6285,N_3155,N_5461);
xor U6286 (N_6286,N_3027,N_5295);
nor U6287 (N_6287,N_5833,N_5521);
nand U6288 (N_6288,N_3240,N_5600);
and U6289 (N_6289,N_5923,N_5373);
nand U6290 (N_6290,N_3006,N_5440);
nor U6291 (N_6291,N_4880,N_3310);
and U6292 (N_6292,N_5272,N_5985);
nand U6293 (N_6293,N_4681,N_3318);
nand U6294 (N_6294,N_4980,N_4425);
and U6295 (N_6295,N_3384,N_4939);
nor U6296 (N_6296,N_5550,N_3123);
nor U6297 (N_6297,N_4191,N_3799);
nor U6298 (N_6298,N_3400,N_3803);
nand U6299 (N_6299,N_4295,N_4959);
or U6300 (N_6300,N_3804,N_3958);
nand U6301 (N_6301,N_3285,N_3059);
or U6302 (N_6302,N_4787,N_3135);
and U6303 (N_6303,N_4618,N_4275);
xnor U6304 (N_6304,N_3353,N_5023);
nand U6305 (N_6305,N_4288,N_4756);
nor U6306 (N_6306,N_3049,N_3842);
xnor U6307 (N_6307,N_5121,N_3272);
and U6308 (N_6308,N_4661,N_5041);
nor U6309 (N_6309,N_3081,N_3429);
or U6310 (N_6310,N_4685,N_3185);
or U6311 (N_6311,N_4032,N_3583);
and U6312 (N_6312,N_4435,N_4458);
or U6313 (N_6313,N_5330,N_5288);
nor U6314 (N_6314,N_3109,N_3747);
nor U6315 (N_6315,N_4256,N_5570);
or U6316 (N_6316,N_4754,N_5703);
nor U6317 (N_6317,N_5251,N_3924);
or U6318 (N_6318,N_4716,N_3236);
or U6319 (N_6319,N_3178,N_5094);
or U6320 (N_6320,N_4795,N_5956);
nor U6321 (N_6321,N_4794,N_4396);
nand U6322 (N_6322,N_3499,N_4684);
nor U6323 (N_6323,N_5692,N_5099);
nor U6324 (N_6324,N_5172,N_3666);
or U6325 (N_6325,N_3302,N_4753);
nand U6326 (N_6326,N_4408,N_4081);
and U6327 (N_6327,N_3615,N_4199);
nand U6328 (N_6328,N_3642,N_5040);
or U6329 (N_6329,N_3452,N_5162);
or U6330 (N_6330,N_4979,N_3352);
or U6331 (N_6331,N_3230,N_3074);
and U6332 (N_6332,N_5848,N_5827);
or U6333 (N_6333,N_3300,N_3542);
nor U6334 (N_6334,N_4790,N_3126);
and U6335 (N_6335,N_5091,N_4690);
and U6336 (N_6336,N_3502,N_3922);
or U6337 (N_6337,N_3889,N_4931);
nand U6338 (N_6338,N_4078,N_3206);
or U6339 (N_6339,N_4299,N_4075);
nor U6340 (N_6340,N_5878,N_4487);
or U6341 (N_6341,N_5635,N_5103);
or U6342 (N_6342,N_3231,N_3182);
and U6343 (N_6343,N_5991,N_5068);
nor U6344 (N_6344,N_3503,N_5335);
nor U6345 (N_6345,N_3569,N_4960);
or U6346 (N_6346,N_4007,N_5797);
or U6347 (N_6347,N_3425,N_4475);
xor U6348 (N_6348,N_3692,N_4076);
xor U6349 (N_6349,N_5089,N_3580);
or U6350 (N_6350,N_3304,N_5751);
and U6351 (N_6351,N_4371,N_3713);
xor U6352 (N_6352,N_3039,N_5139);
nor U6353 (N_6353,N_3745,N_3966);
nor U6354 (N_6354,N_3709,N_5334);
or U6355 (N_6355,N_5171,N_5052);
nand U6356 (N_6356,N_4100,N_4628);
nand U6357 (N_6357,N_3990,N_5656);
or U6358 (N_6358,N_4717,N_3090);
and U6359 (N_6359,N_3370,N_3319);
and U6360 (N_6360,N_3960,N_3348);
nor U6361 (N_6361,N_5919,N_4343);
or U6362 (N_6362,N_3491,N_5810);
and U6363 (N_6363,N_4569,N_3860);
and U6364 (N_6364,N_5939,N_5666);
nor U6365 (N_6365,N_3086,N_5479);
and U6366 (N_6366,N_4895,N_3414);
and U6367 (N_6367,N_5205,N_3867);
or U6368 (N_6368,N_5115,N_5519);
and U6369 (N_6369,N_4485,N_5841);
xor U6370 (N_6370,N_5469,N_4339);
nor U6371 (N_6371,N_3628,N_4889);
xor U6372 (N_6372,N_5090,N_5313);
and U6373 (N_6373,N_3505,N_4934);
nor U6374 (N_6374,N_3037,N_5400);
nor U6375 (N_6375,N_4045,N_4226);
or U6376 (N_6376,N_5704,N_5129);
nor U6377 (N_6377,N_4442,N_5062);
nor U6378 (N_6378,N_5486,N_5220);
nand U6379 (N_6379,N_3180,N_5158);
and U6380 (N_6380,N_5130,N_4677);
xnor U6381 (N_6381,N_5822,N_5065);
or U6382 (N_6382,N_5436,N_3779);
nor U6383 (N_6383,N_3072,N_4544);
or U6384 (N_6384,N_4019,N_4395);
or U6385 (N_6385,N_3711,N_5219);
and U6386 (N_6386,N_3129,N_3112);
nor U6387 (N_6387,N_5332,N_4860);
nand U6388 (N_6388,N_5861,N_4704);
nand U6389 (N_6389,N_4697,N_4558);
and U6390 (N_6390,N_4547,N_3561);
nand U6391 (N_6391,N_5616,N_4996);
nand U6392 (N_6392,N_3515,N_3575);
xnor U6393 (N_6393,N_3309,N_5782);
and U6394 (N_6394,N_4965,N_5714);
nor U6395 (N_6395,N_4382,N_4910);
and U6396 (N_6396,N_4650,N_3186);
or U6397 (N_6397,N_3811,N_4499);
nand U6398 (N_6398,N_4044,N_5609);
or U6399 (N_6399,N_4783,N_4596);
xnor U6400 (N_6400,N_4936,N_4092);
or U6401 (N_6401,N_5725,N_5855);
and U6402 (N_6402,N_4305,N_4080);
xor U6403 (N_6403,N_5488,N_4700);
nand U6404 (N_6404,N_3601,N_4651);
and U6405 (N_6405,N_4463,N_3255);
or U6406 (N_6406,N_3278,N_5230);
and U6407 (N_6407,N_4779,N_3146);
and U6408 (N_6408,N_5042,N_5574);
or U6409 (N_6409,N_5524,N_5340);
nand U6410 (N_6410,N_3220,N_3064);
or U6411 (N_6411,N_4332,N_4925);
and U6412 (N_6412,N_5523,N_5903);
nor U6413 (N_6413,N_4261,N_5559);
and U6414 (N_6414,N_5326,N_4966);
or U6415 (N_6415,N_5299,N_4137);
nand U6416 (N_6416,N_5698,N_4751);
nor U6417 (N_6417,N_5133,N_3620);
nor U6418 (N_6418,N_3568,N_3257);
or U6419 (N_6419,N_4609,N_4405);
or U6420 (N_6420,N_5211,N_5012);
or U6421 (N_6421,N_5881,N_4771);
or U6422 (N_6422,N_5218,N_5934);
nand U6423 (N_6423,N_3986,N_3545);
or U6424 (N_6424,N_4593,N_3547);
and U6425 (N_6425,N_5663,N_5000);
nand U6426 (N_6426,N_5868,N_4894);
or U6427 (N_6427,N_3411,N_3834);
nand U6428 (N_6428,N_3313,N_3038);
and U6429 (N_6429,N_4210,N_4723);
nor U6430 (N_6430,N_3546,N_5320);
nor U6431 (N_6431,N_4099,N_3153);
and U6432 (N_6432,N_3651,N_5322);
nor U6433 (N_6433,N_3172,N_3632);
nor U6434 (N_6434,N_5687,N_3106);
nor U6435 (N_6435,N_4595,N_4269);
nor U6436 (N_6436,N_5899,N_5920);
nor U6437 (N_6437,N_3397,N_3518);
and U6438 (N_6438,N_4538,N_5266);
and U6439 (N_6439,N_3520,N_5571);
or U6440 (N_6440,N_4621,N_4584);
and U6441 (N_6441,N_5186,N_5955);
and U6442 (N_6442,N_3323,N_5774);
and U6443 (N_6443,N_5935,N_5557);
nand U6444 (N_6444,N_3200,N_4202);
and U6445 (N_6445,N_3822,N_4384);
nand U6446 (N_6446,N_3317,N_3725);
or U6447 (N_6447,N_3939,N_4752);
nor U6448 (N_6448,N_5070,N_4390);
nor U6449 (N_6449,N_3169,N_5102);
nand U6450 (N_6450,N_3449,N_5420);
nand U6451 (N_6451,N_4298,N_3043);
and U6452 (N_6452,N_3681,N_5565);
xor U6453 (N_6453,N_5771,N_5481);
nand U6454 (N_6454,N_5003,N_5085);
nor U6455 (N_6455,N_3735,N_3496);
and U6456 (N_6456,N_5924,N_4923);
nor U6457 (N_6457,N_4433,N_4258);
or U6458 (N_6458,N_5979,N_5634);
nor U6459 (N_6459,N_5148,N_4176);
and U6460 (N_6460,N_4373,N_4306);
nand U6461 (N_6461,N_4659,N_3492);
and U6462 (N_6462,N_5772,N_5460);
and U6463 (N_6463,N_5496,N_5549);
or U6464 (N_6464,N_3355,N_3385);
nand U6465 (N_6465,N_3379,N_3347);
xor U6466 (N_6466,N_4468,N_4049);
nand U6467 (N_6467,N_3361,N_5729);
nor U6468 (N_6468,N_4829,N_5796);
nand U6469 (N_6469,N_3523,N_3095);
nor U6470 (N_6470,N_4834,N_5871);
nand U6471 (N_6471,N_5073,N_3879);
or U6472 (N_6472,N_4705,N_4776);
nor U6473 (N_6473,N_3752,N_3833);
nand U6474 (N_6474,N_5021,N_3188);
nand U6475 (N_6475,N_3759,N_4662);
nor U6476 (N_6476,N_3141,N_5228);
nor U6477 (N_6477,N_5530,N_3780);
xor U6478 (N_6478,N_5393,N_4046);
nand U6479 (N_6479,N_3914,N_4760);
and U6480 (N_6480,N_5046,N_5507);
or U6481 (N_6481,N_4243,N_3494);
and U6482 (N_6482,N_5254,N_4899);
xnor U6483 (N_6483,N_5522,N_4271);
or U6484 (N_6484,N_5631,N_4830);
nor U6485 (N_6485,N_4866,N_4872);
nor U6486 (N_6486,N_3837,N_3862);
and U6487 (N_6487,N_4416,N_5755);
or U6488 (N_6488,N_5011,N_5646);
and U6489 (N_6489,N_4869,N_4277);
and U6490 (N_6490,N_4733,N_3042);
and U6491 (N_6491,N_4290,N_3401);
or U6492 (N_6492,N_3020,N_3478);
and U6493 (N_6493,N_3389,N_4160);
and U6494 (N_6494,N_5805,N_5487);
xor U6495 (N_6495,N_4543,N_4465);
and U6496 (N_6496,N_5092,N_5775);
or U6497 (N_6497,N_3647,N_5667);
nor U6498 (N_6498,N_3771,N_5353);
xnor U6499 (N_6499,N_4935,N_4223);
nand U6500 (N_6500,N_4739,N_5384);
nand U6501 (N_6501,N_5717,N_5226);
and U6502 (N_6502,N_4252,N_4971);
nand U6503 (N_6503,N_4179,N_4495);
nand U6504 (N_6504,N_5679,N_4522);
nand U6505 (N_6505,N_5525,N_4027);
nand U6506 (N_6506,N_5328,N_5884);
nor U6507 (N_6507,N_3465,N_3467);
and U6508 (N_6508,N_3426,N_4068);
nand U6509 (N_6509,N_5312,N_3616);
nand U6510 (N_6510,N_4722,N_4800);
nand U6511 (N_6511,N_3160,N_3197);
nor U6512 (N_6512,N_5307,N_3498);
nor U6513 (N_6513,N_3419,N_3117);
nor U6514 (N_6514,N_3063,N_3548);
nor U6515 (N_6515,N_5444,N_4853);
or U6516 (N_6516,N_4879,N_3513);
and U6517 (N_6517,N_5302,N_3367);
or U6518 (N_6518,N_3424,N_3393);
nand U6519 (N_6519,N_3644,N_4337);
and U6520 (N_6520,N_4612,N_4694);
and U6521 (N_6521,N_4023,N_3013);
nand U6522 (N_6522,N_3850,N_4348);
and U6523 (N_6523,N_4906,N_4793);
and U6524 (N_6524,N_4567,N_5947);
or U6525 (N_6525,N_5712,N_5403);
or U6526 (N_6526,N_3820,N_5456);
or U6527 (N_6527,N_4929,N_5203);
or U6528 (N_6528,N_3791,N_5876);
and U6529 (N_6529,N_4379,N_4412);
nor U6530 (N_6530,N_5999,N_3524);
and U6531 (N_6531,N_3490,N_5966);
xnor U6532 (N_6532,N_3242,N_3472);
and U6533 (N_6533,N_4847,N_3599);
or U6534 (N_6534,N_5298,N_3078);
xor U6535 (N_6535,N_5269,N_3965);
nor U6536 (N_6536,N_5136,N_4660);
nand U6537 (N_6537,N_3660,N_4607);
xor U6538 (N_6538,N_4837,N_5192);
or U6539 (N_6539,N_5245,N_3740);
or U6540 (N_6540,N_4691,N_5008);
nand U6541 (N_6541,N_5684,N_3349);
and U6542 (N_6542,N_3210,N_3890);
or U6543 (N_6543,N_3888,N_3704);
nand U6544 (N_6544,N_3455,N_5759);
or U6545 (N_6545,N_3091,N_3439);
and U6546 (N_6546,N_4152,N_3489);
or U6547 (N_6547,N_3314,N_3796);
and U6548 (N_6548,N_5475,N_5387);
or U6549 (N_6549,N_4652,N_5493);
and U6550 (N_6550,N_5516,N_3714);
nor U6551 (N_6551,N_4572,N_3363);
or U6552 (N_6552,N_3423,N_3844);
or U6553 (N_6553,N_5902,N_5636);
or U6554 (N_6554,N_5643,N_4814);
or U6555 (N_6555,N_5503,N_5854);
nand U6556 (N_6556,N_4874,N_4798);
nand U6557 (N_6557,N_3453,N_3102);
and U6558 (N_6558,N_3923,N_3625);
nand U6559 (N_6559,N_3722,N_4422);
nor U6560 (N_6560,N_3915,N_5284);
nand U6561 (N_6561,N_5579,N_3409);
and U6562 (N_6562,N_3556,N_3161);
or U6563 (N_6563,N_3640,N_5286);
nand U6564 (N_6564,N_5142,N_4625);
or U6565 (N_6565,N_5555,N_3654);
and U6566 (N_6566,N_4532,N_4988);
and U6567 (N_6567,N_4670,N_3023);
nand U6568 (N_6568,N_4471,N_4048);
nor U6569 (N_6569,N_5370,N_4734);
nand U6570 (N_6570,N_3328,N_4069);
nand U6571 (N_6571,N_4985,N_4211);
nor U6572 (N_6572,N_3343,N_4819);
or U6573 (N_6573,N_4006,N_4215);
nand U6574 (N_6574,N_5308,N_3964);
or U6575 (N_6575,N_4240,N_3298);
nor U6576 (N_6576,N_3522,N_3018);
nand U6577 (N_6577,N_4856,N_4225);
and U6578 (N_6578,N_5414,N_4370);
and U6579 (N_6579,N_3636,N_3961);
and U6580 (N_6580,N_3578,N_5867);
or U6581 (N_6581,N_3676,N_5159);
or U6582 (N_6582,N_3826,N_5664);
nand U6583 (N_6583,N_5668,N_5161);
nand U6584 (N_6584,N_3192,N_3130);
nand U6585 (N_6585,N_4037,N_3813);
and U6586 (N_6586,N_4424,N_5438);
xor U6587 (N_6587,N_4843,N_3559);
nand U6588 (N_6588,N_4570,N_5497);
or U6589 (N_6589,N_3165,N_4663);
nor U6590 (N_6590,N_4197,N_3708);
xnor U6591 (N_6591,N_4234,N_4172);
and U6592 (N_6592,N_3880,N_5397);
nor U6593 (N_6593,N_3788,N_3396);
nor U6594 (N_6594,N_5341,N_3727);
nor U6595 (N_6595,N_4132,N_5596);
nor U6596 (N_6596,N_4208,N_3854);
and U6597 (N_6597,N_3470,N_4920);
nor U6598 (N_6598,N_5449,N_5399);
and U6599 (N_6599,N_5998,N_5178);
nand U6600 (N_6600,N_4168,N_5959);
and U6601 (N_6601,N_4958,N_4327);
and U6602 (N_6602,N_4004,N_5510);
and U6603 (N_6603,N_4824,N_3592);
nor U6604 (N_6604,N_3329,N_3646);
nor U6605 (N_6605,N_3723,N_5141);
and U6606 (N_6606,N_5873,N_5672);
xor U6607 (N_6607,N_5466,N_5780);
or U6608 (N_6608,N_5281,N_3525);
nand U6609 (N_6609,N_4598,N_5478);
nor U6610 (N_6610,N_3212,N_5050);
nand U6611 (N_6611,N_4013,N_3851);
nor U6612 (N_6612,N_4141,N_4322);
nand U6613 (N_6613,N_4334,N_5834);
nor U6614 (N_6614,N_5427,N_3627);
nand U6615 (N_6615,N_4525,N_3865);
or U6616 (N_6616,N_3237,N_3950);
nor U6617 (N_6617,N_5372,N_5856);
nor U6618 (N_6618,N_4453,N_5880);
and U6619 (N_6619,N_3417,N_4204);
and U6620 (N_6620,N_5674,N_3388);
nand U6621 (N_6621,N_4781,N_3360);
nand U6622 (N_6622,N_3115,N_5732);
xor U6623 (N_6623,N_4566,N_3677);
and U6624 (N_6624,N_4493,N_3098);
xnor U6625 (N_6625,N_3695,N_3277);
or U6626 (N_6626,N_4892,N_5882);
and U6627 (N_6627,N_4698,N_4514);
nand U6628 (N_6628,N_4591,N_3189);
nor U6629 (N_6629,N_3159,N_3299);
nor U6630 (N_6630,N_3814,N_3219);
or U6631 (N_6631,N_5366,N_3797);
nor U6632 (N_6632,N_3917,N_5125);
nor U6633 (N_6633,N_3325,N_4812);
nand U6634 (N_6634,N_3701,N_3191);
and U6635 (N_6635,N_4441,N_5730);
xnor U6636 (N_6636,N_5895,N_5858);
nor U6637 (N_6637,N_5542,N_5336);
nand U6638 (N_6638,N_5467,N_4516);
or U6639 (N_6639,N_4093,N_3963);
or U6640 (N_6640,N_5074,N_3737);
and U6641 (N_6641,N_4840,N_4170);
or U6642 (N_6642,N_3784,N_5252);
and U6643 (N_6643,N_3420,N_5325);
or U6644 (N_6644,N_4675,N_4251);
and U6645 (N_6645,N_3433,N_5007);
nand U6646 (N_6646,N_5035,N_3943);
or U6647 (N_6647,N_4318,N_4010);
nand U6648 (N_6648,N_3500,N_5319);
nand U6649 (N_6649,N_3195,N_3801);
nand U6650 (N_6650,N_4802,N_3843);
or U6651 (N_6651,N_4727,N_3870);
and U6652 (N_6652,N_5371,N_3274);
and U6653 (N_6653,N_5140,N_3440);
xor U6654 (N_6654,N_4120,N_4633);
or U6655 (N_6655,N_3887,N_5015);
xor U6656 (N_6656,N_4744,N_3790);
or U6657 (N_6657,N_3754,N_5323);
or U6658 (N_6658,N_4738,N_3595);
or U6659 (N_6659,N_3335,N_4586);
or U6660 (N_6660,N_5149,N_4655);
nor U6661 (N_6661,N_4653,N_3140);
or U6662 (N_6662,N_4478,N_4627);
nand U6663 (N_6663,N_4055,N_4143);
and U6664 (N_6664,N_4476,N_5014);
and U6665 (N_6665,N_5435,N_5588);
and U6666 (N_6666,N_5830,N_4227);
nor U6667 (N_6667,N_4987,N_3995);
or U6668 (N_6668,N_3002,N_5533);
nand U6669 (N_6669,N_3893,N_3443);
or U6670 (N_6670,N_3877,N_3263);
xor U6671 (N_6671,N_5010,N_4551);
nor U6672 (N_6672,N_5837,N_5807);
nand U6673 (N_6673,N_4398,N_5737);
nor U6674 (N_6674,N_3137,N_4562);
and U6675 (N_6675,N_4826,N_4402);
nand U6676 (N_6676,N_4721,N_3596);
nor U6677 (N_6677,N_4417,N_5064);
and U6678 (N_6678,N_5045,N_3913);
nor U6679 (N_6679,N_5558,N_3124);
or U6680 (N_6680,N_3816,N_5408);
or U6681 (N_6681,N_4610,N_3674);
and U6682 (N_6682,N_3244,N_4028);
or U6683 (N_6683,N_3407,N_3113);
and U6684 (N_6684,N_4428,N_4731);
nor U6685 (N_6685,N_4883,N_4228);
or U6686 (N_6686,N_3984,N_4573);
or U6687 (N_6687,N_4632,N_3897);
or U6688 (N_6688,N_3444,N_4732);
xnor U6689 (N_6689,N_5937,N_5591);
or U6690 (N_6690,N_3466,N_4740);
or U6691 (N_6691,N_5232,N_3693);
nand U6692 (N_6692,N_3730,N_4526);
nand U6693 (N_6693,N_5911,N_4703);
nand U6694 (N_6694,N_3859,N_3217);
nor U6695 (N_6695,N_3945,N_5502);
or U6696 (N_6696,N_3154,N_5303);
or U6697 (N_6697,N_5389,N_5735);
and U6698 (N_6698,N_4873,N_4592);
or U6699 (N_6699,N_5455,N_4296);
nand U6700 (N_6700,N_4165,N_5671);
or U6701 (N_6701,N_5209,N_5276);
and U6702 (N_6702,N_3431,N_4222);
nand U6703 (N_6703,N_3052,N_3566);
and U6704 (N_6704,N_5520,N_4138);
and U6705 (N_6705,N_4260,N_4315);
nor U6706 (N_6706,N_5678,N_3848);
and U6707 (N_6707,N_4512,N_5727);
and U6708 (N_6708,N_5097,N_4308);
and U6709 (N_6709,N_5314,N_5402);
nor U6710 (N_6710,N_5562,N_4190);
xor U6711 (N_6711,N_5241,N_5468);
nor U6712 (N_6712,N_5972,N_5532);
or U6713 (N_6713,N_4410,N_5237);
nor U6714 (N_6714,N_5623,N_3386);
and U6715 (N_6715,N_4745,N_3151);
nor U6716 (N_6716,N_4859,N_4608);
or U6717 (N_6717,N_3276,N_3307);
nand U6718 (N_6718,N_5697,N_3517);
nor U6719 (N_6719,N_3341,N_3650);
and U6720 (N_6720,N_4301,N_4877);
xnor U6721 (N_6721,N_3871,N_5653);
and U6722 (N_6722,N_5889,N_5294);
nor U6723 (N_6723,N_3378,N_3450);
nor U6724 (N_6724,N_4884,N_4324);
nor U6725 (N_6725,N_3832,N_3003);
nand U6726 (N_6726,N_4392,N_3511);
xor U6727 (N_6727,N_3336,N_5819);
nand U6728 (N_6728,N_4648,N_5928);
nor U6729 (N_6729,N_4140,N_4323);
or U6730 (N_6730,N_4095,N_3247);
nor U6731 (N_6731,N_3201,N_5411);
nor U6732 (N_6732,N_4940,N_4918);
nor U6733 (N_6733,N_3689,N_3181);
or U6734 (N_6734,N_5660,N_5517);
nor U6735 (N_6735,N_5229,N_5150);
or U6736 (N_6736,N_3351,N_5201);
nand U6737 (N_6737,N_3746,N_3868);
or U6738 (N_6738,N_5233,N_4580);
or U6739 (N_6739,N_5766,N_3841);
or U6740 (N_6740,N_4903,N_5113);
and U6741 (N_6741,N_5117,N_5086);
or U6742 (N_6742,N_5938,N_3613);
and U6743 (N_6743,N_3672,N_5964);
and U6744 (N_6744,N_4397,N_5898);
nand U6745 (N_6745,N_4436,N_5078);
nand U6746 (N_6746,N_3168,N_4878);
or U6747 (N_6747,N_4022,N_4126);
nor U6748 (N_6748,N_5215,N_3457);
nand U6749 (N_6749,N_4109,N_3157);
xnor U6750 (N_6750,N_4366,N_5904);
xor U6751 (N_6751,N_3662,N_3198);
or U6752 (N_6752,N_5354,N_4999);
or U6753 (N_6753,N_5134,N_3679);
or U6754 (N_6754,N_4553,N_4486);
and U6755 (N_6755,N_5922,N_5002);
nor U6756 (N_6756,N_5707,N_5802);
nor U6757 (N_6757,N_3296,N_5315);
nor U6758 (N_6758,N_4164,N_4438);
xnor U6759 (N_6759,N_4351,N_5626);
or U6760 (N_6760,N_3585,N_5849);
or U6761 (N_6761,N_4446,N_5709);
nand U6762 (N_6762,N_5865,N_4775);
xnor U6763 (N_6763,N_4638,N_4978);
nand U6764 (N_6764,N_3025,N_3065);
or U6765 (N_6765,N_3111,N_4311);
nand U6766 (N_6766,N_4368,N_4702);
nand U6767 (N_6767,N_4919,N_3717);
nor U6768 (N_6768,N_3301,N_4689);
or U6769 (N_6769,N_5681,N_5213);
and U6770 (N_6770,N_3757,N_5693);
xnor U6771 (N_6771,N_3975,N_4206);
and U6772 (N_6772,N_3685,N_5283);
nor U6773 (N_6773,N_3482,N_5506);
xnor U6774 (N_6774,N_3608,N_4498);
nor U6775 (N_6775,N_4611,N_4415);
nand U6776 (N_6776,N_4954,N_5850);
nor U6777 (N_6777,N_4419,N_3835);
or U6778 (N_6778,N_3942,N_4145);
nand U6779 (N_6779,N_5728,N_4947);
or U6780 (N_6780,N_4706,N_3908);
nand U6781 (N_6781,N_5118,N_3731);
nand U6782 (N_6782,N_4714,N_3041);
or U6783 (N_6783,N_5583,N_3823);
and U6784 (N_6784,N_5997,N_4933);
and U6785 (N_6785,N_3069,N_4637);
nor U6786 (N_6786,N_4763,N_3807);
nor U6787 (N_6787,N_3886,N_3919);
nand U6788 (N_6788,N_5196,N_5767);
xnor U6789 (N_6789,N_5946,N_4074);
nor U6790 (N_6790,N_3611,N_4497);
or U6791 (N_6791,N_5127,N_4159);
nor U6792 (N_6792,N_5967,N_3089);
and U6793 (N_6793,N_4993,N_5705);
and U6794 (N_6794,N_3707,N_3184);
or U6795 (N_6795,N_5582,N_3769);
nand U6796 (N_6796,N_3010,N_3895);
nor U6797 (N_6797,N_4528,N_3598);
nand U6798 (N_6798,N_5537,N_5446);
nor U6799 (N_6799,N_3434,N_5360);
nor U6800 (N_6800,N_3447,N_5181);
or U6801 (N_6801,N_4765,N_4777);
nor U6802 (N_6802,N_4534,N_4597);
nor U6803 (N_6803,N_5890,N_4391);
and U6804 (N_6804,N_3907,N_3094);
and U6805 (N_6805,N_3768,N_3404);
nand U6806 (N_6806,N_3639,N_4061);
nand U6807 (N_6807,N_4067,N_5611);
xor U6808 (N_6808,N_3824,N_3214);
xor U6809 (N_6809,N_4770,N_4071);
nand U6810 (N_6810,N_3009,N_4086);
nand U6811 (N_6811,N_5594,N_3445);
and U6812 (N_6812,N_5572,N_3874);
nor U6813 (N_6813,N_3412,N_4406);
or U6814 (N_6814,N_5248,N_3029);
nor U6815 (N_6815,N_3941,N_3526);
nand U6816 (N_6816,N_4282,N_5083);
nor U6817 (N_6817,N_4378,N_3241);
or U6818 (N_6818,N_3235,N_5164);
nand U6819 (N_6819,N_3992,N_3994);
nand U6820 (N_6820,N_3483,N_4976);
nand U6821 (N_6821,N_4374,N_4679);
or U6822 (N_6822,N_3243,N_3825);
or U6823 (N_6823,N_3617,N_3474);
or U6824 (N_6824,N_5419,N_5265);
or U6825 (N_6825,N_3748,N_4970);
nand U6826 (N_6826,N_4852,N_5495);
or U6827 (N_6827,N_3519,N_3532);
nor U6828 (N_6828,N_3577,N_5872);
nand U6829 (N_6829,N_5144,N_5561);
and U6830 (N_6830,N_4668,N_4500);
and U6831 (N_6831,N_4127,N_5777);
xor U6832 (N_6832,N_3934,N_4041);
nand U6833 (N_6833,N_5483,N_5908);
nand U6834 (N_6834,N_3802,N_4130);
nand U6835 (N_6835,N_3334,N_5543);
nor U6836 (N_6836,N_4477,N_3087);
and U6837 (N_6837,N_5992,N_3926);
and U6838 (N_6838,N_4178,N_4088);
and U6839 (N_6839,N_3921,N_5345);
nand U6840 (N_6840,N_4403,N_4649);
nor U6841 (N_6841,N_4294,N_4730);
nor U6842 (N_6842,N_5747,N_3954);
nor U6843 (N_6843,N_5651,N_5926);
or U6844 (N_6844,N_3540,N_3603);
nor U6845 (N_6845,N_3798,N_3782);
and U6846 (N_6846,N_4193,N_3742);
nor U6847 (N_6847,N_4726,N_5888);
nand U6848 (N_6848,N_3667,N_3688);
and U6849 (N_6849,N_4581,N_3202);
nand U6850 (N_6850,N_5124,N_3593);
and U6851 (N_6851,N_3391,N_3700);
or U6852 (N_6852,N_5691,N_4292);
nor U6853 (N_6853,N_5170,N_3326);
nand U6854 (N_6854,N_5001,N_3371);
nor U6855 (N_6855,N_4836,N_4188);
or U6856 (N_6856,N_5806,N_5784);
or U6857 (N_6857,N_5958,N_4357);
or U6858 (N_6858,N_5453,N_4345);
nor U6859 (N_6859,N_4909,N_5417);
and U6860 (N_6860,N_4907,N_4340);
or U6861 (N_6861,N_3073,N_5106);
nor U6862 (N_6862,N_5184,N_5290);
nor U6863 (N_6863,N_4604,N_5374);
and U6864 (N_6864,N_5648,N_3528);
and U6865 (N_6865,N_5677,N_4639);
nand U6866 (N_6866,N_5282,N_4363);
or U6867 (N_6867,N_3581,N_4375);
or U6868 (N_6868,N_4230,N_5597);
xor U6869 (N_6869,N_3162,N_3061);
or U6870 (N_6870,N_3981,N_3508);
and U6871 (N_6871,N_3637,N_4886);
and U6872 (N_6872,N_3552,N_5760);
nand U6873 (N_6873,N_3504,N_4868);
or U6874 (N_6874,N_4297,N_5722);
nor U6875 (N_6875,N_4291,N_4720);
or U6876 (N_6876,N_3432,N_5305);
or U6877 (N_6877,N_4017,N_4481);
or U6878 (N_6878,N_4317,N_3262);
nor U6879 (N_6879,N_4005,N_5592);
nand U6880 (N_6880,N_4114,N_4782);
and U6881 (N_6881,N_4286,N_5071);
xor U6882 (N_6882,N_5563,N_3108);
nor U6883 (N_6883,N_5096,N_5740);
nand U6884 (N_6884,N_4420,N_3132);
or U6885 (N_6885,N_3127,N_4510);
nand U6886 (N_6886,N_3204,N_5109);
xnor U6887 (N_6887,N_5971,N_3597);
or U6888 (N_6888,N_5885,N_3022);
nor U6889 (N_6889,N_4967,N_3028);
and U6890 (N_6890,N_3988,N_3288);
or U6891 (N_6891,N_4302,N_5564);
nand U6892 (N_6892,N_3609,N_4235);
or U6893 (N_6893,N_5785,N_4056);
or U6894 (N_6894,N_4029,N_3589);
nor U6895 (N_6895,N_4372,N_3350);
or U6896 (N_6896,N_3827,N_5188);
nand U6897 (N_6897,N_5982,N_4748);
nand U6898 (N_6898,N_4012,N_3208);
nand U6899 (N_6899,N_5126,N_5662);
nand U6900 (N_6900,N_5801,N_3989);
nor U6901 (N_6901,N_4484,N_5632);
or U6902 (N_6902,N_4828,N_5019);
nor U6903 (N_6903,N_3932,N_4000);
or U6904 (N_6904,N_5199,N_4683);
nor U6905 (N_6905,N_5593,N_3004);
nand U6906 (N_6906,N_5905,N_3959);
and U6907 (N_6907,N_4600,N_5122);
and U6908 (N_6908,N_4713,N_5531);
nand U6909 (N_6909,N_3991,N_5107);
or U6910 (N_6910,N_5137,N_4115);
nor U6911 (N_6911,N_5573,N_3529);
and U6912 (N_6912,N_4352,N_4386);
or U6913 (N_6913,N_5968,N_4052);
nand U6914 (N_6914,N_4561,N_4588);
nand U6915 (N_6915,N_4882,N_3776);
and U6916 (N_6916,N_3289,N_5608);
nand U6917 (N_6917,N_5463,N_5875);
and U6918 (N_6918,N_3297,N_3405);
xnor U6919 (N_6919,N_5482,N_3821);
nor U6920 (N_6920,N_4937,N_5736);
and U6921 (N_6921,N_4577,N_4377);
nor U6922 (N_6922,N_3364,N_5702);
and U6923 (N_6923,N_4039,N_5380);
nand U6924 (N_6924,N_3026,N_4961);
nand U6925 (N_6925,N_3767,N_5377);
nand U6926 (N_6926,N_3594,N_4631);
nor U6927 (N_6927,N_5768,N_4241);
nand U6928 (N_6928,N_3143,N_3454);
nor U6929 (N_6929,N_4455,N_3333);
nand U6930 (N_6930,N_5176,N_4131);
nand U6931 (N_6931,N_4335,N_3935);
xnor U6932 (N_6932,N_5504,N_5620);
or U6933 (N_6933,N_5462,N_3972);
or U6934 (N_6934,N_4811,N_4501);
or U6935 (N_6935,N_5791,N_3805);
nand U6936 (N_6936,N_5870,N_4474);
nand U6937 (N_6937,N_5053,N_5447);
nor U6938 (N_6938,N_3147,N_4862);
and U6939 (N_6939,N_4189,N_4634);
nand U6940 (N_6940,N_3365,N_4342);
or U6941 (N_6941,N_4496,N_5406);
nor U6942 (N_6942,N_5009,N_5816);
xnor U6943 (N_6943,N_5289,N_3268);
nand U6944 (N_6944,N_5499,N_4962);
or U6945 (N_6945,N_5818,N_5261);
nand U6946 (N_6946,N_3332,N_4059);
nor U6947 (N_6947,N_5381,N_4244);
nand U6948 (N_6948,N_3292,N_4142);
or U6949 (N_6949,N_5741,N_5246);
and U6950 (N_6950,N_3092,N_5076);
and U6951 (N_6951,N_4914,N_5206);
or U6952 (N_6952,N_3927,N_5324);
and U6953 (N_6953,N_4192,N_3836);
nor U6954 (N_6954,N_4207,N_3099);
or U6955 (N_6955,N_3743,N_4457);
and U6956 (N_6956,N_5179,N_3227);
or U6957 (N_6957,N_4564,N_4462);
or U6958 (N_6958,N_3394,N_3254);
and U6959 (N_6959,N_3421,N_3327);
nand U6960 (N_6960,N_5800,N_3303);
nand U6961 (N_6961,N_4482,N_4908);
nand U6962 (N_6962,N_3715,N_5969);
xnor U6963 (N_6963,N_3211,N_4529);
nor U6964 (N_6964,N_5190,N_5746);
and U6965 (N_6965,N_4518,N_5647);
nor U6966 (N_6966,N_5669,N_5343);
and U6967 (N_6967,N_3560,N_3398);
or U6968 (N_6968,N_4695,N_3697);
nor U6969 (N_6969,N_3473,N_5913);
nand U6970 (N_6970,N_5359,N_5948);
xnor U6971 (N_6971,N_5275,N_4011);
and U6972 (N_6972,N_3978,N_4255);
or U6973 (N_6973,N_4434,N_4623);
nor U6974 (N_6974,N_5817,N_5072);
nor U6975 (N_6975,N_4620,N_3461);
nor U6976 (N_6976,N_4530,N_3071);
and U6977 (N_6977,N_3891,N_5983);
xnor U6978 (N_6978,N_4003,N_5263);
nor U6979 (N_6979,N_3853,N_3947);
or U6980 (N_6980,N_4121,N_4554);
nor U6981 (N_6981,N_3658,N_5084);
or U6982 (N_6982,N_5311,N_5432);
nor U6983 (N_6983,N_4149,N_5028);
nor U6984 (N_6984,N_5508,N_3509);
and U6985 (N_6985,N_4430,N_4009);
nor U6986 (N_6986,N_5721,N_4503);
nor U6987 (N_6987,N_3339,N_5954);
and U6988 (N_6988,N_3634,N_3881);
nand U6989 (N_6989,N_3900,N_3705);
or U6990 (N_6990,N_5082,N_3716);
nor U6991 (N_6991,N_4839,N_4816);
and U6992 (N_6992,N_5044,N_4759);
nand U6993 (N_6993,N_3521,N_4162);
and U6994 (N_6994,N_5430,N_4912);
or U6995 (N_6995,N_4218,N_5338);
nand U6996 (N_6996,N_5018,N_3911);
and U6997 (N_6997,N_3765,N_4447);
nand U6998 (N_6998,N_5546,N_5143);
and U6999 (N_6999,N_3261,N_3699);
and U7000 (N_7000,N_5025,N_5595);
and U7001 (N_7001,N_5063,N_4278);
nor U7002 (N_7002,N_3680,N_4236);
nand U7003 (N_7003,N_5820,N_3377);
and U7004 (N_7004,N_3678,N_3993);
nand U7005 (N_7005,N_5613,N_5554);
nor U7006 (N_7006,N_3732,N_5216);
and U7007 (N_7007,N_3107,N_4788);
nor U7008 (N_7008,N_5258,N_3764);
and U7009 (N_7009,N_4984,N_4473);
nor U7010 (N_7010,N_3544,N_4293);
nand U7011 (N_7011,N_3983,N_3218);
or U7012 (N_7012,N_4096,N_5491);
nor U7013 (N_7013,N_5398,N_3728);
xor U7014 (N_7014,N_5357,N_5077);
or U7015 (N_7015,N_5363,N_5936);
nor U7016 (N_7016,N_3729,N_4065);
or U7017 (N_7017,N_5792,N_5811);
nand U7018 (N_7018,N_4409,N_5859);
nand U7019 (N_7019,N_4949,N_5165);
nor U7020 (N_7020,N_5576,N_4187);
and U7021 (N_7021,N_4945,N_3564);
nor U7022 (N_7022,N_4089,N_4136);
or U7023 (N_7023,N_4369,N_4603);
nor U7024 (N_7024,N_5688,N_3373);
nand U7025 (N_7025,N_4983,N_5770);
nand U7026 (N_7026,N_3055,N_5645);
and U7027 (N_7027,N_5742,N_4635);
and U7028 (N_7028,N_4718,N_5748);
xor U7029 (N_7029,N_4200,N_3024);
nor U7030 (N_7030,N_3982,N_4394);
nor U7031 (N_7031,N_3539,N_4158);
nand U7032 (N_7032,N_5485,N_3283);
nor U7033 (N_7033,N_5604,N_5713);
and U7034 (N_7034,N_4917,N_3083);
nand U7035 (N_7035,N_5471,N_5316);
nand U7036 (N_7036,N_3815,N_3612);
nand U7037 (N_7037,N_5255,N_5470);
and U7038 (N_7038,N_5452,N_5734);
and U7039 (N_7039,N_5598,N_4968);
nand U7040 (N_7040,N_4504,N_4432);
nand U7041 (N_7041,N_5840,N_4900);
xnor U7042 (N_7042,N_5301,N_5033);
nand U7043 (N_7043,N_4991,N_4186);
xnor U7044 (N_7044,N_4719,N_5425);
xor U7045 (N_7045,N_4119,N_3050);
xnor U7046 (N_7046,N_5738,N_4098);
and U7047 (N_7047,N_4835,N_5580);
nand U7048 (N_7048,N_3435,N_5509);
nor U7049 (N_7049,N_5988,N_4488);
or U7050 (N_7050,N_4134,N_3395);
and U7051 (N_7051,N_4951,N_4008);
nor U7052 (N_7052,N_5424,N_4466);
xor U7053 (N_7053,N_5916,N_5147);
or U7054 (N_7054,N_4213,N_3838);
nand U7055 (N_7055,N_4248,N_3686);
xnor U7056 (N_7056,N_3342,N_4994);
and U7057 (N_7057,N_4768,N_5476);
nor U7058 (N_7058,N_3079,N_5242);
xnor U7059 (N_7059,N_3480,N_3635);
or U7060 (N_7060,N_4571,N_4002);
and U7061 (N_7061,N_4483,N_4276);
or U7062 (N_7062,N_3898,N_4563);
and U7063 (N_7063,N_4272,N_5024);
or U7064 (N_7064,N_5786,N_3275);
and U7065 (N_7065,N_3034,N_3567);
or U7066 (N_7066,N_3484,N_5390);
or U7067 (N_7067,N_4360,N_5244);
or U7068 (N_7068,N_3048,N_5145);
nor U7069 (N_7069,N_4809,N_5404);
nand U7070 (N_7070,N_5963,N_3173);
nor U7071 (N_7071,N_5448,N_3167);
nor U7072 (N_7072,N_4701,N_5177);
nand U7073 (N_7073,N_4326,N_5193);
nand U7074 (N_7074,N_4943,N_4950);
nor U7075 (N_7075,N_4460,N_4166);
and U7076 (N_7076,N_3878,N_4778);
nand U7077 (N_7077,N_3239,N_4891);
nor U7078 (N_7078,N_5477,N_3719);
nor U7079 (N_7079,N_4832,N_3282);
xor U7080 (N_7080,N_4615,N_3011);
and U7081 (N_7081,N_4540,N_5981);
nor U7082 (N_7082,N_3793,N_4890);
or U7083 (N_7083,N_4437,N_4431);
or U7084 (N_7084,N_4472,N_3846);
or U7085 (N_7085,N_3869,N_5719);
nand U7086 (N_7086,N_4805,N_4212);
and U7087 (N_7087,N_4590,N_3260);
xor U7088 (N_7088,N_4273,N_4669);
nor U7089 (N_7089,N_5081,N_3629);
xor U7090 (N_7090,N_4307,N_4686);
nand U7091 (N_7091,N_5318,N_4085);
nand U7092 (N_7092,N_3249,N_3223);
and U7093 (N_7093,N_4729,N_5940);
or U7094 (N_7094,N_4107,N_3570);
nand U7095 (N_7095,N_4887,N_5442);
and U7096 (N_7096,N_4630,N_5851);
or U7097 (N_7097,N_5329,N_5376);
nor U7098 (N_7098,N_5650,N_3806);
and U7099 (N_7099,N_4232,N_5795);
or U7100 (N_7100,N_5347,N_3967);
and U7101 (N_7101,N_3436,N_4710);
or U7102 (N_7102,N_5724,N_3345);
xor U7103 (N_7103,N_3248,N_5182);
nand U7104 (N_7104,N_4280,N_4901);
or U7105 (N_7105,N_4505,N_4682);
or U7106 (N_7106,N_3775,N_4079);
and U7107 (N_7107,N_4385,N_3487);
and U7108 (N_7108,N_5368,N_5860);
or U7109 (N_7109,N_4575,N_5098);
nand U7110 (N_7110,N_4523,N_5829);
and U7111 (N_7111,N_4786,N_4018);
and U7112 (N_7112,N_4253,N_3979);
nand U7113 (N_7113,N_5101,N_3655);
xor U7114 (N_7114,N_3281,N_4489);
or U7115 (N_7115,N_5492,N_3882);
xnor U7116 (N_7116,N_5039,N_5268);
and U7117 (N_7117,N_5778,N_5764);
nor U7118 (N_7118,N_5484,N_3114);
nand U7119 (N_7119,N_3233,N_5441);
nand U7120 (N_7120,N_5762,N_4867);
or U7121 (N_7121,N_4762,N_3551);
or U7122 (N_7122,N_3622,N_4333);
nand U7123 (N_7123,N_5048,N_3331);
xor U7124 (N_7124,N_5174,N_5155);
and U7125 (N_7125,N_4956,N_5652);
or U7126 (N_7126,N_5624,N_5280);
nand U7127 (N_7127,N_4953,N_4040);
and U7128 (N_7128,N_4942,N_5694);
and U7129 (N_7129,N_4804,N_3633);
or U7130 (N_7130,N_3380,N_4321);
and U7131 (N_7131,N_3875,N_4387);
and U7132 (N_7132,N_3269,N_5418);
nor U7133 (N_7133,N_3533,N_4054);
xor U7134 (N_7134,N_4182,N_4101);
nor U7135 (N_7135,N_3164,N_5826);
and U7136 (N_7136,N_4341,N_3944);
or U7137 (N_7137,N_5877,N_4303);
and U7138 (N_7138,N_5941,N_3563);
and U7139 (N_7139,N_5892,N_4042);
nor U7140 (N_7140,N_3402,N_5445);
nor U7141 (N_7141,N_5317,N_5054);
nor U7142 (N_7142,N_3138,N_3555);
and U7143 (N_7143,N_5490,N_3863);
and U7144 (N_7144,N_4404,N_4515);
nand U7145 (N_7145,N_5431,N_4359);
nor U7146 (N_7146,N_5505,N_5682);
nor U7147 (N_7147,N_3382,N_5897);
nor U7148 (N_7148,N_4024,N_5776);
and U7149 (N_7149,N_3550,N_4574);
nor U7150 (N_7150,N_3080,N_4764);
and U7151 (N_7151,N_3584,N_3948);
nor U7152 (N_7152,N_3253,N_4151);
and U7153 (N_7153,N_3015,N_5443);
and U7154 (N_7154,N_4464,N_4674);
nor U7155 (N_7155,N_5914,N_4728);
or U7156 (N_7156,N_3618,N_5185);
nand U7157 (N_7157,N_4309,N_3501);
and U7158 (N_7158,N_5271,N_3706);
and U7159 (N_7159,N_5553,N_3356);
nand U7160 (N_7160,N_4506,N_5874);
and U7161 (N_7161,N_3060,N_3422);
xnor U7162 (N_7162,N_5607,N_4981);
and U7163 (N_7163,N_3016,N_5614);
nand U7164 (N_7164,N_5929,N_4818);
xnor U7165 (N_7165,N_5270,N_5034);
and U7166 (N_7166,N_4712,N_3928);
or U7167 (N_7167,N_4541,N_4552);
and U7168 (N_7168,N_4841,N_5095);
and U7169 (N_7169,N_4817,N_5733);
nand U7170 (N_7170,N_5511,N_5026);
or U7171 (N_7171,N_5250,N_5349);
and U7172 (N_7172,N_5921,N_4090);
and U7173 (N_7173,N_3562,N_5030);
or U7174 (N_7174,N_3845,N_3005);
or U7175 (N_7175,N_4349,N_4216);
nor U7176 (N_7176,N_5556,N_3222);
nor U7177 (N_7177,N_3985,N_5227);
nand U7178 (N_7178,N_3847,N_3669);
and U7179 (N_7179,N_5120,N_5367);
nand U7180 (N_7180,N_4806,N_4440);
nor U7181 (N_7181,N_3469,N_4678);
and U7182 (N_7182,N_4097,N_3855);
or U7183 (N_7183,N_4524,N_4015);
nor U7184 (N_7184,N_4264,N_5950);
nand U7185 (N_7185,N_4263,N_4548);
xnor U7186 (N_7186,N_5214,N_5685);
or U7187 (N_7187,N_5027,N_5673);
or U7188 (N_7188,N_3531,N_3999);
nor U7189 (N_7189,N_4724,N_5909);
nor U7190 (N_7190,N_4094,N_5267);
nor U7191 (N_7191,N_3485,N_5278);
nor U7192 (N_7192,N_3630,N_3103);
and U7193 (N_7193,N_4265,N_4219);
and U7194 (N_7194,N_3828,N_3032);
nand U7195 (N_7195,N_4250,N_3488);
nand U7196 (N_7196,N_3224,N_3987);
and U7197 (N_7197,N_3105,N_5055);
nor U7198 (N_7198,N_5808,N_3294);
nand U7199 (N_7199,N_5392,N_3290);
nor U7200 (N_7200,N_4916,N_3232);
nor U7201 (N_7201,N_4825,N_3084);
or U7202 (N_7202,N_4676,N_3652);
nand U7203 (N_7203,N_3591,N_3750);
and U7204 (N_7204,N_4565,N_5379);
nand U7205 (N_7205,N_3321,N_4735);
and U7206 (N_7206,N_5788,N_4102);
or U7207 (N_7207,N_5886,N_3789);
and U7208 (N_7208,N_4469,N_4082);
and U7209 (N_7209,N_5407,N_4221);
or U7210 (N_7210,N_3101,N_3738);
nand U7211 (N_7211,N_5395,N_5629);
or U7212 (N_7212,N_5239,N_3726);
or U7213 (N_7213,N_3166,N_5696);
nand U7214 (N_7214,N_5581,N_4201);
nand U7215 (N_7215,N_3163,N_3698);
nand U7216 (N_7216,N_5974,N_3406);
nand U7217 (N_7217,N_4769,N_3187);
nand U7218 (N_7218,N_5364,N_4654);
and U7219 (N_7219,N_3293,N_4427);
xor U7220 (N_7220,N_5156,N_5348);
and U7221 (N_7221,N_3925,N_4687);
nand U7222 (N_7222,N_5080,N_4924);
or U7223 (N_7223,N_5217,N_5545);
and U7224 (N_7224,N_5057,N_5602);
and U7225 (N_7225,N_4546,N_5765);
nand U7226 (N_7226,N_3486,N_3145);
nand U7227 (N_7227,N_4858,N_3610);
nand U7228 (N_7228,N_4268,N_5249);
or U7229 (N_7229,N_4870,N_4174);
or U7230 (N_7230,N_3054,N_4559);
or U7231 (N_7231,N_4125,N_3762);
xor U7232 (N_7232,N_3387,N_3506);
and U7233 (N_7233,N_5296,N_5835);
xnor U7234 (N_7234,N_3702,N_4629);
and U7235 (N_7235,N_5458,N_5277);
xnor U7236 (N_7236,N_4646,N_3605);
and U7237 (N_7237,N_5957,N_4320);
nand U7238 (N_7238,N_5813,N_3573);
nor U7239 (N_7239,N_4864,N_3368);
nand U7240 (N_7240,N_4898,N_5273);
or U7241 (N_7241,N_4743,N_5706);
nor U7242 (N_7242,N_3448,N_5059);
nor U7243 (N_7243,N_3631,N_3273);
nor U7244 (N_7244,N_4617,N_3930);
nand U7245 (N_7245,N_5749,N_3663);
and U7246 (N_7246,N_4973,N_4664);
nor U7247 (N_7247,N_3077,N_5416);
nand U7248 (N_7248,N_3997,N_3205);
nor U7249 (N_7249,N_3033,N_4502);
nand U7250 (N_7250,N_4287,N_4807);
nor U7251 (N_7251,N_3974,N_3904);
xor U7252 (N_7252,N_5223,N_4791);
nand U7253 (N_7253,N_3122,N_4035);
or U7254 (N_7254,N_4237,N_4952);
nor U7255 (N_7255,N_3641,N_3286);
and U7256 (N_7256,N_5066,N_5866);
nor U7257 (N_7257,N_5606,N_3653);
nor U7258 (N_7258,N_4173,N_5292);
or U7259 (N_7259,N_4944,N_3495);
and U7260 (N_7260,N_3572,N_4766);
nor U7261 (N_7261,N_5949,N_5846);
nand U7262 (N_7262,N_4490,N_3626);
nor U7263 (N_7263,N_3929,N_4399);
xor U7264 (N_7264,N_4124,N_3691);
or U7265 (N_7265,N_4969,N_5457);
nor U7266 (N_7266,N_5339,N_3437);
nor U7267 (N_7267,N_3458,N_3116);
or U7268 (N_7268,N_4827,N_5773);
xnor U7269 (N_7269,N_5036,N_4589);
nor U7270 (N_7270,N_5932,N_4117);
and U7271 (N_7271,N_5378,N_5321);
or U7272 (N_7272,N_3259,N_4645);
or U7273 (N_7273,N_5197,N_5022);
or U7274 (N_7274,N_4414,N_3468);
nand U7275 (N_7275,N_4568,N_3684);
and U7276 (N_7276,N_3671,N_3068);
nor U7277 (N_7277,N_3410,N_3252);
nand U7278 (N_7278,N_5657,N_4407);
or U7279 (N_7279,N_3056,N_5756);
nor U7280 (N_7280,N_5536,N_4725);
nor U7281 (N_7281,N_4058,N_4358);
nand U7282 (N_7282,N_5853,N_3946);
xor U7283 (N_7283,N_4030,N_5779);
or U7284 (N_7284,N_3507,N_3287);
nor U7285 (N_7285,N_4426,N_4926);
or U7286 (N_7286,N_4606,N_5832);
nor U7287 (N_7287,N_4622,N_3381);
and U7288 (N_7288,N_3858,N_3760);
xor U7289 (N_7289,N_4350,N_3849);
nor U7290 (N_7290,N_5961,N_3035);
or U7291 (N_7291,N_5639,N_4641);
nor U7292 (N_7292,N_3320,N_3250);
nor U7293 (N_7293,N_5644,N_3030);
nor U7294 (N_7294,N_5711,N_5128);
nor U7295 (N_7295,N_3952,N_3229);
nor U7296 (N_7296,N_3864,N_4792);
and U7297 (N_7297,N_3337,N_3638);
nand U7298 (N_7298,N_3021,N_5224);
or U7299 (N_7299,N_4995,N_5037);
nand U7300 (N_7300,N_3171,N_5006);
and U7301 (N_7301,N_3416,N_5526);
xnor U7302 (N_7302,N_3586,N_5287);
and U7303 (N_7303,N_5798,N_5690);
nand U7304 (N_7304,N_4758,N_3758);
nor U7305 (N_7305,N_3346,N_4413);
or U7306 (N_7306,N_3938,N_3774);
or U7307 (N_7307,N_5894,N_5309);
nor U7308 (N_7308,N_4247,N_3100);
or U7309 (N_7309,N_5843,N_4183);
nand U7310 (N_7310,N_5394,N_4902);
and U7311 (N_7311,N_4932,N_3430);
nor U7312 (N_7312,N_3621,N_4084);
xor U7313 (N_7313,N_5538,N_5500);
nor U7314 (N_7314,N_4855,N_4073);
nor U7315 (N_7315,N_5815,N_5454);
and U7316 (N_7316,N_3047,N_3062);
and U7317 (N_7317,N_3558,N_5987);
xnor U7318 (N_7318,N_4245,N_4177);
nand U7319 (N_7319,N_5622,N_5173);
nand U7320 (N_7320,N_4116,N_5047);
and U7321 (N_7321,N_4336,N_3007);
or U7322 (N_7322,N_5051,N_4329);
nand U7323 (N_7323,N_4997,N_4974);
nor U7324 (N_7324,N_4157,N_5627);
xor U7325 (N_7325,N_3590,N_3839);
nor U7326 (N_7326,N_5661,N_5415);
nand U7327 (N_7327,N_4785,N_4169);
or U7328 (N_7328,N_4161,N_4626);
nand U7329 (N_7329,N_3557,N_4057);
and U7330 (N_7330,N_4531,N_5260);
nand U7331 (N_7331,N_4977,N_3142);
xor U7332 (N_7332,N_4016,N_3673);
or U7333 (N_7333,N_3818,N_3724);
nor U7334 (N_7334,N_4820,N_3665);
xnor U7335 (N_7335,N_3901,N_3136);
and U7336 (N_7336,N_5494,N_4599);
nor U7337 (N_7337,N_3479,N_4026);
nand U7338 (N_7338,N_3051,N_3549);
and U7339 (N_7339,N_5803,N_3912);
or U7340 (N_7340,N_5108,N_5618);
and U7341 (N_7341,N_3225,N_3973);
and U7342 (N_7342,N_4346,N_5757);
and U7343 (N_7343,N_3228,N_3664);
or U7344 (N_7344,N_4736,N_4249);
and U7345 (N_7345,N_4797,N_5383);
nand U7346 (N_7346,N_4467,N_4180);
nand U7347 (N_7347,N_4050,N_3481);
and U7348 (N_7348,N_3687,N_4153);
and U7349 (N_7349,N_4815,N_4367);
or U7350 (N_7350,N_3357,N_4312);
or U7351 (N_7351,N_5385,N_5297);
nand U7352 (N_7352,N_5355,N_4636);
or U7353 (N_7353,N_5883,N_5847);
nand U7354 (N_7354,N_3857,N_3213);
or U7355 (N_7355,N_5489,N_4861);
nor U7356 (N_7356,N_3588,N_3817);
or U7357 (N_7357,N_5906,N_4605);
and U7358 (N_7358,N_3088,N_4171);
and U7359 (N_7359,N_4156,N_5901);
and U7360 (N_7360,N_4509,N_4915);
or U7361 (N_7361,N_3661,N_4123);
or U7362 (N_7362,N_3097,N_4613);
or U7363 (N_7363,N_5087,N_5978);
or U7364 (N_7364,N_5031,N_4175);
nand U7365 (N_7365,N_3971,N_3031);
or U7366 (N_7366,N_3053,N_3497);
or U7367 (N_7367,N_4316,N_3795);
or U7368 (N_7368,N_5350,N_4619);
and U7369 (N_7369,N_4539,N_3657);
nor U7370 (N_7370,N_5965,N_3372);
or U7371 (N_7371,N_3916,N_4913);
or U7372 (N_7372,N_3582,N_4550);
and U7373 (N_7373,N_4693,N_5814);
or U7374 (N_7374,N_4110,N_4163);
xor U7375 (N_7375,N_4673,N_4185);
and U7376 (N_7376,N_3366,N_5464);
nand U7377 (N_7377,N_5304,N_5167);
xor U7378 (N_7378,N_5132,N_3493);
nor U7379 (N_7379,N_4850,N_3258);
nand U7380 (N_7380,N_4624,N_3324);
and U7381 (N_7381,N_4205,N_3085);
nand U7382 (N_7382,N_5247,N_5029);
and U7383 (N_7383,N_3918,N_5472);
nand U7384 (N_7384,N_4072,N_4578);
and U7385 (N_7385,N_3280,N_5391);
or U7386 (N_7386,N_3019,N_3012);
nand U7387 (N_7387,N_4231,N_5601);
nand U7388 (N_7388,N_4330,N_5437);
and U7389 (N_7389,N_3014,N_5498);
xnor U7390 (N_7390,N_3179,N_5344);
or U7391 (N_7391,N_5839,N_4746);
and U7392 (N_7392,N_5879,N_5945);
or U7393 (N_7393,N_3464,N_4737);
or U7394 (N_7394,N_5857,N_3295);
nor U7395 (N_7395,N_4229,N_4267);
nor U7396 (N_7396,N_5617,N_4118);
and U7397 (N_7397,N_5032,N_4893);
and U7398 (N_7398,N_3082,N_5869);
and U7399 (N_7399,N_5163,N_4643);
xnor U7400 (N_7400,N_5761,N_5514);
and U7401 (N_7401,N_5175,N_4594);
xor U7402 (N_7402,N_4283,N_5973);
nand U7403 (N_7403,N_5259,N_5918);
and U7404 (N_7404,N_5641,N_4128);
and U7405 (N_7405,N_5465,N_3905);
or U7406 (N_7406,N_5104,N_3199);
nor U7407 (N_7407,N_3476,N_5112);
and U7408 (N_7408,N_3792,N_5166);
nand U7409 (N_7409,N_4576,N_3057);
and U7410 (N_7410,N_4181,N_4238);
nand U7411 (N_7411,N_3176,N_3970);
or U7412 (N_7412,N_5710,N_5293);
or U7413 (N_7413,N_4521,N_5989);
and U7414 (N_7414,N_3902,N_3316);
and U7415 (N_7415,N_3744,N_5331);
and U7416 (N_7416,N_4848,N_5933);
nor U7417 (N_7417,N_3777,N_3516);
and U7418 (N_7418,N_5977,N_3475);
nand U7419 (N_7419,N_5480,N_4289);
nor U7420 (N_7420,N_3696,N_3809);
nand U7421 (N_7421,N_3873,N_3756);
nand U7422 (N_7422,N_5386,N_4203);
and U7423 (N_7423,N_3940,N_3149);
or U7424 (N_7424,N_3830,N_5995);
or U7425 (N_7425,N_4801,N_3576);
and U7426 (N_7426,N_5845,N_4070);
nand U7427 (N_7427,N_3614,N_5605);
nand U7428 (N_7428,N_3772,N_3712);
xor U7429 (N_7429,N_5540,N_5976);
nor U7430 (N_7430,N_5222,N_4060);
and U7431 (N_7431,N_4671,N_4214);
nand U7432 (N_7432,N_4666,N_3471);
nor U7433 (N_7433,N_5896,N_5240);
xor U7434 (N_7434,N_3909,N_3190);
nor U7435 (N_7435,N_3800,N_4656);
xnor U7436 (N_7436,N_5056,N_4749);
or U7437 (N_7437,N_4139,N_4376);
and U7438 (N_7438,N_3773,N_3245);
nand U7439 (N_7439,N_3733,N_5547);
or U7440 (N_7440,N_4083,N_4304);
and U7441 (N_7441,N_3075,N_3794);
nand U7442 (N_7442,N_3216,N_4155);
nor U7443 (N_7443,N_5891,N_4103);
or U7444 (N_7444,N_3291,N_3703);
nor U7445 (N_7445,N_3906,N_3766);
and U7446 (N_7446,N_5996,N_5194);
nor U7447 (N_7447,N_4456,N_5718);
and U7448 (N_7448,N_3375,N_4972);
and U7449 (N_7449,N_5451,N_4963);
and U7450 (N_7450,N_5723,N_4257);
nor U7451 (N_7451,N_3390,N_5473);
nand U7452 (N_7452,N_4557,N_5927);
nor U7453 (N_7453,N_4536,N_5828);
nor U7454 (N_7454,N_5119,N_5804);
nor U7455 (N_7455,N_4715,N_5952);
or U7456 (N_7456,N_5409,N_3734);
or U7457 (N_7457,N_4986,N_5824);
or U7458 (N_7458,N_5100,N_5910);
or U7459 (N_7459,N_4146,N_4905);
or U7460 (N_7460,N_5459,N_4254);
nor U7461 (N_7461,N_5917,N_5146);
nand U7462 (N_7462,N_4672,N_3152);
nand U7463 (N_7463,N_3604,N_5405);
nand U7464 (N_7464,N_5544,N_4062);
nand U7465 (N_7465,N_5234,N_4313);
or U7466 (N_7466,N_3046,N_3308);
nor U7467 (N_7467,N_3829,N_4579);
nand U7468 (N_7468,N_3374,N_5110);
nor U7469 (N_7469,N_3040,N_4854);
nand U7470 (N_7470,N_3998,N_5005);
nand U7471 (N_7471,N_4658,N_4389);
nor U7472 (N_7472,N_4881,N_5783);
or U7473 (N_7473,N_3120,N_3221);
or U7474 (N_7474,N_4896,N_5474);
or U7475 (N_7475,N_3427,N_3980);
xnor U7476 (N_7476,N_4144,N_3656);
and U7477 (N_7477,N_5356,N_3226);
xor U7478 (N_7478,N_3133,N_4537);
and U7479 (N_7479,N_5043,N_3066);
and U7480 (N_7480,N_3121,N_3579);
nand U7481 (N_7481,N_4494,N_5793);
and U7482 (N_7482,N_5986,N_4135);
or U7483 (N_7483,N_3619,N_5243);
or U7484 (N_7484,N_4479,N_3017);
nor U7485 (N_7485,N_4964,N_4813);
nor U7486 (N_7486,N_5337,N_4338);
and U7487 (N_7487,N_4975,N_4259);
nand U7488 (N_7488,N_3193,N_5838);
and U7489 (N_7489,N_4784,N_4846);
or U7490 (N_7490,N_4361,N_3953);
nand U7491 (N_7491,N_4459,N_4300);
and U7492 (N_7492,N_4325,N_5637);
and U7493 (N_7493,N_4353,N_3624);
nor U7494 (N_7494,N_5061,N_5754);
nand U7495 (N_7495,N_4106,N_4928);
nand U7496 (N_7496,N_4527,N_3861);
or U7497 (N_7497,N_5396,N_3446);
xor U7498 (N_7498,N_5539,N_4262);
or U7499 (N_7499,N_5625,N_3852);
or U7500 (N_7500,N_4294,N_5686);
xnor U7501 (N_7501,N_5578,N_3431);
or U7502 (N_7502,N_5751,N_4902);
or U7503 (N_7503,N_5642,N_5948);
nor U7504 (N_7504,N_4794,N_4904);
or U7505 (N_7505,N_4237,N_5354);
or U7506 (N_7506,N_3625,N_5004);
or U7507 (N_7507,N_4975,N_3976);
nand U7508 (N_7508,N_5897,N_5425);
nor U7509 (N_7509,N_3236,N_5662);
and U7510 (N_7510,N_4109,N_3816);
nor U7511 (N_7511,N_5136,N_5497);
xnor U7512 (N_7512,N_5237,N_5335);
or U7513 (N_7513,N_4717,N_3402);
nor U7514 (N_7514,N_3408,N_3760);
or U7515 (N_7515,N_3161,N_5313);
or U7516 (N_7516,N_4959,N_3217);
and U7517 (N_7517,N_4407,N_5779);
nor U7518 (N_7518,N_3954,N_4031);
nand U7519 (N_7519,N_3424,N_3282);
nor U7520 (N_7520,N_3501,N_3225);
and U7521 (N_7521,N_5534,N_4690);
xor U7522 (N_7522,N_5732,N_3533);
xnor U7523 (N_7523,N_4318,N_5551);
xor U7524 (N_7524,N_3634,N_5615);
nand U7525 (N_7525,N_4421,N_4024);
nand U7526 (N_7526,N_5816,N_5068);
nand U7527 (N_7527,N_5290,N_4421);
nor U7528 (N_7528,N_5893,N_4243);
and U7529 (N_7529,N_4968,N_4100);
nor U7530 (N_7530,N_4917,N_5766);
nor U7531 (N_7531,N_4838,N_5394);
nand U7532 (N_7532,N_4754,N_3812);
or U7533 (N_7533,N_5713,N_3121);
xnor U7534 (N_7534,N_3604,N_5098);
nand U7535 (N_7535,N_3072,N_3475);
nand U7536 (N_7536,N_3113,N_5415);
xor U7537 (N_7537,N_5757,N_5192);
or U7538 (N_7538,N_5598,N_3256);
nor U7539 (N_7539,N_3175,N_4437);
nor U7540 (N_7540,N_3465,N_5102);
xnor U7541 (N_7541,N_5524,N_3499);
and U7542 (N_7542,N_4434,N_5729);
and U7543 (N_7543,N_5394,N_4679);
nor U7544 (N_7544,N_3882,N_4626);
and U7545 (N_7545,N_3156,N_4295);
nand U7546 (N_7546,N_5608,N_4025);
xor U7547 (N_7547,N_3011,N_5723);
nand U7548 (N_7548,N_5835,N_3155);
or U7549 (N_7549,N_3536,N_3691);
nand U7550 (N_7550,N_5771,N_3098);
nor U7551 (N_7551,N_3544,N_3417);
nand U7552 (N_7552,N_4467,N_4837);
or U7553 (N_7553,N_5739,N_4503);
nor U7554 (N_7554,N_4805,N_4468);
nand U7555 (N_7555,N_4140,N_3245);
nand U7556 (N_7556,N_3861,N_5220);
and U7557 (N_7557,N_5077,N_5517);
nor U7558 (N_7558,N_4955,N_5768);
nand U7559 (N_7559,N_3511,N_3441);
and U7560 (N_7560,N_4193,N_5563);
or U7561 (N_7561,N_3808,N_5745);
or U7562 (N_7562,N_3227,N_5261);
and U7563 (N_7563,N_5259,N_4176);
and U7564 (N_7564,N_3476,N_4874);
or U7565 (N_7565,N_5615,N_4263);
nor U7566 (N_7566,N_3030,N_5041);
nand U7567 (N_7567,N_4223,N_5309);
nor U7568 (N_7568,N_4275,N_3760);
nand U7569 (N_7569,N_5493,N_3627);
nor U7570 (N_7570,N_3777,N_4826);
nand U7571 (N_7571,N_4196,N_5888);
or U7572 (N_7572,N_3576,N_3942);
xnor U7573 (N_7573,N_3011,N_5963);
nor U7574 (N_7574,N_4785,N_5128);
nor U7575 (N_7575,N_3615,N_5182);
xnor U7576 (N_7576,N_3638,N_3995);
xor U7577 (N_7577,N_4525,N_5622);
or U7578 (N_7578,N_4693,N_3126);
and U7579 (N_7579,N_3642,N_3691);
xnor U7580 (N_7580,N_4977,N_4439);
and U7581 (N_7581,N_4852,N_5712);
nand U7582 (N_7582,N_4601,N_3218);
nor U7583 (N_7583,N_3585,N_3798);
and U7584 (N_7584,N_4662,N_5910);
and U7585 (N_7585,N_3824,N_3169);
nor U7586 (N_7586,N_3732,N_3679);
nand U7587 (N_7587,N_5679,N_4358);
or U7588 (N_7588,N_5398,N_5912);
and U7589 (N_7589,N_5899,N_4556);
and U7590 (N_7590,N_3427,N_4234);
nand U7591 (N_7591,N_3549,N_5593);
and U7592 (N_7592,N_3787,N_4375);
xnor U7593 (N_7593,N_3063,N_5747);
and U7594 (N_7594,N_5142,N_5952);
nand U7595 (N_7595,N_4281,N_3680);
nand U7596 (N_7596,N_5789,N_4759);
or U7597 (N_7597,N_3030,N_4658);
nand U7598 (N_7598,N_4300,N_4841);
nor U7599 (N_7599,N_3863,N_3463);
or U7600 (N_7600,N_5449,N_4427);
or U7601 (N_7601,N_5534,N_4726);
and U7602 (N_7602,N_4045,N_3574);
nor U7603 (N_7603,N_5838,N_4338);
and U7604 (N_7604,N_4140,N_3901);
and U7605 (N_7605,N_4673,N_3092);
or U7606 (N_7606,N_3115,N_4438);
or U7607 (N_7607,N_5711,N_5568);
and U7608 (N_7608,N_4958,N_3518);
and U7609 (N_7609,N_4271,N_3772);
and U7610 (N_7610,N_3827,N_3523);
nor U7611 (N_7611,N_4047,N_4227);
or U7612 (N_7612,N_4446,N_5040);
xor U7613 (N_7613,N_5793,N_3752);
nor U7614 (N_7614,N_3240,N_5411);
and U7615 (N_7615,N_4418,N_3626);
nand U7616 (N_7616,N_5978,N_4784);
or U7617 (N_7617,N_4792,N_5472);
nand U7618 (N_7618,N_4021,N_5239);
nor U7619 (N_7619,N_5179,N_5786);
nor U7620 (N_7620,N_5811,N_5667);
and U7621 (N_7621,N_4562,N_5586);
and U7622 (N_7622,N_4238,N_4504);
nor U7623 (N_7623,N_5631,N_5238);
nor U7624 (N_7624,N_3634,N_5140);
nand U7625 (N_7625,N_3387,N_3937);
and U7626 (N_7626,N_3909,N_4629);
xnor U7627 (N_7627,N_3828,N_3859);
nand U7628 (N_7628,N_5922,N_4257);
or U7629 (N_7629,N_4572,N_3757);
and U7630 (N_7630,N_4294,N_3615);
or U7631 (N_7631,N_5929,N_4091);
xor U7632 (N_7632,N_3324,N_3545);
nor U7633 (N_7633,N_4064,N_5215);
or U7634 (N_7634,N_4134,N_3655);
nor U7635 (N_7635,N_5437,N_3385);
and U7636 (N_7636,N_3096,N_5363);
and U7637 (N_7637,N_3288,N_5933);
nor U7638 (N_7638,N_5237,N_4429);
or U7639 (N_7639,N_3223,N_5655);
or U7640 (N_7640,N_5854,N_5306);
xor U7641 (N_7641,N_5783,N_4276);
nand U7642 (N_7642,N_3016,N_5250);
and U7643 (N_7643,N_4476,N_5432);
or U7644 (N_7644,N_4849,N_5717);
nand U7645 (N_7645,N_4838,N_3748);
xor U7646 (N_7646,N_5400,N_3945);
nand U7647 (N_7647,N_4432,N_5154);
and U7648 (N_7648,N_5733,N_5300);
xor U7649 (N_7649,N_5269,N_5654);
or U7650 (N_7650,N_4888,N_3399);
nand U7651 (N_7651,N_5524,N_4560);
nor U7652 (N_7652,N_4908,N_3162);
nor U7653 (N_7653,N_4798,N_3452);
nand U7654 (N_7654,N_3479,N_5559);
or U7655 (N_7655,N_3781,N_5139);
and U7656 (N_7656,N_3551,N_5994);
or U7657 (N_7657,N_3751,N_4738);
or U7658 (N_7658,N_4463,N_4974);
nand U7659 (N_7659,N_5750,N_4628);
nand U7660 (N_7660,N_5520,N_4671);
or U7661 (N_7661,N_5113,N_4356);
and U7662 (N_7662,N_3676,N_5048);
nand U7663 (N_7663,N_4022,N_5119);
nor U7664 (N_7664,N_3712,N_5700);
and U7665 (N_7665,N_3471,N_4686);
nor U7666 (N_7666,N_4854,N_3006);
and U7667 (N_7667,N_3294,N_3328);
nor U7668 (N_7668,N_4720,N_5703);
or U7669 (N_7669,N_4772,N_3941);
and U7670 (N_7670,N_4040,N_3002);
nand U7671 (N_7671,N_4046,N_5586);
and U7672 (N_7672,N_3916,N_5323);
nand U7673 (N_7673,N_4396,N_4823);
nor U7674 (N_7674,N_5837,N_3069);
or U7675 (N_7675,N_5046,N_3114);
or U7676 (N_7676,N_4365,N_3879);
nor U7677 (N_7677,N_4350,N_3292);
nor U7678 (N_7678,N_4443,N_3200);
xor U7679 (N_7679,N_3397,N_5596);
and U7680 (N_7680,N_5582,N_5545);
or U7681 (N_7681,N_4349,N_5355);
or U7682 (N_7682,N_4737,N_3769);
or U7683 (N_7683,N_4215,N_4789);
or U7684 (N_7684,N_5961,N_4841);
or U7685 (N_7685,N_4596,N_3471);
nand U7686 (N_7686,N_4057,N_4086);
nand U7687 (N_7687,N_5061,N_5792);
or U7688 (N_7688,N_5467,N_3891);
xor U7689 (N_7689,N_3253,N_4441);
or U7690 (N_7690,N_4497,N_5913);
and U7691 (N_7691,N_5841,N_4964);
nand U7692 (N_7692,N_5020,N_4796);
or U7693 (N_7693,N_4789,N_5144);
xor U7694 (N_7694,N_4293,N_5573);
nor U7695 (N_7695,N_5454,N_5432);
nand U7696 (N_7696,N_4206,N_5392);
or U7697 (N_7697,N_5275,N_5250);
nand U7698 (N_7698,N_3482,N_4948);
nor U7699 (N_7699,N_3516,N_3809);
and U7700 (N_7700,N_4635,N_3706);
or U7701 (N_7701,N_4678,N_5922);
and U7702 (N_7702,N_5214,N_4379);
and U7703 (N_7703,N_4583,N_5023);
or U7704 (N_7704,N_4836,N_5707);
or U7705 (N_7705,N_5814,N_4983);
xnor U7706 (N_7706,N_3439,N_5784);
nand U7707 (N_7707,N_3152,N_5802);
nand U7708 (N_7708,N_5427,N_5232);
xor U7709 (N_7709,N_3747,N_3285);
nor U7710 (N_7710,N_3326,N_5342);
nor U7711 (N_7711,N_3667,N_5205);
and U7712 (N_7712,N_5057,N_5291);
and U7713 (N_7713,N_3703,N_4129);
nand U7714 (N_7714,N_5433,N_3462);
and U7715 (N_7715,N_5284,N_4754);
xor U7716 (N_7716,N_4897,N_5493);
xnor U7717 (N_7717,N_5170,N_4739);
xnor U7718 (N_7718,N_4523,N_3564);
nor U7719 (N_7719,N_3370,N_4362);
nand U7720 (N_7720,N_3667,N_3693);
nand U7721 (N_7721,N_5254,N_3969);
and U7722 (N_7722,N_4551,N_3227);
and U7723 (N_7723,N_5366,N_5057);
or U7724 (N_7724,N_3133,N_5425);
or U7725 (N_7725,N_4902,N_4733);
or U7726 (N_7726,N_3097,N_5688);
or U7727 (N_7727,N_4524,N_5900);
and U7728 (N_7728,N_5830,N_5784);
and U7729 (N_7729,N_4916,N_3963);
or U7730 (N_7730,N_4636,N_5043);
nand U7731 (N_7731,N_3807,N_3589);
nand U7732 (N_7732,N_3418,N_3469);
or U7733 (N_7733,N_4147,N_5241);
nor U7734 (N_7734,N_3230,N_4119);
nand U7735 (N_7735,N_5619,N_5589);
xor U7736 (N_7736,N_3053,N_5592);
or U7737 (N_7737,N_3309,N_3660);
nor U7738 (N_7738,N_5486,N_5299);
nand U7739 (N_7739,N_5804,N_3253);
nand U7740 (N_7740,N_4835,N_3778);
or U7741 (N_7741,N_3144,N_4268);
or U7742 (N_7742,N_5588,N_4182);
nor U7743 (N_7743,N_3919,N_5827);
nand U7744 (N_7744,N_4641,N_4315);
or U7745 (N_7745,N_5090,N_4871);
nand U7746 (N_7746,N_4950,N_5799);
nand U7747 (N_7747,N_5815,N_4563);
nand U7748 (N_7748,N_4021,N_4817);
xnor U7749 (N_7749,N_4388,N_5036);
nor U7750 (N_7750,N_3996,N_5830);
or U7751 (N_7751,N_3314,N_5270);
nand U7752 (N_7752,N_5682,N_5713);
nand U7753 (N_7753,N_5763,N_3076);
or U7754 (N_7754,N_4335,N_4525);
nor U7755 (N_7755,N_3729,N_4653);
nand U7756 (N_7756,N_3693,N_5094);
nand U7757 (N_7757,N_4178,N_5425);
or U7758 (N_7758,N_5563,N_4324);
and U7759 (N_7759,N_4448,N_3559);
and U7760 (N_7760,N_5209,N_3057);
and U7761 (N_7761,N_5065,N_4178);
or U7762 (N_7762,N_5541,N_4356);
nor U7763 (N_7763,N_4981,N_4395);
or U7764 (N_7764,N_4592,N_3199);
nand U7765 (N_7765,N_5655,N_4360);
xor U7766 (N_7766,N_5816,N_4162);
nor U7767 (N_7767,N_5088,N_5095);
nand U7768 (N_7768,N_4091,N_3728);
or U7769 (N_7769,N_3948,N_5885);
nand U7770 (N_7770,N_5953,N_3487);
and U7771 (N_7771,N_4381,N_4504);
nand U7772 (N_7772,N_4569,N_3951);
nor U7773 (N_7773,N_4514,N_5511);
nor U7774 (N_7774,N_4771,N_4320);
xnor U7775 (N_7775,N_3749,N_3989);
and U7776 (N_7776,N_5037,N_5122);
nand U7777 (N_7777,N_5069,N_4658);
or U7778 (N_7778,N_4088,N_4587);
or U7779 (N_7779,N_4433,N_5571);
nand U7780 (N_7780,N_4452,N_4100);
or U7781 (N_7781,N_4286,N_5769);
xnor U7782 (N_7782,N_4507,N_5247);
and U7783 (N_7783,N_4801,N_5931);
nor U7784 (N_7784,N_4868,N_3206);
and U7785 (N_7785,N_3507,N_3499);
nand U7786 (N_7786,N_3195,N_4766);
and U7787 (N_7787,N_3331,N_4410);
nand U7788 (N_7788,N_3193,N_5177);
and U7789 (N_7789,N_4977,N_5395);
nor U7790 (N_7790,N_5088,N_5834);
nor U7791 (N_7791,N_5375,N_4452);
nand U7792 (N_7792,N_4829,N_5258);
and U7793 (N_7793,N_3090,N_5092);
or U7794 (N_7794,N_3204,N_4824);
nor U7795 (N_7795,N_3606,N_4882);
and U7796 (N_7796,N_5215,N_3388);
xnor U7797 (N_7797,N_4550,N_5224);
xnor U7798 (N_7798,N_4979,N_4839);
or U7799 (N_7799,N_5884,N_4306);
and U7800 (N_7800,N_5443,N_5782);
and U7801 (N_7801,N_4154,N_4581);
and U7802 (N_7802,N_3157,N_3698);
nand U7803 (N_7803,N_3224,N_3258);
nand U7804 (N_7804,N_4836,N_5220);
or U7805 (N_7805,N_4331,N_5253);
nor U7806 (N_7806,N_5813,N_5109);
xnor U7807 (N_7807,N_5650,N_5766);
nand U7808 (N_7808,N_3939,N_4044);
nor U7809 (N_7809,N_5952,N_4215);
or U7810 (N_7810,N_4401,N_5197);
and U7811 (N_7811,N_3410,N_4201);
or U7812 (N_7812,N_5700,N_4458);
and U7813 (N_7813,N_3260,N_5657);
nand U7814 (N_7814,N_5971,N_5893);
or U7815 (N_7815,N_3067,N_5726);
xnor U7816 (N_7816,N_5237,N_3723);
and U7817 (N_7817,N_4847,N_3694);
nor U7818 (N_7818,N_4226,N_5156);
or U7819 (N_7819,N_3898,N_3912);
nor U7820 (N_7820,N_5715,N_4999);
nor U7821 (N_7821,N_4817,N_3411);
nor U7822 (N_7822,N_5835,N_5711);
nand U7823 (N_7823,N_4920,N_3640);
nor U7824 (N_7824,N_3525,N_3979);
xnor U7825 (N_7825,N_5474,N_4886);
xnor U7826 (N_7826,N_3614,N_5896);
or U7827 (N_7827,N_3434,N_5758);
nor U7828 (N_7828,N_3394,N_3483);
xnor U7829 (N_7829,N_3641,N_4744);
and U7830 (N_7830,N_4641,N_3012);
nor U7831 (N_7831,N_3681,N_5927);
and U7832 (N_7832,N_3468,N_5228);
nor U7833 (N_7833,N_5607,N_4003);
and U7834 (N_7834,N_5849,N_3956);
nor U7835 (N_7835,N_3387,N_5501);
and U7836 (N_7836,N_4972,N_3467);
nand U7837 (N_7837,N_4920,N_5108);
nand U7838 (N_7838,N_5256,N_4408);
or U7839 (N_7839,N_5524,N_4625);
nand U7840 (N_7840,N_3078,N_3625);
and U7841 (N_7841,N_4502,N_3368);
nand U7842 (N_7842,N_5804,N_4762);
nand U7843 (N_7843,N_5749,N_5093);
nor U7844 (N_7844,N_4409,N_5436);
and U7845 (N_7845,N_3875,N_5209);
and U7846 (N_7846,N_3791,N_3141);
nor U7847 (N_7847,N_5572,N_4422);
or U7848 (N_7848,N_3261,N_4753);
nand U7849 (N_7849,N_3289,N_3777);
nand U7850 (N_7850,N_3311,N_3027);
and U7851 (N_7851,N_4346,N_4015);
or U7852 (N_7852,N_3180,N_4900);
nor U7853 (N_7853,N_4191,N_3715);
and U7854 (N_7854,N_4960,N_4197);
nor U7855 (N_7855,N_4767,N_4029);
and U7856 (N_7856,N_3786,N_5556);
nor U7857 (N_7857,N_5604,N_5479);
nand U7858 (N_7858,N_3136,N_5252);
xnor U7859 (N_7859,N_3267,N_5812);
or U7860 (N_7860,N_5479,N_4527);
or U7861 (N_7861,N_4620,N_3155);
nor U7862 (N_7862,N_5386,N_4999);
nand U7863 (N_7863,N_5617,N_5839);
nor U7864 (N_7864,N_3235,N_3532);
nor U7865 (N_7865,N_3898,N_5168);
xnor U7866 (N_7866,N_3784,N_4561);
nand U7867 (N_7867,N_5849,N_3911);
nor U7868 (N_7868,N_5115,N_4342);
and U7869 (N_7869,N_3493,N_5271);
nand U7870 (N_7870,N_3584,N_4375);
xnor U7871 (N_7871,N_4051,N_5791);
nor U7872 (N_7872,N_3309,N_3961);
nor U7873 (N_7873,N_4795,N_3614);
nand U7874 (N_7874,N_5779,N_5463);
nand U7875 (N_7875,N_3733,N_3210);
xnor U7876 (N_7876,N_3227,N_4414);
nor U7877 (N_7877,N_5652,N_3399);
or U7878 (N_7878,N_4110,N_4592);
or U7879 (N_7879,N_3731,N_4104);
and U7880 (N_7880,N_5408,N_5026);
and U7881 (N_7881,N_3402,N_4393);
nor U7882 (N_7882,N_4933,N_4045);
nand U7883 (N_7883,N_3138,N_3243);
and U7884 (N_7884,N_5391,N_3902);
or U7885 (N_7885,N_3893,N_5518);
or U7886 (N_7886,N_4637,N_5859);
nand U7887 (N_7887,N_4676,N_3735);
nor U7888 (N_7888,N_5276,N_5371);
or U7889 (N_7889,N_3002,N_5114);
nor U7890 (N_7890,N_4043,N_3169);
xor U7891 (N_7891,N_5698,N_4680);
and U7892 (N_7892,N_5251,N_5427);
nand U7893 (N_7893,N_3934,N_5229);
and U7894 (N_7894,N_3220,N_4258);
nor U7895 (N_7895,N_3611,N_3840);
nand U7896 (N_7896,N_3767,N_3830);
and U7897 (N_7897,N_4943,N_5359);
or U7898 (N_7898,N_4559,N_5529);
or U7899 (N_7899,N_5115,N_3196);
or U7900 (N_7900,N_5062,N_5322);
nand U7901 (N_7901,N_4140,N_4838);
xor U7902 (N_7902,N_3991,N_5652);
nand U7903 (N_7903,N_4372,N_4290);
nand U7904 (N_7904,N_4795,N_4966);
nand U7905 (N_7905,N_3882,N_3811);
nor U7906 (N_7906,N_5146,N_3579);
and U7907 (N_7907,N_3306,N_3955);
nand U7908 (N_7908,N_4045,N_4089);
nor U7909 (N_7909,N_3929,N_5844);
xor U7910 (N_7910,N_3681,N_3564);
and U7911 (N_7911,N_5840,N_4279);
or U7912 (N_7912,N_5805,N_4497);
nor U7913 (N_7913,N_4213,N_4354);
nor U7914 (N_7914,N_4747,N_4835);
or U7915 (N_7915,N_4501,N_5400);
nor U7916 (N_7916,N_5067,N_5211);
or U7917 (N_7917,N_3228,N_4262);
nor U7918 (N_7918,N_4109,N_5601);
nor U7919 (N_7919,N_5146,N_4073);
and U7920 (N_7920,N_3987,N_3076);
or U7921 (N_7921,N_3997,N_5082);
nor U7922 (N_7922,N_4446,N_4863);
nor U7923 (N_7923,N_3728,N_4259);
nand U7924 (N_7924,N_3185,N_5877);
and U7925 (N_7925,N_4186,N_4636);
xor U7926 (N_7926,N_3972,N_4807);
nor U7927 (N_7927,N_5007,N_4938);
or U7928 (N_7928,N_5253,N_4401);
nand U7929 (N_7929,N_3407,N_4023);
and U7930 (N_7930,N_3313,N_5590);
and U7931 (N_7931,N_4759,N_3399);
or U7932 (N_7932,N_5207,N_5572);
and U7933 (N_7933,N_5170,N_4129);
nand U7934 (N_7934,N_5268,N_4880);
nor U7935 (N_7935,N_3588,N_5437);
and U7936 (N_7936,N_4510,N_3669);
and U7937 (N_7937,N_4896,N_5268);
or U7938 (N_7938,N_3327,N_5509);
or U7939 (N_7939,N_4777,N_4114);
or U7940 (N_7940,N_5461,N_4014);
and U7941 (N_7941,N_5301,N_5690);
nand U7942 (N_7942,N_4782,N_4192);
or U7943 (N_7943,N_5986,N_5513);
nor U7944 (N_7944,N_3734,N_3500);
nor U7945 (N_7945,N_5155,N_5805);
nor U7946 (N_7946,N_5575,N_3182);
nand U7947 (N_7947,N_5876,N_3814);
nor U7948 (N_7948,N_5684,N_5545);
nand U7949 (N_7949,N_3734,N_3516);
and U7950 (N_7950,N_3446,N_4932);
and U7951 (N_7951,N_3180,N_4214);
nor U7952 (N_7952,N_4232,N_4517);
nand U7953 (N_7953,N_3545,N_4049);
and U7954 (N_7954,N_3110,N_5705);
nand U7955 (N_7955,N_3880,N_3093);
nand U7956 (N_7956,N_3952,N_3649);
and U7957 (N_7957,N_4053,N_5650);
nor U7958 (N_7958,N_5453,N_4549);
and U7959 (N_7959,N_3239,N_5807);
and U7960 (N_7960,N_3256,N_4970);
and U7961 (N_7961,N_3464,N_5437);
or U7962 (N_7962,N_3751,N_3481);
nand U7963 (N_7963,N_5349,N_3996);
or U7964 (N_7964,N_4327,N_5639);
or U7965 (N_7965,N_4190,N_3164);
xor U7966 (N_7966,N_5759,N_4319);
nand U7967 (N_7967,N_3982,N_3129);
nor U7968 (N_7968,N_5889,N_4253);
and U7969 (N_7969,N_5368,N_5079);
nor U7970 (N_7970,N_4017,N_4268);
and U7971 (N_7971,N_3224,N_4875);
xnor U7972 (N_7972,N_3379,N_5416);
nor U7973 (N_7973,N_5336,N_5070);
nor U7974 (N_7974,N_3728,N_5637);
xor U7975 (N_7975,N_5656,N_3857);
and U7976 (N_7976,N_4891,N_5761);
or U7977 (N_7977,N_4291,N_5395);
nor U7978 (N_7978,N_3218,N_5693);
and U7979 (N_7979,N_4982,N_3204);
nand U7980 (N_7980,N_4811,N_4727);
and U7981 (N_7981,N_3566,N_3433);
nor U7982 (N_7982,N_3087,N_3398);
nand U7983 (N_7983,N_4910,N_3327);
and U7984 (N_7984,N_3727,N_3861);
nand U7985 (N_7985,N_3856,N_5728);
and U7986 (N_7986,N_4498,N_5252);
or U7987 (N_7987,N_3722,N_3225);
and U7988 (N_7988,N_5052,N_5103);
or U7989 (N_7989,N_4239,N_4612);
or U7990 (N_7990,N_5019,N_4719);
and U7991 (N_7991,N_5835,N_5632);
xnor U7992 (N_7992,N_5488,N_5427);
and U7993 (N_7993,N_3019,N_3454);
or U7994 (N_7994,N_3130,N_5468);
nor U7995 (N_7995,N_4475,N_3091);
and U7996 (N_7996,N_5281,N_4541);
nor U7997 (N_7997,N_5307,N_5524);
xor U7998 (N_7998,N_3499,N_3506);
nor U7999 (N_7999,N_3257,N_3532);
xnor U8000 (N_8000,N_4485,N_4530);
and U8001 (N_8001,N_4711,N_4225);
nor U8002 (N_8002,N_3781,N_4679);
nand U8003 (N_8003,N_4859,N_3670);
or U8004 (N_8004,N_5159,N_5737);
nand U8005 (N_8005,N_4059,N_4186);
or U8006 (N_8006,N_3632,N_3998);
and U8007 (N_8007,N_3312,N_4318);
and U8008 (N_8008,N_4275,N_3419);
xnor U8009 (N_8009,N_3959,N_5078);
or U8010 (N_8010,N_3805,N_4238);
or U8011 (N_8011,N_5727,N_5896);
nand U8012 (N_8012,N_4750,N_3450);
nand U8013 (N_8013,N_3790,N_4352);
xnor U8014 (N_8014,N_5267,N_3746);
nand U8015 (N_8015,N_5397,N_4426);
nor U8016 (N_8016,N_5092,N_3572);
nand U8017 (N_8017,N_4184,N_5081);
or U8018 (N_8018,N_5739,N_4175);
nor U8019 (N_8019,N_3750,N_4857);
or U8020 (N_8020,N_3213,N_4598);
nand U8021 (N_8021,N_4676,N_4204);
nor U8022 (N_8022,N_3383,N_5092);
nand U8023 (N_8023,N_5142,N_3742);
nand U8024 (N_8024,N_5464,N_3981);
nand U8025 (N_8025,N_5535,N_4577);
nor U8026 (N_8026,N_5623,N_3194);
and U8027 (N_8027,N_4952,N_3315);
or U8028 (N_8028,N_3663,N_4207);
or U8029 (N_8029,N_3641,N_5580);
or U8030 (N_8030,N_4412,N_5114);
nor U8031 (N_8031,N_3613,N_5883);
xnor U8032 (N_8032,N_4126,N_5155);
or U8033 (N_8033,N_4612,N_5219);
and U8034 (N_8034,N_5777,N_5753);
and U8035 (N_8035,N_4729,N_4884);
and U8036 (N_8036,N_4404,N_4615);
nor U8037 (N_8037,N_4377,N_3237);
and U8038 (N_8038,N_3739,N_5301);
and U8039 (N_8039,N_3151,N_3856);
nand U8040 (N_8040,N_5490,N_4940);
nand U8041 (N_8041,N_3436,N_3104);
or U8042 (N_8042,N_5251,N_5998);
nand U8043 (N_8043,N_5940,N_5057);
nor U8044 (N_8044,N_5797,N_5047);
nor U8045 (N_8045,N_4833,N_3748);
nand U8046 (N_8046,N_5581,N_5712);
nor U8047 (N_8047,N_5234,N_4399);
or U8048 (N_8048,N_3575,N_3697);
nand U8049 (N_8049,N_5324,N_4512);
nand U8050 (N_8050,N_5870,N_4617);
or U8051 (N_8051,N_5585,N_4797);
and U8052 (N_8052,N_5497,N_3035);
nor U8053 (N_8053,N_4527,N_5354);
or U8054 (N_8054,N_4807,N_4254);
or U8055 (N_8055,N_5298,N_4095);
nand U8056 (N_8056,N_4125,N_5807);
nand U8057 (N_8057,N_4924,N_5310);
nand U8058 (N_8058,N_3296,N_5957);
and U8059 (N_8059,N_5333,N_3432);
and U8060 (N_8060,N_5387,N_4199);
and U8061 (N_8061,N_4347,N_5521);
or U8062 (N_8062,N_5086,N_4749);
or U8063 (N_8063,N_4817,N_3962);
nand U8064 (N_8064,N_3394,N_3165);
nor U8065 (N_8065,N_5851,N_3691);
nor U8066 (N_8066,N_5434,N_4186);
nor U8067 (N_8067,N_5263,N_4795);
nand U8068 (N_8068,N_3309,N_4251);
and U8069 (N_8069,N_5175,N_5749);
or U8070 (N_8070,N_5286,N_4821);
nand U8071 (N_8071,N_5991,N_3115);
nand U8072 (N_8072,N_5454,N_4425);
and U8073 (N_8073,N_3529,N_4574);
and U8074 (N_8074,N_3450,N_4598);
nand U8075 (N_8075,N_5207,N_4696);
nand U8076 (N_8076,N_3231,N_3586);
nor U8077 (N_8077,N_3568,N_4540);
nor U8078 (N_8078,N_3845,N_5408);
or U8079 (N_8079,N_4370,N_5674);
xor U8080 (N_8080,N_4323,N_5167);
and U8081 (N_8081,N_5028,N_5885);
nor U8082 (N_8082,N_3381,N_3071);
and U8083 (N_8083,N_5422,N_3353);
xnor U8084 (N_8084,N_5255,N_5791);
nand U8085 (N_8085,N_5707,N_3345);
nand U8086 (N_8086,N_4179,N_5096);
or U8087 (N_8087,N_3015,N_5712);
nand U8088 (N_8088,N_3947,N_4991);
nand U8089 (N_8089,N_5113,N_5338);
or U8090 (N_8090,N_4964,N_5336);
nor U8091 (N_8091,N_5443,N_5848);
or U8092 (N_8092,N_5832,N_4788);
or U8093 (N_8093,N_3031,N_5630);
or U8094 (N_8094,N_5316,N_3876);
nor U8095 (N_8095,N_3182,N_4335);
nor U8096 (N_8096,N_3508,N_5285);
nor U8097 (N_8097,N_4202,N_4657);
and U8098 (N_8098,N_5973,N_5739);
or U8099 (N_8099,N_3209,N_4515);
nor U8100 (N_8100,N_3668,N_4806);
or U8101 (N_8101,N_4019,N_4194);
or U8102 (N_8102,N_3871,N_5472);
xnor U8103 (N_8103,N_4751,N_3590);
nand U8104 (N_8104,N_3190,N_4338);
or U8105 (N_8105,N_5992,N_3561);
or U8106 (N_8106,N_3986,N_3777);
and U8107 (N_8107,N_4949,N_3075);
nand U8108 (N_8108,N_5772,N_4637);
or U8109 (N_8109,N_5526,N_4691);
and U8110 (N_8110,N_5990,N_5533);
nand U8111 (N_8111,N_5245,N_5976);
xnor U8112 (N_8112,N_4585,N_4215);
xor U8113 (N_8113,N_3510,N_5454);
or U8114 (N_8114,N_5175,N_5297);
nand U8115 (N_8115,N_3544,N_5336);
and U8116 (N_8116,N_5579,N_3722);
nor U8117 (N_8117,N_5141,N_3237);
and U8118 (N_8118,N_4004,N_4804);
nor U8119 (N_8119,N_3611,N_5581);
or U8120 (N_8120,N_4486,N_5354);
nand U8121 (N_8121,N_4018,N_5160);
or U8122 (N_8122,N_3644,N_4088);
or U8123 (N_8123,N_3097,N_4238);
nor U8124 (N_8124,N_4781,N_3058);
nand U8125 (N_8125,N_5312,N_4745);
nor U8126 (N_8126,N_3962,N_3820);
xnor U8127 (N_8127,N_4610,N_3296);
or U8128 (N_8128,N_4546,N_3914);
nor U8129 (N_8129,N_5079,N_4448);
and U8130 (N_8130,N_3165,N_4507);
and U8131 (N_8131,N_5286,N_3617);
and U8132 (N_8132,N_4531,N_3052);
nor U8133 (N_8133,N_5589,N_3050);
and U8134 (N_8134,N_3139,N_3923);
and U8135 (N_8135,N_4734,N_4020);
nor U8136 (N_8136,N_3461,N_3019);
nand U8137 (N_8137,N_3752,N_4336);
nor U8138 (N_8138,N_3176,N_3273);
or U8139 (N_8139,N_4764,N_5783);
nor U8140 (N_8140,N_4927,N_4980);
and U8141 (N_8141,N_4061,N_3294);
or U8142 (N_8142,N_5963,N_4044);
and U8143 (N_8143,N_3945,N_3927);
and U8144 (N_8144,N_5042,N_3504);
or U8145 (N_8145,N_3902,N_4168);
nand U8146 (N_8146,N_3752,N_3936);
xor U8147 (N_8147,N_5891,N_5465);
and U8148 (N_8148,N_5875,N_3212);
or U8149 (N_8149,N_3453,N_4140);
nand U8150 (N_8150,N_4682,N_5573);
nand U8151 (N_8151,N_4534,N_3361);
or U8152 (N_8152,N_4824,N_4799);
or U8153 (N_8153,N_4620,N_4232);
nor U8154 (N_8154,N_4796,N_3621);
xor U8155 (N_8155,N_5152,N_4705);
xnor U8156 (N_8156,N_3064,N_4624);
or U8157 (N_8157,N_5053,N_3707);
or U8158 (N_8158,N_4360,N_4957);
nor U8159 (N_8159,N_5409,N_3105);
or U8160 (N_8160,N_4583,N_4809);
nand U8161 (N_8161,N_3208,N_5375);
and U8162 (N_8162,N_5421,N_3899);
xnor U8163 (N_8163,N_4431,N_4626);
nand U8164 (N_8164,N_4247,N_5111);
or U8165 (N_8165,N_5608,N_5553);
nor U8166 (N_8166,N_5765,N_4277);
nor U8167 (N_8167,N_5948,N_4137);
nor U8168 (N_8168,N_3771,N_4741);
or U8169 (N_8169,N_3755,N_5412);
nand U8170 (N_8170,N_4738,N_4711);
and U8171 (N_8171,N_4638,N_5809);
nor U8172 (N_8172,N_5335,N_4339);
nor U8173 (N_8173,N_5287,N_3680);
nor U8174 (N_8174,N_3633,N_4559);
nor U8175 (N_8175,N_5743,N_4116);
or U8176 (N_8176,N_5537,N_5362);
or U8177 (N_8177,N_5457,N_5989);
nor U8178 (N_8178,N_4250,N_4309);
and U8179 (N_8179,N_3755,N_5371);
nand U8180 (N_8180,N_3021,N_4619);
and U8181 (N_8181,N_4948,N_4034);
xnor U8182 (N_8182,N_3829,N_3379);
or U8183 (N_8183,N_3137,N_5589);
or U8184 (N_8184,N_5834,N_4110);
and U8185 (N_8185,N_4328,N_3176);
and U8186 (N_8186,N_4086,N_3053);
nor U8187 (N_8187,N_3959,N_5120);
nor U8188 (N_8188,N_3778,N_3488);
or U8189 (N_8189,N_5692,N_5253);
nor U8190 (N_8190,N_3586,N_4176);
nand U8191 (N_8191,N_3289,N_5134);
or U8192 (N_8192,N_5789,N_5876);
nor U8193 (N_8193,N_5421,N_5884);
nor U8194 (N_8194,N_3655,N_4149);
nand U8195 (N_8195,N_3671,N_4613);
or U8196 (N_8196,N_3527,N_3086);
and U8197 (N_8197,N_3725,N_4956);
or U8198 (N_8198,N_4537,N_4226);
or U8199 (N_8199,N_3647,N_5036);
nand U8200 (N_8200,N_3254,N_4103);
nand U8201 (N_8201,N_5666,N_4345);
nand U8202 (N_8202,N_4551,N_5724);
nand U8203 (N_8203,N_3222,N_5035);
nand U8204 (N_8204,N_4641,N_3061);
or U8205 (N_8205,N_3375,N_4476);
nor U8206 (N_8206,N_3789,N_4858);
or U8207 (N_8207,N_5109,N_3239);
nor U8208 (N_8208,N_3966,N_4455);
nand U8209 (N_8209,N_5438,N_5249);
and U8210 (N_8210,N_5281,N_5802);
and U8211 (N_8211,N_5455,N_5847);
or U8212 (N_8212,N_4814,N_4622);
nor U8213 (N_8213,N_4460,N_4977);
nor U8214 (N_8214,N_4176,N_5281);
and U8215 (N_8215,N_5326,N_5407);
and U8216 (N_8216,N_3651,N_5909);
xor U8217 (N_8217,N_3652,N_3738);
or U8218 (N_8218,N_3652,N_4576);
nor U8219 (N_8219,N_5789,N_4458);
nor U8220 (N_8220,N_5663,N_4148);
and U8221 (N_8221,N_5886,N_5487);
or U8222 (N_8222,N_5688,N_3858);
nand U8223 (N_8223,N_4224,N_5634);
or U8224 (N_8224,N_3656,N_4446);
nor U8225 (N_8225,N_3707,N_3172);
xnor U8226 (N_8226,N_3092,N_5654);
and U8227 (N_8227,N_5298,N_3438);
nor U8228 (N_8228,N_4732,N_5405);
nand U8229 (N_8229,N_4515,N_5133);
nor U8230 (N_8230,N_3125,N_3872);
nand U8231 (N_8231,N_4190,N_3511);
xnor U8232 (N_8232,N_5921,N_5089);
nor U8233 (N_8233,N_5785,N_4304);
and U8234 (N_8234,N_3341,N_3102);
and U8235 (N_8235,N_4634,N_5780);
nand U8236 (N_8236,N_3086,N_3423);
nor U8237 (N_8237,N_5341,N_4063);
nand U8238 (N_8238,N_3424,N_3320);
nand U8239 (N_8239,N_5510,N_5809);
nand U8240 (N_8240,N_4908,N_5618);
and U8241 (N_8241,N_3512,N_3904);
or U8242 (N_8242,N_4655,N_5288);
or U8243 (N_8243,N_3258,N_5147);
nor U8244 (N_8244,N_4288,N_5580);
and U8245 (N_8245,N_5999,N_4056);
nor U8246 (N_8246,N_5003,N_4904);
nor U8247 (N_8247,N_3301,N_5374);
and U8248 (N_8248,N_5927,N_4053);
and U8249 (N_8249,N_5615,N_5122);
nand U8250 (N_8250,N_4574,N_5459);
and U8251 (N_8251,N_4506,N_4386);
and U8252 (N_8252,N_5112,N_3180);
nand U8253 (N_8253,N_3221,N_4131);
nor U8254 (N_8254,N_4219,N_5819);
nor U8255 (N_8255,N_5474,N_3243);
nor U8256 (N_8256,N_4431,N_4755);
nand U8257 (N_8257,N_4908,N_3911);
nand U8258 (N_8258,N_3057,N_4398);
and U8259 (N_8259,N_4032,N_5195);
and U8260 (N_8260,N_4038,N_3576);
nor U8261 (N_8261,N_3987,N_4481);
nand U8262 (N_8262,N_3724,N_3824);
or U8263 (N_8263,N_3826,N_3675);
nor U8264 (N_8264,N_3460,N_4789);
nand U8265 (N_8265,N_3131,N_5058);
and U8266 (N_8266,N_3731,N_3419);
nand U8267 (N_8267,N_4529,N_4262);
or U8268 (N_8268,N_3316,N_3823);
xor U8269 (N_8269,N_4656,N_4960);
and U8270 (N_8270,N_5636,N_5734);
nor U8271 (N_8271,N_3374,N_3574);
or U8272 (N_8272,N_4288,N_3488);
and U8273 (N_8273,N_4274,N_5099);
or U8274 (N_8274,N_4561,N_4802);
nor U8275 (N_8275,N_5054,N_4948);
and U8276 (N_8276,N_5791,N_4549);
nand U8277 (N_8277,N_5001,N_4690);
nor U8278 (N_8278,N_5357,N_3974);
nor U8279 (N_8279,N_4624,N_4983);
nor U8280 (N_8280,N_3228,N_3904);
and U8281 (N_8281,N_5370,N_3069);
nand U8282 (N_8282,N_3094,N_4424);
nor U8283 (N_8283,N_4024,N_4831);
and U8284 (N_8284,N_4093,N_4189);
nor U8285 (N_8285,N_3114,N_4103);
nor U8286 (N_8286,N_4147,N_5569);
nor U8287 (N_8287,N_3186,N_4408);
nor U8288 (N_8288,N_5472,N_5561);
xnor U8289 (N_8289,N_3006,N_3550);
or U8290 (N_8290,N_4531,N_4532);
and U8291 (N_8291,N_5388,N_4381);
nand U8292 (N_8292,N_5367,N_4553);
and U8293 (N_8293,N_3339,N_4091);
nor U8294 (N_8294,N_3721,N_5463);
nor U8295 (N_8295,N_4038,N_5692);
nand U8296 (N_8296,N_4921,N_5538);
and U8297 (N_8297,N_4254,N_5914);
nor U8298 (N_8298,N_5130,N_3013);
xnor U8299 (N_8299,N_5354,N_4020);
and U8300 (N_8300,N_5738,N_3724);
nand U8301 (N_8301,N_4273,N_4561);
or U8302 (N_8302,N_5237,N_4182);
or U8303 (N_8303,N_4784,N_4752);
nor U8304 (N_8304,N_5979,N_4269);
or U8305 (N_8305,N_3414,N_3993);
and U8306 (N_8306,N_5865,N_4877);
and U8307 (N_8307,N_4400,N_3013);
nor U8308 (N_8308,N_4217,N_5764);
nand U8309 (N_8309,N_4860,N_4622);
xor U8310 (N_8310,N_5328,N_5401);
or U8311 (N_8311,N_3885,N_5931);
xnor U8312 (N_8312,N_4439,N_3884);
or U8313 (N_8313,N_5063,N_5596);
nand U8314 (N_8314,N_5338,N_3901);
or U8315 (N_8315,N_5130,N_5125);
xor U8316 (N_8316,N_4007,N_5059);
nor U8317 (N_8317,N_5502,N_3147);
and U8318 (N_8318,N_5561,N_3727);
nor U8319 (N_8319,N_4489,N_3506);
and U8320 (N_8320,N_3854,N_4732);
xnor U8321 (N_8321,N_5399,N_4927);
nor U8322 (N_8322,N_5457,N_5056);
xor U8323 (N_8323,N_3999,N_3216);
nor U8324 (N_8324,N_3955,N_5595);
nor U8325 (N_8325,N_3010,N_3188);
and U8326 (N_8326,N_5535,N_3911);
or U8327 (N_8327,N_5848,N_4203);
or U8328 (N_8328,N_4542,N_5823);
and U8329 (N_8329,N_4757,N_4482);
nor U8330 (N_8330,N_3584,N_5235);
or U8331 (N_8331,N_5467,N_4207);
and U8332 (N_8332,N_4284,N_3249);
or U8333 (N_8333,N_5355,N_3199);
nand U8334 (N_8334,N_5976,N_4286);
and U8335 (N_8335,N_5729,N_5578);
nand U8336 (N_8336,N_5150,N_5433);
or U8337 (N_8337,N_4487,N_3546);
nor U8338 (N_8338,N_4328,N_5231);
or U8339 (N_8339,N_5938,N_4232);
and U8340 (N_8340,N_5362,N_4097);
and U8341 (N_8341,N_3177,N_5334);
nand U8342 (N_8342,N_3243,N_3638);
xor U8343 (N_8343,N_5578,N_3821);
nand U8344 (N_8344,N_3865,N_4255);
and U8345 (N_8345,N_4261,N_5463);
or U8346 (N_8346,N_5509,N_5698);
or U8347 (N_8347,N_4158,N_4599);
nand U8348 (N_8348,N_5369,N_4250);
or U8349 (N_8349,N_5028,N_4638);
and U8350 (N_8350,N_5894,N_3954);
xor U8351 (N_8351,N_3129,N_3183);
and U8352 (N_8352,N_3672,N_5780);
nor U8353 (N_8353,N_3919,N_4738);
and U8354 (N_8354,N_4613,N_3707);
nand U8355 (N_8355,N_3676,N_5658);
or U8356 (N_8356,N_5021,N_5308);
and U8357 (N_8357,N_3263,N_5654);
nand U8358 (N_8358,N_4806,N_5904);
nor U8359 (N_8359,N_4647,N_5770);
xor U8360 (N_8360,N_5818,N_5120);
or U8361 (N_8361,N_3160,N_4896);
nand U8362 (N_8362,N_5419,N_3603);
nor U8363 (N_8363,N_4860,N_4099);
nor U8364 (N_8364,N_5644,N_3169);
or U8365 (N_8365,N_3650,N_3033);
and U8366 (N_8366,N_3461,N_4158);
nor U8367 (N_8367,N_4222,N_4242);
xor U8368 (N_8368,N_4430,N_5077);
xor U8369 (N_8369,N_5098,N_4908);
or U8370 (N_8370,N_3314,N_5474);
nor U8371 (N_8371,N_5335,N_4105);
and U8372 (N_8372,N_4464,N_3268);
nor U8373 (N_8373,N_3899,N_5811);
nor U8374 (N_8374,N_3212,N_5741);
nand U8375 (N_8375,N_4766,N_4759);
or U8376 (N_8376,N_5368,N_4452);
nor U8377 (N_8377,N_4321,N_5159);
nand U8378 (N_8378,N_4881,N_4867);
nor U8379 (N_8379,N_4559,N_5228);
and U8380 (N_8380,N_3498,N_4386);
or U8381 (N_8381,N_4603,N_5498);
or U8382 (N_8382,N_4956,N_3133);
and U8383 (N_8383,N_3327,N_5257);
nor U8384 (N_8384,N_3280,N_4021);
nand U8385 (N_8385,N_4354,N_3536);
or U8386 (N_8386,N_5981,N_5321);
and U8387 (N_8387,N_3460,N_5767);
and U8388 (N_8388,N_4940,N_4249);
or U8389 (N_8389,N_4128,N_5254);
or U8390 (N_8390,N_3966,N_5728);
and U8391 (N_8391,N_5452,N_3264);
and U8392 (N_8392,N_3239,N_5210);
nand U8393 (N_8393,N_4960,N_3601);
nor U8394 (N_8394,N_5628,N_4426);
nor U8395 (N_8395,N_4082,N_4097);
or U8396 (N_8396,N_3187,N_3035);
xor U8397 (N_8397,N_3688,N_4745);
and U8398 (N_8398,N_4906,N_4366);
xnor U8399 (N_8399,N_4279,N_3548);
nor U8400 (N_8400,N_5290,N_4673);
nor U8401 (N_8401,N_5139,N_3188);
nor U8402 (N_8402,N_4089,N_3357);
and U8403 (N_8403,N_4985,N_3962);
or U8404 (N_8404,N_3685,N_5823);
nor U8405 (N_8405,N_5258,N_4426);
or U8406 (N_8406,N_5037,N_5364);
or U8407 (N_8407,N_5266,N_4799);
and U8408 (N_8408,N_4599,N_5180);
nor U8409 (N_8409,N_5622,N_4795);
nand U8410 (N_8410,N_3234,N_5721);
nor U8411 (N_8411,N_4330,N_4253);
nand U8412 (N_8412,N_5917,N_4100);
xor U8413 (N_8413,N_3455,N_3902);
nor U8414 (N_8414,N_5369,N_4553);
xor U8415 (N_8415,N_3537,N_3687);
and U8416 (N_8416,N_4943,N_4461);
or U8417 (N_8417,N_4575,N_4678);
nand U8418 (N_8418,N_5335,N_4537);
nand U8419 (N_8419,N_4316,N_4026);
nor U8420 (N_8420,N_3119,N_5009);
nor U8421 (N_8421,N_5686,N_4828);
or U8422 (N_8422,N_4771,N_3927);
nor U8423 (N_8423,N_4283,N_4853);
nand U8424 (N_8424,N_5884,N_4984);
and U8425 (N_8425,N_5281,N_5136);
nand U8426 (N_8426,N_4995,N_3221);
or U8427 (N_8427,N_5440,N_5622);
and U8428 (N_8428,N_5413,N_3207);
nor U8429 (N_8429,N_5059,N_3711);
or U8430 (N_8430,N_4798,N_4200);
or U8431 (N_8431,N_4819,N_3750);
nand U8432 (N_8432,N_3325,N_3124);
nor U8433 (N_8433,N_4655,N_4782);
nand U8434 (N_8434,N_5149,N_3404);
and U8435 (N_8435,N_3433,N_3244);
and U8436 (N_8436,N_5220,N_5952);
or U8437 (N_8437,N_4854,N_5800);
or U8438 (N_8438,N_3824,N_3641);
nand U8439 (N_8439,N_4074,N_5739);
nor U8440 (N_8440,N_4150,N_4215);
xor U8441 (N_8441,N_3642,N_4205);
nand U8442 (N_8442,N_3905,N_3534);
nor U8443 (N_8443,N_5852,N_3819);
nor U8444 (N_8444,N_3743,N_4817);
nand U8445 (N_8445,N_5952,N_5554);
nand U8446 (N_8446,N_4831,N_5894);
nand U8447 (N_8447,N_3192,N_3322);
nor U8448 (N_8448,N_3914,N_5469);
or U8449 (N_8449,N_3323,N_5418);
and U8450 (N_8450,N_4045,N_5041);
xnor U8451 (N_8451,N_4429,N_4630);
xor U8452 (N_8452,N_3993,N_3868);
and U8453 (N_8453,N_4372,N_3688);
nand U8454 (N_8454,N_3667,N_5062);
xor U8455 (N_8455,N_5971,N_5970);
nand U8456 (N_8456,N_3193,N_3544);
nand U8457 (N_8457,N_3121,N_3880);
nor U8458 (N_8458,N_4317,N_5292);
xor U8459 (N_8459,N_4097,N_3676);
xor U8460 (N_8460,N_3252,N_5366);
or U8461 (N_8461,N_5091,N_4415);
or U8462 (N_8462,N_3665,N_3836);
xor U8463 (N_8463,N_4889,N_4846);
xnor U8464 (N_8464,N_5121,N_3332);
nor U8465 (N_8465,N_5539,N_3305);
or U8466 (N_8466,N_5191,N_5253);
nand U8467 (N_8467,N_5476,N_4184);
nand U8468 (N_8468,N_4870,N_5667);
or U8469 (N_8469,N_4851,N_4483);
or U8470 (N_8470,N_5265,N_4601);
nor U8471 (N_8471,N_5080,N_3773);
nand U8472 (N_8472,N_3882,N_5793);
xor U8473 (N_8473,N_5565,N_3725);
and U8474 (N_8474,N_5737,N_3038);
nand U8475 (N_8475,N_3026,N_4148);
nor U8476 (N_8476,N_4576,N_3681);
nor U8477 (N_8477,N_4909,N_3828);
or U8478 (N_8478,N_3197,N_5348);
nand U8479 (N_8479,N_5914,N_4710);
nor U8480 (N_8480,N_5332,N_3683);
or U8481 (N_8481,N_4570,N_4299);
nand U8482 (N_8482,N_3211,N_4896);
or U8483 (N_8483,N_3439,N_4484);
nand U8484 (N_8484,N_5417,N_5942);
nand U8485 (N_8485,N_5309,N_5767);
and U8486 (N_8486,N_5871,N_5726);
nor U8487 (N_8487,N_3853,N_5468);
or U8488 (N_8488,N_4617,N_4603);
or U8489 (N_8489,N_4063,N_5994);
or U8490 (N_8490,N_3412,N_4311);
nor U8491 (N_8491,N_3710,N_5159);
and U8492 (N_8492,N_4384,N_3593);
nor U8493 (N_8493,N_5141,N_3260);
or U8494 (N_8494,N_3592,N_4122);
xor U8495 (N_8495,N_3350,N_4518);
and U8496 (N_8496,N_3878,N_3037);
or U8497 (N_8497,N_4772,N_3935);
nor U8498 (N_8498,N_4897,N_5316);
and U8499 (N_8499,N_4495,N_5328);
nor U8500 (N_8500,N_4869,N_4851);
or U8501 (N_8501,N_5366,N_3913);
nor U8502 (N_8502,N_5047,N_5038);
or U8503 (N_8503,N_5871,N_4805);
nand U8504 (N_8504,N_3586,N_3444);
or U8505 (N_8505,N_3821,N_5083);
or U8506 (N_8506,N_5337,N_4567);
and U8507 (N_8507,N_3970,N_4206);
or U8508 (N_8508,N_3766,N_3708);
nand U8509 (N_8509,N_4315,N_3958);
nand U8510 (N_8510,N_3567,N_3539);
nor U8511 (N_8511,N_5143,N_5765);
and U8512 (N_8512,N_3367,N_5463);
or U8513 (N_8513,N_3845,N_4872);
and U8514 (N_8514,N_4924,N_3588);
and U8515 (N_8515,N_4330,N_4123);
and U8516 (N_8516,N_3649,N_3963);
nand U8517 (N_8517,N_4846,N_4274);
or U8518 (N_8518,N_5198,N_4952);
or U8519 (N_8519,N_4410,N_4697);
nor U8520 (N_8520,N_4486,N_3537);
nand U8521 (N_8521,N_4288,N_5792);
xnor U8522 (N_8522,N_4015,N_3789);
or U8523 (N_8523,N_3389,N_4614);
nor U8524 (N_8524,N_4734,N_3572);
and U8525 (N_8525,N_4605,N_5474);
or U8526 (N_8526,N_5363,N_4652);
and U8527 (N_8527,N_3631,N_3105);
nor U8528 (N_8528,N_3550,N_5749);
xor U8529 (N_8529,N_3496,N_3222);
or U8530 (N_8530,N_3667,N_3345);
or U8531 (N_8531,N_4202,N_5145);
nor U8532 (N_8532,N_5317,N_3516);
nand U8533 (N_8533,N_3009,N_4545);
nor U8534 (N_8534,N_4575,N_4093);
or U8535 (N_8535,N_5234,N_5850);
or U8536 (N_8536,N_4304,N_5236);
and U8537 (N_8537,N_5257,N_4937);
or U8538 (N_8538,N_3490,N_3997);
nand U8539 (N_8539,N_5046,N_5189);
or U8540 (N_8540,N_4756,N_4296);
xnor U8541 (N_8541,N_3463,N_5324);
nor U8542 (N_8542,N_3946,N_3374);
nand U8543 (N_8543,N_5982,N_5728);
nand U8544 (N_8544,N_5544,N_4834);
or U8545 (N_8545,N_3191,N_5537);
or U8546 (N_8546,N_3342,N_5123);
nor U8547 (N_8547,N_5573,N_5375);
nor U8548 (N_8548,N_3833,N_3391);
or U8549 (N_8549,N_4313,N_4810);
or U8550 (N_8550,N_5834,N_3708);
or U8551 (N_8551,N_3646,N_4401);
or U8552 (N_8552,N_5526,N_3751);
nor U8553 (N_8553,N_3534,N_3701);
or U8554 (N_8554,N_4999,N_5007);
nor U8555 (N_8555,N_4388,N_4758);
or U8556 (N_8556,N_5399,N_5527);
nor U8557 (N_8557,N_3020,N_5148);
nor U8558 (N_8558,N_3003,N_4967);
nor U8559 (N_8559,N_3052,N_3179);
and U8560 (N_8560,N_3363,N_5805);
nand U8561 (N_8561,N_5200,N_5864);
xor U8562 (N_8562,N_4441,N_4781);
xor U8563 (N_8563,N_4572,N_3577);
and U8564 (N_8564,N_3275,N_3851);
xnor U8565 (N_8565,N_5376,N_4839);
and U8566 (N_8566,N_4096,N_4373);
or U8567 (N_8567,N_4343,N_5921);
or U8568 (N_8568,N_4030,N_4779);
nand U8569 (N_8569,N_5736,N_5898);
or U8570 (N_8570,N_3882,N_3480);
or U8571 (N_8571,N_5410,N_5537);
nand U8572 (N_8572,N_4905,N_3142);
or U8573 (N_8573,N_4993,N_4250);
nor U8574 (N_8574,N_4764,N_5955);
or U8575 (N_8575,N_5610,N_3452);
or U8576 (N_8576,N_4852,N_5884);
nor U8577 (N_8577,N_3001,N_5172);
and U8578 (N_8578,N_5624,N_5177);
or U8579 (N_8579,N_3228,N_3427);
nand U8580 (N_8580,N_5109,N_4556);
nand U8581 (N_8581,N_5265,N_4213);
or U8582 (N_8582,N_4845,N_4338);
or U8583 (N_8583,N_4996,N_5085);
or U8584 (N_8584,N_4782,N_3625);
xnor U8585 (N_8585,N_4661,N_3074);
or U8586 (N_8586,N_4936,N_4200);
nor U8587 (N_8587,N_4104,N_5902);
nor U8588 (N_8588,N_5050,N_4852);
or U8589 (N_8589,N_5767,N_5429);
or U8590 (N_8590,N_4282,N_3664);
xnor U8591 (N_8591,N_5271,N_4655);
and U8592 (N_8592,N_5923,N_3539);
nand U8593 (N_8593,N_4473,N_5568);
and U8594 (N_8594,N_3285,N_3832);
nand U8595 (N_8595,N_4070,N_5887);
nor U8596 (N_8596,N_5845,N_3296);
and U8597 (N_8597,N_3712,N_5307);
and U8598 (N_8598,N_3364,N_4580);
nor U8599 (N_8599,N_5754,N_4339);
nor U8600 (N_8600,N_3153,N_4940);
or U8601 (N_8601,N_4540,N_4886);
nor U8602 (N_8602,N_4528,N_5023);
and U8603 (N_8603,N_3564,N_3646);
or U8604 (N_8604,N_4528,N_3207);
nor U8605 (N_8605,N_5687,N_5803);
nor U8606 (N_8606,N_3838,N_5265);
nand U8607 (N_8607,N_5650,N_5900);
nand U8608 (N_8608,N_5847,N_3552);
xnor U8609 (N_8609,N_4540,N_5870);
nor U8610 (N_8610,N_3089,N_4331);
or U8611 (N_8611,N_3020,N_5984);
nor U8612 (N_8612,N_4925,N_3530);
nor U8613 (N_8613,N_3252,N_5734);
nor U8614 (N_8614,N_4927,N_5225);
nand U8615 (N_8615,N_5220,N_5473);
and U8616 (N_8616,N_5854,N_5859);
or U8617 (N_8617,N_5876,N_4365);
nor U8618 (N_8618,N_5002,N_3381);
xnor U8619 (N_8619,N_3467,N_3343);
and U8620 (N_8620,N_3142,N_4505);
or U8621 (N_8621,N_4414,N_3252);
or U8622 (N_8622,N_5380,N_3397);
nand U8623 (N_8623,N_3181,N_4404);
or U8624 (N_8624,N_4085,N_3997);
nand U8625 (N_8625,N_3319,N_3794);
xnor U8626 (N_8626,N_5384,N_4630);
nand U8627 (N_8627,N_5815,N_5881);
and U8628 (N_8628,N_5673,N_5854);
and U8629 (N_8629,N_3034,N_4761);
nand U8630 (N_8630,N_5302,N_5697);
nand U8631 (N_8631,N_3246,N_5954);
or U8632 (N_8632,N_4343,N_3510);
nand U8633 (N_8633,N_4539,N_4178);
nand U8634 (N_8634,N_5508,N_3044);
or U8635 (N_8635,N_4322,N_4677);
nand U8636 (N_8636,N_5499,N_3226);
nand U8637 (N_8637,N_5487,N_3712);
or U8638 (N_8638,N_4909,N_5132);
or U8639 (N_8639,N_3642,N_4370);
nor U8640 (N_8640,N_5164,N_3162);
and U8641 (N_8641,N_3304,N_5781);
or U8642 (N_8642,N_4084,N_5991);
nor U8643 (N_8643,N_3357,N_5915);
nand U8644 (N_8644,N_5778,N_5671);
or U8645 (N_8645,N_3307,N_5613);
nor U8646 (N_8646,N_3887,N_3976);
and U8647 (N_8647,N_5400,N_5944);
nor U8648 (N_8648,N_4862,N_4564);
nand U8649 (N_8649,N_4598,N_3677);
or U8650 (N_8650,N_3406,N_3056);
nand U8651 (N_8651,N_3700,N_3607);
nand U8652 (N_8652,N_5501,N_3413);
xnor U8653 (N_8653,N_4078,N_4359);
nand U8654 (N_8654,N_4488,N_3664);
nand U8655 (N_8655,N_3573,N_3622);
or U8656 (N_8656,N_3086,N_5659);
or U8657 (N_8657,N_5713,N_5442);
nor U8658 (N_8658,N_4211,N_4578);
and U8659 (N_8659,N_4227,N_4656);
or U8660 (N_8660,N_4439,N_5551);
and U8661 (N_8661,N_4007,N_5776);
or U8662 (N_8662,N_4005,N_4540);
nor U8663 (N_8663,N_5047,N_5894);
nand U8664 (N_8664,N_3058,N_5034);
and U8665 (N_8665,N_4762,N_3730);
and U8666 (N_8666,N_4806,N_4720);
or U8667 (N_8667,N_4005,N_4346);
and U8668 (N_8668,N_3243,N_4055);
nor U8669 (N_8669,N_5360,N_3345);
or U8670 (N_8670,N_4588,N_4436);
and U8671 (N_8671,N_3512,N_5016);
nor U8672 (N_8672,N_4248,N_4796);
nor U8673 (N_8673,N_5816,N_5021);
or U8674 (N_8674,N_3863,N_5933);
nand U8675 (N_8675,N_4522,N_5328);
or U8676 (N_8676,N_3812,N_5298);
xnor U8677 (N_8677,N_5110,N_4498);
and U8678 (N_8678,N_4269,N_4307);
nand U8679 (N_8679,N_3692,N_5666);
and U8680 (N_8680,N_5984,N_3810);
and U8681 (N_8681,N_3452,N_5677);
nor U8682 (N_8682,N_4565,N_4998);
nand U8683 (N_8683,N_3162,N_4462);
or U8684 (N_8684,N_3578,N_4184);
or U8685 (N_8685,N_3364,N_3504);
nand U8686 (N_8686,N_4306,N_4159);
or U8687 (N_8687,N_3057,N_4284);
and U8688 (N_8688,N_4989,N_3620);
nand U8689 (N_8689,N_5878,N_4317);
nor U8690 (N_8690,N_3699,N_3217);
or U8691 (N_8691,N_3920,N_5817);
and U8692 (N_8692,N_4312,N_5030);
nor U8693 (N_8693,N_5055,N_3555);
nor U8694 (N_8694,N_3721,N_3294);
and U8695 (N_8695,N_5049,N_3922);
and U8696 (N_8696,N_3112,N_3194);
or U8697 (N_8697,N_5405,N_4199);
nand U8698 (N_8698,N_3842,N_3912);
nor U8699 (N_8699,N_4245,N_5279);
and U8700 (N_8700,N_4754,N_5871);
and U8701 (N_8701,N_5377,N_5864);
nor U8702 (N_8702,N_5817,N_3917);
nor U8703 (N_8703,N_3086,N_3592);
or U8704 (N_8704,N_3642,N_3868);
nor U8705 (N_8705,N_5573,N_3489);
nor U8706 (N_8706,N_5785,N_4589);
nand U8707 (N_8707,N_3071,N_4349);
nand U8708 (N_8708,N_3174,N_5818);
and U8709 (N_8709,N_4264,N_5166);
or U8710 (N_8710,N_5065,N_5102);
and U8711 (N_8711,N_4285,N_5094);
nor U8712 (N_8712,N_3312,N_3220);
nor U8713 (N_8713,N_5070,N_4808);
nor U8714 (N_8714,N_4223,N_3103);
or U8715 (N_8715,N_5991,N_5772);
and U8716 (N_8716,N_4475,N_3279);
or U8717 (N_8717,N_3201,N_5842);
and U8718 (N_8718,N_3910,N_3846);
and U8719 (N_8719,N_3696,N_4681);
nor U8720 (N_8720,N_4409,N_5903);
nand U8721 (N_8721,N_3251,N_3012);
nor U8722 (N_8722,N_4273,N_3842);
nand U8723 (N_8723,N_4121,N_5611);
or U8724 (N_8724,N_5968,N_4214);
nor U8725 (N_8725,N_5907,N_5477);
or U8726 (N_8726,N_5622,N_5666);
nand U8727 (N_8727,N_4410,N_3954);
or U8728 (N_8728,N_4340,N_4869);
nand U8729 (N_8729,N_3841,N_5909);
nor U8730 (N_8730,N_5113,N_4032);
nand U8731 (N_8731,N_5484,N_5594);
nand U8732 (N_8732,N_5163,N_3554);
and U8733 (N_8733,N_3374,N_4455);
nor U8734 (N_8734,N_4367,N_3630);
nand U8735 (N_8735,N_4043,N_5963);
nand U8736 (N_8736,N_4107,N_5894);
xnor U8737 (N_8737,N_3758,N_4981);
nand U8738 (N_8738,N_5943,N_4689);
nand U8739 (N_8739,N_4489,N_5984);
xnor U8740 (N_8740,N_5696,N_3193);
nor U8741 (N_8741,N_3389,N_5196);
nand U8742 (N_8742,N_3125,N_5474);
or U8743 (N_8743,N_5373,N_5718);
nand U8744 (N_8744,N_5546,N_5894);
and U8745 (N_8745,N_4245,N_5755);
and U8746 (N_8746,N_5544,N_5017);
or U8747 (N_8747,N_4364,N_5166);
or U8748 (N_8748,N_3901,N_4561);
and U8749 (N_8749,N_4268,N_4957);
and U8750 (N_8750,N_3964,N_3903);
or U8751 (N_8751,N_5626,N_3273);
nor U8752 (N_8752,N_4852,N_5225);
nand U8753 (N_8753,N_5176,N_4354);
or U8754 (N_8754,N_4419,N_3646);
or U8755 (N_8755,N_5644,N_5615);
nand U8756 (N_8756,N_3819,N_4016);
nand U8757 (N_8757,N_4448,N_3114);
or U8758 (N_8758,N_4536,N_3492);
nor U8759 (N_8759,N_5991,N_5402);
nor U8760 (N_8760,N_4451,N_4606);
xnor U8761 (N_8761,N_5775,N_5767);
nand U8762 (N_8762,N_3744,N_4911);
or U8763 (N_8763,N_5119,N_4257);
nand U8764 (N_8764,N_3935,N_3865);
and U8765 (N_8765,N_4609,N_4226);
and U8766 (N_8766,N_3160,N_5280);
and U8767 (N_8767,N_4720,N_5294);
or U8768 (N_8768,N_4680,N_3056);
and U8769 (N_8769,N_3590,N_4480);
and U8770 (N_8770,N_3292,N_4324);
or U8771 (N_8771,N_4827,N_5868);
nor U8772 (N_8772,N_5512,N_5585);
nor U8773 (N_8773,N_5740,N_4558);
nor U8774 (N_8774,N_3334,N_4108);
nand U8775 (N_8775,N_5725,N_3716);
nor U8776 (N_8776,N_3924,N_4993);
nand U8777 (N_8777,N_3573,N_5128);
or U8778 (N_8778,N_5996,N_4841);
nand U8779 (N_8779,N_3587,N_5700);
xor U8780 (N_8780,N_4488,N_4399);
and U8781 (N_8781,N_5116,N_5404);
or U8782 (N_8782,N_5687,N_5428);
xor U8783 (N_8783,N_5549,N_4336);
xnor U8784 (N_8784,N_4507,N_4989);
nor U8785 (N_8785,N_3525,N_4872);
nand U8786 (N_8786,N_3178,N_3437);
and U8787 (N_8787,N_4555,N_4019);
xor U8788 (N_8788,N_4836,N_3948);
xor U8789 (N_8789,N_3070,N_4341);
nand U8790 (N_8790,N_4658,N_4503);
or U8791 (N_8791,N_4562,N_3430);
or U8792 (N_8792,N_4928,N_5566);
nand U8793 (N_8793,N_5304,N_3444);
or U8794 (N_8794,N_4547,N_4001);
or U8795 (N_8795,N_4002,N_5854);
and U8796 (N_8796,N_3308,N_5978);
or U8797 (N_8797,N_3440,N_3026);
nor U8798 (N_8798,N_4452,N_3830);
nor U8799 (N_8799,N_3915,N_4361);
or U8800 (N_8800,N_4469,N_3877);
nand U8801 (N_8801,N_5390,N_4551);
xor U8802 (N_8802,N_4616,N_4502);
and U8803 (N_8803,N_3254,N_3894);
or U8804 (N_8804,N_4255,N_5898);
or U8805 (N_8805,N_3277,N_4015);
nand U8806 (N_8806,N_5118,N_3194);
nand U8807 (N_8807,N_5511,N_5345);
nor U8808 (N_8808,N_5295,N_5371);
or U8809 (N_8809,N_5805,N_4114);
xnor U8810 (N_8810,N_5863,N_4085);
nand U8811 (N_8811,N_4685,N_3935);
or U8812 (N_8812,N_4250,N_4317);
nor U8813 (N_8813,N_4921,N_5359);
xor U8814 (N_8814,N_5645,N_3915);
or U8815 (N_8815,N_3319,N_5921);
nor U8816 (N_8816,N_3056,N_5489);
nand U8817 (N_8817,N_3168,N_5821);
nand U8818 (N_8818,N_4941,N_5604);
and U8819 (N_8819,N_4005,N_5042);
nor U8820 (N_8820,N_3073,N_5177);
xnor U8821 (N_8821,N_5827,N_5477);
or U8822 (N_8822,N_4841,N_4295);
or U8823 (N_8823,N_5290,N_5185);
nor U8824 (N_8824,N_3764,N_3676);
or U8825 (N_8825,N_5458,N_3252);
nor U8826 (N_8826,N_4829,N_4871);
xnor U8827 (N_8827,N_5075,N_4781);
and U8828 (N_8828,N_5416,N_4546);
or U8829 (N_8829,N_4135,N_4652);
or U8830 (N_8830,N_5832,N_3090);
xor U8831 (N_8831,N_4291,N_4723);
and U8832 (N_8832,N_3988,N_3165);
nand U8833 (N_8833,N_5535,N_5303);
nand U8834 (N_8834,N_3663,N_5833);
nand U8835 (N_8835,N_4603,N_4567);
nand U8836 (N_8836,N_3915,N_3145);
and U8837 (N_8837,N_3465,N_4994);
xor U8838 (N_8838,N_3795,N_5945);
and U8839 (N_8839,N_4586,N_3066);
xnor U8840 (N_8840,N_5039,N_3751);
or U8841 (N_8841,N_5225,N_4378);
nand U8842 (N_8842,N_3355,N_4597);
nor U8843 (N_8843,N_4690,N_3711);
nand U8844 (N_8844,N_3787,N_4052);
or U8845 (N_8845,N_4677,N_5988);
or U8846 (N_8846,N_4019,N_5278);
nand U8847 (N_8847,N_3677,N_3474);
nand U8848 (N_8848,N_3860,N_4355);
nor U8849 (N_8849,N_5125,N_4949);
or U8850 (N_8850,N_5353,N_3990);
and U8851 (N_8851,N_3229,N_4636);
and U8852 (N_8852,N_3354,N_3489);
and U8853 (N_8853,N_3099,N_3603);
nand U8854 (N_8854,N_5405,N_4386);
and U8855 (N_8855,N_3141,N_4455);
nor U8856 (N_8856,N_3325,N_3383);
or U8857 (N_8857,N_5314,N_4086);
nor U8858 (N_8858,N_3978,N_5077);
or U8859 (N_8859,N_3045,N_4856);
and U8860 (N_8860,N_4774,N_4433);
and U8861 (N_8861,N_4542,N_4998);
xor U8862 (N_8862,N_4982,N_5208);
xnor U8863 (N_8863,N_4786,N_4209);
and U8864 (N_8864,N_5381,N_5140);
nand U8865 (N_8865,N_5378,N_4709);
xnor U8866 (N_8866,N_3495,N_5077);
and U8867 (N_8867,N_3177,N_5802);
or U8868 (N_8868,N_3445,N_4505);
nand U8869 (N_8869,N_5911,N_4276);
and U8870 (N_8870,N_4742,N_5152);
or U8871 (N_8871,N_3704,N_3267);
nor U8872 (N_8872,N_5199,N_3131);
nor U8873 (N_8873,N_5973,N_3786);
and U8874 (N_8874,N_4279,N_3885);
nand U8875 (N_8875,N_3004,N_5160);
or U8876 (N_8876,N_4908,N_4274);
nand U8877 (N_8877,N_5121,N_5688);
nor U8878 (N_8878,N_3462,N_5582);
nor U8879 (N_8879,N_5394,N_5767);
nor U8880 (N_8880,N_5002,N_5712);
or U8881 (N_8881,N_5700,N_4663);
nor U8882 (N_8882,N_5770,N_5427);
nor U8883 (N_8883,N_4454,N_3689);
nor U8884 (N_8884,N_5091,N_3861);
nor U8885 (N_8885,N_3748,N_5008);
nor U8886 (N_8886,N_3871,N_5153);
xor U8887 (N_8887,N_4589,N_5744);
and U8888 (N_8888,N_4548,N_5606);
or U8889 (N_8889,N_3034,N_3363);
or U8890 (N_8890,N_5073,N_4924);
and U8891 (N_8891,N_3337,N_5499);
nor U8892 (N_8892,N_3031,N_5461);
or U8893 (N_8893,N_5914,N_4796);
and U8894 (N_8894,N_3731,N_3763);
or U8895 (N_8895,N_5528,N_3261);
or U8896 (N_8896,N_4760,N_4432);
or U8897 (N_8897,N_3532,N_4652);
nand U8898 (N_8898,N_4980,N_5225);
nand U8899 (N_8899,N_5191,N_3610);
and U8900 (N_8900,N_3898,N_5288);
or U8901 (N_8901,N_3923,N_4040);
nand U8902 (N_8902,N_3985,N_5443);
nand U8903 (N_8903,N_4957,N_4373);
nor U8904 (N_8904,N_4118,N_4228);
nor U8905 (N_8905,N_3615,N_5360);
nand U8906 (N_8906,N_3349,N_3898);
or U8907 (N_8907,N_3943,N_5567);
nor U8908 (N_8908,N_4094,N_3972);
nand U8909 (N_8909,N_5636,N_3016);
or U8910 (N_8910,N_4312,N_4212);
or U8911 (N_8911,N_3749,N_4696);
nor U8912 (N_8912,N_3812,N_4928);
nor U8913 (N_8913,N_5663,N_5907);
nor U8914 (N_8914,N_4077,N_5597);
nand U8915 (N_8915,N_4851,N_4760);
nor U8916 (N_8916,N_4813,N_5466);
nand U8917 (N_8917,N_5613,N_4816);
or U8918 (N_8918,N_3204,N_5814);
nand U8919 (N_8919,N_3785,N_3920);
or U8920 (N_8920,N_5382,N_5173);
and U8921 (N_8921,N_3246,N_4379);
or U8922 (N_8922,N_3798,N_4993);
and U8923 (N_8923,N_5434,N_4831);
or U8924 (N_8924,N_4079,N_4935);
and U8925 (N_8925,N_5282,N_3149);
or U8926 (N_8926,N_4251,N_3435);
nor U8927 (N_8927,N_4814,N_3829);
nand U8928 (N_8928,N_5240,N_3540);
or U8929 (N_8929,N_5697,N_4047);
xor U8930 (N_8930,N_4734,N_5822);
and U8931 (N_8931,N_5665,N_5833);
nor U8932 (N_8932,N_3160,N_3340);
and U8933 (N_8933,N_4979,N_3252);
nor U8934 (N_8934,N_3350,N_5688);
and U8935 (N_8935,N_5095,N_3384);
nand U8936 (N_8936,N_3313,N_5399);
xor U8937 (N_8937,N_3448,N_3643);
nand U8938 (N_8938,N_4240,N_4124);
or U8939 (N_8939,N_3980,N_4712);
xor U8940 (N_8940,N_4027,N_5336);
or U8941 (N_8941,N_5967,N_4296);
and U8942 (N_8942,N_3013,N_5713);
or U8943 (N_8943,N_5054,N_3567);
nand U8944 (N_8944,N_4902,N_3280);
xor U8945 (N_8945,N_4889,N_5568);
xor U8946 (N_8946,N_4972,N_3699);
nand U8947 (N_8947,N_3904,N_5517);
nor U8948 (N_8948,N_4270,N_4129);
and U8949 (N_8949,N_3923,N_5234);
or U8950 (N_8950,N_3670,N_4644);
and U8951 (N_8951,N_5712,N_5229);
and U8952 (N_8952,N_3664,N_4825);
xnor U8953 (N_8953,N_3135,N_3561);
or U8954 (N_8954,N_4722,N_5133);
nand U8955 (N_8955,N_3737,N_3404);
nand U8956 (N_8956,N_4697,N_5272);
nor U8957 (N_8957,N_4699,N_3892);
nand U8958 (N_8958,N_3444,N_3408);
nor U8959 (N_8959,N_5397,N_5547);
or U8960 (N_8960,N_3588,N_3065);
and U8961 (N_8961,N_3293,N_4621);
and U8962 (N_8962,N_4488,N_5022);
or U8963 (N_8963,N_5063,N_3529);
nor U8964 (N_8964,N_5579,N_5058);
xnor U8965 (N_8965,N_5597,N_4096);
and U8966 (N_8966,N_4483,N_5093);
xnor U8967 (N_8967,N_5295,N_5791);
and U8968 (N_8968,N_5090,N_3014);
and U8969 (N_8969,N_5139,N_3201);
and U8970 (N_8970,N_4407,N_3677);
or U8971 (N_8971,N_5108,N_3820);
and U8972 (N_8972,N_4785,N_4708);
nor U8973 (N_8973,N_3952,N_5926);
nand U8974 (N_8974,N_3560,N_4462);
and U8975 (N_8975,N_4361,N_3910);
and U8976 (N_8976,N_5218,N_5309);
xor U8977 (N_8977,N_3425,N_3655);
nor U8978 (N_8978,N_3909,N_4979);
nand U8979 (N_8979,N_3393,N_5540);
or U8980 (N_8980,N_3199,N_5801);
or U8981 (N_8981,N_3085,N_3695);
xor U8982 (N_8982,N_4899,N_5734);
and U8983 (N_8983,N_4441,N_3831);
nand U8984 (N_8984,N_4919,N_5371);
or U8985 (N_8985,N_3794,N_3172);
nor U8986 (N_8986,N_3441,N_3424);
or U8987 (N_8987,N_3482,N_4096);
and U8988 (N_8988,N_4707,N_5235);
and U8989 (N_8989,N_3970,N_3871);
xnor U8990 (N_8990,N_3671,N_5346);
and U8991 (N_8991,N_5265,N_3491);
or U8992 (N_8992,N_4582,N_3189);
or U8993 (N_8993,N_4011,N_5698);
or U8994 (N_8994,N_5338,N_3817);
nand U8995 (N_8995,N_3528,N_4919);
nand U8996 (N_8996,N_5896,N_3216);
and U8997 (N_8997,N_5209,N_4030);
nor U8998 (N_8998,N_4795,N_4529);
nor U8999 (N_8999,N_3866,N_4559);
xor U9000 (N_9000,N_7855,N_7770);
nand U9001 (N_9001,N_6440,N_8471);
nand U9002 (N_9002,N_6303,N_6038);
and U9003 (N_9003,N_6132,N_6137);
nor U9004 (N_9004,N_8050,N_7663);
nor U9005 (N_9005,N_7686,N_7043);
or U9006 (N_9006,N_6689,N_6408);
xor U9007 (N_9007,N_6133,N_8747);
nand U9008 (N_9008,N_7846,N_7916);
nand U9009 (N_9009,N_7774,N_8122);
or U9010 (N_9010,N_8757,N_8054);
nor U9011 (N_9011,N_7531,N_7370);
or U9012 (N_9012,N_6094,N_6631);
nand U9013 (N_9013,N_6144,N_7077);
nor U9014 (N_9014,N_6876,N_8586);
xor U9015 (N_9015,N_6035,N_7853);
or U9016 (N_9016,N_7803,N_8609);
and U9017 (N_9017,N_6007,N_6648);
and U9018 (N_9018,N_6154,N_8269);
or U9019 (N_9019,N_6048,N_6237);
nor U9020 (N_9020,N_8049,N_6432);
nor U9021 (N_9021,N_6337,N_8933);
nor U9022 (N_9022,N_6256,N_7342);
nor U9023 (N_9023,N_7752,N_8378);
and U9024 (N_9024,N_8475,N_8692);
nand U9025 (N_9025,N_6578,N_8233);
or U9026 (N_9026,N_7259,N_6388);
xor U9027 (N_9027,N_8555,N_8034);
xnor U9028 (N_9028,N_8625,N_6386);
or U9029 (N_9029,N_8683,N_6488);
or U9030 (N_9030,N_7690,N_8336);
nor U9031 (N_9031,N_8558,N_7542);
and U9032 (N_9032,N_8077,N_7859);
nor U9033 (N_9033,N_6314,N_6370);
and U9034 (N_9034,N_6204,N_7823);
nor U9035 (N_9035,N_8003,N_8395);
and U9036 (N_9036,N_6188,N_7233);
and U9037 (N_9037,N_7502,N_8789);
or U9038 (N_9038,N_6981,N_7664);
and U9039 (N_9039,N_8944,N_6528);
or U9040 (N_9040,N_8962,N_6008);
or U9041 (N_9041,N_7061,N_8121);
or U9042 (N_9042,N_7889,N_6289);
or U9043 (N_9043,N_7114,N_7813);
or U9044 (N_9044,N_6243,N_6866);
nand U9045 (N_9045,N_7634,N_7909);
nor U9046 (N_9046,N_7503,N_7602);
nand U9047 (N_9047,N_6124,N_7742);
nor U9048 (N_9048,N_8826,N_7331);
or U9049 (N_9049,N_7751,N_8498);
nor U9050 (N_9050,N_6086,N_8744);
and U9051 (N_9051,N_7518,N_7618);
and U9052 (N_9052,N_6993,N_8549);
xor U9053 (N_9053,N_6533,N_6619);
and U9054 (N_9054,N_7661,N_7279);
xor U9055 (N_9055,N_7829,N_6477);
or U9056 (N_9056,N_7950,N_8118);
xor U9057 (N_9057,N_8303,N_8946);
and U9058 (N_9058,N_8705,N_7601);
or U9059 (N_9059,N_8571,N_6496);
nand U9060 (N_9060,N_8527,N_7949);
nor U9061 (N_9061,N_8102,N_6463);
nand U9062 (N_9062,N_8439,N_8635);
or U9063 (N_9063,N_8848,N_6255);
and U9064 (N_9064,N_8063,N_7764);
nand U9065 (N_9065,N_8566,N_8353);
nand U9066 (N_9066,N_8853,N_7595);
nor U9067 (N_9067,N_7217,N_8324);
and U9068 (N_9068,N_6910,N_6711);
nand U9069 (N_9069,N_6239,N_7364);
nor U9070 (N_9070,N_6942,N_8004);
nor U9071 (N_9071,N_7492,N_8682);
nand U9072 (N_9072,N_6655,N_6581);
nand U9073 (N_9073,N_7730,N_8772);
or U9074 (N_9074,N_6653,N_6174);
and U9075 (N_9075,N_8365,N_7188);
or U9076 (N_9076,N_8093,N_8312);
nand U9077 (N_9077,N_7934,N_8714);
nand U9078 (N_9078,N_8074,N_6976);
xor U9079 (N_9079,N_7013,N_8988);
nand U9080 (N_9080,N_6286,N_7867);
xnor U9081 (N_9081,N_8942,N_7406);
nand U9082 (N_9082,N_7184,N_8229);
nor U9083 (N_9083,N_7510,N_6309);
nor U9084 (N_9084,N_6085,N_7347);
nor U9085 (N_9085,N_7472,N_8218);
or U9086 (N_9086,N_7287,N_7306);
and U9087 (N_9087,N_7359,N_7558);
nor U9088 (N_9088,N_8977,N_7588);
nor U9089 (N_9089,N_7957,N_7945);
nor U9090 (N_9090,N_8238,N_6629);
nand U9091 (N_9091,N_6089,N_8443);
and U9092 (N_9092,N_7373,N_6394);
and U9093 (N_9093,N_8830,N_8822);
nor U9094 (N_9094,N_7267,N_6671);
and U9095 (N_9095,N_7509,N_8978);
or U9096 (N_9096,N_8281,N_6425);
xor U9097 (N_9097,N_7850,N_7155);
or U9098 (N_9098,N_6051,N_6898);
nor U9099 (N_9099,N_7317,N_7799);
or U9100 (N_9100,N_8448,N_8051);
nor U9101 (N_9101,N_6078,N_8882);
and U9102 (N_9102,N_7170,N_7394);
or U9103 (N_9103,N_8748,N_6893);
nor U9104 (N_9104,N_6104,N_7562);
xnor U9105 (N_9105,N_8645,N_8596);
nand U9106 (N_9106,N_6067,N_7225);
or U9107 (N_9107,N_8517,N_6766);
and U9108 (N_9108,N_7203,N_6379);
or U9109 (N_9109,N_7231,N_8456);
or U9110 (N_9110,N_7811,N_8831);
nand U9111 (N_9111,N_7091,N_6932);
xnor U9112 (N_9112,N_7513,N_6906);
xnor U9113 (N_9113,N_8937,N_8394);
nand U9114 (N_9114,N_7655,N_8360);
nand U9115 (N_9115,N_7200,N_6355);
and U9116 (N_9116,N_6374,N_7736);
nand U9117 (N_9117,N_8686,N_8184);
or U9118 (N_9118,N_8215,N_6880);
nand U9119 (N_9119,N_6517,N_7837);
xor U9120 (N_9120,N_8026,N_6472);
nand U9121 (N_9121,N_6826,N_8594);
and U9122 (N_9122,N_7658,N_8078);
xnor U9123 (N_9123,N_8923,N_8357);
nand U9124 (N_9124,N_8342,N_6343);
nor U9125 (N_9125,N_7603,N_7870);
or U9126 (N_9126,N_7360,N_8334);
or U9127 (N_9127,N_6665,N_7218);
nor U9128 (N_9128,N_6846,N_7988);
and U9129 (N_9129,N_7694,N_6501);
xor U9130 (N_9130,N_8907,N_8311);
or U9131 (N_9131,N_8987,N_7440);
and U9132 (N_9132,N_8773,N_7906);
or U9133 (N_9133,N_6963,N_7754);
xnor U9134 (N_9134,N_7534,N_6298);
nor U9135 (N_9135,N_6187,N_6365);
and U9136 (N_9136,N_8158,N_7809);
xnor U9137 (N_9137,N_7550,N_6877);
nor U9138 (N_9138,N_7103,N_8719);
xor U9139 (N_9139,N_7180,N_7260);
nand U9140 (N_9140,N_7275,N_8096);
and U9141 (N_9141,N_8701,N_7461);
nand U9142 (N_9142,N_6173,N_7648);
and U9143 (N_9143,N_7445,N_7428);
xnor U9144 (N_9144,N_8217,N_6565);
or U9145 (N_9145,N_8182,N_6372);
and U9146 (N_9146,N_6505,N_6352);
nand U9147 (N_9147,N_7740,N_8029);
or U9148 (N_9148,N_8043,N_7256);
or U9149 (N_9149,N_6946,N_6034);
and U9150 (N_9150,N_7639,N_7289);
and U9151 (N_9151,N_6869,N_7147);
or U9152 (N_9152,N_7997,N_7755);
or U9153 (N_9153,N_6972,N_6192);
nand U9154 (N_9154,N_7483,N_7580);
or U9155 (N_9155,N_7327,N_8011);
xnor U9156 (N_9156,N_8842,N_8825);
nand U9157 (N_9157,N_8990,N_8903);
and U9158 (N_9158,N_8002,N_7884);
and U9159 (N_9159,N_6110,N_7819);
nand U9160 (N_9160,N_8441,N_6549);
or U9161 (N_9161,N_7198,N_7300);
or U9162 (N_9162,N_6740,N_8602);
xor U9163 (N_9163,N_8795,N_6988);
or U9164 (N_9164,N_6485,N_6960);
nor U9165 (N_9165,N_7992,N_8153);
or U9166 (N_9166,N_7790,N_7018);
or U9167 (N_9167,N_7057,N_6604);
nand U9168 (N_9168,N_7137,N_6949);
nor U9169 (N_9169,N_8080,N_7442);
nor U9170 (N_9170,N_7054,N_7913);
and U9171 (N_9171,N_6757,N_7163);
and U9172 (N_9172,N_6109,N_6803);
nand U9173 (N_9173,N_7356,N_6360);
nand U9174 (N_9174,N_6824,N_7786);
or U9175 (N_9175,N_6821,N_7281);
or U9176 (N_9176,N_6551,N_7400);
and U9177 (N_9177,N_8400,N_7741);
xor U9178 (N_9178,N_8604,N_7088);
nor U9179 (N_9179,N_6369,N_6675);
or U9180 (N_9180,N_6262,N_6100);
and U9181 (N_9181,N_8881,N_8700);
nand U9182 (N_9182,N_6597,N_8147);
or U9183 (N_9183,N_8679,N_7581);
xor U9184 (N_9184,N_8626,N_7020);
and U9185 (N_9185,N_7608,N_8272);
nand U9186 (N_9186,N_6116,N_6624);
or U9187 (N_9187,N_7642,N_8436);
and U9188 (N_9188,N_6544,N_6621);
xor U9189 (N_9189,N_6989,N_7041);
and U9190 (N_9190,N_8058,N_6749);
nor U9191 (N_9191,N_8574,N_7473);
nand U9192 (N_9192,N_8313,N_6958);
xnor U9193 (N_9193,N_6342,N_8338);
and U9194 (N_9194,N_7783,N_8173);
xnor U9195 (N_9195,N_8405,N_8099);
and U9196 (N_9196,N_8247,N_8188);
and U9197 (N_9197,N_8454,N_7693);
nor U9198 (N_9198,N_6016,N_7804);
or U9199 (N_9199,N_8290,N_8156);
and U9200 (N_9200,N_8459,N_7700);
nand U9201 (N_9201,N_8514,N_8540);
or U9202 (N_9202,N_7424,N_8824);
or U9203 (N_9203,N_8144,N_7922);
and U9204 (N_9204,N_7169,N_7578);
nand U9205 (N_9205,N_6697,N_7316);
nor U9206 (N_9206,N_7196,N_7351);
and U9207 (N_9207,N_8356,N_8397);
nor U9208 (N_9208,N_7221,N_7926);
and U9209 (N_9209,N_7181,N_8221);
nand U9210 (N_9210,N_7677,N_7879);
nand U9211 (N_9211,N_6199,N_7572);
nand U9212 (N_9212,N_8098,N_8976);
nand U9213 (N_9213,N_7187,N_6759);
or U9214 (N_9214,N_8280,N_8755);
nand U9215 (N_9215,N_7942,N_7499);
or U9216 (N_9216,N_8729,N_8082);
and U9217 (N_9217,N_7277,N_8578);
or U9218 (N_9218,N_6941,N_7905);
or U9219 (N_9219,N_7426,N_7611);
nor U9220 (N_9220,N_8149,N_6075);
and U9221 (N_9221,N_6227,N_8476);
or U9222 (N_9222,N_7678,N_8621);
or U9223 (N_9223,N_6454,N_8091);
and U9224 (N_9224,N_7208,N_8335);
nand U9225 (N_9225,N_6455,N_8119);
and U9226 (N_9226,N_8455,N_7079);
nor U9227 (N_9227,N_6120,N_7051);
and U9228 (N_9228,N_7979,N_7710);
or U9229 (N_9229,N_6471,N_8861);
nand U9230 (N_9230,N_7416,N_7185);
nand U9231 (N_9231,N_7629,N_6070);
nor U9232 (N_9232,N_7524,N_7237);
nor U9233 (N_9233,N_6871,N_8306);
nor U9234 (N_9234,N_7545,N_6944);
nor U9235 (N_9235,N_6524,N_6046);
and U9236 (N_9236,N_6359,N_6205);
or U9237 (N_9237,N_8242,N_7914);
and U9238 (N_9238,N_7702,N_7427);
nand U9239 (N_9239,N_8770,N_6939);
xnor U9240 (N_9240,N_8162,N_7367);
xnor U9241 (N_9241,N_7105,N_6087);
or U9242 (N_9242,N_7767,N_6248);
and U9243 (N_9243,N_6005,N_7235);
and U9244 (N_9244,N_6267,N_6868);
and U9245 (N_9245,N_8369,N_6913);
and U9246 (N_9246,N_7111,N_6783);
xor U9247 (N_9247,N_7273,N_8288);
and U9248 (N_9248,N_7743,N_7030);
nand U9249 (N_9249,N_7563,N_6684);
or U9250 (N_9250,N_8041,N_6829);
nand U9251 (N_9251,N_6159,N_7544);
nor U9252 (N_9252,N_8006,N_7107);
nor U9253 (N_9253,N_6839,N_7007);
xor U9254 (N_9254,N_6742,N_8060);
nor U9255 (N_9255,N_7970,N_8406);
and U9256 (N_9256,N_8135,N_7858);
or U9257 (N_9257,N_6395,N_7506);
nand U9258 (N_9258,N_6206,N_8850);
or U9259 (N_9259,N_8993,N_8320);
nand U9260 (N_9260,N_8298,N_8371);
and U9261 (N_9261,N_6263,N_6231);
nor U9262 (N_9262,N_8348,N_7420);
nand U9263 (N_9263,N_8595,N_7380);
nand U9264 (N_9264,N_6181,N_8833);
and U9265 (N_9265,N_8651,N_6044);
or U9266 (N_9266,N_8477,N_7348);
or U9267 (N_9267,N_6492,N_7075);
xor U9268 (N_9268,N_7869,N_8458);
and U9269 (N_9269,N_7490,N_8435);
nor U9270 (N_9270,N_6093,N_6968);
xor U9271 (N_9271,N_7099,N_7685);
and U9272 (N_9272,N_8847,N_8256);
nand U9273 (N_9273,N_6566,N_7699);
or U9274 (N_9274,N_7717,N_7831);
nand U9275 (N_9275,N_8909,N_7415);
xnor U9276 (N_9276,N_6525,N_8286);
nor U9277 (N_9277,N_7791,N_7994);
xor U9278 (N_9278,N_7726,N_6143);
nand U9279 (N_9279,N_6666,N_6764);
nor U9280 (N_9280,N_7757,N_7094);
nor U9281 (N_9281,N_8680,N_6844);
or U9282 (N_9282,N_7392,N_8160);
and U9283 (N_9283,N_6951,N_7449);
nor U9284 (N_9284,N_7460,N_7928);
nand U9285 (N_9285,N_7112,N_7354);
and U9286 (N_9286,N_6973,N_6073);
nor U9287 (N_9287,N_7032,N_7453);
or U9288 (N_9288,N_7485,N_6383);
nor U9289 (N_9289,N_6322,N_6545);
nand U9290 (N_9290,N_6714,N_7833);
or U9291 (N_9291,N_8743,N_8427);
nor U9292 (N_9292,N_6683,N_8704);
nand U9293 (N_9293,N_8445,N_8857);
or U9294 (N_9294,N_6736,N_8778);
nand U9295 (N_9295,N_8834,N_7881);
and U9296 (N_9296,N_7363,N_7620);
and U9297 (N_9297,N_8409,N_8952);
or U9298 (N_9298,N_6539,N_8001);
and U9299 (N_9299,N_6156,N_8386);
or U9300 (N_9300,N_8127,N_6259);
or U9301 (N_9301,N_7735,N_6668);
and U9302 (N_9302,N_7512,N_6718);
nor U9303 (N_9303,N_6405,N_7211);
nor U9304 (N_9304,N_6815,N_8664);
nor U9305 (N_9305,N_8810,N_7607);
and U9306 (N_9306,N_7939,N_8576);
xor U9307 (N_9307,N_6361,N_8948);
and U9308 (N_9308,N_8349,N_7166);
nand U9309 (N_9309,N_7409,N_7045);
nand U9310 (N_9310,N_6052,N_8316);
nor U9311 (N_9311,N_7109,N_6928);
nand U9312 (N_9312,N_6634,N_8059);
or U9313 (N_9313,N_6664,N_6380);
xor U9314 (N_9314,N_8605,N_7977);
nor U9315 (N_9315,N_8463,N_8681);
or U9316 (N_9316,N_8968,N_7157);
nand U9317 (N_9317,N_6579,N_6606);
nand U9318 (N_9318,N_7766,N_7384);
nand U9319 (N_9319,N_8016,N_7450);
xor U9320 (N_9320,N_7465,N_7223);
nand U9321 (N_9321,N_8044,N_7787);
and U9322 (N_9322,N_8437,N_8543);
nor U9323 (N_9323,N_6936,N_7596);
nand U9324 (N_9324,N_7314,N_6719);
or U9325 (N_9325,N_6332,N_8167);
nor U9326 (N_9326,N_8613,N_7792);
xor U9327 (N_9327,N_7566,N_6638);
nor U9328 (N_9328,N_8854,N_7582);
and U9329 (N_9329,N_6446,N_7817);
or U9330 (N_9330,N_6375,N_6209);
and U9331 (N_9331,N_6688,N_7873);
xor U9332 (N_9332,N_7579,N_7243);
nor U9333 (N_9333,N_8521,N_6253);
nand U9334 (N_9334,N_8532,N_6576);
and U9335 (N_9335,N_8610,N_8859);
and U9336 (N_9336,N_8125,N_8159);
nand U9337 (N_9337,N_8512,N_6475);
nand U9338 (N_9338,N_7397,N_6971);
nand U9339 (N_9339,N_7845,N_8014);
or U9340 (N_9340,N_6594,N_8322);
and U9341 (N_9341,N_7050,N_8835);
nor U9342 (N_9342,N_6961,N_6404);
nor U9343 (N_9343,N_6050,N_8889);
xnor U9344 (N_9344,N_8061,N_7119);
and U9345 (N_9345,N_7507,N_8447);
nor U9346 (N_9346,N_6550,N_7631);
and U9347 (N_9347,N_6569,N_8913);
nand U9348 (N_9348,N_7141,N_7848);
xor U9349 (N_9349,N_8492,N_7643);
nand U9350 (N_9350,N_7610,N_7571);
nand U9351 (N_9351,N_6439,N_7011);
or U9352 (N_9352,N_7594,N_7092);
or U9353 (N_9353,N_6807,N_8032);
and U9354 (N_9354,N_8415,N_6410);
nand U9355 (N_9355,N_8827,N_6837);
and U9356 (N_9356,N_7584,N_6694);
or U9357 (N_9357,N_8749,N_6099);
and U9358 (N_9358,N_8223,N_6362);
and U9359 (N_9359,N_6589,N_8912);
or U9360 (N_9360,N_6516,N_6468);
nor U9361 (N_9361,N_7008,N_7917);
nor U9362 (N_9362,N_6903,N_7446);
nor U9363 (N_9363,N_6908,N_8327);
nor U9364 (N_9364,N_8739,N_6617);
nor U9365 (N_9365,N_6607,N_7753);
or U9366 (N_9366,N_6098,N_8139);
and U9367 (N_9367,N_7820,N_7469);
nor U9368 (N_9368,N_7500,N_6937);
or U9369 (N_9369,N_8511,N_6506);
nand U9370 (N_9370,N_6279,N_7429);
xnor U9371 (N_9371,N_8129,N_6969);
nand U9372 (N_9372,N_6832,N_6312);
nand U9373 (N_9373,N_7715,N_7476);
nor U9374 (N_9374,N_8871,N_8981);
or U9375 (N_9375,N_8361,N_6756);
nor U9376 (N_9376,N_8237,N_7805);
or U9377 (N_9377,N_8685,N_7206);
nor U9378 (N_9378,N_6954,N_7014);
and U9379 (N_9379,N_6084,N_7322);
or U9380 (N_9380,N_6058,N_6938);
nor U9381 (N_9381,N_6065,N_7532);
nor U9382 (N_9382,N_7093,N_6990);
xnor U9383 (N_9383,N_7675,N_8565);
nor U9384 (N_9384,N_8403,N_8323);
nor U9385 (N_9385,N_6458,N_6412);
nand U9386 (N_9386,N_8024,N_7304);
nand U9387 (N_9387,N_8697,N_7568);
nor U9388 (N_9388,N_8766,N_8267);
and U9389 (N_9389,N_8383,N_6271);
nand U9390 (N_9390,N_6509,N_6508);
or U9391 (N_9391,N_8525,N_6457);
or U9392 (N_9392,N_7379,N_8588);
and U9393 (N_9393,N_6117,N_6062);
xnor U9394 (N_9394,N_8257,N_7039);
xor U9395 (N_9395,N_8929,N_6701);
or U9396 (N_9396,N_6233,N_6353);
xor U9397 (N_9397,N_6905,N_7478);
and U9398 (N_9398,N_7656,N_6890);
and U9399 (N_9399,N_8172,N_6669);
nor U9400 (N_9400,N_7311,N_8717);
nand U9401 (N_9401,N_6247,N_7731);
and U9402 (N_9402,N_8112,N_6269);
nand U9403 (N_9403,N_8362,N_6366);
and U9404 (N_9404,N_7435,N_8950);
xnor U9405 (N_9405,N_7960,N_7318);
and U9406 (N_9406,N_6184,N_7529);
and U9407 (N_9407,N_6391,N_6613);
and U9408 (N_9408,N_8449,N_6580);
nand U9409 (N_9409,N_8885,N_7350);
or U9410 (N_9410,N_8984,N_8958);
and U9411 (N_9411,N_7666,N_8639);
xor U9412 (N_9412,N_8883,N_6782);
nor U9413 (N_9413,N_6221,N_6495);
and U9414 (N_9414,N_7302,N_8967);
nor U9415 (N_9415,N_8165,N_7526);
or U9416 (N_9416,N_7272,N_6082);
nand U9417 (N_9417,N_6874,N_8941);
nor U9418 (N_9418,N_8392,N_7431);
xor U9419 (N_9419,N_8318,N_8975);
nor U9420 (N_9420,N_6442,N_6261);
nor U9421 (N_9421,N_7556,N_8385);
nor U9422 (N_9422,N_6705,N_6307);
nand U9423 (N_9423,N_7821,N_7570);
nor U9424 (N_9424,N_8210,N_8259);
nor U9425 (N_9425,N_6507,N_8879);
nor U9426 (N_9426,N_8925,N_7555);
or U9427 (N_9427,N_8746,N_6722);
or U9428 (N_9428,N_6030,N_6825);
nor U9429 (N_9429,N_6816,N_7638);
nand U9430 (N_9430,N_6799,N_8742);
nor U9431 (N_9431,N_7851,N_7025);
and U9432 (N_9432,N_8299,N_7176);
nand U9433 (N_9433,N_6738,N_6559);
nor U9434 (N_9434,N_8617,N_8535);
xnor U9435 (N_9435,N_7222,N_7637);
nand U9436 (N_9436,N_6092,N_8844);
and U9437 (N_9437,N_8894,N_6208);
and U9438 (N_9438,N_8726,N_6418);
or U9439 (N_9439,N_6547,N_6288);
nor U9440 (N_9440,N_8750,N_6965);
and U9441 (N_9441,N_6758,N_7874);
or U9442 (N_9442,N_8354,N_6151);
nand U9443 (N_9443,N_8352,N_6421);
nor U9444 (N_9444,N_8970,N_7719);
or U9445 (N_9445,N_7540,N_7925);
or U9446 (N_9446,N_8563,N_7353);
and U9447 (N_9447,N_8040,N_8343);
and U9448 (N_9448,N_7393,N_6478);
nor U9449 (N_9449,N_6793,N_7430);
nand U9450 (N_9450,N_6608,N_7940);
xnor U9451 (N_9451,N_8841,N_7537);
or U9452 (N_9452,N_6323,N_8786);
and U9453 (N_9453,N_8330,N_6987);
and U9454 (N_9454,N_6693,N_8888);
nor U9455 (N_9455,N_7779,N_8728);
or U9456 (N_9456,N_8111,N_6632);
nor U9457 (N_9457,N_6033,N_6493);
and U9458 (N_9458,N_6315,N_8812);
nor U9459 (N_9459,N_6071,N_8800);
or U9460 (N_9460,N_7860,N_6474);
nand U9461 (N_9461,N_8490,N_7161);
nand U9462 (N_9462,N_6095,N_7636);
nand U9463 (N_9463,N_7718,N_8114);
or U9464 (N_9464,N_6300,N_7371);
nand U9465 (N_9465,N_6039,N_8753);
nor U9466 (N_9466,N_8363,N_7106);
and U9467 (N_9467,N_8577,N_8731);
and U9468 (N_9468,N_6852,N_7258);
or U9469 (N_9469,N_7437,N_6127);
and U9470 (N_9470,N_8481,N_7242);
xor U9471 (N_9471,N_6088,N_7299);
or U9472 (N_9472,N_6847,N_7328);
nand U9473 (N_9473,N_8768,N_6519);
and U9474 (N_9474,N_8101,N_7454);
nand U9475 (N_9475,N_8469,N_6210);
xor U9476 (N_9476,N_7070,N_7332);
and U9477 (N_9477,N_8897,N_8179);
and U9478 (N_9478,N_8009,N_8083);
nor U9479 (N_9479,N_6851,N_7711);
nor U9480 (N_9480,N_6450,N_8674);
nand U9481 (N_9481,N_8460,N_8814);
and U9482 (N_9482,N_7246,N_6568);
or U9483 (N_9483,N_7808,N_8914);
and U9484 (N_9484,N_6685,N_7095);
or U9485 (N_9485,N_8339,N_7857);
and U9486 (N_9486,N_8597,N_7130);
nor U9487 (N_9487,N_7346,N_7885);
nand U9488 (N_9488,N_8025,N_6811);
nand U9489 (N_9489,N_6678,N_7897);
nor U9490 (N_9490,N_7158,N_6326);
nor U9491 (N_9491,N_8434,N_8534);
or U9492 (N_9492,N_7590,N_8630);
nor U9493 (N_9493,N_8030,N_6215);
or U9494 (N_9494,N_8211,N_8329);
or U9495 (N_9495,N_8192,N_6861);
and U9496 (N_9496,N_7871,N_7403);
or U9497 (N_9497,N_6677,N_6703);
or U9498 (N_9498,N_7681,N_7716);
nand U9499 (N_9499,N_7689,N_7480);
nor U9500 (N_9500,N_8315,N_7038);
nor U9501 (N_9501,N_6431,N_7626);
xnor U9502 (N_9502,N_8422,N_8274);
nand U9503 (N_9503,N_7604,N_6356);
and U9504 (N_9504,N_6268,N_8628);
or U9505 (N_9505,N_7797,N_8519);
nand U9506 (N_9506,N_6691,N_6612);
nor U9507 (N_9507,N_8663,N_8891);
or U9508 (N_9508,N_7056,N_6543);
nand U9509 (N_9509,N_7891,N_6892);
nand U9510 (N_9510,N_6681,N_8533);
nand U9511 (N_9511,N_6056,N_6203);
and U9512 (N_9512,N_8774,N_7882);
and U9513 (N_9513,N_8359,N_8887);
and U9514 (N_9514,N_7956,N_7104);
nand U9515 (N_9515,N_8117,N_7978);
nor U9516 (N_9516,N_7861,N_6838);
nand U9517 (N_9517,N_7337,N_6523);
or U9518 (N_9518,N_6567,N_8278);
and U9519 (N_9519,N_6001,N_7971);
or U9520 (N_9520,N_6382,N_6862);
and U9521 (N_9521,N_7876,N_6754);
or U9522 (N_9522,N_7528,N_6006);
and U9523 (N_9523,N_8115,N_6881);
xnor U9524 (N_9524,N_6444,N_6036);
nand U9525 (N_9525,N_6707,N_8372);
nand U9526 (N_9526,N_8904,N_6443);
and U9527 (N_9527,N_7673,N_6334);
and U9528 (N_9528,N_7818,N_6571);
and U9529 (N_9529,N_6226,N_8065);
xor U9530 (N_9530,N_7336,N_8520);
and U9531 (N_9531,N_8972,N_8019);
xnor U9532 (N_9532,N_6223,N_6024);
and U9533 (N_9533,N_6336,N_6385);
and U9534 (N_9534,N_6155,N_8128);
nor U9535 (N_9535,N_7291,N_6294);
nand U9536 (N_9536,N_7153,N_7290);
and U9537 (N_9537,N_6540,N_7935);
nand U9538 (N_9538,N_7888,N_7511);
or U9539 (N_9539,N_7606,N_8983);
xnor U9540 (N_9540,N_6063,N_6590);
nand U9541 (N_9541,N_8707,N_8838);
or U9542 (N_9542,N_6317,N_7413);
nand U9543 (N_9543,N_7625,N_6013);
and U9544 (N_9544,N_8244,N_6435);
or U9545 (N_9545,N_7487,N_8347);
nor U9546 (N_9546,N_6108,N_6232);
or U9547 (N_9547,N_8606,N_8207);
xnor U9548 (N_9548,N_6835,N_6316);
or U9549 (N_9549,N_8271,N_6019);
nand U9550 (N_9550,N_7282,N_6358);
and U9551 (N_9551,N_7197,N_7827);
nand U9552 (N_9552,N_8759,N_8368);
or U9553 (N_9553,N_6611,N_6461);
or U9554 (N_9554,N_6152,N_6138);
or U9555 (N_9555,N_7004,N_7443);
nand U9556 (N_9556,N_8690,N_7521);
xor U9557 (N_9557,N_7411,N_8627);
nor U9558 (N_9558,N_6251,N_7525);
or U9559 (N_9559,N_8052,N_7080);
xor U9560 (N_9560,N_7984,N_8289);
nor U9561 (N_9561,N_6659,N_7175);
and U9562 (N_9562,N_6438,N_6310);
and U9563 (N_9563,N_8784,N_8730);
xor U9564 (N_9564,N_6301,N_7868);
or U9565 (N_9565,N_8505,N_8654);
nand U9566 (N_9566,N_7386,N_8608);
or U9567 (N_9567,N_8661,N_6752);
nand U9568 (N_9568,N_6401,N_8174);
nand U9569 (N_9569,N_6419,N_8495);
nand U9570 (N_9570,N_7033,N_6453);
nand U9571 (N_9571,N_8989,N_7026);
or U9572 (N_9572,N_6022,N_8262);
and U9573 (N_9573,N_7323,N_8884);
xnor U9574 (N_9574,N_6626,N_6119);
or U9575 (N_9575,N_7962,N_8105);
and U9576 (N_9576,N_7477,N_6304);
nand U9577 (N_9577,N_6165,N_6720);
nand U9578 (N_9578,N_8483,N_7100);
or U9579 (N_9579,N_6850,N_8554);
nor U9580 (N_9580,N_6695,N_6333);
xor U9581 (N_9581,N_7422,N_8266);
and U9582 (N_9582,N_8551,N_7705);
nand U9583 (N_9583,N_7167,N_7946);
nand U9584 (N_9584,N_6872,N_8017);
nand U9585 (N_9585,N_8214,N_7362);
xnor U9586 (N_9586,N_7680,N_8056);
nand U9587 (N_9587,N_8875,N_6768);
and U9588 (N_9588,N_8775,N_8837);
and U9589 (N_9589,N_8797,N_8667);
nor U9590 (N_9590,N_8756,N_7768);
and U9591 (N_9591,N_6348,N_8374);
nand U9592 (N_9592,N_6318,N_8767);
nand U9593 (N_9593,N_7295,N_8057);
xor U9594 (N_9594,N_7560,N_7856);
or U9595 (N_9595,N_6922,N_7624);
nor U9596 (N_9596,N_7832,N_8095);
xor U9597 (N_9597,N_6101,N_7973);
nor U9598 (N_9598,N_8293,N_6197);
or U9599 (N_9599,N_8273,N_8136);
xnor U9600 (N_9600,N_8263,N_6797);
nand U9601 (N_9601,N_6296,N_8688);
xnor U9602 (N_9602,N_7746,N_8226);
nand U9603 (N_9603,N_7143,N_8796);
or U9604 (N_9604,N_7261,N_6840);
or U9605 (N_9605,N_7738,N_7900);
or U9606 (N_9606,N_6980,N_6028);
and U9607 (N_9607,N_8716,N_8872);
nor U9608 (N_9608,N_6491,N_7005);
nand U9609 (N_9609,N_6096,N_7670);
and U9610 (N_9610,N_8113,N_7585);
nor U9611 (N_9611,N_6867,N_6107);
or U9612 (N_9612,N_7708,N_7333);
nand U9613 (N_9613,N_7682,N_8585);
or U9614 (N_9614,N_7248,N_7082);
or U9615 (N_9615,N_7676,N_7789);
or U9616 (N_9616,N_6734,N_6999);
and U9617 (N_9617,N_6351,N_8124);
or U9618 (N_9618,N_8340,N_8807);
xnor U9619 (N_9619,N_6784,N_8867);
nand U9620 (N_9620,N_8777,N_7358);
nor U9621 (N_9621,N_6700,N_8297);
nand U9622 (N_9622,N_6934,N_6884);
and U9623 (N_9623,N_8503,N_6526);
or U9624 (N_9624,N_7907,N_8429);
nor U9625 (N_9625,N_6529,N_7313);
xnor U9626 (N_9626,N_8583,N_6820);
nand U9627 (N_9627,N_8924,N_6955);
or U9628 (N_9628,N_7154,N_8131);
and U9629 (N_9629,N_8695,N_7255);
nor U9630 (N_9630,N_7937,N_7470);
nor U9631 (N_9631,N_6692,N_7136);
nor U9632 (N_9632,N_6202,N_8546);
and U9633 (N_9633,N_6465,N_7772);
nand U9634 (N_9634,N_8672,N_7968);
or U9635 (N_9635,N_7912,N_8670);
and U9636 (N_9636,N_6277,N_8504);
and U9637 (N_9637,N_7899,N_8453);
or U9638 (N_9638,N_7669,N_6186);
nor U9639 (N_9639,N_6389,N_6735);
nor U9640 (N_9640,N_6916,N_8013);
xnor U9641 (N_9641,N_8873,N_6555);
nand U9642 (N_9642,N_7640,N_7864);
xnor U9643 (N_9643,N_8696,N_8612);
nor U9644 (N_9644,N_7474,N_6643);
and U9645 (N_9645,N_6328,N_7834);
and U9646 (N_9646,N_8344,N_8246);
or U9647 (N_9647,N_7781,N_6076);
nor U9648 (N_9648,N_8868,N_7191);
and U9649 (N_9649,N_6066,N_8737);
nand U9650 (N_9650,N_8219,N_7815);
nand U9651 (N_9651,N_8564,N_6774);
and U9652 (N_9652,N_7975,N_7278);
xnor U9653 (N_9653,N_6560,N_6586);
nand U9654 (N_9654,N_7046,N_6252);
nor U9655 (N_9655,N_7148,N_6909);
and U9656 (N_9656,N_7653,N_7065);
and U9657 (N_9657,N_7121,N_8264);
xor U9658 (N_9658,N_8039,N_8255);
and U9659 (N_9659,N_8195,N_8931);
nor U9660 (N_9660,N_8880,N_7780);
nand U9661 (N_9661,N_7205,N_8736);
nand U9662 (N_9662,N_8580,N_7650);
nor U9663 (N_9663,N_8196,N_7765);
and U9664 (N_9664,N_6162,N_7116);
or U9665 (N_9665,N_6494,N_6682);
or U9666 (N_9666,N_8428,N_6522);
or U9667 (N_9667,N_8478,N_7965);
or U9668 (N_9668,N_8900,N_6856);
nor U9669 (N_9669,N_7788,N_7140);
and U9670 (N_9670,N_8843,N_7592);
nor U9671 (N_9671,N_7501,N_7006);
and U9672 (N_9672,N_6623,N_6995);
or U9673 (N_9673,N_8225,N_8412);
nor U9674 (N_9674,N_6198,N_7265);
and U9675 (N_9675,N_8738,N_6451);
nand U9676 (N_9676,N_8419,N_7407);
xor U9677 (N_9677,N_6150,N_7623);
nor U9678 (N_9678,N_8377,N_7486);
and U9679 (N_9679,N_8658,N_7574);
or U9680 (N_9680,N_7825,N_7599);
and U9681 (N_9681,N_8722,N_8236);
and U9682 (N_9682,N_6804,N_8793);
nand U9683 (N_9683,N_7172,N_7383);
nand U9684 (N_9684,N_7036,N_8806);
nand U9685 (N_9685,N_6139,N_8325);
and U9686 (N_9686,N_6595,N_7372);
nand U9687 (N_9687,N_8601,N_7382);
and U9688 (N_9688,N_7552,N_6308);
and U9689 (N_9689,N_8097,N_7999);
nor U9690 (N_9690,N_7806,N_8735);
or U9691 (N_9691,N_7319,N_6403);
xor U9692 (N_9692,N_7522,N_6699);
nand U9693 (N_9693,N_6182,N_7551);
xor U9694 (N_9694,N_7872,N_8170);
xor U9695 (N_9695,N_7591,N_6305);
and U9696 (N_9696,N_8677,N_6068);
nand U9697 (N_9697,N_6536,N_6292);
nor U9698 (N_9698,N_7122,N_7844);
and U9699 (N_9699,N_6003,N_7836);
xor U9700 (N_9700,N_6598,N_6956);
and U9701 (N_9701,N_6858,N_7343);
nor U9702 (N_9702,N_6190,N_7178);
or U9703 (N_9703,N_8590,N_7750);
nand U9704 (N_9704,N_7759,N_6064);
and U9705 (N_9705,N_6293,N_6842);
xor U9706 (N_9706,N_8951,N_7060);
nand U9707 (N_9707,N_6662,N_7756);
nand U9708 (N_9708,N_6570,N_6285);
nor U9709 (N_9709,N_8584,N_6020);
or U9710 (N_9710,N_6548,N_7132);
and U9711 (N_9711,N_8222,N_7724);
and U9712 (N_9712,N_7896,N_7762);
or U9713 (N_9713,N_8076,N_7990);
and U9714 (N_9714,N_6373,N_7177);
xnor U9715 (N_9715,N_7587,N_6456);
nor U9716 (N_9716,N_8277,N_7880);
or U9717 (N_9717,N_8529,N_6228);
and U9718 (N_9718,N_7559,N_7763);
nor U9719 (N_9719,N_7438,N_7010);
nor U9720 (N_9720,N_6599,N_8410);
nor U9721 (N_9721,N_6281,N_6585);
nand U9722 (N_9722,N_8846,N_7671);
nor U9723 (N_9723,N_8823,N_6912);
and U9724 (N_9724,N_8497,N_8689);
nor U9725 (N_9725,N_6464,N_7250);
nor U9726 (N_9726,N_7401,N_7687);
nand U9727 (N_9727,N_8877,N_8292);
nor U9728 (N_9728,N_6859,N_8430);
and U9729 (N_9729,N_7234,N_6250);
xor U9730 (N_9730,N_7144,N_8283);
and U9731 (N_9731,N_7933,N_7069);
and U9732 (N_9732,N_7800,N_6499);
and U9733 (N_9733,N_6796,N_8276);
nand U9734 (N_9734,N_6953,N_6521);
or U9735 (N_9735,N_7441,N_6025);
or U9736 (N_9736,N_8963,N_6577);
or U9737 (N_9737,N_8321,N_6962);
nor U9738 (N_9738,N_8591,N_7162);
and U9739 (N_9739,N_8141,N_8104);
nor U9740 (N_9740,N_7019,N_8033);
or U9741 (N_9741,N_6433,N_8971);
and U9742 (N_9742,N_8072,N_6429);
nand U9743 (N_9743,N_8069,N_7182);
and U9744 (N_9744,N_8579,N_8769);
nor U9745 (N_9745,N_6921,N_7536);
or U9746 (N_9746,N_8045,N_8713);
nor U9747 (N_9747,N_6945,N_8802);
and U9748 (N_9748,N_8000,N_8100);
and U9749 (N_9749,N_8553,N_8457);
nand U9750 (N_9750,N_7729,N_7496);
nand U9751 (N_9751,N_7283,N_6557);
or U9752 (N_9752,N_6649,N_6490);
or U9753 (N_9753,N_7436,N_6647);
nor U9754 (N_9754,N_7068,N_6131);
nand U9755 (N_9755,N_6641,N_6584);
xor U9756 (N_9756,N_6582,N_7285);
nor U9757 (N_9757,N_8220,N_8782);
xnor U9758 (N_9758,N_6879,N_8120);
nand U9759 (N_9759,N_7489,N_6166);
and U9760 (N_9760,N_8957,N_8048);
xnor U9761 (N_9761,N_6029,N_8776);
or U9762 (N_9762,N_8408,N_8935);
or U9763 (N_9763,N_6925,N_6633);
nor U9764 (N_9764,N_6140,N_8296);
and U9765 (N_9765,N_8202,N_7459);
nor U9766 (N_9766,N_7508,N_7784);
nand U9767 (N_9767,N_6747,N_8305);
nand U9768 (N_9768,N_7667,N_7843);
nor U9769 (N_9769,N_8388,N_8094);
and U9770 (N_9770,N_6194,N_6480);
nor U9771 (N_9771,N_8465,N_7330);
or U9772 (N_9772,N_8665,N_6416);
and U9773 (N_9773,N_6347,N_7801);
xor U9774 (N_9774,N_6017,N_6575);
and U9775 (N_9775,N_7959,N_7458);
and U9776 (N_9776,N_7516,N_8587);
nor U9777 (N_9777,N_6276,N_7395);
nand U9778 (N_9778,N_6603,N_6327);
or U9779 (N_9779,N_7268,N_8440);
xnor U9780 (N_9780,N_8998,N_8209);
or U9781 (N_9781,N_6855,N_8908);
nor U9782 (N_9782,N_8042,N_7128);
nand U9783 (N_9783,N_7932,N_8845);
and U9784 (N_9784,N_7073,N_8232);
nor U9785 (N_9785,N_6041,N_6257);
and U9786 (N_9786,N_6037,N_7878);
nor U9787 (N_9787,N_7249,N_7696);
nand U9788 (N_9788,N_7548,N_8821);
nor U9789 (N_9789,N_8110,N_8068);
nand U9790 (N_9790,N_6512,N_7627);
or U9791 (N_9791,N_6933,N_8918);
nor U9792 (N_9792,N_8536,N_8550);
nor U9793 (N_9793,N_8275,N_6902);
and U9794 (N_9794,N_8015,N_7001);
and U9795 (N_9795,N_8180,N_7324);
and U9796 (N_9796,N_7423,N_6911);
xor U9797 (N_9797,N_6618,N_8103);
or U9798 (N_9798,N_8928,N_8407);
and U9799 (N_9799,N_6687,N_6860);
and U9800 (N_9800,N_8268,N_7220);
and U9801 (N_9801,N_6422,N_6537);
or U9802 (N_9802,N_8762,N_6436);
and U9803 (N_9803,N_6733,N_7086);
or U9804 (N_9804,N_7455,N_6857);
nand U9805 (N_9805,N_6818,N_8143);
and U9806 (N_9806,N_7775,N_7129);
xnor U9807 (N_9807,N_6964,N_6532);
nor U9808 (N_9808,N_8391,N_6284);
or U9809 (N_9809,N_8706,N_8765);
xnor U9810 (N_9810,N_7520,N_6079);
xnor U9811 (N_9811,N_8624,N_6676);
xnor U9812 (N_9812,N_6773,N_6542);
and U9813 (N_9813,N_7096,N_6147);
nor U9814 (N_9814,N_6853,N_7649);
nor U9815 (N_9815,N_7852,N_7467);
or U9816 (N_9816,N_8376,N_8703);
nor U9817 (N_9817,N_7209,N_7840);
or U9818 (N_9818,N_6015,N_7728);
nor U9819 (N_9819,N_7668,N_6896);
and U9820 (N_9820,N_7842,N_7028);
nand U9821 (N_9821,N_7305,N_6164);
nor U9822 (N_9822,N_6222,N_8253);
nor U9823 (N_9823,N_8758,N_7042);
xnor U9824 (N_9824,N_7981,N_7530);
and U9825 (N_9825,N_8451,N_6926);
xor U9826 (N_9826,N_8614,N_8863);
nand U9827 (N_9827,N_7201,N_7366);
nand U9828 (N_9828,N_8973,N_8656);
nand U9829 (N_9829,N_6899,N_7055);
xnor U9830 (N_9830,N_6054,N_6103);
or U9831 (N_9831,N_6400,N_7118);
nand U9832 (N_9832,N_6427,N_7252);
nand U9833 (N_9833,N_7482,N_8239);
nor U9834 (N_9834,N_7519,N_7034);
nor U9835 (N_9835,N_7739,N_8164);
nor U9836 (N_9836,N_6724,N_7890);
nor U9837 (N_9837,N_8593,N_6663);
nand U9838 (N_9838,N_8390,N_7083);
or U9839 (N_9839,N_8250,N_6541);
and U9840 (N_9840,N_8542,N_6193);
nand U9841 (N_9841,N_8234,N_8038);
or U9842 (N_9842,N_7149,N_6966);
or U9843 (N_9843,N_8249,N_6201);
nor U9844 (N_9844,N_8569,N_6390);
nor U9845 (N_9845,N_8619,N_8418);
nand U9846 (N_9846,N_7139,N_7432);
nor U9847 (N_9847,N_6055,N_7491);
or U9848 (N_9848,N_6081,N_8999);
nand U9849 (N_9849,N_8425,N_6424);
nor U9850 (N_9850,N_7471,N_8607);
or U9851 (N_9851,N_6121,N_8804);
and U9852 (N_9852,N_8864,N_8902);
nand U9853 (N_9853,N_8899,N_6176);
and U9854 (N_9854,N_8573,N_8637);
or U9855 (N_9855,N_6984,N_6207);
or U9856 (N_9856,N_7964,N_7173);
nor U9857 (N_9857,N_6817,N_7953);
and U9858 (N_9858,N_6952,N_8819);
or U9859 (N_9859,N_7284,N_7704);
nand U9860 (N_9860,N_6330,N_8081);
or U9861 (N_9861,N_8611,N_7434);
nor U9862 (N_9862,N_8956,N_6809);
xnor U9863 (N_9863,N_6097,N_8370);
and U9864 (N_9864,N_6417,N_8790);
or U9865 (N_9865,N_8816,N_6324);
nor U9866 (N_9866,N_7727,N_7771);
or U9867 (N_9867,N_8657,N_7645);
or U9868 (N_9868,N_8803,N_8648);
or U9869 (N_9869,N_8832,N_6225);
or U9870 (N_9870,N_7569,N_7993);
xnor U9871 (N_9871,N_6246,N_6822);
and U9872 (N_9872,N_7920,N_8629);
nor U9873 (N_9873,N_6667,N_6510);
xnor U9874 (N_9874,N_7110,N_8720);
and U9875 (N_9875,N_6130,N_7067);
or U9876 (N_9876,N_8206,N_6514);
nor U9877 (N_9877,N_8641,N_6848);
nor U9878 (N_9878,N_8905,N_7543);
nor U9879 (N_9879,N_6335,N_7292);
and U9880 (N_9880,N_6441,N_8598);
nand U9881 (N_9881,N_6843,N_6732);
or U9882 (N_9882,N_6725,N_7982);
nand U9883 (N_9883,N_8431,N_8575);
nor U9884 (N_9884,N_8432,N_7224);
or U9885 (N_9885,N_6957,N_8801);
nor U9886 (N_9886,N_6460,N_7216);
nand U9887 (N_9887,N_6630,N_8161);
nand U9888 (N_9888,N_6026,N_7479);
xnor U9889 (N_9889,N_8364,N_7732);
or U9890 (N_9890,N_6467,N_7807);
or U9891 (N_9891,N_8528,N_7698);
and U9892 (N_9892,N_7795,N_6340);
or U9893 (N_9893,N_8943,N_7308);
and U9894 (N_9894,N_6331,N_8079);
and U9895 (N_9895,N_8071,N_8411);
nand U9896 (N_9896,N_8417,N_8468);
xnor U9897 (N_9897,N_7320,N_7481);
nand U9898 (N_9898,N_7744,N_8687);
and U9899 (N_9899,N_6264,N_7721);
and U9900 (N_9900,N_6721,N_8515);
nor U9901 (N_9901,N_8541,N_7230);
xor U9902 (N_9902,N_8401,N_8581);
nor U9903 (N_9903,N_6706,N_8509);
and U9904 (N_9904,N_6748,N_6834);
xor U9905 (N_9905,N_6142,N_7385);
or U9906 (N_9906,N_7695,N_7254);
or U9907 (N_9907,N_6931,N_7361);
nor U9908 (N_9908,N_7948,N_8531);
nand U9909 (N_9909,N_8927,N_7613);
or U9910 (N_9910,N_7630,N_7269);
or U9911 (N_9911,N_7747,N_7902);
or U9912 (N_9912,N_7017,N_6923);
or U9913 (N_9913,N_8732,N_7089);
nand U9914 (N_9914,N_6180,N_7023);
nor U9915 (N_9915,N_8398,N_7238);
nand U9916 (N_9916,N_7012,N_6831);
and U9917 (N_9917,N_7646,N_8307);
or U9918 (N_9918,N_6563,N_6469);
nor U9919 (N_9919,N_6449,N_7794);
nand U9920 (N_9920,N_8023,N_7404);
nor U9921 (N_9921,N_8906,N_6601);
and U9922 (N_9922,N_6765,N_7024);
or U9923 (N_9923,N_6865,N_7022);
and U9924 (N_9924,N_6191,N_6045);
and U9925 (N_9925,N_8474,N_7127);
and U9926 (N_9926,N_7301,N_8618);
and U9927 (N_9927,N_7183,N_8724);
xnor U9928 (N_9928,N_6278,N_8557);
and U9929 (N_9929,N_7893,N_6368);
or U9930 (N_9930,N_6622,N_6299);
and U9931 (N_9931,N_8866,N_7398);
nor U9932 (N_9932,N_7692,N_7847);
nand U9933 (N_9933,N_7365,N_6220);
nand U9934 (N_9934,N_7910,N_7782);
or U9935 (N_9935,N_6113,N_6778);
nand U9936 (N_9936,N_6153,N_6218);
and U9937 (N_9937,N_7553,N_6136);
nor U9938 (N_9938,N_7101,N_8302);
nor U9939 (N_9939,N_6357,N_6772);
or U9940 (N_9940,N_7150,N_6743);
nor U9941 (N_9941,N_8310,N_7228);
nand U9942 (N_9942,N_6398,N_7564);
nand U9943 (N_9943,N_7293,N_7995);
and U9944 (N_9944,N_7102,N_6982);
and U9945 (N_9945,N_8516,N_8248);
and U9946 (N_9946,N_7901,N_7877);
and U9947 (N_9947,N_7903,N_8284);
and U9948 (N_9948,N_6287,N_8852);
nor U9949 (N_9949,N_8518,N_6275);
and U9950 (N_9950,N_7989,N_6270);
nand U9951 (N_9951,N_7565,N_6106);
and U9952 (N_9952,N_6997,N_7966);
nor U9953 (N_9953,N_7245,N_8181);
nor U9954 (N_9954,N_8781,N_6690);
or U9955 (N_9955,N_6907,N_8502);
xnor U9956 (N_9956,N_8314,N_8496);
nor U9957 (N_9957,N_6325,N_8204);
xor U9958 (N_9958,N_8965,N_7659);
nand U9959 (N_9959,N_7514,N_8603);
xnor U9960 (N_9960,N_8638,N_8133);
and U9961 (N_9961,N_8568,N_6282);
and U9962 (N_9962,N_7961,N_8134);
nor U9963 (N_9963,N_8622,N_7126);
nand U9964 (N_9964,N_7612,N_8792);
xnor U9965 (N_9965,N_8829,N_6053);
or U9966 (N_9966,N_8660,N_7927);
and U9967 (N_9967,N_7841,N_8396);
xor U9968 (N_9968,N_7577,N_6171);
or U9969 (N_9969,N_8116,N_8489);
or U9970 (N_9970,N_7958,N_6996);
nor U9971 (N_9971,N_7189,N_7215);
nand U9972 (N_9972,N_6178,N_6083);
or U9973 (N_9973,N_8493,N_6297);
xnor U9974 (N_9974,N_8171,N_6741);
nor U9975 (N_9975,N_7622,N_6423);
nor U9976 (N_9976,N_7632,N_8926);
nand U9977 (N_9977,N_8012,N_8794);
nor U9978 (N_9978,N_7733,N_7527);
nand U9979 (N_9979,N_8389,N_7497);
and U9980 (N_9980,N_8067,N_8856);
and U9981 (N_9981,N_8358,N_8175);
nor U9982 (N_9982,N_7164,N_6169);
nand U9983 (N_9983,N_8727,N_8954);
and U9984 (N_9984,N_6105,N_6102);
or U9985 (N_9985,N_6530,N_6260);
and U9986 (N_9986,N_8213,N_8245);
xor U9987 (N_9987,N_8169,N_8309);
nor U9988 (N_9988,N_7274,N_8243);
nand U9989 (N_9989,N_6311,N_8659);
and U9990 (N_9990,N_7452,N_8380);
or U9991 (N_9991,N_6798,N_7309);
nor U9992 (N_9992,N_8815,N_6702);
or U9993 (N_9993,N_6644,N_8939);
or U9994 (N_9994,N_8379,N_6849);
nand U9995 (N_9995,N_8849,N_8472);
and U9996 (N_9996,N_6616,N_8754);
nor U9997 (N_9997,N_8560,N_7098);
or U9998 (N_9998,N_8718,N_6175);
nor U9999 (N_9999,N_8037,N_6731);
or U10000 (N_10000,N_6917,N_7204);
or U10001 (N_10001,N_7983,N_6830);
nor U10002 (N_10002,N_6602,N_6605);
nand U10003 (N_10003,N_8995,N_6354);
nand U10004 (N_10004,N_7151,N_7389);
or U10005 (N_10005,N_7113,N_6642);
or U10006 (N_10006,N_8155,N_8524);
or U10007 (N_10007,N_8878,N_6729);
and U10008 (N_10008,N_7345,N_8666);
nor U10009 (N_10009,N_6794,N_8227);
nand U10010 (N_10010,N_7991,N_8055);
or U10011 (N_10011,N_8452,N_6012);
nand U10012 (N_10012,N_8699,N_6888);
nand U10013 (N_10013,N_8387,N_6397);
nor U10014 (N_10014,N_7425,N_6002);
and U10015 (N_10015,N_6235,N_6321);
xnor U10016 (N_10016,N_7190,N_7703);
and U10017 (N_10017,N_7576,N_6273);
nand U10018 (N_10018,N_6593,N_6991);
and U10019 (N_10019,N_8644,N_7071);
nand U10020 (N_10020,N_8200,N_6878);
and U10021 (N_10021,N_8547,N_6503);
nand U10022 (N_10022,N_6710,N_6224);
nor U10023 (N_10023,N_7709,N_7387);
xnor U10024 (N_10024,N_7539,N_7849);
and U10025 (N_10025,N_6069,N_6730);
and U10026 (N_10026,N_6827,N_8522);
nand U10027 (N_10027,N_7097,N_6047);
xor U10028 (N_10028,N_8007,N_7135);
or U10029 (N_10029,N_6091,N_6805);
nor U10030 (N_10030,N_8694,N_6974);
nor U10031 (N_10031,N_6755,N_8241);
nor U10032 (N_10032,N_7123,N_8317);
nand U10033 (N_10033,N_7193,N_8282);
xor U10034 (N_10034,N_8869,N_7619);
or U10035 (N_10035,N_8300,N_7996);
or U10036 (N_10036,N_8561,N_6219);
and U10037 (N_10037,N_8771,N_6708);
nand U10038 (N_10038,N_7396,N_8820);
and U10039 (N_10039,N_8295,N_8702);
nand U10040 (N_10040,N_8142,N_7674);
nor U10041 (N_10041,N_6588,N_8393);
nand U10042 (N_10042,N_8798,N_8231);
nor U10043 (N_10043,N_8752,N_6265);
or U10044 (N_10044,N_8308,N_7257);
and U10045 (N_10045,N_8224,N_8350);
nor U10046 (N_10046,N_8066,N_7195);
nand U10047 (N_10047,N_7251,N_6891);
and U10048 (N_10048,N_7419,N_7192);
and U10049 (N_10049,N_6770,N_7976);
nand U10050 (N_10050,N_6234,N_8808);
nor U10051 (N_10051,N_7199,N_6562);
or U10052 (N_10052,N_8964,N_8537);
nor U10053 (N_10053,N_8668,N_8733);
or U10054 (N_10054,N_7262,N_6200);
or U10055 (N_10055,N_8384,N_8708);
nor U10056 (N_10056,N_8570,N_6709);
and U10057 (N_10057,N_7410,N_8285);
and U10058 (N_10058,N_7156,N_6345);
nand U10059 (N_10059,N_8494,N_6482);
nand U10060 (N_10060,N_8947,N_7597);
or U10061 (N_10061,N_6726,N_8886);
and U10062 (N_10062,N_6500,N_7053);
xor U10063 (N_10063,N_8539,N_8592);
nand U10064 (N_10064,N_6452,N_7561);
nand U10065 (N_10065,N_8673,N_6306);
or U10066 (N_10066,N_6057,N_6646);
nor U10067 (N_10067,N_7412,N_6344);
nor U10068 (N_10068,N_6679,N_6628);
nand U10069 (N_10069,N_6564,N_7688);
nor U10070 (N_10070,N_8991,N_8662);
and U10071 (N_10071,N_8901,N_6511);
and U10072 (N_10072,N_6240,N_7998);
or U10073 (N_10073,N_6534,N_6836);
nor U10074 (N_10074,N_7824,N_6258);
or U10075 (N_10075,N_7583,N_8018);
nor U10076 (N_10076,N_7240,N_6229);
nor U10077 (N_10077,N_6914,N_6637);
nor U10078 (N_10078,N_7785,N_8538);
and U10079 (N_10079,N_6513,N_7468);
nor U10080 (N_10080,N_6761,N_7439);
nand U10081 (N_10081,N_7769,N_8633);
nor U10082 (N_10082,N_7227,N_6806);
xnor U10083 (N_10083,N_7090,N_8636);
nand U10084 (N_10084,N_7462,N_7029);
nand U10085 (N_10085,N_8254,N_7142);
and U10086 (N_10086,N_7835,N_6129);
or U10087 (N_10087,N_6556,N_7883);
or U10088 (N_10088,N_8132,N_7554);
or U10089 (N_10089,N_8734,N_8108);
nor U10090 (N_10090,N_7456,N_8969);
and U10091 (N_10091,N_7027,N_8092);
nand U10092 (N_10092,N_8994,N_8655);
or U10093 (N_10093,N_7186,N_6791);
and U10094 (N_10094,N_7523,N_8326);
or U10095 (N_10095,N_6943,N_8684);
or U10096 (N_10096,N_6812,N_6823);
nor U10097 (N_10097,N_8208,N_6195);
or U10098 (N_10098,N_6600,N_8510);
and U10099 (N_10099,N_6018,N_7494);
xnor U10100 (N_10100,N_8228,N_7854);
nand U10101 (N_10101,N_7830,N_6870);
xor U10102 (N_10102,N_6886,N_7002);
and U10103 (N_10103,N_8194,N_7969);
nand U10104 (N_10104,N_7908,N_6929);
or U10105 (N_10105,N_8106,N_6497);
nor U10106 (N_10106,N_7253,N_6572);
and U10107 (N_10107,N_8028,N_6959);
nor U10108 (N_10108,N_7344,N_6196);
nor U10109 (N_10109,N_7226,N_6745);
nor U10110 (N_10110,N_7947,N_8817);
nor U10111 (N_10111,N_7929,N_6795);
and U10112 (N_10112,N_6518,N_6346);
xor U10113 (N_10113,N_7918,N_6887);
or U10114 (N_10114,N_8761,N_7549);
or U10115 (N_10115,N_6790,N_6371);
nor U10116 (N_10116,N_6489,N_7202);
and U10117 (N_10117,N_6167,N_8148);
and U10118 (N_10118,N_8615,N_7760);
xor U10119 (N_10119,N_6000,N_7660);
xor U10120 (N_10120,N_6112,N_6531);
and U10121 (N_10121,N_6728,N_6515);
nand U10122 (N_10122,N_6483,N_8351);
nor U10123 (N_10123,N_8464,N_8855);
nand U10124 (N_10124,N_6920,N_6712);
nor U10125 (N_10125,N_6527,N_6535);
or U10126 (N_10126,N_8151,N_7276);
and U10127 (N_10127,N_7672,N_8488);
xor U10128 (N_10128,N_8862,N_8818);
or U10129 (N_10129,N_7635,N_7031);
nor U10130 (N_10130,N_8741,N_7915);
nand U10131 (N_10131,N_8895,N_8936);
or U10132 (N_10132,N_8785,N_8916);
or U10133 (N_10133,N_6411,N_6828);
nand U10134 (N_10134,N_6885,N_7444);
or U10135 (N_10135,N_7232,N_6498);
nor U10136 (N_10136,N_7329,N_7980);
or U10137 (N_10137,N_6280,N_6686);
or U10138 (N_10138,N_8152,N_7368);
and U10139 (N_10139,N_7321,N_6462);
nor U10140 (N_10140,N_7778,N_8723);
nor U10141 (N_10141,N_8710,N_7725);
or U10142 (N_10142,N_8053,N_7504);
nor U10143 (N_10143,N_8035,N_6338);
and U10144 (N_10144,N_8642,N_6004);
nand U10145 (N_10145,N_7963,N_6897);
or U10146 (N_10146,N_8291,N_8669);
nand U10147 (N_10147,N_6657,N_7533);
nand U10148 (N_10148,N_7152,N_8764);
nand U10149 (N_10149,N_6767,N_8433);
or U10150 (N_10150,N_6114,N_7081);
and U10151 (N_10151,N_6854,N_6781);
xor U10152 (N_10152,N_8559,N_7761);
or U10153 (N_10153,N_8145,N_7133);
xor U10154 (N_10154,N_7214,N_7706);
and U10155 (N_10155,N_8780,N_7355);
nor U10156 (N_10156,N_7374,N_8036);
nand U10157 (N_10157,N_7352,N_6715);
and U10158 (N_10158,N_8582,N_8230);
nand U10159 (N_10159,N_6845,N_6636);
nor U10160 (N_10160,N_8084,N_8693);
nand U10161 (N_10161,N_7475,N_6779);
nor U10162 (N_10162,N_7171,N_6128);
nand U10163 (N_10163,N_8333,N_8783);
nand U10164 (N_10164,N_8572,N_8840);
or U10165 (N_10165,N_8450,N_7538);
or U10166 (N_10166,N_7773,N_7433);
xnor U10167 (N_10167,N_6031,N_6168);
or U10168 (N_10168,N_6387,N_8381);
nand U10169 (N_10169,N_7058,N_6466);
xor U10170 (N_10170,N_6040,N_6430);
or U10171 (N_10171,N_7072,N_6813);
and U10172 (N_10172,N_6320,N_7447);
and U10173 (N_10173,N_6769,N_6900);
and U10174 (N_10174,N_7408,N_8473);
and U10175 (N_10175,N_7325,N_6978);
xor U10176 (N_10176,N_6042,N_8279);
nor U10177 (N_10177,N_6393,N_7138);
and U10178 (N_10178,N_7388,N_8997);
xor U10179 (N_10179,N_8426,N_8176);
and U10180 (N_10180,N_7654,N_6986);
and U10181 (N_10181,N_7505,N_7134);
and U10182 (N_10182,N_7641,N_7952);
and U10183 (N_10183,N_8992,N_7575);
and U10184 (N_10184,N_7239,N_7326);
and U10185 (N_10185,N_6060,N_8438);
and U10186 (N_10186,N_8945,N_6800);
nor U10187 (N_10187,N_6384,N_7616);
nand U10188 (N_10188,N_7390,N_7495);
and U10189 (N_10189,N_6160,N_8470);
nor U10190 (N_10190,N_6651,N_7930);
or U10191 (N_10191,N_8420,N_7021);
nand U10192 (N_10192,N_7493,N_6553);
and U10193 (N_10193,N_7828,N_6750);
nor U10194 (N_10194,N_8865,N_6216);
and U10195 (N_10195,N_7954,N_7679);
nor U10196 (N_10196,N_8650,N_7967);
nand U10197 (N_10197,N_8870,N_6274);
and U10198 (N_10198,N_6009,N_6407);
or U10199 (N_10199,N_8137,N_7974);
nand U10200 (N_10200,N_7707,N_7816);
or U10201 (N_10201,N_8715,N_6983);
nand U10202 (N_10202,N_8366,N_7044);
xnor U10203 (N_10203,N_8189,N_8199);
or U10204 (N_10204,N_7280,N_7541);
and U10205 (N_10205,N_8966,N_8022);
or U10206 (N_10206,N_6290,N_6011);
nand U10207 (N_10207,N_7798,N_7713);
and U10208 (N_10208,N_8874,N_7294);
nor U10209 (N_10209,N_7040,N_6023);
or U10210 (N_10210,N_7895,N_8949);
nand U10211 (N_10211,N_6185,N_6214);
nor U10212 (N_10212,N_7418,N_7297);
xor U10213 (N_10213,N_7009,N_6737);
nor U10214 (N_10214,N_7339,N_7059);
or U10215 (N_10215,N_8186,N_6470);
xnor U10216 (N_10216,N_8178,N_7951);
nor U10217 (N_10217,N_7335,N_6377);
nor U10218 (N_10218,N_8600,N_6998);
nor U10219 (N_10219,N_6032,N_8461);
nor U10220 (N_10220,N_7593,N_6319);
nand U10221 (N_10221,N_8216,N_8265);
or U10222 (N_10222,N_7125,N_7303);
nor U10223 (N_10223,N_7986,N_8836);
nand U10224 (N_10224,N_7749,N_6894);
nor U10225 (N_10225,N_8986,N_6459);
and U10226 (N_10226,N_7955,N_6409);
nor U10227 (N_10227,N_6043,N_8031);
nand U10228 (N_10228,N_6994,N_6635);
and U10229 (N_10229,N_8809,N_8270);
nand U10230 (N_10230,N_8466,N_7651);
and U10231 (N_10231,N_6918,N_6122);
or U10232 (N_10232,N_6212,N_6118);
or U10233 (N_10233,N_6763,N_6476);
or U10234 (N_10234,N_6080,N_7517);
nor U10235 (N_10235,N_8911,N_6145);
nor U10236 (N_10236,N_6930,N_7567);
or U10237 (N_10237,N_8399,N_8960);
nor U10238 (N_10238,N_6652,N_6378);
and U10239 (N_10239,N_8567,N_8711);
nand U10240 (N_10240,N_7381,N_8491);
and U10241 (N_10241,N_6977,N_7748);
or U10242 (N_10242,N_8544,N_8046);
nand U10243 (N_10243,N_8513,N_7062);
and U10244 (N_10244,N_6970,N_6313);
and U10245 (N_10245,N_8201,N_6437);
nand U10246 (N_10246,N_8915,N_8191);
nand U10247 (N_10247,N_8319,N_8779);
nor U10248 (N_10248,N_7463,N_7391);
or U10249 (N_10249,N_7375,N_6620);
or U10250 (N_10250,N_8653,N_6558);
or U10251 (N_10251,N_7657,N_7919);
or U10252 (N_10252,N_7938,N_6819);
and U10253 (N_10253,N_7621,N_7464);
nor U10254 (N_10254,N_7405,N_7078);
nor U10255 (N_10255,N_8811,N_7684);
and U10256 (N_10256,N_6591,N_6592);
nand U10257 (N_10257,N_6574,N_7812);
or U10258 (N_10258,N_8480,N_7557);
or U10259 (N_10259,N_6538,N_8562);
or U10260 (N_10260,N_8375,N_8760);
or U10261 (N_10261,N_6486,N_7247);
and U10262 (N_10262,N_8917,N_7944);
nor U10263 (N_10263,N_6609,N_8745);
or U10264 (N_10264,N_8955,N_6146);
nand U10265 (N_10265,N_8813,N_6680);
and U10266 (N_10266,N_8839,N_7402);
xnor U10267 (N_10267,N_6935,N_8530);
nand U10268 (N_10268,N_8355,N_8304);
nor U10269 (N_10269,N_6771,N_6792);
nor U10270 (N_10270,N_6583,N_8599);
and U10271 (N_10271,N_7084,N_6049);
or U10272 (N_10272,N_6479,N_7451);
and U10273 (N_10273,N_7886,N_7662);
nor U10274 (N_10274,N_7165,N_6904);
nor U10275 (N_10275,N_7076,N_7035);
nand U10276 (N_10276,N_6406,N_7714);
nand U10277 (N_10277,N_7466,N_6170);
nand U10278 (N_10278,N_6217,N_8212);
nand U10279 (N_10279,N_7369,N_8086);
or U10280 (N_10280,N_8623,N_6674);
nand U10281 (N_10281,N_7904,N_7923);
or U10282 (N_10282,N_8252,N_8647);
and U10283 (N_10283,N_7921,N_6587);
and U10284 (N_10284,N_6801,N_7145);
nor U10285 (N_10285,N_7484,N_8805);
and U10286 (N_10286,N_6615,N_7037);
and U10287 (N_10287,N_8953,N_6673);
nand U10288 (N_10288,N_7898,N_8373);
nand U10289 (N_10289,N_6502,N_6341);
and U10290 (N_10290,N_7697,N_6520);
nor U10291 (N_10291,N_6010,N_7887);
nor U10292 (N_10292,N_6426,N_7535);
and U10293 (N_10293,N_7263,N_8421);
nand U10294 (N_10294,N_6979,N_8258);
and U10295 (N_10295,N_8788,N_7665);
or U10296 (N_10296,N_8698,N_8996);
xor U10297 (N_10297,N_6645,N_7838);
xnor U10298 (N_10298,N_8345,N_8341);
and U10299 (N_10299,N_8346,N_7341);
xor U10300 (N_10300,N_7758,N_7633);
nor U10301 (N_10301,N_6713,N_8892);
nand U10302 (N_10302,N_6266,N_6504);
or U10303 (N_10303,N_6895,N_8073);
or U10304 (N_10304,N_7722,N_8485);
nor U10305 (N_10305,N_7865,N_7160);
nor U10306 (N_10306,N_7615,N_8328);
nor U10307 (N_10307,N_8500,N_6415);
and U10308 (N_10308,N_7972,N_7213);
nor U10309 (N_10309,N_6552,N_8294);
or U10310 (N_10310,N_7875,N_7236);
nor U10311 (N_10311,N_8506,N_6283);
nand U10312 (N_10312,N_6349,N_8138);
nand U10313 (N_10313,N_6717,N_6610);
nand U10314 (N_10314,N_7074,N_6189);
or U10315 (N_10315,N_8508,N_7609);
nor U10316 (N_10316,N_6808,N_7357);
and U10317 (N_10317,N_7600,N_8126);
and U10318 (N_10318,N_6863,N_7052);
nand U10319 (N_10319,N_8631,N_8712);
nor U10320 (N_10320,N_7862,N_8896);
and U10321 (N_10321,N_6392,N_6428);
and U10322 (N_10322,N_7488,N_8675);
and U10323 (N_10323,N_6660,N_6696);
and U10324 (N_10324,N_8193,N_8332);
and U10325 (N_10325,N_7894,N_6339);
nor U10326 (N_10326,N_7399,N_7414);
nand U10327 (N_10327,N_6445,N_6236);
or U10328 (N_10328,N_8620,N_6473);
and U10329 (N_10329,N_6183,N_6841);
or U10330 (N_10330,N_8959,N_8974);
nor U10331 (N_10331,N_7015,N_6786);
nor U10332 (N_10332,N_7179,N_7315);
nor U10333 (N_10333,N_8725,N_6126);
or U10334 (N_10334,N_8075,N_8709);
nor U10335 (N_10335,N_6985,N_7340);
and U10336 (N_10336,N_8423,N_6883);
or U10337 (N_10337,N_8860,N_8691);
or U10338 (N_10338,N_7546,N_8643);
nor U10339 (N_10339,N_8197,N_7108);
and U10340 (N_10340,N_8123,N_6864);
nand U10341 (N_10341,N_7338,N_8676);
nor U10342 (N_10342,N_6546,N_7241);
or U10343 (N_10343,N_7628,N_7087);
nand U10344 (N_10344,N_6402,N_7647);
nand U10345 (N_10345,N_6230,N_6727);
nand U10346 (N_10346,N_8920,N_6272);
nor U10347 (N_10347,N_6915,N_6658);
nand U10348 (N_10348,N_7605,N_7210);
xnor U10349 (N_10349,N_7376,N_6059);
or U10350 (N_10350,N_6448,N_6244);
or U10351 (N_10351,N_8166,N_8416);
nand U10352 (N_10352,N_6661,N_7298);
nand U10353 (N_10353,N_6245,N_7683);
or U10354 (N_10354,N_6650,N_6125);
and U10355 (N_10355,N_8424,N_8010);
and U10356 (N_10356,N_6627,N_6814);
nor U10357 (N_10357,N_6291,N_6149);
nor U10358 (N_10358,N_7286,N_7941);
xor U10359 (N_10359,N_8085,N_6940);
nor U10360 (N_10360,N_8652,N_7334);
and U10361 (N_10361,N_6027,N_8940);
nor U10362 (N_10362,N_8205,N_7777);
or U10363 (N_10363,N_7063,N_8678);
and U10364 (N_10364,N_8235,N_8484);
nand U10365 (N_10365,N_8890,N_6875);
nand U10366 (N_10366,N_6967,N_6148);
or U10367 (N_10367,N_7839,N_8763);
or U10368 (N_10368,N_6484,N_8979);
xor U10369 (N_10369,N_8787,N_8482);
or U10370 (N_10370,N_6111,N_7814);
nand U10371 (N_10371,N_6481,N_6776);
and U10372 (N_10372,N_6302,N_7943);
nor U10373 (N_10373,N_8545,N_8851);
nor U10374 (N_10374,N_7644,N_7987);
nor U10375 (N_10375,N_8190,N_6948);
and U10376 (N_10376,N_7047,N_7288);
nor U10377 (N_10377,N_8985,N_6780);
nor U10378 (N_10378,N_6241,N_7652);
and U10379 (N_10379,N_6367,N_6414);
nor U10380 (N_10380,N_7701,N_8721);
nand U10381 (N_10381,N_8168,N_8414);
and U10382 (N_10382,N_7911,N_6753);
and U10383 (N_10383,N_6123,N_8791);
and U10384 (N_10384,N_6975,N_8005);
nand U10385 (N_10385,N_7115,N_7229);
and U10386 (N_10386,N_7120,N_6420);
or U10387 (N_10387,N_8287,N_7737);
xnor U10388 (N_10388,N_8467,N_8070);
nor U10389 (N_10389,N_7802,N_7936);
and U10390 (N_10390,N_6254,N_6901);
and U10391 (N_10391,N_6723,N_8157);
nand U10392 (N_10392,N_8934,N_7266);
xnor U10393 (N_10393,N_6775,N_8331);
nor U10394 (N_10394,N_8930,N_8616);
and U10395 (N_10395,N_7049,N_6670);
nand U10396 (N_10396,N_8589,N_7016);
or U10397 (N_10397,N_7720,N_8556);
nor U10398 (N_10398,N_6072,N_6172);
nand U10399 (N_10399,N_8640,N_8552);
nand U10400 (N_10400,N_8646,N_8130);
nand U10401 (N_10401,N_6992,N_6399);
xnor U10402 (N_10402,N_6639,N_7003);
nor U10403 (N_10403,N_8062,N_8260);
or U10404 (N_10404,N_7826,N_8442);
nand U10405 (N_10405,N_8523,N_7264);
or U10406 (N_10406,N_7985,N_6238);
and U10407 (N_10407,N_7312,N_7822);
nand U10408 (N_10408,N_7723,N_6074);
xnor U10409 (N_10409,N_7810,N_7712);
or U10410 (N_10410,N_7219,N_6762);
nand U10411 (N_10411,N_8876,N_8444);
and U10412 (N_10412,N_7924,N_8486);
or U10413 (N_10413,N_8367,N_6350);
and U10414 (N_10414,N_7212,N_8261);
and U10415 (N_10415,N_6213,N_7515);
nand U10416 (N_10416,N_7448,N_7589);
nor U10417 (N_10417,N_8938,N_7378);
nor U10418 (N_10418,N_6014,N_8828);
xnor U10419 (N_10419,N_8251,N_6739);
or U10420 (N_10420,N_6157,N_8932);
nor U10421 (N_10421,N_7776,N_6396);
and U10422 (N_10422,N_7498,N_7573);
and U10423 (N_10423,N_6654,N_8240);
or U10424 (N_10424,N_7146,N_7124);
nand U10425 (N_10425,N_8898,N_8008);
or U10426 (N_10426,N_6802,N_7271);
xor U10427 (N_10427,N_8487,N_6787);
nor U10428 (N_10428,N_6746,N_8634);
and U10429 (N_10429,N_6785,N_6434);
nand U10430 (N_10430,N_8858,N_6158);
or U10431 (N_10431,N_6376,N_6573);
nor U10432 (N_10432,N_6810,N_7168);
and U10433 (N_10433,N_8198,N_7349);
or U10434 (N_10434,N_6672,N_6364);
or U10435 (N_10435,N_6090,N_8163);
and U10436 (N_10436,N_6919,N_8064);
or U10437 (N_10437,N_8922,N_6363);
nor U10438 (N_10438,N_6134,N_7421);
and U10439 (N_10439,N_8671,N_8982);
and U10440 (N_10440,N_8921,N_8632);
nand U10441 (N_10441,N_6329,N_6882);
nor U10442 (N_10442,N_7207,N_6596);
nand U10443 (N_10443,N_8185,N_8021);
and U10444 (N_10444,N_7194,N_6413);
xor U10445 (N_10445,N_7863,N_6179);
nand U10446 (N_10446,N_6487,N_7547);
and U10447 (N_10447,N_7131,N_6947);
xnor U10448 (N_10448,N_6242,N_6640);
and U10449 (N_10449,N_8047,N_7691);
nand U10450 (N_10450,N_7174,N_7892);
nor U10451 (N_10451,N_7064,N_7586);
nor U10452 (N_10452,N_8203,N_8446);
nor U10453 (N_10453,N_7244,N_6873);
nor U10454 (N_10454,N_6115,N_7614);
or U10455 (N_10455,N_6447,N_6788);
or U10456 (N_10456,N_6561,N_6789);
nand U10457 (N_10457,N_8150,N_8382);
nor U10458 (N_10458,N_6061,N_7270);
nand U10459 (N_10459,N_8109,N_6950);
nor U10460 (N_10460,N_6698,N_6760);
or U10461 (N_10461,N_6614,N_6249);
or U10462 (N_10462,N_8980,N_8146);
and U10463 (N_10463,N_8337,N_8404);
xor U10464 (N_10464,N_8301,N_8649);
nand U10465 (N_10465,N_8154,N_6163);
nand U10466 (N_10466,N_6021,N_8740);
or U10467 (N_10467,N_7085,N_8088);
or U10468 (N_10468,N_7931,N_8027);
and U10469 (N_10469,N_6177,N_7417);
nor U10470 (N_10470,N_8751,N_7296);
or U10471 (N_10471,N_7066,N_8919);
or U10472 (N_10472,N_8087,N_8183);
nor U10473 (N_10473,N_6554,N_8507);
and U10474 (N_10474,N_8548,N_7117);
xor U10475 (N_10475,N_6777,N_6211);
xnor U10476 (N_10476,N_7598,N_6927);
nand U10477 (N_10477,N_8799,N_6924);
nor U10478 (N_10478,N_7734,N_6295);
and U10479 (N_10479,N_7307,N_8501);
nand U10480 (N_10480,N_7310,N_6889);
nor U10481 (N_10481,N_8479,N_7000);
nand U10482 (N_10482,N_6744,N_6381);
nor U10483 (N_10483,N_6833,N_8462);
nor U10484 (N_10484,N_6704,N_8107);
or U10485 (N_10485,N_8893,N_7048);
nor U10486 (N_10486,N_6656,N_7457);
nand U10487 (N_10487,N_7866,N_8089);
nand U10488 (N_10488,N_8090,N_8402);
nor U10489 (N_10489,N_6625,N_7159);
or U10490 (N_10490,N_7377,N_8526);
xor U10491 (N_10491,N_7745,N_7793);
or U10492 (N_10492,N_8020,N_7617);
nand U10493 (N_10493,N_6077,N_6716);
and U10494 (N_10494,N_8140,N_8499);
nor U10495 (N_10495,N_8910,N_8413);
or U10496 (N_10496,N_6161,N_6141);
nor U10497 (N_10497,N_6135,N_8177);
nand U10498 (N_10498,N_6751,N_8961);
or U10499 (N_10499,N_7796,N_8187);
nand U10500 (N_10500,N_7571,N_8028);
and U10501 (N_10501,N_7522,N_6638);
or U10502 (N_10502,N_6183,N_7777);
and U10503 (N_10503,N_7185,N_6158);
or U10504 (N_10504,N_8408,N_8312);
nor U10505 (N_10505,N_6244,N_8264);
and U10506 (N_10506,N_7790,N_6651);
nand U10507 (N_10507,N_8313,N_7067);
nor U10508 (N_10508,N_7530,N_8400);
or U10509 (N_10509,N_6821,N_6577);
nand U10510 (N_10510,N_6637,N_6854);
or U10511 (N_10511,N_8063,N_6535);
nand U10512 (N_10512,N_6595,N_7037);
nor U10513 (N_10513,N_7038,N_7956);
and U10514 (N_10514,N_8296,N_8485);
nand U10515 (N_10515,N_7340,N_8915);
xor U10516 (N_10516,N_8359,N_7312);
nand U10517 (N_10517,N_6730,N_7505);
nor U10518 (N_10518,N_8479,N_6457);
nand U10519 (N_10519,N_7547,N_6098);
or U10520 (N_10520,N_6769,N_7912);
or U10521 (N_10521,N_6931,N_6442);
or U10522 (N_10522,N_6777,N_6444);
xor U10523 (N_10523,N_7784,N_6466);
nand U10524 (N_10524,N_7068,N_6029);
nand U10525 (N_10525,N_7049,N_8488);
nor U10526 (N_10526,N_8603,N_6243);
or U10527 (N_10527,N_8562,N_7399);
nand U10528 (N_10528,N_8368,N_6304);
nand U10529 (N_10529,N_6152,N_7820);
and U10530 (N_10530,N_7567,N_8724);
and U10531 (N_10531,N_6484,N_6061);
nand U10532 (N_10532,N_7643,N_7980);
or U10533 (N_10533,N_6176,N_8288);
nand U10534 (N_10534,N_6212,N_8219);
nor U10535 (N_10535,N_6091,N_8553);
nor U10536 (N_10536,N_8406,N_7088);
or U10537 (N_10537,N_8610,N_6862);
nor U10538 (N_10538,N_6869,N_6408);
nor U10539 (N_10539,N_6740,N_8710);
or U10540 (N_10540,N_7456,N_7976);
and U10541 (N_10541,N_8611,N_8988);
or U10542 (N_10542,N_7230,N_7766);
or U10543 (N_10543,N_7321,N_7654);
and U10544 (N_10544,N_7995,N_6682);
nand U10545 (N_10545,N_8144,N_6431);
nor U10546 (N_10546,N_7843,N_7774);
nand U10547 (N_10547,N_8240,N_8135);
nor U10548 (N_10548,N_6057,N_8975);
xor U10549 (N_10549,N_6471,N_6804);
and U10550 (N_10550,N_8256,N_8767);
and U10551 (N_10551,N_6980,N_6228);
nor U10552 (N_10552,N_7979,N_8845);
nor U10553 (N_10553,N_8045,N_6313);
and U10554 (N_10554,N_6264,N_8510);
nand U10555 (N_10555,N_8741,N_8906);
and U10556 (N_10556,N_6331,N_6921);
or U10557 (N_10557,N_6036,N_7346);
and U10558 (N_10558,N_7681,N_8478);
or U10559 (N_10559,N_7047,N_6909);
and U10560 (N_10560,N_6422,N_7242);
nor U10561 (N_10561,N_7875,N_8058);
nand U10562 (N_10562,N_6198,N_7735);
or U10563 (N_10563,N_8844,N_6746);
nor U10564 (N_10564,N_6761,N_6698);
or U10565 (N_10565,N_6111,N_8317);
nand U10566 (N_10566,N_8097,N_7903);
nand U10567 (N_10567,N_8325,N_8409);
nand U10568 (N_10568,N_7734,N_6590);
nand U10569 (N_10569,N_8611,N_6419);
nand U10570 (N_10570,N_6608,N_6362);
or U10571 (N_10571,N_7406,N_6536);
or U10572 (N_10572,N_7566,N_8460);
xnor U10573 (N_10573,N_7085,N_6596);
and U10574 (N_10574,N_7411,N_8470);
nor U10575 (N_10575,N_6659,N_6251);
nor U10576 (N_10576,N_6444,N_7557);
xor U10577 (N_10577,N_6910,N_8454);
or U10578 (N_10578,N_7648,N_6992);
nor U10579 (N_10579,N_7962,N_7188);
nand U10580 (N_10580,N_8838,N_6865);
nand U10581 (N_10581,N_7228,N_8691);
and U10582 (N_10582,N_6336,N_8575);
or U10583 (N_10583,N_8507,N_8549);
xor U10584 (N_10584,N_8524,N_6329);
xnor U10585 (N_10585,N_6606,N_8336);
and U10586 (N_10586,N_7563,N_8563);
or U10587 (N_10587,N_7470,N_8533);
and U10588 (N_10588,N_6561,N_8813);
nor U10589 (N_10589,N_6775,N_8389);
and U10590 (N_10590,N_6808,N_7666);
nor U10591 (N_10591,N_6654,N_8367);
xor U10592 (N_10592,N_7569,N_7902);
xor U10593 (N_10593,N_6646,N_8688);
nor U10594 (N_10594,N_6180,N_7320);
and U10595 (N_10595,N_8460,N_6362);
nand U10596 (N_10596,N_7113,N_8353);
xor U10597 (N_10597,N_6026,N_7019);
nor U10598 (N_10598,N_7551,N_6389);
nand U10599 (N_10599,N_7625,N_8566);
and U10600 (N_10600,N_8687,N_7130);
nand U10601 (N_10601,N_6834,N_7661);
nor U10602 (N_10602,N_8742,N_8458);
nand U10603 (N_10603,N_6008,N_6511);
nor U10604 (N_10604,N_6874,N_6151);
nor U10605 (N_10605,N_8190,N_7920);
and U10606 (N_10606,N_8184,N_7217);
xnor U10607 (N_10607,N_6424,N_7953);
and U10608 (N_10608,N_6788,N_8841);
xor U10609 (N_10609,N_8502,N_7498);
and U10610 (N_10610,N_6506,N_8849);
or U10611 (N_10611,N_6312,N_6705);
or U10612 (N_10612,N_7735,N_8941);
nand U10613 (N_10613,N_8685,N_7395);
nand U10614 (N_10614,N_8698,N_6815);
nor U10615 (N_10615,N_7442,N_6345);
or U10616 (N_10616,N_8497,N_8408);
or U10617 (N_10617,N_8233,N_6964);
nand U10618 (N_10618,N_7564,N_6523);
nor U10619 (N_10619,N_7387,N_7113);
nor U10620 (N_10620,N_6333,N_6860);
or U10621 (N_10621,N_8034,N_7704);
xnor U10622 (N_10622,N_8872,N_8463);
nor U10623 (N_10623,N_8984,N_8241);
or U10624 (N_10624,N_6589,N_6407);
nor U10625 (N_10625,N_6756,N_7181);
nor U10626 (N_10626,N_6861,N_7078);
nor U10627 (N_10627,N_6502,N_7169);
xor U10628 (N_10628,N_8446,N_7729);
or U10629 (N_10629,N_6150,N_6794);
or U10630 (N_10630,N_6575,N_8118);
or U10631 (N_10631,N_7891,N_8085);
nor U10632 (N_10632,N_7269,N_8568);
nor U10633 (N_10633,N_8252,N_7550);
xor U10634 (N_10634,N_8381,N_7975);
or U10635 (N_10635,N_7666,N_8955);
or U10636 (N_10636,N_8341,N_8695);
nor U10637 (N_10637,N_7931,N_7710);
nor U10638 (N_10638,N_8421,N_6411);
xnor U10639 (N_10639,N_6028,N_8955);
nor U10640 (N_10640,N_8008,N_6395);
nor U10641 (N_10641,N_7978,N_6230);
nand U10642 (N_10642,N_7289,N_7104);
nand U10643 (N_10643,N_6222,N_6435);
xor U10644 (N_10644,N_6608,N_7688);
nand U10645 (N_10645,N_8638,N_6530);
xnor U10646 (N_10646,N_7093,N_7539);
or U10647 (N_10647,N_7688,N_6207);
xnor U10648 (N_10648,N_8727,N_6883);
nor U10649 (N_10649,N_6494,N_8637);
nor U10650 (N_10650,N_6638,N_8614);
nor U10651 (N_10651,N_6057,N_8358);
and U10652 (N_10652,N_8879,N_6521);
nand U10653 (N_10653,N_8773,N_7563);
xnor U10654 (N_10654,N_7987,N_6242);
or U10655 (N_10655,N_8893,N_6891);
or U10656 (N_10656,N_7132,N_8322);
nor U10657 (N_10657,N_8469,N_7903);
xnor U10658 (N_10658,N_8336,N_6974);
and U10659 (N_10659,N_7477,N_7350);
nand U10660 (N_10660,N_6972,N_8131);
nor U10661 (N_10661,N_6825,N_8359);
and U10662 (N_10662,N_6898,N_7231);
and U10663 (N_10663,N_8594,N_7089);
nand U10664 (N_10664,N_7495,N_7629);
nand U10665 (N_10665,N_8263,N_6502);
and U10666 (N_10666,N_8284,N_7304);
xor U10667 (N_10667,N_6144,N_8372);
and U10668 (N_10668,N_8690,N_8088);
or U10669 (N_10669,N_8895,N_6406);
or U10670 (N_10670,N_8706,N_8094);
or U10671 (N_10671,N_8307,N_8185);
and U10672 (N_10672,N_6464,N_6401);
xnor U10673 (N_10673,N_6860,N_7417);
and U10674 (N_10674,N_7092,N_8508);
and U10675 (N_10675,N_8008,N_7250);
nand U10676 (N_10676,N_6834,N_6247);
or U10677 (N_10677,N_8221,N_6988);
nand U10678 (N_10678,N_8236,N_6435);
and U10679 (N_10679,N_8153,N_7327);
nor U10680 (N_10680,N_6528,N_6054);
or U10681 (N_10681,N_6740,N_6078);
and U10682 (N_10682,N_6677,N_6761);
or U10683 (N_10683,N_7317,N_8869);
xnor U10684 (N_10684,N_6669,N_6361);
and U10685 (N_10685,N_7165,N_7176);
nand U10686 (N_10686,N_7336,N_6588);
nor U10687 (N_10687,N_7425,N_8716);
nand U10688 (N_10688,N_8369,N_6341);
or U10689 (N_10689,N_7241,N_8735);
nor U10690 (N_10690,N_6326,N_8587);
and U10691 (N_10691,N_8666,N_7918);
and U10692 (N_10692,N_7870,N_8854);
nor U10693 (N_10693,N_8756,N_8218);
nor U10694 (N_10694,N_8819,N_6023);
nand U10695 (N_10695,N_6246,N_6699);
or U10696 (N_10696,N_8666,N_6078);
or U10697 (N_10697,N_8825,N_6020);
nand U10698 (N_10698,N_8585,N_8058);
nand U10699 (N_10699,N_8297,N_8303);
nand U10700 (N_10700,N_6728,N_7624);
or U10701 (N_10701,N_6708,N_6053);
nor U10702 (N_10702,N_8242,N_6856);
nand U10703 (N_10703,N_7589,N_8232);
or U10704 (N_10704,N_7625,N_7559);
nor U10705 (N_10705,N_8689,N_8922);
and U10706 (N_10706,N_6223,N_7183);
and U10707 (N_10707,N_8762,N_6021);
nand U10708 (N_10708,N_7762,N_6767);
nor U10709 (N_10709,N_6172,N_8163);
nor U10710 (N_10710,N_7635,N_8281);
nor U10711 (N_10711,N_8732,N_7609);
nor U10712 (N_10712,N_8700,N_6894);
and U10713 (N_10713,N_7522,N_8222);
nand U10714 (N_10714,N_8375,N_6884);
nor U10715 (N_10715,N_7737,N_7618);
nor U10716 (N_10716,N_8470,N_6101);
xnor U10717 (N_10717,N_6166,N_6552);
nor U10718 (N_10718,N_7848,N_7724);
nor U10719 (N_10719,N_8878,N_8669);
and U10720 (N_10720,N_6131,N_7657);
nor U10721 (N_10721,N_7570,N_8571);
nor U10722 (N_10722,N_8545,N_7264);
nor U10723 (N_10723,N_8689,N_6486);
nor U10724 (N_10724,N_6396,N_7870);
nand U10725 (N_10725,N_8180,N_8040);
nand U10726 (N_10726,N_8704,N_6133);
and U10727 (N_10727,N_7054,N_8501);
and U10728 (N_10728,N_7769,N_8568);
xor U10729 (N_10729,N_6720,N_7712);
or U10730 (N_10730,N_7249,N_6498);
xor U10731 (N_10731,N_7172,N_8237);
and U10732 (N_10732,N_7522,N_6895);
nand U10733 (N_10733,N_8768,N_7850);
nand U10734 (N_10734,N_7176,N_7261);
nor U10735 (N_10735,N_6581,N_6245);
or U10736 (N_10736,N_7566,N_6970);
nor U10737 (N_10737,N_8471,N_6915);
nand U10738 (N_10738,N_7806,N_6289);
nand U10739 (N_10739,N_6170,N_6957);
nor U10740 (N_10740,N_6585,N_8669);
nand U10741 (N_10741,N_6928,N_8056);
or U10742 (N_10742,N_6226,N_6180);
and U10743 (N_10743,N_8467,N_6572);
nand U10744 (N_10744,N_6357,N_8475);
nor U10745 (N_10745,N_7343,N_6938);
xnor U10746 (N_10746,N_8461,N_6126);
or U10747 (N_10747,N_7223,N_6053);
nand U10748 (N_10748,N_8055,N_7425);
and U10749 (N_10749,N_6395,N_6552);
nand U10750 (N_10750,N_6176,N_7501);
or U10751 (N_10751,N_7602,N_7994);
nand U10752 (N_10752,N_8123,N_7063);
nand U10753 (N_10753,N_8739,N_6849);
nand U10754 (N_10754,N_6120,N_6082);
nand U10755 (N_10755,N_6865,N_7140);
and U10756 (N_10756,N_7655,N_6315);
and U10757 (N_10757,N_7074,N_8920);
or U10758 (N_10758,N_7619,N_6582);
and U10759 (N_10759,N_8091,N_6831);
or U10760 (N_10760,N_8018,N_7794);
or U10761 (N_10761,N_8839,N_8669);
or U10762 (N_10762,N_7865,N_8989);
and U10763 (N_10763,N_7083,N_8225);
and U10764 (N_10764,N_6531,N_8432);
and U10765 (N_10765,N_6746,N_6796);
and U10766 (N_10766,N_6932,N_8994);
nand U10767 (N_10767,N_7088,N_7600);
and U10768 (N_10768,N_7842,N_7496);
or U10769 (N_10769,N_8891,N_7697);
nor U10770 (N_10770,N_6849,N_6186);
xnor U10771 (N_10771,N_8994,N_8426);
nor U10772 (N_10772,N_7491,N_7425);
nand U10773 (N_10773,N_7489,N_6971);
xor U10774 (N_10774,N_6554,N_7058);
nor U10775 (N_10775,N_6036,N_8566);
or U10776 (N_10776,N_8747,N_8333);
nor U10777 (N_10777,N_8669,N_8507);
and U10778 (N_10778,N_7553,N_7982);
nor U10779 (N_10779,N_6954,N_6787);
nor U10780 (N_10780,N_6279,N_6875);
and U10781 (N_10781,N_7258,N_7843);
xnor U10782 (N_10782,N_7045,N_6805);
and U10783 (N_10783,N_7400,N_8461);
xor U10784 (N_10784,N_7905,N_8294);
nor U10785 (N_10785,N_6122,N_7399);
nand U10786 (N_10786,N_8757,N_8323);
nand U10787 (N_10787,N_7058,N_6060);
nand U10788 (N_10788,N_8516,N_8635);
and U10789 (N_10789,N_8247,N_7491);
nand U10790 (N_10790,N_7386,N_6619);
nand U10791 (N_10791,N_8241,N_7054);
nand U10792 (N_10792,N_6765,N_8336);
or U10793 (N_10793,N_6737,N_6548);
or U10794 (N_10794,N_7697,N_8499);
nand U10795 (N_10795,N_8481,N_7446);
nand U10796 (N_10796,N_8448,N_6360);
nor U10797 (N_10797,N_8921,N_8619);
nand U10798 (N_10798,N_8206,N_8659);
nor U10799 (N_10799,N_6046,N_8267);
and U10800 (N_10800,N_6053,N_6186);
or U10801 (N_10801,N_8873,N_8336);
nor U10802 (N_10802,N_8563,N_6326);
nor U10803 (N_10803,N_7608,N_8793);
or U10804 (N_10804,N_6540,N_7839);
nor U10805 (N_10805,N_6666,N_7144);
nand U10806 (N_10806,N_6533,N_6250);
nand U10807 (N_10807,N_6603,N_6685);
and U10808 (N_10808,N_6151,N_6639);
and U10809 (N_10809,N_8876,N_8152);
nor U10810 (N_10810,N_7108,N_8674);
nand U10811 (N_10811,N_7275,N_8249);
nand U10812 (N_10812,N_7462,N_6556);
and U10813 (N_10813,N_7560,N_7496);
nand U10814 (N_10814,N_8692,N_7574);
xnor U10815 (N_10815,N_6714,N_7821);
or U10816 (N_10816,N_7010,N_7988);
or U10817 (N_10817,N_8678,N_6050);
nor U10818 (N_10818,N_6336,N_7335);
or U10819 (N_10819,N_7458,N_8454);
and U10820 (N_10820,N_7068,N_8227);
xnor U10821 (N_10821,N_7997,N_8479);
or U10822 (N_10822,N_6565,N_6158);
nor U10823 (N_10823,N_6254,N_7879);
nor U10824 (N_10824,N_8784,N_8343);
or U10825 (N_10825,N_8985,N_7574);
nor U10826 (N_10826,N_7868,N_6041);
xor U10827 (N_10827,N_6401,N_6903);
xor U10828 (N_10828,N_6056,N_8707);
or U10829 (N_10829,N_8615,N_6793);
nor U10830 (N_10830,N_7712,N_6721);
nand U10831 (N_10831,N_7787,N_6232);
nand U10832 (N_10832,N_6691,N_8797);
and U10833 (N_10833,N_8371,N_6746);
or U10834 (N_10834,N_6049,N_8964);
nor U10835 (N_10835,N_7564,N_8066);
and U10836 (N_10836,N_7183,N_7827);
nand U10837 (N_10837,N_6969,N_8367);
nand U10838 (N_10838,N_8843,N_8425);
and U10839 (N_10839,N_8193,N_7916);
nor U10840 (N_10840,N_8121,N_7154);
and U10841 (N_10841,N_7062,N_7957);
nand U10842 (N_10842,N_8072,N_6698);
and U10843 (N_10843,N_7237,N_7967);
xnor U10844 (N_10844,N_7551,N_7349);
nand U10845 (N_10845,N_7989,N_6737);
and U10846 (N_10846,N_8917,N_8049);
or U10847 (N_10847,N_7987,N_7660);
or U10848 (N_10848,N_6337,N_7752);
xnor U10849 (N_10849,N_6465,N_7756);
nand U10850 (N_10850,N_7407,N_7121);
and U10851 (N_10851,N_6538,N_7001);
or U10852 (N_10852,N_6742,N_7401);
or U10853 (N_10853,N_6848,N_8607);
or U10854 (N_10854,N_8136,N_7798);
nor U10855 (N_10855,N_7188,N_8437);
nand U10856 (N_10856,N_8358,N_8224);
nand U10857 (N_10857,N_6891,N_8532);
or U10858 (N_10858,N_8181,N_8579);
nand U10859 (N_10859,N_7320,N_7875);
xor U10860 (N_10860,N_8462,N_6639);
xor U10861 (N_10861,N_6661,N_8941);
nand U10862 (N_10862,N_7602,N_6584);
nand U10863 (N_10863,N_7473,N_8453);
nor U10864 (N_10864,N_6501,N_7059);
nand U10865 (N_10865,N_7857,N_6426);
xnor U10866 (N_10866,N_8123,N_8952);
or U10867 (N_10867,N_6727,N_8088);
and U10868 (N_10868,N_8929,N_7325);
or U10869 (N_10869,N_8396,N_6597);
nand U10870 (N_10870,N_6055,N_6326);
or U10871 (N_10871,N_7669,N_6875);
and U10872 (N_10872,N_8183,N_6006);
nand U10873 (N_10873,N_8341,N_8066);
nor U10874 (N_10874,N_8191,N_6008);
or U10875 (N_10875,N_8557,N_8514);
or U10876 (N_10876,N_6867,N_8977);
or U10877 (N_10877,N_8480,N_7017);
nand U10878 (N_10878,N_7558,N_8370);
nand U10879 (N_10879,N_7066,N_7262);
nand U10880 (N_10880,N_6113,N_6768);
and U10881 (N_10881,N_8512,N_6847);
nand U10882 (N_10882,N_7096,N_7572);
or U10883 (N_10883,N_6370,N_7079);
nand U10884 (N_10884,N_7016,N_8084);
nand U10885 (N_10885,N_6338,N_7974);
or U10886 (N_10886,N_8785,N_8469);
nand U10887 (N_10887,N_7795,N_7080);
or U10888 (N_10888,N_6624,N_7132);
or U10889 (N_10889,N_8439,N_8490);
and U10890 (N_10890,N_8342,N_7653);
nor U10891 (N_10891,N_7791,N_7519);
nand U10892 (N_10892,N_6275,N_8657);
and U10893 (N_10893,N_8193,N_6393);
nand U10894 (N_10894,N_8428,N_8694);
or U10895 (N_10895,N_7563,N_7833);
and U10896 (N_10896,N_8246,N_8167);
nand U10897 (N_10897,N_7610,N_6486);
or U10898 (N_10898,N_7458,N_7062);
nand U10899 (N_10899,N_6774,N_6649);
nand U10900 (N_10900,N_7274,N_6491);
or U10901 (N_10901,N_6536,N_8922);
and U10902 (N_10902,N_8929,N_6044);
nor U10903 (N_10903,N_7226,N_7702);
xor U10904 (N_10904,N_6383,N_8065);
nand U10905 (N_10905,N_7469,N_6272);
or U10906 (N_10906,N_8943,N_6238);
or U10907 (N_10907,N_8016,N_6930);
nand U10908 (N_10908,N_6357,N_8133);
nand U10909 (N_10909,N_6114,N_8509);
nor U10910 (N_10910,N_8065,N_8191);
and U10911 (N_10911,N_6684,N_7293);
nand U10912 (N_10912,N_6436,N_7564);
or U10913 (N_10913,N_6821,N_6362);
nor U10914 (N_10914,N_8128,N_7420);
nand U10915 (N_10915,N_8346,N_8639);
nor U10916 (N_10916,N_7641,N_7935);
nor U10917 (N_10917,N_6428,N_6137);
nor U10918 (N_10918,N_6764,N_8228);
nand U10919 (N_10919,N_6551,N_8716);
xnor U10920 (N_10920,N_6768,N_7399);
and U10921 (N_10921,N_8164,N_8730);
or U10922 (N_10922,N_6760,N_6575);
or U10923 (N_10923,N_8509,N_8028);
nor U10924 (N_10924,N_8214,N_6102);
and U10925 (N_10925,N_7143,N_6968);
nand U10926 (N_10926,N_7138,N_6889);
nor U10927 (N_10927,N_7728,N_6376);
nor U10928 (N_10928,N_6011,N_6394);
and U10929 (N_10929,N_7088,N_6822);
and U10930 (N_10930,N_8141,N_6423);
nor U10931 (N_10931,N_6682,N_8955);
nand U10932 (N_10932,N_6493,N_6879);
or U10933 (N_10933,N_8472,N_7855);
nand U10934 (N_10934,N_8247,N_7157);
or U10935 (N_10935,N_7058,N_8153);
nand U10936 (N_10936,N_7775,N_7008);
nor U10937 (N_10937,N_8238,N_6180);
or U10938 (N_10938,N_7837,N_8226);
nor U10939 (N_10939,N_7252,N_7116);
nand U10940 (N_10940,N_8225,N_7584);
nor U10941 (N_10941,N_6483,N_6814);
nor U10942 (N_10942,N_6831,N_8991);
or U10943 (N_10943,N_8996,N_7691);
or U10944 (N_10944,N_7191,N_7662);
nor U10945 (N_10945,N_7661,N_6491);
and U10946 (N_10946,N_6298,N_6837);
nor U10947 (N_10947,N_6336,N_6805);
nor U10948 (N_10948,N_7923,N_6761);
and U10949 (N_10949,N_6997,N_7062);
and U10950 (N_10950,N_8173,N_8474);
nand U10951 (N_10951,N_6216,N_6712);
nor U10952 (N_10952,N_6901,N_6728);
or U10953 (N_10953,N_8546,N_7311);
nand U10954 (N_10954,N_6462,N_6549);
nor U10955 (N_10955,N_6102,N_7228);
or U10956 (N_10956,N_8673,N_8932);
and U10957 (N_10957,N_6973,N_8928);
nand U10958 (N_10958,N_8586,N_7368);
nor U10959 (N_10959,N_7917,N_6436);
and U10960 (N_10960,N_7760,N_6995);
nor U10961 (N_10961,N_6771,N_8312);
nor U10962 (N_10962,N_7371,N_8797);
or U10963 (N_10963,N_8296,N_6276);
or U10964 (N_10964,N_7637,N_6166);
xnor U10965 (N_10965,N_8966,N_7968);
or U10966 (N_10966,N_7029,N_7547);
nand U10967 (N_10967,N_7275,N_8952);
nor U10968 (N_10968,N_8744,N_8814);
and U10969 (N_10969,N_6905,N_8844);
nor U10970 (N_10970,N_8784,N_7840);
or U10971 (N_10971,N_6245,N_8850);
or U10972 (N_10972,N_7024,N_6414);
or U10973 (N_10973,N_8691,N_8111);
or U10974 (N_10974,N_7046,N_8676);
nand U10975 (N_10975,N_8447,N_8064);
nand U10976 (N_10976,N_6452,N_8523);
nand U10977 (N_10977,N_8470,N_7339);
nand U10978 (N_10978,N_7330,N_6876);
xnor U10979 (N_10979,N_8555,N_6660);
or U10980 (N_10980,N_8524,N_6758);
or U10981 (N_10981,N_7377,N_7152);
and U10982 (N_10982,N_7557,N_7630);
nand U10983 (N_10983,N_6245,N_8986);
nand U10984 (N_10984,N_6146,N_8314);
nand U10985 (N_10985,N_8543,N_6094);
nor U10986 (N_10986,N_6746,N_6635);
and U10987 (N_10987,N_6146,N_6906);
nand U10988 (N_10988,N_8456,N_8062);
or U10989 (N_10989,N_8196,N_6921);
or U10990 (N_10990,N_8334,N_6537);
nand U10991 (N_10991,N_7015,N_7065);
or U10992 (N_10992,N_8793,N_7201);
nand U10993 (N_10993,N_6647,N_6461);
or U10994 (N_10994,N_8448,N_7672);
and U10995 (N_10995,N_8802,N_8428);
nand U10996 (N_10996,N_8353,N_8216);
nor U10997 (N_10997,N_6790,N_8122);
nor U10998 (N_10998,N_6227,N_6488);
nor U10999 (N_10999,N_7232,N_7537);
or U11000 (N_11000,N_8426,N_8827);
nor U11001 (N_11001,N_8320,N_8595);
or U11002 (N_11002,N_8507,N_6894);
nand U11003 (N_11003,N_8244,N_8051);
nand U11004 (N_11004,N_7655,N_8301);
or U11005 (N_11005,N_8933,N_8648);
and U11006 (N_11006,N_8308,N_6004);
nor U11007 (N_11007,N_8552,N_6233);
and U11008 (N_11008,N_7614,N_7203);
nand U11009 (N_11009,N_6937,N_6417);
nor U11010 (N_11010,N_6804,N_8051);
and U11011 (N_11011,N_7874,N_8826);
or U11012 (N_11012,N_6765,N_6116);
or U11013 (N_11013,N_7954,N_7851);
nand U11014 (N_11014,N_8598,N_6471);
nor U11015 (N_11015,N_6038,N_6291);
or U11016 (N_11016,N_7148,N_6807);
nand U11017 (N_11017,N_7085,N_6392);
nand U11018 (N_11018,N_6752,N_6076);
nor U11019 (N_11019,N_8531,N_8468);
and U11020 (N_11020,N_8247,N_7924);
or U11021 (N_11021,N_7785,N_8958);
xor U11022 (N_11022,N_7229,N_7584);
and U11023 (N_11023,N_6560,N_7791);
nand U11024 (N_11024,N_6207,N_7683);
nor U11025 (N_11025,N_6338,N_7809);
nor U11026 (N_11026,N_8808,N_6619);
nand U11027 (N_11027,N_7071,N_8725);
nor U11028 (N_11028,N_8874,N_8550);
nand U11029 (N_11029,N_7977,N_7744);
nor U11030 (N_11030,N_8707,N_6044);
nand U11031 (N_11031,N_8393,N_7507);
or U11032 (N_11032,N_6564,N_7140);
nand U11033 (N_11033,N_6641,N_8123);
and U11034 (N_11034,N_7350,N_8544);
or U11035 (N_11035,N_8831,N_8785);
or U11036 (N_11036,N_7336,N_6601);
and U11037 (N_11037,N_6221,N_7741);
nand U11038 (N_11038,N_6534,N_7580);
and U11039 (N_11039,N_7754,N_7001);
nor U11040 (N_11040,N_6024,N_8031);
nand U11041 (N_11041,N_8356,N_8481);
nor U11042 (N_11042,N_7524,N_6881);
and U11043 (N_11043,N_8062,N_7865);
nand U11044 (N_11044,N_8418,N_8873);
or U11045 (N_11045,N_6440,N_8899);
nor U11046 (N_11046,N_8746,N_7652);
nand U11047 (N_11047,N_8185,N_6171);
xnor U11048 (N_11048,N_6817,N_7947);
nor U11049 (N_11049,N_8413,N_7907);
or U11050 (N_11050,N_7423,N_7542);
or U11051 (N_11051,N_6380,N_7999);
or U11052 (N_11052,N_8886,N_7745);
and U11053 (N_11053,N_8665,N_7889);
or U11054 (N_11054,N_7585,N_7545);
or U11055 (N_11055,N_8537,N_8321);
xor U11056 (N_11056,N_8464,N_7126);
xor U11057 (N_11057,N_8686,N_6528);
and U11058 (N_11058,N_8173,N_6715);
or U11059 (N_11059,N_7195,N_6876);
nand U11060 (N_11060,N_8268,N_7276);
nand U11061 (N_11061,N_6096,N_6628);
nor U11062 (N_11062,N_7952,N_7200);
or U11063 (N_11063,N_6571,N_8141);
or U11064 (N_11064,N_6636,N_8713);
and U11065 (N_11065,N_7852,N_8312);
nor U11066 (N_11066,N_6173,N_7647);
nand U11067 (N_11067,N_7172,N_7933);
nor U11068 (N_11068,N_6797,N_6338);
or U11069 (N_11069,N_8404,N_8873);
nor U11070 (N_11070,N_6403,N_6723);
and U11071 (N_11071,N_6308,N_8673);
nor U11072 (N_11072,N_6150,N_6376);
nor U11073 (N_11073,N_8044,N_6057);
or U11074 (N_11074,N_7533,N_8414);
xor U11075 (N_11075,N_8198,N_6186);
and U11076 (N_11076,N_8275,N_6157);
and U11077 (N_11077,N_7031,N_7650);
nand U11078 (N_11078,N_8073,N_6592);
xnor U11079 (N_11079,N_6978,N_7252);
or U11080 (N_11080,N_6938,N_8104);
or U11081 (N_11081,N_6768,N_6571);
nand U11082 (N_11082,N_6711,N_6113);
nor U11083 (N_11083,N_6944,N_8380);
and U11084 (N_11084,N_6826,N_6784);
xnor U11085 (N_11085,N_8545,N_6517);
and U11086 (N_11086,N_8264,N_7118);
nor U11087 (N_11087,N_8636,N_6038);
xor U11088 (N_11088,N_7208,N_8044);
nand U11089 (N_11089,N_6690,N_6578);
nor U11090 (N_11090,N_7329,N_7249);
nor U11091 (N_11091,N_7924,N_8346);
and U11092 (N_11092,N_7107,N_8854);
or U11093 (N_11093,N_7125,N_7013);
and U11094 (N_11094,N_8029,N_8302);
or U11095 (N_11095,N_8497,N_7534);
nor U11096 (N_11096,N_6597,N_6432);
nand U11097 (N_11097,N_8385,N_6146);
nor U11098 (N_11098,N_8118,N_8945);
nand U11099 (N_11099,N_7255,N_6825);
nand U11100 (N_11100,N_7865,N_8484);
and U11101 (N_11101,N_6361,N_7838);
and U11102 (N_11102,N_8209,N_6550);
or U11103 (N_11103,N_6142,N_7982);
or U11104 (N_11104,N_6377,N_8424);
nor U11105 (N_11105,N_8483,N_8807);
nor U11106 (N_11106,N_7141,N_8368);
nand U11107 (N_11107,N_8479,N_7283);
nor U11108 (N_11108,N_8243,N_7415);
nor U11109 (N_11109,N_7316,N_8925);
nor U11110 (N_11110,N_7487,N_6844);
xor U11111 (N_11111,N_6214,N_7169);
nor U11112 (N_11112,N_8488,N_8119);
nand U11113 (N_11113,N_6027,N_6278);
nor U11114 (N_11114,N_6719,N_8360);
or U11115 (N_11115,N_7372,N_7140);
nor U11116 (N_11116,N_6233,N_8597);
nand U11117 (N_11117,N_6619,N_8637);
and U11118 (N_11118,N_7606,N_8744);
nor U11119 (N_11119,N_7282,N_8224);
nor U11120 (N_11120,N_6160,N_8278);
nor U11121 (N_11121,N_6767,N_8131);
nor U11122 (N_11122,N_6875,N_8156);
and U11123 (N_11123,N_7906,N_6875);
and U11124 (N_11124,N_6271,N_6741);
or U11125 (N_11125,N_6330,N_6543);
or U11126 (N_11126,N_6565,N_6547);
nor U11127 (N_11127,N_6341,N_7189);
xor U11128 (N_11128,N_7780,N_7932);
and U11129 (N_11129,N_7542,N_8522);
nand U11130 (N_11130,N_7479,N_6388);
nand U11131 (N_11131,N_7282,N_6559);
xnor U11132 (N_11132,N_7899,N_6348);
or U11133 (N_11133,N_7799,N_8524);
xnor U11134 (N_11134,N_8212,N_6868);
nor U11135 (N_11135,N_6581,N_8242);
or U11136 (N_11136,N_8912,N_8606);
and U11137 (N_11137,N_6797,N_6426);
nand U11138 (N_11138,N_7001,N_6373);
nor U11139 (N_11139,N_7867,N_8013);
or U11140 (N_11140,N_6138,N_6035);
or U11141 (N_11141,N_8113,N_8679);
nor U11142 (N_11142,N_7503,N_7083);
nor U11143 (N_11143,N_6019,N_8935);
or U11144 (N_11144,N_6788,N_7709);
or U11145 (N_11145,N_7523,N_7701);
nor U11146 (N_11146,N_8797,N_6624);
or U11147 (N_11147,N_8157,N_7731);
or U11148 (N_11148,N_8447,N_7805);
nor U11149 (N_11149,N_8097,N_6834);
nand U11150 (N_11150,N_6633,N_6296);
or U11151 (N_11151,N_7885,N_6066);
nor U11152 (N_11152,N_7384,N_6180);
nor U11153 (N_11153,N_6137,N_7536);
nand U11154 (N_11154,N_8120,N_6765);
nor U11155 (N_11155,N_7288,N_6526);
and U11156 (N_11156,N_7327,N_6822);
and U11157 (N_11157,N_7267,N_8568);
or U11158 (N_11158,N_8005,N_6025);
nor U11159 (N_11159,N_8629,N_8925);
or U11160 (N_11160,N_6032,N_6631);
nor U11161 (N_11161,N_8828,N_7671);
or U11162 (N_11162,N_8952,N_8396);
nor U11163 (N_11163,N_7574,N_7134);
nor U11164 (N_11164,N_8429,N_7899);
and U11165 (N_11165,N_7948,N_7325);
and U11166 (N_11166,N_7358,N_7076);
and U11167 (N_11167,N_8578,N_8176);
and U11168 (N_11168,N_8409,N_8028);
and U11169 (N_11169,N_7417,N_7360);
nand U11170 (N_11170,N_7369,N_7558);
or U11171 (N_11171,N_6901,N_7046);
nor U11172 (N_11172,N_7397,N_6060);
nor U11173 (N_11173,N_6141,N_6429);
or U11174 (N_11174,N_6851,N_6687);
nor U11175 (N_11175,N_6460,N_6881);
xnor U11176 (N_11176,N_8609,N_6235);
or U11177 (N_11177,N_8387,N_8345);
xnor U11178 (N_11178,N_6180,N_7284);
nor U11179 (N_11179,N_8083,N_6420);
nand U11180 (N_11180,N_6870,N_6303);
nand U11181 (N_11181,N_8070,N_7781);
or U11182 (N_11182,N_7967,N_7468);
and U11183 (N_11183,N_7545,N_7160);
nor U11184 (N_11184,N_7783,N_8131);
and U11185 (N_11185,N_7146,N_8689);
nor U11186 (N_11186,N_8696,N_6764);
and U11187 (N_11187,N_6590,N_7468);
nor U11188 (N_11188,N_7463,N_6705);
and U11189 (N_11189,N_7170,N_7026);
xor U11190 (N_11190,N_6222,N_6478);
nand U11191 (N_11191,N_8044,N_6168);
and U11192 (N_11192,N_8962,N_6579);
or U11193 (N_11193,N_7206,N_7415);
or U11194 (N_11194,N_8388,N_8760);
and U11195 (N_11195,N_7498,N_7474);
or U11196 (N_11196,N_7339,N_7696);
nor U11197 (N_11197,N_7244,N_7322);
and U11198 (N_11198,N_6050,N_8978);
and U11199 (N_11199,N_6303,N_7924);
or U11200 (N_11200,N_7235,N_7661);
or U11201 (N_11201,N_6162,N_7884);
and U11202 (N_11202,N_7426,N_8748);
and U11203 (N_11203,N_8387,N_8449);
nand U11204 (N_11204,N_6790,N_7897);
nand U11205 (N_11205,N_8482,N_8180);
nand U11206 (N_11206,N_7374,N_8942);
nand U11207 (N_11207,N_8554,N_8900);
nor U11208 (N_11208,N_7118,N_6365);
nand U11209 (N_11209,N_6119,N_6569);
nor U11210 (N_11210,N_6154,N_7385);
xor U11211 (N_11211,N_7121,N_8014);
xor U11212 (N_11212,N_8683,N_8767);
nor U11213 (N_11213,N_7307,N_7732);
nor U11214 (N_11214,N_6937,N_7405);
nand U11215 (N_11215,N_7495,N_7381);
nand U11216 (N_11216,N_7700,N_7491);
nor U11217 (N_11217,N_8575,N_8816);
and U11218 (N_11218,N_8174,N_7098);
nor U11219 (N_11219,N_6353,N_8765);
nand U11220 (N_11220,N_7133,N_7562);
nor U11221 (N_11221,N_8279,N_7197);
or U11222 (N_11222,N_6485,N_8849);
xnor U11223 (N_11223,N_8246,N_7546);
or U11224 (N_11224,N_7161,N_8958);
nand U11225 (N_11225,N_8035,N_6006);
nor U11226 (N_11226,N_7739,N_7066);
nor U11227 (N_11227,N_8771,N_8846);
nand U11228 (N_11228,N_6061,N_8108);
or U11229 (N_11229,N_6066,N_6740);
nand U11230 (N_11230,N_8427,N_7180);
or U11231 (N_11231,N_6532,N_6713);
and U11232 (N_11232,N_7143,N_7241);
or U11233 (N_11233,N_7758,N_6241);
or U11234 (N_11234,N_8000,N_7990);
or U11235 (N_11235,N_8361,N_8258);
nand U11236 (N_11236,N_6729,N_8153);
or U11237 (N_11237,N_7334,N_8489);
nor U11238 (N_11238,N_6133,N_6667);
or U11239 (N_11239,N_6661,N_6361);
and U11240 (N_11240,N_8883,N_8298);
nand U11241 (N_11241,N_6053,N_7923);
or U11242 (N_11242,N_6247,N_6194);
and U11243 (N_11243,N_8306,N_6914);
xnor U11244 (N_11244,N_7225,N_6349);
or U11245 (N_11245,N_8472,N_8767);
nand U11246 (N_11246,N_6425,N_6442);
or U11247 (N_11247,N_7242,N_7774);
and U11248 (N_11248,N_6189,N_7545);
nor U11249 (N_11249,N_7360,N_8397);
or U11250 (N_11250,N_7967,N_8017);
nor U11251 (N_11251,N_6253,N_8499);
nand U11252 (N_11252,N_8805,N_6003);
or U11253 (N_11253,N_6131,N_8614);
and U11254 (N_11254,N_8693,N_8602);
xnor U11255 (N_11255,N_8827,N_6054);
nand U11256 (N_11256,N_8638,N_8509);
and U11257 (N_11257,N_6813,N_6346);
and U11258 (N_11258,N_6867,N_8505);
nor U11259 (N_11259,N_6753,N_6734);
and U11260 (N_11260,N_7506,N_8296);
and U11261 (N_11261,N_7736,N_8096);
nand U11262 (N_11262,N_6909,N_7877);
or U11263 (N_11263,N_7491,N_8479);
nand U11264 (N_11264,N_8280,N_7015);
nor U11265 (N_11265,N_7089,N_8137);
nor U11266 (N_11266,N_7275,N_7661);
or U11267 (N_11267,N_6007,N_7224);
or U11268 (N_11268,N_6948,N_8775);
nor U11269 (N_11269,N_7082,N_8241);
nor U11270 (N_11270,N_8962,N_8633);
nand U11271 (N_11271,N_8509,N_7173);
or U11272 (N_11272,N_7090,N_7931);
nor U11273 (N_11273,N_7900,N_8479);
nor U11274 (N_11274,N_6874,N_7343);
or U11275 (N_11275,N_6616,N_6450);
or U11276 (N_11276,N_8114,N_6200);
and U11277 (N_11277,N_7668,N_7913);
nand U11278 (N_11278,N_8934,N_8840);
nor U11279 (N_11279,N_8957,N_6142);
or U11280 (N_11280,N_6779,N_7488);
nand U11281 (N_11281,N_8298,N_6863);
xor U11282 (N_11282,N_7274,N_7735);
xor U11283 (N_11283,N_6421,N_6497);
xnor U11284 (N_11284,N_7227,N_6115);
nor U11285 (N_11285,N_6784,N_8449);
nor U11286 (N_11286,N_8748,N_7348);
xor U11287 (N_11287,N_8882,N_7833);
or U11288 (N_11288,N_8193,N_7742);
and U11289 (N_11289,N_6017,N_8708);
or U11290 (N_11290,N_8004,N_7317);
nand U11291 (N_11291,N_8386,N_6215);
nor U11292 (N_11292,N_6646,N_8145);
and U11293 (N_11293,N_8248,N_6301);
nor U11294 (N_11294,N_8732,N_6957);
xnor U11295 (N_11295,N_7987,N_6325);
and U11296 (N_11296,N_6190,N_7917);
or U11297 (N_11297,N_7036,N_6682);
and U11298 (N_11298,N_6026,N_8301);
and U11299 (N_11299,N_7122,N_6198);
nor U11300 (N_11300,N_6944,N_8409);
or U11301 (N_11301,N_7415,N_7662);
nor U11302 (N_11302,N_7947,N_7299);
nand U11303 (N_11303,N_8642,N_6937);
and U11304 (N_11304,N_8264,N_7515);
and U11305 (N_11305,N_7242,N_6822);
nand U11306 (N_11306,N_6386,N_6279);
and U11307 (N_11307,N_8909,N_8746);
and U11308 (N_11308,N_7359,N_6817);
nor U11309 (N_11309,N_6126,N_7328);
nor U11310 (N_11310,N_8439,N_6431);
nand U11311 (N_11311,N_7072,N_6098);
or U11312 (N_11312,N_6618,N_7176);
or U11313 (N_11313,N_8741,N_8402);
nand U11314 (N_11314,N_8034,N_7909);
nand U11315 (N_11315,N_8168,N_6441);
nand U11316 (N_11316,N_6973,N_6253);
nor U11317 (N_11317,N_6546,N_7023);
and U11318 (N_11318,N_8250,N_7680);
nor U11319 (N_11319,N_8229,N_8211);
nor U11320 (N_11320,N_7815,N_7831);
and U11321 (N_11321,N_6662,N_7586);
and U11322 (N_11322,N_7089,N_7938);
and U11323 (N_11323,N_6038,N_6286);
and U11324 (N_11324,N_7268,N_7899);
nor U11325 (N_11325,N_8553,N_6717);
nand U11326 (N_11326,N_8785,N_8378);
and U11327 (N_11327,N_7570,N_8209);
nor U11328 (N_11328,N_8755,N_8222);
or U11329 (N_11329,N_8783,N_7047);
nand U11330 (N_11330,N_6344,N_7167);
nand U11331 (N_11331,N_6077,N_6609);
and U11332 (N_11332,N_8715,N_6312);
or U11333 (N_11333,N_6545,N_7103);
nand U11334 (N_11334,N_8374,N_7744);
or U11335 (N_11335,N_8125,N_8416);
nand U11336 (N_11336,N_7624,N_8829);
xor U11337 (N_11337,N_7915,N_6825);
nor U11338 (N_11338,N_7482,N_8512);
nor U11339 (N_11339,N_8417,N_8759);
nor U11340 (N_11340,N_7896,N_8662);
or U11341 (N_11341,N_7755,N_8894);
nor U11342 (N_11342,N_8556,N_6832);
or U11343 (N_11343,N_8573,N_6571);
nor U11344 (N_11344,N_7867,N_8854);
or U11345 (N_11345,N_6077,N_6628);
nor U11346 (N_11346,N_6419,N_7266);
nor U11347 (N_11347,N_6632,N_8027);
or U11348 (N_11348,N_7881,N_8028);
nand U11349 (N_11349,N_7348,N_7341);
and U11350 (N_11350,N_8828,N_8187);
nor U11351 (N_11351,N_7360,N_6102);
nor U11352 (N_11352,N_7015,N_6035);
and U11353 (N_11353,N_7170,N_7407);
nor U11354 (N_11354,N_8204,N_7334);
xnor U11355 (N_11355,N_6719,N_7238);
nand U11356 (N_11356,N_7470,N_6984);
or U11357 (N_11357,N_6843,N_6983);
and U11358 (N_11358,N_6551,N_6457);
or U11359 (N_11359,N_8011,N_8253);
or U11360 (N_11360,N_8205,N_7093);
nor U11361 (N_11361,N_8008,N_6405);
xnor U11362 (N_11362,N_7367,N_7828);
xnor U11363 (N_11363,N_6826,N_8807);
nand U11364 (N_11364,N_6364,N_7912);
nor U11365 (N_11365,N_6263,N_8999);
nor U11366 (N_11366,N_8096,N_6641);
and U11367 (N_11367,N_8803,N_6579);
nand U11368 (N_11368,N_8520,N_7389);
nand U11369 (N_11369,N_6687,N_7238);
and U11370 (N_11370,N_8480,N_8696);
nor U11371 (N_11371,N_7743,N_7345);
or U11372 (N_11372,N_7447,N_6468);
xnor U11373 (N_11373,N_8029,N_6452);
or U11374 (N_11374,N_8623,N_6606);
xnor U11375 (N_11375,N_6195,N_6852);
nor U11376 (N_11376,N_6835,N_7886);
and U11377 (N_11377,N_8044,N_8472);
xnor U11378 (N_11378,N_8322,N_8913);
nand U11379 (N_11379,N_8034,N_7733);
and U11380 (N_11380,N_8128,N_8280);
or U11381 (N_11381,N_6852,N_8169);
and U11382 (N_11382,N_8743,N_6103);
or U11383 (N_11383,N_6922,N_8050);
nor U11384 (N_11384,N_6384,N_8572);
or U11385 (N_11385,N_7810,N_8114);
nand U11386 (N_11386,N_8598,N_6826);
and U11387 (N_11387,N_7550,N_8923);
nand U11388 (N_11388,N_8030,N_8319);
xnor U11389 (N_11389,N_6990,N_7517);
or U11390 (N_11390,N_8754,N_6078);
xor U11391 (N_11391,N_8840,N_6520);
nand U11392 (N_11392,N_7801,N_6536);
nor U11393 (N_11393,N_8436,N_7378);
xnor U11394 (N_11394,N_7428,N_8128);
xor U11395 (N_11395,N_6782,N_7995);
nand U11396 (N_11396,N_8759,N_6117);
or U11397 (N_11397,N_8018,N_8750);
nand U11398 (N_11398,N_7711,N_7482);
nor U11399 (N_11399,N_8281,N_7168);
nor U11400 (N_11400,N_6526,N_6571);
and U11401 (N_11401,N_8280,N_7061);
and U11402 (N_11402,N_6025,N_6361);
or U11403 (N_11403,N_7403,N_8568);
nand U11404 (N_11404,N_8533,N_7413);
and U11405 (N_11405,N_8755,N_7817);
and U11406 (N_11406,N_7791,N_7667);
nor U11407 (N_11407,N_7883,N_8382);
nand U11408 (N_11408,N_8773,N_6416);
and U11409 (N_11409,N_7345,N_7467);
nor U11410 (N_11410,N_8886,N_8343);
nor U11411 (N_11411,N_6522,N_7535);
xnor U11412 (N_11412,N_6702,N_7136);
nand U11413 (N_11413,N_6870,N_6397);
nand U11414 (N_11414,N_7783,N_6299);
nor U11415 (N_11415,N_6939,N_7070);
and U11416 (N_11416,N_8716,N_7786);
or U11417 (N_11417,N_7733,N_6399);
nor U11418 (N_11418,N_6535,N_8103);
nor U11419 (N_11419,N_8747,N_7523);
or U11420 (N_11420,N_6122,N_7097);
or U11421 (N_11421,N_8165,N_8107);
or U11422 (N_11422,N_8691,N_7840);
nor U11423 (N_11423,N_7858,N_7849);
and U11424 (N_11424,N_8434,N_7728);
xor U11425 (N_11425,N_8558,N_6129);
nand U11426 (N_11426,N_8036,N_6410);
and U11427 (N_11427,N_7946,N_6744);
nand U11428 (N_11428,N_8334,N_7629);
or U11429 (N_11429,N_7688,N_7097);
nand U11430 (N_11430,N_8868,N_6112);
nor U11431 (N_11431,N_6408,N_8356);
or U11432 (N_11432,N_7570,N_7645);
nor U11433 (N_11433,N_6270,N_7767);
or U11434 (N_11434,N_8484,N_6935);
nand U11435 (N_11435,N_8310,N_7336);
nand U11436 (N_11436,N_8381,N_8464);
nand U11437 (N_11437,N_6226,N_6068);
nor U11438 (N_11438,N_6679,N_7549);
and U11439 (N_11439,N_6510,N_7396);
xnor U11440 (N_11440,N_6877,N_7788);
and U11441 (N_11441,N_6710,N_8214);
nor U11442 (N_11442,N_7802,N_8787);
or U11443 (N_11443,N_6981,N_7655);
xor U11444 (N_11444,N_6276,N_6996);
and U11445 (N_11445,N_7349,N_7831);
and U11446 (N_11446,N_8330,N_6786);
or U11447 (N_11447,N_6787,N_6922);
nor U11448 (N_11448,N_7463,N_7782);
nand U11449 (N_11449,N_7545,N_7792);
and U11450 (N_11450,N_7116,N_7592);
xor U11451 (N_11451,N_8687,N_7540);
nand U11452 (N_11452,N_7702,N_8659);
and U11453 (N_11453,N_7159,N_6260);
and U11454 (N_11454,N_6035,N_7564);
nor U11455 (N_11455,N_7514,N_7740);
and U11456 (N_11456,N_7590,N_6485);
nor U11457 (N_11457,N_7228,N_8419);
and U11458 (N_11458,N_7833,N_7201);
and U11459 (N_11459,N_7128,N_8530);
or U11460 (N_11460,N_7313,N_6280);
and U11461 (N_11461,N_8603,N_6295);
nand U11462 (N_11462,N_7898,N_8341);
nor U11463 (N_11463,N_8635,N_7048);
nand U11464 (N_11464,N_7676,N_6881);
nand U11465 (N_11465,N_7220,N_8421);
or U11466 (N_11466,N_7587,N_8337);
xnor U11467 (N_11467,N_7507,N_6020);
nor U11468 (N_11468,N_8030,N_8051);
nand U11469 (N_11469,N_8574,N_6046);
and U11470 (N_11470,N_7183,N_6439);
nand U11471 (N_11471,N_6221,N_8615);
xor U11472 (N_11472,N_7622,N_7023);
and U11473 (N_11473,N_6070,N_8790);
or U11474 (N_11474,N_6457,N_8191);
nor U11475 (N_11475,N_6919,N_7049);
or U11476 (N_11476,N_7044,N_7530);
and U11477 (N_11477,N_8651,N_8434);
nand U11478 (N_11478,N_6853,N_6953);
xor U11479 (N_11479,N_6674,N_7964);
or U11480 (N_11480,N_8555,N_6994);
nor U11481 (N_11481,N_6016,N_7576);
nand U11482 (N_11482,N_6132,N_7589);
nand U11483 (N_11483,N_6065,N_8172);
and U11484 (N_11484,N_7484,N_6722);
xor U11485 (N_11485,N_7199,N_6036);
nor U11486 (N_11486,N_7027,N_6151);
xor U11487 (N_11487,N_7905,N_7748);
nor U11488 (N_11488,N_7921,N_8487);
nor U11489 (N_11489,N_8139,N_8629);
nor U11490 (N_11490,N_6167,N_6881);
nor U11491 (N_11491,N_8275,N_6832);
nand U11492 (N_11492,N_6476,N_6146);
or U11493 (N_11493,N_6883,N_6448);
nand U11494 (N_11494,N_7328,N_6757);
xnor U11495 (N_11495,N_7280,N_6714);
xor U11496 (N_11496,N_8584,N_7404);
and U11497 (N_11497,N_7995,N_8642);
and U11498 (N_11498,N_8963,N_6693);
nor U11499 (N_11499,N_7389,N_6509);
nor U11500 (N_11500,N_8897,N_8529);
nand U11501 (N_11501,N_7321,N_7463);
or U11502 (N_11502,N_6458,N_8335);
or U11503 (N_11503,N_6304,N_6306);
or U11504 (N_11504,N_8856,N_7125);
nor U11505 (N_11505,N_7402,N_6900);
nand U11506 (N_11506,N_7229,N_7674);
xor U11507 (N_11507,N_8845,N_8769);
nor U11508 (N_11508,N_6869,N_7429);
xor U11509 (N_11509,N_8434,N_6998);
or U11510 (N_11510,N_6088,N_6338);
nor U11511 (N_11511,N_7309,N_6563);
nand U11512 (N_11512,N_7151,N_8382);
nand U11513 (N_11513,N_8340,N_7498);
nor U11514 (N_11514,N_7060,N_7109);
nand U11515 (N_11515,N_8871,N_6946);
xnor U11516 (N_11516,N_6402,N_6280);
and U11517 (N_11517,N_6769,N_6443);
and U11518 (N_11518,N_6232,N_6135);
or U11519 (N_11519,N_7127,N_8529);
xnor U11520 (N_11520,N_7260,N_7118);
or U11521 (N_11521,N_8383,N_6973);
nor U11522 (N_11522,N_7438,N_6483);
nand U11523 (N_11523,N_7921,N_6743);
and U11524 (N_11524,N_6789,N_8186);
nor U11525 (N_11525,N_6152,N_8856);
xnor U11526 (N_11526,N_7737,N_7778);
or U11527 (N_11527,N_7262,N_8173);
nand U11528 (N_11528,N_8809,N_7444);
nand U11529 (N_11529,N_7034,N_7850);
xor U11530 (N_11530,N_8821,N_7544);
nand U11531 (N_11531,N_7239,N_6710);
or U11532 (N_11532,N_8430,N_8653);
xor U11533 (N_11533,N_7426,N_7907);
or U11534 (N_11534,N_6588,N_6956);
xor U11535 (N_11535,N_8857,N_8314);
nand U11536 (N_11536,N_8262,N_6131);
and U11537 (N_11537,N_6554,N_7768);
nand U11538 (N_11538,N_7360,N_8463);
and U11539 (N_11539,N_8146,N_6275);
and U11540 (N_11540,N_6107,N_8661);
and U11541 (N_11541,N_6824,N_7584);
nand U11542 (N_11542,N_7749,N_8439);
nor U11543 (N_11543,N_8309,N_6851);
or U11544 (N_11544,N_8678,N_7566);
or U11545 (N_11545,N_6203,N_6642);
or U11546 (N_11546,N_7464,N_8706);
or U11547 (N_11547,N_7420,N_7557);
or U11548 (N_11548,N_8277,N_7289);
nand U11549 (N_11549,N_7903,N_8461);
and U11550 (N_11550,N_8938,N_7802);
or U11551 (N_11551,N_8713,N_7172);
nor U11552 (N_11552,N_6273,N_8963);
or U11553 (N_11553,N_8690,N_6728);
and U11554 (N_11554,N_6460,N_6558);
nor U11555 (N_11555,N_7519,N_6708);
or U11556 (N_11556,N_8628,N_6003);
nor U11557 (N_11557,N_6416,N_8294);
nand U11558 (N_11558,N_7229,N_7657);
and U11559 (N_11559,N_7324,N_6827);
nand U11560 (N_11560,N_8983,N_7368);
and U11561 (N_11561,N_8722,N_8901);
nand U11562 (N_11562,N_8313,N_8553);
nor U11563 (N_11563,N_8986,N_7454);
nand U11564 (N_11564,N_6970,N_8558);
nand U11565 (N_11565,N_8703,N_6561);
and U11566 (N_11566,N_7881,N_7153);
nand U11567 (N_11567,N_6575,N_7112);
nand U11568 (N_11568,N_6133,N_8434);
and U11569 (N_11569,N_7115,N_8541);
or U11570 (N_11570,N_7708,N_7583);
nor U11571 (N_11571,N_8881,N_6389);
or U11572 (N_11572,N_6168,N_6105);
and U11573 (N_11573,N_7129,N_6061);
nor U11574 (N_11574,N_8889,N_7506);
and U11575 (N_11575,N_6300,N_8688);
nand U11576 (N_11576,N_8862,N_8133);
nor U11577 (N_11577,N_6183,N_8056);
nor U11578 (N_11578,N_8723,N_7192);
nor U11579 (N_11579,N_8679,N_7085);
nand U11580 (N_11580,N_8183,N_7977);
nor U11581 (N_11581,N_7594,N_7879);
and U11582 (N_11582,N_8814,N_7631);
nand U11583 (N_11583,N_7685,N_7762);
or U11584 (N_11584,N_7469,N_6904);
or U11585 (N_11585,N_7319,N_7379);
nor U11586 (N_11586,N_6304,N_7542);
nor U11587 (N_11587,N_8124,N_6587);
or U11588 (N_11588,N_8327,N_8479);
or U11589 (N_11589,N_7053,N_6354);
nor U11590 (N_11590,N_7043,N_8646);
or U11591 (N_11591,N_7842,N_7706);
xnor U11592 (N_11592,N_7397,N_7875);
or U11593 (N_11593,N_8022,N_6554);
nand U11594 (N_11594,N_7442,N_8698);
or U11595 (N_11595,N_8498,N_6627);
or U11596 (N_11596,N_8781,N_6507);
and U11597 (N_11597,N_6055,N_8278);
nor U11598 (N_11598,N_6846,N_8664);
xnor U11599 (N_11599,N_7337,N_6984);
xnor U11600 (N_11600,N_6433,N_6366);
and U11601 (N_11601,N_8080,N_7633);
or U11602 (N_11602,N_8226,N_7603);
nor U11603 (N_11603,N_6031,N_7073);
or U11604 (N_11604,N_6433,N_8641);
nand U11605 (N_11605,N_8994,N_8762);
and U11606 (N_11606,N_7100,N_7717);
or U11607 (N_11607,N_7514,N_8774);
and U11608 (N_11608,N_8613,N_6803);
or U11609 (N_11609,N_6888,N_7937);
xor U11610 (N_11610,N_7867,N_6043);
or U11611 (N_11611,N_7969,N_7582);
or U11612 (N_11612,N_6312,N_8784);
nand U11613 (N_11613,N_8822,N_7597);
nor U11614 (N_11614,N_7924,N_8231);
nand U11615 (N_11615,N_6503,N_8490);
or U11616 (N_11616,N_6210,N_7014);
nand U11617 (N_11617,N_8640,N_6242);
and U11618 (N_11618,N_7801,N_7346);
nor U11619 (N_11619,N_6948,N_7805);
or U11620 (N_11620,N_7912,N_7401);
or U11621 (N_11621,N_6227,N_8361);
or U11622 (N_11622,N_6675,N_7167);
or U11623 (N_11623,N_7264,N_8132);
and U11624 (N_11624,N_6685,N_6709);
nor U11625 (N_11625,N_6087,N_6867);
nor U11626 (N_11626,N_8915,N_7642);
or U11627 (N_11627,N_8759,N_6611);
or U11628 (N_11628,N_7244,N_7441);
nand U11629 (N_11629,N_7688,N_8029);
nand U11630 (N_11630,N_8749,N_6384);
nand U11631 (N_11631,N_6065,N_6476);
nor U11632 (N_11632,N_7518,N_8468);
nor U11633 (N_11633,N_7785,N_8620);
nor U11634 (N_11634,N_8833,N_6680);
nor U11635 (N_11635,N_6434,N_8146);
nor U11636 (N_11636,N_8800,N_7819);
nand U11637 (N_11637,N_6926,N_8922);
nor U11638 (N_11638,N_6537,N_8293);
nand U11639 (N_11639,N_7568,N_8087);
and U11640 (N_11640,N_7177,N_8611);
xor U11641 (N_11641,N_8539,N_6492);
xnor U11642 (N_11642,N_7687,N_6584);
nand U11643 (N_11643,N_8534,N_6267);
nand U11644 (N_11644,N_8904,N_6887);
nor U11645 (N_11645,N_6408,N_8916);
nor U11646 (N_11646,N_8667,N_8595);
nand U11647 (N_11647,N_7292,N_6715);
or U11648 (N_11648,N_7790,N_8974);
xor U11649 (N_11649,N_8935,N_6921);
or U11650 (N_11650,N_6723,N_8262);
nor U11651 (N_11651,N_6389,N_6613);
or U11652 (N_11652,N_6430,N_7690);
xnor U11653 (N_11653,N_8096,N_7982);
xnor U11654 (N_11654,N_6109,N_8094);
nor U11655 (N_11655,N_6364,N_7150);
xnor U11656 (N_11656,N_6495,N_6333);
nor U11657 (N_11657,N_7756,N_7374);
or U11658 (N_11658,N_8281,N_6780);
and U11659 (N_11659,N_6315,N_7424);
nor U11660 (N_11660,N_7752,N_6111);
nand U11661 (N_11661,N_6124,N_8347);
and U11662 (N_11662,N_7114,N_8182);
nand U11663 (N_11663,N_7339,N_7632);
or U11664 (N_11664,N_8181,N_8089);
nand U11665 (N_11665,N_6114,N_7783);
or U11666 (N_11666,N_8615,N_8962);
and U11667 (N_11667,N_7804,N_8887);
and U11668 (N_11668,N_7371,N_6532);
and U11669 (N_11669,N_6732,N_8085);
and U11670 (N_11670,N_7730,N_7191);
and U11671 (N_11671,N_6339,N_6572);
or U11672 (N_11672,N_7782,N_8707);
nand U11673 (N_11673,N_6488,N_8168);
nand U11674 (N_11674,N_8656,N_7254);
xnor U11675 (N_11675,N_6365,N_6676);
nor U11676 (N_11676,N_6166,N_6261);
nand U11677 (N_11677,N_8652,N_6913);
nor U11678 (N_11678,N_7204,N_6270);
nor U11679 (N_11679,N_8688,N_8245);
xnor U11680 (N_11680,N_6045,N_8599);
and U11681 (N_11681,N_6393,N_6300);
nor U11682 (N_11682,N_6334,N_8192);
nand U11683 (N_11683,N_6080,N_6290);
nor U11684 (N_11684,N_8912,N_8759);
nor U11685 (N_11685,N_8594,N_6911);
xnor U11686 (N_11686,N_8226,N_7419);
and U11687 (N_11687,N_8276,N_8507);
xnor U11688 (N_11688,N_8497,N_7531);
nand U11689 (N_11689,N_7676,N_6020);
or U11690 (N_11690,N_7906,N_8735);
nand U11691 (N_11691,N_7233,N_8015);
nor U11692 (N_11692,N_6148,N_6037);
or U11693 (N_11693,N_6371,N_7293);
and U11694 (N_11694,N_8451,N_6947);
nand U11695 (N_11695,N_7826,N_8409);
and U11696 (N_11696,N_7623,N_8649);
or U11697 (N_11697,N_6567,N_7406);
and U11698 (N_11698,N_6552,N_8394);
or U11699 (N_11699,N_8048,N_8472);
and U11700 (N_11700,N_8081,N_8920);
nor U11701 (N_11701,N_6758,N_7224);
or U11702 (N_11702,N_8933,N_8099);
nor U11703 (N_11703,N_6191,N_8932);
or U11704 (N_11704,N_8933,N_7736);
and U11705 (N_11705,N_8453,N_6258);
or U11706 (N_11706,N_8175,N_7758);
nand U11707 (N_11707,N_7327,N_7893);
nand U11708 (N_11708,N_6780,N_6239);
nor U11709 (N_11709,N_6412,N_6696);
and U11710 (N_11710,N_8174,N_6043);
xnor U11711 (N_11711,N_7440,N_7428);
or U11712 (N_11712,N_7195,N_8337);
or U11713 (N_11713,N_8171,N_6752);
xor U11714 (N_11714,N_8530,N_8962);
nor U11715 (N_11715,N_6262,N_7090);
nor U11716 (N_11716,N_6184,N_6052);
nand U11717 (N_11717,N_7764,N_8324);
and U11718 (N_11718,N_7959,N_6495);
xnor U11719 (N_11719,N_7352,N_8951);
and U11720 (N_11720,N_8349,N_7566);
xnor U11721 (N_11721,N_6236,N_6719);
nor U11722 (N_11722,N_6089,N_8926);
nand U11723 (N_11723,N_8830,N_8865);
nor U11724 (N_11724,N_6956,N_8703);
nor U11725 (N_11725,N_8022,N_7670);
or U11726 (N_11726,N_8951,N_7106);
nand U11727 (N_11727,N_8050,N_7477);
or U11728 (N_11728,N_7621,N_7706);
or U11729 (N_11729,N_7229,N_7447);
nor U11730 (N_11730,N_8122,N_8676);
nor U11731 (N_11731,N_6776,N_8747);
nor U11732 (N_11732,N_7080,N_8021);
and U11733 (N_11733,N_7409,N_7887);
or U11734 (N_11734,N_8229,N_8153);
nor U11735 (N_11735,N_6005,N_6410);
nand U11736 (N_11736,N_6773,N_6508);
nand U11737 (N_11737,N_7475,N_7801);
and U11738 (N_11738,N_8586,N_8708);
or U11739 (N_11739,N_8005,N_6643);
or U11740 (N_11740,N_8696,N_7004);
nand U11741 (N_11741,N_8418,N_8685);
and U11742 (N_11742,N_6959,N_7653);
nor U11743 (N_11743,N_6316,N_6083);
and U11744 (N_11744,N_7159,N_6891);
nand U11745 (N_11745,N_6865,N_6719);
nand U11746 (N_11746,N_6994,N_7677);
nand U11747 (N_11747,N_8936,N_7622);
and U11748 (N_11748,N_7490,N_6523);
and U11749 (N_11749,N_8448,N_8540);
and U11750 (N_11750,N_7975,N_7222);
and U11751 (N_11751,N_7903,N_7369);
nand U11752 (N_11752,N_7493,N_8106);
nand U11753 (N_11753,N_6162,N_6293);
nand U11754 (N_11754,N_6013,N_6113);
or U11755 (N_11755,N_6714,N_6347);
or U11756 (N_11756,N_7094,N_8923);
or U11757 (N_11757,N_8036,N_7350);
nand U11758 (N_11758,N_8655,N_7481);
and U11759 (N_11759,N_7866,N_7069);
nor U11760 (N_11760,N_7427,N_8866);
nor U11761 (N_11761,N_6119,N_8142);
and U11762 (N_11762,N_6122,N_8248);
or U11763 (N_11763,N_7174,N_8687);
and U11764 (N_11764,N_6020,N_7706);
nor U11765 (N_11765,N_6349,N_8745);
nor U11766 (N_11766,N_8060,N_8788);
and U11767 (N_11767,N_6459,N_6280);
nand U11768 (N_11768,N_7510,N_8728);
or U11769 (N_11769,N_6578,N_6269);
nand U11770 (N_11770,N_6130,N_7803);
xnor U11771 (N_11771,N_8018,N_7785);
or U11772 (N_11772,N_7394,N_6389);
nand U11773 (N_11773,N_7014,N_8024);
or U11774 (N_11774,N_7746,N_7823);
or U11775 (N_11775,N_6352,N_6657);
xnor U11776 (N_11776,N_7781,N_8460);
nor U11777 (N_11777,N_7574,N_8102);
nand U11778 (N_11778,N_7729,N_8665);
nor U11779 (N_11779,N_8043,N_6847);
nand U11780 (N_11780,N_8232,N_8970);
nand U11781 (N_11781,N_7496,N_8037);
and U11782 (N_11782,N_7008,N_8014);
and U11783 (N_11783,N_6795,N_7598);
and U11784 (N_11784,N_6062,N_7953);
and U11785 (N_11785,N_6938,N_6168);
and U11786 (N_11786,N_8769,N_7757);
or U11787 (N_11787,N_6992,N_6516);
nand U11788 (N_11788,N_7964,N_7681);
xnor U11789 (N_11789,N_6387,N_7509);
or U11790 (N_11790,N_6769,N_7129);
nor U11791 (N_11791,N_8203,N_8118);
and U11792 (N_11792,N_6990,N_6321);
nor U11793 (N_11793,N_6211,N_7999);
and U11794 (N_11794,N_7058,N_6172);
nand U11795 (N_11795,N_6299,N_8161);
xnor U11796 (N_11796,N_8367,N_6503);
nor U11797 (N_11797,N_6915,N_6905);
and U11798 (N_11798,N_8121,N_7128);
nand U11799 (N_11799,N_8359,N_8068);
and U11800 (N_11800,N_7961,N_8792);
or U11801 (N_11801,N_8113,N_8593);
or U11802 (N_11802,N_8866,N_7480);
nor U11803 (N_11803,N_7839,N_8406);
or U11804 (N_11804,N_7041,N_7027);
nand U11805 (N_11805,N_7953,N_8387);
or U11806 (N_11806,N_7347,N_7883);
and U11807 (N_11807,N_7845,N_8399);
and U11808 (N_11808,N_6966,N_6364);
and U11809 (N_11809,N_7832,N_7631);
and U11810 (N_11810,N_8751,N_7322);
nor U11811 (N_11811,N_7613,N_8018);
and U11812 (N_11812,N_7332,N_6516);
and U11813 (N_11813,N_7943,N_6955);
xor U11814 (N_11814,N_6458,N_7827);
xor U11815 (N_11815,N_7231,N_6239);
and U11816 (N_11816,N_7017,N_6534);
nand U11817 (N_11817,N_6082,N_6479);
nand U11818 (N_11818,N_6894,N_6850);
nand U11819 (N_11819,N_6349,N_7763);
nand U11820 (N_11820,N_7325,N_8025);
or U11821 (N_11821,N_7458,N_6703);
nor U11822 (N_11822,N_8710,N_7503);
nor U11823 (N_11823,N_8643,N_6764);
or U11824 (N_11824,N_6001,N_7734);
nor U11825 (N_11825,N_6414,N_6770);
or U11826 (N_11826,N_7226,N_6460);
nor U11827 (N_11827,N_8557,N_7601);
and U11828 (N_11828,N_6321,N_8698);
and U11829 (N_11829,N_6668,N_8180);
nand U11830 (N_11830,N_8401,N_8566);
nand U11831 (N_11831,N_7714,N_6965);
or U11832 (N_11832,N_6315,N_6487);
or U11833 (N_11833,N_7882,N_6181);
nand U11834 (N_11834,N_8812,N_7550);
or U11835 (N_11835,N_7738,N_7441);
nand U11836 (N_11836,N_8461,N_7228);
nor U11837 (N_11837,N_6803,N_6810);
nor U11838 (N_11838,N_8615,N_8649);
nand U11839 (N_11839,N_6527,N_6350);
and U11840 (N_11840,N_7291,N_7144);
nand U11841 (N_11841,N_6665,N_7430);
or U11842 (N_11842,N_6798,N_6414);
or U11843 (N_11843,N_6273,N_6262);
nor U11844 (N_11844,N_6034,N_8879);
nand U11845 (N_11845,N_8131,N_6608);
nand U11846 (N_11846,N_6762,N_8307);
or U11847 (N_11847,N_6486,N_6485);
or U11848 (N_11848,N_6251,N_6736);
or U11849 (N_11849,N_7990,N_8067);
or U11850 (N_11850,N_7832,N_8439);
or U11851 (N_11851,N_7499,N_8665);
xor U11852 (N_11852,N_7245,N_6545);
xnor U11853 (N_11853,N_6752,N_8689);
nor U11854 (N_11854,N_8838,N_7841);
and U11855 (N_11855,N_8363,N_7558);
and U11856 (N_11856,N_7698,N_8432);
nor U11857 (N_11857,N_6767,N_6175);
nor U11858 (N_11858,N_8936,N_7571);
or U11859 (N_11859,N_6863,N_6303);
nor U11860 (N_11860,N_6955,N_6921);
nor U11861 (N_11861,N_7427,N_6141);
nand U11862 (N_11862,N_7930,N_8272);
xor U11863 (N_11863,N_7987,N_7407);
nand U11864 (N_11864,N_6619,N_6412);
nand U11865 (N_11865,N_8412,N_6534);
nor U11866 (N_11866,N_6547,N_8571);
and U11867 (N_11867,N_6346,N_6980);
nor U11868 (N_11868,N_6554,N_8026);
or U11869 (N_11869,N_6071,N_8042);
nand U11870 (N_11870,N_6814,N_8313);
and U11871 (N_11871,N_8627,N_6253);
nor U11872 (N_11872,N_8849,N_6599);
nor U11873 (N_11873,N_6879,N_7208);
nand U11874 (N_11874,N_8140,N_8044);
nand U11875 (N_11875,N_7485,N_6036);
nand U11876 (N_11876,N_7530,N_6658);
or U11877 (N_11877,N_8728,N_8338);
xor U11878 (N_11878,N_7261,N_7957);
nand U11879 (N_11879,N_8811,N_6622);
or U11880 (N_11880,N_6471,N_8024);
or U11881 (N_11881,N_7358,N_7548);
or U11882 (N_11882,N_6947,N_6657);
or U11883 (N_11883,N_6696,N_7446);
nand U11884 (N_11884,N_6082,N_6930);
and U11885 (N_11885,N_7231,N_6598);
nand U11886 (N_11886,N_8718,N_8881);
nor U11887 (N_11887,N_7024,N_6677);
or U11888 (N_11888,N_8890,N_8532);
and U11889 (N_11889,N_8777,N_6547);
nand U11890 (N_11890,N_8694,N_8719);
nor U11891 (N_11891,N_8534,N_8465);
nor U11892 (N_11892,N_6360,N_8806);
nor U11893 (N_11893,N_6190,N_7483);
nand U11894 (N_11894,N_7431,N_7965);
nand U11895 (N_11895,N_6500,N_8750);
nand U11896 (N_11896,N_8459,N_6371);
or U11897 (N_11897,N_6001,N_6641);
and U11898 (N_11898,N_6769,N_6080);
and U11899 (N_11899,N_8572,N_6348);
and U11900 (N_11900,N_6672,N_8139);
nor U11901 (N_11901,N_8180,N_7275);
or U11902 (N_11902,N_7010,N_7380);
nor U11903 (N_11903,N_7282,N_6202);
nor U11904 (N_11904,N_7752,N_6179);
nand U11905 (N_11905,N_6771,N_8274);
xor U11906 (N_11906,N_6280,N_8195);
and U11907 (N_11907,N_6668,N_8009);
or U11908 (N_11908,N_6037,N_6705);
nand U11909 (N_11909,N_8132,N_7097);
nor U11910 (N_11910,N_6758,N_6125);
nor U11911 (N_11911,N_6361,N_8013);
nor U11912 (N_11912,N_7154,N_8012);
nand U11913 (N_11913,N_8787,N_7429);
nand U11914 (N_11914,N_6538,N_8655);
and U11915 (N_11915,N_7674,N_7990);
or U11916 (N_11916,N_6870,N_6393);
xor U11917 (N_11917,N_7719,N_8791);
nand U11918 (N_11918,N_7843,N_8748);
and U11919 (N_11919,N_6186,N_7725);
xor U11920 (N_11920,N_8881,N_8785);
and U11921 (N_11921,N_7339,N_7570);
or U11922 (N_11922,N_8794,N_7461);
and U11923 (N_11923,N_8577,N_6290);
nor U11924 (N_11924,N_7449,N_6551);
nor U11925 (N_11925,N_7916,N_6917);
nor U11926 (N_11926,N_8570,N_7676);
and U11927 (N_11927,N_7155,N_6512);
nand U11928 (N_11928,N_6134,N_8873);
and U11929 (N_11929,N_7887,N_8754);
nor U11930 (N_11930,N_8250,N_7641);
and U11931 (N_11931,N_6475,N_6299);
or U11932 (N_11932,N_8263,N_7208);
nand U11933 (N_11933,N_6610,N_6559);
nor U11934 (N_11934,N_7056,N_8672);
and U11935 (N_11935,N_6657,N_8691);
nor U11936 (N_11936,N_8712,N_6817);
nand U11937 (N_11937,N_7521,N_6190);
xnor U11938 (N_11938,N_6016,N_8196);
nand U11939 (N_11939,N_6186,N_8381);
nor U11940 (N_11940,N_8122,N_7487);
or U11941 (N_11941,N_7450,N_7922);
or U11942 (N_11942,N_8844,N_8256);
and U11943 (N_11943,N_6260,N_8378);
nor U11944 (N_11944,N_6861,N_6422);
or U11945 (N_11945,N_7126,N_6702);
nand U11946 (N_11946,N_8969,N_6800);
and U11947 (N_11947,N_8549,N_7453);
nor U11948 (N_11948,N_8782,N_6772);
nand U11949 (N_11949,N_7441,N_6670);
or U11950 (N_11950,N_8441,N_6702);
nand U11951 (N_11951,N_8914,N_6853);
nor U11952 (N_11952,N_8828,N_6044);
and U11953 (N_11953,N_8288,N_7449);
nand U11954 (N_11954,N_8964,N_7267);
nand U11955 (N_11955,N_6172,N_7972);
and U11956 (N_11956,N_8789,N_7495);
and U11957 (N_11957,N_6052,N_7112);
nand U11958 (N_11958,N_8566,N_7616);
or U11959 (N_11959,N_7311,N_8374);
and U11960 (N_11960,N_6725,N_8613);
nand U11961 (N_11961,N_8497,N_7091);
or U11962 (N_11962,N_7612,N_8488);
and U11963 (N_11963,N_7630,N_6272);
nor U11964 (N_11964,N_7673,N_8720);
and U11965 (N_11965,N_6928,N_6392);
or U11966 (N_11966,N_7822,N_7480);
nor U11967 (N_11967,N_6460,N_6592);
or U11968 (N_11968,N_7729,N_8342);
nand U11969 (N_11969,N_7235,N_8983);
nand U11970 (N_11970,N_8457,N_8706);
or U11971 (N_11971,N_8250,N_8763);
and U11972 (N_11972,N_8624,N_8465);
xor U11973 (N_11973,N_6414,N_6228);
or U11974 (N_11974,N_6233,N_7449);
and U11975 (N_11975,N_8230,N_7356);
xor U11976 (N_11976,N_7479,N_8093);
and U11977 (N_11977,N_8680,N_6671);
and U11978 (N_11978,N_7476,N_7917);
nor U11979 (N_11979,N_8758,N_7365);
nor U11980 (N_11980,N_8248,N_8243);
nand U11981 (N_11981,N_7741,N_6124);
xor U11982 (N_11982,N_7519,N_6032);
or U11983 (N_11983,N_6843,N_8372);
xnor U11984 (N_11984,N_8579,N_7868);
nor U11985 (N_11985,N_7843,N_8029);
nand U11986 (N_11986,N_6468,N_8332);
xor U11987 (N_11987,N_8855,N_7876);
nor U11988 (N_11988,N_8614,N_7844);
nor U11989 (N_11989,N_6146,N_6239);
and U11990 (N_11990,N_6162,N_8330);
and U11991 (N_11991,N_8441,N_8100);
and U11992 (N_11992,N_7672,N_8548);
or U11993 (N_11993,N_7609,N_8945);
xor U11994 (N_11994,N_8669,N_7982);
and U11995 (N_11995,N_7652,N_7039);
nor U11996 (N_11996,N_7642,N_8030);
nand U11997 (N_11997,N_8608,N_6476);
and U11998 (N_11998,N_6217,N_7054);
or U11999 (N_11999,N_7778,N_7081);
and U12000 (N_12000,N_10883,N_11755);
and U12001 (N_12001,N_11684,N_11121);
nand U12002 (N_12002,N_11826,N_11911);
nand U12003 (N_12003,N_10351,N_10029);
or U12004 (N_12004,N_11073,N_11961);
and U12005 (N_12005,N_11460,N_11405);
or U12006 (N_12006,N_11645,N_10049);
nor U12007 (N_12007,N_10120,N_10422);
nand U12008 (N_12008,N_9930,N_11686);
and U12009 (N_12009,N_10701,N_10340);
xor U12010 (N_12010,N_10128,N_10099);
and U12011 (N_12011,N_10987,N_11011);
or U12012 (N_12012,N_10240,N_11087);
and U12013 (N_12013,N_9540,N_10123);
and U12014 (N_12014,N_9010,N_10745);
or U12015 (N_12015,N_10783,N_9165);
nor U12016 (N_12016,N_11822,N_9907);
nor U12017 (N_12017,N_11900,N_11439);
and U12018 (N_12018,N_9917,N_9266);
and U12019 (N_12019,N_9824,N_9614);
nand U12020 (N_12020,N_11481,N_10589);
or U12021 (N_12021,N_10473,N_11504);
and U12022 (N_12022,N_10568,N_11007);
nand U12023 (N_12023,N_11597,N_11063);
nor U12024 (N_12024,N_9332,N_11507);
and U12025 (N_12025,N_9474,N_10521);
nand U12026 (N_12026,N_11476,N_9626);
nand U12027 (N_12027,N_11190,N_10846);
and U12028 (N_12028,N_10124,N_11308);
and U12029 (N_12029,N_10555,N_9643);
nand U12030 (N_12030,N_9077,N_11834);
nand U12031 (N_12031,N_10694,N_10813);
and U12032 (N_12032,N_9151,N_9591);
or U12033 (N_12033,N_10287,N_10384);
nor U12034 (N_12034,N_10429,N_9167);
xnor U12035 (N_12035,N_10769,N_10188);
nor U12036 (N_12036,N_9523,N_9790);
or U12037 (N_12037,N_11110,N_10986);
xnor U12038 (N_12038,N_10379,N_9796);
and U12039 (N_12039,N_9513,N_10418);
nand U12040 (N_12040,N_10547,N_11039);
nor U12041 (N_12041,N_9473,N_11655);
nor U12042 (N_12042,N_9364,N_9316);
nand U12043 (N_12043,N_10233,N_11934);
or U12044 (N_12044,N_10506,N_10200);
and U12045 (N_12045,N_11554,N_11796);
nand U12046 (N_12046,N_11137,N_11168);
and U12047 (N_12047,N_10198,N_11775);
or U12048 (N_12048,N_9327,N_11029);
xor U12049 (N_12049,N_10945,N_10245);
or U12050 (N_12050,N_9793,N_11606);
xnor U12051 (N_12051,N_11015,N_10228);
and U12052 (N_12052,N_9281,N_10087);
xor U12053 (N_12053,N_10677,N_11562);
nand U12054 (N_12054,N_10576,N_9926);
and U12055 (N_12055,N_10356,N_10281);
nand U12056 (N_12056,N_11511,N_9498);
nor U12057 (N_12057,N_11123,N_9982);
and U12058 (N_12058,N_9497,N_11640);
and U12059 (N_12059,N_10999,N_11624);
nand U12060 (N_12060,N_11618,N_11867);
or U12061 (N_12061,N_9622,N_9426);
or U12062 (N_12062,N_9679,N_11901);
or U12063 (N_12063,N_9652,N_11771);
and U12064 (N_12064,N_9999,N_9115);
nand U12065 (N_12065,N_11727,N_11289);
nand U12066 (N_12066,N_10655,N_9318);
and U12067 (N_12067,N_10827,N_11097);
nand U12068 (N_12068,N_11549,N_10432);
nor U12069 (N_12069,N_11045,N_9604);
or U12070 (N_12070,N_10149,N_11575);
or U12071 (N_12071,N_9965,N_11442);
or U12072 (N_12072,N_9903,N_10131);
and U12073 (N_12073,N_9104,N_10220);
nor U12074 (N_12074,N_10014,N_11300);
and U12075 (N_12075,N_9946,N_10598);
nor U12076 (N_12076,N_11064,N_10681);
and U12077 (N_12077,N_11543,N_10165);
and U12078 (N_12078,N_11099,N_10736);
nand U12079 (N_12079,N_9333,N_9755);
nand U12080 (N_12080,N_11279,N_10262);
or U12081 (N_12081,N_9438,N_11178);
nand U12082 (N_12082,N_9057,N_9600);
or U12083 (N_12083,N_10786,N_9273);
or U12084 (N_12084,N_9725,N_9961);
or U12085 (N_12085,N_9393,N_10800);
or U12086 (N_12086,N_11926,N_11927);
or U12087 (N_12087,N_11733,N_10285);
nand U12088 (N_12088,N_11242,N_11421);
nor U12089 (N_12089,N_9861,N_11695);
nor U12090 (N_12090,N_11333,N_10053);
or U12091 (N_12091,N_11579,N_10454);
and U12092 (N_12092,N_9722,N_10507);
or U12093 (N_12093,N_11102,N_10357);
or U12094 (N_12094,N_11610,N_11372);
nand U12095 (N_12095,N_9306,N_10760);
nand U12096 (N_12096,N_10499,N_11519);
or U12097 (N_12097,N_9532,N_11335);
xor U12098 (N_12098,N_10450,N_11057);
nand U12099 (N_12099,N_10135,N_9298);
nand U12100 (N_12100,N_9014,N_9776);
xor U12101 (N_12101,N_10796,N_10737);
nor U12102 (N_12102,N_10092,N_11125);
or U12103 (N_12103,N_11985,N_9519);
nand U12104 (N_12104,N_11856,N_9241);
and U12105 (N_12105,N_9712,N_9385);
xnor U12106 (N_12106,N_10602,N_10145);
or U12107 (N_12107,N_9501,N_10024);
nor U12108 (N_12108,N_10723,N_11096);
nor U12109 (N_12109,N_9789,N_9065);
nor U12110 (N_12110,N_11227,N_10545);
nand U12111 (N_12111,N_10019,N_11506);
and U12112 (N_12112,N_11729,N_11841);
nand U12113 (N_12113,N_9681,N_11066);
xor U12114 (N_12114,N_11968,N_10525);
and U12115 (N_12115,N_9267,N_10662);
nand U12116 (N_12116,N_9952,N_9527);
and U12117 (N_12117,N_9345,N_10907);
nand U12118 (N_12118,N_9927,N_10704);
nor U12119 (N_12119,N_11812,N_10777);
nand U12120 (N_12120,N_11584,N_9211);
and U12121 (N_12121,N_10970,N_9733);
nand U12122 (N_12122,N_11923,N_10807);
xnor U12123 (N_12123,N_10811,N_10041);
or U12124 (N_12124,N_11909,N_10735);
nor U12125 (N_12125,N_10407,N_11591);
nor U12126 (N_12126,N_9746,N_11441);
and U12127 (N_12127,N_11028,N_10540);
and U12128 (N_12128,N_11262,N_10898);
nor U12129 (N_12129,N_9766,N_10981);
nor U12130 (N_12130,N_11523,N_11356);
nand U12131 (N_12131,N_10226,N_9270);
nor U12132 (N_12132,N_9701,N_10924);
nand U12133 (N_12133,N_11540,N_11484);
nor U12134 (N_12134,N_11570,N_11206);
nand U12135 (N_12135,N_10752,N_9798);
or U12136 (N_12136,N_10366,N_9499);
nor U12137 (N_12137,N_11255,N_9970);
and U12138 (N_12138,N_9670,N_9291);
xor U12139 (N_12139,N_11463,N_11149);
nand U12140 (N_12140,N_10746,N_9063);
nor U12141 (N_12141,N_9598,N_9030);
nand U12142 (N_12142,N_10516,N_9463);
nand U12143 (N_12143,N_9718,N_9434);
nor U12144 (N_12144,N_11889,N_10114);
xor U12145 (N_12145,N_9822,N_11032);
nor U12146 (N_12146,N_11843,N_9160);
xor U12147 (N_12147,N_10191,N_10212);
or U12148 (N_12148,N_11040,N_10111);
or U12149 (N_12149,N_10428,N_9511);
and U12150 (N_12150,N_9539,N_10292);
nand U12151 (N_12151,N_11881,N_11823);
and U12152 (N_12152,N_11427,N_11990);
or U12153 (N_12153,N_11217,N_9794);
nor U12154 (N_12154,N_10596,N_10085);
or U12155 (N_12155,N_10480,N_11311);
xnor U12156 (N_12156,N_9979,N_11737);
or U12157 (N_12157,N_10619,N_9860);
nor U12158 (N_12158,N_11397,N_9613);
and U12159 (N_12159,N_10038,N_10529);
and U12160 (N_12160,N_9747,N_9258);
and U12161 (N_12161,N_10204,N_10588);
nor U12162 (N_12162,N_9753,N_10642);
and U12163 (N_12163,N_9447,N_10819);
and U12164 (N_12164,N_10566,N_10495);
and U12165 (N_12165,N_10624,N_11667);
nor U12166 (N_12166,N_10199,N_11450);
nand U12167 (N_12167,N_9736,N_9308);
nand U12168 (N_12168,N_11574,N_11225);
nor U12169 (N_12169,N_9618,N_10782);
or U12170 (N_12170,N_10923,N_11530);
nor U12171 (N_12171,N_9654,N_9015);
and U12172 (N_12172,N_11013,N_10040);
nand U12173 (N_12173,N_9997,N_9198);
nor U12174 (N_12174,N_9097,N_9778);
and U12175 (N_12175,N_11485,N_11907);
nor U12176 (N_12176,N_9581,N_11842);
nor U12177 (N_12177,N_9131,N_9453);
nand U12178 (N_12178,N_10347,N_9492);
or U12179 (N_12179,N_10140,N_11404);
and U12180 (N_12180,N_9639,N_10951);
xnor U12181 (N_12181,N_9302,N_9212);
xor U12182 (N_12182,N_10098,N_11400);
nand U12183 (N_12183,N_10712,N_9853);
or U12184 (N_12184,N_10150,N_11191);
or U12185 (N_12185,N_11364,N_9577);
or U12186 (N_12186,N_11832,N_9471);
xnor U12187 (N_12187,N_10293,N_9686);
nor U12188 (N_12188,N_10443,N_10471);
nor U12189 (N_12189,N_9374,N_10097);
nand U12190 (N_12190,N_9470,N_10685);
or U12191 (N_12191,N_11384,N_9089);
nand U12192 (N_12192,N_10562,N_9182);
and U12193 (N_12193,N_11041,N_10238);
nand U12194 (N_12194,N_10630,N_11103);
nor U12195 (N_12195,N_11653,N_11112);
nand U12196 (N_12196,N_9294,N_11433);
nor U12197 (N_12197,N_11467,N_10504);
xor U12198 (N_12198,N_9125,N_11316);
or U12199 (N_12199,N_10104,N_9373);
and U12200 (N_12200,N_11209,N_11818);
nand U12201 (N_12201,N_9514,N_9757);
or U12202 (N_12202,N_11557,N_10978);
and U12203 (N_12203,N_10917,N_10444);
xor U12204 (N_12204,N_11902,N_9394);
nor U12205 (N_12205,N_10936,N_9823);
nand U12206 (N_12206,N_9427,N_10420);
nand U12207 (N_12207,N_10882,N_10548);
and U12208 (N_12208,N_10732,N_9574);
nand U12209 (N_12209,N_9816,N_11350);
nor U12210 (N_12210,N_11085,N_9644);
and U12211 (N_12211,N_10872,N_10358);
nor U12212 (N_12212,N_10010,N_11527);
or U12213 (N_12213,N_9428,N_10526);
nand U12214 (N_12214,N_10369,N_11652);
or U12215 (N_12215,N_9887,N_10467);
and U12216 (N_12216,N_10699,N_11194);
or U12217 (N_12217,N_9963,N_11828);
and U12218 (N_12218,N_10860,N_11266);
nand U12219 (N_12219,N_10298,N_10399);
nor U12220 (N_12220,N_9148,N_9484);
nor U12221 (N_12221,N_10308,N_10684);
and U12222 (N_12222,N_11062,N_11231);
nand U12223 (N_12223,N_10136,N_9958);
nand U12224 (N_12224,N_11721,N_10382);
and U12225 (N_12225,N_11688,N_9569);
nand U12226 (N_12226,N_11377,N_10641);
xor U12227 (N_12227,N_9774,N_9017);
or U12228 (N_12228,N_9708,N_11875);
or U12229 (N_12229,N_10478,N_11294);
nor U12230 (N_12230,N_9775,N_10592);
or U12231 (N_12231,N_9410,N_9284);
nand U12232 (N_12232,N_9653,N_11915);
or U12233 (N_12233,N_11830,N_10230);
xnor U12234 (N_12234,N_11366,N_10790);
and U12235 (N_12235,N_11696,N_10673);
and U12236 (N_12236,N_11838,N_10413);
nor U12237 (N_12237,N_9110,N_11494);
nand U12238 (N_12238,N_11496,N_9123);
or U12239 (N_12239,N_11291,N_11583);
xnor U12240 (N_12240,N_9079,N_11556);
and U12241 (N_12241,N_10307,N_11793);
or U12242 (N_12242,N_9183,N_11817);
nand U12243 (N_12243,N_9184,N_9029);
and U12244 (N_12244,N_9376,N_9469);
nor U12245 (N_12245,N_10232,N_11108);
nor U12246 (N_12246,N_11749,N_10580);
nor U12247 (N_12247,N_9922,N_11042);
and U12248 (N_12248,N_9665,N_11001);
or U12249 (N_12249,N_11788,N_11534);
or U12250 (N_12250,N_9781,N_11267);
or U12251 (N_12251,N_9988,N_9756);
nand U12252 (N_12252,N_11341,N_11633);
nand U12253 (N_12253,N_10667,N_10949);
nand U12254 (N_12254,N_11247,N_10629);
nand U12255 (N_12255,N_9924,N_11024);
nand U12256 (N_12256,N_11079,N_11420);
nor U12257 (N_12257,N_11639,N_9632);
or U12258 (N_12258,N_9840,N_10109);
nor U12259 (N_12259,N_11513,N_10391);
and U12260 (N_12260,N_9502,N_10789);
and U12261 (N_12261,N_9889,N_11580);
nand U12262 (N_12262,N_9936,N_11616);
nand U12263 (N_12263,N_10766,N_9769);
nand U12264 (N_12264,N_9950,N_11347);
nor U12265 (N_12265,N_9429,N_9129);
nand U12266 (N_12266,N_9340,N_11252);
and U12267 (N_12267,N_10256,N_9472);
or U12268 (N_12268,N_10785,N_10513);
or U12269 (N_12269,N_11761,N_11569);
nand U12270 (N_12270,N_10964,N_11207);
or U12271 (N_12271,N_10395,N_11179);
nand U12272 (N_12272,N_9667,N_11505);
or U12273 (N_12273,N_11173,N_9865);
nor U12274 (N_12274,N_10415,N_10610);
and U12275 (N_12275,N_9783,N_10608);
nand U12276 (N_12276,N_10631,N_11081);
nand U12277 (N_12277,N_11835,N_10169);
nand U12278 (N_12278,N_11167,N_9899);
nand U12279 (N_12279,N_10721,N_10865);
nor U12280 (N_12280,N_11945,N_10851);
nor U12281 (N_12281,N_11329,N_9704);
and U12282 (N_12282,N_11920,N_9248);
or U12283 (N_12283,N_9649,N_11281);
and U12284 (N_12284,N_11904,N_10421);
nand U12285 (N_12285,N_11177,N_11533);
nor U12286 (N_12286,N_9902,N_11736);
nand U12287 (N_12287,N_11577,N_10605);
and U12288 (N_12288,N_9424,N_9668);
or U12289 (N_12289,N_9877,N_9307);
and U12290 (N_12290,N_9034,N_9638);
or U12291 (N_12291,N_9059,N_10127);
and U12292 (N_12292,N_11687,N_9520);
and U12293 (N_12293,N_10615,N_9159);
nand U12294 (N_12294,N_9720,N_10094);
nor U12295 (N_12295,N_10984,N_9344);
xor U12296 (N_12296,N_11846,N_9478);
nor U12297 (N_12297,N_10916,N_11548);
nor U12298 (N_12298,N_10185,N_9217);
nor U12299 (N_12299,N_9130,N_11192);
and U12300 (N_12300,N_9554,N_10490);
and U12301 (N_12301,N_11808,N_9278);
xnor U12302 (N_12302,N_10877,N_11034);
or U12303 (N_12303,N_10784,N_11813);
xnor U12304 (N_12304,N_9505,N_9326);
and U12305 (N_12305,N_10708,N_9402);
or U12306 (N_12306,N_9039,N_11373);
nand U12307 (N_12307,N_10707,N_10660);
nor U12308 (N_12308,N_11215,N_10470);
or U12309 (N_12309,N_9820,N_11801);
and U12310 (N_12310,N_11600,N_10657);
nor U12311 (N_12311,N_9202,N_10672);
or U12312 (N_12312,N_9342,N_9095);
nand U12313 (N_12313,N_10899,N_10242);
or U12314 (N_12314,N_11762,N_9135);
xor U12315 (N_12315,N_10637,N_10543);
and U12316 (N_12316,N_9830,N_10354);
or U12317 (N_12317,N_9557,N_9337);
nand U12318 (N_12318,N_10816,N_11552);
nor U12319 (N_12319,N_10661,N_10815);
nor U12320 (N_12320,N_10468,N_11665);
nor U12321 (N_12321,N_11868,N_9818);
and U12322 (N_12322,N_11106,N_11620);
nand U12323 (N_12323,N_10034,N_9414);
nand U12324 (N_12324,N_9508,N_11502);
and U12325 (N_12325,N_10886,N_11865);
and U12326 (N_12326,N_9804,N_11969);
and U12327 (N_12327,N_11547,N_10587);
or U12328 (N_12328,N_11387,N_10332);
and U12329 (N_12329,N_10988,N_9698);
nor U12330 (N_12330,N_10156,N_9580);
or U12331 (N_12331,N_11236,N_10100);
nand U12332 (N_12332,N_10828,N_9028);
nor U12333 (N_12333,N_11495,N_11595);
nand U12334 (N_12334,N_11493,N_10007);
nor U12335 (N_12335,N_9204,N_10823);
and U12336 (N_12336,N_9829,N_10244);
nor U12337 (N_12337,N_11148,N_9977);
or U12338 (N_12338,N_10909,N_10950);
and U12339 (N_12339,N_11746,N_11628);
xor U12340 (N_12340,N_10680,N_9423);
and U12341 (N_12341,N_10167,N_10291);
and U12342 (N_12342,N_10457,N_10913);
nand U12343 (N_12343,N_11043,N_9507);
nor U12344 (N_12344,N_9516,N_11848);
or U12345 (N_12345,N_11343,N_9659);
xor U12346 (N_12346,N_9571,N_9283);
and U12347 (N_12347,N_11515,N_10731);
nand U12348 (N_12348,N_9647,N_10973);
nand U12349 (N_12349,N_10265,N_10696);
and U12350 (N_12350,N_11678,N_9603);
and U12351 (N_12351,N_9547,N_9280);
nor U12352 (N_12352,N_10887,N_11139);
or U12353 (N_12353,N_11689,N_9559);
and U12354 (N_12354,N_10843,N_9255);
nand U12355 (N_12355,N_11313,N_11344);
nor U12356 (N_12356,N_9957,N_11629);
or U12357 (N_12357,N_11798,N_10068);
xor U12358 (N_12358,N_10343,N_11951);
nand U12359 (N_12359,N_9700,N_11550);
or U12360 (N_12360,N_9910,N_9617);
or U12361 (N_12361,N_10666,N_11754);
nor U12362 (N_12362,N_10564,N_9465);
or U12363 (N_12363,N_10720,N_11385);
and U12364 (N_12364,N_9150,N_11153);
and U12365 (N_12365,N_9341,N_11949);
nand U12366 (N_12366,N_9244,N_9105);
nor U12367 (N_12367,N_10349,N_9444);
nand U12368 (N_12368,N_11698,N_9091);
or U12369 (N_12369,N_9971,N_9518);
nand U12370 (N_12370,N_10412,N_11122);
and U12371 (N_12371,N_9299,N_11244);
nor U12372 (N_12372,N_9925,N_10552);
nor U12373 (N_12373,N_11470,N_11221);
and U12374 (N_12374,N_10764,N_9949);
nand U12375 (N_12375,N_10016,N_11782);
nand U12376 (N_12376,N_10211,N_10793);
and U12377 (N_12377,N_11141,N_10831);
or U12378 (N_12378,N_10613,N_11458);
xor U12379 (N_12379,N_9611,N_10645);
or U12380 (N_12380,N_11305,N_11748);
or U12381 (N_12381,N_10626,N_9893);
nor U12382 (N_12382,N_11660,N_10956);
and U12383 (N_12383,N_11169,N_10173);
and U12384 (N_12384,N_11457,N_11237);
nor U12385 (N_12385,N_9645,N_9224);
nand U12386 (N_12386,N_11800,N_9646);
nor U12387 (N_12387,N_11571,N_10462);
nand U12388 (N_12388,N_9601,N_10869);
and U12389 (N_12389,N_10152,N_9515);
nand U12390 (N_12390,N_11284,N_10803);
and U12391 (N_12391,N_10890,N_11118);
and U12392 (N_12392,N_11887,N_10215);
nor U12393 (N_12393,N_10779,N_9013);
and U12394 (N_12394,N_9103,N_9509);
or U12395 (N_12395,N_9286,N_11302);
nand U12396 (N_12396,N_9247,N_11675);
and U12397 (N_12397,N_11662,N_11874);
nand U12398 (N_12398,N_10017,N_10814);
or U12399 (N_12399,N_11398,N_11312);
and U12400 (N_12400,N_10558,N_11211);
nand U12401 (N_12401,N_10316,N_11988);
and U12402 (N_12402,N_9964,N_9033);
and U12403 (N_12403,N_11993,N_9324);
xnor U12404 (N_12404,N_9069,N_10690);
nor U12405 (N_12405,N_10751,N_10542);
nor U12406 (N_12406,N_10780,N_9585);
nand U12407 (N_12407,N_10345,N_11938);
xor U12408 (N_12408,N_10288,N_11261);
nand U12409 (N_12409,N_9246,N_11483);
nand U12410 (N_12410,N_10374,N_9590);
nor U12411 (N_12411,N_10711,N_11443);
or U12412 (N_12412,N_9583,N_11590);
nand U12413 (N_12413,N_11625,N_11297);
nor U12414 (N_12414,N_10144,N_10411);
or U12415 (N_12415,N_9289,N_10750);
nand U12416 (N_12416,N_9088,N_10765);
or U12417 (N_12417,N_9588,N_11954);
or U12418 (N_12418,N_10346,N_9185);
nor U12419 (N_12419,N_11829,N_9623);
and U12420 (N_12420,N_9994,N_9627);
and U12421 (N_12421,N_10818,N_9929);
or U12422 (N_12422,N_11205,N_9560);
or U12423 (N_12423,N_11704,N_9397);
nand U12424 (N_12424,N_10182,N_11532);
or U12425 (N_12425,N_11528,N_10404);
and U12426 (N_12426,N_10376,N_11392);
nor U12427 (N_12427,N_11296,N_11608);
and U12428 (N_12428,N_9858,N_10088);
nand U12429 (N_12429,N_11840,N_11650);
xor U12430 (N_12430,N_9319,N_11359);
and U12431 (N_12431,N_10557,N_11976);
and U12432 (N_12432,N_11430,N_10350);
and U12433 (N_12433,N_11987,N_11503);
and U12434 (N_12434,N_11275,N_9062);
nand U12435 (N_12435,N_11589,N_9315);
nand U12436 (N_12436,N_10614,N_10820);
nand U12437 (N_12437,N_10214,N_9205);
or U12438 (N_12438,N_10501,N_11863);
xor U12439 (N_12439,N_9162,N_9261);
or U12440 (N_12440,N_9078,N_10322);
and U12441 (N_12441,N_10020,N_10105);
or U12442 (N_12442,N_9496,N_9064);
nor U12443 (N_12443,N_11399,N_11935);
and U12444 (N_12444,N_10870,N_11958);
nand U12445 (N_12445,N_9245,N_10052);
xor U12446 (N_12446,N_9512,N_11451);
and U12447 (N_12447,N_11986,N_10676);
and U12448 (N_12448,N_10791,N_9593);
nor U12449 (N_12449,N_11280,N_9635);
nand U12450 (N_12450,N_11853,N_10402);
nand U12451 (N_12451,N_9387,N_9196);
nor U12452 (N_12452,N_11060,N_9430);
nor U12453 (N_12453,N_11162,N_9380);
and U12454 (N_12454,N_11202,N_9549);
and U12455 (N_12455,N_11837,N_11539);
and U12456 (N_12456,N_10315,N_11172);
and U12457 (N_12457,N_11204,N_10773);
nand U12458 (N_12458,N_9699,N_9663);
xor U12459 (N_12459,N_9446,N_9537);
nand U12460 (N_12460,N_11322,N_9728);
nor U12461 (N_12461,N_10971,N_10409);
nand U12462 (N_12462,N_9093,N_11315);
or U12463 (N_12463,N_11475,N_10574);
nor U12464 (N_12464,N_10804,N_11324);
nand U12465 (N_12465,N_11369,N_10622);
nand U12466 (N_12466,N_10922,N_11479);
nand U12467 (N_12467,N_11997,N_11637);
and U12468 (N_12468,N_11586,N_9857);
nand U12469 (N_12469,N_10611,N_9368);
or U12470 (N_12470,N_9572,N_11050);
nor U12471 (N_12471,N_10025,N_9096);
nand U12472 (N_12472,N_9875,N_10295);
and U12473 (N_12473,N_10756,N_11488);
or U12474 (N_12474,N_9723,N_9228);
and U12475 (N_12475,N_11107,N_11955);
and U12476 (N_12476,N_11710,N_9032);
nor U12477 (N_12477,N_9814,N_9599);
nand U12478 (N_12478,N_9940,N_10908);
nor U12479 (N_12479,N_9586,N_10320);
and U12480 (N_12480,N_10051,N_9101);
or U12481 (N_12481,N_10845,N_11164);
or U12482 (N_12482,N_9867,N_9792);
nor U12483 (N_12483,N_9163,N_9923);
or U12484 (N_12484,N_10333,N_11456);
nand U12485 (N_12485,N_10586,N_11839);
nand U12486 (N_12486,N_11349,N_9295);
and U12487 (N_12487,N_9522,N_10179);
and U12488 (N_12488,N_11388,N_10604);
nor U12489 (N_12489,N_11517,N_10009);
and U12490 (N_12490,N_10759,N_10161);
or U12491 (N_12491,N_11200,N_11526);
nand U12492 (N_12492,N_10213,N_11567);
nor U12493 (N_12493,N_10153,N_11895);
or U12494 (N_12494,N_10129,N_10703);
and U12495 (N_12495,N_9226,N_9534);
and U12496 (N_12496,N_11025,N_10679);
nand U12497 (N_12497,N_10910,N_10683);
nand U12498 (N_12498,N_10071,N_9362);
and U12499 (N_12499,N_11602,N_9908);
xor U12500 (N_12500,N_10133,N_11445);
nor U12501 (N_12501,N_9144,N_10079);
and U12502 (N_12502,N_11751,N_9730);
nor U12503 (N_12503,N_11642,N_10874);
nor U12504 (N_12504,N_11368,N_9846);
nor U12505 (N_12505,N_10749,N_9597);
and U12506 (N_12506,N_9691,N_11730);
and U12507 (N_12507,N_9637,N_10653);
nand U12508 (N_12508,N_11380,N_11374);
nand U12509 (N_12509,N_11080,N_10015);
xor U12510 (N_12510,N_11760,N_11058);
and U12511 (N_12511,N_11905,N_10748);
nand U12512 (N_12512,N_9542,N_9024);
nor U12513 (N_12513,N_11944,N_9854);
nand U12514 (N_12514,N_11690,N_10113);
nand U12515 (N_12515,N_10342,N_10801);
or U12516 (N_12516,N_11094,N_10095);
xnor U12517 (N_12517,N_9657,N_10493);
and U12518 (N_12518,N_10270,N_9690);
or U12519 (N_12519,N_11896,N_11651);
and U12520 (N_12520,N_9995,N_9561);
nor U12521 (N_12521,N_9445,N_11285);
nand U12522 (N_12522,N_10717,N_11763);
nor U12523 (N_12523,N_11989,N_11016);
xnor U12524 (N_12524,N_11328,N_9071);
nor U12525 (N_12525,N_11588,N_9158);
and U12526 (N_12526,N_11140,N_10483);
nor U12527 (N_12527,N_9146,N_10753);
and U12528 (N_12528,N_10761,N_11018);
or U12529 (N_12529,N_9132,N_9782);
or U12530 (N_12530,N_10888,N_9799);
and U12531 (N_12531,N_11936,N_11464);
xor U12532 (N_12532,N_10560,N_11429);
nand U12533 (N_12533,N_9292,N_10609);
and U12534 (N_12534,N_9739,N_9529);
nand U12535 (N_12535,N_9086,N_10597);
and U12536 (N_12536,N_11082,N_11047);
nand U12537 (N_12537,N_10485,N_9251);
nand U12538 (N_12538,N_11666,N_11129);
and U12539 (N_12539,N_11703,N_9493);
or U12540 (N_12540,N_10072,N_9396);
xnor U12541 (N_12541,N_9227,N_11869);
or U12542 (N_12542,N_11959,N_9099);
nand U12543 (N_12543,N_9486,N_11814);
xnor U12544 (N_12544,N_10519,N_9314);
or U12545 (N_12545,N_10361,N_10334);
nor U12546 (N_12546,N_10508,N_9360);
nor U12547 (N_12547,N_11576,N_10368);
nand U12548 (N_12548,N_11643,N_11171);
nor U12549 (N_12549,N_10590,N_9837);
nor U12550 (N_12550,N_9845,N_11947);
or U12551 (N_12551,N_11594,N_10856);
or U12552 (N_12552,N_10534,N_11535);
or U12553 (N_12553,N_9868,N_10194);
xor U12554 (N_12554,N_11354,N_9441);
nor U12555 (N_12555,N_10252,N_9053);
nand U12556 (N_12556,N_10859,N_11069);
nand U12557 (N_12557,N_11638,N_11409);
or U12558 (N_12558,N_10771,N_10754);
or U12559 (N_12559,N_9176,N_9328);
or U12560 (N_12560,N_11317,N_10084);
nor U12561 (N_12561,N_11520,N_9113);
nand U12562 (N_12562,N_9956,N_9972);
or U12563 (N_12563,N_10891,N_11245);
and U12564 (N_12564,N_9080,N_10193);
xnor U12565 (N_12565,N_10570,N_9788);
or U12566 (N_12566,N_11855,N_9252);
nand U12567 (N_12567,N_9375,N_10031);
nand U12568 (N_12568,N_9981,N_9721);
or U12569 (N_12569,N_9754,N_9399);
or U12570 (N_12570,N_9802,N_10896);
or U12571 (N_12571,N_9628,N_9563);
and U12572 (N_12572,N_10318,N_9467);
or U12573 (N_12573,N_9641,N_9092);
nor U12574 (N_12574,N_11239,N_10317);
nand U12575 (N_12575,N_9349,N_10302);
nor U12576 (N_12576,N_9651,N_11086);
nor U12577 (N_12577,N_11845,N_9455);
xnor U12578 (N_12578,N_10691,N_9386);
and U12579 (N_12579,N_11787,N_9142);
and U12580 (N_12580,N_11790,N_10686);
nand U12581 (N_12581,N_11778,N_10117);
or U12582 (N_12582,N_10181,N_9810);
nand U12583 (N_12583,N_11145,N_11870);
and U12584 (N_12584,N_10830,N_10375);
nor U12585 (N_12585,N_11779,N_11859);
or U12586 (N_12586,N_9938,N_9000);
nor U12587 (N_12587,N_11937,N_10595);
and U12588 (N_12588,N_10788,N_10894);
and U12589 (N_12589,N_9111,N_11339);
or U12590 (N_12590,N_11056,N_10571);
and U12591 (N_12591,N_9450,N_10627);
nor U12592 (N_12592,N_11492,N_9921);
or U12593 (N_12593,N_11440,N_10632);
and U12594 (N_12594,N_10953,N_9216);
xnor U12595 (N_12595,N_9338,N_10235);
nor U12596 (N_12596,N_10942,N_10925);
nor U12597 (N_12597,N_9838,N_9525);
nor U12598 (N_12598,N_10812,N_10011);
or U12599 (N_12599,N_11894,N_10229);
nor U12600 (N_12600,N_11130,N_10044);
or U12601 (N_12601,N_10329,N_9983);
nand U12602 (N_12602,N_11462,N_11005);
xnor U12603 (N_12603,N_10253,N_10665);
xnor U12604 (N_12604,N_9933,N_10983);
and U12605 (N_12605,N_10180,N_11472);
and U12606 (N_12606,N_10567,N_9906);
nand U12607 (N_12607,N_10527,N_11768);
or U12608 (N_12608,N_10702,N_11017);
nor U12609 (N_12609,N_11708,N_9538);
nor U12610 (N_12610,N_10646,N_10163);
or U12611 (N_12611,N_11694,N_9157);
and U12612 (N_12612,N_11711,N_10995);
and U12613 (N_12613,N_11226,N_10006);
nor U12614 (N_12614,N_10359,N_9389);
nand U12615 (N_12615,N_11663,N_9391);
and U12616 (N_12616,N_10578,N_11742);
nand U12617 (N_12617,N_11797,N_10530);
or U12618 (N_12618,N_9931,N_10879);
or U12619 (N_12619,N_11538,N_11299);
nand U12620 (N_12620,N_10075,N_11498);
and U12621 (N_12621,N_9567,N_9795);
nand U12622 (N_12622,N_10108,N_9118);
and U12623 (N_12623,N_9007,N_9801);
nand U12624 (N_12624,N_11072,N_9106);
and U12625 (N_12625,N_10892,N_10082);
or U12626 (N_12626,N_11229,N_9454);
and U12627 (N_12627,N_10931,N_9688);
or U12628 (N_12628,N_11026,N_9147);
nand U12629 (N_12629,N_9166,N_10224);
nor U12630 (N_12630,N_10134,N_10225);
nand U12631 (N_12631,N_10625,N_9173);
and U12632 (N_12632,N_10980,N_9966);
and U12633 (N_12633,N_9238,N_9433);
nand U12634 (N_12634,N_9803,N_10159);
and U12635 (N_12635,N_11750,N_9717);
and U12636 (N_12636,N_10218,N_10234);
nor U12637 (N_12637,N_9729,N_11844);
and U12638 (N_12638,N_9584,N_9031);
nor U12639 (N_12639,N_11941,N_11683);
xnor U12640 (N_12640,N_11357,N_11725);
or U12641 (N_12641,N_10197,N_9592);
nor U12642 (N_12642,N_11862,N_11077);
xnor U12643 (N_12643,N_11559,N_9726);
nor U12644 (N_12644,N_9169,N_10259);
xor U12645 (N_12645,N_9558,N_9951);
and U12646 (N_12646,N_10515,N_10982);
nor U12647 (N_12647,N_10266,N_10839);
or U12648 (N_12648,N_10463,N_9749);
and U12649 (N_12649,N_9296,N_10554);
or U12650 (N_12650,N_10840,N_11033);
nor U12651 (N_12651,N_10960,N_9416);
or U12652 (N_12652,N_11852,N_9256);
nor U12653 (N_12653,N_11286,N_10414);
and U12654 (N_12654,N_11052,N_10652);
nor U12655 (N_12655,N_9460,N_10772);
nand U12656 (N_12656,N_11360,N_10023);
or U12657 (N_12657,N_9329,N_9174);
nor U12658 (N_12658,N_10489,N_11184);
or U12659 (N_12659,N_11700,N_10541);
and U12660 (N_12660,N_11648,N_11890);
xnor U12661 (N_12661,N_11757,N_9197);
nand U12662 (N_12662,N_9909,N_9881);
nand U12663 (N_12663,N_10154,N_10565);
nand U12664 (N_12664,N_10290,N_11410);
xnor U12665 (N_12665,N_9257,N_10321);
and U12666 (N_12666,N_9711,N_9786);
or U12667 (N_12667,N_11213,N_10377);
nand U12668 (N_12668,N_10427,N_11257);
nor U12669 (N_12669,N_9680,N_10852);
nor U12670 (N_12670,N_9528,N_11912);
nor U12671 (N_12671,N_11671,N_11723);
nor U12672 (N_12672,N_10593,N_10434);
nor U12673 (N_12673,N_9685,N_11158);
nor U12674 (N_12674,N_11489,N_10210);
nor U12675 (N_12675,N_10835,N_10955);
nand U12676 (N_12676,N_11522,N_9984);
and U12677 (N_12677,N_11334,N_10503);
or U12678 (N_12678,N_11487,N_9320);
or U12679 (N_12679,N_11031,N_11088);
xor U12680 (N_12680,N_10267,N_10937);
nand U12681 (N_12681,N_11776,N_9083);
nor U12682 (N_12682,N_10762,N_11715);
nand U12683 (N_12683,N_10758,N_11676);
xnor U12684 (N_12684,N_9918,N_11396);
nand U12685 (N_12685,N_10269,N_9962);
nor U12686 (N_12686,N_10001,N_9552);
xnor U12687 (N_12687,N_9869,N_11767);
nand U12688 (N_12688,N_9661,N_11545);
and U12689 (N_12689,N_9939,N_10889);
xnor U12690 (N_12690,N_9141,N_10043);
xor U12691 (N_12691,N_9090,N_10257);
nand U12692 (N_12692,N_9740,N_10741);
or U12693 (N_12693,N_11499,N_10078);
or U12694 (N_12694,N_9553,N_9070);
nor U12695 (N_12695,N_9587,N_10183);
nor U12696 (N_12696,N_9692,N_9102);
nand U12697 (N_12697,N_11230,N_10301);
or U12698 (N_12698,N_10969,N_9170);
and U12699 (N_12699,N_10122,N_9432);
and U12700 (N_12700,N_9347,N_11195);
or U12701 (N_12701,N_11065,N_10822);
nand U12702 (N_12702,N_11971,N_11598);
nand U12703 (N_12703,N_10365,N_11925);
xor U12704 (N_12704,N_10436,N_10651);
nand U12705 (N_12705,N_11996,N_10142);
and U12706 (N_12706,N_11612,N_10687);
nand U12707 (N_12707,N_11174,N_9631);
or U12708 (N_12708,N_11181,N_9656);
or U12709 (N_12709,N_10975,N_10866);
and U12710 (N_12710,N_9275,N_11975);
or U12711 (N_12711,N_11952,N_11784);
or U12712 (N_12712,N_10458,N_10486);
or U12713 (N_12713,N_11789,N_10070);
and U12714 (N_12714,N_11858,N_11820);
nor U12715 (N_12715,N_10722,N_11995);
or U12716 (N_12716,N_9207,N_10512);
or U12717 (N_12717,N_11240,N_11278);
nor U12718 (N_12718,N_9510,N_11111);
xor U12719 (N_12719,N_9108,N_9369);
xor U12720 (N_12720,N_11827,N_9250);
or U12721 (N_12721,N_11319,N_9828);
xor U12722 (N_12722,N_10221,N_10396);
or U12723 (N_12723,N_9011,N_9530);
and U12724 (N_12724,N_11501,N_11635);
and U12725 (N_12725,N_11884,N_10638);
or U12726 (N_12726,N_10972,N_9874);
and U12727 (N_12727,N_10339,N_10591);
xnor U12728 (N_12728,N_11622,N_11919);
or U12729 (N_12729,N_9018,N_11731);
nand U12730 (N_12730,N_9683,N_11717);
nand U12731 (N_12731,N_10195,N_9009);
nand U12732 (N_12732,N_11474,N_9621);
nand U12733 (N_12733,N_11573,N_11799);
xnor U12734 (N_12734,N_11189,N_10905);
and U12735 (N_12735,N_9594,N_10338);
or U12736 (N_12736,N_11417,N_11500);
or U12737 (N_12737,N_11991,N_9061);
or U12738 (N_12738,N_10868,N_11269);
or U12739 (N_12739,N_10809,N_10208);
nand U12740 (N_12740,N_9770,N_11518);
xor U12741 (N_12741,N_10083,N_11438);
nand U12742 (N_12742,N_11059,N_9625);
or U12743 (N_12743,N_9859,N_9866);
nor U12744 (N_12744,N_9264,N_11428);
nand U12745 (N_12745,N_9678,N_10726);
nor U12746 (N_12746,N_9883,N_11471);
nand U12747 (N_12747,N_9282,N_10979);
or U12748 (N_12748,N_9285,N_11753);
nor U12749 (N_12749,N_9260,N_10209);
and U12750 (N_12750,N_11156,N_11525);
nand U12751 (N_12751,N_10744,N_11714);
or U12752 (N_12752,N_9335,N_10927);
or U12753 (N_12753,N_10176,N_10550);
xnor U12754 (N_12754,N_9968,N_10164);
nor U12755 (N_12755,N_9003,N_9975);
nand U12756 (N_12756,N_10438,N_11326);
xor U12757 (N_12757,N_10373,N_9466);
or U12758 (N_12758,N_9745,N_11982);
nand U12759 (N_12759,N_9181,N_10416);
nand U12760 (N_12760,N_10767,N_10177);
nand U12761 (N_12761,N_9480,N_9666);
or U12762 (N_12762,N_10944,N_10855);
nor U12763 (N_12763,N_9221,N_9703);
or U12764 (N_12764,N_11713,N_10027);
and U12765 (N_12765,N_9459,N_9642);
nand U12766 (N_12766,N_11288,N_10058);
nand U12767 (N_12767,N_10065,N_9709);
nand U12768 (N_12768,N_10528,N_9051);
and U12769 (N_12769,N_10740,N_10157);
nor U12770 (N_12770,N_9761,N_11407);
nor U12771 (N_12771,N_10202,N_11159);
nand U12772 (N_12772,N_10985,N_10502);
xor U12773 (N_12773,N_11248,N_10569);
nand U12774 (N_12774,N_10549,N_11712);
nand U12775 (N_12775,N_10206,N_9750);
nor U12776 (N_12776,N_9201,N_9897);
nand U12777 (N_12777,N_10989,N_10618);
and U12778 (N_12778,N_11105,N_9230);
nand U12779 (N_12779,N_9040,N_11878);
nor U12780 (N_12780,N_9138,N_10426);
xor U12781 (N_12781,N_11783,N_11468);
nand U12782 (N_12782,N_11921,N_11791);
or U12783 (N_12783,N_10535,N_9751);
or U12784 (N_12784,N_9974,N_10330);
or U12785 (N_12785,N_10678,N_10271);
xor U12786 (N_12786,N_9888,N_11587);
and U12787 (N_12787,N_11098,N_10030);
nor U12788 (N_12788,N_11752,N_10730);
and U12789 (N_12789,N_9036,N_10616);
nand U12790 (N_12790,N_9054,N_11234);
nand U12791 (N_12791,N_10688,N_9119);
or U12792 (N_12792,N_11253,N_9578);
or U12793 (N_12793,N_9213,N_9073);
or U12794 (N_12794,N_10086,N_10060);
nand U12795 (N_12795,N_11218,N_11899);
and U12796 (N_12796,N_10004,N_9762);
and U12797 (N_12797,N_9942,N_10553);
or U12798 (N_12798,N_9524,N_10066);
nor U12799 (N_12799,N_10160,N_11143);
and U12800 (N_12800,N_10524,N_10362);
xor U12801 (N_12801,N_11824,N_11745);
and U12802 (N_12802,N_9847,N_10294);
nor U12803 (N_12803,N_9180,N_11336);
and U12804 (N_12804,N_11273,N_10216);
and U12805 (N_12805,N_9464,N_10032);
or U12806 (N_12806,N_11461,N_10862);
nand U12807 (N_12807,N_9920,N_9742);
or U12808 (N_12808,N_11546,N_11078);
nand U12809 (N_12809,N_9848,N_11271);
or U12810 (N_12810,N_9764,N_9365);
or U12811 (N_12811,N_9634,N_11379);
nand U12812 (N_12812,N_9477,N_9297);
or U12813 (N_12813,N_10893,N_11537);
nand U12814 (N_12814,N_9892,N_11674);
and U12815 (N_12815,N_9996,N_9087);
nand U12816 (N_12816,N_10273,N_11425);
nand U12817 (N_12817,N_10048,N_11012);
or U12818 (N_12818,N_11282,N_9331);
nor U12819 (N_12819,N_9602,N_9787);
nand U12820 (N_12820,N_10472,N_10810);
xor U12821 (N_12821,N_9177,N_10757);
nor U12822 (N_12822,N_9744,N_11180);
nand U12823 (N_12823,N_10734,N_10370);
or U12824 (N_12824,N_9047,N_9481);
nor U12825 (N_12825,N_9702,N_10465);
or U12826 (N_12826,N_11873,N_9330);
and U12827 (N_12827,N_9215,N_9468);
nor U12828 (N_12828,N_10643,N_11621);
or U12829 (N_12829,N_10431,N_11950);
nand U12830 (N_12830,N_11693,N_11486);
nor U12831 (N_12831,N_11132,N_10996);
nand U12832 (N_12832,N_10654,N_9989);
nand U12833 (N_12833,N_9081,N_10885);
and U12834 (N_12834,N_9640,N_11222);
and U12835 (N_12835,N_9457,N_11061);
nor U12836 (N_12836,N_11565,N_10062);
and U12837 (N_12837,N_11805,N_11833);
or U12838 (N_12838,N_11049,N_10263);
xnor U12839 (N_12839,N_11716,N_11413);
and U12840 (N_12840,N_9916,N_10344);
nor U12841 (N_12841,N_11243,N_10837);
nand U12842 (N_12842,N_10572,N_11473);
xor U12843 (N_12843,N_9379,N_9610);
nor U12844 (N_12844,N_10706,N_9021);
xnor U12845 (N_12845,N_9872,N_9841);
or U12846 (N_12846,N_11857,N_10763);
xor U12847 (N_12847,N_11685,N_11054);
and U12848 (N_12848,N_10090,N_11764);
or U12849 (N_12849,N_11564,N_10055);
or U12850 (N_12850,N_11967,N_11020);
nand U12851 (N_12851,N_9772,N_9312);
and U12852 (N_12852,N_9735,N_10739);
nor U12853 (N_12853,N_10401,N_10328);
and U12854 (N_12854,N_11370,N_11431);
and U12855 (N_12855,N_11466,N_10250);
nand U12856 (N_12856,N_9352,N_9350);
or U12857 (N_12857,N_9813,N_11449);
and U12858 (N_12858,N_11699,N_10921);
or U12859 (N_12859,N_9449,N_11023);
or U12860 (N_12860,N_11003,N_10112);
nor U12861 (N_12861,N_9439,N_11572);
nor U12862 (N_12862,N_9043,N_9808);
and U12863 (N_12863,N_10091,N_10520);
and U12864 (N_12864,N_10451,N_11634);
nor U12865 (N_12865,N_10802,N_11332);
and U12866 (N_12866,N_9864,N_9609);
and U12867 (N_12867,N_11030,N_9716);
nand U12868 (N_12868,N_10057,N_9417);
or U12869 (N_12869,N_11964,N_11292);
xnor U12870 (N_12870,N_10871,N_9126);
nor U12871 (N_12871,N_10063,N_9240);
and U12872 (N_12872,N_11604,N_9991);
or U12873 (N_12873,N_9100,N_9543);
xnor U12874 (N_12874,N_10718,N_10178);
xnor U12875 (N_12875,N_11979,N_11469);
nor U12876 (N_12876,N_10647,N_11448);
or U12877 (N_12877,N_11251,N_11765);
nand U12878 (N_12878,N_10387,N_9879);
nand U12879 (N_12879,N_10963,N_11115);
or U12880 (N_12880,N_10324,N_9200);
and U12881 (N_12881,N_9934,N_11084);
or U12882 (N_12882,N_10037,N_10698);
and U12883 (N_12883,N_11568,N_10408);
nand U12884 (N_12884,N_10858,N_11722);
or U12885 (N_12885,N_9259,N_9253);
nor U12886 (N_12886,N_10255,N_11150);
or U12887 (N_12887,N_11203,N_11337);
nand U12888 (N_12888,N_11160,N_9521);
and U12889 (N_12889,N_11706,N_10174);
nand U12890 (N_12890,N_9896,N_10306);
nor U12891 (N_12891,N_9954,N_10059);
or U12892 (N_12892,N_9696,N_9833);
and U12893 (N_12893,N_10967,N_10669);
nor U12894 (N_12894,N_10623,N_10498);
or U12895 (N_12895,N_9235,N_11946);
nand U12896 (N_12896,N_10475,N_9363);
and U12897 (N_12897,N_9605,N_11561);
xnor U12898 (N_12898,N_11346,N_9682);
xnor U12899 (N_12899,N_9346,N_11719);
or U12900 (N_12900,N_10313,N_9650);
or U12901 (N_12901,N_11807,N_11435);
nor U12902 (N_12902,N_9636,N_10488);
nor U12903 (N_12903,N_9384,N_11816);
or U12904 (N_12904,N_11738,N_10275);
and U12905 (N_12905,N_10260,N_10825);
xnor U12906 (N_12906,N_10579,N_9482);
nand U12907 (N_12907,N_11367,N_10162);
nor U12908 (N_12908,N_11113,N_11630);
nand U12909 (N_12909,N_9544,N_11777);
nand U12910 (N_12910,N_10219,N_11224);
nand U12911 (N_12911,N_11734,N_10064);
nand U12912 (N_12912,N_11283,N_9596);
and U12913 (N_12913,N_11185,N_9619);
and U12914 (N_12914,N_11596,N_10903);
nand U12915 (N_12915,N_10461,N_11142);
and U12916 (N_12916,N_9140,N_11238);
and U12917 (N_12917,N_11720,N_11599);
nand U12918 (N_12918,N_9715,N_9395);
nand U12919 (N_12919,N_11804,N_9356);
and U12920 (N_12920,N_11802,N_10406);
nand U12921 (N_12921,N_11766,N_11127);
nand U12922 (N_12922,N_11806,N_11897);
or U12923 (N_12923,N_10725,N_11914);
and U12924 (N_12924,N_9550,N_9411);
and U12925 (N_12925,N_9491,N_9025);
or U12926 (N_12926,N_11446,N_10130);
xnor U12927 (N_12927,N_10599,N_10042);
nand U12928 (N_12928,N_10537,N_11999);
or U12929 (N_12929,N_10116,N_10808);
nor U12930 (N_12930,N_10289,N_11307);
and U12931 (N_12931,N_9403,N_11880);
xnor U12932 (N_12932,N_11046,N_9825);
and U12933 (N_12933,N_9390,N_10035);
nor U12934 (N_12934,N_10397,N_10533);
and U12935 (N_12935,N_9321,N_11871);
and U12936 (N_12936,N_11670,N_9037);
or U12937 (N_12937,N_11314,N_11154);
nor U12938 (N_12938,N_11293,N_9016);
and U12939 (N_12939,N_10381,N_11119);
or U12940 (N_12940,N_11258,N_11116);
nand U12941 (N_12941,N_11551,N_10236);
nand U12942 (N_12942,N_11138,N_9658);
or U12943 (N_12943,N_11414,N_10634);
nor U12944 (N_12944,N_11432,N_10714);
nand U12945 (N_12945,N_9189,N_9311);
or U12946 (N_12946,N_9856,N_9401);
nand U12947 (N_12947,N_11161,N_9209);
or U12948 (N_12948,N_9456,N_9339);
nor U12949 (N_12949,N_11338,N_9556);
nand U12950 (N_12950,N_10829,N_11592);
or U12951 (N_12951,N_11929,N_11117);
or U12952 (N_12952,N_10585,N_11092);
or U12953 (N_12953,N_10873,N_9743);
nand U12954 (N_12954,N_10459,N_9179);
and U12955 (N_12955,N_10327,N_10582);
nor U12956 (N_12956,N_10449,N_10867);
or U12957 (N_12957,N_9633,N_10125);
xor U12958 (N_12958,N_10961,N_11361);
nand U12959 (N_12959,N_11614,N_10881);
and U12960 (N_12960,N_9831,N_11027);
nand U12961 (N_12961,N_10312,N_10906);
or U12962 (N_12962,N_11705,N_9765);
and U12963 (N_12963,N_10385,N_11365);
and U12964 (N_12964,N_10246,N_10965);
and U12965 (N_12965,N_11885,N_10239);
xnor U12966 (N_12966,N_11623,N_11697);
nand U12967 (N_12967,N_9827,N_9734);
nand U12968 (N_12968,N_11769,N_9199);
or U12969 (N_12969,N_11977,N_9767);
and U12970 (N_12970,N_11163,N_9843);
and U12971 (N_12971,N_9143,N_10151);
and U12972 (N_12972,N_11831,N_10832);
nor U12973 (N_12973,N_10594,N_9741);
or U12974 (N_12974,N_9738,N_10147);
or U12975 (N_12975,N_10047,N_11707);
nand U12976 (N_12976,N_9023,N_11510);
nor U12977 (N_12977,N_11320,N_11555);
and U12978 (N_12978,N_11810,N_11220);
nor U12979 (N_12979,N_11497,N_11542);
or U12980 (N_12980,N_9850,N_10264);
and U12981 (N_12981,N_9067,N_10795);
nor U12982 (N_12982,N_11351,N_11342);
nand U12983 (N_12983,N_9891,N_9672);
nor U12984 (N_12984,N_10081,N_9826);
nand U12985 (N_12985,N_9236,N_9458);
nand U12986 (N_12986,N_10577,N_10311);
and U12987 (N_12987,N_10435,N_11819);
xnor U12988 (N_12988,N_9548,N_10417);
xor U12989 (N_12989,N_11893,N_10393);
nand U12990 (N_12990,N_11391,N_10928);
nand U12991 (N_12991,N_10668,N_9821);
nand U12992 (N_12992,N_9004,N_9461);
nand U12993 (N_12993,N_10948,N_10175);
nor U12994 (N_12994,N_9871,N_11521);
and U12995 (N_12995,N_9490,N_11613);
or U12996 (N_12996,N_9777,N_9046);
and U12997 (N_12997,N_10496,N_11785);
xor U12998 (N_12998,N_11984,N_11773);
nor U12999 (N_12999,N_10103,N_11744);
or U13000 (N_13000,N_10510,N_11673);
nor U13001 (N_13001,N_10433,N_9056);
or U13002 (N_13002,N_10838,N_10190);
and U13003 (N_13003,N_9243,N_10849);
nand U13004 (N_13004,N_9305,N_11067);
nand U13005 (N_13005,N_11114,N_10196);
xnor U13006 (N_13006,N_11983,N_10911);
or U13007 (N_13007,N_10497,N_11478);
nand U13008 (N_13008,N_9759,N_10833);
nand U13009 (N_13009,N_10425,N_11681);
or U13010 (N_13010,N_10805,N_10448);
and U13011 (N_13011,N_11646,N_9359);
nand U13012 (N_13012,N_10670,N_10929);
nand U13013 (N_13013,N_9630,N_11120);
and U13014 (N_13014,N_9780,N_11903);
nor U13015 (N_13015,N_11940,N_11879);
and U13016 (N_13016,N_11759,N_9355);
and U13017 (N_13017,N_10337,N_10674);
and U13018 (N_13018,N_9932,N_11095);
or U13019 (N_13019,N_10268,N_11304);
nand U13020 (N_13020,N_9137,N_10861);
nor U13021 (N_13021,N_11850,N_11383);
nor U13022 (N_13022,N_11636,N_11382);
nor U13023 (N_13023,N_10146,N_9287);
nand U13024 (N_13024,N_9109,N_10900);
and U13025 (N_13025,N_11418,N_11301);
nor U13026 (N_13026,N_11166,N_11401);
nor U13027 (N_13027,N_10442,N_9366);
nand U13028 (N_13028,N_11165,N_10959);
nand U13029 (N_13029,N_11617,N_9664);
and U13030 (N_13030,N_10466,N_9993);
or U13031 (N_13031,N_11290,N_9443);
nor U13032 (N_13032,N_9431,N_10994);
nor U13033 (N_13033,N_10918,N_9714);
nand U13034 (N_13034,N_10158,N_10247);
or U13035 (N_13035,N_11219,N_9768);
nor U13036 (N_13036,N_11459,N_10477);
or U13037 (N_13037,N_9849,N_9948);
or U13038 (N_13038,N_9564,N_11051);
nor U13039 (N_13039,N_11019,N_9785);
and U13040 (N_13040,N_11644,N_10028);
and U13041 (N_13041,N_9412,N_11770);
nor U13042 (N_13042,N_10518,N_10139);
xor U13043 (N_13043,N_9405,N_11412);
or U13044 (N_13044,N_10806,N_11048);
xor U13045 (N_13045,N_11659,N_9980);
and U13046 (N_13046,N_9562,N_11393);
and U13047 (N_13047,N_11957,N_9164);
nand U13048 (N_13048,N_10682,N_10336);
and U13049 (N_13049,N_11035,N_9383);
nor U13050 (N_13050,N_9855,N_10279);
nor U13051 (N_13051,N_11607,N_9807);
xnor U13052 (N_13052,N_10675,N_11216);
or U13053 (N_13053,N_9268,N_11524);
nor U13054 (N_13054,N_10875,N_11724);
nand U13055 (N_13055,N_11891,N_9076);
nor U13056 (N_13056,N_11453,N_9901);
and U13057 (N_13057,N_9817,N_11090);
nand U13058 (N_13058,N_11070,N_11263);
nor U13059 (N_13059,N_11454,N_11994);
nor U13060 (N_13060,N_9309,N_11044);
xnor U13061 (N_13061,N_11147,N_9068);
nand U13062 (N_13062,N_9731,N_10500);
and U13063 (N_13063,N_9323,N_9784);
or U13064 (N_13064,N_10096,N_11781);
nand U13065 (N_13065,N_11186,N_10410);
or U13066 (N_13066,N_11631,N_10544);
nand U13067 (N_13067,N_9900,N_9272);
or U13068 (N_13068,N_9448,N_10299);
and U13069 (N_13069,N_9304,N_11348);
and U13070 (N_13070,N_11924,N_10522);
nand U13071 (N_13071,N_9504,N_10277);
xor U13072 (N_13072,N_9225,N_9839);
nor U13073 (N_13073,N_11402,N_10817);
or U13074 (N_13074,N_9293,N_11876);
nor U13075 (N_13075,N_11864,N_11942);
or U13076 (N_13076,N_11008,N_9959);
nand U13077 (N_13077,N_9048,N_9422);
nand U13078 (N_13078,N_10305,N_11661);
nand U13079 (N_13079,N_11212,N_9973);
nand U13080 (N_13080,N_10957,N_9107);
nor U13081 (N_13081,N_9998,N_10649);
nand U13082 (N_13082,N_11053,N_10372);
nor U13083 (N_13083,N_11241,N_9809);
xnor U13084 (N_13084,N_10297,N_10360);
and U13085 (N_13085,N_9407,N_11424);
and U13086 (N_13086,N_11821,N_10581);
nand U13087 (N_13087,N_11376,N_11183);
nand U13088 (N_13088,N_9060,N_11892);
nor U13089 (N_13089,N_11100,N_9404);
nor U13090 (N_13090,N_10278,N_10254);
and U13091 (N_13091,N_11152,N_10993);
xnor U13092 (N_13092,N_11910,N_10464);
nand U13093 (N_13093,N_10056,N_10441);
nor U13094 (N_13094,N_10943,N_9589);
and U13095 (N_13095,N_10656,N_11641);
or U13096 (N_13096,N_11718,N_9191);
or U13097 (N_13097,N_10456,N_10296);
nand U13098 (N_13098,N_9517,N_10636);
xnor U13099 (N_13099,N_10635,N_9878);
or U13100 (N_13100,N_11861,N_11187);
and U13101 (N_13101,N_9905,N_9382);
xor U13102 (N_13102,N_9541,N_10992);
xnor U13103 (N_13103,N_10912,N_9175);
xor U13104 (N_13104,N_11358,N_9836);
nand U13105 (N_13105,N_11632,N_11295);
and U13106 (N_13106,N_10367,N_10523);
and U13107 (N_13107,N_11603,N_9139);
or U13108 (N_13108,N_11795,N_9254);
nand U13109 (N_13109,N_10768,N_10137);
and U13110 (N_13110,N_9442,N_9400);
and U13111 (N_13111,N_10774,N_9669);
nor U13112 (N_13112,N_11658,N_9495);
or U13113 (N_13113,N_9928,N_10834);
nor U13114 (N_13114,N_9149,N_10045);
nor U13115 (N_13115,N_9050,N_9222);
xnor U13116 (N_13116,N_11170,N_9677);
and U13117 (N_13117,N_11490,N_9452);
and U13118 (N_13118,N_10842,N_9348);
and U13119 (N_13119,N_11176,N_9098);
nor U13120 (N_13120,N_10455,N_10628);
nor U13121 (N_13121,N_11529,N_11091);
or U13122 (N_13122,N_9084,N_9136);
nand U13123 (N_13123,N_10606,N_10107);
nand U13124 (N_13124,N_11447,N_9660);
and U13125 (N_13125,N_9188,N_9582);
and U13126 (N_13126,N_9232,N_10715);
and U13127 (N_13127,N_9760,N_9265);
and U13128 (N_13128,N_11331,N_9392);
and U13129 (N_13129,N_9451,N_10583);
and U13130 (N_13130,N_10021,N_10863);
nor U13131 (N_13131,N_10940,N_9624);
nor U13132 (N_13132,N_10192,N_9607);
nor U13133 (N_13133,N_9124,N_9752);
nor U13134 (N_13134,N_11980,N_10309);
or U13135 (N_13135,N_9190,N_9005);
nor U13136 (N_13136,N_9852,N_10954);
or U13137 (N_13137,N_9955,N_9615);
xnor U13138 (N_13138,N_11375,N_10121);
nand U13139 (N_13139,N_11849,N_11071);
and U13140 (N_13140,N_11953,N_10705);
nor U13141 (N_13141,N_10249,N_9713);
nor U13142 (N_13142,N_9832,N_10392);
nor U13143 (N_13143,N_10794,N_9042);
or U13144 (N_13144,N_11508,N_10743);
nor U13145 (N_13145,N_10419,N_9606);
and U13146 (N_13146,N_11411,N_11038);
or U13147 (N_13147,N_11000,N_10719);
or U13148 (N_13148,N_9882,N_9152);
and U13149 (N_13149,N_11939,N_11426);
nand U13150 (N_13150,N_11815,N_10729);
nor U13151 (N_13151,N_11133,N_10692);
or U13152 (N_13152,N_10248,N_9919);
or U13153 (N_13153,N_11260,N_11553);
or U13154 (N_13154,N_11193,N_11089);
nand U13155 (N_13155,N_11010,N_11512);
nor U13156 (N_13156,N_11847,N_11743);
nand U13157 (N_13157,N_9506,N_11362);
xnor U13158 (N_13158,N_10106,N_10013);
nor U13159 (N_13159,N_11276,N_10386);
nand U13160 (N_13160,N_9231,N_10258);
and U13161 (N_13161,N_10716,N_10847);
or U13162 (N_13162,N_9904,N_9154);
or U13163 (N_13163,N_11131,N_10326);
nor U13164 (N_13164,N_10492,N_9483);
and U13165 (N_13165,N_9406,N_9075);
or U13166 (N_13166,N_10383,N_11615);
xor U13167 (N_13167,N_9353,N_11854);
nand U13168 (N_13168,N_10990,N_9546);
nor U13169 (N_13169,N_11872,N_9263);
xor U13170 (N_13170,N_9579,N_10148);
nor U13171 (N_13171,N_11794,N_10141);
nor U13172 (N_13172,N_10997,N_10138);
nor U13173 (N_13173,N_10474,N_11055);
or U13174 (N_13174,N_11809,N_9689);
nor U13175 (N_13175,N_11482,N_10700);
or U13176 (N_13176,N_9145,N_9354);
xnor U13177 (N_13177,N_10556,N_11306);
and U13178 (N_13178,N_9229,N_10904);
or U13179 (N_13179,N_9116,N_9371);
or U13180 (N_13180,N_10243,N_11437);
nand U13181 (N_13181,N_10283,N_10617);
and U13182 (N_13182,N_9044,N_11679);
nand U13183 (N_13183,N_11330,N_11898);
nand U13184 (N_13184,N_9027,N_9489);
nor U13185 (N_13185,N_10440,N_11477);
or U13186 (N_13186,N_11825,N_10538);
or U13187 (N_13187,N_9462,N_11246);
nand U13188 (N_13188,N_11068,N_11124);
or U13189 (N_13189,N_10479,N_10991);
nand U13190 (N_13190,N_10539,N_9697);
xor U13191 (N_13191,N_11882,N_10460);
nor U13192 (N_13192,N_11386,N_9378);
or U13193 (N_13193,N_11321,N_10939);
and U13194 (N_13194,N_11415,N_10445);
nand U13195 (N_13195,N_9045,N_9551);
nor U13196 (N_13196,N_10061,N_9415);
and U13197 (N_13197,N_11395,N_10482);
xor U13198 (N_13198,N_9503,N_10481);
or U13199 (N_13199,N_11531,N_11188);
nand U13200 (N_13200,N_11692,N_9178);
or U13201 (N_13201,N_9237,N_10110);
or U13202 (N_13202,N_10335,N_9239);
and U13203 (N_13203,N_10089,N_10976);
nand U13204 (N_13204,N_10101,N_11197);
nor U13205 (N_13205,N_11323,N_11917);
nor U13206 (N_13206,N_10659,N_11452);
xor U13207 (N_13207,N_11371,N_9435);
nor U13208 (N_13208,N_10201,N_11965);
or U13209 (N_13209,N_9947,N_10620);
nand U13210 (N_13210,N_11345,N_10282);
nand U13211 (N_13211,N_10119,N_11287);
nor U13212 (N_13212,N_9343,N_9684);
and U13213 (N_13213,N_11611,N_11735);
nor U13214 (N_13214,N_9161,N_10026);
and U13215 (N_13215,N_11669,N_9418);
nor U13216 (N_13216,N_10933,N_10476);
and U13217 (N_13217,N_10046,N_10300);
nor U13218 (N_13218,N_11423,N_9941);
or U13219 (N_13219,N_10509,N_11931);
or U13220 (N_13220,N_11593,N_9870);
or U13221 (N_13221,N_9673,N_10671);
nor U13222 (N_13222,N_11381,N_10484);
and U13223 (N_13223,N_10650,N_11908);
and U13224 (N_13224,N_10077,N_9398);
nand U13225 (N_13225,N_10573,N_11626);
or U13226 (N_13226,N_9674,N_10977);
or U13227 (N_13227,N_10310,N_11352);
nand U13228 (N_13228,N_10132,N_9133);
nand U13229 (N_13229,N_11541,N_9943);
and U13230 (N_13230,N_11228,N_11972);
nand U13231 (N_13231,N_10237,N_9219);
nand U13232 (N_13232,N_11780,N_10713);
nor U13233 (N_13233,N_10423,N_11916);
nor U13234 (N_13234,N_9719,N_9242);
nor U13235 (N_13235,N_9797,N_10303);
nor U13236 (N_13236,N_10600,N_9082);
nor U13237 (N_13237,N_11101,N_10546);
and U13238 (N_13238,N_11109,N_11585);
nor U13239 (N_13239,N_9945,N_10826);
and U13240 (N_13240,N_9990,N_10155);
xnor U13241 (N_13241,N_10018,N_9019);
nand U13242 (N_13242,N_11906,N_9127);
nor U13243 (N_13243,N_10398,N_11973);
or U13244 (N_13244,N_11455,N_9186);
nor U13245 (N_13245,N_11136,N_9262);
nor U13246 (N_13246,N_10934,N_10284);
nor U13247 (N_13247,N_9985,N_11691);
nand U13248 (N_13248,N_11196,N_11403);
or U13249 (N_13249,N_11514,N_9705);
nor U13250 (N_13250,N_10776,N_10920);
and U13251 (N_13251,N_11021,N_10319);
or U13252 (N_13252,N_9214,N_10261);
and U13253 (N_13253,N_10118,N_9361);
nor U13254 (N_13254,N_9863,N_9805);
nor U13255 (N_13255,N_9074,N_9494);
xor U13256 (N_13256,N_9058,N_9595);
nand U13257 (N_13257,N_11664,N_9020);
and U13258 (N_13258,N_11355,N_10469);
and U13259 (N_13259,N_11922,N_11963);
or U13260 (N_13260,N_9687,N_11434);
or U13261 (N_13261,N_9693,N_10799);
xnor U13262 (N_13262,N_9223,N_9912);
and U13263 (N_13263,N_11627,N_10353);
nand U13264 (N_13264,N_11310,N_10168);
or U13265 (N_13265,N_11465,N_9171);
nand U13266 (N_13266,N_9570,N_11654);
or U13267 (N_13267,N_9233,N_10227);
nand U13268 (N_13268,N_11327,N_9812);
nand U13269 (N_13269,N_9873,N_10405);
or U13270 (N_13270,N_9707,N_11277);
nand U13271 (N_13271,N_10074,N_9187);
or U13272 (N_13272,N_10947,N_9475);
nor U13273 (N_13273,N_10584,N_11093);
nor U13274 (N_13274,N_10658,N_9488);
nand U13275 (N_13275,N_10728,N_9322);
nand U13276 (N_13276,N_9935,N_9566);
nor U13277 (N_13277,N_10276,N_11318);
or U13278 (N_13278,N_10223,N_9269);
or U13279 (N_13279,N_10203,N_11609);
xnor U13280 (N_13280,N_11740,N_10693);
and U13281 (N_13281,N_10184,N_11578);
or U13282 (N_13282,N_10189,N_9001);
nor U13283 (N_13283,N_11851,N_11004);
and U13284 (N_13284,N_10878,N_9992);
nand U13285 (N_13285,N_10437,N_11811);
nor U13286 (N_13286,N_9526,N_9022);
or U13287 (N_13287,N_11962,N_10080);
and U13288 (N_13288,N_9937,N_10378);
and U13289 (N_13289,N_10452,N_10439);
nand U13290 (N_13290,N_10430,N_9234);
and U13291 (N_13291,N_11151,N_11866);
or U13292 (N_13292,N_9388,N_10738);
nor U13293 (N_13293,N_11006,N_9206);
and U13294 (N_13294,N_11836,N_10844);
and U13295 (N_13295,N_9193,N_11378);
and U13296 (N_13296,N_9249,N_11943);
nor U13297 (N_13297,N_9565,N_10304);
and U13298 (N_13298,N_11657,N_9545);
nor U13299 (N_13299,N_11558,N_10895);
and U13300 (N_13300,N_10770,N_11918);
and U13301 (N_13301,N_9002,N_9479);
or U13302 (N_13302,N_10389,N_9112);
nand U13303 (N_13303,N_11265,N_10008);
or U13304 (N_13304,N_9531,N_10864);
nand U13305 (N_13305,N_11325,N_10640);
or U13306 (N_13306,N_10926,N_11758);
and U13307 (N_13307,N_9576,N_9533);
xor U13308 (N_13308,N_11560,N_10355);
and U13309 (N_13309,N_9409,N_10069);
and U13310 (N_13310,N_9421,N_9851);
and U13311 (N_13311,N_11182,N_10946);
xor U13312 (N_13312,N_9055,N_10902);
and U13313 (N_13313,N_10446,N_9763);
and U13314 (N_13314,N_9485,N_11656);
and U13315 (N_13315,N_10272,N_9218);
or U13316 (N_13316,N_9676,N_11682);
nand U13317 (N_13317,N_9575,N_11563);
and U13318 (N_13318,N_9271,N_11134);
or U13319 (N_13319,N_9336,N_9876);
nand U13320 (N_13320,N_11298,N_10073);
nand U13321 (N_13321,N_11128,N_10054);
xor U13322 (N_13322,N_9413,N_9351);
nor U13323 (N_13323,N_11741,N_10012);
nor U13324 (N_13324,N_11581,N_10559);
nor U13325 (N_13325,N_11208,N_11036);
nand U13326 (N_13326,N_10935,N_11877);
and U13327 (N_13327,N_10601,N_9819);
nor U13328 (N_13328,N_10787,N_9620);
or U13329 (N_13329,N_11756,N_10280);
nor U13330 (N_13330,N_10514,N_9967);
and U13331 (N_13331,N_10205,N_10884);
and U13332 (N_13332,N_10067,N_9279);
nor U13333 (N_13333,N_11928,N_10695);
nor U13334 (N_13334,N_11536,N_10400);
and U13335 (N_13335,N_9675,N_11566);
nor U13336 (N_13336,N_11647,N_10447);
and U13337 (N_13337,N_9969,N_10505);
nand U13338 (N_13338,N_11233,N_10932);
nand U13339 (N_13339,N_9976,N_10915);
nor U13340 (N_13340,N_10747,N_10331);
and U13341 (N_13341,N_11509,N_10511);
and U13342 (N_13342,N_10857,N_9357);
nand U13343 (N_13343,N_9436,N_9303);
or U13344 (N_13344,N_10251,N_10930);
xor U13345 (N_13345,N_10380,N_9008);
nand U13346 (N_13346,N_10494,N_9052);
xnor U13347 (N_13347,N_11272,N_9274);
or U13348 (N_13348,N_9120,N_10186);
nand U13349 (N_13349,N_9844,N_11948);
xor U13350 (N_13350,N_9911,N_11930);
or U13351 (N_13351,N_11270,N_11075);
nand U13352 (N_13352,N_9834,N_9811);
or U13353 (N_13353,N_10841,N_9153);
and U13354 (N_13354,N_9880,N_11416);
nand U13355 (N_13355,N_10207,N_11009);
xnor U13356 (N_13356,N_9325,N_9913);
xnor U13357 (N_13357,N_11037,N_9117);
nand U13358 (N_13358,N_9300,N_10962);
nor U13359 (N_13359,N_11146,N_9370);
nand U13360 (N_13360,N_9815,N_11157);
nor U13361 (N_13361,N_9573,N_11201);
nor U13362 (N_13362,N_9094,N_10487);
or U13363 (N_13363,N_11860,N_9884);
or U13364 (N_13364,N_11803,N_11250);
or U13365 (N_13365,N_10663,N_9671);
xnor U13366 (N_13366,N_11677,N_10050);
nor U13367 (N_13367,N_9012,N_11340);
nor U13368 (N_13368,N_9317,N_10517);
nor U13369 (N_13369,N_11002,N_9310);
xnor U13370 (N_13370,N_9535,N_11732);
nand U13371 (N_13371,N_10217,N_11883);
or U13372 (N_13372,N_10115,N_10166);
and U13373 (N_13373,N_9114,N_9710);
and U13374 (N_13374,N_10938,N_9655);
and U13375 (N_13375,N_10727,N_9612);
nand U13376 (N_13376,N_9367,N_9437);
and U13377 (N_13377,N_11274,N_10755);
nor U13378 (N_13378,N_9041,N_11888);
or U13379 (N_13379,N_10172,N_9440);
and U13380 (N_13380,N_11104,N_9220);
and U13381 (N_13381,N_10093,N_10798);
nor U13382 (N_13382,N_9377,N_11199);
and U13383 (N_13383,N_10648,N_10836);
nand U13384 (N_13384,N_11214,N_10352);
or U13385 (N_13385,N_10697,N_11970);
xor U13386 (N_13386,N_9066,N_11601);
nand U13387 (N_13387,N_10853,N_9773);
or U13388 (N_13388,N_11363,N_9791);
nand U13389 (N_13389,N_11268,N_10531);
and U13390 (N_13390,N_11254,N_9334);
or U13391 (N_13391,N_9476,N_11303);
xor U13392 (N_13392,N_11390,N_10314);
or U13393 (N_13393,N_10733,N_9372);
nand U13394 (N_13394,N_11309,N_11960);
xnor U13395 (N_13395,N_9835,N_10536);
and U13396 (N_13396,N_9885,N_10724);
nor U13397 (N_13397,N_11772,N_11516);
or U13398 (N_13398,N_9038,N_10532);
nand U13399 (N_13399,N_10639,N_11155);
and U13400 (N_13400,N_9313,N_9381);
nor U13401 (N_13401,N_11422,N_9895);
nand U13402 (N_13402,N_9890,N_10390);
and U13403 (N_13403,N_9156,N_11249);
nor U13404 (N_13404,N_10664,N_11083);
xnor U13405 (N_13405,N_9420,N_10775);
nor U13406 (N_13406,N_10968,N_11264);
or U13407 (N_13407,N_11126,N_11259);
and U13408 (N_13408,N_10914,N_11709);
nand U13409 (N_13409,N_10781,N_10824);
nor U13410 (N_13410,N_10039,N_10000);
nand U13411 (N_13411,N_11210,N_9035);
and U13412 (N_13412,N_9500,N_10689);
xnor U13413 (N_13413,N_11680,N_10854);
and U13414 (N_13414,N_10607,N_11774);
nand U13415 (N_13415,N_10076,N_10033);
nand U13416 (N_13416,N_11014,N_9203);
and U13417 (N_13417,N_10241,N_9085);
or U13418 (N_13418,N_9276,N_9986);
and U13419 (N_13419,N_11256,N_10002);
or U13420 (N_13420,N_11913,N_9894);
nor U13421 (N_13421,N_11974,N_9915);
or U13422 (N_13422,N_11747,N_9737);
nor U13423 (N_13423,N_10348,N_10453);
nor U13424 (N_13424,N_11419,N_11933);
or U13425 (N_13425,N_9886,N_9192);
nor U13426 (N_13426,N_9842,N_9662);
nor U13427 (N_13427,N_9290,N_10797);
and U13428 (N_13428,N_9128,N_9419);
and U13429 (N_13429,N_11491,N_10603);
xor U13430 (N_13430,N_9758,N_10710);
nand U13431 (N_13431,N_9987,N_11144);
and U13432 (N_13432,N_9536,N_10575);
nand U13433 (N_13433,N_10325,N_11198);
xnor U13434 (N_13434,N_9006,N_10187);
or U13435 (N_13435,N_9914,N_9771);
or U13436 (N_13436,N_9072,N_10876);
and U13437 (N_13437,N_9616,N_10919);
nand U13438 (N_13438,N_9953,N_9210);
nor U13439 (N_13439,N_10952,N_11235);
nand U13440 (N_13440,N_11480,N_11353);
and U13441 (N_13441,N_9026,N_9121);
and U13442 (N_13442,N_9277,N_10323);
or U13443 (N_13443,N_9195,N_11406);
nand U13444 (N_13444,N_10958,N_9695);
or U13445 (N_13445,N_11394,N_9301);
and U13446 (N_13446,N_11966,N_9944);
nor U13447 (N_13447,N_11886,N_9960);
and U13448 (N_13448,N_10403,N_10563);
or U13449 (N_13449,N_10005,N_9724);
nand U13450 (N_13450,N_11932,N_9608);
and U13451 (N_13451,N_10897,N_11786);
and U13452 (N_13452,N_11726,N_9358);
and U13453 (N_13453,N_10974,N_11739);
nand U13454 (N_13454,N_10341,N_10551);
and U13455 (N_13455,N_10998,N_10394);
and U13456 (N_13456,N_11408,N_10792);
and U13457 (N_13457,N_10778,N_10612);
and U13458 (N_13458,N_10036,N_10621);
and U13459 (N_13459,N_9694,N_9155);
nor U13460 (N_13460,N_11135,N_9049);
nor U13461 (N_13461,N_11981,N_11668);
nor U13462 (N_13462,N_11998,N_10633);
nor U13463 (N_13463,N_11619,N_11232);
and U13464 (N_13464,N_10126,N_11582);
xor U13465 (N_13465,N_10424,N_10491);
nor U13466 (N_13466,N_10880,N_10371);
nor U13467 (N_13467,N_10231,N_11175);
or U13468 (N_13468,N_11956,N_11074);
nand U13469 (N_13469,N_9408,N_9425);
nor U13470 (N_13470,N_9706,N_11022);
nor U13471 (N_13471,N_9748,N_10022);
and U13472 (N_13472,N_10850,N_10561);
or U13473 (N_13473,N_10848,N_9168);
nor U13474 (N_13474,N_9208,N_10363);
xor U13475 (N_13475,N_9779,N_9732);
nand U13476 (N_13476,N_10364,N_10966);
and U13477 (N_13477,N_9800,N_9555);
and U13478 (N_13478,N_9568,N_11701);
or U13479 (N_13479,N_11436,N_10901);
and U13480 (N_13480,N_10644,N_9978);
or U13481 (N_13481,N_10709,N_11992);
or U13482 (N_13482,N_11389,N_11702);
and U13483 (N_13483,N_11444,N_10102);
and U13484 (N_13484,N_11649,N_9629);
nor U13485 (N_13485,N_11672,N_9862);
xor U13486 (N_13486,N_9122,N_9288);
and U13487 (N_13487,N_9898,N_11544);
and U13488 (N_13488,N_11076,N_10171);
nor U13489 (N_13489,N_11223,N_9487);
nand U13490 (N_13490,N_11728,N_9172);
nor U13491 (N_13491,N_10170,N_9194);
nand U13492 (N_13492,N_10222,N_11605);
and U13493 (N_13493,N_10941,N_10286);
and U13494 (N_13494,N_9134,N_10143);
nand U13495 (N_13495,N_11792,N_9806);
nor U13496 (N_13496,N_9727,N_11978);
nand U13497 (N_13497,N_10821,N_10388);
nand U13498 (N_13498,N_10003,N_10742);
xnor U13499 (N_13499,N_10274,N_9648);
and U13500 (N_13500,N_11335,N_11897);
nor U13501 (N_13501,N_11175,N_9553);
or U13502 (N_13502,N_10538,N_9873);
and U13503 (N_13503,N_10423,N_10798);
nor U13504 (N_13504,N_10160,N_11900);
nor U13505 (N_13505,N_10012,N_11677);
and U13506 (N_13506,N_9244,N_9451);
or U13507 (N_13507,N_9413,N_11950);
or U13508 (N_13508,N_11489,N_11855);
nand U13509 (N_13509,N_11032,N_9933);
nor U13510 (N_13510,N_9964,N_10927);
or U13511 (N_13511,N_11053,N_11489);
and U13512 (N_13512,N_11249,N_9346);
xor U13513 (N_13513,N_9595,N_11399);
nor U13514 (N_13514,N_10740,N_9268);
nand U13515 (N_13515,N_11762,N_10132);
and U13516 (N_13516,N_10887,N_10878);
and U13517 (N_13517,N_9974,N_9517);
or U13518 (N_13518,N_11815,N_11540);
or U13519 (N_13519,N_9641,N_11106);
or U13520 (N_13520,N_11744,N_9232);
nor U13521 (N_13521,N_9419,N_10897);
nand U13522 (N_13522,N_10162,N_9466);
nor U13523 (N_13523,N_10454,N_11123);
xor U13524 (N_13524,N_11088,N_9271);
or U13525 (N_13525,N_10754,N_10358);
nor U13526 (N_13526,N_11750,N_9140);
and U13527 (N_13527,N_9763,N_11337);
nand U13528 (N_13528,N_11447,N_11080);
xnor U13529 (N_13529,N_11593,N_10329);
nand U13530 (N_13530,N_9329,N_11694);
nand U13531 (N_13531,N_10112,N_10771);
and U13532 (N_13532,N_10170,N_9693);
nor U13533 (N_13533,N_9842,N_10078);
and U13534 (N_13534,N_11375,N_9845);
or U13535 (N_13535,N_10992,N_11285);
nand U13536 (N_13536,N_11962,N_11309);
or U13537 (N_13537,N_10510,N_9106);
or U13538 (N_13538,N_9598,N_11085);
or U13539 (N_13539,N_11393,N_9234);
or U13540 (N_13540,N_11654,N_11675);
nor U13541 (N_13541,N_9908,N_10109);
and U13542 (N_13542,N_11042,N_11092);
nand U13543 (N_13543,N_11998,N_10535);
xor U13544 (N_13544,N_11724,N_9005);
or U13545 (N_13545,N_9829,N_10337);
nor U13546 (N_13546,N_10974,N_9981);
and U13547 (N_13547,N_9661,N_11283);
xnor U13548 (N_13548,N_10432,N_9492);
or U13549 (N_13549,N_9824,N_11998);
and U13550 (N_13550,N_11052,N_9877);
nor U13551 (N_13551,N_10023,N_9980);
and U13552 (N_13552,N_10234,N_9804);
and U13553 (N_13553,N_11515,N_9653);
or U13554 (N_13554,N_9466,N_10819);
and U13555 (N_13555,N_11711,N_9857);
nor U13556 (N_13556,N_11810,N_11688);
nor U13557 (N_13557,N_10109,N_10381);
nor U13558 (N_13558,N_9911,N_9152);
nor U13559 (N_13559,N_11604,N_9658);
xnor U13560 (N_13560,N_10192,N_9785);
nor U13561 (N_13561,N_10110,N_11751);
nand U13562 (N_13562,N_10445,N_9066);
xnor U13563 (N_13563,N_11772,N_11770);
nor U13564 (N_13564,N_10391,N_9781);
nor U13565 (N_13565,N_11608,N_10068);
nor U13566 (N_13566,N_9467,N_9217);
nor U13567 (N_13567,N_11577,N_10465);
and U13568 (N_13568,N_11280,N_9477);
nand U13569 (N_13569,N_9915,N_11106);
and U13570 (N_13570,N_10563,N_9951);
or U13571 (N_13571,N_9903,N_11788);
or U13572 (N_13572,N_9975,N_10640);
nor U13573 (N_13573,N_10608,N_9160);
or U13574 (N_13574,N_10557,N_11069);
nor U13575 (N_13575,N_10073,N_11742);
or U13576 (N_13576,N_9353,N_10890);
nand U13577 (N_13577,N_11643,N_11586);
nand U13578 (N_13578,N_9861,N_9478);
or U13579 (N_13579,N_11850,N_9085);
and U13580 (N_13580,N_10954,N_11218);
nand U13581 (N_13581,N_11179,N_10440);
and U13582 (N_13582,N_10508,N_10769);
xor U13583 (N_13583,N_10374,N_11695);
nor U13584 (N_13584,N_11915,N_9929);
and U13585 (N_13585,N_9089,N_10045);
and U13586 (N_13586,N_11246,N_9443);
nand U13587 (N_13587,N_10797,N_10045);
xor U13588 (N_13588,N_9651,N_11811);
and U13589 (N_13589,N_11417,N_9158);
or U13590 (N_13590,N_9928,N_9553);
or U13591 (N_13591,N_11013,N_11702);
xnor U13592 (N_13592,N_9461,N_10281);
and U13593 (N_13593,N_11126,N_11082);
or U13594 (N_13594,N_10123,N_10059);
nor U13595 (N_13595,N_10177,N_10960);
nor U13596 (N_13596,N_11290,N_10772);
nor U13597 (N_13597,N_11306,N_10538);
nor U13598 (N_13598,N_11211,N_9994);
nor U13599 (N_13599,N_10758,N_11100);
nor U13600 (N_13600,N_10243,N_11756);
nand U13601 (N_13601,N_11932,N_11825);
or U13602 (N_13602,N_9033,N_10114);
nand U13603 (N_13603,N_11714,N_10909);
nand U13604 (N_13604,N_10720,N_9957);
xor U13605 (N_13605,N_10337,N_10972);
or U13606 (N_13606,N_10570,N_10080);
nor U13607 (N_13607,N_10959,N_9999);
nor U13608 (N_13608,N_9983,N_10560);
nor U13609 (N_13609,N_9076,N_10671);
nand U13610 (N_13610,N_9937,N_10014);
and U13611 (N_13611,N_10521,N_11960);
or U13612 (N_13612,N_9926,N_9028);
nor U13613 (N_13613,N_9652,N_10211);
nand U13614 (N_13614,N_9966,N_9862);
or U13615 (N_13615,N_10196,N_11510);
and U13616 (N_13616,N_9072,N_11880);
or U13617 (N_13617,N_9110,N_9411);
and U13618 (N_13618,N_10046,N_9556);
nand U13619 (N_13619,N_11925,N_10586);
and U13620 (N_13620,N_11884,N_11532);
or U13621 (N_13621,N_9820,N_9969);
or U13622 (N_13622,N_11632,N_10512);
xor U13623 (N_13623,N_9799,N_10252);
and U13624 (N_13624,N_11996,N_10802);
nor U13625 (N_13625,N_11024,N_9752);
or U13626 (N_13626,N_11025,N_10485);
nor U13627 (N_13627,N_10897,N_10857);
or U13628 (N_13628,N_11952,N_9329);
and U13629 (N_13629,N_10976,N_10412);
and U13630 (N_13630,N_10566,N_10220);
or U13631 (N_13631,N_10530,N_10544);
nand U13632 (N_13632,N_10847,N_10824);
nand U13633 (N_13633,N_10835,N_9125);
nand U13634 (N_13634,N_10486,N_11111);
nand U13635 (N_13635,N_9102,N_11632);
or U13636 (N_13636,N_10520,N_11583);
nor U13637 (N_13637,N_11426,N_10124);
nor U13638 (N_13638,N_11262,N_10233);
nor U13639 (N_13639,N_10561,N_10248);
and U13640 (N_13640,N_9929,N_10134);
and U13641 (N_13641,N_11625,N_11343);
nand U13642 (N_13642,N_11753,N_11170);
and U13643 (N_13643,N_11673,N_9223);
xnor U13644 (N_13644,N_9111,N_11774);
nand U13645 (N_13645,N_9988,N_11229);
xnor U13646 (N_13646,N_10241,N_9690);
or U13647 (N_13647,N_10209,N_11242);
nand U13648 (N_13648,N_11970,N_11170);
and U13649 (N_13649,N_9365,N_9765);
nand U13650 (N_13650,N_9662,N_11736);
or U13651 (N_13651,N_11918,N_11431);
or U13652 (N_13652,N_10514,N_11192);
or U13653 (N_13653,N_9227,N_9589);
nor U13654 (N_13654,N_11713,N_11901);
nand U13655 (N_13655,N_10617,N_9255);
nor U13656 (N_13656,N_10710,N_9446);
and U13657 (N_13657,N_11222,N_9337);
nand U13658 (N_13658,N_11868,N_11834);
and U13659 (N_13659,N_11335,N_11832);
and U13660 (N_13660,N_11557,N_9222);
nor U13661 (N_13661,N_10331,N_9754);
and U13662 (N_13662,N_9201,N_9861);
or U13663 (N_13663,N_9055,N_11099);
nand U13664 (N_13664,N_11579,N_10358);
nand U13665 (N_13665,N_10086,N_11515);
and U13666 (N_13666,N_11677,N_10292);
or U13667 (N_13667,N_9323,N_11837);
nor U13668 (N_13668,N_9821,N_11832);
or U13669 (N_13669,N_11930,N_9620);
nor U13670 (N_13670,N_9775,N_10629);
and U13671 (N_13671,N_10484,N_11377);
nand U13672 (N_13672,N_11709,N_11267);
nor U13673 (N_13673,N_9363,N_11432);
nor U13674 (N_13674,N_11892,N_9926);
xor U13675 (N_13675,N_9681,N_10219);
nor U13676 (N_13676,N_11799,N_9203);
nor U13677 (N_13677,N_10963,N_9355);
nand U13678 (N_13678,N_11301,N_11960);
and U13679 (N_13679,N_9380,N_11879);
or U13680 (N_13680,N_9986,N_11996);
or U13681 (N_13681,N_9815,N_11653);
nand U13682 (N_13682,N_10579,N_10444);
nor U13683 (N_13683,N_11024,N_11073);
and U13684 (N_13684,N_10791,N_10971);
nor U13685 (N_13685,N_10657,N_10644);
or U13686 (N_13686,N_10373,N_9344);
nand U13687 (N_13687,N_9123,N_9570);
and U13688 (N_13688,N_11565,N_9146);
xnor U13689 (N_13689,N_9069,N_10995);
xnor U13690 (N_13690,N_10752,N_11737);
nor U13691 (N_13691,N_9900,N_9210);
or U13692 (N_13692,N_10517,N_10080);
and U13693 (N_13693,N_11853,N_11345);
nor U13694 (N_13694,N_10525,N_9380);
xnor U13695 (N_13695,N_11849,N_11632);
and U13696 (N_13696,N_10211,N_9932);
and U13697 (N_13697,N_10073,N_9764);
nand U13698 (N_13698,N_9334,N_10001);
and U13699 (N_13699,N_11887,N_11925);
nand U13700 (N_13700,N_9667,N_9604);
nor U13701 (N_13701,N_10053,N_10637);
nor U13702 (N_13702,N_10278,N_10486);
nand U13703 (N_13703,N_9232,N_11091);
nand U13704 (N_13704,N_10368,N_11959);
nor U13705 (N_13705,N_11566,N_9695);
or U13706 (N_13706,N_10656,N_9306);
nand U13707 (N_13707,N_10350,N_11526);
nand U13708 (N_13708,N_9763,N_9882);
or U13709 (N_13709,N_11851,N_11681);
nor U13710 (N_13710,N_9910,N_10332);
nor U13711 (N_13711,N_11077,N_11491);
or U13712 (N_13712,N_9982,N_10319);
nand U13713 (N_13713,N_9990,N_9591);
nand U13714 (N_13714,N_9359,N_11693);
nor U13715 (N_13715,N_11107,N_11207);
and U13716 (N_13716,N_9574,N_11828);
and U13717 (N_13717,N_10346,N_11897);
or U13718 (N_13718,N_10438,N_10435);
or U13719 (N_13719,N_11572,N_9838);
nand U13720 (N_13720,N_9162,N_11108);
or U13721 (N_13721,N_11583,N_11349);
nor U13722 (N_13722,N_10832,N_9376);
and U13723 (N_13723,N_10720,N_9434);
or U13724 (N_13724,N_11126,N_11363);
and U13725 (N_13725,N_10184,N_11083);
or U13726 (N_13726,N_10799,N_10096);
nor U13727 (N_13727,N_11870,N_10684);
nor U13728 (N_13728,N_11572,N_10603);
nand U13729 (N_13729,N_11098,N_10011);
nor U13730 (N_13730,N_11498,N_9162);
and U13731 (N_13731,N_10239,N_10388);
or U13732 (N_13732,N_11555,N_11214);
or U13733 (N_13733,N_10372,N_11221);
and U13734 (N_13734,N_9069,N_9806);
and U13735 (N_13735,N_11461,N_9592);
nor U13736 (N_13736,N_10706,N_10301);
nand U13737 (N_13737,N_11995,N_9467);
and U13738 (N_13738,N_9046,N_9988);
or U13739 (N_13739,N_9980,N_9011);
nand U13740 (N_13740,N_11915,N_11979);
nand U13741 (N_13741,N_11804,N_9315);
nor U13742 (N_13742,N_9512,N_10646);
and U13743 (N_13743,N_11696,N_9722);
nor U13744 (N_13744,N_10838,N_11014);
xor U13745 (N_13745,N_11896,N_11159);
or U13746 (N_13746,N_9631,N_10722);
and U13747 (N_13747,N_9463,N_11313);
and U13748 (N_13748,N_9209,N_10995);
or U13749 (N_13749,N_10577,N_11218);
and U13750 (N_13750,N_10129,N_11095);
nor U13751 (N_13751,N_9180,N_9020);
or U13752 (N_13752,N_9939,N_10248);
or U13753 (N_13753,N_10478,N_9755);
or U13754 (N_13754,N_11951,N_10697);
nand U13755 (N_13755,N_10541,N_9439);
and U13756 (N_13756,N_9659,N_9064);
or U13757 (N_13757,N_10555,N_9320);
and U13758 (N_13758,N_10383,N_10690);
nand U13759 (N_13759,N_9778,N_9999);
and U13760 (N_13760,N_9265,N_10429);
nor U13761 (N_13761,N_10606,N_11644);
nand U13762 (N_13762,N_10983,N_10212);
and U13763 (N_13763,N_9713,N_9023);
nor U13764 (N_13764,N_11319,N_10308);
or U13765 (N_13765,N_10883,N_10369);
nor U13766 (N_13766,N_10122,N_11992);
nor U13767 (N_13767,N_9149,N_10055);
nor U13768 (N_13768,N_10552,N_11128);
and U13769 (N_13769,N_11401,N_10131);
nor U13770 (N_13770,N_10282,N_9998);
xnor U13771 (N_13771,N_11699,N_9340);
and U13772 (N_13772,N_10934,N_9819);
nand U13773 (N_13773,N_9165,N_10921);
and U13774 (N_13774,N_10524,N_11818);
nor U13775 (N_13775,N_10403,N_9168);
or U13776 (N_13776,N_10769,N_10926);
and U13777 (N_13777,N_10858,N_11567);
or U13778 (N_13778,N_10063,N_9970);
nor U13779 (N_13779,N_11178,N_11187);
or U13780 (N_13780,N_10922,N_10151);
and U13781 (N_13781,N_10396,N_10074);
xnor U13782 (N_13782,N_10830,N_10517);
and U13783 (N_13783,N_9387,N_11883);
nor U13784 (N_13784,N_9187,N_11490);
nor U13785 (N_13785,N_11680,N_11327);
nand U13786 (N_13786,N_10782,N_9532);
and U13787 (N_13787,N_9432,N_9179);
nor U13788 (N_13788,N_10398,N_9476);
or U13789 (N_13789,N_9900,N_11950);
nor U13790 (N_13790,N_11845,N_9432);
and U13791 (N_13791,N_10255,N_11135);
and U13792 (N_13792,N_10208,N_9900);
or U13793 (N_13793,N_11576,N_9327);
and U13794 (N_13794,N_11668,N_10269);
or U13795 (N_13795,N_11849,N_11794);
nor U13796 (N_13796,N_11604,N_11327);
and U13797 (N_13797,N_9301,N_9191);
nor U13798 (N_13798,N_9488,N_11282);
and U13799 (N_13799,N_10007,N_11303);
nand U13800 (N_13800,N_9842,N_10662);
nand U13801 (N_13801,N_11066,N_11002);
and U13802 (N_13802,N_11860,N_11562);
nor U13803 (N_13803,N_9458,N_10259);
nand U13804 (N_13804,N_9032,N_11739);
and U13805 (N_13805,N_11288,N_11765);
nand U13806 (N_13806,N_9955,N_11921);
nor U13807 (N_13807,N_9196,N_9235);
xor U13808 (N_13808,N_10501,N_11345);
nand U13809 (N_13809,N_11745,N_10645);
nor U13810 (N_13810,N_11647,N_9267);
nand U13811 (N_13811,N_11891,N_11062);
xnor U13812 (N_13812,N_9810,N_11430);
nand U13813 (N_13813,N_9586,N_9976);
or U13814 (N_13814,N_11618,N_10560);
or U13815 (N_13815,N_10108,N_9623);
nor U13816 (N_13816,N_10298,N_10461);
and U13817 (N_13817,N_11558,N_9634);
nand U13818 (N_13818,N_10312,N_9540);
nand U13819 (N_13819,N_10584,N_11614);
xor U13820 (N_13820,N_9846,N_9718);
or U13821 (N_13821,N_9850,N_11487);
and U13822 (N_13822,N_11701,N_9079);
and U13823 (N_13823,N_9273,N_11789);
nor U13824 (N_13824,N_10987,N_10834);
nand U13825 (N_13825,N_11792,N_11531);
nand U13826 (N_13826,N_9050,N_10305);
and U13827 (N_13827,N_9119,N_9680);
nor U13828 (N_13828,N_11855,N_10514);
nand U13829 (N_13829,N_9188,N_11847);
or U13830 (N_13830,N_10983,N_11587);
nand U13831 (N_13831,N_11816,N_11691);
and U13832 (N_13832,N_9369,N_10507);
nor U13833 (N_13833,N_11687,N_11216);
nand U13834 (N_13834,N_9065,N_10038);
and U13835 (N_13835,N_10837,N_11898);
nor U13836 (N_13836,N_9781,N_10765);
nor U13837 (N_13837,N_10158,N_10609);
or U13838 (N_13838,N_9369,N_11610);
nor U13839 (N_13839,N_9058,N_11887);
and U13840 (N_13840,N_10218,N_9414);
nor U13841 (N_13841,N_10928,N_10019);
nor U13842 (N_13842,N_11922,N_11984);
nor U13843 (N_13843,N_10220,N_10514);
and U13844 (N_13844,N_9225,N_10108);
nand U13845 (N_13845,N_9536,N_11364);
nor U13846 (N_13846,N_11541,N_11407);
xnor U13847 (N_13847,N_9267,N_10336);
and U13848 (N_13848,N_9929,N_9623);
or U13849 (N_13849,N_10799,N_9628);
nor U13850 (N_13850,N_9838,N_11481);
nor U13851 (N_13851,N_10105,N_11564);
and U13852 (N_13852,N_11936,N_10348);
nand U13853 (N_13853,N_11701,N_9773);
nor U13854 (N_13854,N_9540,N_11380);
or U13855 (N_13855,N_9895,N_10905);
nor U13856 (N_13856,N_9165,N_11040);
or U13857 (N_13857,N_10541,N_9195);
or U13858 (N_13858,N_11579,N_9966);
nor U13859 (N_13859,N_11749,N_9308);
nand U13860 (N_13860,N_10296,N_11396);
or U13861 (N_13861,N_9388,N_9114);
or U13862 (N_13862,N_9428,N_9312);
nand U13863 (N_13863,N_11339,N_9722);
nor U13864 (N_13864,N_9492,N_11068);
nor U13865 (N_13865,N_11091,N_10103);
nand U13866 (N_13866,N_11111,N_11092);
nor U13867 (N_13867,N_11615,N_11668);
nand U13868 (N_13868,N_9997,N_9785);
and U13869 (N_13869,N_9717,N_10323);
xnor U13870 (N_13870,N_10255,N_9972);
and U13871 (N_13871,N_10771,N_10821);
and U13872 (N_13872,N_9083,N_10320);
and U13873 (N_13873,N_10292,N_9077);
nor U13874 (N_13874,N_9976,N_11272);
nand U13875 (N_13875,N_9352,N_9162);
nand U13876 (N_13876,N_11911,N_11882);
nand U13877 (N_13877,N_11684,N_10190);
or U13878 (N_13878,N_10963,N_10728);
nor U13879 (N_13879,N_10368,N_11130);
or U13880 (N_13880,N_9254,N_9884);
or U13881 (N_13881,N_9540,N_9428);
nand U13882 (N_13882,N_11899,N_9736);
or U13883 (N_13883,N_11205,N_11884);
and U13884 (N_13884,N_10717,N_10955);
nor U13885 (N_13885,N_10674,N_11153);
nor U13886 (N_13886,N_11754,N_9995);
or U13887 (N_13887,N_10729,N_10178);
nor U13888 (N_13888,N_9104,N_11113);
xnor U13889 (N_13889,N_11128,N_11856);
and U13890 (N_13890,N_11371,N_9659);
nor U13891 (N_13891,N_9097,N_11572);
xnor U13892 (N_13892,N_10354,N_9188);
nor U13893 (N_13893,N_9944,N_11990);
xor U13894 (N_13894,N_10932,N_11856);
nor U13895 (N_13895,N_9290,N_10876);
and U13896 (N_13896,N_11336,N_10695);
nor U13897 (N_13897,N_10287,N_11652);
nand U13898 (N_13898,N_11616,N_10194);
xnor U13899 (N_13899,N_9210,N_9734);
nand U13900 (N_13900,N_11947,N_11513);
and U13901 (N_13901,N_10124,N_11085);
or U13902 (N_13902,N_10573,N_11272);
and U13903 (N_13903,N_11666,N_10968);
nand U13904 (N_13904,N_10520,N_11598);
and U13905 (N_13905,N_10568,N_10559);
nor U13906 (N_13906,N_9185,N_11933);
nand U13907 (N_13907,N_11647,N_10115);
or U13908 (N_13908,N_11866,N_11685);
nand U13909 (N_13909,N_10674,N_11108);
nand U13910 (N_13910,N_11793,N_10221);
nor U13911 (N_13911,N_9758,N_9383);
and U13912 (N_13912,N_9279,N_11366);
xnor U13913 (N_13913,N_10749,N_11986);
nor U13914 (N_13914,N_9526,N_10711);
and U13915 (N_13915,N_9502,N_11286);
or U13916 (N_13916,N_11079,N_9681);
or U13917 (N_13917,N_11497,N_9640);
nor U13918 (N_13918,N_10716,N_10811);
nor U13919 (N_13919,N_10539,N_11323);
nor U13920 (N_13920,N_11487,N_10143);
or U13921 (N_13921,N_10183,N_9213);
nor U13922 (N_13922,N_11614,N_11899);
nor U13923 (N_13923,N_11415,N_9718);
nand U13924 (N_13924,N_9982,N_9378);
or U13925 (N_13925,N_9267,N_11564);
nand U13926 (N_13926,N_11017,N_10302);
nor U13927 (N_13927,N_9013,N_9849);
and U13928 (N_13928,N_11671,N_9929);
nand U13929 (N_13929,N_11342,N_10528);
nor U13930 (N_13930,N_9468,N_10256);
nor U13931 (N_13931,N_10516,N_9645);
nand U13932 (N_13932,N_10932,N_9117);
nor U13933 (N_13933,N_11392,N_10861);
or U13934 (N_13934,N_10222,N_10219);
or U13935 (N_13935,N_9054,N_11880);
and U13936 (N_13936,N_9364,N_10318);
and U13937 (N_13937,N_11396,N_11323);
nor U13938 (N_13938,N_11215,N_10420);
or U13939 (N_13939,N_10988,N_11316);
or U13940 (N_13940,N_11476,N_9607);
or U13941 (N_13941,N_10471,N_9475);
nor U13942 (N_13942,N_10608,N_11249);
nand U13943 (N_13943,N_9907,N_10639);
or U13944 (N_13944,N_11794,N_10871);
and U13945 (N_13945,N_9937,N_9466);
or U13946 (N_13946,N_10713,N_10028);
and U13947 (N_13947,N_9038,N_9511);
or U13948 (N_13948,N_11853,N_9446);
nand U13949 (N_13949,N_10042,N_11405);
xnor U13950 (N_13950,N_11418,N_9412);
xor U13951 (N_13951,N_11977,N_9942);
nand U13952 (N_13952,N_9519,N_9091);
and U13953 (N_13953,N_9698,N_10687);
or U13954 (N_13954,N_9528,N_9132);
or U13955 (N_13955,N_11686,N_10392);
or U13956 (N_13956,N_11896,N_10283);
nor U13957 (N_13957,N_10840,N_10889);
or U13958 (N_13958,N_9972,N_9824);
and U13959 (N_13959,N_11296,N_11856);
nand U13960 (N_13960,N_11316,N_10382);
nand U13961 (N_13961,N_9271,N_9029);
nor U13962 (N_13962,N_9991,N_9048);
or U13963 (N_13963,N_11884,N_9133);
and U13964 (N_13964,N_10785,N_10572);
nor U13965 (N_13965,N_10609,N_10233);
and U13966 (N_13966,N_9210,N_9758);
nor U13967 (N_13967,N_10449,N_9758);
and U13968 (N_13968,N_10199,N_9884);
nor U13969 (N_13969,N_9916,N_11310);
nand U13970 (N_13970,N_9135,N_10619);
and U13971 (N_13971,N_10799,N_11614);
nand U13972 (N_13972,N_11665,N_10802);
nor U13973 (N_13973,N_9696,N_11361);
or U13974 (N_13974,N_11018,N_9104);
nor U13975 (N_13975,N_11146,N_11990);
nor U13976 (N_13976,N_11596,N_9570);
nor U13977 (N_13977,N_10476,N_11484);
and U13978 (N_13978,N_11095,N_10519);
and U13979 (N_13979,N_10503,N_10548);
nor U13980 (N_13980,N_10560,N_9352);
nand U13981 (N_13981,N_9336,N_11459);
or U13982 (N_13982,N_10077,N_10939);
nand U13983 (N_13983,N_9296,N_11384);
nand U13984 (N_13984,N_11004,N_9531);
and U13985 (N_13985,N_11573,N_10143);
xnor U13986 (N_13986,N_9769,N_11399);
and U13987 (N_13987,N_11238,N_9469);
nor U13988 (N_13988,N_10880,N_10716);
nand U13989 (N_13989,N_11552,N_11193);
nand U13990 (N_13990,N_10434,N_10752);
nand U13991 (N_13991,N_10179,N_9777);
nand U13992 (N_13992,N_10298,N_9352);
or U13993 (N_13993,N_10230,N_10404);
nand U13994 (N_13994,N_10578,N_11661);
and U13995 (N_13995,N_9224,N_11784);
and U13996 (N_13996,N_11110,N_10141);
and U13997 (N_13997,N_9588,N_11554);
nor U13998 (N_13998,N_11666,N_9969);
xnor U13999 (N_13999,N_10728,N_9672);
and U14000 (N_14000,N_9247,N_11499);
or U14001 (N_14001,N_9240,N_11051);
or U14002 (N_14002,N_9065,N_9944);
xnor U14003 (N_14003,N_9246,N_10181);
and U14004 (N_14004,N_9269,N_10215);
or U14005 (N_14005,N_11267,N_9347);
nand U14006 (N_14006,N_11735,N_9300);
xnor U14007 (N_14007,N_11679,N_10645);
or U14008 (N_14008,N_11299,N_10837);
and U14009 (N_14009,N_10645,N_11790);
or U14010 (N_14010,N_9698,N_11107);
or U14011 (N_14011,N_9216,N_10141);
or U14012 (N_14012,N_10651,N_9012);
or U14013 (N_14013,N_9127,N_10564);
nor U14014 (N_14014,N_10325,N_9560);
xnor U14015 (N_14015,N_10359,N_11918);
xnor U14016 (N_14016,N_11262,N_11593);
or U14017 (N_14017,N_10219,N_9434);
or U14018 (N_14018,N_10947,N_10472);
or U14019 (N_14019,N_11172,N_11704);
and U14020 (N_14020,N_9350,N_9926);
or U14021 (N_14021,N_11704,N_11365);
nand U14022 (N_14022,N_9923,N_9757);
nor U14023 (N_14023,N_9194,N_9024);
or U14024 (N_14024,N_9921,N_9971);
and U14025 (N_14025,N_11217,N_9145);
nor U14026 (N_14026,N_10082,N_10504);
xor U14027 (N_14027,N_10645,N_9645);
nor U14028 (N_14028,N_10990,N_9274);
or U14029 (N_14029,N_9215,N_9110);
xor U14030 (N_14030,N_11614,N_11759);
or U14031 (N_14031,N_10855,N_9216);
nand U14032 (N_14032,N_9784,N_10301);
nor U14033 (N_14033,N_10484,N_10566);
nand U14034 (N_14034,N_10592,N_9562);
xor U14035 (N_14035,N_10234,N_11508);
xor U14036 (N_14036,N_9998,N_9520);
nand U14037 (N_14037,N_9876,N_10562);
xor U14038 (N_14038,N_10382,N_9965);
or U14039 (N_14039,N_10214,N_9547);
and U14040 (N_14040,N_11339,N_11863);
and U14041 (N_14041,N_11941,N_9275);
nand U14042 (N_14042,N_9893,N_10344);
and U14043 (N_14043,N_11176,N_9677);
and U14044 (N_14044,N_11813,N_11385);
xor U14045 (N_14045,N_11598,N_11734);
and U14046 (N_14046,N_9328,N_9926);
and U14047 (N_14047,N_10427,N_9769);
and U14048 (N_14048,N_10479,N_10687);
nand U14049 (N_14049,N_9760,N_9087);
nand U14050 (N_14050,N_10653,N_9268);
nor U14051 (N_14051,N_9997,N_11652);
nor U14052 (N_14052,N_11652,N_9286);
xnor U14053 (N_14053,N_10989,N_10994);
nand U14054 (N_14054,N_9185,N_9896);
and U14055 (N_14055,N_11296,N_10571);
nand U14056 (N_14056,N_9120,N_11513);
nand U14057 (N_14057,N_11316,N_11393);
nand U14058 (N_14058,N_9233,N_11361);
nor U14059 (N_14059,N_9492,N_9868);
or U14060 (N_14060,N_11752,N_9524);
xnor U14061 (N_14061,N_11871,N_9065);
nand U14062 (N_14062,N_9248,N_11821);
nor U14063 (N_14063,N_11550,N_11866);
nand U14064 (N_14064,N_9502,N_11593);
or U14065 (N_14065,N_10687,N_10008);
nand U14066 (N_14066,N_11559,N_10323);
or U14067 (N_14067,N_9707,N_11068);
nor U14068 (N_14068,N_9521,N_10358);
or U14069 (N_14069,N_9136,N_10133);
xor U14070 (N_14070,N_10086,N_11201);
nor U14071 (N_14071,N_11073,N_10700);
or U14072 (N_14072,N_9152,N_10822);
nor U14073 (N_14073,N_9813,N_11308);
or U14074 (N_14074,N_9190,N_11507);
nor U14075 (N_14075,N_11307,N_9663);
nand U14076 (N_14076,N_10564,N_9749);
nand U14077 (N_14077,N_11310,N_11458);
nor U14078 (N_14078,N_10382,N_11577);
and U14079 (N_14079,N_10171,N_10953);
or U14080 (N_14080,N_10966,N_9779);
or U14081 (N_14081,N_10507,N_9406);
or U14082 (N_14082,N_9959,N_11029);
nor U14083 (N_14083,N_11157,N_9684);
nor U14084 (N_14084,N_11922,N_10862);
or U14085 (N_14085,N_10502,N_11379);
or U14086 (N_14086,N_9641,N_10847);
xnor U14087 (N_14087,N_10898,N_11208);
nor U14088 (N_14088,N_11776,N_9175);
nand U14089 (N_14089,N_9058,N_9670);
nand U14090 (N_14090,N_11048,N_10461);
nor U14091 (N_14091,N_11911,N_10913);
nor U14092 (N_14092,N_11041,N_9741);
nor U14093 (N_14093,N_9208,N_9411);
and U14094 (N_14094,N_10626,N_9685);
and U14095 (N_14095,N_11091,N_9196);
or U14096 (N_14096,N_10142,N_9431);
xor U14097 (N_14097,N_9532,N_10177);
xnor U14098 (N_14098,N_9822,N_9554);
nand U14099 (N_14099,N_10298,N_11182);
nand U14100 (N_14100,N_9145,N_10822);
nor U14101 (N_14101,N_9860,N_9142);
nor U14102 (N_14102,N_10819,N_9974);
nand U14103 (N_14103,N_11936,N_11778);
nor U14104 (N_14104,N_11255,N_11354);
nand U14105 (N_14105,N_9166,N_9700);
nand U14106 (N_14106,N_10872,N_10955);
nor U14107 (N_14107,N_9554,N_11097);
nor U14108 (N_14108,N_10084,N_10030);
and U14109 (N_14109,N_10223,N_10598);
nand U14110 (N_14110,N_9623,N_10965);
nor U14111 (N_14111,N_9259,N_10031);
nor U14112 (N_14112,N_11865,N_10841);
nand U14113 (N_14113,N_10663,N_11691);
and U14114 (N_14114,N_9828,N_10386);
and U14115 (N_14115,N_9912,N_11953);
or U14116 (N_14116,N_10499,N_10259);
nand U14117 (N_14117,N_11733,N_9636);
xnor U14118 (N_14118,N_9316,N_10775);
or U14119 (N_14119,N_9109,N_10844);
and U14120 (N_14120,N_9405,N_9064);
nand U14121 (N_14121,N_11705,N_9512);
xor U14122 (N_14122,N_11210,N_9893);
nor U14123 (N_14123,N_10019,N_11056);
and U14124 (N_14124,N_10393,N_11958);
or U14125 (N_14125,N_11948,N_11683);
or U14126 (N_14126,N_9366,N_9117);
or U14127 (N_14127,N_10521,N_9801);
nor U14128 (N_14128,N_9902,N_11855);
nand U14129 (N_14129,N_11943,N_11424);
or U14130 (N_14130,N_9305,N_11727);
and U14131 (N_14131,N_11332,N_9054);
or U14132 (N_14132,N_9480,N_10422);
nand U14133 (N_14133,N_10902,N_11062);
nor U14134 (N_14134,N_11207,N_11434);
or U14135 (N_14135,N_9358,N_11884);
nor U14136 (N_14136,N_10571,N_10202);
and U14137 (N_14137,N_11002,N_11777);
nor U14138 (N_14138,N_10988,N_9911);
nand U14139 (N_14139,N_11049,N_11464);
nand U14140 (N_14140,N_11691,N_9402);
nand U14141 (N_14141,N_10947,N_11154);
nand U14142 (N_14142,N_10485,N_9857);
nand U14143 (N_14143,N_11856,N_11481);
and U14144 (N_14144,N_9694,N_11205);
xnor U14145 (N_14145,N_10188,N_9408);
and U14146 (N_14146,N_9258,N_9319);
or U14147 (N_14147,N_10496,N_11923);
nand U14148 (N_14148,N_10327,N_10471);
and U14149 (N_14149,N_9072,N_9532);
nor U14150 (N_14150,N_9569,N_10639);
nand U14151 (N_14151,N_9388,N_10928);
nor U14152 (N_14152,N_9376,N_9091);
nand U14153 (N_14153,N_10540,N_10018);
nand U14154 (N_14154,N_11060,N_9714);
and U14155 (N_14155,N_10573,N_10133);
or U14156 (N_14156,N_10521,N_11392);
xor U14157 (N_14157,N_10543,N_9757);
xnor U14158 (N_14158,N_9598,N_11672);
and U14159 (N_14159,N_9952,N_9177);
xor U14160 (N_14160,N_10908,N_10171);
or U14161 (N_14161,N_10911,N_10920);
nand U14162 (N_14162,N_9925,N_10430);
nor U14163 (N_14163,N_11675,N_9828);
nor U14164 (N_14164,N_9243,N_9383);
and U14165 (N_14165,N_10200,N_11745);
nand U14166 (N_14166,N_11356,N_11897);
xnor U14167 (N_14167,N_9383,N_10704);
nand U14168 (N_14168,N_11646,N_9341);
or U14169 (N_14169,N_10305,N_11782);
and U14170 (N_14170,N_9373,N_9269);
and U14171 (N_14171,N_9858,N_10715);
nor U14172 (N_14172,N_11085,N_11241);
and U14173 (N_14173,N_11882,N_9839);
and U14174 (N_14174,N_9344,N_10241);
or U14175 (N_14175,N_10857,N_10012);
or U14176 (N_14176,N_9097,N_11446);
nand U14177 (N_14177,N_9323,N_11905);
nand U14178 (N_14178,N_11408,N_9586);
or U14179 (N_14179,N_9554,N_11524);
nor U14180 (N_14180,N_11970,N_9589);
nor U14181 (N_14181,N_9437,N_9738);
and U14182 (N_14182,N_10966,N_10406);
or U14183 (N_14183,N_9628,N_10761);
and U14184 (N_14184,N_10967,N_9739);
nand U14185 (N_14185,N_10723,N_9678);
nor U14186 (N_14186,N_9115,N_9029);
nor U14187 (N_14187,N_11729,N_10491);
nor U14188 (N_14188,N_11461,N_11376);
nor U14189 (N_14189,N_11503,N_9014);
nor U14190 (N_14190,N_10774,N_10918);
nand U14191 (N_14191,N_9553,N_11745);
or U14192 (N_14192,N_10293,N_11245);
nor U14193 (N_14193,N_11967,N_11649);
xnor U14194 (N_14194,N_9473,N_11658);
or U14195 (N_14195,N_9517,N_11740);
and U14196 (N_14196,N_10129,N_10355);
nand U14197 (N_14197,N_11558,N_11054);
or U14198 (N_14198,N_11994,N_9057);
or U14199 (N_14199,N_11742,N_10612);
nand U14200 (N_14200,N_10304,N_10860);
nand U14201 (N_14201,N_10414,N_9757);
xor U14202 (N_14202,N_9344,N_11095);
or U14203 (N_14203,N_11247,N_9304);
or U14204 (N_14204,N_10275,N_10716);
nor U14205 (N_14205,N_10170,N_10056);
nand U14206 (N_14206,N_10827,N_10130);
or U14207 (N_14207,N_9977,N_9275);
nor U14208 (N_14208,N_10174,N_10615);
nor U14209 (N_14209,N_9662,N_11358);
nand U14210 (N_14210,N_11191,N_9080);
or U14211 (N_14211,N_11813,N_9446);
or U14212 (N_14212,N_11350,N_9395);
xor U14213 (N_14213,N_10654,N_9969);
xor U14214 (N_14214,N_10615,N_9054);
nor U14215 (N_14215,N_11634,N_9004);
nor U14216 (N_14216,N_9646,N_9292);
and U14217 (N_14217,N_9533,N_11448);
xor U14218 (N_14218,N_9039,N_10390);
nand U14219 (N_14219,N_9726,N_10110);
and U14220 (N_14220,N_9469,N_10107);
and U14221 (N_14221,N_11246,N_10347);
nor U14222 (N_14222,N_10502,N_11239);
or U14223 (N_14223,N_11921,N_9254);
and U14224 (N_14224,N_11074,N_9115);
nand U14225 (N_14225,N_10097,N_11201);
nor U14226 (N_14226,N_11290,N_9303);
and U14227 (N_14227,N_10144,N_10659);
or U14228 (N_14228,N_11888,N_11592);
xor U14229 (N_14229,N_11987,N_11689);
and U14230 (N_14230,N_11848,N_11406);
nand U14231 (N_14231,N_10205,N_9274);
or U14232 (N_14232,N_9525,N_11910);
nor U14233 (N_14233,N_10704,N_9725);
and U14234 (N_14234,N_11505,N_9132);
and U14235 (N_14235,N_11675,N_11553);
or U14236 (N_14236,N_11593,N_11110);
and U14237 (N_14237,N_10379,N_10319);
nand U14238 (N_14238,N_10099,N_11514);
and U14239 (N_14239,N_11309,N_11570);
nor U14240 (N_14240,N_11590,N_9854);
nor U14241 (N_14241,N_11660,N_11821);
and U14242 (N_14242,N_9752,N_11266);
and U14243 (N_14243,N_10924,N_11567);
xnor U14244 (N_14244,N_9249,N_10773);
and U14245 (N_14245,N_11836,N_10388);
and U14246 (N_14246,N_10456,N_11622);
or U14247 (N_14247,N_9052,N_11302);
and U14248 (N_14248,N_11102,N_11375);
nand U14249 (N_14249,N_11471,N_11407);
nor U14250 (N_14250,N_10485,N_11614);
and U14251 (N_14251,N_11180,N_9671);
nor U14252 (N_14252,N_9711,N_10559);
nor U14253 (N_14253,N_11376,N_9431);
and U14254 (N_14254,N_9942,N_9651);
or U14255 (N_14255,N_10979,N_11862);
or U14256 (N_14256,N_11766,N_11218);
or U14257 (N_14257,N_10058,N_9818);
or U14258 (N_14258,N_9227,N_9243);
nand U14259 (N_14259,N_11958,N_11234);
nor U14260 (N_14260,N_9491,N_11478);
or U14261 (N_14261,N_9202,N_10214);
xnor U14262 (N_14262,N_10623,N_10831);
nand U14263 (N_14263,N_9453,N_11629);
or U14264 (N_14264,N_9754,N_9066);
nand U14265 (N_14265,N_10230,N_9465);
nor U14266 (N_14266,N_11925,N_10058);
nor U14267 (N_14267,N_10764,N_11415);
nand U14268 (N_14268,N_11231,N_11694);
nand U14269 (N_14269,N_10202,N_9449);
and U14270 (N_14270,N_11160,N_10123);
nand U14271 (N_14271,N_9758,N_10844);
and U14272 (N_14272,N_11725,N_10766);
and U14273 (N_14273,N_9095,N_10266);
or U14274 (N_14274,N_9105,N_11809);
and U14275 (N_14275,N_9423,N_11387);
nand U14276 (N_14276,N_10450,N_9234);
or U14277 (N_14277,N_11926,N_9565);
and U14278 (N_14278,N_10223,N_11530);
nand U14279 (N_14279,N_11970,N_11277);
and U14280 (N_14280,N_10094,N_11672);
and U14281 (N_14281,N_11550,N_10249);
nand U14282 (N_14282,N_10415,N_10154);
and U14283 (N_14283,N_9721,N_11461);
or U14284 (N_14284,N_11861,N_11974);
xor U14285 (N_14285,N_10217,N_9657);
nor U14286 (N_14286,N_11020,N_9221);
nand U14287 (N_14287,N_10002,N_11866);
nor U14288 (N_14288,N_10810,N_9547);
or U14289 (N_14289,N_9605,N_9698);
nor U14290 (N_14290,N_11314,N_10883);
nand U14291 (N_14291,N_9965,N_9863);
xor U14292 (N_14292,N_9463,N_9509);
or U14293 (N_14293,N_9763,N_10085);
or U14294 (N_14294,N_10697,N_10176);
and U14295 (N_14295,N_11261,N_11221);
and U14296 (N_14296,N_9727,N_9667);
or U14297 (N_14297,N_9442,N_10126);
and U14298 (N_14298,N_10502,N_10857);
and U14299 (N_14299,N_11903,N_9051);
and U14300 (N_14300,N_10823,N_11219);
nor U14301 (N_14301,N_11313,N_11668);
nor U14302 (N_14302,N_9376,N_11064);
and U14303 (N_14303,N_9430,N_11994);
nand U14304 (N_14304,N_11367,N_11777);
and U14305 (N_14305,N_9053,N_9368);
or U14306 (N_14306,N_11447,N_11753);
or U14307 (N_14307,N_11144,N_9385);
nand U14308 (N_14308,N_9054,N_11347);
nand U14309 (N_14309,N_10642,N_11132);
nand U14310 (N_14310,N_10734,N_11153);
or U14311 (N_14311,N_9765,N_11213);
nand U14312 (N_14312,N_10596,N_9030);
nand U14313 (N_14313,N_11089,N_10176);
and U14314 (N_14314,N_11085,N_11181);
nor U14315 (N_14315,N_10144,N_11206);
nand U14316 (N_14316,N_9508,N_9357);
and U14317 (N_14317,N_9445,N_9464);
or U14318 (N_14318,N_9811,N_9332);
or U14319 (N_14319,N_9226,N_10586);
or U14320 (N_14320,N_10821,N_11114);
and U14321 (N_14321,N_9155,N_10782);
nand U14322 (N_14322,N_10634,N_10995);
nand U14323 (N_14323,N_9447,N_9473);
or U14324 (N_14324,N_10749,N_9872);
nor U14325 (N_14325,N_11122,N_10385);
nor U14326 (N_14326,N_10150,N_10815);
nor U14327 (N_14327,N_9156,N_10972);
nand U14328 (N_14328,N_11497,N_9529);
or U14329 (N_14329,N_11250,N_10363);
xor U14330 (N_14330,N_10812,N_11425);
nand U14331 (N_14331,N_11520,N_9911);
nand U14332 (N_14332,N_9186,N_10257);
and U14333 (N_14333,N_10842,N_11541);
nor U14334 (N_14334,N_10592,N_11238);
or U14335 (N_14335,N_9981,N_11775);
nor U14336 (N_14336,N_10515,N_10575);
nand U14337 (N_14337,N_10373,N_11515);
or U14338 (N_14338,N_10496,N_10134);
nor U14339 (N_14339,N_9183,N_11212);
nor U14340 (N_14340,N_9359,N_9339);
xor U14341 (N_14341,N_11517,N_11631);
nand U14342 (N_14342,N_9386,N_9405);
nor U14343 (N_14343,N_11536,N_10693);
nor U14344 (N_14344,N_10413,N_11099);
nand U14345 (N_14345,N_11076,N_9453);
nor U14346 (N_14346,N_11717,N_11071);
and U14347 (N_14347,N_10786,N_11832);
or U14348 (N_14348,N_9235,N_10398);
nand U14349 (N_14349,N_11755,N_11471);
nand U14350 (N_14350,N_11039,N_10211);
or U14351 (N_14351,N_10396,N_10916);
and U14352 (N_14352,N_10719,N_9374);
nand U14353 (N_14353,N_10814,N_9005);
and U14354 (N_14354,N_10715,N_11033);
nand U14355 (N_14355,N_11385,N_11961);
nor U14356 (N_14356,N_9218,N_11956);
nor U14357 (N_14357,N_11597,N_11048);
and U14358 (N_14358,N_11883,N_9316);
or U14359 (N_14359,N_10437,N_10927);
xnor U14360 (N_14360,N_11219,N_10997);
xnor U14361 (N_14361,N_11192,N_10927);
nand U14362 (N_14362,N_9853,N_9795);
nor U14363 (N_14363,N_10526,N_11496);
and U14364 (N_14364,N_11826,N_11680);
and U14365 (N_14365,N_10386,N_9291);
and U14366 (N_14366,N_11216,N_10782);
nor U14367 (N_14367,N_9428,N_10759);
and U14368 (N_14368,N_9862,N_9539);
and U14369 (N_14369,N_10739,N_10465);
or U14370 (N_14370,N_11627,N_9918);
nand U14371 (N_14371,N_11136,N_10912);
xnor U14372 (N_14372,N_11365,N_11330);
or U14373 (N_14373,N_10577,N_10562);
or U14374 (N_14374,N_9768,N_9104);
xnor U14375 (N_14375,N_10568,N_9124);
nor U14376 (N_14376,N_10691,N_11033);
or U14377 (N_14377,N_11445,N_11847);
nand U14378 (N_14378,N_11548,N_10216);
nand U14379 (N_14379,N_10741,N_9934);
nor U14380 (N_14380,N_11556,N_10915);
nand U14381 (N_14381,N_9157,N_11855);
and U14382 (N_14382,N_9705,N_9970);
nor U14383 (N_14383,N_10797,N_9723);
or U14384 (N_14384,N_9577,N_10283);
nand U14385 (N_14385,N_11003,N_9312);
and U14386 (N_14386,N_11757,N_11975);
and U14387 (N_14387,N_9249,N_9659);
xnor U14388 (N_14388,N_11393,N_11840);
nand U14389 (N_14389,N_11420,N_9848);
xnor U14390 (N_14390,N_10360,N_11171);
and U14391 (N_14391,N_9115,N_10656);
nand U14392 (N_14392,N_9859,N_9833);
nand U14393 (N_14393,N_11363,N_10788);
xor U14394 (N_14394,N_10548,N_10506);
nor U14395 (N_14395,N_11830,N_11198);
and U14396 (N_14396,N_10034,N_10484);
or U14397 (N_14397,N_9746,N_10810);
nor U14398 (N_14398,N_11878,N_11774);
nand U14399 (N_14399,N_9204,N_11635);
or U14400 (N_14400,N_10279,N_10681);
nand U14401 (N_14401,N_10702,N_9746);
and U14402 (N_14402,N_9458,N_11463);
and U14403 (N_14403,N_9368,N_9125);
nand U14404 (N_14404,N_10837,N_10724);
and U14405 (N_14405,N_9507,N_9112);
nand U14406 (N_14406,N_11304,N_9970);
or U14407 (N_14407,N_10437,N_9041);
nor U14408 (N_14408,N_9979,N_11705);
nor U14409 (N_14409,N_11037,N_10467);
or U14410 (N_14410,N_10499,N_10862);
nand U14411 (N_14411,N_10918,N_10612);
nand U14412 (N_14412,N_10956,N_9432);
nand U14413 (N_14413,N_10556,N_10613);
nor U14414 (N_14414,N_10066,N_9838);
nor U14415 (N_14415,N_11154,N_9459);
xor U14416 (N_14416,N_10001,N_10679);
nand U14417 (N_14417,N_11392,N_11345);
nor U14418 (N_14418,N_9969,N_11637);
nand U14419 (N_14419,N_10690,N_9907);
or U14420 (N_14420,N_11754,N_9368);
nand U14421 (N_14421,N_11971,N_10797);
or U14422 (N_14422,N_10445,N_10675);
nand U14423 (N_14423,N_9414,N_10617);
or U14424 (N_14424,N_9185,N_9889);
nand U14425 (N_14425,N_9720,N_10592);
or U14426 (N_14426,N_11283,N_10781);
and U14427 (N_14427,N_9662,N_9440);
or U14428 (N_14428,N_11356,N_11249);
nand U14429 (N_14429,N_11358,N_10244);
nand U14430 (N_14430,N_11848,N_9486);
nand U14431 (N_14431,N_11003,N_10577);
or U14432 (N_14432,N_10240,N_11763);
or U14433 (N_14433,N_11809,N_9261);
or U14434 (N_14434,N_9763,N_9951);
and U14435 (N_14435,N_9647,N_11332);
nor U14436 (N_14436,N_10994,N_11712);
nor U14437 (N_14437,N_10762,N_10390);
nor U14438 (N_14438,N_10705,N_10345);
or U14439 (N_14439,N_9214,N_9752);
nor U14440 (N_14440,N_10521,N_9926);
or U14441 (N_14441,N_11308,N_10320);
nor U14442 (N_14442,N_11992,N_10421);
nand U14443 (N_14443,N_10355,N_11194);
nor U14444 (N_14444,N_11130,N_11628);
nor U14445 (N_14445,N_10357,N_11982);
nor U14446 (N_14446,N_10327,N_11413);
xnor U14447 (N_14447,N_11696,N_10770);
nand U14448 (N_14448,N_9028,N_9776);
nand U14449 (N_14449,N_9680,N_10755);
or U14450 (N_14450,N_11788,N_9465);
nand U14451 (N_14451,N_10115,N_11881);
nor U14452 (N_14452,N_9881,N_10780);
or U14453 (N_14453,N_10669,N_11575);
xor U14454 (N_14454,N_11810,N_11521);
and U14455 (N_14455,N_10175,N_9079);
and U14456 (N_14456,N_9823,N_11439);
and U14457 (N_14457,N_11000,N_11328);
and U14458 (N_14458,N_10903,N_10090);
or U14459 (N_14459,N_10387,N_11838);
xnor U14460 (N_14460,N_9518,N_9145);
nand U14461 (N_14461,N_11114,N_10707);
nor U14462 (N_14462,N_10277,N_10467);
or U14463 (N_14463,N_10679,N_9088);
nand U14464 (N_14464,N_9583,N_11593);
xor U14465 (N_14465,N_9727,N_10219);
and U14466 (N_14466,N_9758,N_11422);
nand U14467 (N_14467,N_10956,N_11453);
and U14468 (N_14468,N_9040,N_11309);
nand U14469 (N_14469,N_10867,N_11300);
or U14470 (N_14470,N_10906,N_9226);
nor U14471 (N_14471,N_9131,N_10660);
or U14472 (N_14472,N_10820,N_9776);
nand U14473 (N_14473,N_10009,N_9997);
and U14474 (N_14474,N_9373,N_11565);
nand U14475 (N_14475,N_11736,N_10432);
nor U14476 (N_14476,N_11704,N_11932);
and U14477 (N_14477,N_10061,N_9748);
or U14478 (N_14478,N_11199,N_9988);
nor U14479 (N_14479,N_9038,N_9968);
or U14480 (N_14480,N_10738,N_10681);
or U14481 (N_14481,N_9735,N_10616);
nand U14482 (N_14482,N_11665,N_10253);
or U14483 (N_14483,N_10933,N_9985);
nor U14484 (N_14484,N_10636,N_9206);
and U14485 (N_14485,N_9255,N_10880);
nand U14486 (N_14486,N_10265,N_10453);
nor U14487 (N_14487,N_9071,N_9237);
or U14488 (N_14488,N_9284,N_10717);
nor U14489 (N_14489,N_11261,N_10668);
nand U14490 (N_14490,N_9441,N_11226);
nor U14491 (N_14491,N_9581,N_11343);
nand U14492 (N_14492,N_11177,N_11666);
nand U14493 (N_14493,N_11419,N_11265);
and U14494 (N_14494,N_10994,N_9807);
nor U14495 (N_14495,N_10030,N_9745);
nor U14496 (N_14496,N_11913,N_9833);
xor U14497 (N_14497,N_9147,N_11956);
and U14498 (N_14498,N_11985,N_9883);
xnor U14499 (N_14499,N_9574,N_10796);
nor U14500 (N_14500,N_10474,N_11762);
and U14501 (N_14501,N_10662,N_10343);
nor U14502 (N_14502,N_11523,N_9223);
or U14503 (N_14503,N_11157,N_9715);
nor U14504 (N_14504,N_11747,N_10090);
or U14505 (N_14505,N_10578,N_10698);
or U14506 (N_14506,N_10227,N_10149);
and U14507 (N_14507,N_9474,N_9915);
nand U14508 (N_14508,N_11501,N_9871);
xnor U14509 (N_14509,N_9271,N_11714);
and U14510 (N_14510,N_10750,N_9738);
nand U14511 (N_14511,N_11624,N_9353);
xor U14512 (N_14512,N_9369,N_11570);
xor U14513 (N_14513,N_9365,N_9832);
or U14514 (N_14514,N_11333,N_9208);
nor U14515 (N_14515,N_11325,N_9664);
nand U14516 (N_14516,N_9870,N_11948);
nand U14517 (N_14517,N_11283,N_11301);
or U14518 (N_14518,N_10703,N_10445);
nor U14519 (N_14519,N_10510,N_11776);
or U14520 (N_14520,N_10876,N_10988);
or U14521 (N_14521,N_9658,N_9118);
xor U14522 (N_14522,N_10328,N_9149);
or U14523 (N_14523,N_9690,N_10674);
xnor U14524 (N_14524,N_9763,N_10618);
and U14525 (N_14525,N_9836,N_11717);
nor U14526 (N_14526,N_11434,N_9113);
or U14527 (N_14527,N_11977,N_11537);
or U14528 (N_14528,N_10013,N_10450);
nor U14529 (N_14529,N_9074,N_10660);
nor U14530 (N_14530,N_9293,N_9954);
xnor U14531 (N_14531,N_10262,N_10473);
or U14532 (N_14532,N_10081,N_11122);
or U14533 (N_14533,N_11268,N_10892);
or U14534 (N_14534,N_11136,N_10575);
and U14535 (N_14535,N_11080,N_10370);
nor U14536 (N_14536,N_10548,N_9592);
or U14537 (N_14537,N_11432,N_9775);
nor U14538 (N_14538,N_9220,N_9521);
nor U14539 (N_14539,N_11907,N_11977);
and U14540 (N_14540,N_10586,N_9441);
nor U14541 (N_14541,N_11385,N_11707);
and U14542 (N_14542,N_10220,N_9283);
or U14543 (N_14543,N_11102,N_9305);
nor U14544 (N_14544,N_9857,N_11966);
and U14545 (N_14545,N_10652,N_10355);
and U14546 (N_14546,N_11750,N_10922);
and U14547 (N_14547,N_9516,N_10010);
and U14548 (N_14548,N_11103,N_10525);
or U14549 (N_14549,N_10617,N_9375);
nor U14550 (N_14550,N_9535,N_9338);
or U14551 (N_14551,N_11811,N_11829);
and U14552 (N_14552,N_10052,N_11246);
nand U14553 (N_14553,N_9968,N_11177);
xor U14554 (N_14554,N_11601,N_10831);
or U14555 (N_14555,N_11953,N_11747);
or U14556 (N_14556,N_10047,N_9221);
nor U14557 (N_14557,N_11033,N_11558);
or U14558 (N_14558,N_10843,N_11750);
nor U14559 (N_14559,N_10815,N_11322);
or U14560 (N_14560,N_11979,N_9529);
and U14561 (N_14561,N_9446,N_9376);
and U14562 (N_14562,N_11711,N_10393);
xnor U14563 (N_14563,N_9077,N_9494);
or U14564 (N_14564,N_10778,N_9646);
or U14565 (N_14565,N_11506,N_10066);
nor U14566 (N_14566,N_11596,N_9697);
nor U14567 (N_14567,N_11325,N_10102);
or U14568 (N_14568,N_9110,N_10163);
or U14569 (N_14569,N_9827,N_11119);
and U14570 (N_14570,N_11495,N_10380);
nand U14571 (N_14571,N_11602,N_9445);
or U14572 (N_14572,N_9290,N_10617);
nand U14573 (N_14573,N_9059,N_10025);
and U14574 (N_14574,N_9846,N_11405);
or U14575 (N_14575,N_10022,N_9106);
and U14576 (N_14576,N_10358,N_10407);
and U14577 (N_14577,N_10367,N_11473);
and U14578 (N_14578,N_9654,N_10532);
or U14579 (N_14579,N_11817,N_11869);
or U14580 (N_14580,N_10944,N_10017);
or U14581 (N_14581,N_9908,N_10039);
nand U14582 (N_14582,N_11776,N_9026);
nand U14583 (N_14583,N_10386,N_11119);
xor U14584 (N_14584,N_9805,N_11381);
nor U14585 (N_14585,N_10075,N_10562);
and U14586 (N_14586,N_9565,N_9038);
or U14587 (N_14587,N_9025,N_11720);
nand U14588 (N_14588,N_10123,N_9128);
nand U14589 (N_14589,N_10942,N_10731);
nor U14590 (N_14590,N_9944,N_10926);
or U14591 (N_14591,N_11784,N_11412);
or U14592 (N_14592,N_11779,N_11016);
or U14593 (N_14593,N_9585,N_11072);
or U14594 (N_14594,N_10840,N_10422);
and U14595 (N_14595,N_10954,N_9358);
nor U14596 (N_14596,N_11184,N_11836);
nor U14597 (N_14597,N_10738,N_10074);
or U14598 (N_14598,N_9248,N_9862);
or U14599 (N_14599,N_11273,N_11890);
nor U14600 (N_14600,N_10675,N_9329);
nor U14601 (N_14601,N_10336,N_11646);
nor U14602 (N_14602,N_11923,N_10862);
xor U14603 (N_14603,N_11834,N_10566);
or U14604 (N_14604,N_11020,N_9090);
and U14605 (N_14605,N_11600,N_11378);
and U14606 (N_14606,N_10642,N_11963);
xor U14607 (N_14607,N_9149,N_9747);
and U14608 (N_14608,N_9645,N_9327);
or U14609 (N_14609,N_11901,N_9702);
or U14610 (N_14610,N_10232,N_9517);
nor U14611 (N_14611,N_9180,N_9114);
and U14612 (N_14612,N_10411,N_10817);
or U14613 (N_14613,N_9924,N_10522);
and U14614 (N_14614,N_10367,N_11806);
nand U14615 (N_14615,N_9059,N_11430);
nor U14616 (N_14616,N_11805,N_10399);
or U14617 (N_14617,N_9563,N_9500);
nand U14618 (N_14618,N_9648,N_10035);
nand U14619 (N_14619,N_10044,N_9250);
nand U14620 (N_14620,N_11562,N_10534);
and U14621 (N_14621,N_10745,N_11730);
or U14622 (N_14622,N_11114,N_9030);
and U14623 (N_14623,N_9725,N_10081);
and U14624 (N_14624,N_10268,N_10403);
nor U14625 (N_14625,N_9348,N_9439);
nor U14626 (N_14626,N_11438,N_10413);
and U14627 (N_14627,N_10677,N_9966);
or U14628 (N_14628,N_11600,N_11129);
or U14629 (N_14629,N_9984,N_11482);
and U14630 (N_14630,N_9930,N_10203);
or U14631 (N_14631,N_11475,N_11408);
and U14632 (N_14632,N_9517,N_9707);
nor U14633 (N_14633,N_11275,N_10169);
nor U14634 (N_14634,N_9570,N_9695);
and U14635 (N_14635,N_11454,N_9188);
or U14636 (N_14636,N_10431,N_11259);
or U14637 (N_14637,N_10760,N_11853);
nor U14638 (N_14638,N_11319,N_10501);
nand U14639 (N_14639,N_10778,N_9928);
nor U14640 (N_14640,N_10177,N_10831);
or U14641 (N_14641,N_10312,N_11731);
nor U14642 (N_14642,N_11712,N_9969);
xnor U14643 (N_14643,N_10071,N_9754);
nor U14644 (N_14644,N_11064,N_9263);
nor U14645 (N_14645,N_11820,N_10794);
nand U14646 (N_14646,N_10547,N_11983);
nand U14647 (N_14647,N_11575,N_9145);
nor U14648 (N_14648,N_11498,N_11596);
and U14649 (N_14649,N_9621,N_9093);
or U14650 (N_14650,N_11210,N_10730);
and U14651 (N_14651,N_9431,N_9212);
or U14652 (N_14652,N_10627,N_10572);
nor U14653 (N_14653,N_11408,N_9108);
nand U14654 (N_14654,N_11215,N_9693);
nand U14655 (N_14655,N_10589,N_11726);
xnor U14656 (N_14656,N_11365,N_9366);
nand U14657 (N_14657,N_9984,N_11485);
or U14658 (N_14658,N_10602,N_9286);
nor U14659 (N_14659,N_11874,N_11017);
or U14660 (N_14660,N_10758,N_11703);
and U14661 (N_14661,N_10898,N_11582);
and U14662 (N_14662,N_10434,N_9326);
nor U14663 (N_14663,N_9523,N_11083);
nor U14664 (N_14664,N_11529,N_9777);
nand U14665 (N_14665,N_11710,N_9534);
and U14666 (N_14666,N_9068,N_9287);
and U14667 (N_14667,N_9537,N_10430);
nor U14668 (N_14668,N_10166,N_11472);
or U14669 (N_14669,N_9179,N_9134);
xnor U14670 (N_14670,N_10483,N_10890);
or U14671 (N_14671,N_9208,N_10831);
or U14672 (N_14672,N_10844,N_9942);
nor U14673 (N_14673,N_9144,N_10500);
nand U14674 (N_14674,N_11290,N_10176);
xor U14675 (N_14675,N_9287,N_11126);
and U14676 (N_14676,N_11611,N_11782);
or U14677 (N_14677,N_11785,N_11310);
nor U14678 (N_14678,N_11685,N_9771);
or U14679 (N_14679,N_9455,N_10889);
and U14680 (N_14680,N_10109,N_10523);
and U14681 (N_14681,N_11282,N_11216);
and U14682 (N_14682,N_9092,N_9341);
and U14683 (N_14683,N_9745,N_9735);
xnor U14684 (N_14684,N_9908,N_11354);
nand U14685 (N_14685,N_11838,N_11649);
and U14686 (N_14686,N_10724,N_10894);
or U14687 (N_14687,N_10140,N_9096);
or U14688 (N_14688,N_11579,N_9143);
or U14689 (N_14689,N_10754,N_10192);
nor U14690 (N_14690,N_9665,N_10217);
nand U14691 (N_14691,N_9944,N_11418);
or U14692 (N_14692,N_9869,N_10241);
nor U14693 (N_14693,N_10623,N_9652);
nand U14694 (N_14694,N_11966,N_11491);
nor U14695 (N_14695,N_9654,N_10711);
nand U14696 (N_14696,N_11113,N_10957);
nand U14697 (N_14697,N_10943,N_9027);
or U14698 (N_14698,N_9091,N_10026);
nor U14699 (N_14699,N_9071,N_11181);
nor U14700 (N_14700,N_10561,N_11223);
nand U14701 (N_14701,N_11433,N_11558);
xnor U14702 (N_14702,N_9887,N_9047);
and U14703 (N_14703,N_9021,N_9684);
xnor U14704 (N_14704,N_11332,N_11920);
or U14705 (N_14705,N_9144,N_9301);
or U14706 (N_14706,N_10200,N_9593);
nand U14707 (N_14707,N_10994,N_11912);
and U14708 (N_14708,N_11398,N_10053);
nor U14709 (N_14709,N_9446,N_10559);
and U14710 (N_14710,N_11780,N_10220);
nor U14711 (N_14711,N_9043,N_9943);
or U14712 (N_14712,N_10899,N_10608);
or U14713 (N_14713,N_10527,N_9693);
or U14714 (N_14714,N_11685,N_10267);
nor U14715 (N_14715,N_9582,N_11998);
nand U14716 (N_14716,N_10538,N_11112);
and U14717 (N_14717,N_10183,N_10569);
or U14718 (N_14718,N_10494,N_9766);
and U14719 (N_14719,N_9339,N_10202);
or U14720 (N_14720,N_10532,N_9484);
or U14721 (N_14721,N_11812,N_10007);
nand U14722 (N_14722,N_10594,N_11411);
and U14723 (N_14723,N_9603,N_11932);
nor U14724 (N_14724,N_11425,N_10280);
or U14725 (N_14725,N_9070,N_9984);
nand U14726 (N_14726,N_9416,N_11898);
and U14727 (N_14727,N_10482,N_9211);
and U14728 (N_14728,N_10433,N_9640);
nor U14729 (N_14729,N_9758,N_11749);
or U14730 (N_14730,N_11165,N_11197);
and U14731 (N_14731,N_9471,N_9996);
nor U14732 (N_14732,N_10763,N_9102);
and U14733 (N_14733,N_10139,N_10241);
or U14734 (N_14734,N_9743,N_9347);
nand U14735 (N_14735,N_10673,N_9944);
or U14736 (N_14736,N_11143,N_9972);
or U14737 (N_14737,N_10760,N_10292);
nand U14738 (N_14738,N_11373,N_9468);
or U14739 (N_14739,N_10045,N_11522);
nor U14740 (N_14740,N_9438,N_11286);
and U14741 (N_14741,N_10103,N_9294);
nor U14742 (N_14742,N_10749,N_11055);
or U14743 (N_14743,N_11328,N_11356);
and U14744 (N_14744,N_11032,N_10554);
xor U14745 (N_14745,N_11522,N_11715);
xor U14746 (N_14746,N_9840,N_10326);
xnor U14747 (N_14747,N_10556,N_9153);
nand U14748 (N_14748,N_9804,N_9575);
or U14749 (N_14749,N_9433,N_9516);
xor U14750 (N_14750,N_10338,N_11912);
or U14751 (N_14751,N_11678,N_9073);
and U14752 (N_14752,N_10478,N_10971);
nand U14753 (N_14753,N_9298,N_9449);
and U14754 (N_14754,N_9800,N_9691);
and U14755 (N_14755,N_10647,N_9697);
or U14756 (N_14756,N_10585,N_9180);
or U14757 (N_14757,N_9526,N_10361);
nand U14758 (N_14758,N_9094,N_9270);
and U14759 (N_14759,N_11052,N_10216);
xnor U14760 (N_14760,N_11768,N_10073);
nor U14761 (N_14761,N_9395,N_11117);
nor U14762 (N_14762,N_10964,N_9261);
xor U14763 (N_14763,N_11130,N_10662);
or U14764 (N_14764,N_11920,N_11302);
or U14765 (N_14765,N_9845,N_10984);
nand U14766 (N_14766,N_11894,N_11192);
and U14767 (N_14767,N_11140,N_11078);
and U14768 (N_14768,N_10514,N_10573);
nand U14769 (N_14769,N_11867,N_11639);
or U14770 (N_14770,N_11497,N_10126);
nand U14771 (N_14771,N_9304,N_11786);
nor U14772 (N_14772,N_10927,N_11261);
nor U14773 (N_14773,N_10182,N_10362);
and U14774 (N_14774,N_9952,N_10058);
or U14775 (N_14775,N_10361,N_11236);
xnor U14776 (N_14776,N_10320,N_10605);
and U14777 (N_14777,N_11773,N_10186);
nand U14778 (N_14778,N_9819,N_11173);
or U14779 (N_14779,N_11710,N_9117);
nor U14780 (N_14780,N_11781,N_11080);
xnor U14781 (N_14781,N_10772,N_11076);
and U14782 (N_14782,N_9077,N_11655);
xor U14783 (N_14783,N_10798,N_11595);
and U14784 (N_14784,N_11172,N_9838);
nand U14785 (N_14785,N_10297,N_10923);
nand U14786 (N_14786,N_11971,N_10831);
and U14787 (N_14787,N_10872,N_9201);
or U14788 (N_14788,N_11627,N_9853);
or U14789 (N_14789,N_10319,N_9300);
nor U14790 (N_14790,N_9162,N_10869);
xor U14791 (N_14791,N_11725,N_11939);
xnor U14792 (N_14792,N_9001,N_11550);
and U14793 (N_14793,N_9169,N_11007);
nand U14794 (N_14794,N_10061,N_9072);
nand U14795 (N_14795,N_9525,N_9338);
nor U14796 (N_14796,N_9575,N_11767);
or U14797 (N_14797,N_11935,N_9956);
and U14798 (N_14798,N_11046,N_11100);
nand U14799 (N_14799,N_9065,N_10536);
and U14800 (N_14800,N_10918,N_11802);
and U14801 (N_14801,N_10405,N_10418);
and U14802 (N_14802,N_11526,N_10851);
or U14803 (N_14803,N_10966,N_9101);
nand U14804 (N_14804,N_10219,N_11999);
or U14805 (N_14805,N_11903,N_10400);
nor U14806 (N_14806,N_10895,N_10958);
nand U14807 (N_14807,N_10827,N_9705);
nand U14808 (N_14808,N_11367,N_10044);
and U14809 (N_14809,N_10521,N_10284);
nand U14810 (N_14810,N_9801,N_9942);
or U14811 (N_14811,N_11381,N_10684);
and U14812 (N_14812,N_10041,N_9356);
or U14813 (N_14813,N_11119,N_10591);
nand U14814 (N_14814,N_11483,N_11140);
and U14815 (N_14815,N_9755,N_10399);
or U14816 (N_14816,N_9324,N_10512);
nor U14817 (N_14817,N_11947,N_9580);
nor U14818 (N_14818,N_9977,N_10987);
nand U14819 (N_14819,N_9529,N_9667);
nand U14820 (N_14820,N_10538,N_11106);
or U14821 (N_14821,N_11121,N_9619);
or U14822 (N_14822,N_10978,N_10525);
or U14823 (N_14823,N_10778,N_10010);
and U14824 (N_14824,N_11097,N_9616);
nor U14825 (N_14825,N_11416,N_11362);
nand U14826 (N_14826,N_11836,N_11835);
nor U14827 (N_14827,N_11724,N_11917);
xnor U14828 (N_14828,N_10373,N_11278);
nor U14829 (N_14829,N_10864,N_10439);
nand U14830 (N_14830,N_9523,N_11660);
or U14831 (N_14831,N_11403,N_9579);
xor U14832 (N_14832,N_10519,N_11424);
or U14833 (N_14833,N_9517,N_9365);
xnor U14834 (N_14834,N_10922,N_11239);
nor U14835 (N_14835,N_11696,N_9890);
nand U14836 (N_14836,N_9114,N_11193);
and U14837 (N_14837,N_10586,N_11420);
and U14838 (N_14838,N_10412,N_11065);
or U14839 (N_14839,N_11358,N_10798);
and U14840 (N_14840,N_10881,N_11901);
and U14841 (N_14841,N_10849,N_11644);
nor U14842 (N_14842,N_9069,N_10861);
xnor U14843 (N_14843,N_10610,N_10010);
nand U14844 (N_14844,N_9171,N_10401);
and U14845 (N_14845,N_11774,N_10992);
and U14846 (N_14846,N_9610,N_9423);
and U14847 (N_14847,N_10845,N_10503);
nand U14848 (N_14848,N_11032,N_10594);
and U14849 (N_14849,N_9412,N_9539);
nor U14850 (N_14850,N_10624,N_9280);
and U14851 (N_14851,N_9387,N_10347);
nand U14852 (N_14852,N_10957,N_10055);
nor U14853 (N_14853,N_9600,N_11001);
and U14854 (N_14854,N_9685,N_11753);
nand U14855 (N_14855,N_11483,N_11848);
nand U14856 (N_14856,N_11159,N_9546);
nand U14857 (N_14857,N_10355,N_10570);
nand U14858 (N_14858,N_9756,N_9897);
nor U14859 (N_14859,N_10638,N_10850);
and U14860 (N_14860,N_9551,N_11038);
and U14861 (N_14861,N_9943,N_11821);
nor U14862 (N_14862,N_11045,N_10867);
nand U14863 (N_14863,N_9080,N_9378);
nor U14864 (N_14864,N_10861,N_9821);
and U14865 (N_14865,N_11435,N_10084);
nor U14866 (N_14866,N_9626,N_9483);
xnor U14867 (N_14867,N_9679,N_10031);
nand U14868 (N_14868,N_11704,N_9455);
nand U14869 (N_14869,N_9826,N_10146);
xor U14870 (N_14870,N_9329,N_10409);
xnor U14871 (N_14871,N_9556,N_9877);
nor U14872 (N_14872,N_10666,N_10078);
nor U14873 (N_14873,N_9911,N_9133);
xnor U14874 (N_14874,N_10547,N_9238);
nand U14875 (N_14875,N_11988,N_10127);
nor U14876 (N_14876,N_10829,N_10079);
and U14877 (N_14877,N_10093,N_9739);
nor U14878 (N_14878,N_10575,N_9338);
or U14879 (N_14879,N_10978,N_9114);
nor U14880 (N_14880,N_10185,N_9283);
or U14881 (N_14881,N_11677,N_10776);
nand U14882 (N_14882,N_9072,N_10955);
and U14883 (N_14883,N_9882,N_10219);
nor U14884 (N_14884,N_9905,N_9443);
nor U14885 (N_14885,N_10751,N_10873);
or U14886 (N_14886,N_10207,N_10426);
nor U14887 (N_14887,N_10734,N_9215);
or U14888 (N_14888,N_11819,N_11642);
and U14889 (N_14889,N_10964,N_10327);
nor U14890 (N_14890,N_9257,N_9864);
nor U14891 (N_14891,N_9691,N_9467);
nand U14892 (N_14892,N_9016,N_11973);
nor U14893 (N_14893,N_11366,N_11212);
or U14894 (N_14894,N_9810,N_11198);
and U14895 (N_14895,N_10061,N_10038);
nand U14896 (N_14896,N_9446,N_9887);
nand U14897 (N_14897,N_10943,N_10676);
and U14898 (N_14898,N_9697,N_11903);
nand U14899 (N_14899,N_11803,N_10904);
xnor U14900 (N_14900,N_11176,N_11868);
xnor U14901 (N_14901,N_10860,N_10110);
nor U14902 (N_14902,N_9637,N_9757);
nand U14903 (N_14903,N_10096,N_9189);
and U14904 (N_14904,N_11398,N_10631);
nand U14905 (N_14905,N_9158,N_10897);
nand U14906 (N_14906,N_9548,N_9770);
nand U14907 (N_14907,N_11884,N_9866);
nand U14908 (N_14908,N_11013,N_11609);
nor U14909 (N_14909,N_9251,N_10508);
nand U14910 (N_14910,N_11207,N_9399);
and U14911 (N_14911,N_10420,N_10532);
nor U14912 (N_14912,N_11265,N_11902);
nand U14913 (N_14913,N_9688,N_10946);
and U14914 (N_14914,N_10254,N_10385);
xnor U14915 (N_14915,N_9175,N_10538);
nor U14916 (N_14916,N_10016,N_11084);
nand U14917 (N_14917,N_10693,N_9633);
or U14918 (N_14918,N_10679,N_10866);
nand U14919 (N_14919,N_9945,N_9905);
and U14920 (N_14920,N_9561,N_9371);
nor U14921 (N_14921,N_11470,N_9474);
xor U14922 (N_14922,N_10350,N_11444);
nor U14923 (N_14923,N_10352,N_10239);
nor U14924 (N_14924,N_10967,N_9235);
nor U14925 (N_14925,N_11436,N_9856);
and U14926 (N_14926,N_11218,N_11461);
nand U14927 (N_14927,N_9182,N_10129);
and U14928 (N_14928,N_9499,N_10548);
or U14929 (N_14929,N_11950,N_11884);
nor U14930 (N_14930,N_10139,N_11677);
nand U14931 (N_14931,N_9752,N_11778);
nand U14932 (N_14932,N_11442,N_11713);
nor U14933 (N_14933,N_10057,N_10853);
or U14934 (N_14934,N_11528,N_10277);
xnor U14935 (N_14935,N_9324,N_11562);
xnor U14936 (N_14936,N_10710,N_10163);
nand U14937 (N_14937,N_11229,N_10505);
or U14938 (N_14938,N_9718,N_11743);
and U14939 (N_14939,N_10177,N_9914);
nor U14940 (N_14940,N_10728,N_10522);
or U14941 (N_14941,N_9977,N_11917);
nor U14942 (N_14942,N_11784,N_9990);
nand U14943 (N_14943,N_11780,N_11334);
nor U14944 (N_14944,N_10224,N_9731);
nand U14945 (N_14945,N_9488,N_9673);
xor U14946 (N_14946,N_10549,N_10231);
and U14947 (N_14947,N_10320,N_9072);
nand U14948 (N_14948,N_9185,N_10605);
xnor U14949 (N_14949,N_10825,N_9223);
nand U14950 (N_14950,N_10971,N_10939);
and U14951 (N_14951,N_11542,N_9763);
nand U14952 (N_14952,N_9785,N_10358);
nand U14953 (N_14953,N_9533,N_11500);
nor U14954 (N_14954,N_11299,N_10576);
xor U14955 (N_14955,N_11744,N_11575);
nor U14956 (N_14956,N_9865,N_10067);
or U14957 (N_14957,N_9934,N_9147);
and U14958 (N_14958,N_11208,N_9056);
and U14959 (N_14959,N_11831,N_11181);
or U14960 (N_14960,N_11988,N_11532);
or U14961 (N_14961,N_11858,N_9502);
and U14962 (N_14962,N_11901,N_9778);
and U14963 (N_14963,N_11689,N_9427);
and U14964 (N_14964,N_11525,N_11705);
or U14965 (N_14965,N_9860,N_10680);
and U14966 (N_14966,N_10685,N_11500);
nand U14967 (N_14967,N_9355,N_10392);
nand U14968 (N_14968,N_11590,N_10875);
nor U14969 (N_14969,N_9966,N_10713);
nor U14970 (N_14970,N_11965,N_10527);
nor U14971 (N_14971,N_11027,N_9491);
or U14972 (N_14972,N_11463,N_11253);
or U14973 (N_14973,N_11097,N_11400);
nor U14974 (N_14974,N_11466,N_11247);
and U14975 (N_14975,N_9131,N_10306);
nand U14976 (N_14976,N_11982,N_9986);
xnor U14977 (N_14977,N_10823,N_9062);
and U14978 (N_14978,N_9969,N_11449);
xnor U14979 (N_14979,N_10284,N_10557);
nand U14980 (N_14980,N_10176,N_10705);
nor U14981 (N_14981,N_11630,N_11682);
and U14982 (N_14982,N_10576,N_10401);
nand U14983 (N_14983,N_11765,N_9674);
nand U14984 (N_14984,N_9310,N_11896);
or U14985 (N_14985,N_9624,N_9967);
and U14986 (N_14986,N_11270,N_10479);
and U14987 (N_14987,N_10981,N_9878);
or U14988 (N_14988,N_10868,N_11580);
and U14989 (N_14989,N_11953,N_11655);
nor U14990 (N_14990,N_10233,N_9449);
and U14991 (N_14991,N_10232,N_11739);
nand U14992 (N_14992,N_10205,N_9205);
nand U14993 (N_14993,N_9976,N_11858);
xor U14994 (N_14994,N_11171,N_11537);
nor U14995 (N_14995,N_9086,N_9053);
or U14996 (N_14996,N_11808,N_9839);
and U14997 (N_14997,N_10494,N_11901);
or U14998 (N_14998,N_9415,N_10150);
or U14999 (N_14999,N_9196,N_11589);
nor U15000 (N_15000,N_13572,N_12757);
nand U15001 (N_15001,N_14641,N_12470);
nor U15002 (N_15002,N_14992,N_13034);
nand U15003 (N_15003,N_14249,N_13608);
nand U15004 (N_15004,N_14300,N_14807);
nand U15005 (N_15005,N_14773,N_13318);
nand U15006 (N_15006,N_14377,N_13407);
nand U15007 (N_15007,N_14663,N_13039);
or U15008 (N_15008,N_12129,N_13718);
or U15009 (N_15009,N_12662,N_13459);
nand U15010 (N_15010,N_13184,N_13835);
nor U15011 (N_15011,N_14699,N_13732);
nand U15012 (N_15012,N_14533,N_12814);
nor U15013 (N_15013,N_12257,N_12824);
and U15014 (N_15014,N_13522,N_14809);
or U15015 (N_15015,N_12748,N_14906);
or U15016 (N_15016,N_13719,N_13766);
nand U15017 (N_15017,N_14778,N_13383);
nor U15018 (N_15018,N_13616,N_14870);
or U15019 (N_15019,N_14536,N_12039);
xnor U15020 (N_15020,N_12144,N_14787);
xor U15021 (N_15021,N_14475,N_13514);
and U15022 (N_15022,N_12977,N_12058);
nor U15023 (N_15023,N_12013,N_14147);
nor U15024 (N_15024,N_13912,N_12186);
and U15025 (N_15025,N_14597,N_12961);
and U15026 (N_15026,N_12167,N_13689);
and U15027 (N_15027,N_12951,N_12958);
nand U15028 (N_15028,N_14901,N_14605);
or U15029 (N_15029,N_14935,N_13927);
and U15030 (N_15030,N_13907,N_14666);
nor U15031 (N_15031,N_13177,N_14818);
nor U15032 (N_15032,N_12028,N_12721);
and U15033 (N_15033,N_12934,N_12469);
and U15034 (N_15034,N_13294,N_14329);
and U15035 (N_15035,N_14980,N_14683);
nor U15036 (N_15036,N_12691,N_13140);
nor U15037 (N_15037,N_14640,N_14917);
nor U15038 (N_15038,N_14211,N_13623);
and U15039 (N_15039,N_13391,N_12648);
nor U15040 (N_15040,N_13588,N_14722);
nand U15041 (N_15041,N_12114,N_13811);
xnor U15042 (N_15042,N_13883,N_14301);
and U15043 (N_15043,N_13631,N_13108);
nand U15044 (N_15044,N_12932,N_14647);
nand U15045 (N_15045,N_12917,N_13508);
or U15046 (N_15046,N_13743,N_13581);
xnor U15047 (N_15047,N_12450,N_14355);
nor U15048 (N_15048,N_14658,N_14631);
or U15049 (N_15049,N_12991,N_13001);
xnor U15050 (N_15050,N_14720,N_14462);
nor U15051 (N_15051,N_12635,N_12248);
and U15052 (N_15052,N_14039,N_13491);
nand U15053 (N_15053,N_12338,N_14817);
nand U15054 (N_15054,N_12707,N_12295);
nand U15055 (N_15055,N_14276,N_14841);
and U15056 (N_15056,N_13392,N_12240);
or U15057 (N_15057,N_13528,N_12610);
xnor U15058 (N_15058,N_12014,N_13729);
nand U15059 (N_15059,N_13535,N_14823);
nand U15060 (N_15060,N_12441,N_13541);
and U15061 (N_15061,N_12092,N_13710);
or U15062 (N_15062,N_13244,N_13401);
nand U15063 (N_15063,N_13022,N_13991);
xor U15064 (N_15064,N_13076,N_13339);
nand U15065 (N_15065,N_14503,N_14168);
and U15066 (N_15066,N_12145,N_12698);
and U15067 (N_15067,N_13409,N_14714);
nand U15068 (N_15068,N_14950,N_13788);
nand U15069 (N_15069,N_12916,N_13837);
nand U15070 (N_15070,N_13063,N_12402);
nor U15071 (N_15071,N_12359,N_13791);
nand U15072 (N_15072,N_12363,N_14471);
xor U15073 (N_15073,N_14520,N_13727);
and U15074 (N_15074,N_13798,N_13029);
nor U15075 (N_15075,N_13259,N_12084);
nand U15076 (N_15076,N_14534,N_14375);
xnor U15077 (N_15077,N_14087,N_13361);
nor U15078 (N_15078,N_12633,N_12752);
or U15079 (N_15079,N_13266,N_12802);
or U15080 (N_15080,N_14280,N_14441);
nor U15081 (N_15081,N_14885,N_12876);
nor U15082 (N_15082,N_14439,N_14248);
and U15083 (N_15083,N_14975,N_14508);
nor U15084 (N_15084,N_13537,N_13260);
or U15085 (N_15085,N_13525,N_14042);
nand U15086 (N_15086,N_14972,N_13114);
nor U15087 (N_15087,N_14483,N_12930);
and U15088 (N_15088,N_14794,N_14660);
nor U15089 (N_15089,N_14379,N_13340);
nand U15090 (N_15090,N_13810,N_14584);
nand U15091 (N_15091,N_12526,N_12592);
or U15092 (N_15092,N_13834,N_12121);
or U15093 (N_15093,N_12063,N_13731);
nand U15094 (N_15094,N_12712,N_14792);
nor U15095 (N_15095,N_14112,N_12866);
or U15096 (N_15096,N_12361,N_12858);
nor U15097 (N_15097,N_12787,N_13609);
nand U15098 (N_15098,N_13355,N_14900);
nor U15099 (N_15099,N_12751,N_12534);
nor U15100 (N_15100,N_12889,N_14532);
nor U15101 (N_15101,N_14299,N_13128);
nand U15102 (N_15102,N_13571,N_14389);
or U15103 (N_15103,N_12139,N_13136);
nand U15104 (N_15104,N_14550,N_14850);
or U15105 (N_15105,N_12856,N_14421);
or U15106 (N_15106,N_13901,N_14590);
or U15107 (N_15107,N_13526,N_12815);
and U15108 (N_15108,N_14799,N_12126);
and U15109 (N_15109,N_12180,N_13078);
or U15110 (N_15110,N_14037,N_12510);
or U15111 (N_15111,N_13456,N_14750);
nor U15112 (N_15112,N_12496,N_13990);
and U15113 (N_15113,N_14925,N_12176);
nand U15114 (N_15114,N_13319,N_12501);
or U15115 (N_15115,N_12461,N_12324);
nor U15116 (N_15116,N_14303,N_12262);
nor U15117 (N_15117,N_12973,N_14965);
and U15118 (N_15118,N_14227,N_12807);
or U15119 (N_15119,N_14706,N_13431);
nor U15120 (N_15120,N_14738,N_12946);
nor U15121 (N_15121,N_12996,N_14108);
nor U15122 (N_15122,N_12250,N_13441);
xor U15123 (N_15123,N_13378,N_13538);
or U15124 (N_15124,N_12445,N_14611);
nor U15125 (N_15125,N_13612,N_13484);
and U15126 (N_15126,N_13750,N_12577);
nor U15127 (N_15127,N_13062,N_13212);
nand U15128 (N_15128,N_12275,N_13500);
and U15129 (N_15129,N_13911,N_14382);
or U15130 (N_15130,N_14247,N_14707);
xnor U15131 (N_15131,N_13498,N_13782);
and U15132 (N_15132,N_13347,N_12320);
and U15133 (N_15133,N_14951,N_14292);
nand U15134 (N_15134,N_13317,N_14320);
or U15135 (N_15135,N_13278,N_14907);
and U15136 (N_15136,N_14139,N_14190);
nand U15137 (N_15137,N_14419,N_13692);
nor U15138 (N_15138,N_12796,N_14411);
nor U15139 (N_15139,N_12997,N_13799);
xor U15140 (N_15140,N_13116,N_14863);
xnor U15141 (N_15141,N_13688,N_12485);
xnor U15142 (N_15142,N_12972,N_13478);
nor U15143 (N_15143,N_12286,N_14749);
and U15144 (N_15144,N_13221,N_12774);
and U15145 (N_15145,N_12953,N_12553);
nor U15146 (N_15146,N_14819,N_13956);
xor U15147 (N_15147,N_13726,N_13112);
nor U15148 (N_15148,N_12102,N_13171);
and U15149 (N_15149,N_13950,N_13234);
and U15150 (N_15150,N_14369,N_14592);
nor U15151 (N_15151,N_12556,N_13295);
and U15152 (N_15152,N_12411,N_14163);
and U15153 (N_15153,N_13371,N_12602);
nand U15154 (N_15154,N_12971,N_14480);
nor U15155 (N_15155,N_13671,N_12886);
xor U15156 (N_15156,N_14137,N_12723);
and U15157 (N_15157,N_14994,N_13125);
nor U15158 (N_15158,N_12127,N_13453);
nor U15159 (N_15159,N_12990,N_13965);
nor U15160 (N_15160,N_12799,N_14099);
and U15161 (N_15161,N_13951,N_14180);
or U15162 (N_15162,N_14103,N_14467);
nand U15163 (N_15163,N_14395,N_12056);
nor U15164 (N_15164,N_13669,N_14089);
and U15165 (N_15165,N_12331,N_12509);
or U15166 (N_15166,N_14846,N_14322);
and U15167 (N_15167,N_13293,N_12277);
xor U15168 (N_15168,N_13473,N_14542);
nor U15169 (N_15169,N_13229,N_14776);
nor U15170 (N_15170,N_14406,N_14889);
or U15171 (N_15171,N_12835,N_13971);
or U15172 (N_15172,N_13496,N_14058);
and U15173 (N_15173,N_14772,N_13479);
or U15174 (N_15174,N_14277,N_12498);
nor U15175 (N_15175,N_13326,N_14884);
or U15176 (N_15176,N_13379,N_12689);
nor U15177 (N_15177,N_12021,N_14635);
or U15178 (N_15178,N_13751,N_12863);
and U15179 (N_15179,N_14685,N_12097);
and U15180 (N_15180,N_13232,N_12829);
xor U15181 (N_15181,N_13399,N_14495);
nor U15182 (N_15182,N_13226,N_12902);
nor U15183 (N_15183,N_12370,N_12066);
or U15184 (N_15184,N_13341,N_14861);
and U15185 (N_15185,N_12692,N_14189);
or U15186 (N_15186,N_12920,N_14426);
or U15187 (N_15187,N_12706,N_14555);
and U15188 (N_15188,N_13625,N_13792);
nand U15189 (N_15189,N_12182,N_12316);
nand U15190 (N_15190,N_14668,N_12900);
or U15191 (N_15191,N_12348,N_12962);
nor U15192 (N_15192,N_14252,N_14518);
nand U15193 (N_15193,N_13497,N_14468);
and U15194 (N_15194,N_14804,N_14624);
and U15195 (N_15195,N_14024,N_12952);
or U15196 (N_15196,N_13010,N_13312);
or U15197 (N_15197,N_14902,N_14830);
and U15198 (N_15198,N_12598,N_13027);
nor U15199 (N_15199,N_14517,N_14877);
and U15200 (N_15200,N_13539,N_12836);
nor U15201 (N_15201,N_14387,N_14438);
nor U15202 (N_15202,N_12614,N_13178);
and U15203 (N_15203,N_14044,N_14654);
and U15204 (N_15204,N_14283,N_14110);
nand U15205 (N_15205,N_12789,N_14754);
nor U15206 (N_15206,N_14485,N_12529);
nand U15207 (N_15207,N_12593,N_14378);
and U15208 (N_15208,N_13734,N_13845);
nor U15209 (N_15209,N_12711,N_13404);
or U15210 (N_15210,N_12516,N_12290);
nand U15211 (N_15211,N_12371,N_13676);
or U15212 (N_15212,N_13198,N_14558);
nand U15213 (N_15213,N_13635,N_14373);
or U15214 (N_15214,N_14852,N_13569);
or U15215 (N_15215,N_14404,N_14847);
nand U15216 (N_15216,N_14497,N_12899);
or U15217 (N_15217,N_13793,N_12263);
and U15218 (N_15218,N_12232,N_14899);
nor U15219 (N_15219,N_12327,N_12417);
nand U15220 (N_15220,N_13250,N_14523);
and U15221 (N_15221,N_13652,N_13947);
or U15222 (N_15222,N_14444,N_12718);
and U15223 (N_15223,N_12009,N_14549);
and U15224 (N_15224,N_14594,N_13704);
nor U15225 (N_15225,N_12185,N_12631);
nand U15226 (N_15226,N_13060,N_13637);
and U15227 (N_15227,N_12680,N_14729);
nor U15228 (N_15228,N_13418,N_13813);
and U15229 (N_15229,N_14000,N_13315);
or U15230 (N_15230,N_12430,N_13053);
or U15231 (N_15231,N_12770,N_12568);
nand U15232 (N_15232,N_12089,N_13654);
nor U15233 (N_15233,N_14077,N_13309);
nand U15234 (N_15234,N_13520,N_14559);
or U15235 (N_15235,N_14129,N_12744);
and U15236 (N_15236,N_14392,N_14422);
xor U15237 (N_15237,N_12439,N_13576);
nor U15238 (N_15238,N_14878,N_12574);
nand U15239 (N_15239,N_12080,N_13931);
nor U15240 (N_15240,N_13282,N_14046);
nand U15241 (N_15241,N_13882,N_13096);
nor U15242 (N_15242,N_12898,N_12463);
and U15243 (N_15243,N_14451,N_12607);
or U15244 (N_15244,N_12840,N_14843);
nand U15245 (N_15245,N_14642,N_14431);
nor U15246 (N_15246,N_13725,N_13223);
nor U15247 (N_15247,N_13744,N_14756);
and U15248 (N_15248,N_13626,N_14747);
nor U15249 (N_15249,N_12304,N_14203);
and U15250 (N_15250,N_14837,N_14418);
nor U15251 (N_15251,N_12609,N_12563);
or U15252 (N_15252,N_13553,N_12270);
and U15253 (N_15253,N_14505,N_12685);
or U15254 (N_15254,N_14927,N_12674);
or U15255 (N_15255,N_12995,N_12002);
nand U15256 (N_15256,N_12606,N_14181);
nand U15257 (N_15257,N_13083,N_14834);
or U15258 (N_15258,N_12280,N_12847);
nand U15259 (N_15259,N_13833,N_12714);
nor U15260 (N_15260,N_13408,N_14101);
and U15261 (N_15261,N_12345,N_12012);
and U15262 (N_15262,N_12927,N_12538);
or U15263 (N_15263,N_13237,N_12551);
xnor U15264 (N_15264,N_14401,N_14115);
xor U15265 (N_15265,N_12850,N_14606);
or U15266 (N_15266,N_12964,N_13899);
and U15267 (N_15267,N_14097,N_12184);
nor U15268 (N_15268,N_13316,N_12095);
nor U15269 (N_15269,N_12825,N_13356);
nor U15270 (N_15270,N_14987,N_13893);
xor U15271 (N_15271,N_12346,N_12735);
and U15272 (N_15272,N_14038,N_14083);
xnor U15273 (N_15273,N_12423,N_12347);
nand U15274 (N_15274,N_13587,N_13860);
or U15275 (N_15275,N_14630,N_12699);
and U15276 (N_15276,N_14579,N_12765);
or U15277 (N_15277,N_12843,N_14019);
nand U15278 (N_15278,N_12208,N_14669);
or U15279 (N_15279,N_12006,N_13026);
or U15280 (N_15280,N_14610,N_14775);
and U15281 (N_15281,N_13998,N_14760);
and U15282 (N_15282,N_14002,N_13439);
and U15283 (N_15283,N_12435,N_14319);
and U15284 (N_15284,N_13677,N_13066);
or U15285 (N_15285,N_12851,N_14531);
nand U15286 (N_15286,N_14740,N_12895);
and U15287 (N_15287,N_12800,N_12151);
and U15288 (N_15288,N_12999,N_14457);
nand U15289 (N_15289,N_14161,N_13800);
nand U15290 (N_15290,N_12030,N_14687);
or U15291 (N_15291,N_14470,N_12554);
nor U15292 (N_15292,N_13072,N_12746);
nor U15293 (N_15293,N_14297,N_12918);
or U15294 (N_15294,N_13281,N_12414);
and U15295 (N_15295,N_12169,N_14356);
xnor U15296 (N_15296,N_12224,N_12104);
or U15297 (N_15297,N_14763,N_14570);
xor U15298 (N_15298,N_13402,N_13310);
and U15299 (N_15299,N_13209,N_12508);
or U15300 (N_15300,N_14318,N_14943);
nand U15301 (N_15301,N_13368,N_13832);
nand U15302 (N_15302,N_12955,N_14578);
and U15303 (N_15303,N_12437,N_12933);
or U15304 (N_15304,N_12237,N_13132);
or U15305 (N_15305,N_13573,N_12213);
or U15306 (N_15306,N_12358,N_14091);
or U15307 (N_15307,N_13030,N_13272);
xor U15308 (N_15308,N_14123,N_12111);
xnor U15309 (N_15309,N_14028,N_12626);
or U15310 (N_15310,N_13284,N_13297);
nor U15311 (N_15311,N_12659,N_13196);
and U15312 (N_15312,N_13103,N_13094);
nor U15313 (N_15313,N_14017,N_14638);
nor U15314 (N_15314,N_14400,N_14936);
and U15315 (N_15315,N_14674,N_13425);
nand U15316 (N_15316,N_13040,N_14814);
nor U15317 (N_15317,N_13546,N_14170);
nor U15318 (N_15318,N_13583,N_13119);
nand U15319 (N_15319,N_13976,N_14246);
and U15320 (N_15320,N_13959,N_12289);
and U15321 (N_15321,N_13055,N_12885);
or U15322 (N_15322,N_12078,N_12987);
or U15323 (N_15323,N_12645,N_14472);
nor U15324 (N_15324,N_14636,N_12291);
or U15325 (N_15325,N_14095,N_13507);
nor U15326 (N_15326,N_13896,N_14589);
nor U15327 (N_15327,N_13476,N_14164);
nand U15328 (N_15328,N_12809,N_13830);
or U15329 (N_15329,N_14151,N_12732);
xor U15330 (N_15330,N_13149,N_14969);
and U15331 (N_15331,N_14239,N_14420);
nand U15332 (N_15332,N_13088,N_13274);
and U15333 (N_15333,N_12585,N_12451);
or U15334 (N_15334,N_14234,N_12623);
and U15335 (N_15335,N_13011,N_12937);
nor U15336 (N_15336,N_13445,N_12644);
and U15337 (N_15337,N_12785,N_13376);
and U15338 (N_15338,N_13906,N_12688);
xor U15339 (N_15339,N_12130,N_14285);
nor U15340 (N_15340,N_14715,N_13017);
or U15341 (N_15341,N_13005,N_13280);
nand U15342 (N_15342,N_14782,N_14547);
nand U15343 (N_15343,N_14713,N_12019);
and U15344 (N_15344,N_12088,N_13268);
nor U15345 (N_15345,N_13201,N_14703);
nand U15346 (N_15346,N_13164,N_14996);
nand U15347 (N_15347,N_14326,N_13643);
or U15348 (N_15348,N_13869,N_13106);
xnor U15349 (N_15349,N_12513,N_14662);
and U15350 (N_15350,N_12118,N_13336);
or U15351 (N_15351,N_14460,N_14810);
nand U15352 (N_15352,N_14348,N_14025);
xor U15353 (N_15353,N_13262,N_14509);
and U15354 (N_15354,N_13449,N_12373);
or U15355 (N_15355,N_14551,N_13924);
or U15356 (N_15356,N_14376,N_14898);
and U15357 (N_15357,N_13759,N_14096);
and U15358 (N_15358,N_12369,N_14801);
nor U15359 (N_15359,N_14036,N_13414);
nor U15360 (N_15360,N_14682,N_13602);
and U15361 (N_15361,N_14539,N_13464);
nand U15362 (N_15362,N_14204,N_14323);
or U15363 (N_15363,N_12293,N_12005);
nand U15364 (N_15364,N_13985,N_13968);
nand U15365 (N_15365,N_12632,N_13458);
nor U15366 (N_15366,N_14245,N_13279);
or U15367 (N_15367,N_12068,N_13821);
xor U15368 (N_15368,N_13708,N_14043);
nor U15369 (N_15369,N_12427,N_12093);
or U15370 (N_15370,N_13429,N_14835);
nand U15371 (N_15371,N_12945,N_13645);
nor U15372 (N_15372,N_13735,N_14689);
or U15373 (N_15373,N_13121,N_12702);
nor U15374 (N_15374,N_14655,N_13475);
or U15375 (N_15375,N_12242,N_13486);
and U15376 (N_15376,N_14466,N_12569);
or U15377 (N_15377,N_14120,N_12203);
nor U15378 (N_15378,N_14781,N_14868);
nor U15379 (N_15379,N_14327,N_13621);
and U15380 (N_15380,N_14060,N_14619);
nor U15381 (N_15381,N_12797,N_14106);
nand U15382 (N_15382,N_14603,N_13655);
and U15383 (N_15383,N_14477,N_13999);
nand U15384 (N_15384,N_13518,N_13885);
and U15385 (N_15385,N_13542,N_13286);
and U15386 (N_15386,N_13974,N_13059);
or U15387 (N_15387,N_12247,N_12708);
nor U15388 (N_15388,N_14399,N_12868);
nor U15389 (N_15389,N_13217,N_12460);
nor U15390 (N_15390,N_12818,N_13624);
or U15391 (N_15391,N_12500,N_12806);
nand U15392 (N_15392,N_14514,N_12199);
nand U15393 (N_15393,N_13276,N_14939);
nand U15394 (N_15394,N_14072,N_13977);
nand U15395 (N_15395,N_14691,N_13243);
xnor U15396 (N_15396,N_13829,N_14014);
nor U15397 (N_15397,N_13195,N_13737);
nor U15398 (N_15398,N_12064,N_14521);
or U15399 (N_15399,N_12288,N_12709);
nand U15400 (N_15400,N_14366,N_14312);
or U15401 (N_15401,N_13713,N_12236);
nor U15402 (N_15402,N_13109,N_12742);
nand U15403 (N_15403,N_13031,N_12517);
nand U15404 (N_15404,N_12312,N_13663);
or U15405 (N_15405,N_12812,N_12488);
or U15406 (N_15406,N_14187,N_12808);
and U15407 (N_15407,N_14704,N_13041);
or U15408 (N_15408,N_14815,N_13787);
or U15409 (N_15409,N_13018,N_12070);
and U15410 (N_15410,N_13712,N_14694);
nor U15411 (N_15411,N_13185,N_14891);
and U15412 (N_15412,N_14803,N_14117);
nand U15413 (N_15413,N_14922,N_13002);
nand U15414 (N_15414,N_14063,N_12911);
and U15415 (N_15415,N_13721,N_14183);
xor U15416 (N_15416,N_14914,N_14342);
and U15417 (N_15417,N_14344,N_13920);
and U15418 (N_15418,N_14228,N_14908);
nand U15419 (N_15419,N_13930,N_12261);
nor U15420 (N_15420,N_12399,N_12368);
xor U15421 (N_15421,N_13334,N_14769);
nor U15422 (N_15422,N_13870,N_13323);
xnor U15423 (N_15423,N_14450,N_13079);
nor U15424 (N_15424,N_12073,N_13170);
and U15425 (N_15425,N_13775,N_14136);
or U15426 (N_15426,N_13137,N_14800);
xor U15427 (N_15427,N_14127,N_12693);
and U15428 (N_15428,N_12595,N_12940);
nand U15429 (N_15429,N_12099,N_12781);
and U15430 (N_15430,N_12573,N_13390);
nand U15431 (N_15431,N_14933,N_12136);
or U15432 (N_15432,N_14263,N_12724);
nor U15433 (N_15433,N_14384,N_13501);
or U15434 (N_15434,N_13599,N_12094);
nor U15435 (N_15435,N_12310,N_13093);
or U15436 (N_15436,N_14684,N_12342);
or U15437 (N_15437,N_13740,N_14459);
or U15438 (N_15438,N_13955,N_14338);
and U15439 (N_15439,N_12533,N_13267);
and U15440 (N_15440,N_12067,N_14545);
nand U15441 (N_15441,N_12337,N_13736);
xor U15442 (N_15442,N_13159,N_12542);
or U15443 (N_15443,N_12518,N_13204);
nand U15444 (N_15444,N_13398,N_14313);
and U15445 (N_15445,N_12357,N_14573);
and U15446 (N_15446,N_14371,N_14930);
nor U15447 (N_15447,N_12846,N_14009);
or U15448 (N_15448,N_12321,N_12673);
or U15449 (N_15449,N_13642,N_13598);
and U15450 (N_15450,N_13898,N_14278);
or U15451 (N_15451,N_12650,N_13091);
xnor U15452 (N_15452,N_13585,N_14572);
or U15453 (N_15453,N_12323,N_12157);
nor U15454 (N_15454,N_13086,N_12256);
nand U15455 (N_15455,N_12612,N_13176);
or U15456 (N_15456,N_14945,N_13988);
and U15457 (N_15457,N_12069,N_14725);
or U15458 (N_15458,N_13586,N_12497);
or U15459 (N_15459,N_14047,N_14308);
or U15460 (N_15460,N_14116,N_14496);
nand U15461 (N_15461,N_13873,N_13304);
nor U15462 (N_15462,N_14162,N_12436);
and U15463 (N_15463,N_14774,N_12570);
and U15464 (N_15464,N_13761,N_13480);
and U15465 (N_15465,N_12487,N_13995);
nor U15466 (N_15466,N_13241,N_13056);
and U15467 (N_15467,N_12663,N_13722);
or U15468 (N_15468,N_14100,N_12837);
xor U15469 (N_15469,N_14620,N_12384);
xnor U15470 (N_15470,N_13224,N_13756);
or U15471 (N_15471,N_13469,N_13842);
and U15472 (N_15472,N_13194,N_13477);
xnor U15473 (N_15473,N_13820,N_12753);
or U15474 (N_15474,N_13021,N_13245);
or U15475 (N_15475,N_13597,N_13807);
nor U15476 (N_15476,N_13742,N_12040);
or U15477 (N_15477,N_12113,N_14960);
nand U15478 (N_15478,N_12378,N_13747);
nor U15479 (N_15479,N_12939,N_14561);
nand U15480 (N_15480,N_13711,N_14434);
or U15481 (N_15481,N_13314,N_14090);
nor U15482 (N_15482,N_13487,N_12383);
or U15483 (N_15483,N_12020,N_12172);
and U15484 (N_15484,N_13848,N_14881);
nand U15485 (N_15485,N_14895,N_14793);
or U15486 (N_15486,N_13351,N_14331);
and U15487 (N_15487,N_13650,N_14981);
and U15488 (N_15488,N_13894,N_12737);
and U15489 (N_15489,N_12216,N_13292);
and U15490 (N_15490,N_13242,N_13269);
xnor U15491 (N_15491,N_12502,N_14500);
or U15492 (N_15492,N_13993,N_12311);
nor U15493 (N_15493,N_14499,N_14256);
and U15494 (N_15494,N_14385,N_13815);
nor U15495 (N_15495,N_14458,N_14946);
nor U15496 (N_15496,N_13000,N_13622);
xor U15497 (N_15497,N_13329,N_13472);
and U15498 (N_15498,N_14985,N_14753);
xor U15499 (N_15499,N_14932,N_12985);
or U15500 (N_15500,N_14757,N_14109);
and U15501 (N_15501,N_14616,N_12052);
nand U15502 (N_15502,N_14836,N_13192);
nand U15503 (N_15503,N_14690,N_12238);
or U15504 (N_15504,N_13206,N_14944);
and U15505 (N_15505,N_14104,N_13972);
or U15506 (N_15506,N_13778,N_12697);
or U15507 (N_15507,N_14380,N_12119);
and U15508 (N_15508,N_13424,N_12771);
or U15509 (N_15509,N_12634,N_12394);
and U15510 (N_15510,N_14295,N_14209);
nor U15511 (N_15511,N_13270,N_12483);
nor U15512 (N_15512,N_12074,N_13337);
and U15513 (N_15513,N_13389,N_13181);
and U15514 (N_15514,N_14507,N_12171);
or U15515 (N_15515,N_14525,N_14731);
nand U15516 (N_15516,N_13413,N_14848);
xor U15517 (N_15517,N_12893,N_14207);
nand U15518 (N_15518,N_13890,N_13646);
nand U15519 (N_15519,N_13207,N_14343);
and U15520 (N_15520,N_12221,N_13554);
nand U15521 (N_15521,N_13437,N_14673);
and U15522 (N_15522,N_14968,N_14436);
and U15523 (N_15523,N_14242,N_13174);
xnor U15524 (N_15524,N_12228,N_12936);
nor U15525 (N_15525,N_13303,N_12532);
nand U15526 (N_15526,N_14031,N_14440);
xnor U15527 (N_15527,N_12967,N_12860);
and U15528 (N_15528,N_12076,N_12421);
nor U15529 (N_15529,N_13455,N_14449);
or U15530 (N_15530,N_13611,N_14258);
nor U15531 (N_15531,N_13948,N_12950);
or U15532 (N_15532,N_12656,N_13190);
xnor U15533 (N_15533,N_12234,N_12731);
nor U15534 (N_15534,N_14791,N_13104);
or U15535 (N_15535,N_14330,N_13914);
xor U15536 (N_15536,N_12811,N_12993);
and U15537 (N_15537,N_12528,N_12670);
nor U15538 (N_15538,N_12974,N_13962);
or U15539 (N_15539,N_14955,N_14931);
nand U15540 (N_15540,N_14425,N_14688);
or U15541 (N_15541,N_14219,N_13460);
nand U15542 (N_15542,N_14529,N_14569);
or U15543 (N_15543,N_13916,N_13210);
nor U15544 (N_15544,N_12443,N_12214);
and U15545 (N_15545,N_12315,N_13366);
or U15546 (N_15546,N_13023,N_14332);
or U15547 (N_15547,N_13098,N_13511);
nor U15548 (N_15548,N_13717,N_13981);
and U15549 (N_15549,N_12923,N_12302);
nand U15550 (N_15550,N_14055,N_12385);
and U15551 (N_15551,N_14264,N_14954);
or U15552 (N_15552,N_13570,N_14512);
nand U15553 (N_15553,N_13289,N_14705);
nor U15554 (N_15554,N_14273,N_13416);
nand U15555 (N_15555,N_13462,N_14541);
nor U15556 (N_15556,N_13384,N_14006);
and U15557 (N_15557,N_12629,N_14563);
and U15558 (N_15558,N_13189,N_13222);
nor U15559 (N_15559,N_14625,N_13805);
nor U15560 (N_15560,N_14210,N_13047);
nand U15561 (N_15561,N_12643,N_13372);
nor U15562 (N_15562,N_14494,N_12174);
nor U15563 (N_15563,N_13836,N_14957);
nand U15564 (N_15564,N_12531,N_13360);
and U15565 (N_15565,N_13730,N_12166);
nand U15566 (N_15566,N_14953,N_14990);
and U15567 (N_15567,N_13105,N_14410);
and U15568 (N_15568,N_13794,N_14347);
or U15569 (N_15569,N_12832,N_12332);
and U15570 (N_15570,N_12148,N_12292);
and U15571 (N_15571,N_12026,N_13929);
and U15572 (N_15572,N_14172,N_13328);
nor U15573 (N_15573,N_13783,N_12764);
xnor U15574 (N_15574,N_12319,N_12202);
nand U15575 (N_15575,N_12890,N_12010);
nor U15576 (N_15576,N_12654,N_12980);
nand U15577 (N_15577,N_13754,N_14243);
nor U15578 (N_15578,N_14700,N_13773);
nor U15579 (N_15579,N_12854,N_12701);
and U15580 (N_15580,N_14702,N_13239);
and U15581 (N_15581,N_13809,N_12160);
or U15582 (N_15582,N_14150,N_14309);
or U15583 (N_15583,N_14598,N_13917);
nor U15584 (N_15584,N_14762,N_13135);
or U15585 (N_15585,N_13175,N_12273);
nor U15586 (N_15586,N_14719,N_12562);
nor U15587 (N_15587,N_12083,N_13296);
nand U15588 (N_15588,N_13670,N_12027);
or U15589 (N_15589,N_13253,N_13330);
xnor U15590 (N_15590,N_13186,N_14200);
or U15591 (N_15591,N_12804,N_12492);
nor U15592 (N_15592,N_13589,N_14405);
or U15593 (N_15593,N_14306,N_13780);
and U15594 (N_15594,N_12284,N_12908);
and U15595 (N_15595,N_13065,N_14298);
nor U15596 (N_15596,N_12845,N_14304);
xor U15597 (N_15597,N_12416,N_12888);
nand U15598 (N_15598,N_13377,N_12493);
and U15599 (N_15599,N_13679,N_12550);
nand U15600 (N_15600,N_12354,N_14317);
and U15601 (N_15601,N_13305,N_13935);
nor U15602 (N_15602,N_13338,N_14888);
nor U15603 (N_15603,N_13246,N_12722);
and U15604 (N_15604,N_13524,N_14676);
nand U15605 (N_15605,N_12527,N_14515);
and U15606 (N_15606,N_13849,N_12072);
and U15607 (N_15607,N_13534,N_14926);
nand U15608 (N_15608,N_14354,N_13205);
nand U15609 (N_15609,N_12328,N_14244);
or U15610 (N_15610,N_12769,N_14238);
or U15611 (N_15611,N_14808,N_13941);
xor U15612 (N_15612,N_13665,N_12106);
or U15613 (N_15613,N_14328,N_13651);
or U15614 (N_15614,N_14911,N_13871);
nor U15615 (N_15615,N_13866,N_12376);
nor U15616 (N_15616,N_13666,N_13502);
and U15617 (N_15617,N_12060,N_14958);
or U15618 (N_15618,N_14126,N_12398);
or U15619 (N_15619,N_14949,N_12455);
and U15620 (N_15620,N_14634,N_12857);
or U15621 (N_15621,N_14748,N_13126);
nand U15622 (N_15622,N_14146,N_12963);
nand U15623 (N_15623,N_13036,N_12669);
xnor U15624 (N_15624,N_12037,N_14742);
nor U15625 (N_15625,N_14093,N_13447);
nand U15626 (N_15626,N_13016,N_13275);
and U15627 (N_15627,N_13880,N_13179);
or U15628 (N_15628,N_13827,N_13966);
and U15629 (N_15629,N_14053,N_14482);
or U15630 (N_15630,N_13331,N_12719);
and U15631 (N_15631,N_12791,N_14580);
nor U15632 (N_15632,N_13373,N_13162);
nor U15633 (N_15633,N_12446,N_12728);
nor U15634 (N_15634,N_12684,N_14827);
or U15635 (N_15635,N_12035,N_14250);
nor U15636 (N_15636,N_12390,N_14272);
nor U15637 (N_15637,N_13661,N_14621);
or U15638 (N_15638,N_13919,N_14461);
or U15639 (N_15639,N_12274,N_12143);
or U15640 (N_15640,N_12849,N_14920);
and U15641 (N_15641,N_12264,N_14718);
nor U15642 (N_15642,N_14959,N_13320);
nor U15643 (N_15643,N_12395,N_14595);
nand U15644 (N_15644,N_12474,N_12874);
nor U15645 (N_15645,N_12565,N_14838);
nand U15646 (N_15646,N_13878,N_14066);
xor U15647 (N_15647,N_14184,N_14553);
xnor U15648 (N_15648,N_12181,N_14081);
xor U15649 (N_15649,N_12658,N_14288);
or U15650 (N_15650,N_14140,N_14374);
and U15651 (N_15651,N_12298,N_12449);
nand U15652 (N_15652,N_12560,N_13219);
and U15653 (N_15653,N_13193,N_14941);
or U15654 (N_15654,N_12341,N_12330);
nor U15655 (N_15655,N_14156,N_12008);
nand U15656 (N_15656,N_13240,N_13367);
nand U15657 (N_15657,N_14255,N_14565);
and U15658 (N_15658,N_12220,N_14266);
or U15659 (N_15659,N_14644,N_12218);
xor U15660 (N_15660,N_14362,N_13607);
nor U15661 (N_15661,N_12704,N_12472);
and U15662 (N_15662,N_12981,N_13515);
nand U15663 (N_15663,N_14453,N_14628);
and U15664 (N_15664,N_14078,N_14904);
nor U15665 (N_15665,N_13523,N_13509);
and U15666 (N_15666,N_13471,N_12826);
or U15667 (N_15667,N_12738,N_13134);
and U15668 (N_15668,N_14839,N_12434);
and U15669 (N_15669,N_12473,N_14730);
or U15670 (N_15670,N_13427,N_14284);
or U15671 (N_15671,N_12459,N_14289);
and U15672 (N_15672,N_14335,N_14122);
or U15673 (N_15673,N_12407,N_14586);
and U15674 (N_15674,N_12834,N_14132);
nand U15675 (N_15675,N_13892,N_13442);
nand U15676 (N_15676,N_13388,N_13403);
or U15677 (N_15677,N_13872,N_14692);
nand U15678 (N_15678,N_12081,N_14604);
xor U15679 (N_15679,N_13024,N_12740);
and U15680 (N_15680,N_12230,N_12161);
nand U15681 (N_15681,N_14386,N_12029);
and U15682 (N_15682,N_13913,N_12642);
nand U15683 (N_15683,N_12882,N_14314);
nor U15684 (N_15684,N_13806,N_14381);
and U15685 (N_15685,N_12480,N_14217);
and U15686 (N_15686,N_13864,N_12988);
and U15687 (N_15687,N_12599,N_14587);
nor U15688 (N_15688,N_12803,N_13853);
nand U15689 (N_15689,N_13618,N_14812);
or U15690 (N_15690,N_12576,N_13987);
nor U15691 (N_15691,N_13038,N_13760);
nor U15692 (N_15692,N_13139,N_12676);
or U15693 (N_15693,N_13967,N_13693);
nand U15694 (N_15694,N_14745,N_13879);
and U15695 (N_15695,N_12620,N_13746);
or U15696 (N_15696,N_13703,N_13236);
or U15697 (N_15697,N_12559,N_13601);
or U15698 (N_15698,N_14648,N_13680);
or U15699 (N_15699,N_13166,N_14918);
or U15700 (N_15700,N_13513,N_12672);
xnor U15701 (N_15701,N_14882,N_14057);
nor U15702 (N_15702,N_12283,N_12581);
nor U15703 (N_15703,N_13838,N_14346);
and U15704 (N_15704,N_14510,N_12255);
nand U15705 (N_15705,N_13290,N_14564);
nor U15706 (N_15706,N_13548,N_14806);
nor U15707 (N_15707,N_12969,N_13172);
xor U15708 (N_15708,N_14004,N_12821);
and U15709 (N_15709,N_12521,N_14853);
or U15710 (N_15710,N_13659,N_13037);
nor U15711 (N_15711,N_12831,N_12252);
nor U15712 (N_15712,N_12087,N_12314);
nand U15713 (N_15713,N_13200,N_13343);
and U15714 (N_15714,N_12226,N_13225);
nor U15715 (N_15715,N_13167,N_14615);
xnor U15716 (N_15716,N_13709,N_13374);
or U15717 (N_15717,N_13249,N_12720);
nor U15718 (N_15718,N_13235,N_14240);
nand U15719 (N_15719,N_13123,N_13938);
and U15720 (N_15720,N_12909,N_13077);
nor U15721 (N_15721,N_12405,N_14223);
or U15722 (N_15722,N_14670,N_13949);
or U15723 (N_15723,N_13578,N_13900);
or U15724 (N_15724,N_12432,N_12536);
xor U15725 (N_15725,N_14613,N_13946);
or U15726 (N_15726,N_14741,N_13157);
nand U15727 (N_15727,N_14982,N_13795);
nand U15728 (N_15728,N_12217,N_13996);
nor U15729 (N_15729,N_13574,N_13215);
nor U15730 (N_15730,N_12050,N_14999);
or U15731 (N_15731,N_12715,N_13396);
and U15732 (N_15732,N_13169,N_13851);
nor U15733 (N_15733,N_12142,N_13432);
nand U15734 (N_15734,N_13007,N_12869);
nand U15735 (N_15735,N_14260,N_13092);
and U15736 (N_15736,N_14113,N_14397);
or U15737 (N_15737,N_13521,N_13859);
and U15738 (N_15738,N_12100,N_12784);
nand U15739 (N_15739,N_12668,N_12992);
nand U15740 (N_15740,N_13633,N_12098);
nand U15741 (N_15741,N_13359,N_12947);
nor U15742 (N_15742,N_13020,N_13506);
or U15743 (N_15743,N_12647,N_13889);
and U15744 (N_15744,N_14862,N_14402);
and U15745 (N_15745,N_13577,N_14464);
or U15746 (N_15746,N_12360,N_12317);
and U15747 (N_15747,N_12586,N_14412);
or U15748 (N_15748,N_13781,N_13342);
nand U15749 (N_15749,N_14746,N_14048);
nor U15750 (N_15750,N_13888,N_13954);
xor U15751 (N_15751,N_13348,N_12269);
and U15752 (N_15752,N_14535,N_12839);
nand U15753 (N_15753,N_12392,N_13579);
or U15754 (N_15754,N_14964,N_13461);
or U15755 (N_15755,N_12032,N_13620);
or U15756 (N_15756,N_14721,N_13748);
nand U15757 (N_15757,N_12031,N_12022);
nor U15758 (N_15758,N_14216,N_12418);
xnor U15759 (N_15759,N_13258,N_12075);
or U15760 (N_15760,N_12420,N_14575);
or U15761 (N_15761,N_13875,N_12096);
nand U15762 (N_15762,N_13014,N_12308);
nor U15763 (N_15763,N_12057,N_12910);
or U15764 (N_15764,N_14588,N_14259);
nor U15765 (N_15765,N_13915,N_14241);
or U15766 (N_15766,N_12755,N_12705);
nor U15767 (N_15767,N_14678,N_13543);
nand U15768 (N_15768,N_14526,N_14049);
xor U15769 (N_15769,N_13050,N_14732);
xor U15770 (N_15770,N_13154,N_12490);
and U15771 (N_15771,N_12079,N_13333);
nand U15772 (N_15772,N_12281,N_13214);
or U15773 (N_15773,N_14784,N_12380);
and U15774 (N_15774,N_14583,N_14639);
nand U15775 (N_15775,N_12641,N_13454);
nor U15776 (N_15776,N_13682,N_12925);
and U15777 (N_15777,N_13084,N_14398);
and U15778 (N_15778,N_13153,N_14321);
nor U15779 (N_15779,N_14915,N_14428);
and U15780 (N_15780,N_12747,N_14267);
nand U15781 (N_15781,N_14865,N_12520);
or U15782 (N_15782,N_13979,N_13433);
nor U15783 (N_15783,N_13435,N_12892);
nor U15784 (N_15784,N_12219,N_12381);
xor U15785 (N_15785,N_12164,N_12594);
nor U15786 (N_15786,N_14723,N_13208);
xor U15787 (N_15787,N_14873,N_14653);
nor U15788 (N_15788,N_13385,N_13686);
or U15789 (N_15789,N_12805,N_12188);
nor U15790 (N_15790,N_12003,N_13980);
xnor U15791 (N_15791,N_12646,N_12245);
nor U15792 (N_15792,N_14728,N_12244);
and U15793 (N_15793,N_13004,N_12539);
or U15794 (N_15794,N_13165,N_14826);
xnor U15795 (N_15795,N_14767,N_14649);
or U15796 (N_15796,N_13228,N_12484);
or U15797 (N_15797,N_12567,N_14360);
or U15798 (N_15798,N_13075,N_13550);
and U15799 (N_15799,N_13512,N_14855);
and U15800 (N_15800,N_12547,N_12223);
xor U15801 (N_15801,N_14027,N_12864);
nor U15802 (N_15802,N_14152,N_14271);
or U15803 (N_15803,N_14608,N_13551);
and U15804 (N_15804,N_12272,N_12522);
nand U15805 (N_15805,N_14339,N_13816);
or U15806 (N_15806,N_14443,N_14423);
xnor U15807 (N_15807,N_13685,N_13146);
xnor U15808 (N_15808,N_14350,N_12733);
or U15809 (N_15809,N_14766,N_14432);
nor U15810 (N_15810,N_14537,N_14540);
and U15811 (N_15811,N_13393,N_12975);
or U15812 (N_15812,N_13531,N_14851);
nand U15813 (N_15813,N_13264,N_14858);
nand U15814 (N_15814,N_12051,N_14928);
and U15815 (N_15815,N_12779,N_13610);
nor U15816 (N_15816,N_13961,N_14854);
or U15817 (N_15817,N_12926,N_14887);
nor U15818 (N_15818,N_13203,N_13745);
nor U15819 (N_15819,N_14390,N_13008);
nand U15820 (N_15820,N_14059,N_14768);
or U15821 (N_15821,N_13558,N_12017);
nand U15822 (N_15822,N_12433,N_12422);
nor U15823 (N_15823,N_13428,N_14221);
and U15824 (N_15824,N_12034,N_13064);
or U15825 (N_15825,N_14617,N_14977);
nor U15826 (N_15826,N_14978,N_13715);
nor U15827 (N_15827,N_12505,N_12651);
nand U15828 (N_15828,N_13723,N_12904);
nor U15829 (N_15829,N_12458,N_13406);
xnor U15830 (N_15830,N_12555,N_14192);
nor U15831 (N_15831,N_12428,N_14388);
or U15832 (N_15832,N_13101,N_12128);
and U15833 (N_15833,N_13964,N_13335);
or U15834 (N_15834,N_14224,N_13277);
nand U15835 (N_15835,N_14157,N_14491);
and U15836 (N_15836,N_13273,N_13673);
xor U15837 (N_15837,N_14844,N_14212);
or U15838 (N_15838,N_12178,N_13248);
nor U15839 (N_15839,N_12396,N_14208);
nand U15840 (N_15840,N_12700,N_12540);
nand U15841 (N_15841,N_13032,N_12457);
or U15842 (N_15842,N_12625,N_13989);
nor U15843 (N_15843,N_14056,N_13230);
nand U15844 (N_15844,N_13354,N_13690);
nand U15845 (N_15845,N_12571,N_12410);
nor U15846 (N_15846,N_14403,N_12822);
nand U15847 (N_15847,N_13797,N_13346);
or U15848 (N_15848,N_12334,N_12884);
or U15849 (N_15849,N_12603,N_12425);
nand U15850 (N_15850,N_13922,N_13095);
and U15851 (N_15851,N_12287,N_12870);
and U15852 (N_15852,N_13739,N_14396);
nor U15853 (N_15853,N_12303,N_14909);
xor U15854 (N_15854,N_13353,N_12730);
xnor U15855 (N_15855,N_13352,N_13557);
or U15856 (N_15856,N_13465,N_12678);
nand U15857 (N_15857,N_12476,N_13142);
and U15858 (N_15858,N_13928,N_12965);
or U15859 (N_15859,N_14294,N_12611);
or U15860 (N_15860,N_12545,N_14478);
or U15861 (N_15861,N_12943,N_12653);
nor U15862 (N_15862,N_13881,N_12322);
nand U15863 (N_15863,N_12896,N_12830);
nor U15864 (N_15864,N_12038,N_14370);
xor U15865 (N_15865,N_13188,N_12638);
nand U15866 (N_15866,N_14998,N_14903);
or U15867 (N_15867,N_13127,N_12170);
or U15868 (N_15868,N_14391,N_12149);
nand U15869 (N_15869,N_12941,N_13265);
nand U15870 (N_15870,N_12454,N_12023);
or U15871 (N_15871,N_14084,N_13182);
nor U15872 (N_15872,N_12156,N_14859);
nor U15873 (N_15873,N_13308,N_12352);
nand U15874 (N_15874,N_13369,N_14897);
or U15875 (N_15875,N_12786,N_14566);
nand U15876 (N_15876,N_14661,N_13753);
and U15877 (N_15877,N_14351,N_14337);
xor U15878 (N_15878,N_12758,N_13908);
and U15879 (N_15879,N_12844,N_14269);
nand U15880 (N_15880,N_14734,N_13953);
or U15881 (N_15881,N_13647,N_14128);
xor U15882 (N_15882,N_14568,N_14359);
and U15883 (N_15883,N_12198,N_14765);
xor U15884 (N_15884,N_12025,N_12793);
or U15885 (N_15885,N_12124,N_13080);
nor U15886 (N_15886,N_13852,N_14824);
and U15887 (N_15887,N_13613,N_14310);
and U15888 (N_15888,N_13043,N_14811);
and U15889 (N_15889,N_12276,N_14222);
nor U15890 (N_15890,N_12353,N_12001);
and U15891 (N_15891,N_13555,N_12133);
nand U15892 (N_15892,N_12743,N_12489);
nor U15893 (N_15893,N_12552,N_13307);
and U15894 (N_15894,N_12313,N_12514);
or U15895 (N_15895,N_13288,N_14429);
nor U15896 (N_15896,N_12683,N_14574);
xnor U15897 (N_15897,N_14869,N_14874);
xor U15898 (N_15898,N_12624,N_13752);
and U15899 (N_15899,N_14974,N_12447);
and U15900 (N_15900,N_14643,N_14600);
or U15901 (N_15901,N_12364,N_12954);
and U15902 (N_15902,N_13986,N_14020);
nor U15903 (N_15903,N_13764,N_14105);
or U15904 (N_15904,N_12696,N_14735);
or U15905 (N_15905,N_14833,N_13874);
nor U15906 (N_15906,N_12138,N_12235);
and U15907 (N_15907,N_12666,N_14934);
or U15908 (N_15908,N_13233,N_13493);
and U15909 (N_15909,N_13662,N_12499);
or U15910 (N_15910,N_14991,N_14143);
and U15911 (N_15911,N_14237,N_12667);
and U15912 (N_15912,N_12741,N_12426);
or U15913 (N_15913,N_14680,N_14825);
and U15914 (N_15914,N_14196,N_12137);
nor U15915 (N_15915,N_12375,N_14134);
nor U15916 (N_15916,N_13696,N_13067);
or U15917 (N_15917,N_13593,N_12584);
nand U15918 (N_15918,N_12135,N_12389);
and U15919 (N_15919,N_14805,N_12622);
nor U15920 (N_15920,N_13846,N_13489);
and U15921 (N_15921,N_14363,N_14165);
nand U15922 (N_15922,N_14229,N_14073);
or U15923 (N_15923,N_14469,N_12865);
nand U15924 (N_15924,N_12931,N_14995);
xnor U15925 (N_15925,N_14712,N_14124);
xor U15926 (N_15926,N_12596,N_14711);
nand U15927 (N_15927,N_13009,N_12453);
and U15928 (N_15928,N_12333,N_14973);
xnor U15929 (N_15929,N_14956,N_13120);
nor U15930 (N_15930,N_14035,N_14188);
or U15931 (N_15931,N_12193,N_13311);
or U15932 (N_15932,N_14633,N_14012);
xnor U15933 (N_15933,N_12047,N_12086);
or U15934 (N_15934,N_12970,N_13504);
nand U15935 (N_15935,N_14612,N_13943);
or U15936 (N_15936,N_14679,N_12621);
nor U15937 (N_15937,N_12984,N_13028);
and U15938 (N_15938,N_13482,N_13287);
and U15939 (N_15939,N_12179,N_13463);
nor U15940 (N_15940,N_13124,N_12935);
and U15941 (N_15941,N_13467,N_13527);
and U15942 (N_15942,N_12855,N_13817);
nand U15943 (N_15943,N_13926,N_12792);
xnor U15944 (N_15944,N_14102,N_14709);
or U15945 (N_15945,N_12880,N_12326);
and U15946 (N_15946,N_12343,N_12828);
nand U15947 (N_15947,N_14970,N_14966);
nor U15948 (N_15948,N_14876,N_14357);
nand U15949 (N_15949,N_12155,N_14281);
nand U15950 (N_15950,N_13697,N_14567);
and U15951 (N_15951,N_12112,N_13657);
nor U15952 (N_15952,N_14751,N_12887);
or U15953 (N_15953,N_13173,N_12873);
or U15954 (N_15954,N_14979,N_12780);
nor U15955 (N_15955,N_12442,N_12117);
and U15956 (N_15956,N_13769,N_13344);
nor U15957 (N_15957,N_12838,N_12462);
nor U15958 (N_15958,N_14296,N_12852);
and U15959 (N_15959,N_12503,N_14665);
nand U15960 (N_15960,N_12726,N_12816);
nor U15961 (N_15961,N_13891,N_14910);
nor U15962 (N_15962,N_13045,N_12246);
nor U15963 (N_15963,N_12150,N_13044);
or U15964 (N_15964,N_13405,N_13627);
nand U15965 (N_15965,N_14785,N_13934);
and U15966 (N_15966,N_12278,N_13876);
nor U15967 (N_15967,N_12491,N_13560);
nand U15968 (N_15968,N_13803,N_12665);
xor U15969 (N_15969,N_13263,N_13012);
xor U15970 (N_15970,N_12894,N_14365);
nor U15971 (N_15971,N_12285,N_13561);
and U15972 (N_15972,N_12041,N_12848);
xor U15973 (N_15973,N_13145,N_14492);
xnor U15974 (N_15974,N_14409,N_14905);
nand U15975 (N_15975,N_14199,N_14759);
nor U15976 (N_15976,N_13660,N_13668);
nand U15977 (N_15977,N_14119,N_12015);
nor U15978 (N_15978,N_12597,N_14779);
and U15979 (N_15979,N_12374,N_14454);
or U15980 (N_15980,N_12403,N_14912);
nand U15981 (N_15981,N_13345,N_12147);
nor U15982 (N_15982,N_13636,N_12982);
or U15983 (N_15983,N_14867,N_12131);
or U15984 (N_15984,N_13978,N_13089);
xnor U15985 (N_15985,N_14214,N_14489);
nand U15986 (N_15986,N_13755,N_13868);
nand U15987 (N_15987,N_12546,N_14315);
or U15988 (N_15988,N_13254,N_12657);
xnor U15989 (N_15989,N_12675,N_12132);
nand U15990 (N_15990,N_13594,N_13687);
nand U15991 (N_15991,N_13452,N_12511);
or U15992 (N_15992,N_14230,N_14316);
nor U15993 (N_15993,N_13826,N_12871);
or U15994 (N_15994,N_14138,N_12300);
or U15995 (N_15995,N_12661,N_14487);
and U15996 (N_15996,N_13450,N_12801);
or U15997 (N_15997,N_12589,N_13070);
xor U15998 (N_15998,N_13150,N_13470);
nor U15999 (N_15999,N_13133,N_14614);
nand U16000 (N_16000,N_14758,N_12519);
nor U16001 (N_16001,N_14820,N_14724);
or U16002 (N_16002,N_12942,N_14198);
nor U16003 (N_16003,N_13698,N_13327);
nand U16004 (N_16004,N_14821,N_12209);
and U16005 (N_16005,N_12966,N_13048);
nor U16006 (N_16006,N_14530,N_14727);
and U16007 (N_16007,N_13495,N_13672);
nor U16008 (N_16008,N_14032,N_14424);
nand U16009 (N_16009,N_14447,N_14916);
nand U16010 (N_16010,N_14484,N_14186);
or U16011 (N_16011,N_13936,N_14860);
nand U16012 (N_16012,N_13419,N_14050);
and U16013 (N_16013,N_13227,N_13867);
and U16014 (N_16014,N_13332,N_14023);
nand U16015 (N_16015,N_12754,N_12196);
nor U16016 (N_16016,N_12448,N_14088);
or U16017 (N_16017,N_14546,N_14771);
nor U16018 (N_16018,N_12158,N_14976);
or U16019 (N_16019,N_13131,N_13492);
and U16020 (N_16020,N_12391,N_12431);
or U16021 (N_16021,N_12366,N_12543);
nor U16022 (N_16022,N_14696,N_12605);
and U16023 (N_16023,N_13828,N_14018);
nand U16024 (N_16024,N_12703,N_13863);
or U16025 (N_16025,N_12959,N_14148);
xnor U16026 (N_16026,N_13958,N_13061);
nor U16027 (N_16027,N_13862,N_12122);
nor U16028 (N_16028,N_14637,N_14194);
nor U16029 (N_16029,N_14177,N_13937);
or U16030 (N_16030,N_14452,N_12351);
nand U16031 (N_16031,N_13051,N_14393);
xnor U16032 (N_16032,N_13562,N_12438);
nand U16033 (N_16033,N_12109,N_14287);
or U16034 (N_16034,N_14474,N_14693);
and U16035 (N_16035,N_12192,N_14098);
nor U16036 (N_16036,N_14010,N_13944);
and U16037 (N_16037,N_13211,N_12249);
and U16038 (N_16038,N_14333,N_14627);
nand U16039 (N_16039,N_12061,N_13299);
nand U16040 (N_16040,N_13457,N_12168);
and U16041 (N_16041,N_12082,N_14845);
xnor U16042 (N_16042,N_14875,N_14717);
nor U16043 (N_16043,N_12504,N_12120);
nand U16044 (N_16044,N_12767,N_12515);
and U16045 (N_16045,N_13905,N_12429);
nand U16046 (N_16046,N_13420,N_13706);
nor U16047 (N_16047,N_13683,N_13547);
nand U16048 (N_16048,N_14141,N_12055);
nor U16049 (N_16049,N_14591,N_12761);
and U16050 (N_16050,N_14167,N_14498);
and U16051 (N_16051,N_12254,N_14788);
nor U16052 (N_16052,N_14651,N_12071);
nand U16053 (N_16053,N_13370,N_12141);
nor U16054 (N_16054,N_12525,N_13897);
and U16055 (N_16055,N_12788,N_14524);
xor U16056 (N_16056,N_14275,N_13381);
nor U16057 (N_16057,N_12877,N_12409);
nor U16058 (N_16058,N_14554,N_14892);
xor U16059 (N_16059,N_12979,N_12694);
nor U16060 (N_16060,N_12231,N_12046);
nor U16061 (N_16061,N_13895,N_14415);
or U16062 (N_16062,N_14052,N_13887);
and U16063 (N_16063,N_13549,N_14516);
nor U16064 (N_16064,N_12397,N_14013);
xnor U16065 (N_16065,N_12481,N_13444);
nand U16066 (N_16066,N_13111,N_14790);
nand U16067 (N_16067,N_12018,N_14522);
and U16068 (N_16068,N_13649,N_14435);
or U16069 (N_16069,N_13231,N_12090);
and U16070 (N_16070,N_14963,N_12587);
and U16071 (N_16071,N_13802,N_13155);
nand U16072 (N_16072,N_13436,N_13054);
nor U16073 (N_16073,N_12790,N_13090);
or U16074 (N_16074,N_13147,N_14919);
nand U16075 (N_16075,N_14265,N_13544);
nor U16076 (N_16076,N_12464,N_13430);
nor U16077 (N_16077,N_13530,N_13566);
or U16078 (N_16078,N_14182,N_12197);
nor U16079 (N_16079,N_13733,N_13261);
nand U16080 (N_16080,N_14197,N_14270);
nand U16081 (N_16081,N_12627,N_13850);
nand U16082 (N_16082,N_14345,N_14481);
and U16083 (N_16083,N_14880,N_14650);
nand U16084 (N_16084,N_12875,N_12827);
nor U16085 (N_16085,N_12782,N_14797);
xnor U16086 (N_16086,N_14414,N_12891);
and U16087 (N_16087,N_13069,N_12265);
nor U16088 (N_16088,N_12024,N_12335);
or U16089 (N_16089,N_12413,N_13386);
or U16090 (N_16090,N_12928,N_14602);
nor U16091 (N_16091,N_12048,N_12059);
nor U16092 (N_16092,N_13395,N_13918);
or U16093 (N_16093,N_13042,N_12566);
and U16094 (N_16094,N_14737,N_13394);
or U16095 (N_16095,N_13152,N_12207);
nor U16096 (N_16096,N_14153,N_13035);
nor U16097 (N_16097,N_12467,N_13667);
nand U16098 (N_16098,N_13854,N_12507);
and U16099 (N_16099,N_13191,N_12336);
or U16100 (N_16100,N_13183,N_13681);
nor U16101 (N_16101,N_14233,N_12465);
and U16102 (N_16102,N_13855,N_14984);
and U16103 (N_16103,N_12725,N_14086);
nand U16104 (N_16104,N_14034,N_14291);
or U16105 (N_16105,N_13823,N_13632);
nor U16106 (N_16106,N_14581,N_13325);
nor U16107 (N_16107,N_14866,N_14130);
or U16108 (N_16108,N_14864,N_14446);
or U16109 (N_16109,N_12640,N_14761);
and U16110 (N_16110,N_14353,N_14571);
nand U16111 (N_16111,N_12444,N_14832);
xnor U16112 (N_16112,N_13640,N_14133);
nand U16113 (N_16113,N_12687,N_14796);
and U16114 (N_16114,N_12604,N_12110);
nor U16115 (N_16115,N_13350,N_13257);
and U16116 (N_16116,N_14082,N_13438);
nand U16117 (N_16117,N_12388,N_14822);
nand U16118 (N_16118,N_13656,N_14894);
xor U16119 (N_16119,N_13019,N_13771);
and U16120 (N_16120,N_12305,N_12976);
or U16121 (N_16121,N_13982,N_12279);
and U16122 (N_16122,N_14726,N_14940);
xor U16123 (N_16123,N_14872,N_13786);
or U16124 (N_16124,N_13738,N_13364);
and U16125 (N_16125,N_13540,N_13481);
or U16126 (N_16126,N_14593,N_14560);
nand U16127 (N_16127,N_13757,N_12406);
xor U16128 (N_16128,N_12907,N_12608);
and U16129 (N_16129,N_14427,N_13796);
xnor U16130 (N_16130,N_12544,N_14279);
and U16131 (N_16131,N_13324,N_12810);
nor U16132 (N_16132,N_12710,N_12530);
or U16133 (N_16133,N_14011,N_13644);
and U16134 (N_16134,N_12377,N_12146);
and U16135 (N_16135,N_13068,N_13777);
and U16136 (N_16136,N_13963,N_14506);
nor U16137 (N_16137,N_13291,N_14607);
or U16138 (N_16138,N_14857,N_12494);
or U16139 (N_16139,N_12578,N_12591);
nand U16140 (N_16140,N_13397,N_14744);
nor U16141 (N_16141,N_14486,N_14511);
and U16142 (N_16142,N_14001,N_12191);
or U16143 (N_16143,N_14176,N_13903);
and U16144 (N_16144,N_12613,N_14040);
or U16145 (N_16145,N_12986,N_12187);
nor U16146 (N_16146,N_12615,N_14075);
or U16147 (N_16147,N_14923,N_13584);
nand U16148 (N_16148,N_14502,N_13707);
and U16149 (N_16149,N_13148,N_12382);
or U16150 (N_16150,N_14005,N_12881);
or U16151 (N_16151,N_14118,N_12210);
xor U16152 (N_16152,N_12091,N_13564);
or U16153 (N_16153,N_12750,N_12905);
and U16154 (N_16154,N_13251,N_13033);
nor U16155 (N_16155,N_12325,N_12572);
and U16156 (N_16156,N_13580,N_14340);
and U16157 (N_16157,N_13485,N_14770);
and U16158 (N_16158,N_13674,N_13216);
or U16159 (N_16159,N_13886,N_13074);
nor U16160 (N_16160,N_12745,N_13603);
nor U16161 (N_16161,N_13785,N_12512);
nand U16162 (N_16162,N_14191,N_13144);
and U16163 (N_16163,N_12906,N_14986);
and U16164 (N_16164,N_14802,N_12763);
nand U16165 (N_16165,N_13451,N_14305);
nand U16166 (N_16166,N_14501,N_13143);
xnor U16167 (N_16167,N_12103,N_14997);
and U16168 (N_16168,N_13199,N_14367);
or U16169 (N_16169,N_14262,N_12679);
and U16170 (N_16170,N_12200,N_13151);
nor U16171 (N_16171,N_14629,N_12456);
or U16172 (N_16172,N_13382,N_14282);
and U16173 (N_16173,N_12872,N_14937);
or U16174 (N_16174,N_13255,N_12077);
xnor U16175 (N_16175,N_13932,N_13358);
and U16176 (N_16176,N_14543,N_13115);
and U16177 (N_16177,N_13552,N_12042);
nor U16178 (N_16178,N_14890,N_12306);
and U16179 (N_16179,N_12154,N_14736);
nand U16180 (N_16180,N_13861,N_14179);
nand U16181 (N_16181,N_12766,N_12583);
and U16182 (N_16182,N_13724,N_12773);
nand U16183 (N_16183,N_12671,N_13957);
or U16184 (N_16184,N_12408,N_12557);
or U16185 (N_16185,N_12729,N_13494);
nor U16186 (N_16186,N_14739,N_13285);
nand U16187 (N_16187,N_13925,N_12762);
xor U16188 (N_16188,N_13812,N_14215);
nand U16189 (N_16189,N_14577,N_12165);
xnor U16190 (N_16190,N_13691,N_12205);
nor U16191 (N_16191,N_14971,N_12775);
nor U16192 (N_16192,N_14465,N_12681);
or U16193 (N_16193,N_14205,N_14752);
nor U16194 (N_16194,N_14552,N_13824);
nand U16195 (N_16195,N_14158,N_14026);
and U16196 (N_16196,N_13779,N_12739);
and U16197 (N_16197,N_12628,N_13619);
nand U16198 (N_16198,N_14372,N_13130);
and U16199 (N_16199,N_12768,N_12134);
nand U16200 (N_16200,N_13213,N_12600);
or U16201 (N_16201,N_14173,N_13141);
nand U16202 (N_16202,N_13082,N_12297);
or U16203 (N_16203,N_13006,N_13772);
nand U16204 (N_16204,N_13749,N_12795);
nand U16205 (N_16205,N_13490,N_14879);
and U16206 (N_16206,N_13100,N_14166);
nor U16207 (N_16207,N_12233,N_14456);
nor U16208 (N_16208,N_14599,N_14068);
nor U16209 (N_16209,N_12717,N_13448);
or U16210 (N_16210,N_14849,N_13113);
or U16211 (N_16211,N_13728,N_12924);
nand U16212 (N_16212,N_13720,N_12664);
nor U16213 (N_16213,N_13252,N_14675);
nand U16214 (N_16214,N_12794,N_14311);
nor U16215 (N_16215,N_13639,N_13099);
nand U16216 (N_16216,N_12948,N_14236);
or U16217 (N_16217,N_14257,N_12229);
and U16218 (N_16218,N_14094,N_12736);
nor U16219 (N_16219,N_13628,N_13410);
nand U16220 (N_16220,N_14947,N_14556);
or U16221 (N_16221,N_12195,N_13161);
or U16222 (N_16222,N_12350,N_12415);
and U16223 (N_16223,N_14493,N_13638);
xor U16224 (N_16224,N_13256,N_12903);
nand U16225 (N_16225,N_12541,N_13933);
or U16226 (N_16226,N_14952,N_13536);
nor U16227 (N_16227,N_14967,N_12404);
nor U16228 (N_16228,N_14701,N_13298);
nor U16229 (N_16229,N_13923,N_13300);
or U16230 (N_16230,N_14125,N_12616);
nor U16231 (N_16231,N_12190,N_14656);
nor U16232 (N_16232,N_14828,N_14107);
nor U16233 (N_16233,N_12820,N_12749);
nand U16234 (N_16234,N_14290,N_13412);
or U16235 (N_16235,N_13417,N_14254);
nor U16236 (N_16236,N_13218,N_13614);
and U16237 (N_16237,N_12471,N_12201);
nand U16238 (N_16238,N_13505,N_13466);
nand U16239 (N_16239,N_14942,N_13238);
nor U16240 (N_16240,N_14473,N_13819);
and U16241 (N_16241,N_14293,N_14220);
xor U16242 (N_16242,N_14448,N_12468);
and U16243 (N_16243,N_13400,N_13202);
nor U16244 (N_16244,N_13421,N_14789);
nand U16245 (N_16245,N_13565,N_14413);
and U16246 (N_16246,N_12239,N_13071);
or U16247 (N_16247,N_14003,N_13695);
and U16248 (N_16248,N_12819,N_13592);
xor U16249 (N_16249,N_14325,N_13567);
nor U16250 (N_16250,N_13768,N_14829);
and U16251 (N_16251,N_14302,N_12734);
and U16252 (N_16252,N_13474,N_13784);
nor U16253 (N_16253,N_13160,N_12823);
nand U16254 (N_16254,N_14131,N_12011);
nor U16255 (N_16255,N_12495,N_14195);
and U16256 (N_16256,N_12299,N_13322);
nor U16257 (N_16257,N_13847,N_14921);
nor U16258 (N_16258,N_12211,N_13700);
xnor U16259 (N_16259,N_12878,N_14445);
and U16260 (N_16260,N_12862,N_14022);
nor U16261 (N_16261,N_14154,N_12362);
nand U16262 (N_16262,N_13301,N_13789);
nor U16263 (N_16263,N_14476,N_13362);
nor U16264 (N_16264,N_14324,N_12452);
and U16265 (N_16265,N_12879,N_12601);
nor U16266 (N_16266,N_13904,N_12535);
xor U16267 (N_16267,N_12841,N_13365);
xor U16268 (N_16268,N_13415,N_13997);
nor U16269 (N_16269,N_13046,N_12919);
nor U16270 (N_16270,N_14948,N_14544);
and U16271 (N_16271,N_13058,N_12105);
and U16272 (N_16272,N_13582,N_14045);
and U16273 (N_16273,N_13057,N_13615);
xnor U16274 (N_16274,N_13822,N_14596);
nand U16275 (N_16275,N_12309,N_12915);
or U16276 (N_16276,N_14527,N_12727);
and U16277 (N_16277,N_14585,N_14733);
nor U16278 (N_16278,N_14813,N_12000);
nor U16279 (N_16279,N_14015,N_13630);
nor U16280 (N_16280,N_12372,N_13568);
nor U16281 (N_16281,N_13902,N_13118);
nand U16282 (N_16282,N_14618,N_14664);
nand U16283 (N_16283,N_13702,N_12241);
nor U16284 (N_16284,N_13488,N_13705);
xor U16285 (N_16285,N_13519,N_14144);
nor U16286 (N_16286,N_13675,N_12340);
and U16287 (N_16287,N_12085,N_14364);
or U16288 (N_16288,N_13545,N_14490);
or U16289 (N_16289,N_13648,N_14169);
and U16290 (N_16290,N_13831,N_13499);
and U16291 (N_16291,N_14652,N_14121);
nor U16292 (N_16292,N_12222,N_14672);
nor U16293 (N_16293,N_12251,N_14623);
nand U16294 (N_16294,N_13563,N_13992);
or U16295 (N_16295,N_14174,N_14201);
nor U16296 (N_16296,N_13970,N_14051);
nor U16297 (N_16297,N_12175,N_13804);
nand U16298 (N_16298,N_13909,N_12318);
and U16299 (N_16299,N_14225,N_12695);
nand U16300 (N_16300,N_14021,N_12401);
or U16301 (N_16301,N_14924,N_14455);
and U16302 (N_16302,N_14764,N_14557);
nand U16303 (N_16303,N_13664,N_12778);
and U16304 (N_16304,N_13283,N_14341);
or U16305 (N_16305,N_14856,N_13049);
nor U16306 (N_16306,N_12419,N_14145);
or U16307 (N_16307,N_12798,N_12561);
or U16308 (N_16308,N_14226,N_12994);
xor U16309 (N_16309,N_13529,N_14528);
nor U16310 (N_16310,N_12978,N_14430);
and U16311 (N_16311,N_12162,N_14896);
nor U16312 (N_16312,N_12204,N_14274);
nand U16313 (N_16313,N_13168,N_12065);
nor U16314 (N_16314,N_14071,N_13110);
nor U16315 (N_16315,N_14538,N_14334);
or U16316 (N_16316,N_13003,N_13443);
nand U16317 (N_16317,N_12901,N_13013);
nand U16318 (N_16318,N_14716,N_13983);
and U16319 (N_16319,N_14016,N_12989);
or U16320 (N_16320,N_12152,N_12580);
and U16321 (N_16321,N_13939,N_12588);
and U16322 (N_16322,N_12356,N_13446);
nand U16323 (N_16323,N_13363,N_12125);
nor U16324 (N_16324,N_14061,N_13087);
nand U16325 (N_16325,N_13306,N_13973);
and U16326 (N_16326,N_13434,N_14609);
nor U16327 (N_16327,N_14062,N_12033);
and U16328 (N_16328,N_12107,N_13052);
or U16329 (N_16329,N_12506,N_14708);
and U16330 (N_16330,N_14030,N_14336);
or U16331 (N_16331,N_13357,N_14433);
and U16332 (N_16332,N_14114,N_12921);
xnor U16333 (N_16333,N_14962,N_12258);
nand U16334 (N_16334,N_12466,N_12759);
xnor U16335 (N_16335,N_14710,N_12582);
nor U16336 (N_16336,N_13699,N_14160);
nor U16337 (N_16337,N_12478,N_12548);
nand U16338 (N_16338,N_13945,N_12477);
nor U16339 (N_16339,N_13163,N_12301);
and U16340 (N_16340,N_14659,N_12968);
nor U16341 (N_16341,N_12833,N_12393);
nor U16342 (N_16342,N_13975,N_14671);
nor U16343 (N_16343,N_13843,N_14008);
xor U16344 (N_16344,N_12558,N_14307);
nor U16345 (N_16345,N_13857,N_12859);
or U16346 (N_16346,N_13716,N_13839);
and U16347 (N_16347,N_12386,N_12682);
or U16348 (N_16348,N_12649,N_12206);
xor U16349 (N_16349,N_12549,N_14155);
and U16350 (N_16350,N_13641,N_14206);
and U16351 (N_16351,N_12523,N_14632);
nand U16352 (N_16352,N_13271,N_12294);
or U16353 (N_16353,N_14070,N_13825);
and U16354 (N_16354,N_14548,N_12177);
and U16355 (N_16355,N_12108,N_12271);
xor U16356 (N_16356,N_14513,N_14231);
or U16357 (N_16357,N_12677,N_13411);
nand U16358 (N_16358,N_14667,N_13969);
nand U16359 (N_16359,N_12267,N_13940);
nand U16360 (N_16360,N_12140,N_12183);
and U16361 (N_16361,N_12617,N_13884);
or U16362 (N_16362,N_14755,N_14149);
xnor U16363 (N_16363,N_12776,N_12007);
or U16364 (N_16364,N_14085,N_14743);
nand U16365 (N_16365,N_14352,N_14893);
xor U16366 (N_16366,N_12867,N_12817);
and U16367 (N_16367,N_12365,N_12116);
or U16368 (N_16368,N_14286,N_14582);
or U16369 (N_16369,N_14111,N_14135);
and U16370 (N_16370,N_14268,N_12639);
nand U16371 (N_16371,N_13533,N_12412);
nor U16372 (N_16372,N_14079,N_13591);
and U16373 (N_16373,N_12049,N_13081);
or U16374 (N_16374,N_13468,N_13856);
or U16375 (N_16375,N_14786,N_14622);
nor U16376 (N_16376,N_13380,N_14261);
xor U16377 (N_16377,N_14033,N_13559);
nand U16378 (N_16378,N_14213,N_12349);
and U16379 (N_16379,N_14657,N_14988);
nand U16380 (N_16380,N_13770,N_14798);
nor U16381 (N_16381,N_13129,N_13302);
nand U16382 (N_16382,N_14646,N_14780);
nor U16383 (N_16383,N_14361,N_13634);
nor U16384 (N_16384,N_12296,N_13790);
nor U16385 (N_16385,N_14831,N_14989);
nor U16386 (N_16386,N_12440,N_14993);
and U16387 (N_16387,N_14645,N_12756);
nor U16388 (N_16388,N_14488,N_13138);
nor U16389 (N_16389,N_14519,N_12655);
nor U16390 (N_16390,N_14417,N_14074);
and U16391 (N_16391,N_14576,N_13776);
nor U16392 (N_16392,N_14795,N_12212);
nor U16393 (N_16393,N_12266,N_13122);
and U16394 (N_16394,N_12575,N_12486);
and U16395 (N_16395,N_12897,N_14251);
nand U16396 (N_16396,N_12387,N_12475);
nor U16397 (N_16397,N_14076,N_14408);
and U16398 (N_16398,N_12813,N_13694);
and U16399 (N_16399,N_12215,N_14938);
nand U16400 (N_16400,N_14842,N_12716);
nand U16401 (N_16401,N_13556,N_12883);
nor U16402 (N_16402,N_13960,N_12842);
or U16403 (N_16403,N_14504,N_12938);
nor U16404 (N_16404,N_13984,N_13952);
nor U16405 (N_16405,N_12914,N_13085);
nor U16406 (N_16406,N_12660,N_12957);
and U16407 (N_16407,N_12652,N_13758);
nand U16408 (N_16408,N_13440,N_13596);
and U16409 (N_16409,N_14442,N_13422);
nand U16410 (N_16410,N_12016,N_14437);
and U16411 (N_16411,N_12983,N_13097);
or U16412 (N_16412,N_14871,N_13517);
or U16413 (N_16413,N_14626,N_13942);
xnor U16414 (N_16414,N_13321,N_14067);
nor U16415 (N_16415,N_13483,N_14983);
or U16416 (N_16416,N_12036,N_12253);
and U16417 (N_16417,N_13575,N_12344);
or U16418 (N_16418,N_12367,N_12159);
nand U16419 (N_16419,N_12618,N_13117);
nor U16420 (N_16420,N_13774,N_14394);
nor U16421 (N_16421,N_13910,N_12922);
or U16422 (N_16422,N_12713,N_12227);
or U16423 (N_16423,N_12307,N_13025);
and U16424 (N_16424,N_12424,N_12960);
xor U16425 (N_16425,N_12783,N_12054);
nand U16426 (N_16426,N_13765,N_13684);
nand U16427 (N_16427,N_13629,N_14681);
nand U16428 (N_16428,N_12101,N_12062);
nor U16429 (N_16429,N_13387,N_13604);
and U16430 (N_16430,N_13426,N_13107);
and U16431 (N_16431,N_13187,N_14349);
nand U16432 (N_16432,N_13994,N_13073);
and U16433 (N_16433,N_13423,N_12929);
and U16434 (N_16434,N_12949,N_12912);
and U16435 (N_16435,N_13714,N_14069);
xor U16436 (N_16436,N_12524,N_13921);
xor U16437 (N_16437,N_14054,N_14368);
nand U16438 (N_16438,N_14253,N_12590);
nand U16439 (N_16439,N_12282,N_14883);
or U16440 (N_16440,N_14783,N_14171);
and U16441 (N_16441,N_13877,N_14698);
and U16442 (N_16442,N_14840,N_13510);
nand U16443 (N_16443,N_14064,N_12944);
nand U16444 (N_16444,N_13844,N_14065);
or U16445 (N_16445,N_12853,N_13678);
and U16446 (N_16446,N_13617,N_13653);
xor U16447 (N_16447,N_12777,N_13102);
and U16448 (N_16448,N_14562,N_13814);
nor U16449 (N_16449,N_13595,N_12115);
or U16450 (N_16450,N_14695,N_13841);
and U16451 (N_16451,N_12637,N_14007);
nor U16452 (N_16452,N_13220,N_13818);
and U16453 (N_16453,N_12479,N_14029);
nand U16454 (N_16454,N_12259,N_12225);
and U16455 (N_16455,N_13375,N_13741);
and U16456 (N_16456,N_14777,N_12329);
or U16457 (N_16457,N_14416,N_13532);
nand U16458 (N_16458,N_13015,N_12564);
or U16459 (N_16459,N_12194,N_14816);
or U16460 (N_16460,N_12004,N_12956);
nand U16461 (N_16461,N_14193,N_12260);
or U16462 (N_16462,N_14159,N_12861);
xor U16463 (N_16463,N_13858,N_13865);
nor U16464 (N_16464,N_12686,N_14601);
nor U16465 (N_16465,N_13349,N_13503);
nor U16466 (N_16466,N_14178,N_12690);
nand U16467 (N_16467,N_13180,N_13767);
xnor U16468 (N_16468,N_13197,N_14479);
nand U16469 (N_16469,N_12163,N_12189);
or U16470 (N_16470,N_14929,N_14697);
nor U16471 (N_16471,N_12379,N_14185);
and U16472 (N_16472,N_14235,N_14080);
or U16473 (N_16473,N_12913,N_13763);
and U16474 (N_16474,N_14677,N_14142);
xnor U16475 (N_16475,N_12053,N_14202);
nor U16476 (N_16476,N_13605,N_12482);
nor U16477 (N_16477,N_13156,N_12630);
and U16478 (N_16478,N_12339,N_13701);
xnor U16479 (N_16479,N_14041,N_14092);
or U16480 (N_16480,N_13590,N_12619);
xnor U16481 (N_16481,N_14407,N_13606);
nand U16482 (N_16482,N_12043,N_13808);
and U16483 (N_16483,N_12772,N_12636);
and U16484 (N_16484,N_12537,N_13762);
or U16485 (N_16485,N_12243,N_13600);
nand U16486 (N_16486,N_12579,N_12173);
xnor U16487 (N_16487,N_14686,N_14886);
or U16488 (N_16488,N_14383,N_13801);
nand U16489 (N_16489,N_12123,N_14358);
or U16490 (N_16490,N_14232,N_13158);
and U16491 (N_16491,N_14463,N_14913);
nand U16492 (N_16492,N_12355,N_12998);
or U16493 (N_16493,N_14961,N_12268);
nand U16494 (N_16494,N_12760,N_14218);
or U16495 (N_16495,N_13247,N_13840);
nor U16496 (N_16496,N_12044,N_12045);
or U16497 (N_16497,N_12153,N_12400);
nor U16498 (N_16498,N_13313,N_13658);
nand U16499 (N_16499,N_13516,N_14175);
nand U16500 (N_16500,N_12922,N_14655);
nor U16501 (N_16501,N_13828,N_12890);
or U16502 (N_16502,N_13580,N_13931);
and U16503 (N_16503,N_14164,N_14276);
nand U16504 (N_16504,N_13801,N_14041);
nor U16505 (N_16505,N_12055,N_12478);
nor U16506 (N_16506,N_13378,N_13526);
nor U16507 (N_16507,N_12610,N_13928);
nand U16508 (N_16508,N_13493,N_13685);
nor U16509 (N_16509,N_12115,N_14262);
nor U16510 (N_16510,N_13579,N_14431);
nor U16511 (N_16511,N_13839,N_14491);
or U16512 (N_16512,N_12939,N_12972);
nor U16513 (N_16513,N_13788,N_14964);
or U16514 (N_16514,N_12620,N_14794);
nor U16515 (N_16515,N_14375,N_13359);
and U16516 (N_16516,N_12362,N_12042);
or U16517 (N_16517,N_13187,N_13324);
and U16518 (N_16518,N_14108,N_14011);
and U16519 (N_16519,N_12021,N_12235);
nand U16520 (N_16520,N_13965,N_13187);
xnor U16521 (N_16521,N_14557,N_13079);
and U16522 (N_16522,N_13180,N_12734);
or U16523 (N_16523,N_12163,N_13976);
nor U16524 (N_16524,N_12233,N_14746);
nand U16525 (N_16525,N_13983,N_13363);
and U16526 (N_16526,N_14616,N_14194);
nand U16527 (N_16527,N_14625,N_12396);
or U16528 (N_16528,N_12116,N_14483);
and U16529 (N_16529,N_13488,N_12774);
or U16530 (N_16530,N_12405,N_14226);
nor U16531 (N_16531,N_12459,N_13214);
or U16532 (N_16532,N_13543,N_12958);
nand U16533 (N_16533,N_14350,N_12553);
xor U16534 (N_16534,N_14721,N_12818);
and U16535 (N_16535,N_14684,N_13253);
nor U16536 (N_16536,N_13173,N_13241);
nor U16537 (N_16537,N_14319,N_12360);
nand U16538 (N_16538,N_12431,N_14035);
nand U16539 (N_16539,N_12430,N_13820);
nand U16540 (N_16540,N_12992,N_13853);
or U16541 (N_16541,N_12561,N_14391);
nor U16542 (N_16542,N_12999,N_13210);
xnor U16543 (N_16543,N_12285,N_13488);
and U16544 (N_16544,N_12161,N_13073);
and U16545 (N_16545,N_12188,N_12005);
nor U16546 (N_16546,N_13547,N_12136);
and U16547 (N_16547,N_14862,N_13455);
nor U16548 (N_16548,N_12350,N_13966);
nor U16549 (N_16549,N_12751,N_12431);
or U16550 (N_16550,N_12255,N_12152);
nand U16551 (N_16551,N_12568,N_14668);
nand U16552 (N_16552,N_12163,N_12489);
xor U16553 (N_16553,N_12633,N_13353);
and U16554 (N_16554,N_13710,N_12116);
nor U16555 (N_16555,N_12603,N_14558);
xor U16556 (N_16556,N_13695,N_14291);
nand U16557 (N_16557,N_14401,N_12211);
and U16558 (N_16558,N_12509,N_14468);
nor U16559 (N_16559,N_14696,N_12839);
nor U16560 (N_16560,N_12651,N_12260);
or U16561 (N_16561,N_13040,N_13595);
nor U16562 (N_16562,N_14349,N_14602);
or U16563 (N_16563,N_13774,N_12367);
nor U16564 (N_16564,N_12678,N_13998);
nor U16565 (N_16565,N_13004,N_13891);
nand U16566 (N_16566,N_14978,N_14776);
or U16567 (N_16567,N_13084,N_12740);
or U16568 (N_16568,N_13553,N_14876);
and U16569 (N_16569,N_13027,N_14056);
nor U16570 (N_16570,N_13843,N_13127);
or U16571 (N_16571,N_12940,N_14925);
or U16572 (N_16572,N_12834,N_12478);
nor U16573 (N_16573,N_13445,N_13391);
or U16574 (N_16574,N_12628,N_12077);
xor U16575 (N_16575,N_13042,N_14145);
xor U16576 (N_16576,N_14292,N_12845);
or U16577 (N_16577,N_14774,N_14525);
and U16578 (N_16578,N_14441,N_12177);
nand U16579 (N_16579,N_14272,N_14463);
or U16580 (N_16580,N_12095,N_13181);
nor U16581 (N_16581,N_13808,N_12968);
or U16582 (N_16582,N_12225,N_14187);
nor U16583 (N_16583,N_13584,N_13406);
nand U16584 (N_16584,N_12469,N_13057);
and U16585 (N_16585,N_13983,N_14560);
and U16586 (N_16586,N_12898,N_12239);
nor U16587 (N_16587,N_13487,N_14979);
or U16588 (N_16588,N_13478,N_12443);
and U16589 (N_16589,N_14695,N_13201);
and U16590 (N_16590,N_12927,N_14249);
or U16591 (N_16591,N_12578,N_14425);
and U16592 (N_16592,N_14410,N_12253);
and U16593 (N_16593,N_13769,N_13487);
nor U16594 (N_16594,N_12971,N_12071);
and U16595 (N_16595,N_13909,N_12226);
nand U16596 (N_16596,N_14401,N_12372);
nor U16597 (N_16597,N_13585,N_14491);
or U16598 (N_16598,N_14653,N_12439);
nand U16599 (N_16599,N_14159,N_13145);
or U16600 (N_16600,N_14179,N_13279);
xor U16601 (N_16601,N_12769,N_14035);
nor U16602 (N_16602,N_14685,N_13399);
nor U16603 (N_16603,N_12312,N_12544);
or U16604 (N_16604,N_14143,N_13278);
or U16605 (N_16605,N_14522,N_14007);
nand U16606 (N_16606,N_13039,N_14731);
or U16607 (N_16607,N_14104,N_13379);
xnor U16608 (N_16608,N_12851,N_14840);
and U16609 (N_16609,N_14384,N_12908);
and U16610 (N_16610,N_14104,N_14495);
or U16611 (N_16611,N_14101,N_13577);
and U16612 (N_16612,N_14893,N_14473);
and U16613 (N_16613,N_12956,N_13955);
and U16614 (N_16614,N_13532,N_13792);
and U16615 (N_16615,N_14683,N_13030);
nand U16616 (N_16616,N_12140,N_12486);
nand U16617 (N_16617,N_13757,N_12678);
nand U16618 (N_16618,N_13028,N_12777);
and U16619 (N_16619,N_13691,N_12640);
xnor U16620 (N_16620,N_14743,N_13443);
nor U16621 (N_16621,N_13518,N_14257);
nand U16622 (N_16622,N_12758,N_12051);
and U16623 (N_16623,N_13902,N_13790);
and U16624 (N_16624,N_14089,N_13908);
xor U16625 (N_16625,N_14289,N_12981);
and U16626 (N_16626,N_13109,N_12552);
or U16627 (N_16627,N_14455,N_12371);
or U16628 (N_16628,N_14201,N_13735);
or U16629 (N_16629,N_14852,N_12737);
xor U16630 (N_16630,N_13833,N_13918);
or U16631 (N_16631,N_12158,N_14027);
xor U16632 (N_16632,N_13474,N_14627);
or U16633 (N_16633,N_13083,N_12712);
or U16634 (N_16634,N_13777,N_14304);
xor U16635 (N_16635,N_12969,N_12870);
nand U16636 (N_16636,N_14500,N_13473);
nand U16637 (N_16637,N_12971,N_12809);
nand U16638 (N_16638,N_14977,N_12118);
nand U16639 (N_16639,N_13475,N_14088);
nand U16640 (N_16640,N_12819,N_13665);
and U16641 (N_16641,N_12782,N_14700);
or U16642 (N_16642,N_13480,N_14321);
nand U16643 (N_16643,N_13064,N_12566);
nor U16644 (N_16644,N_14766,N_12501);
and U16645 (N_16645,N_12761,N_13663);
and U16646 (N_16646,N_13985,N_14301);
nand U16647 (N_16647,N_13337,N_14810);
xnor U16648 (N_16648,N_12607,N_14744);
and U16649 (N_16649,N_13997,N_12280);
nor U16650 (N_16650,N_12471,N_14635);
xnor U16651 (N_16651,N_12997,N_13757);
or U16652 (N_16652,N_14503,N_13891);
or U16653 (N_16653,N_13373,N_14661);
and U16654 (N_16654,N_12138,N_12146);
and U16655 (N_16655,N_12429,N_13587);
nor U16656 (N_16656,N_12407,N_13605);
nor U16657 (N_16657,N_14016,N_14088);
and U16658 (N_16658,N_13980,N_12903);
nand U16659 (N_16659,N_14533,N_12862);
and U16660 (N_16660,N_14781,N_14198);
nand U16661 (N_16661,N_13247,N_12598);
nand U16662 (N_16662,N_12968,N_12377);
and U16663 (N_16663,N_12591,N_13781);
nor U16664 (N_16664,N_12028,N_13758);
xor U16665 (N_16665,N_14503,N_12635);
or U16666 (N_16666,N_14980,N_14992);
nor U16667 (N_16667,N_14155,N_13776);
nand U16668 (N_16668,N_12031,N_12157);
nor U16669 (N_16669,N_14088,N_12050);
or U16670 (N_16670,N_12081,N_12729);
and U16671 (N_16671,N_14217,N_12699);
nor U16672 (N_16672,N_12130,N_12779);
or U16673 (N_16673,N_12817,N_13294);
nand U16674 (N_16674,N_13070,N_12603);
and U16675 (N_16675,N_13051,N_14552);
nor U16676 (N_16676,N_13777,N_12865);
nand U16677 (N_16677,N_13790,N_12965);
nor U16678 (N_16678,N_13699,N_12634);
and U16679 (N_16679,N_12973,N_12179);
and U16680 (N_16680,N_13219,N_12740);
nand U16681 (N_16681,N_14633,N_12037);
and U16682 (N_16682,N_14100,N_14089);
or U16683 (N_16683,N_14305,N_12508);
and U16684 (N_16684,N_12664,N_13572);
and U16685 (N_16685,N_12832,N_12296);
nand U16686 (N_16686,N_13129,N_14694);
or U16687 (N_16687,N_13361,N_12109);
and U16688 (N_16688,N_12799,N_13393);
nor U16689 (N_16689,N_13766,N_14440);
nand U16690 (N_16690,N_14212,N_14449);
xor U16691 (N_16691,N_13986,N_14824);
xor U16692 (N_16692,N_12535,N_12353);
and U16693 (N_16693,N_12201,N_14475);
nor U16694 (N_16694,N_14244,N_14473);
nand U16695 (N_16695,N_14041,N_14134);
nor U16696 (N_16696,N_13731,N_12119);
or U16697 (N_16697,N_13230,N_13061);
and U16698 (N_16698,N_12637,N_14762);
nor U16699 (N_16699,N_13975,N_12276);
or U16700 (N_16700,N_13616,N_12343);
nor U16701 (N_16701,N_13676,N_14812);
and U16702 (N_16702,N_14692,N_12584);
nand U16703 (N_16703,N_14576,N_14118);
and U16704 (N_16704,N_13139,N_14219);
xor U16705 (N_16705,N_14506,N_13526);
nor U16706 (N_16706,N_12936,N_12889);
or U16707 (N_16707,N_12050,N_13440);
xnor U16708 (N_16708,N_12086,N_14276);
and U16709 (N_16709,N_12945,N_14400);
or U16710 (N_16710,N_12996,N_12406);
xor U16711 (N_16711,N_14118,N_14310);
and U16712 (N_16712,N_12624,N_14991);
or U16713 (N_16713,N_13999,N_14800);
and U16714 (N_16714,N_12288,N_13795);
or U16715 (N_16715,N_13312,N_14242);
nand U16716 (N_16716,N_14721,N_13598);
nand U16717 (N_16717,N_13146,N_12436);
and U16718 (N_16718,N_13952,N_14102);
nor U16719 (N_16719,N_13502,N_14135);
or U16720 (N_16720,N_14568,N_14959);
and U16721 (N_16721,N_13725,N_12403);
nor U16722 (N_16722,N_14867,N_13116);
and U16723 (N_16723,N_12989,N_12600);
nor U16724 (N_16724,N_12562,N_13408);
nor U16725 (N_16725,N_14359,N_14531);
xnor U16726 (N_16726,N_14614,N_13983);
nand U16727 (N_16727,N_12929,N_12881);
xnor U16728 (N_16728,N_14946,N_12593);
nand U16729 (N_16729,N_12025,N_12854);
nand U16730 (N_16730,N_13574,N_12679);
or U16731 (N_16731,N_13381,N_14759);
xnor U16732 (N_16732,N_13437,N_13339);
nand U16733 (N_16733,N_14437,N_13776);
and U16734 (N_16734,N_14690,N_12631);
nand U16735 (N_16735,N_13888,N_13534);
and U16736 (N_16736,N_12648,N_13383);
nand U16737 (N_16737,N_14807,N_12547);
or U16738 (N_16738,N_14707,N_12272);
and U16739 (N_16739,N_13205,N_13533);
and U16740 (N_16740,N_14610,N_14792);
nand U16741 (N_16741,N_12031,N_12494);
nand U16742 (N_16742,N_12580,N_14581);
nor U16743 (N_16743,N_12951,N_14335);
nor U16744 (N_16744,N_13655,N_14291);
nor U16745 (N_16745,N_12323,N_13283);
nand U16746 (N_16746,N_12925,N_12982);
nor U16747 (N_16747,N_12431,N_14046);
or U16748 (N_16748,N_14860,N_14166);
nand U16749 (N_16749,N_14031,N_12755);
xnor U16750 (N_16750,N_14083,N_12106);
or U16751 (N_16751,N_12217,N_14667);
nand U16752 (N_16752,N_13005,N_13560);
or U16753 (N_16753,N_12322,N_12522);
nor U16754 (N_16754,N_12300,N_13545);
and U16755 (N_16755,N_14702,N_13985);
or U16756 (N_16756,N_13458,N_12348);
or U16757 (N_16757,N_14061,N_14497);
or U16758 (N_16758,N_13528,N_12914);
nor U16759 (N_16759,N_13524,N_13947);
nor U16760 (N_16760,N_14883,N_12742);
nand U16761 (N_16761,N_12668,N_12188);
and U16762 (N_16762,N_12870,N_12087);
xnor U16763 (N_16763,N_14218,N_14639);
nand U16764 (N_16764,N_14147,N_14334);
nor U16765 (N_16765,N_13439,N_14504);
nand U16766 (N_16766,N_13610,N_14937);
xor U16767 (N_16767,N_13924,N_13447);
and U16768 (N_16768,N_14440,N_13103);
nand U16769 (N_16769,N_13957,N_12730);
nor U16770 (N_16770,N_12211,N_13211);
xor U16771 (N_16771,N_13258,N_12494);
xor U16772 (N_16772,N_12588,N_12085);
nor U16773 (N_16773,N_13979,N_14254);
xnor U16774 (N_16774,N_12940,N_13263);
nand U16775 (N_16775,N_13015,N_13792);
nor U16776 (N_16776,N_13894,N_14309);
and U16777 (N_16777,N_13138,N_12855);
or U16778 (N_16778,N_12277,N_12173);
nor U16779 (N_16779,N_13006,N_14724);
nor U16780 (N_16780,N_13622,N_14267);
nor U16781 (N_16781,N_14842,N_14188);
or U16782 (N_16782,N_14057,N_13143);
xor U16783 (N_16783,N_14466,N_12500);
nand U16784 (N_16784,N_13217,N_14431);
and U16785 (N_16785,N_13334,N_13039);
nand U16786 (N_16786,N_14733,N_14566);
xnor U16787 (N_16787,N_12040,N_12905);
and U16788 (N_16788,N_12595,N_14954);
nor U16789 (N_16789,N_12491,N_12508);
or U16790 (N_16790,N_14320,N_13466);
or U16791 (N_16791,N_14581,N_14565);
xnor U16792 (N_16792,N_12224,N_12598);
nand U16793 (N_16793,N_12160,N_14540);
nor U16794 (N_16794,N_13285,N_12066);
xnor U16795 (N_16795,N_14073,N_12941);
or U16796 (N_16796,N_13227,N_14456);
nor U16797 (N_16797,N_12502,N_13322);
nand U16798 (N_16798,N_13981,N_13645);
nor U16799 (N_16799,N_14355,N_13522);
and U16800 (N_16800,N_12626,N_12074);
or U16801 (N_16801,N_14073,N_12133);
nor U16802 (N_16802,N_14707,N_13159);
nor U16803 (N_16803,N_12687,N_12925);
nand U16804 (N_16804,N_13097,N_12635);
nor U16805 (N_16805,N_12885,N_14663);
nor U16806 (N_16806,N_12449,N_12742);
nand U16807 (N_16807,N_12296,N_12511);
and U16808 (N_16808,N_14863,N_14318);
and U16809 (N_16809,N_13661,N_13378);
xor U16810 (N_16810,N_14351,N_14324);
nor U16811 (N_16811,N_13864,N_13608);
nor U16812 (N_16812,N_13955,N_14581);
nor U16813 (N_16813,N_14049,N_14091);
or U16814 (N_16814,N_14576,N_13127);
nand U16815 (N_16815,N_12281,N_12531);
nor U16816 (N_16816,N_13493,N_13257);
and U16817 (N_16817,N_12707,N_14630);
and U16818 (N_16818,N_14240,N_12105);
nor U16819 (N_16819,N_14308,N_13658);
and U16820 (N_16820,N_14512,N_13044);
and U16821 (N_16821,N_13568,N_13051);
nor U16822 (N_16822,N_14120,N_12608);
nor U16823 (N_16823,N_12334,N_13078);
and U16824 (N_16824,N_13228,N_12739);
and U16825 (N_16825,N_14548,N_14123);
xnor U16826 (N_16826,N_14912,N_13138);
and U16827 (N_16827,N_14053,N_12523);
nand U16828 (N_16828,N_12074,N_12338);
or U16829 (N_16829,N_13970,N_14576);
nand U16830 (N_16830,N_13901,N_12299);
nor U16831 (N_16831,N_14333,N_13242);
and U16832 (N_16832,N_14402,N_12063);
or U16833 (N_16833,N_12891,N_14230);
or U16834 (N_16834,N_13167,N_12455);
or U16835 (N_16835,N_14698,N_12864);
nor U16836 (N_16836,N_14191,N_13086);
nor U16837 (N_16837,N_12430,N_12436);
xor U16838 (N_16838,N_13510,N_12263);
or U16839 (N_16839,N_12441,N_13064);
nor U16840 (N_16840,N_12836,N_13294);
and U16841 (N_16841,N_12489,N_13619);
nor U16842 (N_16842,N_14288,N_14674);
nor U16843 (N_16843,N_13497,N_13335);
nand U16844 (N_16844,N_13764,N_13311);
nand U16845 (N_16845,N_14739,N_14185);
nor U16846 (N_16846,N_14530,N_13257);
or U16847 (N_16847,N_12263,N_12775);
nand U16848 (N_16848,N_12725,N_14238);
and U16849 (N_16849,N_12614,N_12365);
and U16850 (N_16850,N_14854,N_14068);
nor U16851 (N_16851,N_14033,N_14941);
or U16852 (N_16852,N_12502,N_12536);
nor U16853 (N_16853,N_12690,N_14794);
and U16854 (N_16854,N_13477,N_14676);
nor U16855 (N_16855,N_12406,N_14376);
and U16856 (N_16856,N_14856,N_14237);
nand U16857 (N_16857,N_13712,N_14240);
and U16858 (N_16858,N_12810,N_14622);
or U16859 (N_16859,N_14901,N_13851);
or U16860 (N_16860,N_12964,N_12649);
nand U16861 (N_16861,N_14750,N_13316);
nand U16862 (N_16862,N_14263,N_12374);
xnor U16863 (N_16863,N_12774,N_14219);
nor U16864 (N_16864,N_13832,N_14120);
and U16865 (N_16865,N_13006,N_13596);
or U16866 (N_16866,N_12432,N_14605);
nor U16867 (N_16867,N_14821,N_14228);
nand U16868 (N_16868,N_13175,N_12922);
xor U16869 (N_16869,N_14220,N_12882);
nor U16870 (N_16870,N_14118,N_14883);
nand U16871 (N_16871,N_14160,N_12469);
nand U16872 (N_16872,N_12087,N_13903);
and U16873 (N_16873,N_13690,N_13280);
and U16874 (N_16874,N_14302,N_13115);
xnor U16875 (N_16875,N_14480,N_12796);
nor U16876 (N_16876,N_13736,N_13681);
nand U16877 (N_16877,N_13509,N_13644);
xor U16878 (N_16878,N_13030,N_12343);
and U16879 (N_16879,N_13349,N_12810);
or U16880 (N_16880,N_12226,N_14099);
nand U16881 (N_16881,N_14029,N_13322);
nand U16882 (N_16882,N_12478,N_13309);
or U16883 (N_16883,N_12549,N_14801);
nand U16884 (N_16884,N_14722,N_14216);
nor U16885 (N_16885,N_13120,N_13402);
and U16886 (N_16886,N_14728,N_14205);
nor U16887 (N_16887,N_12657,N_13846);
or U16888 (N_16888,N_14468,N_12939);
nand U16889 (N_16889,N_12223,N_12861);
and U16890 (N_16890,N_13004,N_13942);
and U16891 (N_16891,N_14247,N_12702);
xnor U16892 (N_16892,N_12134,N_14850);
nand U16893 (N_16893,N_14635,N_14807);
xnor U16894 (N_16894,N_13172,N_13948);
xnor U16895 (N_16895,N_12733,N_13212);
nor U16896 (N_16896,N_12257,N_13574);
or U16897 (N_16897,N_13744,N_12365);
and U16898 (N_16898,N_12976,N_12308);
nor U16899 (N_16899,N_13364,N_13163);
nand U16900 (N_16900,N_13078,N_13352);
nor U16901 (N_16901,N_13560,N_12853);
and U16902 (N_16902,N_13978,N_13658);
nor U16903 (N_16903,N_14215,N_14226);
or U16904 (N_16904,N_14121,N_12950);
nor U16905 (N_16905,N_12227,N_12434);
nand U16906 (N_16906,N_13892,N_14134);
xnor U16907 (N_16907,N_13968,N_12376);
nand U16908 (N_16908,N_14758,N_13043);
and U16909 (N_16909,N_12212,N_12546);
and U16910 (N_16910,N_14811,N_12922);
and U16911 (N_16911,N_14766,N_13887);
and U16912 (N_16912,N_12526,N_12375);
and U16913 (N_16913,N_13286,N_12818);
xor U16914 (N_16914,N_12217,N_12925);
nor U16915 (N_16915,N_14560,N_13779);
nor U16916 (N_16916,N_13473,N_13616);
nand U16917 (N_16917,N_14820,N_12023);
nor U16918 (N_16918,N_13508,N_13796);
xor U16919 (N_16919,N_14378,N_12864);
nor U16920 (N_16920,N_14547,N_12033);
or U16921 (N_16921,N_14893,N_14990);
or U16922 (N_16922,N_12322,N_14334);
nand U16923 (N_16923,N_13813,N_14287);
or U16924 (N_16924,N_14650,N_14177);
nor U16925 (N_16925,N_14472,N_12475);
nand U16926 (N_16926,N_13366,N_13135);
and U16927 (N_16927,N_12229,N_12953);
xor U16928 (N_16928,N_12518,N_13584);
or U16929 (N_16929,N_13817,N_13312);
nand U16930 (N_16930,N_14891,N_12977);
and U16931 (N_16931,N_12795,N_12289);
and U16932 (N_16932,N_13319,N_14132);
and U16933 (N_16933,N_14765,N_12011);
nand U16934 (N_16934,N_14931,N_13377);
xor U16935 (N_16935,N_13283,N_12790);
and U16936 (N_16936,N_13204,N_12975);
or U16937 (N_16937,N_12543,N_13012);
or U16938 (N_16938,N_12807,N_14562);
nand U16939 (N_16939,N_13721,N_13144);
or U16940 (N_16940,N_13889,N_12490);
nor U16941 (N_16941,N_12649,N_13277);
nor U16942 (N_16942,N_12428,N_14589);
nand U16943 (N_16943,N_13735,N_14955);
and U16944 (N_16944,N_13293,N_14822);
and U16945 (N_16945,N_14487,N_14053);
xor U16946 (N_16946,N_12831,N_12505);
nand U16947 (N_16947,N_14138,N_12830);
or U16948 (N_16948,N_12912,N_13272);
nand U16949 (N_16949,N_13299,N_14134);
and U16950 (N_16950,N_14526,N_13273);
and U16951 (N_16951,N_12648,N_13596);
and U16952 (N_16952,N_12489,N_14044);
and U16953 (N_16953,N_14236,N_13716);
nand U16954 (N_16954,N_14926,N_14675);
nor U16955 (N_16955,N_14473,N_12553);
nand U16956 (N_16956,N_13217,N_14143);
or U16957 (N_16957,N_12347,N_14432);
and U16958 (N_16958,N_14962,N_14073);
and U16959 (N_16959,N_13542,N_14348);
nor U16960 (N_16960,N_12029,N_13690);
nand U16961 (N_16961,N_13979,N_14755);
nand U16962 (N_16962,N_13693,N_13314);
or U16963 (N_16963,N_12764,N_12930);
and U16964 (N_16964,N_13062,N_14085);
and U16965 (N_16965,N_13776,N_12522);
xnor U16966 (N_16966,N_14180,N_13562);
and U16967 (N_16967,N_12270,N_14222);
or U16968 (N_16968,N_13084,N_14202);
nor U16969 (N_16969,N_13393,N_13974);
nand U16970 (N_16970,N_14245,N_13777);
nand U16971 (N_16971,N_13340,N_13053);
nand U16972 (N_16972,N_13906,N_12132);
and U16973 (N_16973,N_12872,N_13307);
nor U16974 (N_16974,N_14980,N_12034);
nand U16975 (N_16975,N_14473,N_12776);
and U16976 (N_16976,N_13807,N_12944);
or U16977 (N_16977,N_12714,N_14559);
and U16978 (N_16978,N_12519,N_13497);
nand U16979 (N_16979,N_12392,N_12142);
or U16980 (N_16980,N_12743,N_14259);
nor U16981 (N_16981,N_13570,N_13300);
nor U16982 (N_16982,N_14277,N_13891);
and U16983 (N_16983,N_14755,N_13221);
nand U16984 (N_16984,N_13045,N_13299);
nand U16985 (N_16985,N_14262,N_12731);
nor U16986 (N_16986,N_12129,N_13124);
or U16987 (N_16987,N_14287,N_13350);
or U16988 (N_16988,N_14919,N_13582);
or U16989 (N_16989,N_12423,N_14229);
and U16990 (N_16990,N_14517,N_13909);
or U16991 (N_16991,N_14693,N_12403);
nand U16992 (N_16992,N_14187,N_14722);
nor U16993 (N_16993,N_14997,N_13754);
nand U16994 (N_16994,N_12970,N_13702);
nand U16995 (N_16995,N_14896,N_13397);
or U16996 (N_16996,N_12798,N_12685);
nand U16997 (N_16997,N_14681,N_12500);
or U16998 (N_16998,N_12462,N_13897);
nand U16999 (N_16999,N_14006,N_14297);
nand U17000 (N_17000,N_12896,N_13955);
or U17001 (N_17001,N_13120,N_14232);
or U17002 (N_17002,N_14192,N_13560);
or U17003 (N_17003,N_13642,N_12181);
and U17004 (N_17004,N_13714,N_12416);
and U17005 (N_17005,N_13432,N_12594);
and U17006 (N_17006,N_12283,N_12047);
nor U17007 (N_17007,N_12179,N_13305);
xnor U17008 (N_17008,N_13897,N_14211);
and U17009 (N_17009,N_12209,N_12418);
nor U17010 (N_17010,N_12767,N_14654);
and U17011 (N_17011,N_12245,N_13220);
or U17012 (N_17012,N_12097,N_14115);
and U17013 (N_17013,N_13475,N_13053);
and U17014 (N_17014,N_13176,N_13069);
or U17015 (N_17015,N_14073,N_12323);
and U17016 (N_17016,N_14137,N_12792);
or U17017 (N_17017,N_14146,N_13066);
nand U17018 (N_17018,N_13182,N_12195);
and U17019 (N_17019,N_12295,N_14061);
nand U17020 (N_17020,N_13745,N_12563);
or U17021 (N_17021,N_12292,N_14939);
xor U17022 (N_17022,N_14958,N_12486);
and U17023 (N_17023,N_14745,N_14894);
xor U17024 (N_17024,N_14969,N_14762);
nor U17025 (N_17025,N_14577,N_14663);
or U17026 (N_17026,N_14424,N_13055);
nor U17027 (N_17027,N_13162,N_13071);
nor U17028 (N_17028,N_12976,N_13500);
or U17029 (N_17029,N_14539,N_12688);
xnor U17030 (N_17030,N_14180,N_13940);
nand U17031 (N_17031,N_13405,N_14447);
xor U17032 (N_17032,N_12650,N_12199);
nand U17033 (N_17033,N_14228,N_14760);
nand U17034 (N_17034,N_12462,N_13770);
and U17035 (N_17035,N_14014,N_13254);
xnor U17036 (N_17036,N_14143,N_13594);
xor U17037 (N_17037,N_14661,N_12744);
or U17038 (N_17038,N_12089,N_13791);
or U17039 (N_17039,N_13717,N_14058);
and U17040 (N_17040,N_14424,N_14177);
xor U17041 (N_17041,N_12507,N_12048);
nor U17042 (N_17042,N_12148,N_13648);
nand U17043 (N_17043,N_14161,N_13049);
or U17044 (N_17044,N_13658,N_14436);
nand U17045 (N_17045,N_14162,N_14687);
or U17046 (N_17046,N_12702,N_14648);
and U17047 (N_17047,N_12813,N_14938);
nor U17048 (N_17048,N_12247,N_13551);
and U17049 (N_17049,N_13340,N_14661);
and U17050 (N_17050,N_13627,N_14629);
or U17051 (N_17051,N_14110,N_13176);
xor U17052 (N_17052,N_14436,N_12629);
nor U17053 (N_17053,N_14372,N_14109);
or U17054 (N_17054,N_14218,N_12024);
or U17055 (N_17055,N_12037,N_14225);
nor U17056 (N_17056,N_13500,N_12046);
nor U17057 (N_17057,N_12307,N_12243);
and U17058 (N_17058,N_12791,N_14880);
nand U17059 (N_17059,N_14564,N_12960);
and U17060 (N_17060,N_13224,N_13098);
or U17061 (N_17061,N_13843,N_13460);
xnor U17062 (N_17062,N_13706,N_12036);
nand U17063 (N_17063,N_12038,N_12324);
and U17064 (N_17064,N_13387,N_14951);
nor U17065 (N_17065,N_12129,N_12670);
xnor U17066 (N_17066,N_13938,N_14634);
nor U17067 (N_17067,N_13422,N_14041);
nor U17068 (N_17068,N_12518,N_13282);
nor U17069 (N_17069,N_12245,N_13639);
or U17070 (N_17070,N_13603,N_14165);
or U17071 (N_17071,N_13282,N_14759);
and U17072 (N_17072,N_14487,N_12202);
xnor U17073 (N_17073,N_12603,N_13274);
and U17074 (N_17074,N_13215,N_12079);
xor U17075 (N_17075,N_12371,N_13029);
or U17076 (N_17076,N_14648,N_14601);
and U17077 (N_17077,N_13374,N_14208);
nand U17078 (N_17078,N_13892,N_13846);
nand U17079 (N_17079,N_13365,N_14423);
nand U17080 (N_17080,N_14206,N_13548);
nor U17081 (N_17081,N_12150,N_14989);
nand U17082 (N_17082,N_12192,N_13897);
nand U17083 (N_17083,N_13218,N_12476);
and U17084 (N_17084,N_13414,N_13363);
nor U17085 (N_17085,N_13345,N_14061);
nor U17086 (N_17086,N_14488,N_14431);
or U17087 (N_17087,N_13709,N_13821);
nor U17088 (N_17088,N_14739,N_13551);
and U17089 (N_17089,N_13067,N_13260);
or U17090 (N_17090,N_14777,N_12506);
or U17091 (N_17091,N_12968,N_14885);
nand U17092 (N_17092,N_14811,N_13196);
or U17093 (N_17093,N_12612,N_12364);
and U17094 (N_17094,N_13888,N_12176);
nor U17095 (N_17095,N_12834,N_13294);
or U17096 (N_17096,N_14027,N_14251);
xor U17097 (N_17097,N_12000,N_12672);
nand U17098 (N_17098,N_12889,N_13409);
nor U17099 (N_17099,N_14887,N_14712);
and U17100 (N_17100,N_13601,N_13054);
nand U17101 (N_17101,N_14905,N_14423);
or U17102 (N_17102,N_14701,N_13954);
or U17103 (N_17103,N_12769,N_12616);
xnor U17104 (N_17104,N_12541,N_13350);
xor U17105 (N_17105,N_13539,N_12518);
xor U17106 (N_17106,N_12418,N_13079);
xor U17107 (N_17107,N_12438,N_13545);
nor U17108 (N_17108,N_14595,N_13016);
or U17109 (N_17109,N_14861,N_14820);
and U17110 (N_17110,N_14317,N_13001);
and U17111 (N_17111,N_14289,N_13378);
nor U17112 (N_17112,N_13275,N_14902);
nand U17113 (N_17113,N_14019,N_12128);
nand U17114 (N_17114,N_13662,N_13836);
and U17115 (N_17115,N_13338,N_14878);
nor U17116 (N_17116,N_12385,N_13586);
or U17117 (N_17117,N_12699,N_14268);
nand U17118 (N_17118,N_12652,N_12157);
nor U17119 (N_17119,N_14043,N_13949);
and U17120 (N_17120,N_12380,N_12733);
and U17121 (N_17121,N_12937,N_14637);
nor U17122 (N_17122,N_14551,N_12019);
nor U17123 (N_17123,N_14750,N_13754);
and U17124 (N_17124,N_13195,N_13112);
nand U17125 (N_17125,N_13681,N_14951);
nand U17126 (N_17126,N_12721,N_12412);
and U17127 (N_17127,N_12298,N_13514);
nor U17128 (N_17128,N_14849,N_14417);
nor U17129 (N_17129,N_13060,N_14588);
nand U17130 (N_17130,N_12136,N_12943);
nor U17131 (N_17131,N_13254,N_14118);
and U17132 (N_17132,N_14017,N_14241);
and U17133 (N_17133,N_13040,N_12473);
nor U17134 (N_17134,N_12512,N_12991);
nor U17135 (N_17135,N_14199,N_12171);
xor U17136 (N_17136,N_13294,N_14336);
or U17137 (N_17137,N_12534,N_14017);
nand U17138 (N_17138,N_12563,N_13658);
or U17139 (N_17139,N_13185,N_14162);
or U17140 (N_17140,N_13243,N_12894);
nand U17141 (N_17141,N_14116,N_14651);
or U17142 (N_17142,N_12875,N_13669);
nor U17143 (N_17143,N_14443,N_13918);
and U17144 (N_17144,N_12847,N_12495);
and U17145 (N_17145,N_12056,N_13327);
nor U17146 (N_17146,N_14812,N_14582);
nand U17147 (N_17147,N_14715,N_13156);
nor U17148 (N_17148,N_14338,N_13891);
xor U17149 (N_17149,N_12346,N_12343);
and U17150 (N_17150,N_14514,N_14997);
or U17151 (N_17151,N_14489,N_12116);
nand U17152 (N_17152,N_13955,N_13840);
and U17153 (N_17153,N_13732,N_13488);
and U17154 (N_17154,N_12835,N_14743);
nor U17155 (N_17155,N_14568,N_12991);
nand U17156 (N_17156,N_12272,N_13125);
xnor U17157 (N_17157,N_13380,N_14936);
and U17158 (N_17158,N_12070,N_13557);
or U17159 (N_17159,N_13385,N_12378);
nand U17160 (N_17160,N_12578,N_14543);
xnor U17161 (N_17161,N_14526,N_14332);
nor U17162 (N_17162,N_12309,N_12434);
or U17163 (N_17163,N_12268,N_13084);
and U17164 (N_17164,N_13569,N_14577);
nand U17165 (N_17165,N_14821,N_12619);
xnor U17166 (N_17166,N_12057,N_13286);
or U17167 (N_17167,N_12576,N_13133);
nand U17168 (N_17168,N_14345,N_14565);
and U17169 (N_17169,N_12247,N_13623);
xnor U17170 (N_17170,N_14974,N_12985);
nand U17171 (N_17171,N_13196,N_13859);
nor U17172 (N_17172,N_12212,N_14469);
or U17173 (N_17173,N_12825,N_12374);
nor U17174 (N_17174,N_12393,N_13086);
nor U17175 (N_17175,N_14359,N_13336);
nand U17176 (N_17176,N_14698,N_12201);
nand U17177 (N_17177,N_12556,N_14135);
xnor U17178 (N_17178,N_14701,N_13447);
nor U17179 (N_17179,N_13547,N_14439);
and U17180 (N_17180,N_14083,N_14341);
or U17181 (N_17181,N_13388,N_13630);
nor U17182 (N_17182,N_13330,N_13879);
or U17183 (N_17183,N_14153,N_14700);
nand U17184 (N_17184,N_12082,N_14577);
and U17185 (N_17185,N_12959,N_12753);
nand U17186 (N_17186,N_13489,N_12575);
or U17187 (N_17187,N_13332,N_13901);
and U17188 (N_17188,N_12144,N_14883);
and U17189 (N_17189,N_14427,N_12969);
nor U17190 (N_17190,N_13610,N_14177);
nand U17191 (N_17191,N_13734,N_14413);
nor U17192 (N_17192,N_14038,N_13394);
and U17193 (N_17193,N_12303,N_13861);
nand U17194 (N_17194,N_13636,N_14870);
and U17195 (N_17195,N_12280,N_14665);
nand U17196 (N_17196,N_14920,N_13433);
nand U17197 (N_17197,N_12737,N_13344);
nand U17198 (N_17198,N_14160,N_12572);
nor U17199 (N_17199,N_12279,N_14660);
and U17200 (N_17200,N_12558,N_13951);
nand U17201 (N_17201,N_13830,N_14110);
nand U17202 (N_17202,N_12389,N_13382);
and U17203 (N_17203,N_13048,N_13119);
nand U17204 (N_17204,N_14017,N_12645);
and U17205 (N_17205,N_13416,N_13170);
nand U17206 (N_17206,N_14201,N_12888);
and U17207 (N_17207,N_13924,N_13711);
nor U17208 (N_17208,N_14290,N_14283);
xor U17209 (N_17209,N_14954,N_12816);
nor U17210 (N_17210,N_12828,N_12173);
nor U17211 (N_17211,N_14350,N_13593);
and U17212 (N_17212,N_13266,N_14392);
nor U17213 (N_17213,N_12411,N_14865);
nor U17214 (N_17214,N_14893,N_14296);
nor U17215 (N_17215,N_13957,N_14254);
xor U17216 (N_17216,N_13377,N_12451);
and U17217 (N_17217,N_14895,N_12433);
or U17218 (N_17218,N_12553,N_14799);
nand U17219 (N_17219,N_13396,N_14052);
and U17220 (N_17220,N_13619,N_14352);
nor U17221 (N_17221,N_14034,N_12851);
nor U17222 (N_17222,N_14370,N_14726);
nor U17223 (N_17223,N_14868,N_12492);
or U17224 (N_17224,N_13513,N_14033);
nand U17225 (N_17225,N_14862,N_13107);
nand U17226 (N_17226,N_13291,N_12492);
nor U17227 (N_17227,N_12742,N_14081);
nor U17228 (N_17228,N_14880,N_13193);
nand U17229 (N_17229,N_12897,N_14684);
nor U17230 (N_17230,N_14236,N_14975);
nor U17231 (N_17231,N_14045,N_12638);
xor U17232 (N_17232,N_14691,N_13838);
and U17233 (N_17233,N_13387,N_14467);
nand U17234 (N_17234,N_12916,N_12450);
nor U17235 (N_17235,N_14544,N_12422);
nand U17236 (N_17236,N_12349,N_12623);
or U17237 (N_17237,N_14501,N_13349);
nand U17238 (N_17238,N_12294,N_13732);
nor U17239 (N_17239,N_12451,N_13241);
or U17240 (N_17240,N_13141,N_14738);
nand U17241 (N_17241,N_12861,N_12181);
nand U17242 (N_17242,N_14776,N_12147);
nor U17243 (N_17243,N_14786,N_12780);
or U17244 (N_17244,N_14192,N_13896);
and U17245 (N_17245,N_12490,N_14702);
nand U17246 (N_17246,N_14500,N_14715);
nand U17247 (N_17247,N_13692,N_14258);
nor U17248 (N_17248,N_13984,N_14202);
nand U17249 (N_17249,N_14258,N_13753);
nor U17250 (N_17250,N_12851,N_14417);
and U17251 (N_17251,N_13450,N_14887);
and U17252 (N_17252,N_14649,N_12244);
nor U17253 (N_17253,N_14711,N_14371);
nor U17254 (N_17254,N_12434,N_13742);
xnor U17255 (N_17255,N_13935,N_12536);
and U17256 (N_17256,N_13822,N_12550);
or U17257 (N_17257,N_14424,N_13320);
or U17258 (N_17258,N_12354,N_13826);
nand U17259 (N_17259,N_12416,N_13186);
or U17260 (N_17260,N_13433,N_12509);
xor U17261 (N_17261,N_14680,N_12615);
and U17262 (N_17262,N_13821,N_14684);
nor U17263 (N_17263,N_14041,N_13683);
nand U17264 (N_17264,N_14666,N_13273);
nand U17265 (N_17265,N_13898,N_12696);
nor U17266 (N_17266,N_13370,N_13934);
xnor U17267 (N_17267,N_14128,N_13587);
nand U17268 (N_17268,N_14953,N_14984);
nand U17269 (N_17269,N_13545,N_13998);
or U17270 (N_17270,N_14427,N_14622);
nand U17271 (N_17271,N_13586,N_14930);
nor U17272 (N_17272,N_12402,N_13184);
nand U17273 (N_17273,N_12803,N_13787);
nor U17274 (N_17274,N_13430,N_13138);
and U17275 (N_17275,N_14326,N_14061);
xnor U17276 (N_17276,N_14613,N_14938);
or U17277 (N_17277,N_13767,N_12843);
xnor U17278 (N_17278,N_13781,N_13754);
nor U17279 (N_17279,N_12340,N_14111);
and U17280 (N_17280,N_12289,N_12279);
nand U17281 (N_17281,N_14385,N_12217);
xnor U17282 (N_17282,N_14701,N_14582);
nand U17283 (N_17283,N_12248,N_12823);
nor U17284 (N_17284,N_14430,N_14550);
and U17285 (N_17285,N_14137,N_14530);
nor U17286 (N_17286,N_14324,N_13488);
and U17287 (N_17287,N_14790,N_14968);
nand U17288 (N_17288,N_14817,N_14304);
or U17289 (N_17289,N_13457,N_12857);
nand U17290 (N_17290,N_12423,N_13500);
nor U17291 (N_17291,N_12451,N_13095);
nor U17292 (N_17292,N_13350,N_14833);
and U17293 (N_17293,N_14053,N_12370);
nand U17294 (N_17294,N_14750,N_12658);
and U17295 (N_17295,N_14782,N_12837);
and U17296 (N_17296,N_13662,N_14737);
xor U17297 (N_17297,N_14509,N_14260);
or U17298 (N_17298,N_14581,N_14739);
nor U17299 (N_17299,N_14922,N_14125);
and U17300 (N_17300,N_12209,N_12212);
and U17301 (N_17301,N_12411,N_12174);
or U17302 (N_17302,N_12484,N_12630);
or U17303 (N_17303,N_13193,N_14871);
nand U17304 (N_17304,N_13656,N_12735);
or U17305 (N_17305,N_14068,N_13606);
xnor U17306 (N_17306,N_12592,N_13005);
xor U17307 (N_17307,N_14717,N_12290);
or U17308 (N_17308,N_13934,N_13340);
or U17309 (N_17309,N_14424,N_14642);
and U17310 (N_17310,N_13510,N_14719);
or U17311 (N_17311,N_14223,N_13320);
and U17312 (N_17312,N_14283,N_12572);
or U17313 (N_17313,N_14937,N_12506);
and U17314 (N_17314,N_14605,N_13085);
and U17315 (N_17315,N_12719,N_13895);
nand U17316 (N_17316,N_12759,N_14422);
or U17317 (N_17317,N_14599,N_13109);
xnor U17318 (N_17318,N_12529,N_13620);
nand U17319 (N_17319,N_12145,N_14835);
xnor U17320 (N_17320,N_14210,N_14168);
nand U17321 (N_17321,N_13936,N_14061);
or U17322 (N_17322,N_14840,N_14323);
nand U17323 (N_17323,N_13934,N_13757);
and U17324 (N_17324,N_14205,N_13354);
nor U17325 (N_17325,N_14534,N_13764);
xnor U17326 (N_17326,N_14402,N_14503);
nor U17327 (N_17327,N_14437,N_12842);
and U17328 (N_17328,N_12686,N_12934);
nor U17329 (N_17329,N_13753,N_14358);
and U17330 (N_17330,N_14070,N_13849);
nand U17331 (N_17331,N_12670,N_12740);
xnor U17332 (N_17332,N_14162,N_14521);
and U17333 (N_17333,N_13432,N_13380);
xnor U17334 (N_17334,N_13406,N_13604);
nor U17335 (N_17335,N_14056,N_12449);
nand U17336 (N_17336,N_14589,N_12675);
nand U17337 (N_17337,N_13971,N_12060);
and U17338 (N_17338,N_14111,N_13371);
nor U17339 (N_17339,N_12123,N_14081);
nor U17340 (N_17340,N_12202,N_13062);
nor U17341 (N_17341,N_13174,N_13617);
xnor U17342 (N_17342,N_14998,N_12278);
or U17343 (N_17343,N_12466,N_13692);
or U17344 (N_17344,N_13233,N_13701);
or U17345 (N_17345,N_14265,N_12041);
nand U17346 (N_17346,N_12826,N_13552);
and U17347 (N_17347,N_14741,N_14830);
nand U17348 (N_17348,N_13766,N_14568);
xor U17349 (N_17349,N_12492,N_13264);
and U17350 (N_17350,N_14212,N_14811);
nor U17351 (N_17351,N_12191,N_14072);
nand U17352 (N_17352,N_12030,N_13048);
and U17353 (N_17353,N_13018,N_13714);
and U17354 (N_17354,N_12659,N_12461);
nor U17355 (N_17355,N_13554,N_12299);
xnor U17356 (N_17356,N_14382,N_13821);
nand U17357 (N_17357,N_13351,N_12173);
or U17358 (N_17358,N_12328,N_12531);
nor U17359 (N_17359,N_12617,N_13724);
xor U17360 (N_17360,N_12326,N_13693);
nor U17361 (N_17361,N_13768,N_12620);
and U17362 (N_17362,N_13452,N_12253);
nand U17363 (N_17363,N_13633,N_14653);
nand U17364 (N_17364,N_14305,N_14476);
nand U17365 (N_17365,N_14158,N_14616);
xnor U17366 (N_17366,N_13029,N_13352);
nor U17367 (N_17367,N_12664,N_13096);
nor U17368 (N_17368,N_14340,N_14816);
or U17369 (N_17369,N_12834,N_14984);
nand U17370 (N_17370,N_13400,N_12465);
xor U17371 (N_17371,N_14420,N_12383);
or U17372 (N_17372,N_14402,N_14118);
nand U17373 (N_17373,N_14616,N_12921);
nand U17374 (N_17374,N_14293,N_13449);
nand U17375 (N_17375,N_12270,N_14609);
or U17376 (N_17376,N_12243,N_12212);
and U17377 (N_17377,N_14069,N_14864);
xor U17378 (N_17378,N_14054,N_13401);
and U17379 (N_17379,N_14329,N_14459);
and U17380 (N_17380,N_13386,N_14129);
nor U17381 (N_17381,N_14982,N_13186);
or U17382 (N_17382,N_14329,N_14286);
nor U17383 (N_17383,N_14136,N_13292);
nor U17384 (N_17384,N_13636,N_12727);
or U17385 (N_17385,N_13676,N_14834);
nor U17386 (N_17386,N_13532,N_12228);
and U17387 (N_17387,N_13471,N_13831);
xnor U17388 (N_17388,N_14413,N_13232);
nand U17389 (N_17389,N_13087,N_14295);
nor U17390 (N_17390,N_12722,N_12179);
nor U17391 (N_17391,N_12163,N_12299);
nor U17392 (N_17392,N_13903,N_14152);
nor U17393 (N_17393,N_13644,N_13160);
and U17394 (N_17394,N_14729,N_14973);
nor U17395 (N_17395,N_14908,N_14937);
nor U17396 (N_17396,N_14435,N_13503);
nand U17397 (N_17397,N_12488,N_13503);
nor U17398 (N_17398,N_13040,N_12177);
or U17399 (N_17399,N_14410,N_14108);
xnor U17400 (N_17400,N_13722,N_14105);
or U17401 (N_17401,N_13842,N_14208);
or U17402 (N_17402,N_12519,N_12550);
and U17403 (N_17403,N_14590,N_14581);
and U17404 (N_17404,N_12036,N_12658);
or U17405 (N_17405,N_13838,N_12413);
xor U17406 (N_17406,N_14617,N_13383);
xor U17407 (N_17407,N_13263,N_13194);
xnor U17408 (N_17408,N_13903,N_13585);
and U17409 (N_17409,N_12103,N_14128);
nand U17410 (N_17410,N_13946,N_13145);
and U17411 (N_17411,N_13172,N_13633);
and U17412 (N_17412,N_12505,N_13857);
or U17413 (N_17413,N_13891,N_12003);
nand U17414 (N_17414,N_14320,N_12220);
and U17415 (N_17415,N_12352,N_13399);
nand U17416 (N_17416,N_13680,N_12492);
nor U17417 (N_17417,N_13097,N_13460);
and U17418 (N_17418,N_14975,N_12877);
or U17419 (N_17419,N_14147,N_13137);
and U17420 (N_17420,N_13327,N_14026);
xnor U17421 (N_17421,N_12617,N_14898);
nor U17422 (N_17422,N_12573,N_12072);
nor U17423 (N_17423,N_13095,N_14454);
xor U17424 (N_17424,N_13586,N_12607);
and U17425 (N_17425,N_14273,N_13925);
and U17426 (N_17426,N_13830,N_12422);
nand U17427 (N_17427,N_12294,N_12989);
or U17428 (N_17428,N_13417,N_12868);
or U17429 (N_17429,N_12489,N_14473);
and U17430 (N_17430,N_14210,N_14252);
nand U17431 (N_17431,N_13796,N_14642);
and U17432 (N_17432,N_13099,N_14170);
xnor U17433 (N_17433,N_12106,N_12035);
or U17434 (N_17434,N_14399,N_14447);
nand U17435 (N_17435,N_12224,N_14150);
and U17436 (N_17436,N_12472,N_13349);
or U17437 (N_17437,N_12038,N_13313);
nor U17438 (N_17438,N_13449,N_13311);
nand U17439 (N_17439,N_14717,N_13356);
and U17440 (N_17440,N_13837,N_12185);
or U17441 (N_17441,N_14939,N_12002);
nor U17442 (N_17442,N_13769,N_14585);
nor U17443 (N_17443,N_13125,N_12613);
and U17444 (N_17444,N_14245,N_14233);
and U17445 (N_17445,N_13386,N_12755);
or U17446 (N_17446,N_13661,N_14219);
and U17447 (N_17447,N_12846,N_14105);
or U17448 (N_17448,N_13236,N_12886);
nand U17449 (N_17449,N_14636,N_13642);
nand U17450 (N_17450,N_14876,N_12398);
and U17451 (N_17451,N_14431,N_13274);
xor U17452 (N_17452,N_12745,N_12401);
or U17453 (N_17453,N_12405,N_12117);
nand U17454 (N_17454,N_14408,N_14592);
or U17455 (N_17455,N_13239,N_13244);
xnor U17456 (N_17456,N_14432,N_14097);
nor U17457 (N_17457,N_14963,N_13908);
or U17458 (N_17458,N_12170,N_14527);
and U17459 (N_17459,N_12423,N_14368);
or U17460 (N_17460,N_14570,N_14688);
or U17461 (N_17461,N_13108,N_13132);
xnor U17462 (N_17462,N_13708,N_12394);
nor U17463 (N_17463,N_13703,N_12870);
and U17464 (N_17464,N_14083,N_12180);
xnor U17465 (N_17465,N_13701,N_13969);
nor U17466 (N_17466,N_12749,N_14836);
nand U17467 (N_17467,N_14288,N_13262);
nor U17468 (N_17468,N_12989,N_14716);
nand U17469 (N_17469,N_13014,N_14017);
and U17470 (N_17470,N_14988,N_14235);
nand U17471 (N_17471,N_13226,N_13588);
nor U17472 (N_17472,N_12394,N_13493);
or U17473 (N_17473,N_14045,N_12079);
nand U17474 (N_17474,N_14967,N_13413);
nor U17475 (N_17475,N_12168,N_12631);
nand U17476 (N_17476,N_14836,N_12329);
nor U17477 (N_17477,N_14823,N_13656);
and U17478 (N_17478,N_13950,N_14088);
nor U17479 (N_17479,N_14275,N_14621);
or U17480 (N_17480,N_12990,N_14732);
or U17481 (N_17481,N_14507,N_12196);
nor U17482 (N_17482,N_14317,N_14432);
or U17483 (N_17483,N_12657,N_12271);
or U17484 (N_17484,N_14993,N_14229);
nor U17485 (N_17485,N_12625,N_12031);
nand U17486 (N_17486,N_12493,N_14482);
or U17487 (N_17487,N_14972,N_12740);
nand U17488 (N_17488,N_12265,N_14280);
and U17489 (N_17489,N_14742,N_12841);
xnor U17490 (N_17490,N_13222,N_12430);
or U17491 (N_17491,N_12130,N_12014);
or U17492 (N_17492,N_14056,N_13955);
or U17493 (N_17493,N_13754,N_12820);
xor U17494 (N_17494,N_14860,N_14403);
and U17495 (N_17495,N_13113,N_13851);
and U17496 (N_17496,N_14550,N_13155);
nor U17497 (N_17497,N_13497,N_13881);
or U17498 (N_17498,N_13690,N_12172);
nand U17499 (N_17499,N_14388,N_14091);
and U17500 (N_17500,N_12687,N_14519);
and U17501 (N_17501,N_13312,N_13927);
nand U17502 (N_17502,N_14559,N_13117);
and U17503 (N_17503,N_14511,N_14954);
nor U17504 (N_17504,N_12039,N_13788);
or U17505 (N_17505,N_13435,N_13769);
and U17506 (N_17506,N_13319,N_12964);
nand U17507 (N_17507,N_12019,N_13204);
nor U17508 (N_17508,N_14806,N_14089);
xnor U17509 (N_17509,N_13523,N_12716);
nand U17510 (N_17510,N_12884,N_14702);
and U17511 (N_17511,N_13654,N_13737);
nor U17512 (N_17512,N_14063,N_14545);
and U17513 (N_17513,N_14220,N_14756);
nor U17514 (N_17514,N_13486,N_12989);
xor U17515 (N_17515,N_14946,N_12542);
nor U17516 (N_17516,N_12458,N_14645);
nand U17517 (N_17517,N_13947,N_14271);
or U17518 (N_17518,N_14220,N_12354);
nor U17519 (N_17519,N_12718,N_12035);
xor U17520 (N_17520,N_13289,N_12958);
nand U17521 (N_17521,N_14501,N_12478);
nor U17522 (N_17522,N_13562,N_12602);
nor U17523 (N_17523,N_14581,N_12680);
and U17524 (N_17524,N_13675,N_13727);
or U17525 (N_17525,N_13238,N_12380);
or U17526 (N_17526,N_13790,N_13392);
or U17527 (N_17527,N_13912,N_12747);
or U17528 (N_17528,N_14357,N_14772);
nor U17529 (N_17529,N_14805,N_14869);
nor U17530 (N_17530,N_14207,N_12280);
and U17531 (N_17531,N_14736,N_14516);
nor U17532 (N_17532,N_13549,N_13586);
nand U17533 (N_17533,N_12269,N_12671);
nand U17534 (N_17534,N_14176,N_14478);
nor U17535 (N_17535,N_14142,N_14123);
nor U17536 (N_17536,N_12790,N_14518);
nor U17537 (N_17537,N_13687,N_13462);
and U17538 (N_17538,N_12387,N_12535);
or U17539 (N_17539,N_12423,N_14858);
and U17540 (N_17540,N_13598,N_14529);
nand U17541 (N_17541,N_13218,N_12603);
nor U17542 (N_17542,N_14930,N_12838);
nor U17543 (N_17543,N_12782,N_13004);
or U17544 (N_17544,N_13830,N_12320);
nor U17545 (N_17545,N_13479,N_13008);
nand U17546 (N_17546,N_14772,N_13389);
nand U17547 (N_17547,N_12885,N_12075);
nor U17548 (N_17548,N_12233,N_14451);
and U17549 (N_17549,N_14299,N_12331);
and U17550 (N_17550,N_12955,N_12500);
or U17551 (N_17551,N_13958,N_14933);
nor U17552 (N_17552,N_14157,N_12584);
nand U17553 (N_17553,N_14852,N_12469);
or U17554 (N_17554,N_14767,N_14093);
xor U17555 (N_17555,N_14840,N_13413);
and U17556 (N_17556,N_13099,N_14932);
or U17557 (N_17557,N_13856,N_14762);
nand U17558 (N_17558,N_14247,N_13530);
and U17559 (N_17559,N_13990,N_14304);
nor U17560 (N_17560,N_14789,N_12143);
or U17561 (N_17561,N_13998,N_14656);
nor U17562 (N_17562,N_12229,N_14934);
nor U17563 (N_17563,N_14240,N_14359);
nor U17564 (N_17564,N_13358,N_13795);
or U17565 (N_17565,N_13295,N_14022);
nand U17566 (N_17566,N_12600,N_13592);
nand U17567 (N_17567,N_12905,N_14011);
or U17568 (N_17568,N_13343,N_14044);
or U17569 (N_17569,N_13705,N_14883);
nand U17570 (N_17570,N_13575,N_14607);
and U17571 (N_17571,N_12175,N_14203);
and U17572 (N_17572,N_13605,N_14416);
nand U17573 (N_17573,N_13307,N_14605);
nand U17574 (N_17574,N_12419,N_13325);
or U17575 (N_17575,N_12552,N_12868);
or U17576 (N_17576,N_14666,N_12364);
xor U17577 (N_17577,N_13870,N_14991);
nand U17578 (N_17578,N_14529,N_14720);
or U17579 (N_17579,N_13934,N_13119);
nor U17580 (N_17580,N_12473,N_13616);
or U17581 (N_17581,N_12576,N_14629);
nor U17582 (N_17582,N_12860,N_14062);
or U17583 (N_17583,N_12630,N_13437);
and U17584 (N_17584,N_12620,N_12532);
nand U17585 (N_17585,N_13284,N_13189);
nand U17586 (N_17586,N_13466,N_14937);
or U17587 (N_17587,N_12467,N_14895);
and U17588 (N_17588,N_14279,N_13178);
and U17589 (N_17589,N_14031,N_14626);
nand U17590 (N_17590,N_13852,N_13462);
and U17591 (N_17591,N_14102,N_13357);
or U17592 (N_17592,N_12771,N_14270);
and U17593 (N_17593,N_14908,N_12778);
and U17594 (N_17594,N_14485,N_13430);
nand U17595 (N_17595,N_14038,N_14804);
and U17596 (N_17596,N_12776,N_12488);
and U17597 (N_17597,N_12017,N_12172);
xor U17598 (N_17598,N_14535,N_12395);
nand U17599 (N_17599,N_13621,N_12944);
xor U17600 (N_17600,N_14010,N_13333);
or U17601 (N_17601,N_13458,N_12346);
nor U17602 (N_17602,N_12387,N_13708);
nand U17603 (N_17603,N_14512,N_12493);
nor U17604 (N_17604,N_12109,N_12736);
nand U17605 (N_17605,N_13845,N_12072);
nor U17606 (N_17606,N_14523,N_12821);
nor U17607 (N_17607,N_12690,N_12204);
nor U17608 (N_17608,N_13832,N_13066);
xnor U17609 (N_17609,N_13760,N_14498);
and U17610 (N_17610,N_13788,N_12473);
or U17611 (N_17611,N_12510,N_14585);
nor U17612 (N_17612,N_12399,N_13920);
nor U17613 (N_17613,N_14073,N_13461);
nand U17614 (N_17614,N_14361,N_13454);
nor U17615 (N_17615,N_12279,N_12709);
and U17616 (N_17616,N_13456,N_14775);
nand U17617 (N_17617,N_12804,N_13277);
or U17618 (N_17618,N_12682,N_12359);
nand U17619 (N_17619,N_14382,N_13533);
nand U17620 (N_17620,N_12430,N_12258);
or U17621 (N_17621,N_14361,N_12987);
xnor U17622 (N_17622,N_12634,N_14881);
nand U17623 (N_17623,N_12211,N_13348);
nor U17624 (N_17624,N_13447,N_14891);
and U17625 (N_17625,N_14257,N_14939);
or U17626 (N_17626,N_12649,N_12188);
nand U17627 (N_17627,N_12914,N_14631);
nand U17628 (N_17628,N_12947,N_12770);
or U17629 (N_17629,N_12795,N_12858);
nor U17630 (N_17630,N_13441,N_13996);
nand U17631 (N_17631,N_12501,N_14181);
and U17632 (N_17632,N_12559,N_12745);
nor U17633 (N_17633,N_13440,N_14005);
nand U17634 (N_17634,N_12085,N_12372);
or U17635 (N_17635,N_13145,N_14427);
nand U17636 (N_17636,N_12382,N_12984);
nor U17637 (N_17637,N_14233,N_14751);
nor U17638 (N_17638,N_12778,N_12313);
nand U17639 (N_17639,N_13866,N_14443);
and U17640 (N_17640,N_14278,N_13239);
and U17641 (N_17641,N_12350,N_14570);
or U17642 (N_17642,N_13992,N_14133);
and U17643 (N_17643,N_14234,N_13630);
nand U17644 (N_17644,N_14371,N_13229);
nand U17645 (N_17645,N_14211,N_14107);
and U17646 (N_17646,N_12991,N_14857);
or U17647 (N_17647,N_14350,N_12799);
or U17648 (N_17648,N_12759,N_14203);
nand U17649 (N_17649,N_13783,N_13658);
xor U17650 (N_17650,N_14549,N_13024);
or U17651 (N_17651,N_13000,N_13250);
or U17652 (N_17652,N_13500,N_14647);
or U17653 (N_17653,N_13794,N_13333);
xnor U17654 (N_17654,N_13825,N_14150);
nor U17655 (N_17655,N_13975,N_12065);
or U17656 (N_17656,N_13501,N_14951);
xnor U17657 (N_17657,N_13273,N_13727);
nor U17658 (N_17658,N_12815,N_14053);
and U17659 (N_17659,N_12332,N_13966);
xnor U17660 (N_17660,N_12118,N_12996);
nor U17661 (N_17661,N_14620,N_12847);
or U17662 (N_17662,N_13870,N_14714);
nor U17663 (N_17663,N_14507,N_12946);
or U17664 (N_17664,N_12592,N_14495);
or U17665 (N_17665,N_12558,N_14239);
nand U17666 (N_17666,N_13616,N_12082);
and U17667 (N_17667,N_12303,N_13022);
nand U17668 (N_17668,N_14391,N_14287);
nand U17669 (N_17669,N_12332,N_12706);
nand U17670 (N_17670,N_14050,N_12486);
nand U17671 (N_17671,N_13982,N_12247);
and U17672 (N_17672,N_14247,N_13078);
xnor U17673 (N_17673,N_14368,N_12996);
and U17674 (N_17674,N_13180,N_13654);
xor U17675 (N_17675,N_12716,N_13315);
and U17676 (N_17676,N_13860,N_14501);
nor U17677 (N_17677,N_12832,N_14213);
and U17678 (N_17678,N_13548,N_12902);
or U17679 (N_17679,N_12581,N_12237);
nor U17680 (N_17680,N_12685,N_14217);
and U17681 (N_17681,N_14835,N_12452);
or U17682 (N_17682,N_14030,N_12246);
nand U17683 (N_17683,N_13783,N_12567);
and U17684 (N_17684,N_14952,N_14124);
and U17685 (N_17685,N_12643,N_14858);
nand U17686 (N_17686,N_13355,N_12978);
nand U17687 (N_17687,N_12643,N_13630);
nand U17688 (N_17688,N_13067,N_13102);
or U17689 (N_17689,N_12500,N_12878);
nand U17690 (N_17690,N_13672,N_12436);
or U17691 (N_17691,N_14881,N_14228);
or U17692 (N_17692,N_13758,N_12097);
nand U17693 (N_17693,N_14046,N_12239);
nand U17694 (N_17694,N_14005,N_14431);
xor U17695 (N_17695,N_13133,N_14665);
nand U17696 (N_17696,N_13708,N_12216);
xnor U17697 (N_17697,N_13768,N_14288);
nand U17698 (N_17698,N_13274,N_12368);
nor U17699 (N_17699,N_14816,N_14848);
and U17700 (N_17700,N_12524,N_12847);
and U17701 (N_17701,N_13966,N_13510);
or U17702 (N_17702,N_12261,N_12383);
or U17703 (N_17703,N_13473,N_12443);
or U17704 (N_17704,N_14450,N_13768);
nor U17705 (N_17705,N_12324,N_12034);
and U17706 (N_17706,N_13874,N_13875);
or U17707 (N_17707,N_13897,N_12834);
or U17708 (N_17708,N_12256,N_13674);
and U17709 (N_17709,N_14379,N_14753);
nand U17710 (N_17710,N_13916,N_13808);
nor U17711 (N_17711,N_12421,N_13616);
nor U17712 (N_17712,N_12822,N_13885);
or U17713 (N_17713,N_12862,N_12263);
nand U17714 (N_17714,N_13766,N_13858);
xnor U17715 (N_17715,N_12234,N_14857);
and U17716 (N_17716,N_14470,N_14841);
nor U17717 (N_17717,N_14770,N_13079);
nor U17718 (N_17718,N_14435,N_13725);
nor U17719 (N_17719,N_12973,N_13066);
or U17720 (N_17720,N_12415,N_13507);
nor U17721 (N_17721,N_12600,N_13170);
nor U17722 (N_17722,N_13261,N_13993);
or U17723 (N_17723,N_14621,N_13712);
or U17724 (N_17724,N_13426,N_12515);
xnor U17725 (N_17725,N_14346,N_13948);
xnor U17726 (N_17726,N_13205,N_14743);
nor U17727 (N_17727,N_12150,N_14582);
and U17728 (N_17728,N_14210,N_13551);
nor U17729 (N_17729,N_12354,N_12055);
nor U17730 (N_17730,N_13180,N_14908);
and U17731 (N_17731,N_12866,N_14618);
nor U17732 (N_17732,N_14647,N_14016);
nor U17733 (N_17733,N_13379,N_13094);
nand U17734 (N_17734,N_14153,N_13104);
or U17735 (N_17735,N_14461,N_12199);
and U17736 (N_17736,N_13201,N_14125);
and U17737 (N_17737,N_13993,N_12334);
xor U17738 (N_17738,N_12689,N_14371);
nand U17739 (N_17739,N_12705,N_13445);
nand U17740 (N_17740,N_14754,N_13746);
nor U17741 (N_17741,N_14482,N_13649);
or U17742 (N_17742,N_13415,N_14061);
nor U17743 (N_17743,N_14123,N_12706);
or U17744 (N_17744,N_14966,N_14480);
or U17745 (N_17745,N_12366,N_14973);
or U17746 (N_17746,N_14943,N_14087);
or U17747 (N_17747,N_12632,N_14417);
nand U17748 (N_17748,N_14223,N_12673);
xnor U17749 (N_17749,N_13779,N_13885);
xnor U17750 (N_17750,N_13471,N_12311);
nor U17751 (N_17751,N_12023,N_14882);
or U17752 (N_17752,N_14623,N_14472);
nand U17753 (N_17753,N_12708,N_14054);
and U17754 (N_17754,N_13930,N_12833);
or U17755 (N_17755,N_14732,N_12965);
or U17756 (N_17756,N_12658,N_14341);
nand U17757 (N_17757,N_14856,N_14164);
or U17758 (N_17758,N_12980,N_14034);
nor U17759 (N_17759,N_12943,N_13669);
and U17760 (N_17760,N_13601,N_14694);
nand U17761 (N_17761,N_12586,N_12546);
xor U17762 (N_17762,N_13442,N_12729);
nand U17763 (N_17763,N_14412,N_14995);
nand U17764 (N_17764,N_14885,N_12675);
nor U17765 (N_17765,N_13800,N_12546);
nor U17766 (N_17766,N_12950,N_12396);
or U17767 (N_17767,N_13031,N_12168);
nor U17768 (N_17768,N_12181,N_13326);
and U17769 (N_17769,N_14507,N_14847);
nor U17770 (N_17770,N_14252,N_13432);
nor U17771 (N_17771,N_12986,N_12719);
nor U17772 (N_17772,N_14168,N_13070);
nor U17773 (N_17773,N_13927,N_13673);
nand U17774 (N_17774,N_12022,N_13017);
or U17775 (N_17775,N_12554,N_13375);
xor U17776 (N_17776,N_13588,N_13487);
nor U17777 (N_17777,N_13373,N_12549);
and U17778 (N_17778,N_12388,N_13163);
nand U17779 (N_17779,N_12441,N_13733);
and U17780 (N_17780,N_14190,N_12167);
nand U17781 (N_17781,N_12130,N_14194);
and U17782 (N_17782,N_14406,N_14878);
or U17783 (N_17783,N_13190,N_13729);
nor U17784 (N_17784,N_14612,N_12214);
and U17785 (N_17785,N_13791,N_12898);
and U17786 (N_17786,N_14875,N_13826);
or U17787 (N_17787,N_14037,N_14601);
nor U17788 (N_17788,N_14684,N_12576);
or U17789 (N_17789,N_12406,N_12898);
nor U17790 (N_17790,N_14025,N_14065);
or U17791 (N_17791,N_13189,N_12445);
nand U17792 (N_17792,N_13141,N_14568);
or U17793 (N_17793,N_13812,N_12697);
nor U17794 (N_17794,N_13028,N_12740);
or U17795 (N_17795,N_12486,N_13106);
nor U17796 (N_17796,N_12123,N_12634);
and U17797 (N_17797,N_13623,N_12577);
nor U17798 (N_17798,N_13780,N_12480);
nand U17799 (N_17799,N_14941,N_12041);
nor U17800 (N_17800,N_14296,N_13613);
and U17801 (N_17801,N_12285,N_14972);
nor U17802 (N_17802,N_12746,N_13280);
or U17803 (N_17803,N_14126,N_13289);
nor U17804 (N_17804,N_13976,N_13474);
or U17805 (N_17805,N_14949,N_13521);
nand U17806 (N_17806,N_14389,N_12848);
or U17807 (N_17807,N_12496,N_12935);
nand U17808 (N_17808,N_12223,N_14341);
nor U17809 (N_17809,N_12856,N_13267);
and U17810 (N_17810,N_13023,N_14017);
nand U17811 (N_17811,N_13575,N_13210);
nand U17812 (N_17812,N_14902,N_13284);
and U17813 (N_17813,N_14678,N_14046);
xor U17814 (N_17814,N_12484,N_13339);
nand U17815 (N_17815,N_14894,N_14248);
and U17816 (N_17816,N_13433,N_12844);
nand U17817 (N_17817,N_12110,N_13220);
nor U17818 (N_17818,N_13378,N_14957);
nand U17819 (N_17819,N_12490,N_14132);
or U17820 (N_17820,N_13744,N_14595);
xor U17821 (N_17821,N_12057,N_14257);
nand U17822 (N_17822,N_12864,N_13424);
nand U17823 (N_17823,N_13736,N_13834);
and U17824 (N_17824,N_13040,N_14898);
and U17825 (N_17825,N_14974,N_12411);
xor U17826 (N_17826,N_12897,N_13306);
or U17827 (N_17827,N_12138,N_14649);
nand U17828 (N_17828,N_13621,N_14966);
xnor U17829 (N_17829,N_14209,N_12880);
or U17830 (N_17830,N_12307,N_14297);
and U17831 (N_17831,N_12212,N_14355);
and U17832 (N_17832,N_12165,N_13159);
nand U17833 (N_17833,N_13616,N_13947);
nor U17834 (N_17834,N_13626,N_14732);
xnor U17835 (N_17835,N_13975,N_12728);
nand U17836 (N_17836,N_14886,N_13192);
and U17837 (N_17837,N_12314,N_14611);
and U17838 (N_17838,N_14021,N_14442);
and U17839 (N_17839,N_12070,N_12425);
nor U17840 (N_17840,N_14651,N_12572);
or U17841 (N_17841,N_14155,N_12471);
and U17842 (N_17842,N_12562,N_13356);
nor U17843 (N_17843,N_14798,N_12391);
and U17844 (N_17844,N_12887,N_12140);
nand U17845 (N_17845,N_14617,N_14429);
or U17846 (N_17846,N_13826,N_12817);
and U17847 (N_17847,N_12217,N_14235);
xor U17848 (N_17848,N_13524,N_13119);
and U17849 (N_17849,N_14119,N_12423);
nand U17850 (N_17850,N_14071,N_12998);
xnor U17851 (N_17851,N_13802,N_14767);
and U17852 (N_17852,N_12402,N_14696);
and U17853 (N_17853,N_13310,N_13762);
or U17854 (N_17854,N_12606,N_12359);
nand U17855 (N_17855,N_13074,N_12008);
nand U17856 (N_17856,N_13193,N_13263);
nand U17857 (N_17857,N_13512,N_14627);
nand U17858 (N_17858,N_14627,N_14069);
or U17859 (N_17859,N_14673,N_13868);
nor U17860 (N_17860,N_12317,N_13056);
xor U17861 (N_17861,N_13797,N_12986);
nand U17862 (N_17862,N_12786,N_13811);
nand U17863 (N_17863,N_12013,N_14960);
nand U17864 (N_17864,N_14212,N_12419);
xor U17865 (N_17865,N_14682,N_13474);
and U17866 (N_17866,N_13632,N_13714);
and U17867 (N_17867,N_14509,N_14821);
nand U17868 (N_17868,N_13045,N_14437);
and U17869 (N_17869,N_12840,N_13837);
and U17870 (N_17870,N_14766,N_12080);
or U17871 (N_17871,N_14025,N_14883);
and U17872 (N_17872,N_12265,N_12674);
nor U17873 (N_17873,N_14369,N_12421);
and U17874 (N_17874,N_13669,N_12560);
nand U17875 (N_17875,N_14946,N_14166);
or U17876 (N_17876,N_12831,N_13122);
or U17877 (N_17877,N_13009,N_14889);
xnor U17878 (N_17878,N_14396,N_14096);
nand U17879 (N_17879,N_14837,N_14410);
or U17880 (N_17880,N_14256,N_13177);
and U17881 (N_17881,N_12849,N_12327);
and U17882 (N_17882,N_13893,N_12428);
or U17883 (N_17883,N_12638,N_13264);
nand U17884 (N_17884,N_13788,N_12654);
xor U17885 (N_17885,N_13745,N_14375);
nand U17886 (N_17886,N_14665,N_14191);
or U17887 (N_17887,N_14117,N_14999);
nand U17888 (N_17888,N_12868,N_12930);
nand U17889 (N_17889,N_13114,N_14551);
nand U17890 (N_17890,N_13238,N_12313);
and U17891 (N_17891,N_12766,N_14799);
and U17892 (N_17892,N_14034,N_12511);
or U17893 (N_17893,N_12552,N_13257);
xor U17894 (N_17894,N_12291,N_12801);
or U17895 (N_17895,N_12673,N_14156);
and U17896 (N_17896,N_12391,N_14802);
nand U17897 (N_17897,N_13065,N_14497);
and U17898 (N_17898,N_13190,N_13721);
nor U17899 (N_17899,N_14649,N_12100);
nor U17900 (N_17900,N_14919,N_14719);
and U17901 (N_17901,N_12543,N_13999);
or U17902 (N_17902,N_12427,N_12648);
nand U17903 (N_17903,N_13395,N_14090);
or U17904 (N_17904,N_14020,N_12574);
or U17905 (N_17905,N_14954,N_12847);
or U17906 (N_17906,N_12732,N_13161);
nand U17907 (N_17907,N_13142,N_13949);
xor U17908 (N_17908,N_13270,N_13589);
or U17909 (N_17909,N_12521,N_13427);
and U17910 (N_17910,N_12232,N_13556);
or U17911 (N_17911,N_13210,N_14143);
or U17912 (N_17912,N_12166,N_12423);
nor U17913 (N_17913,N_12935,N_14951);
nand U17914 (N_17914,N_14998,N_12428);
xnor U17915 (N_17915,N_14006,N_13155);
nand U17916 (N_17916,N_12835,N_14861);
or U17917 (N_17917,N_12269,N_13846);
or U17918 (N_17918,N_13716,N_13325);
nor U17919 (N_17919,N_12991,N_12148);
or U17920 (N_17920,N_12827,N_13472);
xnor U17921 (N_17921,N_13484,N_14993);
xor U17922 (N_17922,N_14467,N_12156);
nand U17923 (N_17923,N_12898,N_13720);
nand U17924 (N_17924,N_14803,N_12856);
xnor U17925 (N_17925,N_14680,N_12538);
xnor U17926 (N_17926,N_14619,N_12373);
or U17927 (N_17927,N_13083,N_14605);
nor U17928 (N_17928,N_14239,N_14302);
and U17929 (N_17929,N_13200,N_12003);
and U17930 (N_17930,N_13129,N_14778);
or U17931 (N_17931,N_12605,N_13154);
nor U17932 (N_17932,N_13180,N_13957);
nor U17933 (N_17933,N_12822,N_12326);
xnor U17934 (N_17934,N_14321,N_13273);
nor U17935 (N_17935,N_14900,N_13932);
nor U17936 (N_17936,N_14010,N_13300);
and U17937 (N_17937,N_13367,N_12859);
or U17938 (N_17938,N_12346,N_13935);
nor U17939 (N_17939,N_12712,N_14164);
nor U17940 (N_17940,N_13732,N_14579);
nand U17941 (N_17941,N_12561,N_14383);
xnor U17942 (N_17942,N_12319,N_12087);
nand U17943 (N_17943,N_13975,N_13698);
or U17944 (N_17944,N_12302,N_14442);
and U17945 (N_17945,N_13322,N_12427);
and U17946 (N_17946,N_12690,N_14469);
or U17947 (N_17947,N_12510,N_12935);
and U17948 (N_17948,N_14064,N_14284);
and U17949 (N_17949,N_12705,N_13344);
and U17950 (N_17950,N_12533,N_13602);
nand U17951 (N_17951,N_12959,N_12644);
or U17952 (N_17952,N_14467,N_14893);
and U17953 (N_17953,N_13830,N_13297);
and U17954 (N_17954,N_14083,N_12356);
nand U17955 (N_17955,N_14512,N_12108);
and U17956 (N_17956,N_13939,N_12997);
or U17957 (N_17957,N_13800,N_14151);
or U17958 (N_17958,N_14530,N_12761);
and U17959 (N_17959,N_14711,N_13950);
nand U17960 (N_17960,N_14900,N_14092);
nor U17961 (N_17961,N_12648,N_13613);
and U17962 (N_17962,N_14779,N_14857);
or U17963 (N_17963,N_12575,N_14981);
and U17964 (N_17964,N_13473,N_13507);
nand U17965 (N_17965,N_12050,N_12300);
nand U17966 (N_17966,N_14044,N_13757);
xor U17967 (N_17967,N_14957,N_14173);
or U17968 (N_17968,N_12837,N_14213);
or U17969 (N_17969,N_12856,N_14848);
nand U17970 (N_17970,N_14478,N_12703);
nor U17971 (N_17971,N_12856,N_12695);
nor U17972 (N_17972,N_13315,N_14085);
or U17973 (N_17973,N_12992,N_14373);
or U17974 (N_17974,N_12644,N_13913);
nor U17975 (N_17975,N_12266,N_12530);
nand U17976 (N_17976,N_12689,N_14980);
nor U17977 (N_17977,N_13442,N_14709);
nand U17978 (N_17978,N_14662,N_13424);
nor U17979 (N_17979,N_12597,N_12275);
nor U17980 (N_17980,N_14014,N_13795);
and U17981 (N_17981,N_14481,N_12705);
nand U17982 (N_17982,N_14111,N_13919);
or U17983 (N_17983,N_12849,N_14723);
xor U17984 (N_17984,N_12019,N_13768);
nand U17985 (N_17985,N_13863,N_14324);
nor U17986 (N_17986,N_14043,N_14754);
and U17987 (N_17987,N_13064,N_13426);
nand U17988 (N_17988,N_12578,N_13088);
xor U17989 (N_17989,N_12565,N_14280);
and U17990 (N_17990,N_14280,N_13867);
and U17991 (N_17991,N_14402,N_13705);
and U17992 (N_17992,N_13218,N_14169);
nor U17993 (N_17993,N_12823,N_12785);
and U17994 (N_17994,N_12641,N_12877);
nand U17995 (N_17995,N_12682,N_14161);
nand U17996 (N_17996,N_13043,N_13606);
or U17997 (N_17997,N_12895,N_12490);
and U17998 (N_17998,N_13038,N_13243);
nand U17999 (N_17999,N_13221,N_12440);
nor U18000 (N_18000,N_15325,N_17610);
xor U18001 (N_18001,N_17026,N_15583);
and U18002 (N_18002,N_15605,N_17218);
xor U18003 (N_18003,N_16447,N_16771);
and U18004 (N_18004,N_16528,N_16444);
xnor U18005 (N_18005,N_16638,N_16492);
nor U18006 (N_18006,N_16632,N_15007);
or U18007 (N_18007,N_16039,N_16933);
xor U18008 (N_18008,N_17533,N_17867);
or U18009 (N_18009,N_17875,N_16740);
or U18010 (N_18010,N_17028,N_15611);
nand U18011 (N_18011,N_15627,N_17107);
or U18012 (N_18012,N_15827,N_15271);
and U18013 (N_18013,N_17190,N_15927);
nor U18014 (N_18014,N_16355,N_16089);
or U18015 (N_18015,N_16563,N_15392);
and U18016 (N_18016,N_16366,N_15490);
xnor U18017 (N_18017,N_15242,N_17520);
and U18018 (N_18018,N_16251,N_15130);
xor U18019 (N_18019,N_16195,N_17542);
nand U18020 (N_18020,N_15747,N_17863);
or U18021 (N_18021,N_16892,N_17512);
nor U18022 (N_18022,N_16266,N_17650);
nor U18023 (N_18023,N_17247,N_15525);
or U18024 (N_18024,N_17984,N_16985);
nor U18025 (N_18025,N_17581,N_16363);
and U18026 (N_18026,N_17594,N_17000);
nand U18027 (N_18027,N_17742,N_15069);
or U18028 (N_18028,N_15400,N_17041);
or U18029 (N_18029,N_16412,N_17325);
and U18030 (N_18030,N_16486,N_15235);
and U18031 (N_18031,N_15132,N_17280);
nor U18032 (N_18032,N_17001,N_17705);
or U18033 (N_18033,N_16175,N_17458);
or U18034 (N_18034,N_16243,N_17595);
or U18035 (N_18035,N_15011,N_17873);
or U18036 (N_18036,N_16147,N_15497);
nand U18037 (N_18037,N_15680,N_16280);
and U18038 (N_18038,N_16664,N_17270);
xor U18039 (N_18039,N_16864,N_15214);
xor U18040 (N_18040,N_15879,N_16821);
nand U18041 (N_18041,N_16518,N_16454);
nor U18042 (N_18042,N_15134,N_16644);
xor U18043 (N_18043,N_15360,N_16795);
nor U18044 (N_18044,N_16183,N_17010);
and U18045 (N_18045,N_16799,N_15170);
nand U18046 (N_18046,N_15424,N_16180);
and U18047 (N_18047,N_15893,N_16670);
and U18048 (N_18048,N_16306,N_16205);
nand U18049 (N_18049,N_16372,N_15565);
nor U18050 (N_18050,N_17017,N_15157);
nor U18051 (N_18051,N_17996,N_16860);
xor U18052 (N_18052,N_15390,N_17489);
and U18053 (N_18053,N_17024,N_16559);
and U18054 (N_18054,N_16357,N_16582);
and U18055 (N_18055,N_16718,N_16116);
nand U18056 (N_18056,N_15279,N_17055);
xnor U18057 (N_18057,N_15382,N_15180);
nor U18058 (N_18058,N_17668,N_16449);
nand U18059 (N_18059,N_16055,N_15908);
and U18060 (N_18060,N_15821,N_16904);
and U18061 (N_18061,N_16971,N_17367);
or U18062 (N_18062,N_17663,N_15287);
or U18063 (N_18063,N_16943,N_16703);
nor U18064 (N_18064,N_15707,N_17356);
or U18065 (N_18065,N_15910,N_17661);
xnor U18066 (N_18066,N_17105,N_15362);
and U18067 (N_18067,N_16430,N_16207);
nor U18068 (N_18068,N_15735,N_15898);
or U18069 (N_18069,N_17314,N_15266);
nor U18070 (N_18070,N_17279,N_17108);
nand U18071 (N_18071,N_16513,N_16229);
and U18072 (N_18072,N_15558,N_15272);
nand U18073 (N_18073,N_15010,N_15146);
nor U18074 (N_18074,N_16438,N_16869);
or U18075 (N_18075,N_16035,N_16370);
and U18076 (N_18076,N_15785,N_17069);
nor U18077 (N_18077,N_17008,N_15509);
xnor U18078 (N_18078,N_16717,N_17456);
nand U18079 (N_18079,N_15318,N_16351);
or U18080 (N_18080,N_16396,N_15521);
or U18081 (N_18081,N_15001,N_17540);
nor U18082 (N_18082,N_15819,N_15120);
nor U18083 (N_18083,N_17640,N_15169);
or U18084 (N_18084,N_16191,N_16090);
nor U18085 (N_18085,N_16543,N_15489);
nor U18086 (N_18086,N_17973,N_16930);
and U18087 (N_18087,N_16897,N_17783);
nor U18088 (N_18088,N_17558,N_16509);
and U18089 (N_18089,N_17819,N_16046);
nor U18090 (N_18090,N_17032,N_17119);
or U18091 (N_18091,N_15080,N_15687);
xor U18092 (N_18092,N_16666,N_16157);
nor U18093 (N_18093,N_15957,N_17766);
nor U18094 (N_18094,N_16096,N_17227);
nor U18095 (N_18095,N_15951,N_17543);
or U18096 (N_18096,N_17267,N_15301);
xnor U18097 (N_18097,N_17529,N_17803);
nor U18098 (N_18098,N_17848,N_17160);
xor U18099 (N_18099,N_17934,N_16526);
nand U18100 (N_18100,N_17490,N_15450);
xnor U18101 (N_18101,N_15777,N_17246);
xnor U18102 (N_18102,N_17833,N_17333);
and U18103 (N_18103,N_17158,N_16298);
or U18104 (N_18104,N_15442,N_15637);
and U18105 (N_18105,N_15161,N_17752);
or U18106 (N_18106,N_17004,N_17199);
or U18107 (N_18107,N_15330,N_15966);
or U18108 (N_18108,N_16197,N_17413);
or U18109 (N_18109,N_17449,N_17236);
nand U18110 (N_18110,N_17588,N_17322);
and U18111 (N_18111,N_17198,N_17839);
or U18112 (N_18112,N_17173,N_17619);
and U18113 (N_18113,N_17301,N_17743);
or U18114 (N_18114,N_15028,N_15840);
nor U18115 (N_18115,N_16099,N_17877);
and U18116 (N_18116,N_15111,N_15987);
and U18117 (N_18117,N_16667,N_16552);
nor U18118 (N_18118,N_15800,N_15977);
nand U18119 (N_18119,N_16798,N_15261);
nand U18120 (N_18120,N_17880,N_15173);
or U18121 (N_18121,N_17676,N_15589);
nand U18122 (N_18122,N_16658,N_16735);
nand U18123 (N_18123,N_17541,N_17941);
or U18124 (N_18124,N_17787,N_15776);
and U18125 (N_18125,N_17556,N_17976);
and U18126 (N_18126,N_15705,N_16020);
nand U18127 (N_18127,N_15869,N_15892);
xnor U18128 (N_18128,N_17933,N_16086);
nand U18129 (N_18129,N_17061,N_17336);
xnor U18130 (N_18130,N_16262,N_15665);
xnor U18131 (N_18131,N_15619,N_17254);
nor U18132 (N_18132,N_15854,N_16383);
and U18133 (N_18133,N_15556,N_17185);
xor U18134 (N_18134,N_17259,N_15254);
xor U18135 (N_18135,N_17067,N_15040);
or U18136 (N_18136,N_16271,N_17776);
nor U18137 (N_18137,N_15948,N_17037);
xnor U18138 (N_18138,N_16504,N_15406);
and U18139 (N_18139,N_15181,N_17756);
nor U18140 (N_18140,N_15479,N_17097);
nor U18141 (N_18141,N_15058,N_15522);
nand U18142 (N_18142,N_16053,N_16103);
xnor U18143 (N_18143,N_15802,N_15095);
nand U18144 (N_18144,N_17828,N_15804);
or U18145 (N_18145,N_15575,N_15176);
and U18146 (N_18146,N_16669,N_17011);
nand U18147 (N_18147,N_17256,N_16336);
and U18148 (N_18148,N_15354,N_16401);
or U18149 (N_18149,N_17388,N_15823);
nand U18150 (N_18150,N_17799,N_16219);
xnor U18151 (N_18151,N_17036,N_16810);
nor U18152 (N_18152,N_16951,N_16825);
or U18153 (N_18153,N_15813,N_17746);
and U18154 (N_18154,N_15016,N_16209);
nand U18155 (N_18155,N_15062,N_17870);
and U18156 (N_18156,N_15286,N_16646);
nor U18157 (N_18157,N_15668,N_15784);
xnor U18158 (N_18158,N_16601,N_16373);
nor U18159 (N_18159,N_15002,N_16161);
nand U18160 (N_18160,N_16113,N_17826);
or U18161 (N_18161,N_16312,N_16495);
nand U18162 (N_18162,N_17321,N_15303);
and U18163 (N_18163,N_15013,N_17806);
or U18164 (N_18164,N_17950,N_17044);
nand U18165 (N_18165,N_15876,N_15024);
nor U18166 (N_18166,N_16862,N_16642);
xnor U18167 (N_18167,N_15227,N_17887);
and U18168 (N_18168,N_15328,N_17981);
or U18169 (N_18169,N_15851,N_17441);
nand U18170 (N_18170,N_15061,N_17077);
nor U18171 (N_18171,N_16389,N_16080);
and U18172 (N_18172,N_16142,N_17118);
nor U18173 (N_18173,N_16626,N_16338);
nor U18174 (N_18174,N_15409,N_16101);
and U18175 (N_18175,N_16174,N_15918);
nor U18176 (N_18176,N_15131,N_15493);
nand U18177 (N_18177,N_15604,N_15787);
xor U18178 (N_18178,N_17444,N_16166);
nor U18179 (N_18179,N_15573,N_17644);
and U18180 (N_18180,N_17271,N_17244);
or U18181 (N_18181,N_16696,N_17035);
xor U18182 (N_18182,N_15098,N_17491);
and U18183 (N_18183,N_15774,N_16091);
nand U18184 (N_18184,N_16405,N_15388);
nand U18185 (N_18185,N_17944,N_15515);
nor U18186 (N_18186,N_16540,N_17850);
or U18187 (N_18187,N_15222,N_17514);
nor U18188 (N_18188,N_15794,N_17825);
or U18189 (N_18189,N_16478,N_17946);
or U18190 (N_18190,N_17122,N_17189);
nor U18191 (N_18191,N_17416,N_16094);
and U18192 (N_18192,N_17911,N_16838);
or U18193 (N_18193,N_16006,N_15825);
nor U18194 (N_18194,N_16034,N_15445);
and U18195 (N_18195,N_15306,N_15591);
nand U18196 (N_18196,N_17149,N_16906);
nor U18197 (N_18197,N_15427,N_17781);
and U18198 (N_18198,N_16616,N_17103);
nor U18199 (N_18199,N_16846,N_17398);
or U18200 (N_18200,N_16077,N_17841);
nor U18201 (N_18201,N_16313,N_16952);
or U18202 (N_18202,N_15809,N_16259);
nor U18203 (N_18203,N_15834,N_15398);
and U18204 (N_18204,N_17597,N_15996);
xor U18205 (N_18205,N_16352,N_16177);
nand U18206 (N_18206,N_17862,N_17507);
nor U18207 (N_18207,N_15403,N_15077);
xor U18208 (N_18208,N_16988,N_16976);
and U18209 (N_18209,N_16295,N_16759);
nand U18210 (N_18210,N_16204,N_15249);
nand U18211 (N_18211,N_16571,N_15372);
and U18212 (N_18212,N_17736,N_17019);
and U18213 (N_18213,N_16296,N_15791);
nand U18214 (N_18214,N_15658,N_17229);
nor U18215 (N_18215,N_16932,N_17219);
nand U18216 (N_18216,N_16996,N_17345);
nand U18217 (N_18217,N_16858,N_16480);
nand U18218 (N_18218,N_15965,N_16460);
or U18219 (N_18219,N_15609,N_16138);
nand U18220 (N_18220,N_17616,N_15389);
xor U18221 (N_18221,N_17665,N_16661);
xor U18222 (N_18222,N_15625,N_17224);
or U18223 (N_18223,N_17424,N_16434);
or U18224 (N_18224,N_15128,N_15711);
nor U18225 (N_18225,N_16456,N_16580);
nand U18226 (N_18226,N_17732,N_16765);
nor U18227 (N_18227,N_16467,N_17057);
and U18228 (N_18228,N_16865,N_16607);
or U18229 (N_18229,N_15508,N_16994);
or U18230 (N_18230,N_16645,N_17142);
nand U18231 (N_18231,N_16671,N_17562);
nor U18232 (N_18232,N_17846,N_16514);
nor U18233 (N_18233,N_16049,N_16741);
and U18234 (N_18234,N_17778,N_17276);
nand U18235 (N_18235,N_17673,N_15454);
nor U18236 (N_18236,N_17517,N_15725);
nor U18237 (N_18237,N_16657,N_15381);
and U18238 (N_18238,N_16832,N_16755);
nand U18239 (N_18239,N_17559,N_16800);
or U18240 (N_18240,N_15218,N_17250);
and U18241 (N_18241,N_16889,N_16284);
nor U18242 (N_18242,N_17741,N_16485);
nor U18243 (N_18243,N_15216,N_15968);
and U18244 (N_18244,N_16210,N_15140);
nand U18245 (N_18245,N_15021,N_16446);
or U18246 (N_18246,N_17178,N_17092);
or U18247 (N_18247,N_17920,N_16630);
nand U18248 (N_18248,N_15590,N_15278);
or U18249 (N_18249,N_17786,N_17731);
and U18250 (N_18250,N_16025,N_15596);
xnor U18251 (N_18251,N_17053,N_16767);
and U18252 (N_18252,N_17426,N_16653);
nand U18253 (N_18253,N_17384,N_15566);
and U18254 (N_18254,N_15920,N_17379);
and U18255 (N_18255,N_15849,N_15642);
and U18256 (N_18256,N_16894,N_15672);
nor U18257 (N_18257,N_17411,N_17427);
and U18258 (N_18258,N_17855,N_17241);
nand U18259 (N_18259,N_16005,N_15749);
or U18260 (N_18260,N_16127,N_17547);
and U18261 (N_18261,N_15315,N_15692);
nor U18262 (N_18262,N_16544,N_17994);
or U18263 (N_18263,N_17615,N_15481);
nor U18264 (N_18264,N_16534,N_17740);
or U18265 (N_18265,N_16004,N_15626);
nand U18266 (N_18266,N_15820,N_17470);
nor U18267 (N_18267,N_16967,N_15555);
and U18268 (N_18268,N_16835,N_15344);
or U18269 (N_18269,N_16376,N_15178);
or U18270 (N_18270,N_17265,N_17997);
or U18271 (N_18271,N_17724,N_15171);
nand U18272 (N_18272,N_15729,N_16844);
or U18273 (N_18273,N_17837,N_17085);
and U18274 (N_18274,N_15006,N_17773);
nand U18275 (N_18275,N_16867,N_17425);
nor U18276 (N_18276,N_15934,N_15796);
and U18277 (N_18277,N_15211,N_16065);
nand U18278 (N_18278,N_16409,N_16201);
or U18279 (N_18279,N_17461,N_16359);
or U18280 (N_18280,N_16981,N_17153);
or U18281 (N_18281,N_16947,N_16317);
or U18282 (N_18282,N_15523,N_17194);
or U18283 (N_18283,N_15746,N_17145);
nor U18284 (N_18284,N_16685,N_16304);
or U18285 (N_18285,N_17633,N_15886);
nand U18286 (N_18286,N_17159,N_16712);
nor U18287 (N_18287,N_17370,N_17907);
nor U18288 (N_18288,N_16407,N_17601);
nand U18289 (N_18289,N_16109,N_15505);
and U18290 (N_18290,N_16520,N_16877);
xnor U18291 (N_18291,N_16908,N_15401);
nor U18292 (N_18292,N_16322,N_16707);
xnor U18293 (N_18293,N_17751,N_15004);
nand U18294 (N_18294,N_16564,N_16477);
and U18295 (N_18295,N_17402,N_15338);
and U18296 (N_18296,N_17947,N_17400);
nand U18297 (N_18297,N_16690,N_16168);
xnor U18298 (N_18298,N_16081,N_17910);
and U18299 (N_18299,N_15909,N_17226);
or U18300 (N_18300,N_17523,N_15538);
xnor U18301 (N_18301,N_16746,N_15750);
nor U18302 (N_18302,N_17471,N_16484);
or U18303 (N_18303,N_15663,N_17972);
nand U18304 (N_18304,N_16457,N_16315);
and U18305 (N_18305,N_15488,N_15941);
and U18306 (N_18306,N_17039,N_17078);
or U18307 (N_18307,N_17038,N_17641);
or U18308 (N_18308,N_17928,N_16185);
or U18309 (N_18309,N_17631,N_17963);
xor U18310 (N_18310,N_17366,N_15017);
or U18311 (N_18311,N_15913,N_16292);
xor U18312 (N_18312,N_16387,N_16935);
nor U18313 (N_18313,N_17729,N_16682);
or U18314 (N_18314,N_16772,N_16708);
nor U18315 (N_18315,N_15858,N_15230);
nor U18316 (N_18316,N_15789,N_16382);
nand U18317 (N_18317,N_16057,N_17094);
nand U18318 (N_18318,N_15081,N_15906);
and U18319 (N_18319,N_16913,N_15492);
and U18320 (N_18320,N_17175,N_15105);
or U18321 (N_18321,N_16870,N_15340);
nor U18322 (N_18322,N_16018,N_16303);
xnor U18323 (N_18323,N_16036,N_15929);
nand U18324 (N_18324,N_16915,N_15086);
and U18325 (N_18325,N_15498,N_17062);
and U18326 (N_18326,N_17669,N_17580);
nand U18327 (N_18327,N_16538,N_16165);
nor U18328 (N_18328,N_15195,N_15981);
xor U18329 (N_18329,N_17027,N_17790);
nand U18330 (N_18330,N_17454,N_16794);
and U18331 (N_18331,N_16074,N_17434);
or U18332 (N_18332,N_17701,N_16960);
nand U18333 (N_18333,N_16662,N_16880);
or U18334 (N_18334,N_15548,N_15032);
or U18335 (N_18335,N_16660,N_16546);
and U18336 (N_18336,N_17999,N_16061);
nor U18337 (N_18337,N_15598,N_15666);
nor U18338 (N_18338,N_15837,N_17304);
and U18339 (N_18339,N_15363,N_15064);
and U18340 (N_18340,N_15262,N_15563);
nor U18341 (N_18341,N_16128,N_17212);
or U18342 (N_18342,N_16419,N_17674);
and U18343 (N_18343,N_17252,N_16997);
and U18344 (N_18344,N_17283,N_17769);
nor U18345 (N_18345,N_16882,N_16143);
or U18346 (N_18346,N_16631,N_15138);
nand U18347 (N_18347,N_15654,N_15615);
nand U18348 (N_18348,N_15686,N_15894);
and U18349 (N_18349,N_15978,N_16819);
and U18350 (N_18350,N_16406,N_17853);
xnor U18351 (N_18351,N_16170,N_17086);
and U18352 (N_18352,N_16737,N_16466);
and U18353 (N_18353,N_16393,N_17912);
and U18354 (N_18354,N_16745,N_17221);
nor U18355 (N_18355,N_15135,N_17504);
xor U18356 (N_18356,N_17519,N_17628);
nor U18357 (N_18357,N_15712,N_16663);
or U18358 (N_18358,N_16784,N_17792);
xnor U18359 (N_18359,N_17180,N_17613);
and U18360 (N_18360,N_15585,N_17445);
nand U18361 (N_18361,N_17121,N_15925);
nand U18362 (N_18362,N_16610,N_16624);
or U18363 (N_18363,N_17621,N_15145);
or U18364 (N_18364,N_16803,N_17710);
or U18365 (N_18365,N_16443,N_15453);
nor U18366 (N_18366,N_16367,N_17156);
nand U18367 (N_18367,N_16069,N_16151);
and U18368 (N_18368,N_17550,N_16278);
nor U18369 (N_18369,N_16714,N_17524);
nand U18370 (N_18370,N_17515,N_17191);
or U18371 (N_18371,N_16876,N_16008);
or U18372 (N_18372,N_15501,N_15539);
and U18373 (N_18373,N_15190,N_16182);
xnor U18374 (N_18374,N_16744,N_15467);
nor U18375 (N_18375,N_17587,N_15477);
or U18376 (N_18376,N_15592,N_15434);
or U18377 (N_18377,N_17312,N_17734);
and U18378 (N_18378,N_17483,N_16250);
nor U18379 (N_18379,N_17949,N_16026);
nor U18380 (N_18380,N_17805,N_16426);
nand U18381 (N_18381,N_16600,N_15352);
nor U18382 (N_18382,N_17840,N_15265);
nand U18383 (N_18383,N_16281,N_15657);
nor U18384 (N_18384,N_16796,N_15150);
and U18385 (N_18385,N_17137,N_17617);
and U18386 (N_18386,N_16581,N_16112);
and U18387 (N_18387,N_16169,N_16340);
xnor U18388 (N_18388,N_17930,N_17048);
nand U18389 (N_18389,N_15659,N_17022);
xnor U18390 (N_18390,N_15034,N_15056);
nand U18391 (N_18391,N_16684,N_16288);
or U18392 (N_18392,N_15418,N_16458);
or U18393 (N_18393,N_17498,N_16321);
nor U18394 (N_18394,N_17744,N_16102);
nand U18395 (N_18395,N_17087,N_16156);
or U18396 (N_18396,N_17624,N_16299);
nand U18397 (N_18397,N_16589,N_17808);
or U18398 (N_18398,N_16872,N_15865);
nand U18399 (N_18399,N_17390,N_16941);
and U18400 (N_18400,N_15194,N_16378);
and U18401 (N_18401,N_15755,N_17553);
nand U18402 (N_18402,N_16959,N_15739);
nand U18403 (N_18403,N_17856,N_17249);
xnor U18404 (N_18404,N_17438,N_17147);
nor U18405 (N_18405,N_15970,N_17653);
and U18406 (N_18406,N_17374,N_15387);
xnor U18407 (N_18407,N_17866,N_15250);
or U18408 (N_18408,N_15859,N_16989);
nor U18409 (N_18409,N_15644,N_15507);
or U18410 (N_18410,N_17109,N_17832);
nand U18411 (N_18411,N_17295,N_16539);
xor U18412 (N_18412,N_16792,N_17623);
and U18413 (N_18413,N_15166,N_17054);
or U18414 (N_18414,N_16119,N_16731);
and U18415 (N_18415,N_16476,N_17499);
nor U18416 (N_18416,N_15866,N_16859);
and U18417 (N_18417,N_17914,N_17754);
nand U18418 (N_18418,N_16747,N_15989);
nor U18419 (N_18419,N_16473,N_15233);
nand U18420 (N_18420,N_15843,N_15206);
or U18421 (N_18421,N_17956,N_17719);
or U18422 (N_18422,N_16542,N_16963);
nand U18423 (N_18423,N_16318,N_15950);
nor U18424 (N_18424,N_15341,N_15149);
nand U18425 (N_18425,N_15133,N_16845);
and U18426 (N_18426,N_15332,N_17566);
and U18427 (N_18427,N_15737,N_15196);
and U18428 (N_18428,N_17117,N_17365);
nor U18429 (N_18429,N_17404,N_15026);
nand U18430 (N_18430,N_16075,N_17788);
or U18431 (N_18431,N_15917,N_16556);
nor U18432 (N_18432,N_17183,N_17363);
nand U18433 (N_18433,N_16071,N_16834);
or U18434 (N_18434,N_17590,N_17859);
nor U18435 (N_18435,N_15848,N_15482);
or U18436 (N_18436,N_17392,N_17484);
and U18437 (N_18437,N_15667,N_16385);
nand U18438 (N_18438,N_16399,N_17018);
and U18439 (N_18439,N_16045,N_16962);
nand U18440 (N_18440,N_16087,N_16332);
nand U18441 (N_18441,N_16381,N_16585);
nor U18442 (N_18442,N_16417,N_15259);
nand U18443 (N_18443,N_17687,N_15736);
nand U18444 (N_18444,N_16983,N_15972);
nand U18445 (N_18445,N_16519,N_17935);
nor U18446 (N_18446,N_15048,N_17785);
or U18447 (N_18447,N_15901,N_17899);
and U18448 (N_18448,N_17273,N_15374);
nand U18449 (N_18449,N_15610,N_15142);
and U18450 (N_18450,N_16788,N_17937);
nand U18451 (N_18451,N_16415,N_15309);
nand U18452 (N_18452,N_17381,N_15769);
nand U18453 (N_18453,N_17962,N_17480);
nand U18454 (N_18454,N_15714,N_17612);
and U18455 (N_18455,N_17591,N_17154);
and U18456 (N_18456,N_15480,N_17535);
or U18457 (N_18457,N_17764,N_17672);
and U18458 (N_18458,N_17992,N_16541);
nand U18459 (N_18459,N_16629,N_16575);
and U18460 (N_18460,N_16124,N_15179);
nand U18461 (N_18461,N_15393,N_15203);
nor U18462 (N_18462,N_15386,N_15472);
xor U18463 (N_18463,N_16354,N_16294);
nor U18464 (N_18464,N_17182,N_17327);
nand U18465 (N_18465,N_16905,N_17263);
nor U18466 (N_18466,N_16612,N_15455);
nand U18467 (N_18467,N_16608,N_16676);
nor U18468 (N_18468,N_16625,N_15762);
nor U18469 (N_18469,N_16452,N_16380);
xnor U18470 (N_18470,N_16293,N_16475);
nor U18471 (N_18471,N_16153,N_15616);
and U18472 (N_18472,N_15009,N_16672);
and U18473 (N_18473,N_15108,N_16900);
nand U18474 (N_18474,N_15991,N_17380);
nand U18475 (N_18475,N_17407,N_16011);
nand U18476 (N_18476,N_16070,N_17371);
nand U18477 (N_18477,N_16568,N_15655);
nand U18478 (N_18478,N_17686,N_16890);
nand U18479 (N_18479,N_16141,N_17251);
nand U18480 (N_18480,N_16029,N_15955);
nand U18481 (N_18481,N_17305,N_15810);
xor U18482 (N_18482,N_17487,N_15973);
nor U18483 (N_18483,N_16936,N_16085);
or U18484 (N_18484,N_16469,N_15995);
or U18485 (N_18485,N_17917,N_15246);
nand U18486 (N_18486,N_15877,N_15432);
nand U18487 (N_18487,N_15188,N_15491);
nor U18488 (N_18488,N_15109,N_17780);
xnor U18489 (N_18489,N_15676,N_15121);
nor U18490 (N_18490,N_16993,N_17029);
and U18491 (N_18491,N_17485,N_17376);
nand U18492 (N_18492,N_17217,N_15413);
and U18493 (N_18493,N_17261,N_15158);
or U18494 (N_18494,N_16488,N_17353);
and U18495 (N_18495,N_17155,N_16275);
and U18496 (N_18496,N_17608,N_15051);
or U18497 (N_18497,N_16948,N_16232);
or U18498 (N_18498,N_16896,N_17135);
nor U18499 (N_18499,N_17702,N_17794);
nand U18500 (N_18500,N_16374,N_16964);
and U18501 (N_18501,N_16565,N_16957);
nor U18502 (N_18502,N_17106,N_16365);
or U18503 (N_18503,N_15961,N_17339);
nand U18504 (N_18504,N_16384,N_15231);
or U18505 (N_18505,N_15027,N_15148);
nor U18506 (N_18506,N_17014,N_17372);
xor U18507 (N_18507,N_15461,N_17889);
nand U18508 (N_18508,N_15815,N_17927);
nand U18509 (N_18509,N_17481,N_15457);
or U18510 (N_18510,N_16961,N_17496);
or U18511 (N_18511,N_16748,N_15473);
and U18512 (N_18512,N_16200,N_16940);
and U18513 (N_18513,N_17288,N_17876);
nand U18514 (N_18514,N_16269,N_15500);
and U18515 (N_18515,N_15225,N_16335);
and U18516 (N_18516,N_17294,N_17095);
and U18517 (N_18517,N_17609,N_15838);
nor U18518 (N_18518,N_15656,N_16028);
and U18519 (N_18519,N_17651,N_17505);
nand U18520 (N_18520,N_15940,N_15074);
xnor U18521 (N_18521,N_15041,N_17569);
and U18522 (N_18522,N_16290,N_15971);
and U18523 (N_18523,N_15759,N_17648);
and U18524 (N_18524,N_16463,N_16598);
nor U18525 (N_18525,N_15799,N_16902);
and U18526 (N_18526,N_16573,N_17486);
nor U18527 (N_18527,N_17300,N_17688);
xor U18528 (N_18528,N_16781,N_16211);
nor U18529 (N_18529,N_17412,N_15976);
and U18530 (N_18530,N_15175,N_15685);
nor U18531 (N_18531,N_17695,N_15648);
and U18532 (N_18532,N_16263,N_16595);
or U18533 (N_18533,N_17214,N_15650);
nand U18534 (N_18534,N_16618,N_16358);
nor U18535 (N_18535,N_15209,N_15559);
and U18536 (N_18536,N_15740,N_17045);
or U18537 (N_18537,N_16802,N_15471);
or U18538 (N_18538,N_15752,N_17638);
nand U18539 (N_18539,N_17891,N_16226);
and U18540 (N_18540,N_17838,N_15914);
nand U18541 (N_18541,N_16193,N_15285);
or U18542 (N_18542,N_17269,N_16079);
nand U18543 (N_18543,N_15545,N_15783);
nand U18544 (N_18544,N_15806,N_16007);
or U18545 (N_18545,N_17552,N_16786);
nor U18546 (N_18546,N_16909,N_15669);
nand U18547 (N_18547,N_15094,N_16939);
or U18548 (N_18548,N_17671,N_16686);
xnor U18549 (N_18549,N_16235,N_16809);
xor U18550 (N_18550,N_16596,N_16522);
or U18551 (N_18551,N_17429,N_17448);
nand U18552 (N_18552,N_17316,N_17330);
nand U18553 (N_18553,N_17723,N_15839);
nor U18554 (N_18554,N_16000,N_16041);
or U18555 (N_18555,N_15606,N_17549);
nor U18556 (N_18556,N_17871,N_15738);
nand U18557 (N_18557,N_15417,N_16246);
xnor U18558 (N_18558,N_16619,N_15091);
and U18559 (N_18559,N_17532,N_16054);
and U18560 (N_18560,N_17664,N_16056);
or U18561 (N_18561,N_16349,N_17816);
xor U18562 (N_18562,N_16603,N_17652);
and U18563 (N_18563,N_15113,N_17422);
nand U18564 (N_18564,N_15571,N_15316);
and U18565 (N_18565,N_15141,N_15293);
or U18566 (N_18566,N_16181,N_16224);
nor U18567 (N_18567,N_17457,N_17500);
or U18568 (N_18568,N_16532,N_15517);
xor U18569 (N_18569,N_15574,N_16030);
nand U18570 (N_18570,N_17771,N_15456);
and U18571 (N_18571,N_15770,N_16023);
xnor U18572 (N_18572,N_17302,N_15295);
and U18573 (N_18573,N_17451,N_15552);
and U18574 (N_18574,N_17111,N_16445);
nand U18575 (N_18575,N_16888,N_17768);
nand U18576 (N_18576,N_15629,N_15673);
and U18577 (N_18577,N_17796,N_16885);
nor U18578 (N_18578,N_15294,N_16377);
nand U18579 (N_18579,N_15063,N_16010);
and U18580 (N_18580,N_17123,N_15678);
and U18581 (N_18581,N_17459,N_15767);
nor U18582 (N_18582,N_15670,N_15014);
or U18583 (N_18583,N_15347,N_16946);
xor U18584 (N_18584,N_15912,N_16950);
and U18585 (N_18585,N_17923,N_15535);
or U18586 (N_18586,N_17394,N_17146);
and U18587 (N_18587,N_15369,N_17116);
or U18588 (N_18588,N_15857,N_17073);
or U18589 (N_18589,N_16145,N_15323);
nand U18590 (N_18590,N_16068,N_15057);
nor U18591 (N_18591,N_16032,N_15775);
and U18592 (N_18592,N_15734,N_15284);
xor U18593 (N_18593,N_16945,N_16360);
nor U18594 (N_18594,N_17238,N_15071);
nor U18595 (N_18595,N_15743,N_16258);
nor U18596 (N_18596,N_15412,N_15334);
nand U18597 (N_18597,N_16098,N_16789);
and U18598 (N_18598,N_15942,N_17593);
and U18599 (N_18599,N_15828,N_16697);
or U18600 (N_18600,N_15617,N_17681);
nand U18601 (N_18601,N_17240,N_15786);
and U18602 (N_18602,N_17278,N_16841);
nand U18603 (N_18603,N_16031,N_17222);
nor U18604 (N_18604,N_16929,N_16024);
nand U18605 (N_18605,N_17636,N_16436);
and U18606 (N_18606,N_16451,N_16561);
nand U18607 (N_18607,N_16190,N_17675);
nand U18608 (N_18608,N_16852,N_15296);
xnor U18609 (N_18609,N_17174,N_17760);
nand U18610 (N_18610,N_17967,N_16461);
nand U18611 (N_18611,N_17344,N_15537);
or U18612 (N_18612,N_17980,N_15751);
or U18613 (N_18613,N_17555,N_17645);
and U18614 (N_18614,N_15102,N_15460);
xor U18615 (N_18615,N_17319,N_15329);
nand U18616 (N_18616,N_15554,N_15870);
and U18617 (N_18617,N_17823,N_17656);
nand U18618 (N_18618,N_16678,N_16154);
nand U18619 (N_18619,N_17357,N_17013);
nor U18620 (N_18620,N_16198,N_17296);
or U18621 (N_18621,N_16255,N_15012);
nor U18622 (N_18622,N_15671,N_17310);
and U18623 (N_18623,N_16404,N_16924);
and U18624 (N_18624,N_16493,N_15862);
nand U18625 (N_18625,N_17245,N_15724);
nand U18626 (N_18626,N_15983,N_16325);
nand U18627 (N_18627,N_15576,N_15217);
xor U18628 (N_18628,N_17307,N_15029);
or U18629 (N_18629,N_16826,N_17083);
nor U18630 (N_18630,N_17931,N_16766);
or U18631 (N_18631,N_16713,N_15070);
xor U18632 (N_18632,N_16414,N_16136);
or U18633 (N_18633,N_17753,N_17443);
and U18634 (N_18634,N_17034,N_16769);
nand U18635 (N_18635,N_15832,N_15969);
and U18636 (N_18636,N_17757,N_17739);
or U18637 (N_18637,N_16824,N_16044);
nand U18638 (N_18638,N_16973,N_15486);
nand U18639 (N_18639,N_17205,N_17409);
nand U18640 (N_18640,N_15582,N_15599);
or U18641 (N_18641,N_15385,N_16857);
nand U18642 (N_18642,N_16591,N_15847);
or U18643 (N_18643,N_15201,N_17058);
nand U18644 (N_18644,N_16337,N_15924);
nor U18645 (N_18645,N_16705,N_17802);
and U18646 (N_18646,N_15088,N_16059);
or U18647 (N_18647,N_15115,N_17797);
and U18648 (N_18648,N_16225,N_15163);
nand U18649 (N_18649,N_15706,N_16562);
nor U18650 (N_18650,N_17810,N_16222);
nor U18651 (N_18651,N_15634,N_15238);
and U18652 (N_18652,N_16550,N_16027);
and U18653 (N_18653,N_15241,N_15496);
and U18654 (N_18654,N_17368,N_16777);
nand U18655 (N_18655,N_15760,N_15139);
and U18656 (N_18656,N_17358,N_17176);
or U18657 (N_18657,N_16881,N_16987);
and U18658 (N_18658,N_16578,N_15540);
or U18659 (N_18659,N_17925,N_15561);
or U18660 (N_18660,N_15090,N_17157);
and U18661 (N_18661,N_17986,N_15232);
nor U18662 (N_18662,N_15485,N_16060);
nand U18663 (N_18663,N_16428,N_17005);
xor U18664 (N_18664,N_16273,N_16289);
nand U18665 (N_18665,N_15874,N_15407);
or U18666 (N_18666,N_15727,N_15184);
or U18667 (N_18667,N_16613,N_17355);
and U18668 (N_18668,N_15584,N_16464);
nand U18669 (N_18669,N_16974,N_15549);
nor U18670 (N_18670,N_15930,N_16651);
nand U18671 (N_18671,N_15159,N_17204);
and U18672 (N_18672,N_15059,N_17258);
xnor U18673 (N_18673,N_17632,N_16196);
nand U18674 (N_18674,N_15376,N_17530);
and U18675 (N_18675,N_15204,N_17618);
nor U18676 (N_18676,N_17346,N_15975);
or U18677 (N_18677,N_15274,N_17905);
nand U18678 (N_18678,N_15322,N_17908);
or U18679 (N_18679,N_15005,N_15962);
nor U18680 (N_18680,N_15939,N_16206);
nor U18681 (N_18681,N_17306,N_17959);
or U18682 (N_18682,N_17290,N_15337);
nand U18683 (N_18683,N_17033,N_16627);
nor U18684 (N_18684,N_16758,N_15185);
and U18685 (N_18685,N_15137,N_16743);
and U18686 (N_18686,N_16978,N_17161);
nand U18687 (N_18687,N_17080,N_16931);
and U18688 (N_18688,N_15875,N_16115);
or U18689 (N_18689,N_15364,N_17059);
nor U18690 (N_18690,N_17639,N_17919);
and U18691 (N_18691,N_15361,N_16634);
or U18692 (N_18692,N_17679,N_15156);
nor U18693 (N_18693,N_17395,N_15431);
nand U18694 (N_18694,N_17172,N_16536);
nand U18695 (N_18695,N_15885,N_16330);
nand U18696 (N_18696,N_16435,N_15199);
nand U18697 (N_18697,N_16328,N_15436);
or U18698 (N_18698,N_16455,N_16511);
or U18699 (N_18699,N_16067,N_15635);
or U18700 (N_18700,N_16652,N_16868);
nor U18701 (N_18701,N_17707,N_17466);
or U18702 (N_18702,N_17228,N_17408);
or U18703 (N_18703,N_15822,N_17942);
and U18704 (N_18704,N_16639,N_16602);
nand U18705 (N_18705,N_15256,N_15160);
or U18706 (N_18706,N_16347,N_16604);
xnor U18707 (N_18707,N_17938,N_16064);
nor U18708 (N_18708,N_16261,N_16567);
nor U18709 (N_18709,N_15331,N_16621);
or U18710 (N_18710,N_16817,N_17909);
or U18711 (N_18711,N_15990,N_15420);
or U18712 (N_18712,N_17560,N_16131);
nor U18713 (N_18713,N_15623,N_16920);
nand U18714 (N_18714,N_17446,N_17521);
nand U18715 (N_18715,N_17488,N_16052);
nor U18716 (N_18716,N_16609,N_15551);
nor U18717 (N_18717,N_16503,N_17264);
and U18718 (N_18718,N_15757,N_17405);
or U18719 (N_18719,N_17475,N_17298);
nor U18720 (N_18720,N_17577,N_16572);
and U18721 (N_18721,N_16228,N_15411);
nand U18722 (N_18722,N_15607,N_15647);
or U18723 (N_18723,N_15495,N_17065);
nor U18724 (N_18724,N_15154,N_16213);
and U18725 (N_18725,N_16139,N_16411);
and U18726 (N_18726,N_16848,N_17579);
and U18727 (N_18727,N_15096,N_15536);
nor U18728 (N_18728,N_16287,N_17913);
and U18729 (N_18729,N_17012,N_17793);
nand U18730 (N_18730,N_16242,N_17704);
and U18731 (N_18731,N_17574,N_15100);
nor U18732 (N_18732,N_17534,N_15778);
or U18733 (N_18733,N_17557,N_15855);
nor U18734 (N_18734,N_17737,N_17148);
and U18735 (N_18735,N_15985,N_16732);
and U18736 (N_18736,N_16734,N_17351);
and U18737 (N_18737,N_15192,N_15674);
nor U18738 (N_18738,N_17572,N_15503);
or U18739 (N_18739,N_15314,N_16855);
or U18740 (N_18740,N_15856,N_17334);
and U18741 (N_18741,N_16106,N_17337);
nand U18742 (N_18742,N_15816,N_17326);
and U18743 (N_18743,N_15689,N_17755);
nand U18744 (N_18744,N_15476,N_17983);
nor U18745 (N_18745,N_16728,N_17452);
and U18746 (N_18746,N_16914,N_16736);
or U18747 (N_18747,N_16309,N_16082);
nand U18748 (N_18748,N_16083,N_15888);
nor U18749 (N_18749,N_16334,N_15097);
xnor U18750 (N_18750,N_15075,N_16674);
xor U18751 (N_18751,N_15652,N_15891);
nor U18752 (N_18752,N_16992,N_16216);
nand U18753 (N_18753,N_17952,N_16977);
nand U18754 (N_18754,N_15000,N_16108);
and U18755 (N_18755,N_17099,N_15311);
nor U18756 (N_18756,N_15038,N_15541);
nor U18757 (N_18757,N_15949,N_15391);
xnor U18758 (N_18758,N_17511,N_17343);
and U18759 (N_18759,N_16129,N_16346);
or U18760 (N_18760,N_16729,N_17501);
or U18761 (N_18761,N_17043,N_16413);
nor U18762 (N_18762,N_15126,N_15569);
and U18763 (N_18763,N_17655,N_17926);
and U18764 (N_18764,N_17139,N_16570);
and U18765 (N_18765,N_16711,N_16958);
nand U18766 (N_18766,N_15353,N_16291);
nor U18767 (N_18767,N_17396,N_15107);
and U18768 (N_18768,N_17361,N_16822);
nand U18769 (N_18769,N_15220,N_17076);
nand U18770 (N_18770,N_16923,N_17722);
nor U18771 (N_18771,N_17009,N_16342);
xnor U18772 (N_18772,N_16017,N_15694);
nand U18773 (N_18773,N_17406,N_15730);
or U18774 (N_18774,N_15164,N_15550);
nor U18775 (N_18775,N_16012,N_16423);
nand U18776 (N_18776,N_17260,N_16866);
nor U18777 (N_18777,N_15974,N_17684);
nand U18778 (N_18778,N_16706,N_17421);
and U18779 (N_18779,N_16353,N_15622);
nor U18780 (N_18780,N_15186,N_16212);
or U18781 (N_18781,N_17385,N_17063);
or U18782 (N_18782,N_15722,N_15421);
nand U18783 (N_18783,N_15880,N_15979);
or U18784 (N_18784,N_15720,N_16260);
and U18785 (N_18785,N_17266,N_17694);
nor U18786 (N_18786,N_15543,N_15698);
nor U18787 (N_18787,N_15719,N_15597);
or U18788 (N_18788,N_17888,N_15326);
nand U18789 (N_18789,N_15753,N_17626);
xor U18790 (N_18790,N_15008,N_15527);
nor U18791 (N_18791,N_16331,N_17373);
nand U18792 (N_18792,N_16853,N_17382);
and U18793 (N_18793,N_17829,N_16254);
nand U18794 (N_18794,N_16237,N_16301);
nand U18795 (N_18795,N_15082,N_16348);
nor U18796 (N_18796,N_15905,N_17031);
and U18797 (N_18797,N_17678,N_16150);
nor U18798 (N_18798,N_15465,N_17812);
nand U18799 (N_18799,N_15696,N_16675);
nor U18800 (N_18800,N_16548,N_15405);
nor U18801 (N_18801,N_15452,N_15302);
nor U18802 (N_18802,N_15036,N_17800);
nand U18803 (N_18803,N_15359,N_16763);
nand U18804 (N_18804,N_17433,N_16163);
nand U18805 (N_18805,N_16110,N_16648);
or U18806 (N_18806,N_17614,N_16042);
xor U18807 (N_18807,N_16040,N_15697);
xor U18808 (N_18808,N_15531,N_17255);
and U18809 (N_18809,N_16450,N_17822);
and U18810 (N_18810,N_15127,N_16779);
and U18811 (N_18811,N_16531,N_15494);
or U18812 (N_18812,N_15922,N_17893);
nand U18813 (N_18813,N_17169,N_16323);
xor U18814 (N_18814,N_16785,N_15812);
and U18815 (N_18815,N_16551,N_17528);
nand U18816 (N_18816,N_17857,N_17629);
or U18817 (N_18817,N_16773,N_15723);
nor U18818 (N_18818,N_17332,N_15844);
and U18819 (N_18819,N_16341,N_17971);
or U18820 (N_18820,N_15200,N_16019);
nand U18821 (N_18821,N_15771,N_17081);
or U18822 (N_18822,N_17021,N_15933);
and U18823 (N_18823,N_17918,N_15093);
or U18824 (N_18824,N_16283,N_16938);
nor U18825 (N_18825,N_17197,N_16680);
and U18826 (N_18826,N_15076,N_16202);
and U18827 (N_18827,N_17758,N_17397);
or U18828 (N_18828,N_17845,N_17943);
or U18829 (N_18829,N_15954,N_15754);
nor U18830 (N_18830,N_17220,N_15700);
nand U18831 (N_18831,N_15470,N_15240);
or U18832 (N_18832,N_17020,N_16424);
and U18833 (N_18833,N_17242,N_16831);
or U18834 (N_18834,N_16368,N_17921);
nand U18835 (N_18835,N_15110,N_16919);
or U18836 (N_18836,N_17717,N_16649);
nand U18837 (N_18837,N_17939,N_15884);
or U18838 (N_18838,N_16267,N_17414);
and U18839 (N_18839,N_16021,N_17874);
nand U18840 (N_18840,N_16517,N_16244);
or U18841 (N_18841,N_15921,N_16107);
or U18842 (N_18842,N_17463,N_15520);
or U18843 (N_18843,N_16907,N_17464);
and U18844 (N_18844,N_15683,N_17210);
xor U18845 (N_18845,N_15443,N_16566);
or U18846 (N_18846,N_15620,N_17088);
nand U18847 (N_18847,N_16956,N_17733);
or U18848 (N_18848,N_17884,N_15395);
and U18849 (N_18849,N_15383,N_16879);
or U18850 (N_18850,N_17584,N_16916);
nand U18851 (N_18851,N_16910,N_16236);
or U18852 (N_18852,N_16972,N_16816);
nor U18853 (N_18853,N_17186,N_15451);
nand U18854 (N_18854,N_16557,N_15861);
and U18855 (N_18855,N_15852,N_15675);
nand U18856 (N_18856,N_15084,N_15277);
or U18857 (N_18857,N_16327,N_15144);
nand U18858 (N_18858,N_17383,N_17082);
nand U18859 (N_18859,N_15860,N_16489);
xnor U18860 (N_18860,N_15643,N_15043);
nand U18861 (N_18861,N_16474,N_16847);
nor U18862 (N_18862,N_16078,N_15936);
and U18863 (N_18863,N_17418,N_16234);
nor U18864 (N_18864,N_15718,N_17565);
and U18865 (N_18865,N_17974,N_15679);
or U18866 (N_18866,N_16814,N_16130);
and U18867 (N_18867,N_16203,N_17127);
nor U18868 (N_18868,N_15346,N_15928);
xnor U18869 (N_18869,N_15474,N_17209);
and U18870 (N_18870,N_16084,N_15304);
xor U18871 (N_18871,N_17901,N_16668);
xnor U18872 (N_18872,N_16537,N_17750);
nor U18873 (N_18873,N_15267,N_17620);
nor U18874 (N_18874,N_15958,N_16586);
or U18875 (N_18875,N_15684,N_17084);
nand U18876 (N_18876,N_15189,N_15817);
nand U18877 (N_18877,N_16775,N_15484);
and U18878 (N_18878,N_17328,N_16453);
or U18879 (N_18879,N_17435,N_17842);
and U18880 (N_18880,N_17399,N_15276);
nand U18881 (N_18881,N_17213,N_16727);
and U18882 (N_18882,N_16693,N_17936);
nand U18883 (N_18883,N_15899,N_16874);
nand U18884 (N_18884,N_15365,N_16953);
nand U18885 (N_18885,N_16527,N_17852);
and U18886 (N_18886,N_16326,N_15695);
nand U18887 (N_18887,N_17342,N_17450);
or U18888 (N_18888,N_16599,N_17975);
xnor U18889 (N_18889,N_15378,N_17125);
nor U18890 (N_18890,N_16158,N_17243);
or U18891 (N_18891,N_16037,N_16375);
nand U18892 (N_18892,N_17347,N_15292);
and U18893 (N_18893,N_15602,N_17195);
nor U18894 (N_18894,N_16369,N_16022);
and U18895 (N_18895,N_16553,N_17714);
nand U18896 (N_18896,N_16698,N_16220);
or U18897 (N_18897,N_17320,N_17537);
or U18898 (N_18898,N_15324,N_17257);
nand U18899 (N_18899,N_17352,N_16014);
nand U18900 (N_18900,N_16683,N_16521);
nor U18901 (N_18901,N_17728,N_16710);
and U18902 (N_18902,N_16233,N_15018);
nor U18903 (N_18903,N_17978,N_17492);
nand U18904 (N_18904,N_15601,N_16949);
and U18905 (N_18905,N_17948,N_17090);
and U18906 (N_18906,N_15464,N_16757);
nor U18907 (N_18907,N_15313,N_15356);
and U18908 (N_18908,N_17847,N_15380);
or U18909 (N_18909,N_16215,N_15741);
nand U18910 (N_18910,N_15570,N_16873);
xnor U18911 (N_18911,N_15136,N_17932);
or U18912 (N_18912,N_15693,N_15044);
or U18913 (N_18913,N_15513,N_15068);
or U18914 (N_18914,N_16754,N_16937);
nor U18915 (N_18915,N_17115,N_15568);
nand U18916 (N_18916,N_15245,N_15841);
and U18917 (N_18917,N_17713,N_16167);
and U18918 (N_18918,N_16836,N_17813);
nand U18919 (N_18919,N_15833,N_15066);
xor U18920 (N_18920,N_15052,N_16015);
nor U18921 (N_18921,N_15980,N_17896);
nor U18922 (N_18922,N_17696,N_16230);
xor U18923 (N_18923,N_15312,N_17954);
nand U18924 (N_18924,N_17364,N_17430);
or U18925 (N_18925,N_15015,N_15191);
or U18926 (N_18926,N_17275,N_16724);
nand U18927 (N_18927,N_17046,N_15953);
nand U18928 (N_18928,N_16525,N_17166);
nor U18929 (N_18929,N_15618,N_16410);
or U18930 (N_18930,N_15628,N_15904);
xor U18931 (N_18931,N_16679,N_15193);
nand U18932 (N_18932,N_16922,N_15943);
nand U18933 (N_18933,N_17977,N_17789);
or U18934 (N_18934,N_17814,N_16465);
nor U18935 (N_18935,N_16545,N_16583);
xor U18936 (N_18936,N_17253,N_15524);
nor U18937 (N_18937,N_15197,N_17795);
nor U18938 (N_18938,N_15257,N_17235);
or U18939 (N_18939,N_16726,N_15042);
or U18940 (N_18940,N_16188,N_15305);
nor U18941 (N_18941,N_17469,N_15600);
nand U18942 (N_18942,N_15699,N_16491);
nor U18943 (N_18943,N_17827,N_17649);
and U18944 (N_18944,N_17292,N_16605);
and U18945 (N_18945,N_15728,N_16427);
nor U18946 (N_18946,N_15483,N_16975);
nand U18947 (N_18947,N_16482,N_17101);
or U18948 (N_18948,N_17985,N_17465);
or U18949 (N_18949,N_16628,N_16100);
xnor U18950 (N_18950,N_17582,N_17362);
nor U18951 (N_18951,N_17583,N_15049);
or U18952 (N_18952,N_17970,N_17677);
and U18953 (N_18953,N_17879,N_17646);
nor U18954 (N_18954,N_15506,N_15662);
nand U18955 (N_18955,N_16155,N_15152);
and U18956 (N_18956,N_17303,N_17890);
nor U18957 (N_18957,N_17144,N_15247);
and U18958 (N_18958,N_16665,N_17460);
nand U18959 (N_18959,N_15682,N_15544);
or U18960 (N_18960,N_17341,N_15404);
or U18961 (N_18961,N_16811,N_16448);
nor U18962 (N_18962,N_16695,N_16160);
or U18963 (N_18963,N_16850,N_16481);
and U18964 (N_18964,N_16111,N_17598);
or U18965 (N_18965,N_16320,N_17164);
xor U18966 (N_18966,N_17377,N_17171);
nor U18967 (N_18967,N_17697,N_15808);
nor U18968 (N_18968,N_16217,N_15264);
and U18969 (N_18969,N_15221,N_16982);
or U18970 (N_18970,N_15283,N_16887);
or U18971 (N_18971,N_15731,N_15758);
or U18972 (N_18972,N_16311,N_17299);
and U18973 (N_18973,N_16472,N_15342);
nand U18974 (N_18974,N_17202,N_16752);
nand U18975 (N_18975,N_17881,N_17110);
xor U18976 (N_18976,N_16350,N_17215);
nor U18977 (N_18977,N_15745,N_15801);
or U18978 (N_18978,N_15165,N_17807);
or U18979 (N_18979,N_17129,N_15123);
nor U18980 (N_18980,N_16126,N_16760);
nand U18981 (N_18981,N_17991,N_17130);
and U18982 (N_18982,N_16911,N_15350);
nor U18983 (N_18983,N_16687,N_16345);
nor U18984 (N_18984,N_15715,N_15297);
and U18985 (N_18985,N_15428,N_15122);
and U18986 (N_18986,N_17216,N_17965);
nand U18987 (N_18987,N_17389,N_15019);
nor U18988 (N_18988,N_15594,N_16498);
or U18989 (N_18989,N_17551,N_15830);
nand U18990 (N_18990,N_15099,N_15415);
nor U18991 (N_18991,N_15422,N_16970);
nor U18992 (N_18992,N_15210,N_16117);
nand U18993 (N_18993,N_17447,N_15748);
nand U18994 (N_18994,N_15463,N_17526);
and U18995 (N_18995,N_16742,N_17331);
xor U18996 (N_18996,N_17849,N_17544);
or U18997 (N_18997,N_16420,N_15499);
nor U18998 (N_18998,N_15773,N_15681);
or U18999 (N_18999,N_16555,N_16891);
or U19000 (N_19000,N_16620,N_17462);
or U19001 (N_19001,N_17104,N_16942);
xor U19002 (N_19002,N_17239,N_17040);
xor U19003 (N_19003,N_15560,N_16659);
xnor U19004 (N_19004,N_17730,N_17772);
nor U19005 (N_19005,N_15588,N_16400);
xnor U19006 (N_19006,N_17354,N_15781);
nor U19007 (N_19007,N_17835,N_16768);
nor U19008 (N_19008,N_16051,N_16506);
nand U19009 (N_19009,N_16761,N_16829);
nor U19010 (N_19010,N_16002,N_15534);
xnor U19011 (N_19011,N_17030,N_15299);
nand U19012 (N_19012,N_15782,N_17900);
nand U19013 (N_19013,N_16431,N_16790);
or U19014 (N_19014,N_17904,N_15031);
or U19015 (N_19015,N_17693,N_17141);
nand U19016 (N_19016,N_17348,N_15645);
or U19017 (N_19017,N_16934,N_16140);
and U19018 (N_19018,N_16148,N_17573);
nor U19019 (N_19019,N_15638,N_16702);
and U19020 (N_19020,N_17323,N_17297);
nand U19021 (N_19021,N_17804,N_17720);
xor U19022 (N_19022,N_16871,N_17168);
nor U19023 (N_19023,N_16849,N_17015);
xnor U19024 (N_19024,N_17865,N_16379);
or U19025 (N_19025,N_16483,N_16533);
nor U19026 (N_19026,N_16408,N_15932);
or U19027 (N_19027,N_16494,N_17711);
and U19028 (N_19028,N_17968,N_17642);
or U19029 (N_19029,N_15053,N_17575);
and U19030 (N_19030,N_16247,N_15766);
or U19031 (N_19031,N_16257,N_16146);
or U19032 (N_19032,N_17126,N_16459);
or U19033 (N_19033,N_15317,N_17563);
nand U19034 (N_19034,N_17670,N_15807);
nand U19035 (N_19035,N_15938,N_15631);
or U19036 (N_19036,N_17765,N_15079);
nand U19037 (N_19037,N_15726,N_16199);
nor U19038 (N_19038,N_16132,N_17234);
xor U19039 (N_19039,N_17538,N_15717);
xnor U19040 (N_19040,N_15343,N_16194);
nand U19041 (N_19041,N_16364,N_16339);
nor U19042 (N_19042,N_16048,N_17903);
xnor U19043 (N_19043,N_16076,N_17989);
nand U19044 (N_19044,N_16912,N_15733);
nor U19045 (N_19045,N_15275,N_17635);
nand U19046 (N_19046,N_17497,N_15268);
xnor U19047 (N_19047,N_15183,N_16954);
nor U19048 (N_19048,N_15613,N_17091);
nand U19049 (N_19049,N_17576,N_16898);
nor U19050 (N_19050,N_17767,N_16801);
nor U19051 (N_19051,N_17886,N_17606);
nand U19052 (N_19052,N_16300,N_16187);
and U19053 (N_19053,N_17248,N_16432);
or U19054 (N_19054,N_17506,N_15721);
or U19055 (N_19055,N_17432,N_15710);
or U19056 (N_19056,N_16991,N_15444);
or U19057 (N_19057,N_17513,N_16001);
or U19058 (N_19058,N_15959,N_17775);
nand U19059 (N_19059,N_15651,N_17953);
nor U19060 (N_19060,N_17467,N_16227);
nor U19061 (N_19061,N_15788,N_17883);
nand U19062 (N_19062,N_16343,N_16588);
or U19063 (N_19063,N_17622,N_17120);
nand U19064 (N_19064,N_16928,N_16500);
and U19065 (N_19065,N_15003,N_15947);
xor U19066 (N_19066,N_15067,N_15333);
and U19067 (N_19067,N_15182,N_17152);
xor U19068 (N_19068,N_15603,N_17098);
nor U19069 (N_19069,N_16279,N_15586);
or U19070 (N_19070,N_15814,N_17509);
nor U19071 (N_19071,N_15237,N_17071);
and U19072 (N_19072,N_15640,N_15931);
and U19073 (N_19073,N_16529,N_16058);
or U19074 (N_19074,N_17150,N_17151);
nor U19075 (N_19075,N_15867,N_15532);
and U19076 (N_19076,N_16739,N_15511);
nand U19077 (N_19077,N_15020,N_16878);
and U19078 (N_19078,N_17725,N_16787);
and U19079 (N_19079,N_16092,N_15829);
xnor U19080 (N_19080,N_15916,N_17193);
or U19081 (N_19081,N_17987,N_15842);
nor U19082 (N_19082,N_16584,N_17821);
or U19083 (N_19083,N_17929,N_16643);
nor U19084 (N_19084,N_16105,N_16636);
nand U19085 (N_19085,N_15690,N_16333);
and U19086 (N_19086,N_17634,N_15702);
xor U19087 (N_19087,N_15308,N_15300);
nor U19088 (N_19088,N_16192,N_16756);
nor U19089 (N_19089,N_15155,N_15595);
and U19090 (N_19090,N_16791,N_17049);
nor U19091 (N_19091,N_15881,N_15937);
nor U19092 (N_19092,N_17546,N_15384);
or U19093 (N_19093,N_17525,N_17510);
xor U19094 (N_19094,N_15367,N_17112);
or U19095 (N_19095,N_15999,N_16700);
xnor U19096 (N_19096,N_15366,N_17647);
nand U19097 (N_19097,N_16927,N_16362);
or U19098 (N_19098,N_15504,N_16783);
and U19099 (N_19099,N_17727,N_15764);
nor U19100 (N_19100,N_16471,N_17188);
nand U19101 (N_19101,N_17502,N_15593);
nand U19102 (N_19102,N_16861,N_17131);
nor U19103 (N_19103,N_16122,N_16921);
or U19104 (N_19104,N_16391,N_17915);
nor U19105 (N_19105,N_16635,N_16223);
nor U19106 (N_19106,N_16808,N_15907);
nor U19107 (N_19107,N_15882,N_17192);
nor U19108 (N_19108,N_15440,N_16386);
nand U19109 (N_19109,N_15935,N_17340);
and U19110 (N_19110,N_17335,N_17784);
xnor U19111 (N_19111,N_15425,N_17683);
nor U19112 (N_19112,N_16282,N_17637);
nand U19113 (N_19113,N_15915,N_17423);
nand U19114 (N_19114,N_15244,N_15624);
nand U19115 (N_19115,N_16253,N_15224);
nand U19116 (N_19116,N_17993,N_15229);
nor U19117 (N_19117,N_16650,N_17167);
nor U19118 (N_19118,N_15873,N_16966);
or U19119 (N_19119,N_17955,N_17567);
nor U19120 (N_19120,N_16884,N_15060);
nor U19121 (N_19121,N_15251,N_16063);
or U19122 (N_19122,N_16329,N_16125);
nand U19123 (N_19123,N_15104,N_15072);
nand U19124 (N_19124,N_15037,N_15219);
or U19125 (N_19125,N_15528,N_17128);
nand U19126 (N_19126,N_15371,N_16135);
nand U19127 (N_19127,N_16388,N_15466);
nand U19128 (N_19128,N_16694,N_17564);
or U19129 (N_19129,N_17401,N_15744);
nor U19130 (N_19130,N_16721,N_15047);
nand U19131 (N_19131,N_17060,N_16549);
nor U19132 (N_19132,N_15430,N_15116);
nand U19133 (N_19133,N_15336,N_17897);
and U19134 (N_19134,N_16265,N_15289);
xnor U19135 (N_19135,N_17437,N_15805);
or U19136 (N_19136,N_17349,N_16371);
nor U19137 (N_19137,N_16114,N_16149);
and U19138 (N_19138,N_15125,N_15713);
nor U19139 (N_19139,N_16137,N_17420);
and U19140 (N_19140,N_15952,N_17700);
and U19141 (N_19141,N_17181,N_16016);
and U19142 (N_19142,N_16812,N_17957);
and U19143 (N_19143,N_17478,N_16895);
nor U19144 (N_19144,N_17503,N_17324);
and U19145 (N_19145,N_16403,N_15795);
nor U19146 (N_19146,N_16437,N_17042);
nor U19147 (N_19147,N_16270,N_17378);
and U19148 (N_19148,N_15273,N_15793);
nand U19149 (N_19149,N_17417,N_15845);
nand U19150 (N_19150,N_15963,N_15030);
or U19151 (N_19151,N_17350,N_17415);
nor U19152 (N_19152,N_17056,N_16009);
nor U19153 (N_19153,N_16753,N_16274);
nand U19154 (N_19154,N_15399,N_17869);
nor U19155 (N_19155,N_16248,N_15441);
or U19156 (N_19156,N_17479,N_16268);
nor U19157 (N_19157,N_15124,N_17138);
or U19158 (N_19158,N_15437,N_15790);
or U19159 (N_19159,N_17387,N_16512);
xnor U19160 (N_19160,N_17735,N_17100);
and U19161 (N_19161,N_15883,N_16615);
nor U19162 (N_19162,N_15065,N_17284);
xnor U19163 (N_19163,N_16178,N_15688);
or U19164 (N_19164,N_16003,N_17237);
nand U19165 (N_19165,N_16715,N_17578);
nand U19166 (N_19166,N_17468,N_17851);
nor U19167 (N_19167,N_17685,N_16497);
nor U19168 (N_19168,N_15850,N_16780);
nor U19169 (N_19169,N_15402,N_16264);
or U19170 (N_19170,N_15468,N_16593);
and U19171 (N_19171,N_16501,N_15377);
or U19172 (N_19172,N_15307,N_17770);
nor U19173 (N_19173,N_17177,N_17531);
nand U19174 (N_19174,N_17836,N_17763);
or U19175 (N_19175,N_16569,N_17184);
nor U19176 (N_19176,N_17777,N_17208);
and U19177 (N_19177,N_16171,N_16252);
nand U19178 (N_19178,N_16121,N_16487);
nand U19179 (N_19179,N_15234,N_16965);
nor U19180 (N_19180,N_16173,N_17233);
nand U19181 (N_19181,N_17782,N_16062);
or U19182 (N_19182,N_15119,N_16159);
or U19183 (N_19183,N_15994,N_17482);
nor U19184 (N_19184,N_16249,N_15351);
or U19185 (N_19185,N_17666,N_15319);
xor U19186 (N_19186,N_17140,N_16093);
nor U19187 (N_19187,N_17516,N_15478);
nand U19188 (N_19188,N_16969,N_16856);
and U19189 (N_19189,N_17428,N_17885);
and U19190 (N_19190,N_15103,N_15167);
nand U19191 (N_19191,N_16496,N_16984);
or U19192 (N_19192,N_16749,N_16899);
nor U19193 (N_19193,N_17114,N_15243);
nor U19194 (N_19194,N_17995,N_16479);
and U19195 (N_19195,N_17359,N_16397);
nand U19196 (N_19196,N_15579,N_17643);
nor U19197 (N_19197,N_17165,N_16998);
nand U19198 (N_19198,N_17599,N_15357);
nor U19199 (N_19199,N_15519,N_17074);
and U19200 (N_19200,N_17047,N_15291);
nand U19201 (N_19201,N_16305,N_17132);
nand U19202 (N_19202,N_17654,N_17712);
nor U19203 (N_19203,N_15228,N_16218);
nor U19204 (N_19204,N_15379,N_16558);
xnor U19205 (N_19205,N_15085,N_15997);
or U19206 (N_19206,N_16677,N_17003);
xor U19207 (N_19207,N_17124,N_17052);
nor U19208 (N_19208,N_17289,N_16730);
or U19209 (N_19209,N_17882,N_15846);
xor U19210 (N_19210,N_15824,N_15327);
or U19211 (N_19211,N_16827,N_16704);
nand U19212 (N_19212,N_17473,N_15426);
and U19213 (N_19213,N_15447,N_16073);
nand U19214 (N_19214,N_15677,N_15988);
nor U19215 (N_19215,N_17738,N_16606);
or U19216 (N_19216,N_16681,N_17969);
and U19217 (N_19217,N_15811,N_17716);
nand U19218 (N_19218,N_17958,N_17230);
xor U19219 (N_19219,N_15797,N_17761);
or U19220 (N_19220,N_17493,N_16072);
and U19221 (N_19221,N_17660,N_15542);
nor U19222 (N_19222,N_16709,N_17277);
or U19223 (N_19223,N_17924,N_15349);
nor U19224 (N_19224,N_15708,N_15153);
or U19225 (N_19225,N_15023,N_16118);
or U19226 (N_19226,N_17064,N_16925);
or U19227 (N_19227,N_15368,N_17680);
and U19228 (N_19228,N_15614,N_15818);
or U19229 (N_19229,N_16535,N_16470);
or U19230 (N_19230,N_15803,N_15512);
and U19231 (N_19231,N_15516,N_16995);
and U19232 (N_19232,N_15831,N_16574);
and U19233 (N_19233,N_17603,N_15281);
and U19234 (N_19234,N_15438,N_15716);
or U19235 (N_19235,N_15321,N_17231);
nand U19236 (N_19236,N_17824,N_17016);
nor U19237 (N_19237,N_17006,N_16297);
nor U19238 (N_19238,N_15792,N_16733);
and U19239 (N_19239,N_17369,N_16577);
or U19240 (N_19240,N_17604,N_16104);
and U19241 (N_19241,N_17536,N_15903);
xor U19242 (N_19242,N_16179,N_15641);
or U19243 (N_19243,N_17834,N_15639);
nand U19244 (N_19244,N_17596,N_15895);
or U19245 (N_19245,N_15419,N_16505);
xnor U19246 (N_19246,N_16238,N_16324);
nand U19247 (N_19247,N_15553,N_17391);
or U19248 (N_19248,N_16805,N_16214);
nor U19249 (N_19249,N_16770,N_16673);
nand U19250 (N_19250,N_16316,N_15853);
nand U19251 (N_19251,N_17611,N_15664);
and U19252 (N_19252,N_15703,N_15756);
and U19253 (N_19253,N_16691,N_17699);
nor U19254 (N_19254,N_16875,N_17691);
or U19255 (N_19255,N_15798,N_15078);
xor U19256 (N_19256,N_17206,N_17586);
nand U19257 (N_19257,N_16688,N_16344);
or U19258 (N_19258,N_17706,N_17861);
or U19259 (N_19259,N_17436,N_15087);
or U19260 (N_19260,N_15458,N_16806);
nand U19261 (N_19261,N_15147,N_15252);
nor U19262 (N_19262,N_17393,N_15998);
or U19263 (N_19263,N_15253,N_16398);
or U19264 (N_19264,N_17170,N_15960);
and U19265 (N_19265,N_15207,N_15035);
and U19266 (N_19266,N_17232,N_16692);
nand U19267 (N_19267,N_17801,N_16839);
nor U19268 (N_19268,N_15902,N_15396);
nor U19269 (N_19269,N_17708,N_17527);
or U19270 (N_19270,N_17223,N_16637);
nand U19271 (N_19271,N_16356,N_15114);
nor U19272 (N_19272,N_15335,N_15054);
or U19273 (N_19273,N_15101,N_15546);
nand U19274 (N_19274,N_17187,N_15572);
nor U19275 (N_19275,N_15433,N_16804);
nor U19276 (N_19276,N_16088,N_15208);
or U19277 (N_19277,N_15868,N_16979);
xnor U19278 (N_19278,N_15779,N_17698);
nor U19279 (N_19279,N_17522,N_15982);
nor U19280 (N_19280,N_17774,N_17311);
or U19281 (N_19281,N_16725,N_16640);
or U19282 (N_19282,N_16186,N_16286);
xor U19283 (N_19283,N_15871,N_17102);
or U19284 (N_19284,N_17518,N_17658);
nor U19285 (N_19285,N_15887,N_15945);
xnor U19286 (N_19286,N_15863,N_17715);
or U19287 (N_19287,N_15587,N_15967);
or U19288 (N_19288,N_17477,N_15704);
nand U19289 (N_19289,N_17410,N_15168);
and U19290 (N_19290,N_15761,N_17657);
nand U19291 (N_19291,N_15129,N_15772);
and U19292 (N_19292,N_15763,N_17895);
and U19293 (N_19293,N_15557,N_15212);
or U19294 (N_19294,N_15112,N_15514);
or U19295 (N_19295,N_17830,N_16782);
xor U19296 (N_19296,N_16614,N_16592);
nand U19297 (N_19297,N_17818,N_16307);
nor U19298 (N_19298,N_17225,N_17762);
nor U19299 (N_19299,N_17403,N_17075);
nor U19300 (N_19300,N_15836,N_17023);
nand U19301 (N_19301,N_16439,N_17317);
or U19302 (N_19302,N_17203,N_17200);
nor U19303 (N_19303,N_17201,N_17089);
xnor U19304 (N_19304,N_16622,N_15661);
nor U19305 (N_19305,N_15646,N_17831);
nand U19306 (N_19306,N_16828,N_17455);
or U19307 (N_19307,N_16689,N_16395);
nand U19308 (N_19308,N_16429,N_16764);
and U19309 (N_19309,N_16837,N_15984);
or U19310 (N_19310,N_17318,N_15397);
or U19311 (N_19311,N_16830,N_17682);
nor U19312 (N_19312,N_15926,N_15089);
and U19313 (N_19313,N_16038,N_15198);
nand U19314 (N_19314,N_16418,N_16617);
or U19315 (N_19315,N_16508,N_17285);
and U19316 (N_19316,N_17748,N_15564);
or U19317 (N_19317,N_17539,N_16240);
nand U19318 (N_19318,N_17902,N_17979);
and U19319 (N_19319,N_17592,N_15872);
or U19320 (N_19320,N_15310,N_17386);
or U19321 (N_19321,N_17338,N_16390);
or U19322 (N_19322,N_16462,N_17749);
nor U19323 (N_19323,N_16050,N_16576);
or U19324 (N_19324,N_17872,N_17709);
nor U19325 (N_19325,N_17922,N_17561);
xor U19326 (N_19326,N_15358,N_15213);
and U19327 (N_19327,N_15177,N_16442);
or U19328 (N_19328,N_17179,N_16579);
and U19329 (N_19329,N_17607,N_17589);
and U19330 (N_19330,N_16095,N_15270);
and U19331 (N_19331,N_15986,N_16043);
or U19332 (N_19332,N_15964,N_16394);
and U19333 (N_19333,N_16886,N_16134);
nand U19334 (N_19334,N_16813,N_15580);
and U19335 (N_19335,N_17440,N_16164);
or U19336 (N_19336,N_16999,N_17375);
xor U19337 (N_19337,N_17050,N_17282);
and U19338 (N_19338,N_15487,N_17268);
or U19339 (N_19339,N_16655,N_17007);
nand U19340 (N_19340,N_15429,N_17982);
or U19341 (N_19341,N_16245,N_17439);
xor U19342 (N_19342,N_17811,N_17051);
and U19343 (N_19343,N_15992,N_17940);
nor U19344 (N_19344,N_16820,N_17627);
or U19345 (N_19345,N_15826,N_15577);
or U19346 (N_19346,N_17079,N_16176);
nor U19347 (N_19347,N_15050,N_15765);
nor U19348 (N_19348,N_16231,N_16776);
or U19349 (N_19349,N_15923,N_16308);
and U19350 (N_19350,N_15630,N_16440);
nand U19351 (N_19351,N_17602,N_15280);
xor U19352 (N_19352,N_16723,N_17291);
nand U19353 (N_19353,N_17571,N_17072);
and U19354 (N_19354,N_17964,N_17864);
nand U19355 (N_19355,N_15236,N_16944);
xnor U19356 (N_19356,N_17093,N_15239);
and U19357 (N_19357,N_17262,N_15260);
nand U19358 (N_19358,N_16441,N_15469);
and U19359 (N_19359,N_17945,N_15355);
nand U19360 (N_19360,N_17630,N_16239);
or U19361 (N_19361,N_16285,N_17747);
nand U19362 (N_19362,N_17843,N_17718);
or U19363 (N_19363,N_15919,N_15459);
and U19364 (N_19364,N_17211,N_16507);
and U19365 (N_19365,N_16918,N_17286);
or U19366 (N_19366,N_16523,N_16701);
or U19367 (N_19367,N_15022,N_17315);
or U19368 (N_19368,N_16510,N_16863);
and U19369 (N_19369,N_17568,N_16716);
and U19370 (N_19370,N_15993,N_17329);
xor U19371 (N_19371,N_17951,N_16893);
nor U19372 (N_19372,N_16980,N_17858);
nor U19373 (N_19373,N_16990,N_15900);
nand U19374 (N_19374,N_16722,N_16955);
nand U19375 (N_19375,N_16926,N_17815);
or U19376 (N_19376,N_15518,N_16818);
or U19377 (N_19377,N_15636,N_16807);
or U19378 (N_19378,N_17659,N_15348);
nand U19379 (N_19379,N_16241,N_15410);
or U19380 (N_19380,N_15174,N_15653);
or U19381 (N_19381,N_15187,N_15612);
nand U19382 (N_19382,N_16843,N_15897);
nand U19383 (N_19383,N_15288,N_16641);
nor U19384 (N_19384,N_15632,N_17281);
or U19385 (N_19385,N_17779,N_17274);
nor U19386 (N_19386,N_16499,N_16402);
and U19387 (N_19387,N_15172,N_17143);
and U19388 (N_19388,N_16901,N_15255);
and U19389 (N_19389,N_16597,N_16815);
and U19390 (N_19390,N_16530,N_15944);
nor U19391 (N_19391,N_17916,N_17854);
and U19392 (N_19392,N_16144,N_16611);
and U19393 (N_19393,N_17360,N_15408);
nand U19394 (N_19394,N_15911,N_15701);
or U19395 (N_19395,N_16123,N_15282);
nor U19396 (N_19396,N_17844,N_15946);
and U19397 (N_19397,N_15226,N_16738);
and U19398 (N_19398,N_17878,N_15526);
or U19399 (N_19399,N_15039,N_16774);
or U19400 (N_19400,N_16361,N_17025);
nand U19401 (N_19401,N_17703,N_17476);
xnor U19402 (N_19402,N_17966,N_16319);
nand U19403 (N_19403,N_15768,N_16633);
or U19404 (N_19404,N_15025,N_15864);
nand U19405 (N_19405,N_15202,N_15449);
or U19406 (N_19406,N_17453,N_15956);
nor U19407 (N_19407,N_15345,N_17207);
and U19408 (N_19408,N_15633,N_17721);
or U19409 (N_19409,N_16162,N_17554);
and U19410 (N_19410,N_16778,N_17309);
or U19411 (N_19411,N_16047,N_17474);
xnor U19412 (N_19412,N_16793,N_15732);
and U19413 (N_19413,N_16560,N_17162);
or U19414 (N_19414,N_17070,N_15046);
and U19415 (N_19415,N_16594,N_17585);
nand U19416 (N_19416,N_16013,N_15423);
xnor U19417 (N_19417,N_15223,N_17472);
and U19418 (N_19418,N_16277,N_17196);
xor U19419 (N_19419,N_16120,N_17096);
or U19420 (N_19420,N_15339,N_16272);
or U19421 (N_19421,N_16314,N_16208);
xnor U19422 (N_19422,N_15462,N_16762);
nor U19423 (N_19423,N_15835,N_15533);
xnor U19424 (N_19424,N_15691,N_16547);
or U19425 (N_19425,N_15205,N_16623);
nor U19426 (N_19426,N_16433,N_16421);
and U19427 (N_19427,N_17726,N_17419);
nand U19428 (N_19428,N_15215,N_15448);
nor U19429 (N_19429,N_16256,N_16751);
nand U19430 (N_19430,N_17791,N_15394);
or U19431 (N_19431,N_16184,N_15581);
and U19432 (N_19432,N_16490,N_16425);
nor U19433 (N_19433,N_15649,N_15896);
xor U19434 (N_19434,N_16968,N_16554);
nand U19435 (N_19435,N_15660,N_17809);
nand U19436 (N_19436,N_15621,N_16422);
or U19437 (N_19437,N_17961,N_16515);
nor U19438 (N_19438,N_15083,N_17494);
nand U19439 (N_19439,N_15742,N_16033);
or U19440 (N_19440,N_16416,N_17689);
nand U19441 (N_19441,N_16833,N_15162);
and U19442 (N_19442,N_16883,N_17308);
or U19443 (N_19443,N_15502,N_15446);
nand U19444 (N_19444,N_15439,N_17998);
nor U19445 (N_19445,N_17163,N_16590);
or U19446 (N_19446,N_17545,N_16392);
nand U19447 (N_19447,N_16066,N_17442);
or U19448 (N_19448,N_16699,N_17798);
nor U19449 (N_19449,N_17293,N_17990);
and U19450 (N_19450,N_16133,N_15055);
and U19451 (N_19451,N_16516,N_17960);
nor U19452 (N_19452,N_16750,N_15298);
or U19453 (N_19453,N_15320,N_17868);
xor U19454 (N_19454,N_17508,N_17892);
nand U19455 (N_19455,N_15889,N_16502);
or U19456 (N_19456,N_16917,N_16172);
or U19457 (N_19457,N_17133,N_16854);
and U19458 (N_19458,N_17134,N_15118);
or U19459 (N_19459,N_17667,N_17988);
or U19460 (N_19460,N_15033,N_15890);
nor U19461 (N_19461,N_16524,N_17431);
nor U19462 (N_19462,N_15263,N_15106);
or U19463 (N_19463,N_15578,N_17690);
xnor U19464 (N_19464,N_16851,N_15510);
xor U19465 (N_19465,N_15248,N_15143);
or U19466 (N_19466,N_17287,N_17860);
nand U19467 (N_19467,N_17272,N_17898);
xnor U19468 (N_19468,N_15117,N_16647);
nor U19469 (N_19469,N_17548,N_15269);
nor U19470 (N_19470,N_15475,N_17570);
and U19471 (N_19471,N_16720,N_15709);
nand U19472 (N_19472,N_15547,N_16654);
nor U19473 (N_19473,N_16310,N_17662);
nor U19474 (N_19474,N_17625,N_16152);
and U19475 (N_19475,N_16823,N_15258);
xor U19476 (N_19476,N_15375,N_16840);
nand U19477 (N_19477,N_15092,N_15529);
and U19478 (N_19478,N_17113,N_17495);
nor U19479 (N_19479,N_16986,N_16719);
nor U19480 (N_19480,N_17745,N_17906);
nor U19481 (N_19481,N_16189,N_16903);
or U19482 (N_19482,N_17136,N_17066);
nand U19483 (N_19483,N_15151,N_15878);
nor U19484 (N_19484,N_15562,N_16587);
nor U19485 (N_19485,N_17605,N_15290);
or U19486 (N_19486,N_15370,N_15045);
nand U19487 (N_19487,N_17313,N_15373);
or U19488 (N_19488,N_17002,N_17692);
and U19489 (N_19489,N_16221,N_17600);
and U19490 (N_19490,N_16276,N_15414);
and U19491 (N_19491,N_17894,N_17820);
and U19492 (N_19492,N_15435,N_15073);
and U19493 (N_19493,N_16302,N_15567);
nand U19494 (N_19494,N_17759,N_17068);
nor U19495 (N_19495,N_16842,N_16656);
nand U19496 (N_19496,N_16097,N_16468);
nor U19497 (N_19497,N_15530,N_15780);
xor U19498 (N_19498,N_17817,N_15608);
xnor U19499 (N_19499,N_15416,N_16797);
xor U19500 (N_19500,N_15455,N_15079);
or U19501 (N_19501,N_16743,N_17350);
and U19502 (N_19502,N_16003,N_16897);
xnor U19503 (N_19503,N_15676,N_15729);
nor U19504 (N_19504,N_15752,N_16485);
nor U19505 (N_19505,N_17665,N_15905);
nand U19506 (N_19506,N_17657,N_15750);
nand U19507 (N_19507,N_16139,N_17928);
nor U19508 (N_19508,N_17335,N_17821);
nand U19509 (N_19509,N_15711,N_15138);
nand U19510 (N_19510,N_16804,N_15575);
nand U19511 (N_19511,N_15664,N_17936);
nor U19512 (N_19512,N_16007,N_15481);
or U19513 (N_19513,N_17520,N_15661);
nand U19514 (N_19514,N_17864,N_17355);
nor U19515 (N_19515,N_15982,N_16882);
nand U19516 (N_19516,N_17569,N_17458);
and U19517 (N_19517,N_17830,N_16274);
xor U19518 (N_19518,N_16744,N_17448);
or U19519 (N_19519,N_16982,N_17378);
or U19520 (N_19520,N_15652,N_16706);
nand U19521 (N_19521,N_17673,N_16063);
xor U19522 (N_19522,N_15620,N_15317);
or U19523 (N_19523,N_16399,N_16155);
nor U19524 (N_19524,N_17925,N_17483);
nor U19525 (N_19525,N_17350,N_16228);
and U19526 (N_19526,N_17225,N_17280);
and U19527 (N_19527,N_16317,N_17366);
xnor U19528 (N_19528,N_15306,N_15054);
and U19529 (N_19529,N_16572,N_16322);
nand U19530 (N_19530,N_17062,N_17634);
nor U19531 (N_19531,N_17535,N_16494);
xnor U19532 (N_19532,N_17326,N_17617);
nor U19533 (N_19533,N_15198,N_17335);
xnor U19534 (N_19534,N_16494,N_17829);
nor U19535 (N_19535,N_17729,N_15808);
and U19536 (N_19536,N_16436,N_15700);
xnor U19537 (N_19537,N_17412,N_16226);
and U19538 (N_19538,N_17491,N_15864);
or U19539 (N_19539,N_15004,N_17283);
nor U19540 (N_19540,N_16885,N_16089);
or U19541 (N_19541,N_17316,N_17817);
nor U19542 (N_19542,N_16751,N_16521);
nand U19543 (N_19543,N_15569,N_16382);
and U19544 (N_19544,N_16103,N_15595);
and U19545 (N_19545,N_16265,N_17558);
nand U19546 (N_19546,N_17523,N_15886);
or U19547 (N_19547,N_16692,N_15713);
and U19548 (N_19548,N_15119,N_15570);
or U19549 (N_19549,N_15911,N_17050);
and U19550 (N_19550,N_15143,N_16554);
or U19551 (N_19551,N_16320,N_15198);
nor U19552 (N_19552,N_17783,N_17469);
or U19553 (N_19553,N_16610,N_17036);
or U19554 (N_19554,N_16845,N_15851);
and U19555 (N_19555,N_17587,N_17847);
or U19556 (N_19556,N_17627,N_15134);
nor U19557 (N_19557,N_17406,N_16614);
and U19558 (N_19558,N_16256,N_16032);
or U19559 (N_19559,N_15226,N_15178);
and U19560 (N_19560,N_16507,N_15632);
and U19561 (N_19561,N_16059,N_15465);
or U19562 (N_19562,N_15649,N_16217);
nor U19563 (N_19563,N_16849,N_16244);
nor U19564 (N_19564,N_15184,N_17207);
and U19565 (N_19565,N_15494,N_17631);
and U19566 (N_19566,N_15712,N_16084);
or U19567 (N_19567,N_15681,N_16327);
nand U19568 (N_19568,N_16892,N_15990);
xnor U19569 (N_19569,N_16886,N_17481);
and U19570 (N_19570,N_16394,N_15664);
xor U19571 (N_19571,N_16069,N_16730);
nor U19572 (N_19572,N_16535,N_17473);
xnor U19573 (N_19573,N_15651,N_16591);
nand U19574 (N_19574,N_16056,N_15821);
nand U19575 (N_19575,N_17275,N_17819);
and U19576 (N_19576,N_15937,N_17532);
and U19577 (N_19577,N_16516,N_15038);
nand U19578 (N_19578,N_17414,N_17408);
nand U19579 (N_19579,N_16200,N_17693);
or U19580 (N_19580,N_17034,N_17130);
nor U19581 (N_19581,N_15897,N_15687);
nor U19582 (N_19582,N_15071,N_17163);
nand U19583 (N_19583,N_15756,N_15415);
and U19584 (N_19584,N_16708,N_16101);
and U19585 (N_19585,N_17812,N_17054);
nor U19586 (N_19586,N_15758,N_17330);
nor U19587 (N_19587,N_17802,N_15728);
xor U19588 (N_19588,N_17360,N_16625);
and U19589 (N_19589,N_17487,N_16399);
and U19590 (N_19590,N_15339,N_17380);
nand U19591 (N_19591,N_17425,N_17998);
nor U19592 (N_19592,N_17069,N_17400);
and U19593 (N_19593,N_16538,N_15365);
nand U19594 (N_19594,N_15537,N_17637);
xnor U19595 (N_19595,N_17420,N_16066);
or U19596 (N_19596,N_15719,N_17536);
and U19597 (N_19597,N_17805,N_17833);
or U19598 (N_19598,N_16325,N_17199);
nand U19599 (N_19599,N_17938,N_16143);
xnor U19600 (N_19600,N_17119,N_15933);
nor U19601 (N_19601,N_16723,N_17537);
xor U19602 (N_19602,N_16200,N_17510);
or U19603 (N_19603,N_15729,N_16953);
or U19604 (N_19604,N_17047,N_15412);
nand U19605 (N_19605,N_17561,N_16024);
or U19606 (N_19606,N_15608,N_15726);
xnor U19607 (N_19607,N_15036,N_16107);
nor U19608 (N_19608,N_15741,N_15947);
xnor U19609 (N_19609,N_15575,N_15412);
and U19610 (N_19610,N_16011,N_15587);
nand U19611 (N_19611,N_16870,N_17554);
nor U19612 (N_19612,N_16319,N_17895);
nand U19613 (N_19613,N_15451,N_17386);
xor U19614 (N_19614,N_16255,N_17431);
nor U19615 (N_19615,N_15549,N_17257);
and U19616 (N_19616,N_15031,N_17339);
and U19617 (N_19617,N_17552,N_17894);
and U19618 (N_19618,N_17236,N_17528);
and U19619 (N_19619,N_15097,N_17692);
nand U19620 (N_19620,N_17043,N_15898);
nand U19621 (N_19621,N_16708,N_17406);
nor U19622 (N_19622,N_16340,N_17397);
or U19623 (N_19623,N_15831,N_16495);
nor U19624 (N_19624,N_15077,N_16105);
nor U19625 (N_19625,N_15589,N_16820);
nor U19626 (N_19626,N_15476,N_15358);
nor U19627 (N_19627,N_17540,N_16887);
or U19628 (N_19628,N_16985,N_15118);
or U19629 (N_19629,N_16503,N_15146);
and U19630 (N_19630,N_15591,N_17389);
xnor U19631 (N_19631,N_16394,N_17796);
nor U19632 (N_19632,N_15195,N_15052);
or U19633 (N_19633,N_17249,N_15997);
or U19634 (N_19634,N_16449,N_16859);
nand U19635 (N_19635,N_17525,N_17898);
nand U19636 (N_19636,N_17546,N_16901);
and U19637 (N_19637,N_15648,N_15644);
nor U19638 (N_19638,N_17400,N_15935);
or U19639 (N_19639,N_15390,N_17222);
nand U19640 (N_19640,N_17723,N_17845);
nand U19641 (N_19641,N_15283,N_17623);
xor U19642 (N_19642,N_17447,N_16341);
nand U19643 (N_19643,N_16146,N_15994);
and U19644 (N_19644,N_15770,N_15913);
nor U19645 (N_19645,N_17044,N_16162);
or U19646 (N_19646,N_17301,N_16261);
and U19647 (N_19647,N_15728,N_15083);
and U19648 (N_19648,N_16142,N_15700);
and U19649 (N_19649,N_15955,N_17144);
nand U19650 (N_19650,N_17007,N_17728);
nor U19651 (N_19651,N_16886,N_17588);
nand U19652 (N_19652,N_17552,N_15733);
nor U19653 (N_19653,N_16055,N_15397);
nor U19654 (N_19654,N_16855,N_17632);
nand U19655 (N_19655,N_15968,N_17504);
and U19656 (N_19656,N_15547,N_15280);
and U19657 (N_19657,N_16573,N_15516);
nand U19658 (N_19658,N_17837,N_15900);
or U19659 (N_19659,N_15364,N_15957);
nor U19660 (N_19660,N_17491,N_17153);
nand U19661 (N_19661,N_16181,N_17822);
or U19662 (N_19662,N_16682,N_17509);
and U19663 (N_19663,N_15137,N_15278);
nand U19664 (N_19664,N_16456,N_17278);
nand U19665 (N_19665,N_15680,N_17167);
or U19666 (N_19666,N_16147,N_15958);
xor U19667 (N_19667,N_16545,N_15110);
xnor U19668 (N_19668,N_17708,N_15858);
nor U19669 (N_19669,N_16044,N_17969);
and U19670 (N_19670,N_16358,N_16381);
nand U19671 (N_19671,N_15634,N_17825);
and U19672 (N_19672,N_16198,N_16310);
nor U19673 (N_19673,N_16241,N_15613);
nor U19674 (N_19674,N_15341,N_17123);
and U19675 (N_19675,N_17894,N_16911);
and U19676 (N_19676,N_16873,N_15707);
or U19677 (N_19677,N_17506,N_17580);
nand U19678 (N_19678,N_16421,N_15485);
and U19679 (N_19679,N_16502,N_16670);
nand U19680 (N_19680,N_17113,N_16192);
xor U19681 (N_19681,N_16211,N_16127);
nand U19682 (N_19682,N_16345,N_16654);
nand U19683 (N_19683,N_17566,N_16411);
or U19684 (N_19684,N_17580,N_15942);
and U19685 (N_19685,N_16882,N_16439);
nand U19686 (N_19686,N_17115,N_16258);
nor U19687 (N_19687,N_17287,N_17696);
and U19688 (N_19688,N_15818,N_16700);
nor U19689 (N_19689,N_17192,N_16387);
nand U19690 (N_19690,N_16107,N_15911);
nand U19691 (N_19691,N_15482,N_16692);
nor U19692 (N_19692,N_17994,N_16829);
xnor U19693 (N_19693,N_17286,N_16669);
and U19694 (N_19694,N_17604,N_17859);
nand U19695 (N_19695,N_16167,N_16523);
and U19696 (N_19696,N_16445,N_15000);
nand U19697 (N_19697,N_16630,N_16867);
and U19698 (N_19698,N_17424,N_16114);
and U19699 (N_19699,N_16226,N_17627);
or U19700 (N_19700,N_17628,N_15933);
nand U19701 (N_19701,N_15426,N_17810);
and U19702 (N_19702,N_16241,N_16908);
nor U19703 (N_19703,N_17600,N_16234);
nand U19704 (N_19704,N_17732,N_16796);
nand U19705 (N_19705,N_16155,N_16094);
nor U19706 (N_19706,N_17515,N_15168);
xnor U19707 (N_19707,N_15128,N_16031);
nor U19708 (N_19708,N_16411,N_16408);
or U19709 (N_19709,N_17228,N_15076);
and U19710 (N_19710,N_16772,N_16528);
nor U19711 (N_19711,N_15613,N_17760);
nand U19712 (N_19712,N_16795,N_16912);
or U19713 (N_19713,N_17496,N_15077);
nand U19714 (N_19714,N_15236,N_17714);
xor U19715 (N_19715,N_15987,N_15711);
nand U19716 (N_19716,N_17978,N_15120);
nor U19717 (N_19717,N_15969,N_17135);
or U19718 (N_19718,N_15246,N_17763);
nor U19719 (N_19719,N_15430,N_15478);
or U19720 (N_19720,N_16735,N_17542);
nor U19721 (N_19721,N_16395,N_15047);
xnor U19722 (N_19722,N_15589,N_16967);
or U19723 (N_19723,N_16577,N_15368);
and U19724 (N_19724,N_16020,N_17332);
and U19725 (N_19725,N_15821,N_16524);
and U19726 (N_19726,N_15974,N_15739);
nand U19727 (N_19727,N_16741,N_15165);
and U19728 (N_19728,N_15596,N_17549);
nand U19729 (N_19729,N_17466,N_16137);
and U19730 (N_19730,N_17206,N_15083);
xnor U19731 (N_19731,N_17463,N_15875);
and U19732 (N_19732,N_17554,N_17707);
and U19733 (N_19733,N_15593,N_17201);
nor U19734 (N_19734,N_15438,N_17137);
and U19735 (N_19735,N_17886,N_17913);
and U19736 (N_19736,N_15511,N_17141);
or U19737 (N_19737,N_16214,N_15839);
nand U19738 (N_19738,N_17654,N_17316);
or U19739 (N_19739,N_17511,N_15116);
xnor U19740 (N_19740,N_16440,N_15138);
nand U19741 (N_19741,N_15026,N_15641);
nor U19742 (N_19742,N_16969,N_17912);
and U19743 (N_19743,N_16786,N_17868);
nor U19744 (N_19744,N_16826,N_15445);
nand U19745 (N_19745,N_17357,N_15801);
or U19746 (N_19746,N_17266,N_16825);
nor U19747 (N_19747,N_17754,N_17490);
and U19748 (N_19748,N_17688,N_16368);
or U19749 (N_19749,N_17979,N_15155);
nand U19750 (N_19750,N_15642,N_15314);
and U19751 (N_19751,N_15905,N_15664);
or U19752 (N_19752,N_17880,N_15950);
and U19753 (N_19753,N_15022,N_16120);
or U19754 (N_19754,N_15624,N_16316);
xnor U19755 (N_19755,N_15253,N_16149);
nand U19756 (N_19756,N_16915,N_15978);
or U19757 (N_19757,N_15787,N_17229);
nor U19758 (N_19758,N_16692,N_16435);
nand U19759 (N_19759,N_15627,N_17521);
nand U19760 (N_19760,N_15861,N_16305);
or U19761 (N_19761,N_16476,N_16369);
nor U19762 (N_19762,N_17656,N_16740);
and U19763 (N_19763,N_15930,N_16512);
and U19764 (N_19764,N_16546,N_16668);
and U19765 (N_19765,N_16919,N_15620);
and U19766 (N_19766,N_15726,N_15634);
nand U19767 (N_19767,N_17888,N_15969);
nand U19768 (N_19768,N_15406,N_15208);
and U19769 (N_19769,N_16125,N_17920);
and U19770 (N_19770,N_17018,N_17313);
and U19771 (N_19771,N_17424,N_16141);
nand U19772 (N_19772,N_15413,N_17383);
nand U19773 (N_19773,N_17310,N_15675);
nor U19774 (N_19774,N_15820,N_15346);
nand U19775 (N_19775,N_15452,N_17549);
nor U19776 (N_19776,N_17342,N_17455);
nor U19777 (N_19777,N_16285,N_16435);
nand U19778 (N_19778,N_15991,N_17374);
or U19779 (N_19779,N_15115,N_16017);
nand U19780 (N_19780,N_15056,N_17853);
nor U19781 (N_19781,N_15196,N_16989);
and U19782 (N_19782,N_16161,N_17435);
and U19783 (N_19783,N_15677,N_17697);
and U19784 (N_19784,N_17008,N_16994);
xnor U19785 (N_19785,N_15583,N_15617);
nor U19786 (N_19786,N_16318,N_16243);
nand U19787 (N_19787,N_15831,N_15555);
nand U19788 (N_19788,N_17040,N_16363);
or U19789 (N_19789,N_15752,N_16773);
nor U19790 (N_19790,N_17671,N_16416);
and U19791 (N_19791,N_15825,N_17818);
nand U19792 (N_19792,N_16435,N_16371);
nor U19793 (N_19793,N_16960,N_15420);
nor U19794 (N_19794,N_16187,N_16646);
nor U19795 (N_19795,N_15207,N_15467);
or U19796 (N_19796,N_16792,N_17597);
nand U19797 (N_19797,N_17945,N_17814);
and U19798 (N_19798,N_15005,N_16531);
nor U19799 (N_19799,N_16353,N_15944);
and U19800 (N_19800,N_16679,N_16251);
nor U19801 (N_19801,N_15809,N_15521);
xnor U19802 (N_19802,N_16227,N_15393);
nand U19803 (N_19803,N_17084,N_17902);
or U19804 (N_19804,N_17317,N_16919);
nor U19805 (N_19805,N_17885,N_17486);
or U19806 (N_19806,N_15653,N_15207);
nand U19807 (N_19807,N_15891,N_15900);
and U19808 (N_19808,N_15257,N_16252);
and U19809 (N_19809,N_17492,N_16850);
or U19810 (N_19810,N_16041,N_17838);
nor U19811 (N_19811,N_17752,N_16743);
and U19812 (N_19812,N_15586,N_17421);
xor U19813 (N_19813,N_15781,N_15969);
or U19814 (N_19814,N_16060,N_15806);
and U19815 (N_19815,N_16354,N_16987);
xnor U19816 (N_19816,N_16382,N_17019);
nor U19817 (N_19817,N_17928,N_15644);
xnor U19818 (N_19818,N_15006,N_16446);
nor U19819 (N_19819,N_15300,N_17270);
or U19820 (N_19820,N_15450,N_15444);
or U19821 (N_19821,N_17660,N_15881);
nand U19822 (N_19822,N_17542,N_17933);
nand U19823 (N_19823,N_17657,N_16089);
nor U19824 (N_19824,N_17381,N_16691);
xnor U19825 (N_19825,N_17839,N_15609);
and U19826 (N_19826,N_16208,N_17629);
nand U19827 (N_19827,N_15505,N_16038);
and U19828 (N_19828,N_17826,N_17161);
nor U19829 (N_19829,N_15960,N_17477);
xor U19830 (N_19830,N_15874,N_17190);
nor U19831 (N_19831,N_16049,N_16057);
nor U19832 (N_19832,N_17258,N_15702);
and U19833 (N_19833,N_17818,N_16413);
or U19834 (N_19834,N_15960,N_17200);
nand U19835 (N_19835,N_15840,N_15661);
nor U19836 (N_19836,N_16438,N_17549);
or U19837 (N_19837,N_15673,N_15278);
nor U19838 (N_19838,N_15052,N_17426);
and U19839 (N_19839,N_16150,N_16034);
nor U19840 (N_19840,N_16974,N_16099);
and U19841 (N_19841,N_16856,N_17484);
or U19842 (N_19842,N_17818,N_16170);
and U19843 (N_19843,N_16422,N_16244);
xnor U19844 (N_19844,N_17333,N_16000);
and U19845 (N_19845,N_16759,N_16884);
or U19846 (N_19846,N_16063,N_17089);
nor U19847 (N_19847,N_15103,N_17147);
nor U19848 (N_19848,N_15450,N_16002);
or U19849 (N_19849,N_15344,N_15252);
nor U19850 (N_19850,N_16032,N_17700);
nor U19851 (N_19851,N_15400,N_15314);
nor U19852 (N_19852,N_15742,N_15641);
or U19853 (N_19853,N_17882,N_16078);
or U19854 (N_19854,N_15641,N_15539);
xnor U19855 (N_19855,N_17093,N_15088);
and U19856 (N_19856,N_17309,N_15615);
or U19857 (N_19857,N_15584,N_17494);
nor U19858 (N_19858,N_17224,N_16602);
xor U19859 (N_19859,N_15365,N_16588);
nor U19860 (N_19860,N_15565,N_16029);
nand U19861 (N_19861,N_17771,N_17073);
nor U19862 (N_19862,N_15553,N_16762);
or U19863 (N_19863,N_17919,N_15567);
nand U19864 (N_19864,N_16741,N_15111);
nor U19865 (N_19865,N_17949,N_17123);
nor U19866 (N_19866,N_15079,N_17755);
and U19867 (N_19867,N_16249,N_17145);
or U19868 (N_19868,N_15140,N_17519);
nor U19869 (N_19869,N_16837,N_17049);
or U19870 (N_19870,N_17827,N_17327);
and U19871 (N_19871,N_16544,N_17359);
and U19872 (N_19872,N_15409,N_16593);
or U19873 (N_19873,N_17008,N_15352);
and U19874 (N_19874,N_17169,N_15465);
or U19875 (N_19875,N_15560,N_15527);
and U19876 (N_19876,N_15497,N_17037);
nand U19877 (N_19877,N_16461,N_16209);
nand U19878 (N_19878,N_17950,N_15119);
and U19879 (N_19879,N_16301,N_15889);
or U19880 (N_19880,N_15951,N_15221);
and U19881 (N_19881,N_15542,N_15409);
xnor U19882 (N_19882,N_17006,N_15988);
and U19883 (N_19883,N_16625,N_15400);
or U19884 (N_19884,N_17667,N_15302);
nand U19885 (N_19885,N_16151,N_15698);
nand U19886 (N_19886,N_16775,N_17391);
or U19887 (N_19887,N_16995,N_15101);
nand U19888 (N_19888,N_16999,N_15411);
or U19889 (N_19889,N_15143,N_15258);
nand U19890 (N_19890,N_17008,N_15522);
nor U19891 (N_19891,N_17853,N_17574);
or U19892 (N_19892,N_17496,N_15221);
nor U19893 (N_19893,N_16912,N_15711);
nor U19894 (N_19894,N_17050,N_15270);
nand U19895 (N_19895,N_16984,N_16060);
nor U19896 (N_19896,N_16773,N_15538);
nand U19897 (N_19897,N_17771,N_16297);
and U19898 (N_19898,N_16338,N_15384);
and U19899 (N_19899,N_16740,N_16737);
nand U19900 (N_19900,N_16640,N_16033);
or U19901 (N_19901,N_16667,N_17575);
and U19902 (N_19902,N_17434,N_17922);
and U19903 (N_19903,N_16834,N_15452);
nor U19904 (N_19904,N_15298,N_17127);
nand U19905 (N_19905,N_17978,N_15587);
and U19906 (N_19906,N_16953,N_15670);
or U19907 (N_19907,N_17575,N_15374);
nor U19908 (N_19908,N_15570,N_16527);
or U19909 (N_19909,N_15434,N_15414);
nor U19910 (N_19910,N_16994,N_15306);
or U19911 (N_19911,N_15887,N_15473);
nand U19912 (N_19912,N_17035,N_15972);
nand U19913 (N_19913,N_15815,N_16648);
nor U19914 (N_19914,N_17102,N_15829);
and U19915 (N_19915,N_16003,N_15272);
and U19916 (N_19916,N_16339,N_16854);
and U19917 (N_19917,N_16384,N_17739);
or U19918 (N_19918,N_15904,N_16198);
nand U19919 (N_19919,N_15307,N_17933);
nor U19920 (N_19920,N_15145,N_16872);
nand U19921 (N_19921,N_15480,N_17291);
nand U19922 (N_19922,N_17326,N_16330);
xnor U19923 (N_19923,N_17155,N_16898);
nand U19924 (N_19924,N_17207,N_16148);
xor U19925 (N_19925,N_15157,N_16893);
and U19926 (N_19926,N_16907,N_17728);
nand U19927 (N_19927,N_17144,N_17916);
or U19928 (N_19928,N_15191,N_16558);
nor U19929 (N_19929,N_16339,N_15989);
or U19930 (N_19930,N_16161,N_15963);
nor U19931 (N_19931,N_15443,N_15131);
or U19932 (N_19932,N_15107,N_15598);
and U19933 (N_19933,N_16593,N_17751);
nor U19934 (N_19934,N_17714,N_17924);
xnor U19935 (N_19935,N_15406,N_16977);
nor U19936 (N_19936,N_17986,N_17912);
and U19937 (N_19937,N_17062,N_15980);
nor U19938 (N_19938,N_15627,N_17600);
nand U19939 (N_19939,N_15433,N_16744);
nand U19940 (N_19940,N_16948,N_15529);
or U19941 (N_19941,N_17253,N_17028);
nand U19942 (N_19942,N_15321,N_17058);
and U19943 (N_19943,N_16891,N_16448);
or U19944 (N_19944,N_17031,N_16718);
and U19945 (N_19945,N_16363,N_15320);
nor U19946 (N_19946,N_16805,N_17111);
nand U19947 (N_19947,N_15300,N_17903);
nand U19948 (N_19948,N_16978,N_16615);
and U19949 (N_19949,N_16289,N_15356);
nor U19950 (N_19950,N_17567,N_15181);
nor U19951 (N_19951,N_15739,N_16159);
or U19952 (N_19952,N_16897,N_16406);
and U19953 (N_19953,N_15470,N_16171);
and U19954 (N_19954,N_16200,N_16093);
or U19955 (N_19955,N_17014,N_17446);
xnor U19956 (N_19956,N_15355,N_15283);
or U19957 (N_19957,N_16991,N_17764);
and U19958 (N_19958,N_15737,N_15914);
and U19959 (N_19959,N_15133,N_16512);
nand U19960 (N_19960,N_17764,N_16781);
and U19961 (N_19961,N_16829,N_16804);
nor U19962 (N_19962,N_17195,N_17018);
or U19963 (N_19963,N_16843,N_16818);
or U19964 (N_19964,N_15734,N_17432);
or U19965 (N_19965,N_16309,N_15647);
nand U19966 (N_19966,N_15621,N_15654);
nor U19967 (N_19967,N_15679,N_16634);
nor U19968 (N_19968,N_16983,N_15942);
and U19969 (N_19969,N_16535,N_17269);
nand U19970 (N_19970,N_17175,N_17299);
or U19971 (N_19971,N_15282,N_15880);
xor U19972 (N_19972,N_15427,N_16479);
xnor U19973 (N_19973,N_15429,N_16648);
nor U19974 (N_19974,N_16632,N_15547);
nor U19975 (N_19975,N_16264,N_17411);
nand U19976 (N_19976,N_15138,N_17192);
or U19977 (N_19977,N_15959,N_15066);
and U19978 (N_19978,N_17268,N_17049);
or U19979 (N_19979,N_17040,N_15799);
nor U19980 (N_19980,N_16443,N_15300);
or U19981 (N_19981,N_15304,N_16740);
or U19982 (N_19982,N_17648,N_15365);
nand U19983 (N_19983,N_16727,N_16073);
or U19984 (N_19984,N_15094,N_16069);
xor U19985 (N_19985,N_15455,N_15659);
nand U19986 (N_19986,N_15572,N_16720);
nor U19987 (N_19987,N_16500,N_17313);
nand U19988 (N_19988,N_16208,N_16530);
nor U19989 (N_19989,N_17053,N_16242);
nor U19990 (N_19990,N_15783,N_15738);
or U19991 (N_19991,N_15594,N_16290);
or U19992 (N_19992,N_15480,N_16201);
nand U19993 (N_19993,N_16340,N_17823);
nor U19994 (N_19994,N_17928,N_15713);
nor U19995 (N_19995,N_16933,N_17264);
nor U19996 (N_19996,N_16337,N_17683);
nor U19997 (N_19997,N_16442,N_17850);
or U19998 (N_19998,N_16504,N_16978);
nand U19999 (N_19999,N_16045,N_16426);
and U20000 (N_20000,N_16144,N_15594);
xnor U20001 (N_20001,N_16447,N_16125);
nand U20002 (N_20002,N_17078,N_16007);
nor U20003 (N_20003,N_16259,N_17853);
nor U20004 (N_20004,N_16724,N_16830);
nor U20005 (N_20005,N_16741,N_17266);
nor U20006 (N_20006,N_17586,N_15665);
nor U20007 (N_20007,N_16070,N_15135);
nor U20008 (N_20008,N_17755,N_16312);
and U20009 (N_20009,N_16559,N_16827);
and U20010 (N_20010,N_16410,N_15611);
nor U20011 (N_20011,N_17784,N_15782);
or U20012 (N_20012,N_16657,N_16459);
and U20013 (N_20013,N_16177,N_16575);
nand U20014 (N_20014,N_17745,N_15262);
and U20015 (N_20015,N_15622,N_17623);
nor U20016 (N_20016,N_17926,N_17600);
and U20017 (N_20017,N_16739,N_15124);
nand U20018 (N_20018,N_16861,N_16275);
and U20019 (N_20019,N_15295,N_17376);
and U20020 (N_20020,N_16389,N_15775);
nand U20021 (N_20021,N_17576,N_15349);
or U20022 (N_20022,N_16504,N_16313);
nor U20023 (N_20023,N_16423,N_15488);
and U20024 (N_20024,N_17106,N_16730);
xnor U20025 (N_20025,N_15372,N_17787);
nand U20026 (N_20026,N_15454,N_15179);
nand U20027 (N_20027,N_15726,N_15437);
or U20028 (N_20028,N_16994,N_16500);
nand U20029 (N_20029,N_17684,N_16335);
or U20030 (N_20030,N_17161,N_16494);
nor U20031 (N_20031,N_16687,N_16192);
or U20032 (N_20032,N_15994,N_17178);
nand U20033 (N_20033,N_17524,N_15587);
nand U20034 (N_20034,N_17708,N_17040);
and U20035 (N_20035,N_16945,N_15552);
or U20036 (N_20036,N_15986,N_16762);
nand U20037 (N_20037,N_17987,N_15454);
nand U20038 (N_20038,N_16049,N_16595);
or U20039 (N_20039,N_16725,N_17501);
or U20040 (N_20040,N_16893,N_15093);
and U20041 (N_20041,N_17718,N_17650);
nand U20042 (N_20042,N_17330,N_17647);
and U20043 (N_20043,N_16901,N_17940);
xor U20044 (N_20044,N_16648,N_17417);
or U20045 (N_20045,N_17171,N_17924);
nand U20046 (N_20046,N_15917,N_15582);
or U20047 (N_20047,N_15830,N_17853);
nand U20048 (N_20048,N_15315,N_16368);
nand U20049 (N_20049,N_15285,N_16998);
and U20050 (N_20050,N_16440,N_17355);
nand U20051 (N_20051,N_15342,N_15824);
and U20052 (N_20052,N_15351,N_15478);
and U20053 (N_20053,N_17636,N_17021);
nor U20054 (N_20054,N_15642,N_17216);
xor U20055 (N_20055,N_17970,N_16289);
nor U20056 (N_20056,N_16100,N_16473);
and U20057 (N_20057,N_16794,N_16039);
nor U20058 (N_20058,N_15093,N_17270);
or U20059 (N_20059,N_15897,N_17340);
nand U20060 (N_20060,N_17151,N_16043);
and U20061 (N_20061,N_16499,N_15306);
nor U20062 (N_20062,N_16185,N_15066);
nand U20063 (N_20063,N_16480,N_16134);
and U20064 (N_20064,N_15928,N_15373);
or U20065 (N_20065,N_17890,N_16530);
nor U20066 (N_20066,N_15178,N_17056);
and U20067 (N_20067,N_15509,N_17834);
xor U20068 (N_20068,N_16972,N_15813);
nor U20069 (N_20069,N_17933,N_17529);
nor U20070 (N_20070,N_16005,N_17016);
nor U20071 (N_20071,N_16254,N_17070);
nor U20072 (N_20072,N_16694,N_15097);
nor U20073 (N_20073,N_16498,N_15585);
and U20074 (N_20074,N_17704,N_16043);
nor U20075 (N_20075,N_16602,N_15615);
and U20076 (N_20076,N_15907,N_16236);
nor U20077 (N_20077,N_16503,N_15704);
xnor U20078 (N_20078,N_16084,N_16983);
nor U20079 (N_20079,N_15127,N_17977);
or U20080 (N_20080,N_15658,N_17947);
and U20081 (N_20081,N_17028,N_16765);
nor U20082 (N_20082,N_16735,N_17332);
and U20083 (N_20083,N_16951,N_15288);
nor U20084 (N_20084,N_15465,N_15298);
and U20085 (N_20085,N_15365,N_15754);
or U20086 (N_20086,N_17119,N_15908);
nor U20087 (N_20087,N_16006,N_15839);
and U20088 (N_20088,N_15106,N_15121);
xnor U20089 (N_20089,N_17133,N_15463);
xnor U20090 (N_20090,N_16455,N_15006);
or U20091 (N_20091,N_15846,N_17687);
nor U20092 (N_20092,N_15915,N_15615);
xor U20093 (N_20093,N_17709,N_17387);
nor U20094 (N_20094,N_16895,N_16839);
nor U20095 (N_20095,N_15557,N_15597);
nor U20096 (N_20096,N_17376,N_17467);
nor U20097 (N_20097,N_16343,N_17629);
nor U20098 (N_20098,N_17697,N_16988);
and U20099 (N_20099,N_15339,N_15147);
nor U20100 (N_20100,N_15816,N_16295);
nor U20101 (N_20101,N_16436,N_15232);
or U20102 (N_20102,N_15975,N_17923);
nand U20103 (N_20103,N_16941,N_16425);
nor U20104 (N_20104,N_15334,N_15647);
and U20105 (N_20105,N_17410,N_16307);
and U20106 (N_20106,N_16387,N_17586);
nand U20107 (N_20107,N_15493,N_17543);
nor U20108 (N_20108,N_16562,N_15189);
nor U20109 (N_20109,N_17104,N_17681);
nand U20110 (N_20110,N_16638,N_17471);
nand U20111 (N_20111,N_16716,N_15760);
or U20112 (N_20112,N_16415,N_16014);
and U20113 (N_20113,N_17655,N_17095);
nand U20114 (N_20114,N_16121,N_16916);
nor U20115 (N_20115,N_16459,N_15309);
xnor U20116 (N_20116,N_16585,N_17302);
and U20117 (N_20117,N_16888,N_17284);
nand U20118 (N_20118,N_15759,N_17169);
and U20119 (N_20119,N_17160,N_17657);
and U20120 (N_20120,N_17932,N_16047);
or U20121 (N_20121,N_17960,N_16968);
xor U20122 (N_20122,N_16311,N_16607);
or U20123 (N_20123,N_16981,N_16056);
and U20124 (N_20124,N_17506,N_16161);
nand U20125 (N_20125,N_17375,N_15552);
nand U20126 (N_20126,N_15662,N_16263);
nor U20127 (N_20127,N_17868,N_16991);
nor U20128 (N_20128,N_16672,N_15396);
and U20129 (N_20129,N_15483,N_15475);
nor U20130 (N_20130,N_15374,N_16705);
and U20131 (N_20131,N_16877,N_16023);
nand U20132 (N_20132,N_15021,N_16791);
nor U20133 (N_20133,N_17023,N_16903);
nor U20134 (N_20134,N_15477,N_15346);
and U20135 (N_20135,N_15073,N_16356);
nor U20136 (N_20136,N_15721,N_16425);
or U20137 (N_20137,N_16758,N_17589);
nor U20138 (N_20138,N_15536,N_16004);
nor U20139 (N_20139,N_15240,N_16743);
nand U20140 (N_20140,N_17250,N_17986);
or U20141 (N_20141,N_15193,N_15899);
xnor U20142 (N_20142,N_16779,N_15035);
and U20143 (N_20143,N_16183,N_16843);
nand U20144 (N_20144,N_17825,N_17864);
and U20145 (N_20145,N_17846,N_16451);
nor U20146 (N_20146,N_15758,N_17870);
and U20147 (N_20147,N_16920,N_17470);
nor U20148 (N_20148,N_16188,N_15128);
or U20149 (N_20149,N_15601,N_15470);
nand U20150 (N_20150,N_16950,N_15525);
and U20151 (N_20151,N_16679,N_17699);
or U20152 (N_20152,N_15437,N_17495);
and U20153 (N_20153,N_15515,N_15672);
nor U20154 (N_20154,N_17158,N_17773);
and U20155 (N_20155,N_17007,N_15674);
and U20156 (N_20156,N_15371,N_15161);
nand U20157 (N_20157,N_17243,N_15469);
and U20158 (N_20158,N_17287,N_15451);
or U20159 (N_20159,N_15264,N_17858);
or U20160 (N_20160,N_15552,N_17191);
and U20161 (N_20161,N_15957,N_17852);
and U20162 (N_20162,N_17449,N_16151);
and U20163 (N_20163,N_17052,N_15805);
and U20164 (N_20164,N_16501,N_17221);
nor U20165 (N_20165,N_16591,N_17160);
nor U20166 (N_20166,N_15250,N_15677);
and U20167 (N_20167,N_15499,N_16403);
and U20168 (N_20168,N_15933,N_16288);
or U20169 (N_20169,N_15402,N_15412);
xor U20170 (N_20170,N_17070,N_16347);
xor U20171 (N_20171,N_17214,N_15944);
nor U20172 (N_20172,N_16763,N_17073);
and U20173 (N_20173,N_17527,N_15789);
or U20174 (N_20174,N_17622,N_15817);
and U20175 (N_20175,N_16603,N_16068);
and U20176 (N_20176,N_15970,N_17514);
and U20177 (N_20177,N_17248,N_17776);
nor U20178 (N_20178,N_16836,N_17371);
and U20179 (N_20179,N_17566,N_15155);
nor U20180 (N_20180,N_16188,N_15115);
or U20181 (N_20181,N_16963,N_17928);
nor U20182 (N_20182,N_16021,N_17907);
and U20183 (N_20183,N_16038,N_16515);
and U20184 (N_20184,N_17543,N_15351);
nor U20185 (N_20185,N_16048,N_15628);
nor U20186 (N_20186,N_17991,N_15832);
nor U20187 (N_20187,N_17869,N_16286);
nand U20188 (N_20188,N_17558,N_17124);
or U20189 (N_20189,N_16043,N_16193);
nor U20190 (N_20190,N_16673,N_15602);
xor U20191 (N_20191,N_15713,N_15836);
nor U20192 (N_20192,N_17044,N_16520);
or U20193 (N_20193,N_16348,N_16814);
and U20194 (N_20194,N_15168,N_16651);
xnor U20195 (N_20195,N_16743,N_17833);
nor U20196 (N_20196,N_17388,N_15897);
nand U20197 (N_20197,N_16296,N_17644);
and U20198 (N_20198,N_17299,N_16993);
or U20199 (N_20199,N_17131,N_15425);
and U20200 (N_20200,N_16381,N_15328);
nor U20201 (N_20201,N_15020,N_17255);
xnor U20202 (N_20202,N_16664,N_15773);
xnor U20203 (N_20203,N_17455,N_17550);
and U20204 (N_20204,N_15888,N_17645);
nand U20205 (N_20205,N_15308,N_16964);
or U20206 (N_20206,N_15007,N_16494);
nor U20207 (N_20207,N_16187,N_17926);
nand U20208 (N_20208,N_17363,N_16953);
and U20209 (N_20209,N_17849,N_16216);
nand U20210 (N_20210,N_17336,N_15676);
nand U20211 (N_20211,N_15983,N_15885);
nor U20212 (N_20212,N_17591,N_15466);
nand U20213 (N_20213,N_15508,N_16716);
and U20214 (N_20214,N_17982,N_16568);
nor U20215 (N_20215,N_17771,N_16566);
nand U20216 (N_20216,N_16093,N_15868);
nand U20217 (N_20217,N_16235,N_15974);
nand U20218 (N_20218,N_15949,N_17550);
nand U20219 (N_20219,N_16244,N_15539);
nand U20220 (N_20220,N_16390,N_15266);
nor U20221 (N_20221,N_15104,N_16242);
or U20222 (N_20222,N_16028,N_17124);
or U20223 (N_20223,N_16094,N_17825);
nand U20224 (N_20224,N_15794,N_15108);
xor U20225 (N_20225,N_16961,N_16553);
and U20226 (N_20226,N_17805,N_17240);
nand U20227 (N_20227,N_16261,N_16208);
or U20228 (N_20228,N_16452,N_17374);
xor U20229 (N_20229,N_16701,N_17164);
and U20230 (N_20230,N_16780,N_15852);
or U20231 (N_20231,N_16279,N_17445);
nor U20232 (N_20232,N_15869,N_17403);
nand U20233 (N_20233,N_16828,N_17860);
nor U20234 (N_20234,N_17673,N_16057);
nor U20235 (N_20235,N_17459,N_16004);
or U20236 (N_20236,N_15986,N_16428);
or U20237 (N_20237,N_15704,N_16335);
nor U20238 (N_20238,N_15931,N_17004);
nand U20239 (N_20239,N_16648,N_16301);
or U20240 (N_20240,N_15322,N_16189);
nor U20241 (N_20241,N_15715,N_15456);
nand U20242 (N_20242,N_16793,N_16585);
nor U20243 (N_20243,N_16307,N_17602);
or U20244 (N_20244,N_16045,N_15856);
and U20245 (N_20245,N_17650,N_16941);
nor U20246 (N_20246,N_17995,N_17547);
or U20247 (N_20247,N_15097,N_17866);
and U20248 (N_20248,N_17235,N_16555);
nand U20249 (N_20249,N_16100,N_17190);
nor U20250 (N_20250,N_17621,N_17719);
or U20251 (N_20251,N_16995,N_17946);
nand U20252 (N_20252,N_15243,N_17294);
and U20253 (N_20253,N_17076,N_15495);
or U20254 (N_20254,N_17508,N_16557);
and U20255 (N_20255,N_17251,N_15803);
nand U20256 (N_20256,N_16675,N_17808);
xor U20257 (N_20257,N_16363,N_15840);
xor U20258 (N_20258,N_16991,N_17102);
and U20259 (N_20259,N_16162,N_16950);
nand U20260 (N_20260,N_16399,N_17618);
or U20261 (N_20261,N_16143,N_15112);
nor U20262 (N_20262,N_17349,N_17094);
and U20263 (N_20263,N_15976,N_16014);
and U20264 (N_20264,N_16630,N_16869);
nand U20265 (N_20265,N_15301,N_16285);
nand U20266 (N_20266,N_16193,N_17193);
nor U20267 (N_20267,N_17256,N_16422);
or U20268 (N_20268,N_17533,N_17424);
xnor U20269 (N_20269,N_17265,N_15550);
or U20270 (N_20270,N_17039,N_17092);
or U20271 (N_20271,N_17467,N_17641);
and U20272 (N_20272,N_15578,N_15379);
nand U20273 (N_20273,N_17408,N_17936);
or U20274 (N_20274,N_16729,N_15785);
nand U20275 (N_20275,N_15512,N_15694);
and U20276 (N_20276,N_16479,N_16397);
nor U20277 (N_20277,N_17311,N_16145);
nor U20278 (N_20278,N_16682,N_16092);
or U20279 (N_20279,N_17262,N_15665);
nor U20280 (N_20280,N_16829,N_15676);
nor U20281 (N_20281,N_16054,N_15702);
and U20282 (N_20282,N_16406,N_17083);
or U20283 (N_20283,N_15617,N_16418);
or U20284 (N_20284,N_16088,N_16120);
xnor U20285 (N_20285,N_17191,N_16610);
nor U20286 (N_20286,N_16838,N_15921);
nand U20287 (N_20287,N_17795,N_17504);
nor U20288 (N_20288,N_17274,N_15972);
and U20289 (N_20289,N_15887,N_15216);
xnor U20290 (N_20290,N_16087,N_15288);
and U20291 (N_20291,N_15668,N_17768);
and U20292 (N_20292,N_16080,N_17598);
nor U20293 (N_20293,N_15388,N_17652);
nor U20294 (N_20294,N_17180,N_16537);
nor U20295 (N_20295,N_17848,N_15021);
nand U20296 (N_20296,N_15462,N_15684);
nor U20297 (N_20297,N_16305,N_16780);
xnor U20298 (N_20298,N_16981,N_15956);
and U20299 (N_20299,N_15516,N_15048);
and U20300 (N_20300,N_15794,N_15956);
nor U20301 (N_20301,N_16576,N_15399);
and U20302 (N_20302,N_17452,N_15920);
nor U20303 (N_20303,N_15386,N_15763);
nor U20304 (N_20304,N_17002,N_17492);
nand U20305 (N_20305,N_17015,N_16680);
or U20306 (N_20306,N_15251,N_15480);
xnor U20307 (N_20307,N_17750,N_16141);
xor U20308 (N_20308,N_17285,N_16389);
nor U20309 (N_20309,N_17070,N_17876);
nand U20310 (N_20310,N_15636,N_15508);
and U20311 (N_20311,N_17854,N_17494);
nor U20312 (N_20312,N_15348,N_15769);
or U20313 (N_20313,N_15509,N_16121);
or U20314 (N_20314,N_15935,N_16317);
or U20315 (N_20315,N_15527,N_16148);
and U20316 (N_20316,N_15839,N_15453);
or U20317 (N_20317,N_15676,N_17307);
nor U20318 (N_20318,N_15409,N_17551);
nor U20319 (N_20319,N_15131,N_16678);
nand U20320 (N_20320,N_15393,N_15742);
xor U20321 (N_20321,N_17652,N_16187);
or U20322 (N_20322,N_16927,N_15671);
nand U20323 (N_20323,N_17034,N_15865);
or U20324 (N_20324,N_15035,N_17382);
nand U20325 (N_20325,N_15535,N_16389);
and U20326 (N_20326,N_17044,N_17893);
xor U20327 (N_20327,N_16054,N_15198);
or U20328 (N_20328,N_15493,N_15650);
nand U20329 (N_20329,N_17701,N_15632);
and U20330 (N_20330,N_17822,N_17542);
nor U20331 (N_20331,N_16099,N_16554);
nor U20332 (N_20332,N_15405,N_16403);
nand U20333 (N_20333,N_16644,N_16879);
or U20334 (N_20334,N_16913,N_16333);
and U20335 (N_20335,N_16322,N_16196);
nand U20336 (N_20336,N_15729,N_15484);
xnor U20337 (N_20337,N_17331,N_17577);
nor U20338 (N_20338,N_17789,N_15953);
and U20339 (N_20339,N_17280,N_15974);
or U20340 (N_20340,N_17572,N_17352);
nand U20341 (N_20341,N_17234,N_17230);
nor U20342 (N_20342,N_15085,N_15866);
nor U20343 (N_20343,N_17811,N_15577);
or U20344 (N_20344,N_15174,N_15625);
or U20345 (N_20345,N_16151,N_16122);
and U20346 (N_20346,N_17547,N_16047);
nand U20347 (N_20347,N_15933,N_16279);
nor U20348 (N_20348,N_17520,N_17084);
xnor U20349 (N_20349,N_15182,N_15335);
or U20350 (N_20350,N_15753,N_17559);
and U20351 (N_20351,N_16190,N_16408);
or U20352 (N_20352,N_15957,N_16827);
nor U20353 (N_20353,N_16116,N_17832);
nand U20354 (N_20354,N_17734,N_16237);
and U20355 (N_20355,N_15825,N_17233);
xnor U20356 (N_20356,N_16979,N_15391);
or U20357 (N_20357,N_17626,N_15205);
or U20358 (N_20358,N_16120,N_16577);
nand U20359 (N_20359,N_15174,N_15333);
nor U20360 (N_20360,N_17784,N_16648);
and U20361 (N_20361,N_16361,N_16817);
and U20362 (N_20362,N_16895,N_17120);
nor U20363 (N_20363,N_15517,N_15785);
or U20364 (N_20364,N_17480,N_17976);
and U20365 (N_20365,N_16371,N_16999);
and U20366 (N_20366,N_17008,N_15890);
and U20367 (N_20367,N_17628,N_17023);
nand U20368 (N_20368,N_17907,N_17538);
and U20369 (N_20369,N_16679,N_15450);
nand U20370 (N_20370,N_17560,N_16568);
xor U20371 (N_20371,N_17452,N_16857);
and U20372 (N_20372,N_15841,N_17569);
or U20373 (N_20373,N_15400,N_15305);
xor U20374 (N_20374,N_17550,N_16934);
nor U20375 (N_20375,N_15807,N_16074);
nor U20376 (N_20376,N_17539,N_16992);
nor U20377 (N_20377,N_17191,N_17625);
and U20378 (N_20378,N_16784,N_15259);
nand U20379 (N_20379,N_17997,N_15493);
and U20380 (N_20380,N_17352,N_17391);
and U20381 (N_20381,N_15892,N_17548);
nor U20382 (N_20382,N_15565,N_15882);
or U20383 (N_20383,N_16017,N_16973);
or U20384 (N_20384,N_15221,N_15674);
nand U20385 (N_20385,N_15128,N_16690);
or U20386 (N_20386,N_17610,N_16427);
or U20387 (N_20387,N_17034,N_16792);
or U20388 (N_20388,N_15107,N_15152);
nor U20389 (N_20389,N_16111,N_16115);
xor U20390 (N_20390,N_16110,N_15260);
or U20391 (N_20391,N_17886,N_16247);
nor U20392 (N_20392,N_15970,N_15921);
nor U20393 (N_20393,N_16552,N_15293);
and U20394 (N_20394,N_16968,N_17034);
nand U20395 (N_20395,N_16605,N_15878);
or U20396 (N_20396,N_16631,N_17927);
and U20397 (N_20397,N_15071,N_15030);
and U20398 (N_20398,N_17508,N_17547);
nor U20399 (N_20399,N_16163,N_17265);
nor U20400 (N_20400,N_16769,N_16146);
nor U20401 (N_20401,N_16585,N_15882);
nor U20402 (N_20402,N_17164,N_15298);
nor U20403 (N_20403,N_16099,N_16715);
nor U20404 (N_20404,N_15852,N_17006);
and U20405 (N_20405,N_15957,N_16782);
or U20406 (N_20406,N_15268,N_15914);
or U20407 (N_20407,N_15009,N_15139);
nor U20408 (N_20408,N_16476,N_17263);
nor U20409 (N_20409,N_16138,N_16927);
nor U20410 (N_20410,N_17065,N_17816);
and U20411 (N_20411,N_16966,N_17661);
nor U20412 (N_20412,N_17560,N_15158);
nand U20413 (N_20413,N_16659,N_16973);
or U20414 (N_20414,N_16803,N_17683);
xnor U20415 (N_20415,N_15727,N_16402);
and U20416 (N_20416,N_15775,N_15400);
xnor U20417 (N_20417,N_15963,N_17650);
nand U20418 (N_20418,N_17410,N_17279);
or U20419 (N_20419,N_16206,N_17781);
nand U20420 (N_20420,N_16463,N_17708);
and U20421 (N_20421,N_15328,N_17721);
nor U20422 (N_20422,N_15640,N_16333);
nand U20423 (N_20423,N_15219,N_17330);
nand U20424 (N_20424,N_15458,N_15725);
nor U20425 (N_20425,N_15650,N_15275);
nor U20426 (N_20426,N_17163,N_17961);
or U20427 (N_20427,N_15176,N_17189);
nor U20428 (N_20428,N_17889,N_16544);
or U20429 (N_20429,N_17276,N_16526);
and U20430 (N_20430,N_17848,N_15492);
nor U20431 (N_20431,N_17841,N_15792);
nor U20432 (N_20432,N_15902,N_16156);
nand U20433 (N_20433,N_16475,N_17605);
nor U20434 (N_20434,N_15267,N_15596);
nand U20435 (N_20435,N_16767,N_15148);
and U20436 (N_20436,N_16769,N_15005);
xnor U20437 (N_20437,N_16732,N_16202);
nand U20438 (N_20438,N_15635,N_16351);
or U20439 (N_20439,N_15434,N_17900);
nand U20440 (N_20440,N_16076,N_16626);
nand U20441 (N_20441,N_15406,N_16466);
nand U20442 (N_20442,N_17380,N_15188);
xnor U20443 (N_20443,N_17133,N_17433);
xnor U20444 (N_20444,N_15305,N_15366);
nor U20445 (N_20445,N_15845,N_16659);
nand U20446 (N_20446,N_15882,N_17837);
nor U20447 (N_20447,N_17254,N_16838);
nor U20448 (N_20448,N_16577,N_15753);
nand U20449 (N_20449,N_15280,N_17473);
nand U20450 (N_20450,N_17814,N_15150);
or U20451 (N_20451,N_15037,N_15855);
and U20452 (N_20452,N_16808,N_17559);
and U20453 (N_20453,N_17732,N_16116);
and U20454 (N_20454,N_17561,N_15158);
nor U20455 (N_20455,N_16376,N_16821);
and U20456 (N_20456,N_16670,N_15338);
nor U20457 (N_20457,N_15113,N_15461);
xnor U20458 (N_20458,N_15593,N_15050);
and U20459 (N_20459,N_16094,N_17315);
xor U20460 (N_20460,N_15387,N_17880);
nor U20461 (N_20461,N_17501,N_15148);
or U20462 (N_20462,N_16373,N_15027);
nand U20463 (N_20463,N_16864,N_16241);
or U20464 (N_20464,N_16562,N_15266);
xor U20465 (N_20465,N_15625,N_15921);
nand U20466 (N_20466,N_15180,N_15301);
nand U20467 (N_20467,N_15867,N_15621);
or U20468 (N_20468,N_15576,N_16389);
or U20469 (N_20469,N_17652,N_15113);
or U20470 (N_20470,N_16536,N_17670);
or U20471 (N_20471,N_17124,N_15988);
nor U20472 (N_20472,N_15764,N_15783);
and U20473 (N_20473,N_17592,N_16942);
or U20474 (N_20474,N_16939,N_17981);
or U20475 (N_20475,N_17317,N_15018);
and U20476 (N_20476,N_16730,N_16828);
or U20477 (N_20477,N_17216,N_15794);
or U20478 (N_20478,N_17504,N_16843);
or U20479 (N_20479,N_15055,N_15336);
and U20480 (N_20480,N_17725,N_15493);
nor U20481 (N_20481,N_17862,N_15606);
nand U20482 (N_20482,N_16300,N_17155);
or U20483 (N_20483,N_15663,N_17998);
xor U20484 (N_20484,N_15375,N_15662);
nand U20485 (N_20485,N_15963,N_15627);
or U20486 (N_20486,N_16159,N_16742);
and U20487 (N_20487,N_15088,N_15270);
and U20488 (N_20488,N_15152,N_16732);
nand U20489 (N_20489,N_15230,N_16226);
nor U20490 (N_20490,N_15120,N_16396);
or U20491 (N_20491,N_17573,N_16474);
or U20492 (N_20492,N_17682,N_16204);
nor U20493 (N_20493,N_17519,N_15697);
nand U20494 (N_20494,N_16312,N_16662);
and U20495 (N_20495,N_16189,N_17063);
nor U20496 (N_20496,N_15099,N_15522);
nor U20497 (N_20497,N_17519,N_17625);
and U20498 (N_20498,N_16361,N_16484);
nor U20499 (N_20499,N_17167,N_16322);
nor U20500 (N_20500,N_16620,N_17819);
and U20501 (N_20501,N_17484,N_15248);
or U20502 (N_20502,N_16218,N_15593);
and U20503 (N_20503,N_16999,N_17214);
and U20504 (N_20504,N_15415,N_16563);
or U20505 (N_20505,N_16306,N_16066);
nor U20506 (N_20506,N_16840,N_15421);
nor U20507 (N_20507,N_16941,N_17922);
and U20508 (N_20508,N_16485,N_17669);
or U20509 (N_20509,N_16338,N_16464);
or U20510 (N_20510,N_17851,N_16797);
xnor U20511 (N_20511,N_17243,N_16961);
nand U20512 (N_20512,N_15262,N_17484);
xor U20513 (N_20513,N_17961,N_17045);
nand U20514 (N_20514,N_17301,N_15957);
and U20515 (N_20515,N_15471,N_17073);
nand U20516 (N_20516,N_17813,N_17846);
and U20517 (N_20517,N_17333,N_17825);
and U20518 (N_20518,N_17530,N_17452);
and U20519 (N_20519,N_16832,N_16372);
and U20520 (N_20520,N_16391,N_17843);
or U20521 (N_20521,N_16956,N_16692);
nor U20522 (N_20522,N_17282,N_15361);
or U20523 (N_20523,N_15247,N_15185);
nand U20524 (N_20524,N_15413,N_15712);
and U20525 (N_20525,N_15893,N_15857);
nand U20526 (N_20526,N_16365,N_17447);
and U20527 (N_20527,N_15631,N_15917);
nand U20528 (N_20528,N_16048,N_16575);
or U20529 (N_20529,N_15785,N_17119);
nand U20530 (N_20530,N_17137,N_16970);
nor U20531 (N_20531,N_17038,N_15765);
or U20532 (N_20532,N_16383,N_15793);
and U20533 (N_20533,N_15519,N_17202);
nor U20534 (N_20534,N_15146,N_17743);
and U20535 (N_20535,N_17568,N_16923);
xor U20536 (N_20536,N_15346,N_15777);
nor U20537 (N_20537,N_17347,N_16928);
and U20538 (N_20538,N_17497,N_17254);
or U20539 (N_20539,N_15074,N_17187);
or U20540 (N_20540,N_17882,N_17787);
and U20541 (N_20541,N_17654,N_15242);
and U20542 (N_20542,N_17095,N_17826);
and U20543 (N_20543,N_15273,N_17166);
or U20544 (N_20544,N_15884,N_15261);
nor U20545 (N_20545,N_15654,N_16246);
xnor U20546 (N_20546,N_16919,N_15807);
and U20547 (N_20547,N_16286,N_16509);
nor U20548 (N_20548,N_15341,N_16557);
or U20549 (N_20549,N_16670,N_17211);
nor U20550 (N_20550,N_16494,N_15845);
nand U20551 (N_20551,N_17329,N_17070);
or U20552 (N_20552,N_17954,N_15969);
or U20553 (N_20553,N_16494,N_16027);
and U20554 (N_20554,N_17626,N_17181);
nand U20555 (N_20555,N_17677,N_17840);
nor U20556 (N_20556,N_15515,N_16946);
nor U20557 (N_20557,N_16287,N_17751);
nor U20558 (N_20558,N_17628,N_16878);
nor U20559 (N_20559,N_17685,N_16170);
or U20560 (N_20560,N_16651,N_17845);
nand U20561 (N_20561,N_17079,N_15973);
nand U20562 (N_20562,N_16097,N_17177);
xor U20563 (N_20563,N_15514,N_16304);
and U20564 (N_20564,N_17038,N_16435);
nand U20565 (N_20565,N_16978,N_17042);
xor U20566 (N_20566,N_15356,N_15583);
and U20567 (N_20567,N_15386,N_17944);
and U20568 (N_20568,N_15891,N_17368);
xnor U20569 (N_20569,N_17505,N_15285);
nand U20570 (N_20570,N_15540,N_17081);
nor U20571 (N_20571,N_15226,N_17069);
and U20572 (N_20572,N_17549,N_16294);
nor U20573 (N_20573,N_16505,N_15625);
nor U20574 (N_20574,N_16050,N_17168);
xor U20575 (N_20575,N_17431,N_17713);
xnor U20576 (N_20576,N_17203,N_16465);
and U20577 (N_20577,N_17123,N_17318);
and U20578 (N_20578,N_15746,N_15339);
nand U20579 (N_20579,N_15611,N_17332);
or U20580 (N_20580,N_17633,N_15461);
nand U20581 (N_20581,N_17340,N_16084);
or U20582 (N_20582,N_15322,N_16609);
or U20583 (N_20583,N_17057,N_16668);
and U20584 (N_20584,N_17992,N_17696);
nor U20585 (N_20585,N_15222,N_16493);
or U20586 (N_20586,N_16804,N_15430);
nand U20587 (N_20587,N_15882,N_15020);
nand U20588 (N_20588,N_15108,N_15451);
xnor U20589 (N_20589,N_17508,N_16866);
nand U20590 (N_20590,N_16243,N_17928);
and U20591 (N_20591,N_15087,N_15062);
and U20592 (N_20592,N_17049,N_15906);
nor U20593 (N_20593,N_15100,N_15368);
xnor U20594 (N_20594,N_15473,N_17664);
nand U20595 (N_20595,N_17881,N_17891);
and U20596 (N_20596,N_17409,N_15973);
nand U20597 (N_20597,N_17419,N_15353);
nand U20598 (N_20598,N_15481,N_17914);
or U20599 (N_20599,N_17663,N_16256);
or U20600 (N_20600,N_17309,N_15810);
and U20601 (N_20601,N_16437,N_15519);
nand U20602 (N_20602,N_17389,N_16446);
or U20603 (N_20603,N_16657,N_16575);
xor U20604 (N_20604,N_16754,N_17640);
and U20605 (N_20605,N_17806,N_17836);
or U20606 (N_20606,N_15664,N_17691);
nor U20607 (N_20607,N_17276,N_17576);
or U20608 (N_20608,N_16161,N_15111);
nor U20609 (N_20609,N_16769,N_15977);
or U20610 (N_20610,N_17220,N_17789);
nand U20611 (N_20611,N_16220,N_16216);
or U20612 (N_20612,N_17018,N_16240);
xor U20613 (N_20613,N_17456,N_15516);
nand U20614 (N_20614,N_16274,N_17567);
or U20615 (N_20615,N_16061,N_17564);
and U20616 (N_20616,N_16569,N_17857);
and U20617 (N_20617,N_16747,N_17276);
and U20618 (N_20618,N_15143,N_17373);
nor U20619 (N_20619,N_15466,N_15818);
and U20620 (N_20620,N_15710,N_17586);
or U20621 (N_20621,N_15077,N_17933);
nand U20622 (N_20622,N_15426,N_17242);
xnor U20623 (N_20623,N_16266,N_17310);
nand U20624 (N_20624,N_17639,N_17980);
nor U20625 (N_20625,N_17690,N_15223);
or U20626 (N_20626,N_15230,N_17961);
and U20627 (N_20627,N_17789,N_17390);
and U20628 (N_20628,N_16475,N_15653);
and U20629 (N_20629,N_16687,N_17171);
and U20630 (N_20630,N_15157,N_15746);
and U20631 (N_20631,N_15693,N_15723);
nand U20632 (N_20632,N_15120,N_16471);
or U20633 (N_20633,N_16096,N_16213);
nor U20634 (N_20634,N_16636,N_17241);
nand U20635 (N_20635,N_15880,N_17953);
nand U20636 (N_20636,N_15935,N_17568);
nand U20637 (N_20637,N_17419,N_16746);
or U20638 (N_20638,N_15088,N_15531);
nor U20639 (N_20639,N_16434,N_16041);
or U20640 (N_20640,N_15672,N_15248);
xor U20641 (N_20641,N_15077,N_15522);
nor U20642 (N_20642,N_16876,N_16063);
nor U20643 (N_20643,N_16051,N_16913);
and U20644 (N_20644,N_17127,N_17424);
nor U20645 (N_20645,N_16242,N_17253);
or U20646 (N_20646,N_15883,N_15845);
nor U20647 (N_20647,N_16466,N_17841);
or U20648 (N_20648,N_16169,N_15532);
nor U20649 (N_20649,N_15644,N_16818);
nand U20650 (N_20650,N_17468,N_15671);
or U20651 (N_20651,N_17689,N_17783);
and U20652 (N_20652,N_15394,N_15410);
or U20653 (N_20653,N_17536,N_16591);
nor U20654 (N_20654,N_15712,N_15505);
xnor U20655 (N_20655,N_16041,N_17321);
or U20656 (N_20656,N_17631,N_17656);
nor U20657 (N_20657,N_15407,N_15875);
or U20658 (N_20658,N_15633,N_16024);
and U20659 (N_20659,N_17121,N_16983);
nand U20660 (N_20660,N_15758,N_17317);
and U20661 (N_20661,N_16870,N_16340);
nor U20662 (N_20662,N_16400,N_17987);
or U20663 (N_20663,N_17162,N_15205);
or U20664 (N_20664,N_17455,N_15706);
or U20665 (N_20665,N_15992,N_16552);
nor U20666 (N_20666,N_16006,N_17338);
nand U20667 (N_20667,N_16697,N_15807);
and U20668 (N_20668,N_16286,N_16652);
or U20669 (N_20669,N_16887,N_15797);
nand U20670 (N_20670,N_17922,N_17314);
and U20671 (N_20671,N_17786,N_17339);
or U20672 (N_20672,N_16814,N_16152);
nand U20673 (N_20673,N_17898,N_17141);
nor U20674 (N_20674,N_15764,N_17176);
nand U20675 (N_20675,N_16880,N_15424);
and U20676 (N_20676,N_17739,N_15307);
or U20677 (N_20677,N_15066,N_15211);
or U20678 (N_20678,N_15377,N_15869);
xor U20679 (N_20679,N_16347,N_16423);
nand U20680 (N_20680,N_17659,N_16814);
nor U20681 (N_20681,N_16613,N_17630);
and U20682 (N_20682,N_16989,N_15040);
nand U20683 (N_20683,N_17691,N_16491);
and U20684 (N_20684,N_15416,N_16425);
nor U20685 (N_20685,N_16284,N_15451);
nor U20686 (N_20686,N_17218,N_16812);
and U20687 (N_20687,N_16906,N_15680);
nor U20688 (N_20688,N_15719,N_17584);
or U20689 (N_20689,N_17222,N_15436);
and U20690 (N_20690,N_16032,N_16479);
xnor U20691 (N_20691,N_16384,N_17973);
nand U20692 (N_20692,N_16640,N_16667);
and U20693 (N_20693,N_17858,N_17250);
and U20694 (N_20694,N_17261,N_17672);
nand U20695 (N_20695,N_17779,N_15260);
nand U20696 (N_20696,N_15576,N_17480);
xor U20697 (N_20697,N_15609,N_15005);
xor U20698 (N_20698,N_16872,N_17055);
nand U20699 (N_20699,N_16058,N_16657);
nand U20700 (N_20700,N_15317,N_17111);
and U20701 (N_20701,N_16434,N_15381);
nor U20702 (N_20702,N_16043,N_16153);
nor U20703 (N_20703,N_17654,N_17608);
nor U20704 (N_20704,N_17475,N_15139);
or U20705 (N_20705,N_15508,N_15264);
nand U20706 (N_20706,N_17079,N_15474);
or U20707 (N_20707,N_15116,N_16973);
nor U20708 (N_20708,N_17222,N_17039);
and U20709 (N_20709,N_15276,N_17270);
xor U20710 (N_20710,N_15988,N_15696);
nor U20711 (N_20711,N_15981,N_17868);
nor U20712 (N_20712,N_16583,N_16257);
or U20713 (N_20713,N_16243,N_16272);
or U20714 (N_20714,N_15094,N_16674);
or U20715 (N_20715,N_16829,N_16222);
or U20716 (N_20716,N_16271,N_17947);
and U20717 (N_20717,N_17733,N_16273);
nor U20718 (N_20718,N_15845,N_16357);
and U20719 (N_20719,N_17521,N_17512);
nand U20720 (N_20720,N_15907,N_15847);
nand U20721 (N_20721,N_16429,N_17052);
nand U20722 (N_20722,N_17278,N_15725);
or U20723 (N_20723,N_16497,N_16685);
nand U20724 (N_20724,N_15355,N_17987);
xor U20725 (N_20725,N_16616,N_17190);
nor U20726 (N_20726,N_16674,N_15829);
or U20727 (N_20727,N_17451,N_17966);
and U20728 (N_20728,N_16813,N_17469);
and U20729 (N_20729,N_15958,N_16289);
and U20730 (N_20730,N_16196,N_17450);
or U20731 (N_20731,N_16285,N_15022);
nand U20732 (N_20732,N_17346,N_16828);
nor U20733 (N_20733,N_16458,N_15231);
or U20734 (N_20734,N_17947,N_15463);
or U20735 (N_20735,N_17047,N_17507);
nand U20736 (N_20736,N_15534,N_17190);
or U20737 (N_20737,N_15345,N_15407);
or U20738 (N_20738,N_16093,N_16483);
nor U20739 (N_20739,N_17540,N_15347);
and U20740 (N_20740,N_15361,N_16914);
nand U20741 (N_20741,N_17247,N_16371);
nor U20742 (N_20742,N_16892,N_17469);
nor U20743 (N_20743,N_15272,N_17993);
nor U20744 (N_20744,N_16746,N_16160);
or U20745 (N_20745,N_16009,N_15006);
and U20746 (N_20746,N_15024,N_17019);
or U20747 (N_20747,N_17216,N_17162);
nand U20748 (N_20748,N_17955,N_16520);
nor U20749 (N_20749,N_15428,N_16199);
and U20750 (N_20750,N_17233,N_16587);
and U20751 (N_20751,N_17865,N_17041);
and U20752 (N_20752,N_15251,N_17871);
xor U20753 (N_20753,N_16365,N_15137);
nor U20754 (N_20754,N_17192,N_15886);
or U20755 (N_20755,N_15679,N_15513);
nand U20756 (N_20756,N_16674,N_17221);
and U20757 (N_20757,N_17628,N_17364);
and U20758 (N_20758,N_16882,N_17315);
and U20759 (N_20759,N_15781,N_16140);
or U20760 (N_20760,N_15373,N_16936);
or U20761 (N_20761,N_15632,N_16853);
and U20762 (N_20762,N_16470,N_17166);
nor U20763 (N_20763,N_15357,N_17534);
nor U20764 (N_20764,N_15199,N_17148);
xor U20765 (N_20765,N_17547,N_17697);
nand U20766 (N_20766,N_15102,N_17444);
xnor U20767 (N_20767,N_16012,N_16239);
nor U20768 (N_20768,N_15970,N_17965);
and U20769 (N_20769,N_15605,N_17820);
nand U20770 (N_20770,N_16002,N_17861);
xnor U20771 (N_20771,N_17135,N_15614);
nand U20772 (N_20772,N_17768,N_16700);
and U20773 (N_20773,N_15528,N_16421);
nor U20774 (N_20774,N_17767,N_17552);
nor U20775 (N_20775,N_17328,N_16287);
and U20776 (N_20776,N_17304,N_17492);
nor U20777 (N_20777,N_17540,N_16557);
nand U20778 (N_20778,N_17994,N_15071);
nor U20779 (N_20779,N_15024,N_15748);
or U20780 (N_20780,N_16114,N_17263);
nor U20781 (N_20781,N_15971,N_17445);
xor U20782 (N_20782,N_17264,N_16201);
nand U20783 (N_20783,N_16139,N_16155);
nor U20784 (N_20784,N_16278,N_16761);
nor U20785 (N_20785,N_17482,N_16940);
nand U20786 (N_20786,N_15705,N_15648);
and U20787 (N_20787,N_17101,N_15008);
xor U20788 (N_20788,N_16858,N_17162);
or U20789 (N_20789,N_15760,N_17052);
nor U20790 (N_20790,N_15106,N_17654);
nor U20791 (N_20791,N_16951,N_16872);
nor U20792 (N_20792,N_15361,N_16433);
and U20793 (N_20793,N_16886,N_15958);
nand U20794 (N_20794,N_17128,N_17968);
and U20795 (N_20795,N_16331,N_16223);
and U20796 (N_20796,N_17009,N_16429);
or U20797 (N_20797,N_15556,N_16854);
or U20798 (N_20798,N_16521,N_15602);
nand U20799 (N_20799,N_16009,N_17944);
or U20800 (N_20800,N_15814,N_15759);
nor U20801 (N_20801,N_15952,N_15131);
or U20802 (N_20802,N_17903,N_15042);
nor U20803 (N_20803,N_15625,N_15827);
and U20804 (N_20804,N_16682,N_15915);
nor U20805 (N_20805,N_16207,N_17475);
nor U20806 (N_20806,N_15232,N_17942);
nor U20807 (N_20807,N_17032,N_16421);
xor U20808 (N_20808,N_17549,N_15767);
or U20809 (N_20809,N_17976,N_16800);
or U20810 (N_20810,N_15956,N_16539);
and U20811 (N_20811,N_17693,N_16777);
nor U20812 (N_20812,N_17689,N_15423);
nor U20813 (N_20813,N_16001,N_17878);
xor U20814 (N_20814,N_17905,N_16933);
and U20815 (N_20815,N_17771,N_15931);
nand U20816 (N_20816,N_15927,N_15626);
or U20817 (N_20817,N_15034,N_15914);
and U20818 (N_20818,N_15788,N_17225);
nand U20819 (N_20819,N_17060,N_16074);
nor U20820 (N_20820,N_17795,N_17555);
nand U20821 (N_20821,N_17793,N_17346);
nor U20822 (N_20822,N_15478,N_17447);
nand U20823 (N_20823,N_15249,N_16078);
or U20824 (N_20824,N_17905,N_16920);
xor U20825 (N_20825,N_17853,N_15037);
nor U20826 (N_20826,N_17213,N_15126);
xnor U20827 (N_20827,N_16780,N_15294);
nand U20828 (N_20828,N_17267,N_15665);
or U20829 (N_20829,N_17960,N_17255);
or U20830 (N_20830,N_15947,N_15621);
xnor U20831 (N_20831,N_17278,N_16278);
nand U20832 (N_20832,N_16679,N_15904);
nor U20833 (N_20833,N_15823,N_15428);
and U20834 (N_20834,N_15305,N_16802);
nor U20835 (N_20835,N_17159,N_15954);
and U20836 (N_20836,N_15140,N_15579);
nor U20837 (N_20837,N_16466,N_17992);
and U20838 (N_20838,N_15100,N_15325);
and U20839 (N_20839,N_16247,N_15670);
xnor U20840 (N_20840,N_15555,N_16344);
nand U20841 (N_20841,N_15891,N_16614);
nand U20842 (N_20842,N_15186,N_15588);
nand U20843 (N_20843,N_17426,N_17212);
nand U20844 (N_20844,N_16894,N_15800);
or U20845 (N_20845,N_17585,N_15122);
or U20846 (N_20846,N_15849,N_15405);
nand U20847 (N_20847,N_16712,N_17856);
nand U20848 (N_20848,N_15143,N_17943);
nand U20849 (N_20849,N_16365,N_16815);
or U20850 (N_20850,N_16180,N_17895);
or U20851 (N_20851,N_15464,N_17399);
nor U20852 (N_20852,N_17987,N_16060);
and U20853 (N_20853,N_16601,N_16430);
nor U20854 (N_20854,N_15797,N_16315);
nor U20855 (N_20855,N_15595,N_15676);
nor U20856 (N_20856,N_16276,N_17630);
or U20857 (N_20857,N_17742,N_17690);
nor U20858 (N_20858,N_15798,N_16168);
and U20859 (N_20859,N_15905,N_17046);
nor U20860 (N_20860,N_16157,N_16828);
nor U20861 (N_20861,N_17191,N_15322);
and U20862 (N_20862,N_17935,N_17372);
nor U20863 (N_20863,N_16024,N_17366);
nor U20864 (N_20864,N_15068,N_15851);
or U20865 (N_20865,N_17155,N_17620);
and U20866 (N_20866,N_15446,N_17819);
nor U20867 (N_20867,N_16988,N_17662);
xor U20868 (N_20868,N_17040,N_17532);
nand U20869 (N_20869,N_16193,N_15700);
and U20870 (N_20870,N_17018,N_15711);
or U20871 (N_20871,N_17714,N_17736);
nand U20872 (N_20872,N_15778,N_15591);
nor U20873 (N_20873,N_16922,N_16329);
nor U20874 (N_20874,N_15304,N_16205);
or U20875 (N_20875,N_15225,N_17979);
nor U20876 (N_20876,N_15986,N_15150);
or U20877 (N_20877,N_17793,N_17648);
xnor U20878 (N_20878,N_17059,N_16123);
or U20879 (N_20879,N_16533,N_15113);
and U20880 (N_20880,N_16402,N_16805);
nor U20881 (N_20881,N_16572,N_15606);
or U20882 (N_20882,N_15862,N_16606);
nand U20883 (N_20883,N_15364,N_15413);
or U20884 (N_20884,N_16057,N_15068);
or U20885 (N_20885,N_16174,N_15348);
or U20886 (N_20886,N_17904,N_17880);
nor U20887 (N_20887,N_17152,N_17884);
or U20888 (N_20888,N_16376,N_15314);
nor U20889 (N_20889,N_15344,N_17124);
nor U20890 (N_20890,N_16926,N_17355);
nor U20891 (N_20891,N_17170,N_17246);
nor U20892 (N_20892,N_17608,N_17592);
and U20893 (N_20893,N_16962,N_17448);
and U20894 (N_20894,N_16421,N_15083);
or U20895 (N_20895,N_15073,N_17288);
xor U20896 (N_20896,N_16841,N_15797);
nand U20897 (N_20897,N_15999,N_15827);
and U20898 (N_20898,N_17184,N_15179);
nand U20899 (N_20899,N_17454,N_16225);
and U20900 (N_20900,N_17527,N_16248);
nor U20901 (N_20901,N_15413,N_16382);
xor U20902 (N_20902,N_15471,N_17189);
nor U20903 (N_20903,N_15432,N_17122);
or U20904 (N_20904,N_16746,N_16315);
and U20905 (N_20905,N_16249,N_16341);
nor U20906 (N_20906,N_16055,N_17234);
and U20907 (N_20907,N_15043,N_16270);
or U20908 (N_20908,N_15431,N_17062);
and U20909 (N_20909,N_17705,N_15179);
nor U20910 (N_20910,N_17749,N_16434);
and U20911 (N_20911,N_16378,N_15266);
nor U20912 (N_20912,N_16078,N_17719);
nand U20913 (N_20913,N_15965,N_16287);
nand U20914 (N_20914,N_16867,N_15801);
nor U20915 (N_20915,N_17930,N_16606);
nand U20916 (N_20916,N_15475,N_17598);
nand U20917 (N_20917,N_15953,N_16249);
and U20918 (N_20918,N_16534,N_17215);
nand U20919 (N_20919,N_16117,N_15339);
and U20920 (N_20920,N_17134,N_16046);
or U20921 (N_20921,N_15482,N_15554);
or U20922 (N_20922,N_15956,N_15337);
nand U20923 (N_20923,N_17478,N_16993);
nand U20924 (N_20924,N_17542,N_16152);
nor U20925 (N_20925,N_16734,N_17017);
nand U20926 (N_20926,N_17810,N_17733);
or U20927 (N_20927,N_15113,N_17418);
nor U20928 (N_20928,N_15007,N_17344);
nor U20929 (N_20929,N_15340,N_15284);
nand U20930 (N_20930,N_15013,N_15845);
and U20931 (N_20931,N_16336,N_15145);
and U20932 (N_20932,N_16961,N_15684);
nor U20933 (N_20933,N_16546,N_15884);
or U20934 (N_20934,N_17322,N_16970);
xor U20935 (N_20935,N_16630,N_16993);
and U20936 (N_20936,N_16098,N_15818);
and U20937 (N_20937,N_17174,N_15598);
and U20938 (N_20938,N_15609,N_15031);
and U20939 (N_20939,N_16616,N_16583);
nand U20940 (N_20940,N_15310,N_17450);
and U20941 (N_20941,N_15840,N_15350);
nand U20942 (N_20942,N_15670,N_17512);
and U20943 (N_20943,N_17268,N_16572);
nor U20944 (N_20944,N_17457,N_17815);
or U20945 (N_20945,N_15002,N_17362);
and U20946 (N_20946,N_17919,N_15409);
nor U20947 (N_20947,N_15083,N_15443);
xnor U20948 (N_20948,N_16197,N_15113);
nor U20949 (N_20949,N_15070,N_17510);
and U20950 (N_20950,N_16586,N_15902);
or U20951 (N_20951,N_15459,N_17667);
xor U20952 (N_20952,N_17148,N_17829);
and U20953 (N_20953,N_16555,N_15958);
nor U20954 (N_20954,N_15367,N_16245);
or U20955 (N_20955,N_16112,N_15494);
xnor U20956 (N_20956,N_15668,N_15832);
nand U20957 (N_20957,N_17124,N_17615);
nand U20958 (N_20958,N_17958,N_15246);
and U20959 (N_20959,N_17940,N_17715);
xnor U20960 (N_20960,N_15005,N_17833);
xnor U20961 (N_20961,N_15502,N_16296);
xnor U20962 (N_20962,N_16070,N_16255);
nand U20963 (N_20963,N_17687,N_17056);
nor U20964 (N_20964,N_15862,N_17830);
and U20965 (N_20965,N_17530,N_15214);
or U20966 (N_20966,N_16397,N_15577);
nor U20967 (N_20967,N_16751,N_17419);
nand U20968 (N_20968,N_15280,N_17523);
nor U20969 (N_20969,N_15934,N_17382);
and U20970 (N_20970,N_15700,N_15438);
nand U20971 (N_20971,N_16291,N_16284);
or U20972 (N_20972,N_15303,N_17747);
xnor U20973 (N_20973,N_15104,N_15827);
or U20974 (N_20974,N_16582,N_17555);
or U20975 (N_20975,N_17504,N_16919);
nor U20976 (N_20976,N_16924,N_17592);
and U20977 (N_20977,N_15369,N_16298);
xor U20978 (N_20978,N_16671,N_16770);
or U20979 (N_20979,N_16730,N_16288);
nor U20980 (N_20980,N_17337,N_17833);
and U20981 (N_20981,N_15246,N_17110);
or U20982 (N_20982,N_16652,N_15539);
nor U20983 (N_20983,N_15069,N_15496);
nor U20984 (N_20984,N_15773,N_16063);
nand U20985 (N_20985,N_15884,N_15510);
nor U20986 (N_20986,N_16669,N_15925);
nor U20987 (N_20987,N_15835,N_15663);
nand U20988 (N_20988,N_15992,N_15149);
xnor U20989 (N_20989,N_15817,N_16126);
nor U20990 (N_20990,N_16337,N_16379);
or U20991 (N_20991,N_16268,N_17147);
nor U20992 (N_20992,N_15193,N_16519);
xor U20993 (N_20993,N_17944,N_17479);
and U20994 (N_20994,N_15501,N_17656);
nand U20995 (N_20995,N_17317,N_17682);
nand U20996 (N_20996,N_15193,N_15573);
nand U20997 (N_20997,N_17285,N_17514);
and U20998 (N_20998,N_17839,N_15600);
nor U20999 (N_20999,N_15168,N_16284);
and U21000 (N_21000,N_18382,N_19295);
or U21001 (N_21001,N_20436,N_19056);
nand U21002 (N_21002,N_19106,N_19840);
or U21003 (N_21003,N_19336,N_20309);
or U21004 (N_21004,N_20983,N_20329);
and U21005 (N_21005,N_19745,N_19967);
and U21006 (N_21006,N_20172,N_18396);
nor U21007 (N_21007,N_20252,N_19079);
nand U21008 (N_21008,N_20775,N_19096);
and U21009 (N_21009,N_20072,N_20641);
nand U21010 (N_21010,N_19319,N_19981);
nor U21011 (N_21011,N_18459,N_19726);
xnor U21012 (N_21012,N_19899,N_18939);
and U21013 (N_21013,N_19758,N_20743);
or U21014 (N_21014,N_18812,N_20842);
or U21015 (N_21015,N_19493,N_19135);
nand U21016 (N_21016,N_20690,N_19437);
nand U21017 (N_21017,N_19152,N_20941);
nand U21018 (N_21018,N_18371,N_20210);
or U21019 (N_21019,N_18690,N_19577);
xnor U21020 (N_21020,N_19980,N_18881);
nor U21021 (N_21021,N_18608,N_20532);
nor U21022 (N_21022,N_20076,N_18346);
nor U21023 (N_21023,N_20556,N_19140);
nand U21024 (N_21024,N_18452,N_19146);
and U21025 (N_21025,N_20707,N_18302);
nand U21026 (N_21026,N_18402,N_18518);
or U21027 (N_21027,N_18101,N_19894);
xor U21028 (N_21028,N_18900,N_18029);
or U21029 (N_21029,N_19795,N_18246);
or U21030 (N_21030,N_20365,N_20134);
and U21031 (N_21031,N_20129,N_19272);
nand U21032 (N_21032,N_18805,N_20531);
nand U21033 (N_21033,N_19053,N_19728);
or U21034 (N_21034,N_19603,N_18128);
nor U21035 (N_21035,N_18352,N_20725);
or U21036 (N_21036,N_19667,N_18222);
nor U21037 (N_21037,N_18619,N_20428);
nand U21038 (N_21038,N_18543,N_18033);
nand U21039 (N_21039,N_18449,N_18969);
nand U21040 (N_21040,N_18430,N_19507);
nor U21041 (N_21041,N_18625,N_19622);
or U21042 (N_21042,N_19123,N_18853);
nand U21043 (N_21043,N_18023,N_19306);
xnor U21044 (N_21044,N_20798,N_18290);
nand U21045 (N_21045,N_18549,N_19904);
and U21046 (N_21046,N_20986,N_20332);
nor U21047 (N_21047,N_19033,N_19486);
nor U21048 (N_21048,N_18976,N_19928);
xor U21049 (N_21049,N_18924,N_19343);
and U21050 (N_21050,N_19551,N_19270);
or U21051 (N_21051,N_18068,N_19235);
nand U21052 (N_21052,N_18126,N_20821);
or U21053 (N_21053,N_18523,N_19464);
nand U21054 (N_21054,N_18506,N_19470);
and U21055 (N_21055,N_19640,N_20173);
nor U21056 (N_21056,N_20489,N_18330);
and U21057 (N_21057,N_20876,N_20561);
and U21058 (N_21058,N_18666,N_19202);
xnor U21059 (N_21059,N_20978,N_19003);
nor U21060 (N_21060,N_20931,N_18771);
nand U21061 (N_21061,N_20139,N_19528);
and U21062 (N_21062,N_20853,N_20406);
nor U21063 (N_21063,N_19584,N_20482);
or U21064 (N_21064,N_20936,N_18561);
nor U21065 (N_21065,N_20075,N_19711);
or U21066 (N_21066,N_19410,N_18059);
or U21067 (N_21067,N_19816,N_19345);
nand U21068 (N_21068,N_20011,N_20766);
nor U21069 (N_21069,N_18836,N_18591);
and U21070 (N_21070,N_18806,N_19426);
and U21071 (N_21071,N_19991,N_19597);
or U21072 (N_21072,N_18992,N_20396);
or U21073 (N_21073,N_19301,N_20148);
and U21074 (N_21074,N_18753,N_18626);
or U21075 (N_21075,N_19349,N_19596);
or U21076 (N_21076,N_19124,N_18337);
and U21077 (N_21077,N_18929,N_19230);
or U21078 (N_21078,N_18675,N_20687);
nand U21079 (N_21079,N_20717,N_18892);
nand U21080 (N_21080,N_19269,N_19378);
and U21081 (N_21081,N_20156,N_18709);
nand U21082 (N_21082,N_19309,N_20926);
and U21083 (N_21083,N_18269,N_18750);
nand U21084 (N_21084,N_19685,N_20238);
or U21085 (N_21085,N_18254,N_18963);
nor U21086 (N_21086,N_19273,N_19327);
or U21087 (N_21087,N_19141,N_20657);
nand U21088 (N_21088,N_20003,N_19875);
xor U21089 (N_21089,N_20473,N_18032);
and U21090 (N_21090,N_19495,N_19340);
nor U21091 (N_21091,N_18846,N_19794);
nor U21092 (N_21092,N_19290,N_19885);
and U21093 (N_21093,N_19595,N_20426);
and U21094 (N_21094,N_19455,N_20455);
nand U21095 (N_21095,N_18581,N_20814);
nor U21096 (N_21096,N_20940,N_18741);
or U21097 (N_21097,N_20783,N_20987);
nand U21098 (N_21098,N_20680,N_19258);
or U21099 (N_21099,N_20155,N_18738);
xnor U21100 (N_21100,N_19449,N_20086);
nand U21101 (N_21101,N_20189,N_20184);
nand U21102 (N_21102,N_18163,N_18260);
and U21103 (N_21103,N_19751,N_20419);
and U21104 (N_21104,N_18184,N_19600);
or U21105 (N_21105,N_19709,N_18973);
nand U21106 (N_21106,N_20614,N_18258);
nor U21107 (N_21107,N_19281,N_19617);
and U21108 (N_21108,N_18011,N_19203);
nor U21109 (N_21109,N_19854,N_19147);
xor U21110 (N_21110,N_20738,N_20168);
xnor U21111 (N_21111,N_20515,N_18948);
nor U21112 (N_21112,N_18162,N_18340);
xor U21113 (N_21113,N_19847,N_20327);
nand U21114 (N_21114,N_18880,N_20079);
or U21115 (N_21115,N_19534,N_20703);
nand U21116 (N_21116,N_20899,N_19761);
and U21117 (N_21117,N_20035,N_20626);
or U21118 (N_21118,N_18253,N_19246);
nand U21119 (N_21119,N_18996,N_20767);
nand U21120 (N_21120,N_20729,N_20277);
nand U21121 (N_21121,N_19939,N_20866);
or U21122 (N_21122,N_19965,N_19490);
or U21123 (N_21123,N_19253,N_18610);
nand U21124 (N_21124,N_19628,N_19353);
nand U21125 (N_21125,N_18531,N_18102);
and U21126 (N_21126,N_19564,N_20742);
nor U21127 (N_21127,N_19805,N_19484);
nor U21128 (N_21128,N_18325,N_18431);
nor U21129 (N_21129,N_19744,N_19477);
or U21130 (N_21130,N_19959,N_19282);
and U21131 (N_21131,N_19362,N_19589);
xnor U21132 (N_21132,N_20207,N_19641);
xor U21133 (N_21133,N_19606,N_18151);
xor U21134 (N_21134,N_19245,N_18870);
and U21135 (N_21135,N_18063,N_19837);
nor U21136 (N_21136,N_18949,N_18400);
or U21137 (N_21137,N_18558,N_18796);
nor U21138 (N_21138,N_20163,N_18329);
or U21139 (N_21139,N_19896,N_18886);
and U21140 (N_21140,N_18021,N_19408);
or U21141 (N_21141,N_18009,N_18694);
nand U21142 (N_21142,N_19749,N_20991);
nor U21143 (N_21143,N_18208,N_18377);
nand U21144 (N_21144,N_18732,N_20666);
nor U21145 (N_21145,N_19307,N_18131);
and U21146 (N_21146,N_20678,N_18974);
or U21147 (N_21147,N_20143,N_18994);
xnor U21148 (N_21148,N_19344,N_20387);
nand U21149 (N_21149,N_18448,N_19673);
or U21150 (N_21150,N_20824,N_20340);
or U21151 (N_21151,N_19357,N_18108);
nor U21152 (N_21152,N_19873,N_20362);
xnor U21153 (N_21153,N_19262,N_18091);
and U21154 (N_21154,N_20985,N_19839);
or U21155 (N_21155,N_18483,N_18294);
or U21156 (N_21156,N_18706,N_18327);
nor U21157 (N_21157,N_19738,N_18259);
xnor U21158 (N_21158,N_19347,N_20637);
and U21159 (N_21159,N_20648,N_18687);
nand U21160 (N_21160,N_18217,N_20115);
or U21161 (N_21161,N_20398,N_20120);
and U21162 (N_21162,N_18354,N_18562);
nor U21163 (N_21163,N_20583,N_18257);
xnor U21164 (N_21164,N_18262,N_20967);
or U21165 (N_21165,N_20881,N_19650);
nand U21166 (N_21166,N_18692,N_19583);
and U21167 (N_21167,N_19724,N_20417);
nor U21168 (N_21168,N_19655,N_20551);
and U21169 (N_21169,N_19030,N_18708);
nor U21170 (N_21170,N_18792,N_20322);
nand U21171 (N_21171,N_18095,N_18857);
nor U21172 (N_21172,N_20476,N_19718);
and U21173 (N_21173,N_20787,N_20060);
nand U21174 (N_21174,N_18946,N_19260);
nor U21175 (N_21175,N_18953,N_18803);
or U21176 (N_21176,N_18952,N_20534);
nand U21177 (N_21177,N_18555,N_19624);
or U21178 (N_21178,N_19500,N_20921);
nand U21179 (N_21179,N_19571,N_18175);
and U21180 (N_21180,N_20144,N_20696);
nand U21181 (N_21181,N_18736,N_18422);
nor U21182 (N_21182,N_19924,N_20355);
and U21183 (N_21183,N_19883,N_19292);
or U21184 (N_21184,N_19429,N_19304);
nor U21185 (N_21185,N_20470,N_19774);
and U21186 (N_21186,N_18441,N_19215);
xnor U21187 (N_21187,N_20465,N_19494);
or U21188 (N_21188,N_18264,N_19457);
and U21189 (N_21189,N_20167,N_20984);
nand U21190 (N_21190,N_18829,N_18757);
nor U21191 (N_21191,N_18985,N_18092);
and U21192 (N_21192,N_18006,N_18094);
nor U21193 (N_21193,N_18243,N_19663);
nor U21194 (N_21194,N_20747,N_19513);
nor U21195 (N_21195,N_19782,N_20286);
nor U21196 (N_21196,N_20023,N_18931);
nor U21197 (N_21197,N_18800,N_20585);
nor U21198 (N_21198,N_18845,N_18837);
or U21199 (N_21199,N_20835,N_18779);
or U21200 (N_21200,N_20812,N_19586);
xnor U21201 (N_21201,N_19293,N_19403);
nor U21202 (N_21202,N_20067,N_20834);
or U21203 (N_21203,N_19083,N_19958);
and U21204 (N_21204,N_18461,N_19392);
and U21205 (N_21205,N_18417,N_18535);
xnor U21206 (N_21206,N_19069,N_20545);
and U21207 (N_21207,N_19374,N_19601);
or U21208 (N_21208,N_19447,N_20508);
and U21209 (N_21209,N_18471,N_20728);
or U21210 (N_21210,N_18825,N_20395);
and U21211 (N_21211,N_20536,N_19112);
nand U21212 (N_21212,N_18312,N_18274);
or U21213 (N_21213,N_18442,N_19328);
and U21214 (N_21214,N_19972,N_18936);
nor U21215 (N_21215,N_19004,N_19983);
xor U21216 (N_21216,N_18576,N_18170);
nor U21217 (N_21217,N_20377,N_19912);
xnor U21218 (N_21218,N_19120,N_20682);
nand U21219 (N_21219,N_18744,N_18678);
or U21220 (N_21220,N_20212,N_20069);
nor U21221 (N_21221,N_19961,N_18760);
nor U21222 (N_21222,N_20042,N_19330);
xor U21223 (N_21223,N_19434,N_18632);
and U21224 (N_21224,N_20056,N_18901);
or U21225 (N_21225,N_20304,N_19370);
or U21226 (N_21226,N_19799,N_19969);
nand U21227 (N_21227,N_18194,N_19405);
nor U21228 (N_21228,N_19868,N_20381);
and U21229 (N_21229,N_19436,N_18199);
or U21230 (N_21230,N_18154,N_19395);
or U21231 (N_21231,N_18315,N_19066);
or U21232 (N_21232,N_19974,N_19504);
and U21233 (N_21233,N_20851,N_18293);
xor U21234 (N_21234,N_19103,N_19765);
nand U21235 (N_21235,N_19017,N_19629);
nor U21236 (N_21236,N_20723,N_19067);
or U21237 (N_21237,N_20865,N_18823);
and U21238 (N_21238,N_18276,N_20468);
or U21239 (N_21239,N_20226,N_18201);
or U21240 (N_21240,N_20629,N_20861);
and U21241 (N_21241,N_20801,N_20625);
nand U21242 (N_21242,N_18482,N_18215);
nor U21243 (N_21243,N_20907,N_19978);
nor U21244 (N_21244,N_18305,N_18532);
or U21245 (N_21245,N_20839,N_19278);
nand U21246 (N_21246,N_18727,N_18462);
xor U21247 (N_21247,N_18964,N_18956);
and U21248 (N_21248,N_19942,N_19148);
nor U21249 (N_21249,N_19248,N_19680);
nor U21250 (N_21250,N_19028,N_18841);
and U21251 (N_21251,N_19737,N_19212);
and U21252 (N_21252,N_18255,N_20638);
nor U21253 (N_21253,N_20669,N_19948);
or U21254 (N_21254,N_19401,N_18070);
nor U21255 (N_21255,N_20177,N_18832);
and U21256 (N_21256,N_20361,N_19393);
and U21257 (N_21257,N_20517,N_18500);
and U21258 (N_21258,N_20720,N_20898);
nor U21259 (N_21259,N_20333,N_19802);
nand U21260 (N_21260,N_19946,N_18489);
nand U21261 (N_21261,N_18782,N_20374);
and U21262 (N_21262,N_19042,N_18238);
or U21263 (N_21263,N_19296,N_20371);
nor U21264 (N_21264,N_18465,N_20160);
or U21265 (N_21265,N_19492,N_19989);
and U21266 (N_21266,N_19804,N_19377);
nand U21267 (N_21267,N_19741,N_20591);
nand U21268 (N_21268,N_19386,N_20855);
or U21269 (N_21269,N_18527,N_18013);
and U21270 (N_21270,N_18115,N_20415);
nor U21271 (N_21271,N_20380,N_20486);
nand U21272 (N_21272,N_19529,N_18177);
and U21273 (N_21273,N_19676,N_19322);
nor U21274 (N_21274,N_19545,N_20518);
nor U21275 (N_21275,N_20873,N_20947);
and U21276 (N_21276,N_20151,N_20871);
xor U21277 (N_21277,N_19478,N_19381);
nor U21278 (N_21278,N_19136,N_19199);
nand U21279 (N_21279,N_18181,N_18844);
nor U21280 (N_21280,N_19118,N_18096);
or U21281 (N_21281,N_18767,N_20231);
or U21282 (N_21282,N_19329,N_18848);
or U21283 (N_21283,N_19018,N_20126);
or U21284 (N_21284,N_20099,N_18428);
or U21285 (N_21285,N_18456,N_18401);
or U21286 (N_21286,N_19530,N_19591);
nand U21287 (N_21287,N_19797,N_18838);
and U21288 (N_21288,N_18569,N_19735);
nor U21289 (N_21289,N_18959,N_20593);
or U21290 (N_21290,N_18460,N_18999);
xor U21291 (N_21291,N_19976,N_19001);
nand U21292 (N_21292,N_20150,N_18686);
and U21293 (N_21293,N_19131,N_18475);
nor U21294 (N_21294,N_18394,N_20499);
and U21295 (N_21295,N_19697,N_19732);
nor U21296 (N_21296,N_20968,N_18391);
and U21297 (N_21297,N_18157,N_19111);
nand U21298 (N_21298,N_19178,N_20457);
or U21299 (N_21299,N_20636,N_19602);
nand U21300 (N_21300,N_20521,N_19389);
and U21301 (N_21301,N_20062,N_20647);
and U21302 (N_21302,N_20575,N_20430);
nor U21303 (N_21303,N_19369,N_19055);
nor U21304 (N_21304,N_19009,N_20284);
or U21305 (N_21305,N_18214,N_19119);
and U21306 (N_21306,N_20495,N_19649);
nand U21307 (N_21307,N_18719,N_18652);
and U21308 (N_21308,N_18883,N_18918);
xor U21309 (N_21309,N_19787,N_20002);
nor U21310 (N_21310,N_18122,N_19396);
nand U21311 (N_21311,N_20171,N_19716);
or U21312 (N_21312,N_19932,N_18634);
or U21313 (N_21313,N_18057,N_20410);
nor U21314 (N_21314,N_19021,N_18689);
and U21315 (N_21315,N_18539,N_20832);
nor U21316 (N_21316,N_19471,N_20217);
nor U21317 (N_21317,N_20911,N_20253);
nor U21318 (N_21318,N_18542,N_18876);
and U21319 (N_21319,N_18144,N_20559);
nand U21320 (N_21320,N_18896,N_20019);
xor U21321 (N_21321,N_20127,N_19472);
nand U21322 (N_21322,N_20758,N_19714);
nand U21323 (N_21323,N_19320,N_20892);
nor U21324 (N_21324,N_19700,N_19285);
nand U21325 (N_21325,N_19354,N_20093);
nand U21326 (N_21326,N_19998,N_20951);
nor U21327 (N_21327,N_20768,N_20979);
nor U21328 (N_21328,N_18715,N_19954);
or U21329 (N_21329,N_20000,N_18587);
nand U21330 (N_21330,N_19913,N_19300);
nor U21331 (N_21331,N_20234,N_20193);
and U21332 (N_21332,N_19257,N_18839);
and U21333 (N_21333,N_20826,N_20825);
xnor U21334 (N_21334,N_18646,N_20346);
nand U21335 (N_21335,N_20675,N_19893);
and U21336 (N_21336,N_18613,N_20731);
nand U21337 (N_21337,N_19962,N_18373);
nor U21338 (N_21338,N_18830,N_20100);
or U21339 (N_21339,N_18510,N_19771);
and U21340 (N_21340,N_20740,N_18849);
and U21341 (N_21341,N_20845,N_20563);
nand U21342 (N_21342,N_19171,N_19866);
nand U21343 (N_21343,N_19621,N_20528);
nand U21344 (N_21344,N_20670,N_19944);
nand U21345 (N_21345,N_20256,N_19139);
or U21346 (N_21346,N_18917,N_19590);
nor U21347 (N_21347,N_20524,N_18043);
and U21348 (N_21348,N_19678,N_18357);
or U21349 (N_21349,N_19214,N_18130);
or U21350 (N_21350,N_18004,N_20822);
nor U21351 (N_21351,N_18798,N_18065);
xor U21352 (N_21352,N_20818,N_18724);
and U21353 (N_21353,N_19323,N_19815);
or U21354 (N_21354,N_20512,N_20982);
or U21355 (N_21355,N_20401,N_18287);
xor U21356 (N_21356,N_20481,N_20992);
nand U21357 (N_21357,N_20359,N_18421);
nand U21358 (N_21358,N_18336,N_19722);
xnor U21359 (N_21359,N_20664,N_18622);
nand U21360 (N_21360,N_19071,N_18178);
or U21361 (N_21361,N_20658,N_20450);
nor U21362 (N_21362,N_18477,N_18685);
nand U21363 (N_21363,N_19427,N_19996);
nand U21364 (N_21364,N_20527,N_19853);
and U21365 (N_21365,N_18790,N_18047);
and U21366 (N_21366,N_18867,N_19878);
nand U21367 (N_21367,N_18758,N_18618);
and U21368 (N_21368,N_20706,N_19216);
nor U21369 (N_21369,N_19747,N_20045);
nor U21370 (N_21370,N_18306,N_20581);
and U21371 (N_21371,N_19388,N_18875);
nand U21372 (N_21372,N_18654,N_19243);
nor U21373 (N_21373,N_20015,N_19731);
xor U21374 (N_21374,N_20026,N_18761);
and U21375 (N_21375,N_19196,N_20878);
nor U21376 (N_21376,N_19190,N_20420);
nor U21377 (N_21377,N_19635,N_18291);
nand U21378 (N_21378,N_18814,N_20884);
nand U21379 (N_21379,N_19713,N_20860);
nor U21380 (N_21380,N_19646,N_18676);
nand U21381 (N_21381,N_20954,N_18042);
nor U21382 (N_21382,N_19011,N_20055);
and U21383 (N_21383,N_19218,N_18544);
and U21384 (N_21384,N_19918,N_20973);
nor U21385 (N_21385,N_20004,N_20616);
or U21386 (N_21386,N_19525,N_20070);
nor U21387 (N_21387,N_19770,N_18801);
or U21388 (N_21388,N_18797,N_18932);
nand U21389 (N_21389,N_19776,N_19811);
nand U21390 (N_21390,N_19515,N_18025);
or U21391 (N_21391,N_19609,N_19085);
or U21392 (N_21392,N_20196,N_18112);
or U21393 (N_21393,N_18049,N_20145);
nor U21394 (N_21394,N_18568,N_19582);
nand U21395 (N_21395,N_19952,N_20789);
and U21396 (N_21396,N_18769,N_18145);
xor U21397 (N_21397,N_20872,N_18987);
and U21398 (N_21398,N_20570,N_18602);
nor U21399 (N_21399,N_18223,N_19647);
and U21400 (N_21400,N_19445,N_20033);
nand U21401 (N_21401,N_18376,N_20667);
nand U21402 (N_21402,N_18388,N_20584);
nor U21403 (N_21403,N_18642,N_18479);
nor U21404 (N_21404,N_19409,N_19791);
nand U21405 (N_21405,N_19435,N_19173);
nor U21406 (N_21406,N_20312,N_19608);
and U21407 (N_21407,N_20988,N_20057);
or U21408 (N_21408,N_19326,N_20749);
and U21409 (N_21409,N_20507,N_19242);
xnor U21410 (N_21410,N_19933,N_19817);
or U21411 (N_21411,N_18756,N_18713);
or U21412 (N_21412,N_20452,N_19143);
and U21413 (N_21413,N_20710,N_20413);
and U21414 (N_21414,N_18893,N_20888);
nor U21415 (N_21415,N_20170,N_20848);
xnor U21416 (N_21416,N_20552,N_18051);
xor U21417 (N_21417,N_18055,N_20542);
nor U21418 (N_21418,N_18473,N_18824);
nand U21419 (N_21419,N_18366,N_19546);
nand U21420 (N_21420,N_19479,N_19007);
and U21421 (N_21421,N_18906,N_18316);
nand U21422 (N_21422,N_19180,N_20554);
and U21423 (N_21423,N_20034,N_18504);
and U21424 (N_21424,N_18795,N_20761);
nor U21425 (N_21425,N_18370,N_20192);
nor U21426 (N_21426,N_20314,N_19054);
and U21427 (N_21427,N_18908,N_18943);
and U21428 (N_21428,N_19047,N_20128);
nand U21429 (N_21429,N_18450,N_19929);
and U21430 (N_21430,N_18139,N_20378);
or U21431 (N_21431,N_18445,N_18574);
and U21432 (N_21432,N_20830,N_18491);
and U21433 (N_21433,N_20005,N_18429);
nor U21434 (N_21434,N_20777,N_19497);
and U21435 (N_21435,N_19556,N_19454);
nand U21436 (N_21436,N_18989,N_20258);
and U21437 (N_21437,N_19938,N_19879);
and U21438 (N_21438,N_18755,N_18530);
nand U21439 (N_21439,N_19580,N_20772);
nor U21440 (N_21440,N_18044,N_20024);
and U21441 (N_21441,N_19049,N_20477);
xor U21442 (N_21442,N_18559,N_19955);
nand U21443 (N_21443,N_20358,N_18747);
xor U21444 (N_21444,N_18285,N_18409);
and U21445 (N_21445,N_18603,N_19852);
nand U21446 (N_21446,N_18146,N_19174);
nor U21447 (N_21447,N_19578,N_19544);
and U21448 (N_21448,N_19828,N_19516);
and U21449 (N_21449,N_19982,N_18640);
and U21450 (N_21450,N_20750,N_18171);
or U21451 (N_21451,N_20923,N_19366);
nand U21452 (N_21452,N_20118,N_20633);
nor U21453 (N_21453,N_18458,N_19145);
and U21454 (N_21454,N_20997,N_20108);
nand U21455 (N_21455,N_19964,N_20449);
and U21456 (N_21456,N_19756,N_19268);
nand U21457 (N_21457,N_18638,N_18239);
or U21458 (N_21458,N_19211,N_19267);
and U21459 (N_21459,N_18089,N_20964);
nand U21460 (N_21460,N_19587,N_19460);
nor U21461 (N_21461,N_18564,N_19082);
nand U21462 (N_21462,N_20714,N_18677);
and U21463 (N_21463,N_18451,N_19537);
nand U21464 (N_21464,N_19754,N_20367);
and U21465 (N_21465,N_20928,N_20908);
and U21466 (N_21466,N_20604,N_18586);
nor U21467 (N_21467,N_20813,N_20513);
nand U21468 (N_21468,N_19917,N_20891);
nor U21469 (N_21469,N_20573,N_19517);
and U21470 (N_21470,N_20245,N_19090);
and U21471 (N_21471,N_19360,N_18863);
and U21472 (N_21472,N_18804,N_19630);
nor U21473 (N_21473,N_18833,N_20886);
nand U21474 (N_21474,N_18362,N_20922);
or U21475 (N_21475,N_18879,N_20297);
or U21476 (N_21476,N_20819,N_20390);
nor U21477 (N_21477,N_18350,N_20976);
nand U21478 (N_21478,N_20858,N_18842);
xor U21479 (N_21479,N_19559,N_19683);
and U21480 (N_21480,N_18873,N_18311);
nand U21481 (N_21481,N_19681,N_20175);
or U21482 (N_21482,N_19213,N_20338);
xor U21483 (N_21483,N_19598,N_19999);
nor U21484 (N_21484,N_20001,N_19541);
or U21485 (N_21485,N_18161,N_19176);
and U21486 (N_21486,N_20577,N_20257);
and U21487 (N_21487,N_20356,N_18907);
and U21488 (N_21488,N_18134,N_20971);
and U21489 (N_21489,N_20123,N_19153);
or U21490 (N_21490,N_18501,N_18748);
or U21491 (N_21491,N_18960,N_18598);
and U21492 (N_21492,N_19480,N_20538);
xnor U21493 (N_21493,N_20927,N_18765);
and U21494 (N_21494,N_19674,N_18817);
nand U21495 (N_21495,N_20588,N_18572);
nand U21496 (N_21496,N_18016,N_20915);
or U21497 (N_21497,N_18874,N_18275);
xnor U21498 (N_21498,N_19032,N_20278);
or U21499 (N_21499,N_18653,N_19702);
nand U21500 (N_21500,N_20236,N_19666);
and U21501 (N_21501,N_18843,N_19125);
or U21502 (N_21502,N_19276,N_18183);
nor U21503 (N_21503,N_20601,N_20533);
or U21504 (N_21504,N_20628,N_19834);
nor U21505 (N_21505,N_19593,N_19192);
nand U21506 (N_21506,N_20182,N_18540);
nand U21507 (N_21507,N_19704,N_19499);
nor U21508 (N_21508,N_20909,N_18811);
or U21509 (N_21509,N_20662,N_18176);
and U21510 (N_21510,N_19299,N_20400);
nand U21511 (N_21511,N_19692,N_19155);
nor U21512 (N_21512,N_18639,N_20882);
nor U21513 (N_21513,N_20646,N_18623);
nand U21514 (N_21514,N_18359,N_20681);
xnor U21515 (N_21515,N_18298,N_18935);
xnor U21516 (N_21516,N_19458,N_19807);
nor U21517 (N_21517,N_20315,N_18237);
or U21518 (N_21518,N_20068,N_20956);
nor U21519 (N_21519,N_19669,N_18152);
nand U21520 (N_21520,N_19019,N_18123);
xor U21521 (N_21521,N_19059,N_18854);
xnor U21522 (N_21522,N_18067,N_18488);
nand U21523 (N_21523,N_19158,N_18364);
nor U21524 (N_21524,N_19391,N_19519);
nand U21525 (N_21525,N_19755,N_18365);
nor U21526 (N_21526,N_20305,N_20544);
nand U21527 (N_21527,N_18615,N_18045);
nor U21528 (N_21528,N_18594,N_18981);
and U21529 (N_21529,N_18135,N_19129);
nor U21530 (N_21530,N_20530,N_20924);
or U21531 (N_21531,N_19832,N_20014);
and U21532 (N_21532,N_18075,N_18344);
and U21533 (N_21533,N_20339,N_20247);
nor U21534 (N_21534,N_18397,N_20043);
and U21535 (N_21535,N_19303,N_20649);
nor U21536 (N_21536,N_19289,N_19407);
and U21537 (N_21537,N_18072,N_19316);
nor U21538 (N_21538,N_19956,N_18210);
nor U21539 (N_21539,N_18381,N_18551);
and U21540 (N_21540,N_18813,N_20856);
nand U21541 (N_21541,N_18313,N_20602);
and U21542 (N_21542,N_20183,N_18984);
nor U21543 (N_21543,N_20291,N_20894);
or U21544 (N_21544,N_18148,N_18138);
or U21545 (N_21545,N_19126,N_19696);
and U21546 (N_21546,N_18000,N_18179);
nand U21547 (N_21547,N_19318,N_19557);
or U21548 (N_21548,N_20125,N_20030);
xnor U21549 (N_21549,N_19931,N_20008);
nor U21550 (N_21550,N_20464,N_19833);
or U21551 (N_21551,N_20509,N_18725);
and U21552 (N_21552,N_18492,N_20500);
and U21553 (N_21553,N_19183,N_20820);
nand U21554 (N_21554,N_18073,N_19725);
and U21555 (N_21555,N_20135,N_18926);
and U21556 (N_21556,N_20065,N_18571);
or U21557 (N_21557,N_19197,N_18665);
nor U21558 (N_21558,N_19233,N_19467);
nand U21559 (N_21559,N_20603,N_20098);
nand U21560 (N_21560,N_20590,N_20440);
and U21561 (N_21561,N_20523,N_20061);
nand U21562 (N_21562,N_18556,N_19489);
xnor U21563 (N_21563,N_19984,N_20849);
and U21564 (N_21564,N_18174,N_19168);
or U21565 (N_21565,N_19073,N_18778);
and U21566 (N_21566,N_20689,N_20439);
or U21567 (N_21567,N_19845,N_18310);
or U21568 (N_21568,N_18256,N_18036);
nor U21569 (N_21569,N_18751,N_20560);
and U21570 (N_21570,N_20555,N_20833);
and U21571 (N_21571,N_18802,N_20009);
or U21572 (N_21572,N_18722,N_20897);
nand U21573 (N_21573,N_19652,N_18395);
xor U21574 (N_21574,N_18425,N_19539);
nor U21575 (N_21575,N_20101,N_20792);
nor U21576 (N_21576,N_18229,N_18991);
nor U21577 (N_21577,N_19540,N_19874);
or U21578 (N_21578,N_19461,N_18386);
xnor U21579 (N_21579,N_20421,N_20427);
nor U21580 (N_21580,N_19599,N_20977);
nor U21581 (N_21581,N_18662,N_20739);
nand U21582 (N_21582,N_19463,N_19166);
or U21583 (N_21583,N_18904,N_18443);
or U21584 (N_21584,N_20576,N_20230);
nor U21585 (N_21585,N_20916,N_18191);
and U21586 (N_21586,N_20393,N_18143);
nand U21587 (N_21587,N_18140,N_18383);
and U21588 (N_21588,N_19757,N_20587);
nand U21589 (N_21589,N_20655,N_19228);
nor U21590 (N_21590,N_19160,N_20963);
or U21591 (N_21591,N_19800,N_20595);
nor U21592 (N_21592,N_20132,N_20350);
nand U21593 (N_21593,N_20096,N_18499);
or U21594 (N_21594,N_18859,N_18216);
or U21595 (N_21595,N_18783,N_18743);
xnor U21596 (N_21596,N_19104,N_20771);
and U21597 (N_21597,N_19312,N_19671);
nand U21598 (N_21598,N_19058,N_18599);
nor U21599 (N_21599,N_18659,N_20970);
nand U21600 (N_21600,N_18137,N_18196);
or U21601 (N_21601,N_18552,N_19365);
xor U21602 (N_21602,N_20698,N_18292);
and U21603 (N_21603,N_19167,N_20569);
nor U21604 (N_21604,N_19132,N_18707);
nor U21605 (N_21605,N_18922,N_20607);
and U21606 (N_21606,N_19000,N_18525);
and U21607 (N_21607,N_20879,N_20321);
or U21608 (N_21608,N_19512,N_19266);
nand U21609 (N_21609,N_19568,N_19572);
nor U21610 (N_21610,N_19223,N_18050);
nand U21611 (N_21611,N_18058,N_20474);
or U21612 (N_21612,N_20402,N_20080);
nand U21613 (N_21613,N_19550,N_19415);
nor U21614 (N_21614,N_19498,N_18641);
or U21615 (N_21615,N_18721,N_20444);
or U21616 (N_21616,N_18084,N_18681);
nand U21617 (N_21617,N_20857,N_19565);
nand U21618 (N_21618,N_19194,N_20535);
or U21619 (N_21619,N_18606,N_18232);
nor U21620 (N_21620,N_20756,N_19821);
nor U21621 (N_21621,N_20282,N_18596);
nand U21622 (N_21622,N_19567,N_19514);
nor U21623 (N_21623,N_19170,N_18090);
nor U21624 (N_21624,N_20046,N_19995);
or U21625 (N_21625,N_18524,N_18774);
and U21626 (N_21626,N_19626,N_18384);
and U21627 (N_21627,N_20716,N_18934);
nand U21628 (N_21628,N_19705,N_19172);
xor U21629 (N_21629,N_18056,N_19502);
nor U21630 (N_21630,N_19960,N_18584);
nor U21631 (N_21631,N_18498,N_19051);
nor U21632 (N_21632,N_20319,N_20582);
or U21633 (N_21633,N_20249,N_18322);
nand U21634 (N_21634,N_20197,N_19997);
and U21635 (N_21635,N_18041,N_20425);
nand U21636 (N_21636,N_20691,N_20594);
or U21637 (N_21637,N_20222,N_18704);
and U21638 (N_21638,N_18248,N_19115);
or U21639 (N_21639,N_20264,N_19936);
nor U21640 (N_21640,N_20142,N_19219);
and U21641 (N_21641,N_18787,N_19739);
or U21642 (N_21642,N_19819,N_18731);
nor U21643 (N_21643,N_19727,N_19050);
nand U21644 (N_21644,N_19902,N_20617);
and U21645 (N_21645,N_19656,N_18745);
nand U21646 (N_21646,N_19075,N_19473);
nand U21647 (N_21647,N_19232,N_19008);
nor U21648 (N_21648,N_20275,N_20945);
nor U21649 (N_21649,N_19835,N_19510);
nor U21650 (N_21650,N_19693,N_18597);
nand U21651 (N_21651,N_19860,N_18655);
nand U21652 (N_21652,N_20935,N_19450);
nor U21653 (N_21653,N_19826,N_18895);
or U21654 (N_21654,N_20867,N_19107);
nor U21655 (N_21655,N_18864,N_18231);
or U21656 (N_21656,N_20730,N_19092);
nand U21657 (N_21657,N_18950,N_20325);
and U21658 (N_21658,N_20955,N_19298);
xnor U21659 (N_21659,N_18111,N_18478);
or U21660 (N_21660,N_19046,N_18822);
nand U21661 (N_21661,N_19308,N_18627);
nor U21662 (N_21662,N_18104,N_19100);
nand U21663 (N_21663,N_20273,N_19616);
nand U21664 (N_21664,N_18988,N_20791);
nor U21665 (N_21665,N_20786,N_19549);
nor U21666 (N_21666,N_20235,N_18005);
nor U21667 (N_21667,N_20082,N_20382);
xor U21668 (N_21668,N_19070,N_20206);
and U21669 (N_21669,N_18034,N_18621);
nand U21670 (N_21670,N_20240,N_18010);
and U21671 (N_21671,N_18752,N_18669);
nand U21672 (N_21672,N_20007,N_20392);
or U21673 (N_21673,N_18204,N_19425);
nand U21674 (N_21674,N_18107,N_18263);
or U21675 (N_21675,N_18351,N_19923);
nor U21676 (N_21676,N_20572,N_20650);
nand U21677 (N_21677,N_19283,N_20456);
xnor U21678 (N_21678,N_19777,N_20423);
nor U21679 (N_21679,N_18710,N_19247);
and U21680 (N_21680,N_19352,N_19768);
or U21681 (N_21681,N_20343,N_19715);
xor U21682 (N_21682,N_19803,N_18119);
and U21683 (N_21683,N_18407,N_20794);
nor U21684 (N_21684,N_18775,N_18297);
and U21685 (N_21685,N_18776,N_20066);
nand U21686 (N_21686,N_20216,N_19193);
or U21687 (N_21687,N_19687,N_19733);
and U21688 (N_21688,N_20962,N_18136);
nor U21689 (N_21689,N_19064,N_20461);
or U21690 (N_21690,N_19341,N_18106);
and U21691 (N_21691,N_20121,N_18320);
and U21692 (N_21692,N_18712,N_19116);
nand U21693 (N_21693,N_18763,N_19610);
nor U21694 (N_21694,N_20021,N_20251);
and U21695 (N_21695,N_18589,N_20353);
nand U21696 (N_21696,N_19506,N_20154);
or U21697 (N_21697,N_19849,N_19639);
and U21698 (N_21698,N_18496,N_19291);
and U21699 (N_21699,N_18242,N_19521);
and U21700 (N_21700,N_18970,N_20492);
or U21701 (N_21701,N_20232,N_20686);
nor U21702 (N_21702,N_18512,N_18087);
nor U21703 (N_21703,N_18508,N_19734);
and U21704 (N_21704,N_18423,N_20422);
or U21705 (N_21705,N_19249,N_19518);
and U21706 (N_21706,N_20215,N_18912);
or U21707 (N_21707,N_20627,N_20178);
nand U21708 (N_21708,N_20162,N_18573);
or U21709 (N_21709,N_18536,N_19846);
xnor U21710 (N_21710,N_19689,N_20980);
xnor U21711 (N_21711,N_19977,N_18052);
and U21712 (N_21712,N_20870,N_20445);
or U21713 (N_21713,N_20567,N_20063);
nand U21714 (N_21714,N_18278,N_19558);
xor U21715 (N_21715,N_19444,N_20213);
nor U21716 (N_21716,N_18167,N_18986);
nand U21717 (N_21717,N_20656,N_18379);
nor U21718 (N_21718,N_20755,N_18563);
nand U21719 (N_21719,N_18700,N_20201);
or U21720 (N_21720,N_18200,N_20780);
nor U21721 (N_21721,N_20209,N_20285);
nor U21722 (N_21722,N_19710,N_19637);
nor U21723 (N_21723,N_20903,N_19036);
and U21724 (N_21724,N_19563,N_19331);
nor U21725 (N_21725,N_19830,N_20272);
or U21726 (N_21726,N_18318,N_20146);
xnor U21727 (N_21727,N_20516,N_19188);
and U21728 (N_21728,N_18645,N_19763);
nand U21729 (N_21729,N_18509,N_19022);
or U21730 (N_21730,N_20869,N_20225);
nand U21731 (N_21731,N_18928,N_20562);
nor U21732 (N_21732,N_19632,N_18674);
and U21733 (N_21733,N_20608,N_19466);
nand U21734 (N_21734,N_19095,N_20885);
and U21735 (N_21735,N_19279,N_18548);
and U21736 (N_21736,N_20246,N_19723);
and U21737 (N_21737,N_18249,N_19682);
and U21738 (N_21738,N_20250,N_19287);
or U21739 (N_21739,N_20293,N_20391);
or U21740 (N_21740,N_18003,N_19332);
and U21741 (N_21741,N_20153,N_20949);
or U21742 (N_21742,N_18913,N_19350);
nor U21743 (N_21743,N_18233,N_18635);
xor U21744 (N_21744,N_18300,N_19576);
nor U21745 (N_21745,N_18995,N_19333);
nor U21746 (N_21746,N_20995,N_19334);
nor U21747 (N_21747,N_18961,N_18399);
nor U21748 (N_21748,N_20902,N_20180);
or U21749 (N_21749,N_20462,N_19448);
or U21750 (N_21750,N_20942,N_18319);
xor U21751 (N_21751,N_20759,N_18835);
nand U21752 (N_21752,N_18324,N_19138);
nor U21753 (N_21753,N_18098,N_20248);
or U21754 (N_21754,N_19773,N_20701);
xor U21755 (N_21755,N_20384,N_18808);
nor U21756 (N_21756,N_19200,N_19179);
or U21757 (N_21757,N_20149,N_19859);
or U21758 (N_21758,N_19536,N_19824);
nor U21759 (N_21759,N_19522,N_19108);
nand U21760 (N_21760,N_20038,N_20799);
and U21761 (N_21761,N_19088,N_19078);
and U21762 (N_21762,N_19788,N_19130);
nor U21763 (N_21763,N_18203,N_18513);
and U21764 (N_21764,N_20394,N_20910);
and U21765 (N_21765,N_19098,N_19363);
or U21766 (N_21766,N_18172,N_20580);
and U21767 (N_21767,N_19421,N_18374);
and U21768 (N_21768,N_18282,N_18650);
nor U21769 (N_21769,N_20317,N_19086);
nand U21770 (N_21770,N_20635,N_19317);
nand U21771 (N_21771,N_18369,N_18405);
or U21772 (N_21772,N_18494,N_20796);
and U21773 (N_21773,N_18125,N_19708);
nand U21774 (N_21774,N_18766,N_18342);
nor U21775 (N_21775,N_18455,N_18955);
nand U21776 (N_21776,N_20218,N_19339);
and U21777 (N_21777,N_18234,N_19182);
nand U21778 (N_21778,N_19742,N_20943);
xnor U21779 (N_21779,N_18093,N_20200);
or U21780 (N_21780,N_19670,N_20809);
or U21781 (N_21781,N_18580,N_18547);
and U21782 (N_21782,N_18476,N_19627);
nand U21783 (N_21783,N_20974,N_19523);
and U21784 (N_21784,N_18529,N_18150);
xnor U21785 (N_21785,N_18467,N_20543);
or U21786 (N_21786,N_20416,N_20326);
and U21787 (N_21787,N_19814,N_20836);
or U21788 (N_21788,N_20663,N_18729);
nor U21789 (N_21789,N_18206,N_18326);
nor U21790 (N_21790,N_18915,N_18941);
or U21791 (N_21791,N_19748,N_20467);
or U21792 (N_21792,N_18667,N_19052);
or U21793 (N_21793,N_20630,N_20357);
xnor U21794 (N_21794,N_20078,N_19169);
nand U21795 (N_21795,N_18267,N_20883);
xor U21796 (N_21796,N_18533,N_20827);
or U21797 (N_21797,N_19538,N_19775);
and U21798 (N_21798,N_18133,N_19412);
and U21799 (N_21799,N_20741,N_18164);
nand U21800 (N_21800,N_18550,N_19259);
and U21801 (N_21801,N_19134,N_19175);
or U21802 (N_21802,N_18903,N_19288);
nand U21803 (N_21803,N_20279,N_18132);
nor U21804 (N_21804,N_18420,N_19686);
and U21805 (N_21805,N_19356,N_18426);
nor U21806 (N_21806,N_18169,N_18749);
xor U21807 (N_21807,N_18165,N_20161);
nor U21808 (N_21808,N_19302,N_18224);
nand U21809 (N_21809,N_20048,N_18617);
and U21810 (N_21810,N_20204,N_19790);
or U21811 (N_21811,N_18277,N_20969);
nor U21812 (N_21812,N_19657,N_20036);
or U21813 (N_21813,N_20795,N_18890);
or U21814 (N_21814,N_20930,N_19441);
nor U21815 (N_21815,N_19462,N_20383);
xnor U21816 (N_21816,N_19951,N_19979);
nor U21817 (N_21817,N_18071,N_20094);
and U21818 (N_21818,N_20539,N_18611);
nand U21819 (N_21819,N_18840,N_20762);
nor U21820 (N_21820,N_18040,N_19068);
and U21821 (N_21821,N_19150,N_19207);
and U21822 (N_21822,N_18195,N_19481);
nor U21823 (N_21823,N_20237,N_20434);
nor U21824 (N_21824,N_18077,N_18444);
or U21825 (N_21825,N_18688,N_20642);
nor U21826 (N_21826,N_20404,N_20596);
nor U21827 (N_21827,N_18037,N_20950);
xor U21828 (N_21828,N_18888,N_20110);
and U21829 (N_21829,N_20514,N_20185);
and U21830 (N_21830,N_19604,N_19940);
or U21831 (N_21831,N_18211,N_19850);
or U21832 (N_21832,N_20179,N_18155);
nand U21833 (N_21833,N_18480,N_20345);
nor U21834 (N_21834,N_20397,N_20880);
and U21835 (N_21835,N_20674,N_18339);
nor U21836 (N_21836,N_19045,N_18885);
and U21837 (N_21837,N_18578,N_20166);
or U21838 (N_21838,N_20877,N_20547);
and U21839 (N_21839,N_18288,N_18008);
nand U21840 (N_21840,N_20271,N_20194);
and U21841 (N_21841,N_18153,N_18411);
or U21842 (N_21842,N_20239,N_18945);
xnor U21843 (N_21843,N_19084,N_18244);
nor U21844 (N_21844,N_18514,N_18644);
nor U21845 (N_21845,N_18251,N_20574);
nor U21846 (N_21846,N_20779,N_19569);
or U21847 (N_21847,N_19390,N_19672);
and U21848 (N_21848,N_18236,N_19581);
or U21849 (N_21849,N_18404,N_20084);
xor U21850 (N_21850,N_19375,N_19930);
and U21851 (N_21851,N_19876,N_19061);
nor U21852 (N_21852,N_18735,N_18697);
nand U21853 (N_21853,N_20448,N_19443);
and U21854 (N_21854,N_18980,N_20913);
xnor U21855 (N_21855,N_18296,N_19149);
or U21856 (N_21856,N_20920,N_19870);
and U21857 (N_21857,N_18612,N_19430);
or U21858 (N_21858,N_19623,N_19113);
xnor U21859 (N_21859,N_19820,N_20432);
nand U21860 (N_21860,N_19970,N_18668);
or U21861 (N_21861,N_19122,N_20044);
and U21862 (N_21862,N_20748,N_19346);
nor U21863 (N_21863,N_18661,N_20157);
nand U21864 (N_21864,N_18180,N_20778);
or U21865 (N_21865,N_18015,N_19740);
and U21866 (N_21866,N_19935,N_18605);
and U21867 (N_21867,N_19891,N_20223);
xnor U21868 (N_21868,N_18097,N_18702);
nand U21869 (N_21869,N_18469,N_20016);
nand U21870 (N_21870,N_19994,N_18882);
nor U21871 (N_21871,N_19712,N_18517);
and U21872 (N_21872,N_20996,N_18850);
and U21873 (N_21873,N_19526,N_20360);
nand U21874 (N_21874,N_19533,N_18914);
nor U21875 (N_21875,N_20087,N_19102);
nand U21876 (N_21876,N_19250,N_20460);
nand U21877 (N_21877,N_19222,N_20300);
nor U21878 (N_21878,N_20896,N_19428);
or U21879 (N_21879,N_19719,N_20083);
nand U21880 (N_21880,N_19048,N_20712);
or U21881 (N_21881,N_19121,N_18649);
xnor U21882 (N_21882,N_19025,N_18198);
or U21883 (N_21883,N_20754,N_19204);
and U21884 (N_21884,N_19261,N_20296);
and U21885 (N_21885,N_20274,N_19527);
nor U21886 (N_21886,N_19091,N_18630);
nand U21887 (N_21887,N_20433,N_20323);
nor U21888 (N_21888,N_18368,N_18643);
nand U21889 (N_21889,N_18281,N_20965);
nand U21890 (N_21890,N_19620,N_20403);
and U21891 (N_21891,N_19431,N_18768);
or U21892 (N_21892,N_18304,N_20550);
nor U21893 (N_21893,N_18947,N_18553);
or U21894 (N_21894,N_19785,N_20519);
or U21895 (N_21895,N_19117,N_18737);
nor U21896 (N_21896,N_18799,N_18209);
nor U21897 (N_21897,N_19439,N_20815);
or U21898 (N_21898,N_20085,N_20373);
nor U21899 (N_21899,N_20431,N_20624);
nor U21900 (N_21900,N_18616,N_20411);
and U21901 (N_21901,N_18930,N_18349);
or U21902 (N_21902,N_18614,N_20564);
or U21903 (N_21903,N_18784,N_20620);
nand U21904 (N_21904,N_19217,N_19241);
nand U21905 (N_21905,N_19865,N_18592);
nand U21906 (N_21906,N_19220,N_20165);
xor U21907 (N_21907,N_20939,N_18503);
and U21908 (N_21908,N_20205,N_20025);
and U21909 (N_21909,N_20702,N_18884);
nor U21910 (N_21910,N_19881,N_20281);
or U21911 (N_21911,N_18156,N_18265);
or U21912 (N_21912,N_19373,N_18588);
xor U21913 (N_21913,N_19154,N_18408);
nor U21914 (N_21914,N_20441,N_19806);
xnor U21915 (N_21915,N_19311,N_19908);
xnor U21916 (N_21916,N_20159,N_18781);
or U21917 (N_21917,N_18889,N_20537);
and U21918 (N_21918,N_20504,N_18861);
nor U21919 (N_21919,N_18647,N_20276);
xor U21920 (N_21920,N_19372,N_19675);
and U21921 (N_21921,N_18188,N_20887);
nand U21922 (N_21922,N_19779,N_19524);
nor U21923 (N_21923,N_19063,N_20242);
xnor U21924 (N_21924,N_18245,N_18393);
or U21925 (N_21925,N_19274,N_19566);
nor U21926 (N_21926,N_19137,N_19297);
and U21927 (N_21927,N_18764,N_20540);
nand U21928 (N_21928,N_18815,N_18899);
or U21929 (N_21929,N_19842,N_18268);
and U21930 (N_21930,N_20505,N_20295);
and U21931 (N_21931,N_19271,N_18022);
xnor U21932 (N_21932,N_18247,N_19746);
xor U21933 (N_21933,N_20485,N_20619);
and U21934 (N_21934,N_19065,N_19483);
and U21935 (N_21935,N_19383,N_19020);
nor U21936 (N_21936,N_19417,N_19901);
and U21937 (N_21937,N_19256,N_18990);
nor U21938 (N_21938,N_19926,N_18821);
xor U21939 (N_21939,N_18528,N_20270);
xor U21940 (N_21940,N_19313,N_19949);
or U21941 (N_21941,N_18308,N_20106);
nand U21942 (N_21942,N_18317,N_20032);
nand U21943 (N_21943,N_19128,N_20221);
or U21944 (N_21944,N_18567,N_18028);
nor U21945 (N_21945,N_19015,N_20746);
nand U21946 (N_21946,N_18590,N_18851);
nand U21947 (N_21947,N_20724,N_18159);
xor U21948 (N_21948,N_19189,N_18024);
and U21949 (N_21949,N_20265,N_19813);
or U21950 (N_21950,N_18862,N_19368);
or U21951 (N_21951,N_18786,N_18048);
nor U21952 (N_21952,N_20893,N_18925);
xor U21953 (N_21953,N_18967,N_20342);
or U21954 (N_21954,N_20443,N_19474);
nor U21955 (N_21955,N_20186,N_20301);
and U21956 (N_21956,N_19456,N_18852);
nand U21957 (N_21957,N_18027,N_20677);
nand U21958 (N_21958,N_20837,N_19809);
and U21959 (N_21959,N_18378,N_19110);
and U21960 (N_21960,N_18457,N_18754);
or U21961 (N_21961,N_20241,N_18633);
and U21962 (N_21962,N_20568,N_19614);
xnor U21963 (N_21963,N_20028,N_19035);
nor U21964 (N_21964,N_19906,N_18149);
nor U21965 (N_21965,N_19482,N_18703);
xnor U21966 (N_21966,N_19206,N_18250);
nand U21967 (N_21967,N_19438,N_19553);
and U21968 (N_21968,N_19201,N_19552);
or U21969 (N_21969,N_18121,N_20652);
nand U21970 (N_21970,N_20844,N_20037);
and U21971 (N_21971,N_18185,N_18810);
or U21972 (N_21972,N_20463,N_18053);
nand U21973 (N_21973,N_20722,N_20631);
nand U21974 (N_21974,N_20679,N_20685);
or U21975 (N_21975,N_19920,N_18168);
nor U21976 (N_21976,N_20289,N_18919);
or U21977 (N_21977,N_20900,N_19848);
nand U21978 (N_21978,N_19385,N_18723);
and U21979 (N_21979,N_19440,N_18147);
and U21980 (N_21980,N_19922,N_18332);
xor U21981 (N_21981,N_18356,N_19101);
or U21982 (N_21982,N_20615,N_19575);
nand U21983 (N_21983,N_18289,N_18695);
nand U21984 (N_21984,N_18490,N_20990);
and U21985 (N_21985,N_19877,N_19611);
nand U21986 (N_21986,N_20364,N_18740);
nand U21987 (N_21987,N_19937,N_18966);
nor U21988 (N_21988,N_20408,N_20981);
nand U21989 (N_21989,N_18847,N_19177);
nor U21990 (N_21990,N_20447,N_20169);
or U21991 (N_21991,N_20174,N_20303);
and U21992 (N_21992,N_19953,N_18307);
xnor U21993 (N_21993,N_18345,N_19905);
or U21994 (N_21994,N_18019,N_20097);
and U21995 (N_21995,N_20868,N_20895);
xnor U21996 (N_21996,N_18566,N_19818);
nor U21997 (N_21997,N_20017,N_19792);
nor U21998 (N_21998,N_20494,N_19419);
nor U21999 (N_21999,N_19823,N_19643);
or U22000 (N_22000,N_19034,N_19433);
and U22001 (N_22001,N_19314,N_20774);
nor U22002 (N_22002,N_19284,N_18218);
nand U22003 (N_22003,N_19691,N_19914);
and U22004 (N_22004,N_18438,N_19029);
xor U22005 (N_22005,N_20262,N_18673);
and U22006 (N_22006,N_20484,N_19543);
and U22007 (N_22007,N_20366,N_18372);
or U22008 (N_22008,N_20546,N_19796);
nand U22009 (N_22009,N_19947,N_19265);
nand U22010 (N_22010,N_19986,N_18205);
and U22011 (N_22011,N_19503,N_18299);
or U22012 (N_22012,N_18074,N_20111);
and U22013 (N_22013,N_18190,N_20483);
or U22014 (N_22014,N_18463,N_19638);
and U22015 (N_22015,N_18637,N_19074);
or U22016 (N_22016,N_18252,N_20841);
nand U22017 (N_22017,N_18398,N_19186);
nand U22018 (N_22018,N_18173,N_18083);
and U22019 (N_22019,N_19072,N_18435);
and U22020 (N_22020,N_20609,N_19645);
nor U22021 (N_22021,N_18333,N_18628);
and U22022 (N_22022,N_20379,N_20334);
nor U22023 (N_22023,N_20283,N_20854);
and U22024 (N_22024,N_18392,N_18620);
nor U22025 (N_22025,N_19841,N_19161);
or U22026 (N_22026,N_19165,N_18521);
nand U22027 (N_22027,N_18940,N_19355);
and U22028 (N_22028,N_19402,N_19535);
or U22029 (N_22029,N_20727,N_19759);
nor U22030 (N_22030,N_20711,N_20446);
nand U22031 (N_22031,N_20618,N_18972);
and U22032 (N_22032,N_18515,N_20059);
and U22033 (N_22033,N_19040,N_20254);
nand U22034 (N_22034,N_18820,N_20704);
xnor U22035 (N_22035,N_19764,N_18734);
nand U22036 (N_22036,N_19185,N_18331);
and U22037 (N_22037,N_18240,N_18511);
nand U22038 (N_22038,N_20376,N_18202);
or U22039 (N_22039,N_20164,N_18454);
xor U22040 (N_22040,N_18375,N_18338);
nor U22041 (N_22041,N_18538,N_20874);
or U22042 (N_22042,N_20058,N_20368);
or U22043 (N_22043,N_20788,N_19909);
nor U22044 (N_22044,N_18502,N_18220);
or U22045 (N_22045,N_19634,N_18658);
nor U22046 (N_22046,N_19221,N_19897);
nor U22047 (N_22047,N_20632,N_18579);
xor U22048 (N_22048,N_19766,N_20520);
nor U22049 (N_22049,N_19789,N_18909);
nor U22050 (N_22050,N_20176,N_19338);
nand U22051 (N_22051,N_20914,N_19406);
nor U22052 (N_22052,N_19413,N_18363);
xor U22053 (N_22053,N_18129,N_19886);
or U22054 (N_22054,N_18360,N_18868);
and U22055 (N_22055,N_20280,N_20136);
nand U22056 (N_22056,N_20859,N_20726);
or U22057 (N_22057,N_18968,N_19348);
xor U22058 (N_22058,N_20490,N_20901);
xor U22059 (N_22059,N_20122,N_19382);
or U22060 (N_22060,N_19547,N_19459);
and U22061 (N_22061,N_20336,N_18228);
nand U22062 (N_22062,N_20558,N_19827);
and U22063 (N_22063,N_19142,N_18230);
xnor U22064 (N_22064,N_18920,N_20199);
and U22065 (N_22065,N_20292,N_18416);
and U22066 (N_22066,N_19181,N_20612);
and U22067 (N_22067,N_18726,N_19941);
nand U22068 (N_22068,N_19225,N_19367);
and U22069 (N_22069,N_19887,N_18975);
and U22070 (N_22070,N_20850,N_20354);
nand U22071 (N_22071,N_20610,N_18911);
or U22072 (N_22072,N_20103,N_19862);
nor U22073 (N_22073,N_19562,N_19900);
or U22074 (N_22074,N_20793,N_19229);
or U22075 (N_22075,N_18437,N_19701);
nor U22076 (N_22076,N_20831,N_20233);
and U22077 (N_22077,N_18520,N_19520);
and U22078 (N_22078,N_18944,N_18341);
nor U22079 (N_22079,N_20668,N_18818);
and U22080 (N_22080,N_19688,N_18012);
nand U22081 (N_22081,N_20852,N_20027);
or U22082 (N_22082,N_18554,N_20503);
nand U22083 (N_22083,N_20480,N_20904);
nand U22084 (N_22084,N_18937,N_20385);
xnor U22085 (N_22085,N_19414,N_18497);
and U22086 (N_22086,N_19044,N_20653);
and U22087 (N_22087,N_18670,N_20260);
nor U22088 (N_22088,N_19236,N_18235);
or U22089 (N_22089,N_19162,N_20442);
and U22090 (N_22090,N_19294,N_20623);
nor U22091 (N_22091,N_18537,N_20890);
xnor U22092 (N_22092,N_19858,N_19864);
or U22093 (N_22093,N_20586,N_20310);
and U22094 (N_22094,N_18651,N_18225);
or U22095 (N_22095,N_19975,N_18759);
nor U22096 (N_22096,N_19487,N_20605);
or U22097 (N_22097,N_18403,N_20266);
xor U22098 (N_22098,N_20683,N_20957);
or U22099 (N_22099,N_18295,N_18271);
and U22100 (N_22100,N_19957,N_19475);
xnor U22101 (N_22101,N_19379,N_18585);
nand U22102 (N_22102,N_19423,N_18916);
nor U22103 (N_22103,N_18860,N_19254);
and U22104 (N_22104,N_20006,N_18062);
nand U22105 (N_22105,N_20511,N_19863);
and U22106 (N_22106,N_20734,N_20994);
or U22107 (N_22107,N_20181,N_19925);
nor U22108 (N_22108,N_19031,N_19703);
nand U22109 (N_22109,N_19342,N_20829);
and U22110 (N_22110,N_20959,N_20744);
or U22111 (N_22111,N_19570,N_20298);
xor U22112 (N_22112,N_19851,N_19315);
nand U22113 (N_22113,N_20335,N_19432);
and U22114 (N_22114,N_18878,N_19012);
or U22115 (N_22115,N_20713,N_19488);
nand U22116 (N_22116,N_19966,N_19720);
and U22117 (N_22117,N_18733,N_19684);
and U22118 (N_22118,N_19416,N_20639);
nor U22119 (N_22119,N_19184,N_20661);
nor U22120 (N_22120,N_18577,N_18962);
nor U22121 (N_22121,N_18105,N_20763);
or U22122 (N_22122,N_18046,N_20688);
nor U22123 (N_22123,N_20579,N_19151);
and U22124 (N_22124,N_20487,N_19619);
nand U22125 (N_22125,N_19164,N_18117);
or U22126 (N_22126,N_20925,N_19062);
or U22127 (N_22127,N_18328,N_20116);
or U22128 (N_22128,N_18739,N_18413);
nand U22129 (N_22129,N_18826,N_20131);
and U22130 (N_22130,N_19613,N_19451);
nor U22131 (N_22131,N_19736,N_18595);
nor U22132 (N_22132,N_18894,N_20501);
or U22133 (N_22133,N_18711,N_18440);
nor U22134 (N_22134,N_20773,N_20104);
nor U22135 (N_22135,N_18007,N_20571);
and U22136 (N_22136,N_18516,N_20671);
and U22137 (N_22137,N_19910,N_20320);
or U22138 (N_22138,N_18831,N_20337);
nand U22139 (N_22139,N_20243,N_18794);
nand U22140 (N_22140,N_18321,N_19943);
nor U22141 (N_22141,N_18213,N_20828);
nand U22142 (N_22142,N_19880,N_18361);
and U22143 (N_22143,N_19653,N_18957);
and U22144 (N_22144,N_18657,N_20770);
and U22145 (N_22145,N_20018,N_19324);
xor U22146 (N_22146,N_19255,N_19784);
nor U22147 (N_22147,N_19335,N_20805);
nor U22148 (N_22148,N_19945,N_19469);
or U22149 (N_22149,N_18978,N_19027);
or U22150 (N_22150,N_19127,N_18993);
nand U22151 (N_22151,N_20684,N_19277);
and U22152 (N_22152,N_18309,N_18466);
nand U22153 (N_22153,N_19508,N_18166);
nand U22154 (N_22154,N_20047,N_20130);
and U22155 (N_22155,N_19496,N_20565);
nand U22156 (N_22156,N_18788,N_19485);
nand U22157 (N_22157,N_20330,N_19156);
or U22158 (N_22158,N_19861,N_19252);
and U22159 (N_22159,N_20261,N_18698);
nand U22160 (N_22160,N_20191,N_20692);
xor U22161 (N_22161,N_20324,N_19452);
and U22162 (N_22162,N_18280,N_19424);
and U22163 (N_22163,N_19767,N_20147);
nand U22164 (N_22164,N_20597,N_20889);
and U22165 (N_22165,N_18453,N_19934);
nor U22166 (N_22166,N_20107,N_19446);
nand U22167 (N_22167,N_18656,N_20052);
nand U22168 (N_22168,N_20673,N_18730);
or U22169 (N_22169,N_19810,N_18887);
nor U22170 (N_22170,N_19081,N_18663);
or U22171 (N_22171,N_19793,N_20948);
nand U22172 (N_22172,N_18965,N_20290);
and U22173 (N_22173,N_18227,N_18828);
and U22174 (N_22174,N_19919,N_19625);
or U22175 (N_22175,N_20050,N_19191);
nor U22176 (N_22176,N_19275,N_18684);
or U22177 (N_22177,N_20733,N_20117);
xor U22178 (N_22178,N_19615,N_18958);
nor U22179 (N_22179,N_18951,N_19642);
nor U22180 (N_22180,N_20211,N_19607);
or U22181 (N_22181,N_20732,N_20932);
nor U22182 (N_22182,N_20074,N_18785);
nor U22183 (N_22183,N_20736,N_18192);
nor U22184 (N_22184,N_18714,N_20375);
nor U22185 (N_22185,N_18604,N_18418);
or U22186 (N_22186,N_19163,N_18565);
nor U22187 (N_22187,N_18834,N_18439);
nor U22188 (N_22188,N_20352,N_19420);
nor U22189 (N_22189,N_18780,N_20389);
or U22190 (N_22190,N_19060,N_19903);
and U22191 (N_22191,N_20958,N_19144);
nand U22192 (N_22192,N_19109,N_20412);
nor U22193 (N_22193,N_19721,N_20875);
or U22194 (N_22194,N_19548,N_19836);
xnor U22195 (N_22195,N_18570,N_19772);
or U22196 (N_22196,N_18545,N_19892);
and U22197 (N_22197,N_19661,N_20944);
nor U22198 (N_22198,N_20790,N_20557);
and U22199 (N_22199,N_18272,N_19753);
nand U22200 (N_22200,N_20363,N_19855);
nor U22201 (N_22201,N_18485,N_19585);
nor U22202 (N_22202,N_18270,N_18189);
or U22203 (N_22203,N_19592,N_19898);
and U22204 (N_22204,N_18607,N_18672);
and U22205 (N_22205,N_20219,N_18600);
nand U22206 (N_22206,N_20370,N_20418);
xnor U22207 (N_22207,N_20506,N_18160);
xnor U22208 (N_22208,N_18241,N_20526);
and U22209 (N_22209,N_18187,N_19993);
or U22210 (N_22210,N_18142,N_19337);
nand U22211 (N_22211,N_18347,N_20525);
and U22212 (N_22212,N_20013,N_18526);
xor U22213 (N_22213,N_18546,N_18816);
and U22214 (N_22214,N_18158,N_18998);
or U22215 (N_22215,N_20141,N_19016);
nand U22216 (N_22216,N_18468,N_19963);
nor U22217 (N_22217,N_20438,N_18226);
and U22218 (N_22218,N_18273,N_20372);
nor U22219 (N_22219,N_18076,N_20119);
xnor U22220 (N_22220,N_20695,N_18927);
or U22221 (N_22221,N_18601,N_19973);
nor U22222 (N_22222,N_20705,N_20905);
nor U22223 (N_22223,N_20784,N_19077);
or U22224 (N_22224,N_19882,N_20039);
and U22225 (N_22225,N_20488,N_19781);
or U22226 (N_22226,N_19468,N_20553);
nand U22227 (N_22227,N_20697,N_20802);
and U22228 (N_22228,N_20152,N_20808);
nand U22229 (N_22229,N_19227,N_19554);
nor U22230 (N_22230,N_20294,N_19884);
and U22231 (N_22231,N_19097,N_18921);
xnor U22232 (N_22232,N_20807,N_20549);
or U22233 (N_22233,N_20719,N_18534);
xor U22234 (N_22234,N_20228,N_20054);
and U22235 (N_22235,N_19384,N_18286);
nor U22236 (N_22236,N_20091,N_19361);
and U22237 (N_22237,N_19867,N_19014);
xor U22238 (N_22238,N_18284,N_18541);
or U22239 (N_22239,N_20810,N_18086);
and U22240 (N_22240,N_19397,N_19665);
nand U22241 (N_22241,N_20088,N_20158);
or U22242 (N_22242,N_20548,N_19730);
and U22243 (N_22243,N_20451,N_20751);
xor U22244 (N_22244,N_20919,N_19579);
nor U22245 (N_22245,N_18026,N_19024);
nand U22246 (N_22246,N_18910,N_20259);
or U22247 (N_22247,N_20424,N_19231);
nor U22248 (N_22248,N_20064,N_19411);
nor U22249 (N_22249,N_18522,N_18693);
nand U22250 (N_22250,N_18124,N_18905);
or U22251 (N_22251,N_20244,N_20966);
and U22252 (N_22252,N_18412,N_19251);
nand U22253 (N_22253,N_19907,N_18113);
or U22254 (N_22254,N_18410,N_18348);
or U22255 (N_22255,N_19760,N_19418);
or U22256 (N_22256,N_18433,N_20737);
nand U22257 (N_22257,N_19677,N_19769);
and U22258 (N_22258,N_20811,N_18557);
nand U22259 (N_22259,N_19133,N_18701);
xnor U22260 (N_22260,N_19198,N_19043);
or U22261 (N_22261,N_18100,N_20049);
and U22262 (N_22262,N_18118,N_20934);
nand U22263 (N_22263,N_19010,N_20529);
and U22264 (N_22264,N_19264,N_18066);
nand U22265 (N_22265,N_20347,N_18424);
nor U22266 (N_22266,N_19209,N_18358);
or U22267 (N_22267,N_19690,N_18447);
nor U22268 (N_22268,N_19026,N_18897);
nor U22269 (N_22269,N_20459,N_19099);
nand U22270 (N_22270,N_18182,N_20715);
nand U22271 (N_22271,N_18127,N_19644);
or U22272 (N_22272,N_19659,N_20472);
or U22273 (N_22273,N_19783,N_19660);
xnor U22274 (N_22274,N_20863,N_19786);
and U22275 (N_22275,N_20220,N_20203);
nand U22276 (N_22276,N_20399,N_18942);
xor U22277 (N_22277,N_18038,N_18683);
nor U22278 (N_22278,N_18078,N_18079);
or U22279 (N_22279,N_20843,N_20953);
or U22280 (N_22280,N_19808,N_18902);
and U22281 (N_22281,N_20644,N_19238);
nor U22282 (N_22282,N_18464,N_18069);
or U22283 (N_22283,N_20208,N_18807);
and U22284 (N_22284,N_18103,N_18114);
nand U22285 (N_22285,N_18560,N_20479);
nand U22286 (N_22286,N_19801,N_20765);
and U22287 (N_22287,N_19089,N_20435);
nor U22288 (N_22288,N_18141,N_19105);
nor U22289 (N_22289,N_19843,N_19310);
nor U22290 (N_22290,N_18682,N_18390);
nand U22291 (N_22291,N_20010,N_20369);
or U22292 (N_22292,N_20952,N_19911);
nor U22293 (N_22293,N_19555,N_18770);
or U22294 (N_22294,N_19422,N_19717);
nor U22295 (N_22295,N_20502,N_18116);
nor U22296 (N_22296,N_20993,N_20313);
xor U22297 (N_22297,N_20041,N_20906);
or U22298 (N_22298,N_20598,N_18018);
or U22299 (N_22299,N_20331,N_18933);
or U22300 (N_22300,N_19371,N_20676);
and U22301 (N_22301,N_18809,N_20454);
or U22302 (N_22302,N_20351,N_18696);
nor U22303 (N_22303,N_19205,N_18720);
or U22304 (N_22304,N_18856,N_19729);
nand U22305 (N_22305,N_20961,N_20634);
and U22306 (N_22306,N_18898,N_18977);
and U22307 (N_22307,N_19916,N_20081);
nand U22308 (N_22308,N_18746,N_18419);
or U22309 (N_22309,N_19505,N_18624);
or U22310 (N_22310,N_20846,N_18609);
and U22311 (N_22311,N_20022,N_20946);
nor U22312 (N_22312,N_18777,N_18109);
and U22313 (N_22313,N_19825,N_18355);
nand U22314 (N_22314,N_18207,N_20769);
and U22315 (N_22315,N_19239,N_18470);
or U22316 (N_22316,N_20651,N_20227);
nand U22317 (N_22317,N_19968,N_20757);
nand U22318 (N_22318,N_20760,N_20409);
nor U22319 (N_22319,N_20109,N_20823);
and U22320 (N_22320,N_20137,N_19325);
and U22321 (N_22321,N_19041,N_18343);
or U22322 (N_22322,N_18380,N_19872);
and U22323 (N_22323,N_19511,N_18434);
nor U22324 (N_22324,N_19501,N_19364);
nand U22325 (N_22325,N_19560,N_20718);
nand U22326 (N_22326,N_19658,N_20721);
nor U22327 (N_22327,N_20589,N_20803);
and U22328 (N_22328,N_19234,N_18415);
nor U22329 (N_22329,N_20709,N_19080);
or U22330 (N_22330,N_19476,N_18495);
xor U22331 (N_22331,N_20138,N_20491);
nor U22332 (N_22332,N_20124,N_20785);
nor U22333 (N_22333,N_18099,N_20437);
xnor U22334 (N_22334,N_19224,N_18871);
and U22335 (N_22335,N_18314,N_20816);
nor U22336 (N_22336,N_20341,N_20114);
nor U22337 (N_22337,N_20092,N_20198);
nand U22338 (N_22338,N_18014,N_20522);
and U22339 (N_22339,N_19263,N_18631);
and U22340 (N_22340,N_18085,N_20781);
and U22341 (N_22341,N_18983,N_19005);
nand U22342 (N_22342,N_18186,N_19542);
nand U22343 (N_22343,N_20694,N_18791);
nand U22344 (N_22344,N_18427,N_19380);
or U22345 (N_22345,N_19888,N_18866);
xor U22346 (N_22346,N_20613,N_18035);
nor U22347 (N_22347,N_20287,N_18474);
nand U22348 (N_22348,N_18773,N_18334);
and U22349 (N_22349,N_18636,N_20862);
nor U22350 (N_22350,N_18487,N_20776);
xnor U22351 (N_22351,N_20847,N_20659);
and U22352 (N_22352,N_20269,N_20188);
or U22353 (N_22353,N_18691,N_19561);
or U22354 (N_22354,N_19210,N_19465);
and U22355 (N_22355,N_19664,N_19491);
or U22356 (N_22356,N_20592,N_20202);
nand U22357 (N_22357,N_19992,N_19358);
or U22358 (N_22358,N_18762,N_19743);
and U22359 (N_22359,N_20302,N_20140);
and U22360 (N_22360,N_19573,N_20975);
or U22361 (N_22361,N_19394,N_18671);
nand U22362 (N_22362,N_20864,N_18020);
or U22363 (N_22363,N_19856,N_20349);
or U22364 (N_22364,N_20817,N_18353);
or U22365 (N_22365,N_20316,N_18827);
nand U22366 (N_22366,N_20838,N_20187);
or U22367 (N_22367,N_18582,N_20095);
nand U22368 (N_22368,N_18772,N_20255);
or U22369 (N_22369,N_20288,N_18877);
and U22370 (N_22370,N_18481,N_20541);
nand U22371 (N_22371,N_19087,N_19895);
nor U22372 (N_22372,N_18493,N_20105);
nor U22373 (N_22373,N_18387,N_19889);
nor U22374 (N_22374,N_19159,N_20073);
nor U22375 (N_22375,N_20999,N_18335);
nand U22376 (N_22376,N_20496,N_20640);
xor U22377 (N_22377,N_20782,N_18446);
or U22378 (N_22378,N_19778,N_20077);
and U22379 (N_22379,N_18017,N_19636);
nand U22380 (N_22380,N_18088,N_20040);
and U22381 (N_22381,N_20020,N_20471);
and U22382 (N_22382,N_19871,N_20606);
nor U22383 (N_22383,N_18660,N_19351);
or U22384 (N_22384,N_18505,N_19013);
nor U22385 (N_22385,N_20133,N_20645);
and U22386 (N_22386,N_20654,N_20308);
and U22387 (N_22387,N_20053,N_20429);
nor U22388 (N_22388,N_18728,N_18872);
xnor U22389 (N_22389,N_19990,N_18742);
or U22390 (N_22390,N_18064,N_18997);
or U22391 (N_22391,N_19915,N_18212);
nand U22392 (N_22392,N_18002,N_20318);
and U22393 (N_22393,N_20566,N_20622);
nor U22394 (N_22394,N_20458,N_19114);
nor U22395 (N_22395,N_19240,N_19698);
nand U22396 (N_22396,N_19400,N_19094);
xor U22397 (N_22397,N_19588,N_19244);
and U22398 (N_22398,N_20497,N_19707);
or U22399 (N_22399,N_19699,N_19662);
nor U22400 (N_22400,N_18472,N_20299);
and U22401 (N_22401,N_18923,N_18679);
nor U22402 (N_22402,N_18716,N_19057);
and U22403 (N_22403,N_19442,N_18279);
nor U22404 (N_22404,N_18303,N_18414);
or U22405 (N_22405,N_18060,N_18789);
nand U22406 (N_22406,N_18971,N_18110);
nor U22407 (N_22407,N_19023,N_20386);
xnor U22408 (N_22408,N_19605,N_18855);
xor U22409 (N_22409,N_18219,N_18699);
and U22410 (N_22410,N_18054,N_19869);
nor U22411 (N_22411,N_20933,N_19321);
or U22412 (N_22412,N_20031,N_19618);
nor U22413 (N_22413,N_19752,N_18869);
xnor U22414 (N_22414,N_18865,N_20611);
and U22415 (N_22415,N_19812,N_19798);
nor U22416 (N_22416,N_18323,N_18648);
or U22417 (N_22417,N_18432,N_20510);
xnor U22418 (N_22418,N_20190,N_20917);
nor U22419 (N_22419,N_18717,N_20102);
nor U22420 (N_22420,N_18197,N_20089);
or U22421 (N_22421,N_18680,N_19037);
nor U22422 (N_22422,N_20929,N_19399);
nor U22423 (N_22423,N_20989,N_20071);
nand U22424 (N_22424,N_18001,N_18082);
nor U22425 (N_22425,N_19187,N_18061);
or U22426 (N_22426,N_19453,N_20800);
or U22427 (N_22427,N_19822,N_18664);
and U22428 (N_22428,N_20693,N_18367);
nand U22429 (N_22429,N_20753,N_19594);
xor U22430 (N_22430,N_19376,N_19002);
nand U22431 (N_22431,N_18954,N_18266);
xnor U22432 (N_22432,N_19679,N_20840);
and U22433 (N_22433,N_20752,N_20797);
and U22434 (N_22434,N_19695,N_20307);
nor U22435 (N_22435,N_18030,N_20708);
xnor U22436 (N_22436,N_19668,N_18120);
xor U22437 (N_22437,N_20498,N_19633);
nand U22438 (N_22438,N_18718,N_18283);
xnor U22439 (N_22439,N_18938,N_18793);
or U22440 (N_22440,N_18261,N_20937);
nand U22441 (N_22441,N_20311,N_19237);
nand U22442 (N_22442,N_20918,N_18406);
and U22443 (N_22443,N_18486,N_20388);
or U22444 (N_22444,N_18583,N_18575);
xor U22445 (N_22445,N_19927,N_20224);
or U22446 (N_22446,N_19750,N_20665);
nand U22447 (N_22447,N_19280,N_19076);
and U22448 (N_22448,N_18858,N_20599);
or U22449 (N_22449,N_19890,N_19838);
or U22450 (N_22450,N_19286,N_19762);
nand U22451 (N_22451,N_19006,N_18080);
nand U22452 (N_22452,N_19651,N_19509);
and U22453 (N_22453,N_20699,N_20621);
nand U22454 (N_22454,N_20960,N_19404);
nor U22455 (N_22455,N_18629,N_19574);
nor U22456 (N_22456,N_20600,N_18389);
or U22457 (N_22457,N_18031,N_20478);
nor U22458 (N_22458,N_20113,N_18385);
nand U22459 (N_22459,N_20672,N_20090);
or U22460 (N_22460,N_18301,N_19612);
and U22461 (N_22461,N_20407,N_20806);
and U22462 (N_22462,N_20735,N_20012);
nand U22463 (N_22463,N_20214,N_19195);
and U22464 (N_22464,N_19971,N_19305);
or U22465 (N_22465,N_20804,N_19631);
and U22466 (N_22466,N_19844,N_18519);
or U22467 (N_22467,N_18705,N_20700);
nand U22468 (N_22468,N_18982,N_19857);
or U22469 (N_22469,N_18507,N_19780);
nand U22470 (N_22470,N_20348,N_18979);
xor U22471 (N_22471,N_19226,N_19038);
and U22472 (N_22472,N_18593,N_18891);
or U22473 (N_22473,N_20112,N_20764);
nand U22474 (N_22474,N_20029,N_19987);
nor U22475 (N_22475,N_19921,N_20578);
xnor U22476 (N_22476,N_19831,N_20745);
nand U22477 (N_22477,N_20912,N_19398);
or U22478 (N_22478,N_20938,N_20972);
and U22479 (N_22479,N_18819,N_20344);
xnor U22480 (N_22480,N_20414,N_20453);
or U22481 (N_22481,N_18436,N_18484);
xnor U22482 (N_22482,N_20469,N_20263);
and U22483 (N_22483,N_18221,N_19988);
or U22484 (N_22484,N_19950,N_20998);
xor U22485 (N_22485,N_19359,N_19157);
or U22486 (N_22486,N_20328,N_18039);
nand U22487 (N_22487,N_19694,N_20475);
and U22488 (N_22488,N_20493,N_19706);
nor U22489 (N_22489,N_20306,N_20268);
or U22490 (N_22490,N_19985,N_20405);
or U22491 (N_22491,N_19648,N_19654);
nor U22492 (N_22492,N_19208,N_19531);
or U22493 (N_22493,N_20643,N_19387);
nor U22494 (N_22494,N_20195,N_19829);
nor U22495 (N_22495,N_18081,N_20051);
and U22496 (N_22496,N_19093,N_18193);
or U22497 (N_22497,N_20466,N_19532);
xor U22498 (N_22498,N_19039,N_20267);
nand U22499 (N_22499,N_20660,N_20229);
and U22500 (N_22500,N_19414,N_18984);
nor U22501 (N_22501,N_20307,N_18571);
xnor U22502 (N_22502,N_20099,N_19073);
or U22503 (N_22503,N_20903,N_20344);
nor U22504 (N_22504,N_20137,N_19148);
nor U22505 (N_22505,N_20204,N_20510);
or U22506 (N_22506,N_20139,N_18634);
and U22507 (N_22507,N_19724,N_19476);
and U22508 (N_22508,N_19773,N_20239);
and U22509 (N_22509,N_20623,N_18302);
nor U22510 (N_22510,N_19582,N_19045);
or U22511 (N_22511,N_20879,N_19520);
nor U22512 (N_22512,N_20563,N_19085);
nand U22513 (N_22513,N_19336,N_20222);
or U22514 (N_22514,N_18388,N_20987);
nor U22515 (N_22515,N_20787,N_20120);
and U22516 (N_22516,N_19511,N_19821);
xnor U22517 (N_22517,N_19532,N_18692);
or U22518 (N_22518,N_19230,N_20993);
nand U22519 (N_22519,N_18254,N_18053);
or U22520 (N_22520,N_19382,N_19607);
nand U22521 (N_22521,N_20142,N_19571);
nand U22522 (N_22522,N_18680,N_18500);
or U22523 (N_22523,N_18547,N_19262);
nor U22524 (N_22524,N_20209,N_18331);
nand U22525 (N_22525,N_19510,N_20542);
nand U22526 (N_22526,N_20572,N_20237);
and U22527 (N_22527,N_19493,N_18988);
nand U22528 (N_22528,N_20681,N_18870);
and U22529 (N_22529,N_20260,N_19571);
and U22530 (N_22530,N_18283,N_20497);
nor U22531 (N_22531,N_19568,N_18197);
and U22532 (N_22532,N_18165,N_20940);
and U22533 (N_22533,N_20711,N_18250);
xor U22534 (N_22534,N_18325,N_20491);
nand U22535 (N_22535,N_20859,N_20918);
xnor U22536 (N_22536,N_18634,N_18098);
nand U22537 (N_22537,N_20626,N_20294);
or U22538 (N_22538,N_20060,N_19051);
or U22539 (N_22539,N_20516,N_19268);
nor U22540 (N_22540,N_19764,N_19858);
and U22541 (N_22541,N_20674,N_20656);
and U22542 (N_22542,N_20439,N_20408);
nand U22543 (N_22543,N_18726,N_20991);
or U22544 (N_22544,N_19413,N_20824);
or U22545 (N_22545,N_18151,N_19389);
nand U22546 (N_22546,N_18529,N_18450);
xor U22547 (N_22547,N_20384,N_20649);
nor U22548 (N_22548,N_18639,N_20122);
or U22549 (N_22549,N_19947,N_20584);
or U22550 (N_22550,N_19988,N_19836);
nand U22551 (N_22551,N_18350,N_18116);
nand U22552 (N_22552,N_19051,N_20375);
nand U22553 (N_22553,N_19883,N_18335);
nand U22554 (N_22554,N_18449,N_19785);
nand U22555 (N_22555,N_18019,N_20188);
or U22556 (N_22556,N_20489,N_18734);
nand U22557 (N_22557,N_20152,N_20342);
nor U22558 (N_22558,N_19205,N_19580);
nor U22559 (N_22559,N_18320,N_20071);
nor U22560 (N_22560,N_20578,N_19250);
or U22561 (N_22561,N_18839,N_19514);
xor U22562 (N_22562,N_18953,N_19937);
nand U22563 (N_22563,N_19583,N_19842);
nor U22564 (N_22564,N_18319,N_18689);
and U22565 (N_22565,N_18170,N_19669);
and U22566 (N_22566,N_18621,N_18934);
nor U22567 (N_22567,N_19093,N_18532);
xnor U22568 (N_22568,N_18003,N_18912);
nand U22569 (N_22569,N_20478,N_18640);
and U22570 (N_22570,N_20805,N_20559);
and U22571 (N_22571,N_18370,N_19113);
xor U22572 (N_22572,N_18907,N_20367);
or U22573 (N_22573,N_18709,N_20968);
nor U22574 (N_22574,N_18702,N_19142);
nand U22575 (N_22575,N_19570,N_20982);
and U22576 (N_22576,N_19780,N_20823);
and U22577 (N_22577,N_20426,N_20380);
or U22578 (N_22578,N_19968,N_18576);
and U22579 (N_22579,N_20731,N_18177);
and U22580 (N_22580,N_18185,N_19609);
and U22581 (N_22581,N_20992,N_18924);
and U22582 (N_22582,N_20405,N_19807);
nor U22583 (N_22583,N_19135,N_18414);
xor U22584 (N_22584,N_19205,N_18987);
xnor U22585 (N_22585,N_20497,N_20397);
or U22586 (N_22586,N_20062,N_18096);
and U22587 (N_22587,N_18038,N_20424);
xor U22588 (N_22588,N_20336,N_19739);
or U22589 (N_22589,N_19434,N_18838);
or U22590 (N_22590,N_19147,N_20559);
and U22591 (N_22591,N_19401,N_20414);
nor U22592 (N_22592,N_19780,N_19517);
or U22593 (N_22593,N_20040,N_19731);
and U22594 (N_22594,N_18132,N_18328);
nand U22595 (N_22595,N_18232,N_18735);
nand U22596 (N_22596,N_18696,N_20491);
or U22597 (N_22597,N_18447,N_18874);
and U22598 (N_22598,N_20911,N_19823);
and U22599 (N_22599,N_20538,N_20241);
and U22600 (N_22600,N_20617,N_20662);
nand U22601 (N_22601,N_19526,N_19495);
xnor U22602 (N_22602,N_20223,N_20831);
xnor U22603 (N_22603,N_20626,N_20006);
nand U22604 (N_22604,N_18394,N_20083);
and U22605 (N_22605,N_19710,N_20559);
or U22606 (N_22606,N_20847,N_20064);
nand U22607 (N_22607,N_18004,N_20668);
and U22608 (N_22608,N_20655,N_19315);
nand U22609 (N_22609,N_18352,N_19384);
xor U22610 (N_22610,N_18998,N_20712);
nand U22611 (N_22611,N_18486,N_18588);
nor U22612 (N_22612,N_20449,N_18198);
and U22613 (N_22613,N_19039,N_18032);
or U22614 (N_22614,N_19649,N_18872);
and U22615 (N_22615,N_19915,N_20561);
or U22616 (N_22616,N_18998,N_19542);
or U22617 (N_22617,N_20971,N_20390);
or U22618 (N_22618,N_18196,N_19420);
xnor U22619 (N_22619,N_18394,N_19344);
nor U22620 (N_22620,N_20386,N_18372);
and U22621 (N_22621,N_20569,N_18955);
or U22622 (N_22622,N_20912,N_18000);
or U22623 (N_22623,N_19683,N_19749);
or U22624 (N_22624,N_20091,N_20201);
and U22625 (N_22625,N_18579,N_19421);
nor U22626 (N_22626,N_20047,N_20254);
nand U22627 (N_22627,N_20378,N_18626);
nor U22628 (N_22628,N_19968,N_18029);
nand U22629 (N_22629,N_20771,N_19576);
or U22630 (N_22630,N_19289,N_20714);
or U22631 (N_22631,N_18955,N_20884);
or U22632 (N_22632,N_20257,N_20657);
nor U22633 (N_22633,N_18426,N_19132);
and U22634 (N_22634,N_19976,N_19877);
nand U22635 (N_22635,N_18920,N_19782);
nand U22636 (N_22636,N_20937,N_19758);
nand U22637 (N_22637,N_20413,N_18854);
nand U22638 (N_22638,N_20660,N_20631);
or U22639 (N_22639,N_20785,N_19486);
nor U22640 (N_22640,N_19818,N_20097);
and U22641 (N_22641,N_18089,N_18339);
xnor U22642 (N_22642,N_18787,N_18466);
xor U22643 (N_22643,N_20475,N_18708);
and U22644 (N_22644,N_19815,N_18796);
and U22645 (N_22645,N_18883,N_20958);
and U22646 (N_22646,N_20330,N_18630);
or U22647 (N_22647,N_20485,N_18883);
nor U22648 (N_22648,N_19960,N_20438);
nor U22649 (N_22649,N_18752,N_19125);
and U22650 (N_22650,N_20342,N_20903);
nor U22651 (N_22651,N_19468,N_19378);
and U22652 (N_22652,N_19105,N_20485);
nand U22653 (N_22653,N_20756,N_18892);
and U22654 (N_22654,N_19464,N_19847);
nand U22655 (N_22655,N_20794,N_19966);
nand U22656 (N_22656,N_19159,N_19272);
and U22657 (N_22657,N_19428,N_20649);
nor U22658 (N_22658,N_18758,N_18047);
and U22659 (N_22659,N_18392,N_20341);
and U22660 (N_22660,N_20880,N_18947);
nor U22661 (N_22661,N_19502,N_20176);
or U22662 (N_22662,N_18558,N_20277);
nand U22663 (N_22663,N_18237,N_18960);
xnor U22664 (N_22664,N_19690,N_18135);
nor U22665 (N_22665,N_18149,N_20122);
or U22666 (N_22666,N_19425,N_19132);
or U22667 (N_22667,N_18459,N_19713);
and U22668 (N_22668,N_20526,N_20887);
nand U22669 (N_22669,N_18875,N_19480);
nand U22670 (N_22670,N_18723,N_18819);
and U22671 (N_22671,N_18892,N_18623);
and U22672 (N_22672,N_19096,N_19075);
nor U22673 (N_22673,N_20041,N_20726);
or U22674 (N_22674,N_19222,N_20158);
and U22675 (N_22675,N_18547,N_19778);
nand U22676 (N_22676,N_19092,N_18278);
nor U22677 (N_22677,N_20440,N_18091);
xnor U22678 (N_22678,N_20629,N_18665);
nand U22679 (N_22679,N_20896,N_20359);
nand U22680 (N_22680,N_20302,N_20304);
xor U22681 (N_22681,N_19908,N_18187);
nor U22682 (N_22682,N_20648,N_20890);
or U22683 (N_22683,N_20874,N_19462);
nand U22684 (N_22684,N_19618,N_18497);
or U22685 (N_22685,N_19284,N_18822);
nand U22686 (N_22686,N_20537,N_20207);
or U22687 (N_22687,N_18518,N_18154);
nand U22688 (N_22688,N_18571,N_18099);
nand U22689 (N_22689,N_20314,N_19892);
and U22690 (N_22690,N_18652,N_19668);
nor U22691 (N_22691,N_18486,N_20212);
nor U22692 (N_22692,N_19043,N_20395);
nor U22693 (N_22693,N_18563,N_18597);
nor U22694 (N_22694,N_18873,N_20914);
nor U22695 (N_22695,N_19090,N_19538);
and U22696 (N_22696,N_20833,N_20954);
or U22697 (N_22697,N_19116,N_19589);
or U22698 (N_22698,N_20183,N_20786);
xor U22699 (N_22699,N_20491,N_18076);
nor U22700 (N_22700,N_20675,N_18336);
nand U22701 (N_22701,N_20856,N_20689);
nor U22702 (N_22702,N_18944,N_18975);
nand U22703 (N_22703,N_18799,N_19983);
or U22704 (N_22704,N_19856,N_18211);
and U22705 (N_22705,N_20456,N_20695);
nor U22706 (N_22706,N_20505,N_20664);
or U22707 (N_22707,N_19269,N_18062);
or U22708 (N_22708,N_20254,N_20577);
or U22709 (N_22709,N_20725,N_20468);
xnor U22710 (N_22710,N_19324,N_19315);
or U22711 (N_22711,N_18232,N_19861);
nor U22712 (N_22712,N_18356,N_20966);
nand U22713 (N_22713,N_18418,N_20902);
and U22714 (N_22714,N_18575,N_19103);
or U22715 (N_22715,N_20363,N_19762);
and U22716 (N_22716,N_19797,N_18702);
nand U22717 (N_22717,N_20928,N_18283);
nor U22718 (N_22718,N_18172,N_20694);
or U22719 (N_22719,N_18316,N_18444);
and U22720 (N_22720,N_18573,N_20834);
nand U22721 (N_22721,N_18730,N_19309);
nor U22722 (N_22722,N_20437,N_19900);
nand U22723 (N_22723,N_19492,N_20046);
nand U22724 (N_22724,N_18461,N_20734);
nand U22725 (N_22725,N_18356,N_18327);
and U22726 (N_22726,N_18466,N_18919);
nand U22727 (N_22727,N_19517,N_18556);
or U22728 (N_22728,N_19951,N_20783);
and U22729 (N_22729,N_20246,N_19193);
nor U22730 (N_22730,N_20908,N_18803);
nand U22731 (N_22731,N_19671,N_18024);
and U22732 (N_22732,N_20188,N_18389);
nand U22733 (N_22733,N_18778,N_19310);
and U22734 (N_22734,N_18234,N_18503);
nand U22735 (N_22735,N_20226,N_20383);
or U22736 (N_22736,N_18978,N_19531);
nand U22737 (N_22737,N_18929,N_20417);
nor U22738 (N_22738,N_20561,N_20680);
nor U22739 (N_22739,N_18479,N_19122);
or U22740 (N_22740,N_19996,N_20055);
nand U22741 (N_22741,N_20153,N_19269);
nand U22742 (N_22742,N_20108,N_20891);
and U22743 (N_22743,N_19462,N_20731);
xnor U22744 (N_22744,N_19334,N_19736);
or U22745 (N_22745,N_19500,N_19283);
or U22746 (N_22746,N_20782,N_19676);
nand U22747 (N_22747,N_20886,N_18928);
nor U22748 (N_22748,N_18626,N_18733);
nor U22749 (N_22749,N_18311,N_19244);
nand U22750 (N_22750,N_19458,N_20579);
or U22751 (N_22751,N_20684,N_19248);
nand U22752 (N_22752,N_19169,N_19161);
and U22753 (N_22753,N_20422,N_18041);
nand U22754 (N_22754,N_18893,N_20719);
and U22755 (N_22755,N_19796,N_20805);
or U22756 (N_22756,N_20396,N_19409);
nand U22757 (N_22757,N_19523,N_19317);
xor U22758 (N_22758,N_18628,N_18522);
nand U22759 (N_22759,N_20449,N_19405);
and U22760 (N_22760,N_19636,N_18378);
or U22761 (N_22761,N_18729,N_20739);
nor U22762 (N_22762,N_18739,N_18705);
or U22763 (N_22763,N_18826,N_18010);
and U22764 (N_22764,N_19942,N_19039);
or U22765 (N_22765,N_19774,N_19310);
or U22766 (N_22766,N_20640,N_20884);
nor U22767 (N_22767,N_20775,N_18953);
xor U22768 (N_22768,N_20609,N_20814);
xnor U22769 (N_22769,N_18327,N_18183);
nor U22770 (N_22770,N_18780,N_18129);
and U22771 (N_22771,N_18998,N_19389);
or U22772 (N_22772,N_20100,N_18240);
nand U22773 (N_22773,N_19861,N_19939);
nand U22774 (N_22774,N_19174,N_18337);
nand U22775 (N_22775,N_19854,N_20850);
and U22776 (N_22776,N_20599,N_19459);
nor U22777 (N_22777,N_20421,N_19381);
nand U22778 (N_22778,N_19967,N_18379);
or U22779 (N_22779,N_18102,N_20034);
nand U22780 (N_22780,N_19433,N_19021);
or U22781 (N_22781,N_19908,N_18984);
nor U22782 (N_22782,N_18656,N_18754);
and U22783 (N_22783,N_18694,N_18445);
nor U22784 (N_22784,N_20698,N_20562);
nand U22785 (N_22785,N_20817,N_18164);
and U22786 (N_22786,N_19730,N_20129);
nor U22787 (N_22787,N_19179,N_19723);
nor U22788 (N_22788,N_19218,N_19878);
nor U22789 (N_22789,N_18995,N_20651);
and U22790 (N_22790,N_18530,N_20134);
and U22791 (N_22791,N_19978,N_18842);
nand U22792 (N_22792,N_19342,N_18041);
and U22793 (N_22793,N_18920,N_19168);
nor U22794 (N_22794,N_18468,N_18408);
or U22795 (N_22795,N_20123,N_19417);
nand U22796 (N_22796,N_19762,N_19514);
nor U22797 (N_22797,N_20392,N_20014);
nor U22798 (N_22798,N_19039,N_19485);
nand U22799 (N_22799,N_19008,N_20664);
and U22800 (N_22800,N_20323,N_19203);
and U22801 (N_22801,N_20264,N_20689);
nor U22802 (N_22802,N_19441,N_19891);
nor U22803 (N_22803,N_19184,N_19460);
and U22804 (N_22804,N_19397,N_18668);
nand U22805 (N_22805,N_19607,N_18147);
or U22806 (N_22806,N_18028,N_20322);
and U22807 (N_22807,N_18991,N_19006);
and U22808 (N_22808,N_18729,N_18809);
or U22809 (N_22809,N_19886,N_19603);
xor U22810 (N_22810,N_18148,N_20850);
and U22811 (N_22811,N_20935,N_19208);
and U22812 (N_22812,N_18580,N_19193);
and U22813 (N_22813,N_19020,N_18490);
or U22814 (N_22814,N_20139,N_20557);
nand U22815 (N_22815,N_19091,N_19559);
and U22816 (N_22816,N_20396,N_20222);
and U22817 (N_22817,N_18367,N_20962);
and U22818 (N_22818,N_20306,N_20499);
nor U22819 (N_22819,N_19052,N_18819);
nor U22820 (N_22820,N_20759,N_20139);
or U22821 (N_22821,N_18840,N_18060);
or U22822 (N_22822,N_18531,N_18437);
xnor U22823 (N_22823,N_19017,N_20456);
xnor U22824 (N_22824,N_18566,N_18923);
nand U22825 (N_22825,N_20864,N_18819);
nand U22826 (N_22826,N_18562,N_20599);
nand U22827 (N_22827,N_18446,N_20033);
nor U22828 (N_22828,N_18836,N_18637);
and U22829 (N_22829,N_18656,N_18611);
and U22830 (N_22830,N_19576,N_20433);
nand U22831 (N_22831,N_20623,N_20967);
xor U22832 (N_22832,N_19513,N_18540);
and U22833 (N_22833,N_18042,N_18681);
and U22834 (N_22834,N_19234,N_20219);
nor U22835 (N_22835,N_19256,N_18152);
and U22836 (N_22836,N_19478,N_19513);
nand U22837 (N_22837,N_19925,N_20305);
nand U22838 (N_22838,N_18163,N_18417);
nand U22839 (N_22839,N_19132,N_20783);
and U22840 (N_22840,N_19536,N_18548);
or U22841 (N_22841,N_19947,N_20944);
nor U22842 (N_22842,N_18855,N_18413);
nand U22843 (N_22843,N_18430,N_19387);
and U22844 (N_22844,N_20714,N_20017);
nand U22845 (N_22845,N_18027,N_18412);
or U22846 (N_22846,N_19739,N_18920);
nand U22847 (N_22847,N_20713,N_18637);
and U22848 (N_22848,N_19013,N_18878);
or U22849 (N_22849,N_20378,N_20925);
and U22850 (N_22850,N_19937,N_19917);
nor U22851 (N_22851,N_18952,N_19703);
or U22852 (N_22852,N_20168,N_18151);
or U22853 (N_22853,N_18462,N_19112);
nand U22854 (N_22854,N_18177,N_19220);
nor U22855 (N_22855,N_20730,N_20245);
and U22856 (N_22856,N_20146,N_18648);
nor U22857 (N_22857,N_18752,N_18726);
and U22858 (N_22858,N_18831,N_19416);
and U22859 (N_22859,N_18172,N_19603);
xnor U22860 (N_22860,N_20761,N_19241);
and U22861 (N_22861,N_20931,N_20057);
xor U22862 (N_22862,N_20230,N_19864);
nor U22863 (N_22863,N_19604,N_19035);
nand U22864 (N_22864,N_19825,N_19305);
nand U22865 (N_22865,N_18733,N_19747);
nand U22866 (N_22866,N_20937,N_18170);
or U22867 (N_22867,N_20931,N_19594);
and U22868 (N_22868,N_19451,N_18086);
xor U22869 (N_22869,N_19090,N_20870);
or U22870 (N_22870,N_18532,N_19151);
or U22871 (N_22871,N_19091,N_18314);
and U22872 (N_22872,N_19378,N_20794);
and U22873 (N_22873,N_20221,N_19328);
nor U22874 (N_22874,N_20229,N_20241);
nand U22875 (N_22875,N_19386,N_20820);
or U22876 (N_22876,N_19963,N_19201);
and U22877 (N_22877,N_20909,N_18840);
and U22878 (N_22878,N_20790,N_20518);
or U22879 (N_22879,N_18768,N_19274);
and U22880 (N_22880,N_18150,N_18067);
and U22881 (N_22881,N_19820,N_20523);
xnor U22882 (N_22882,N_19387,N_20510);
xor U22883 (N_22883,N_19277,N_19270);
xor U22884 (N_22884,N_20882,N_19224);
nor U22885 (N_22885,N_18215,N_20778);
or U22886 (N_22886,N_19433,N_18371);
nor U22887 (N_22887,N_19508,N_20330);
and U22888 (N_22888,N_19724,N_18888);
and U22889 (N_22889,N_19631,N_19161);
nand U22890 (N_22890,N_18278,N_18661);
nor U22891 (N_22891,N_18538,N_20542);
nor U22892 (N_22892,N_20079,N_18557);
xnor U22893 (N_22893,N_20248,N_19263);
nand U22894 (N_22894,N_19531,N_18671);
xnor U22895 (N_22895,N_20071,N_19932);
and U22896 (N_22896,N_19222,N_20092);
nand U22897 (N_22897,N_19524,N_19623);
or U22898 (N_22898,N_19567,N_19345);
xor U22899 (N_22899,N_20769,N_20638);
nand U22900 (N_22900,N_20253,N_20915);
or U22901 (N_22901,N_20779,N_18791);
nor U22902 (N_22902,N_19842,N_19252);
xnor U22903 (N_22903,N_20856,N_19505);
nand U22904 (N_22904,N_20881,N_19856);
nand U22905 (N_22905,N_18633,N_19207);
nor U22906 (N_22906,N_20102,N_20979);
or U22907 (N_22907,N_19939,N_18189);
nor U22908 (N_22908,N_19970,N_18884);
nor U22909 (N_22909,N_20538,N_18007);
nor U22910 (N_22910,N_20075,N_20043);
nand U22911 (N_22911,N_20210,N_19446);
xnor U22912 (N_22912,N_18251,N_20923);
or U22913 (N_22913,N_19392,N_18168);
nor U22914 (N_22914,N_19749,N_18633);
nor U22915 (N_22915,N_18108,N_19816);
nor U22916 (N_22916,N_20852,N_20426);
or U22917 (N_22917,N_20640,N_19361);
and U22918 (N_22918,N_20087,N_20652);
nor U22919 (N_22919,N_19946,N_18247);
and U22920 (N_22920,N_18670,N_18045);
or U22921 (N_22921,N_20233,N_18413);
xnor U22922 (N_22922,N_20767,N_19144);
or U22923 (N_22923,N_19221,N_20340);
nor U22924 (N_22924,N_18771,N_18859);
xnor U22925 (N_22925,N_18191,N_20165);
nor U22926 (N_22926,N_19230,N_19862);
nand U22927 (N_22927,N_18476,N_20378);
or U22928 (N_22928,N_20502,N_20264);
or U22929 (N_22929,N_18580,N_18044);
xnor U22930 (N_22930,N_19943,N_20742);
or U22931 (N_22931,N_18333,N_18520);
nand U22932 (N_22932,N_18125,N_20389);
and U22933 (N_22933,N_20882,N_19906);
and U22934 (N_22934,N_19471,N_19127);
and U22935 (N_22935,N_19285,N_18860);
nand U22936 (N_22936,N_20012,N_18172);
and U22937 (N_22937,N_20802,N_18798);
xor U22938 (N_22938,N_19995,N_20638);
or U22939 (N_22939,N_18502,N_18867);
xnor U22940 (N_22940,N_18178,N_18547);
nand U22941 (N_22941,N_19838,N_20144);
or U22942 (N_22942,N_18024,N_18734);
nand U22943 (N_22943,N_19020,N_20036);
nand U22944 (N_22944,N_18590,N_18546);
nor U22945 (N_22945,N_18519,N_20622);
and U22946 (N_22946,N_19385,N_19709);
and U22947 (N_22947,N_20064,N_19732);
xor U22948 (N_22948,N_19951,N_19164);
and U22949 (N_22949,N_20799,N_20411);
nor U22950 (N_22950,N_20513,N_18575);
nand U22951 (N_22951,N_20984,N_18353);
nand U22952 (N_22952,N_18503,N_18428);
nor U22953 (N_22953,N_18313,N_20497);
nand U22954 (N_22954,N_20350,N_19521);
nor U22955 (N_22955,N_18260,N_19070);
nand U22956 (N_22956,N_20775,N_18072);
xor U22957 (N_22957,N_18309,N_18099);
or U22958 (N_22958,N_20480,N_20761);
xnor U22959 (N_22959,N_20712,N_20951);
and U22960 (N_22960,N_20217,N_19300);
nand U22961 (N_22961,N_19457,N_19682);
and U22962 (N_22962,N_18898,N_19314);
and U22963 (N_22963,N_20013,N_20945);
xor U22964 (N_22964,N_19094,N_19705);
or U22965 (N_22965,N_18376,N_19912);
or U22966 (N_22966,N_20978,N_19671);
nand U22967 (N_22967,N_20656,N_20692);
nor U22968 (N_22968,N_19849,N_19003);
xor U22969 (N_22969,N_19679,N_19939);
and U22970 (N_22970,N_20627,N_18090);
and U22971 (N_22971,N_19426,N_18912);
and U22972 (N_22972,N_20509,N_19560);
xor U22973 (N_22973,N_18970,N_20362);
nor U22974 (N_22974,N_20370,N_18809);
xor U22975 (N_22975,N_19114,N_20617);
xnor U22976 (N_22976,N_19759,N_20892);
and U22977 (N_22977,N_20723,N_18699);
or U22978 (N_22978,N_19862,N_18262);
and U22979 (N_22979,N_18936,N_19674);
xnor U22980 (N_22980,N_19172,N_18455);
nand U22981 (N_22981,N_20714,N_20013);
or U22982 (N_22982,N_19363,N_18661);
or U22983 (N_22983,N_20147,N_19315);
or U22984 (N_22984,N_20024,N_18430);
nand U22985 (N_22985,N_19598,N_20844);
nor U22986 (N_22986,N_20353,N_20330);
or U22987 (N_22987,N_20252,N_20418);
nand U22988 (N_22988,N_19412,N_18822);
or U22989 (N_22989,N_19613,N_20828);
or U22990 (N_22990,N_20266,N_20002);
nor U22991 (N_22991,N_20760,N_20493);
or U22992 (N_22992,N_18907,N_20934);
nand U22993 (N_22993,N_18951,N_18373);
and U22994 (N_22994,N_20892,N_18416);
and U22995 (N_22995,N_18625,N_20115);
or U22996 (N_22996,N_19212,N_19416);
nand U22997 (N_22997,N_19252,N_20773);
and U22998 (N_22998,N_18808,N_20327);
xor U22999 (N_22999,N_18280,N_20507);
nor U23000 (N_23000,N_19694,N_20971);
or U23001 (N_23001,N_19650,N_18893);
and U23002 (N_23002,N_20562,N_19087);
nand U23003 (N_23003,N_18862,N_20237);
and U23004 (N_23004,N_20654,N_18173);
nand U23005 (N_23005,N_20689,N_19646);
or U23006 (N_23006,N_18430,N_20585);
and U23007 (N_23007,N_19740,N_20141);
xor U23008 (N_23008,N_18879,N_20555);
nor U23009 (N_23009,N_19461,N_20198);
nor U23010 (N_23010,N_18764,N_18892);
or U23011 (N_23011,N_19424,N_19866);
nand U23012 (N_23012,N_20784,N_18375);
nor U23013 (N_23013,N_20343,N_20280);
nor U23014 (N_23014,N_19866,N_18787);
nand U23015 (N_23015,N_19127,N_18460);
and U23016 (N_23016,N_19334,N_19824);
and U23017 (N_23017,N_18240,N_19733);
and U23018 (N_23018,N_20176,N_20320);
and U23019 (N_23019,N_19073,N_19659);
nand U23020 (N_23020,N_19539,N_19803);
and U23021 (N_23021,N_19452,N_19207);
or U23022 (N_23022,N_20140,N_20409);
and U23023 (N_23023,N_19799,N_20679);
nor U23024 (N_23024,N_20038,N_19728);
or U23025 (N_23025,N_19887,N_20538);
nand U23026 (N_23026,N_19110,N_20156);
xnor U23027 (N_23027,N_19569,N_20031);
or U23028 (N_23028,N_18806,N_19844);
nor U23029 (N_23029,N_19166,N_18847);
or U23030 (N_23030,N_20507,N_20063);
nand U23031 (N_23031,N_20101,N_19404);
xor U23032 (N_23032,N_19406,N_19802);
or U23033 (N_23033,N_20900,N_20179);
xor U23034 (N_23034,N_18469,N_18435);
or U23035 (N_23035,N_18351,N_19917);
nand U23036 (N_23036,N_18591,N_20642);
nor U23037 (N_23037,N_18902,N_20229);
and U23038 (N_23038,N_19261,N_18140);
nand U23039 (N_23039,N_19099,N_20366);
and U23040 (N_23040,N_19229,N_18616);
nand U23041 (N_23041,N_19157,N_19959);
or U23042 (N_23042,N_19299,N_19611);
or U23043 (N_23043,N_19847,N_20019);
or U23044 (N_23044,N_18784,N_18546);
nor U23045 (N_23045,N_20923,N_20379);
and U23046 (N_23046,N_19538,N_18138);
nor U23047 (N_23047,N_20680,N_19619);
nor U23048 (N_23048,N_20573,N_19421);
nor U23049 (N_23049,N_20333,N_19125);
xnor U23050 (N_23050,N_19753,N_19543);
nor U23051 (N_23051,N_20810,N_20726);
nand U23052 (N_23052,N_20945,N_19083);
and U23053 (N_23053,N_19864,N_20575);
nand U23054 (N_23054,N_18527,N_19786);
nand U23055 (N_23055,N_18164,N_20288);
xnor U23056 (N_23056,N_20975,N_18899);
xnor U23057 (N_23057,N_20050,N_19664);
nand U23058 (N_23058,N_19903,N_20622);
or U23059 (N_23059,N_20587,N_18625);
and U23060 (N_23060,N_18140,N_19335);
nor U23061 (N_23061,N_18003,N_18590);
or U23062 (N_23062,N_19386,N_20938);
nand U23063 (N_23063,N_19162,N_20096);
nor U23064 (N_23064,N_20836,N_18810);
nand U23065 (N_23065,N_20318,N_18673);
nand U23066 (N_23066,N_18401,N_19600);
nor U23067 (N_23067,N_20200,N_19279);
nand U23068 (N_23068,N_20189,N_18424);
nor U23069 (N_23069,N_19096,N_18322);
or U23070 (N_23070,N_20325,N_20563);
xor U23071 (N_23071,N_18004,N_18608);
and U23072 (N_23072,N_20938,N_19471);
nand U23073 (N_23073,N_20203,N_19939);
or U23074 (N_23074,N_20110,N_18127);
or U23075 (N_23075,N_19308,N_18317);
nor U23076 (N_23076,N_19607,N_20077);
and U23077 (N_23077,N_18130,N_18281);
and U23078 (N_23078,N_19650,N_19221);
xnor U23079 (N_23079,N_19286,N_20957);
and U23080 (N_23080,N_20022,N_18671);
and U23081 (N_23081,N_19528,N_19466);
or U23082 (N_23082,N_19466,N_20008);
nand U23083 (N_23083,N_19714,N_18244);
xor U23084 (N_23084,N_18441,N_18912);
nor U23085 (N_23085,N_18849,N_19629);
or U23086 (N_23086,N_19131,N_18037);
or U23087 (N_23087,N_19898,N_20649);
nor U23088 (N_23088,N_18269,N_19407);
nor U23089 (N_23089,N_18457,N_19039);
xnor U23090 (N_23090,N_18884,N_18163);
nand U23091 (N_23091,N_20494,N_20105);
and U23092 (N_23092,N_18080,N_19601);
nand U23093 (N_23093,N_18183,N_19668);
nand U23094 (N_23094,N_19639,N_18383);
nand U23095 (N_23095,N_18003,N_19108);
nand U23096 (N_23096,N_18972,N_18822);
nor U23097 (N_23097,N_19373,N_19831);
or U23098 (N_23098,N_19244,N_19823);
nand U23099 (N_23099,N_19954,N_18867);
or U23100 (N_23100,N_18978,N_18033);
or U23101 (N_23101,N_20031,N_18881);
nand U23102 (N_23102,N_18963,N_18827);
and U23103 (N_23103,N_19998,N_18922);
nor U23104 (N_23104,N_19885,N_18338);
or U23105 (N_23105,N_18351,N_20305);
xnor U23106 (N_23106,N_19516,N_20590);
nor U23107 (N_23107,N_19929,N_19103);
nor U23108 (N_23108,N_20201,N_19707);
xor U23109 (N_23109,N_18978,N_20445);
nand U23110 (N_23110,N_20495,N_20058);
xor U23111 (N_23111,N_18478,N_19999);
or U23112 (N_23112,N_18905,N_20612);
xnor U23113 (N_23113,N_20885,N_20437);
or U23114 (N_23114,N_19097,N_19386);
nand U23115 (N_23115,N_18367,N_20131);
or U23116 (N_23116,N_20396,N_18878);
or U23117 (N_23117,N_19605,N_18801);
nand U23118 (N_23118,N_18197,N_18146);
or U23119 (N_23119,N_18616,N_19300);
nor U23120 (N_23120,N_18848,N_19684);
nor U23121 (N_23121,N_20236,N_19457);
and U23122 (N_23122,N_18824,N_20956);
or U23123 (N_23123,N_20863,N_18187);
and U23124 (N_23124,N_19499,N_19379);
nand U23125 (N_23125,N_18645,N_19015);
nand U23126 (N_23126,N_20065,N_19251);
and U23127 (N_23127,N_19692,N_20976);
xor U23128 (N_23128,N_19594,N_19591);
xnor U23129 (N_23129,N_19749,N_19129);
or U23130 (N_23130,N_20198,N_20016);
and U23131 (N_23131,N_19174,N_18062);
or U23132 (N_23132,N_18548,N_18786);
nand U23133 (N_23133,N_18986,N_18873);
nor U23134 (N_23134,N_19313,N_19678);
and U23135 (N_23135,N_18695,N_18478);
and U23136 (N_23136,N_18189,N_18547);
xor U23137 (N_23137,N_20003,N_20804);
and U23138 (N_23138,N_20536,N_18593);
nand U23139 (N_23139,N_19581,N_19516);
and U23140 (N_23140,N_20121,N_18247);
nand U23141 (N_23141,N_20900,N_20167);
nand U23142 (N_23142,N_20849,N_18051);
nor U23143 (N_23143,N_20709,N_19660);
nand U23144 (N_23144,N_20659,N_20777);
xnor U23145 (N_23145,N_20440,N_18446);
nand U23146 (N_23146,N_19547,N_18898);
nor U23147 (N_23147,N_18648,N_20003);
nand U23148 (N_23148,N_18390,N_19095);
nor U23149 (N_23149,N_19149,N_18880);
and U23150 (N_23150,N_19933,N_20295);
nor U23151 (N_23151,N_19573,N_18860);
nand U23152 (N_23152,N_20862,N_18771);
or U23153 (N_23153,N_20242,N_19836);
nand U23154 (N_23154,N_19476,N_20737);
or U23155 (N_23155,N_18501,N_19476);
and U23156 (N_23156,N_19998,N_18502);
nand U23157 (N_23157,N_19059,N_19728);
xnor U23158 (N_23158,N_19106,N_18823);
nand U23159 (N_23159,N_18438,N_19969);
or U23160 (N_23160,N_18993,N_18021);
and U23161 (N_23161,N_20178,N_18208);
nand U23162 (N_23162,N_19883,N_19678);
and U23163 (N_23163,N_20995,N_19708);
and U23164 (N_23164,N_20601,N_18771);
nand U23165 (N_23165,N_18953,N_18488);
nand U23166 (N_23166,N_18321,N_18780);
and U23167 (N_23167,N_19701,N_19521);
and U23168 (N_23168,N_18080,N_20846);
or U23169 (N_23169,N_19617,N_19140);
or U23170 (N_23170,N_18071,N_20207);
nand U23171 (N_23171,N_19399,N_20464);
and U23172 (N_23172,N_19966,N_18178);
nand U23173 (N_23173,N_18632,N_20660);
and U23174 (N_23174,N_19428,N_19148);
nand U23175 (N_23175,N_20802,N_19444);
and U23176 (N_23176,N_19908,N_19332);
nand U23177 (N_23177,N_18067,N_20714);
xor U23178 (N_23178,N_18025,N_19014);
or U23179 (N_23179,N_19032,N_20143);
nor U23180 (N_23180,N_20361,N_19395);
and U23181 (N_23181,N_19314,N_18793);
or U23182 (N_23182,N_20843,N_19890);
nor U23183 (N_23183,N_20334,N_20538);
nor U23184 (N_23184,N_20560,N_18029);
nor U23185 (N_23185,N_20270,N_19921);
xor U23186 (N_23186,N_19774,N_18248);
nand U23187 (N_23187,N_20650,N_20679);
xnor U23188 (N_23188,N_19599,N_19973);
nand U23189 (N_23189,N_18692,N_20951);
or U23190 (N_23190,N_19855,N_18091);
nand U23191 (N_23191,N_20833,N_19298);
nand U23192 (N_23192,N_19908,N_18295);
or U23193 (N_23193,N_20586,N_19394);
nand U23194 (N_23194,N_19704,N_18817);
and U23195 (N_23195,N_18222,N_19717);
nor U23196 (N_23196,N_19599,N_20337);
nor U23197 (N_23197,N_19701,N_20581);
nand U23198 (N_23198,N_18288,N_19445);
or U23199 (N_23199,N_18106,N_20950);
or U23200 (N_23200,N_20081,N_19253);
nor U23201 (N_23201,N_18878,N_18072);
nand U23202 (N_23202,N_18845,N_18318);
and U23203 (N_23203,N_18277,N_20421);
nand U23204 (N_23204,N_18692,N_20734);
nor U23205 (N_23205,N_20960,N_20731);
and U23206 (N_23206,N_19977,N_18528);
or U23207 (N_23207,N_19215,N_19964);
or U23208 (N_23208,N_20646,N_18178);
or U23209 (N_23209,N_19394,N_20792);
nor U23210 (N_23210,N_20719,N_19509);
nand U23211 (N_23211,N_20474,N_20030);
nand U23212 (N_23212,N_19415,N_19160);
and U23213 (N_23213,N_19874,N_19512);
and U23214 (N_23214,N_18660,N_20472);
nor U23215 (N_23215,N_20472,N_19726);
and U23216 (N_23216,N_20257,N_20550);
nor U23217 (N_23217,N_18962,N_19722);
nand U23218 (N_23218,N_18753,N_19081);
and U23219 (N_23219,N_20334,N_18019);
nand U23220 (N_23220,N_20552,N_18047);
and U23221 (N_23221,N_18400,N_20750);
or U23222 (N_23222,N_18448,N_18113);
nand U23223 (N_23223,N_19790,N_19386);
nor U23224 (N_23224,N_20731,N_18089);
nand U23225 (N_23225,N_20035,N_19110);
or U23226 (N_23226,N_19245,N_20250);
and U23227 (N_23227,N_19250,N_18302);
or U23228 (N_23228,N_20366,N_18990);
nor U23229 (N_23229,N_20136,N_19781);
nor U23230 (N_23230,N_18710,N_18415);
nor U23231 (N_23231,N_18330,N_19961);
nor U23232 (N_23232,N_20855,N_18704);
or U23233 (N_23233,N_19985,N_18252);
xnor U23234 (N_23234,N_20670,N_19496);
nand U23235 (N_23235,N_18991,N_20436);
nor U23236 (N_23236,N_19967,N_20209);
or U23237 (N_23237,N_18443,N_20633);
and U23238 (N_23238,N_19977,N_20782);
and U23239 (N_23239,N_20696,N_20652);
and U23240 (N_23240,N_19595,N_18428);
or U23241 (N_23241,N_19490,N_20588);
nand U23242 (N_23242,N_20193,N_18922);
nand U23243 (N_23243,N_19314,N_18031);
xor U23244 (N_23244,N_20996,N_19128);
or U23245 (N_23245,N_19023,N_19718);
and U23246 (N_23246,N_18787,N_19730);
xor U23247 (N_23247,N_20167,N_19846);
nor U23248 (N_23248,N_19823,N_20315);
nor U23249 (N_23249,N_20964,N_18209);
nor U23250 (N_23250,N_18971,N_19415);
xnor U23251 (N_23251,N_19131,N_18998);
nor U23252 (N_23252,N_20030,N_19918);
nand U23253 (N_23253,N_19782,N_19231);
xor U23254 (N_23254,N_20282,N_20237);
nor U23255 (N_23255,N_19866,N_18758);
nor U23256 (N_23256,N_19449,N_19225);
xnor U23257 (N_23257,N_19200,N_18042);
and U23258 (N_23258,N_20280,N_19431);
nand U23259 (N_23259,N_20880,N_18107);
nand U23260 (N_23260,N_19667,N_18781);
nor U23261 (N_23261,N_19596,N_19018);
nand U23262 (N_23262,N_19527,N_19305);
xnor U23263 (N_23263,N_18171,N_19475);
or U23264 (N_23264,N_20424,N_20040);
xnor U23265 (N_23265,N_18283,N_18637);
and U23266 (N_23266,N_20834,N_18003);
nand U23267 (N_23267,N_19507,N_18183);
or U23268 (N_23268,N_18627,N_20707);
nor U23269 (N_23269,N_20318,N_19075);
or U23270 (N_23270,N_18360,N_20455);
nand U23271 (N_23271,N_20471,N_20787);
nor U23272 (N_23272,N_19471,N_20195);
xor U23273 (N_23273,N_20463,N_18892);
or U23274 (N_23274,N_20392,N_19373);
nand U23275 (N_23275,N_18653,N_18120);
nand U23276 (N_23276,N_20873,N_19468);
nand U23277 (N_23277,N_20166,N_18952);
or U23278 (N_23278,N_19274,N_19534);
xnor U23279 (N_23279,N_18012,N_19052);
nand U23280 (N_23280,N_20274,N_20233);
xor U23281 (N_23281,N_20205,N_20440);
nor U23282 (N_23282,N_20987,N_19772);
or U23283 (N_23283,N_18043,N_19386);
xor U23284 (N_23284,N_19403,N_20452);
nor U23285 (N_23285,N_20467,N_20648);
nand U23286 (N_23286,N_18432,N_20343);
nand U23287 (N_23287,N_20644,N_18494);
or U23288 (N_23288,N_19103,N_19557);
nor U23289 (N_23289,N_20689,N_19837);
nor U23290 (N_23290,N_20446,N_20633);
and U23291 (N_23291,N_20875,N_19684);
nand U23292 (N_23292,N_18606,N_19778);
nand U23293 (N_23293,N_19744,N_20782);
and U23294 (N_23294,N_18610,N_19099);
nand U23295 (N_23295,N_18148,N_19491);
nand U23296 (N_23296,N_18110,N_18117);
and U23297 (N_23297,N_19771,N_20905);
or U23298 (N_23298,N_18283,N_18406);
nor U23299 (N_23299,N_18771,N_18388);
nor U23300 (N_23300,N_19083,N_18221);
and U23301 (N_23301,N_18312,N_20433);
nor U23302 (N_23302,N_18698,N_18183);
xor U23303 (N_23303,N_18271,N_19687);
nand U23304 (N_23304,N_19856,N_19253);
nand U23305 (N_23305,N_20820,N_18952);
nor U23306 (N_23306,N_18575,N_18677);
xnor U23307 (N_23307,N_20158,N_20753);
nand U23308 (N_23308,N_18833,N_18683);
nand U23309 (N_23309,N_19814,N_18089);
nand U23310 (N_23310,N_20453,N_18575);
or U23311 (N_23311,N_19127,N_20507);
and U23312 (N_23312,N_18620,N_18339);
nand U23313 (N_23313,N_18767,N_20584);
nand U23314 (N_23314,N_19952,N_18463);
xnor U23315 (N_23315,N_18883,N_18298);
nor U23316 (N_23316,N_18278,N_20917);
nand U23317 (N_23317,N_20413,N_19755);
nor U23318 (N_23318,N_20865,N_20977);
and U23319 (N_23319,N_19672,N_18054);
and U23320 (N_23320,N_19222,N_18128);
xnor U23321 (N_23321,N_18660,N_20140);
and U23322 (N_23322,N_19929,N_20307);
xor U23323 (N_23323,N_19854,N_19830);
and U23324 (N_23324,N_20444,N_19908);
nand U23325 (N_23325,N_18502,N_20642);
and U23326 (N_23326,N_20515,N_19514);
or U23327 (N_23327,N_19365,N_19680);
nor U23328 (N_23328,N_18510,N_19893);
nand U23329 (N_23329,N_20046,N_19665);
nor U23330 (N_23330,N_20489,N_20687);
xor U23331 (N_23331,N_19236,N_18988);
or U23332 (N_23332,N_20480,N_18937);
and U23333 (N_23333,N_19606,N_20320);
nand U23334 (N_23334,N_20713,N_19369);
nand U23335 (N_23335,N_20220,N_18090);
nor U23336 (N_23336,N_19410,N_18221);
nor U23337 (N_23337,N_18124,N_18277);
nand U23338 (N_23338,N_19207,N_20659);
or U23339 (N_23339,N_20894,N_20767);
nand U23340 (N_23340,N_19072,N_19195);
and U23341 (N_23341,N_20420,N_19029);
or U23342 (N_23342,N_20051,N_18944);
or U23343 (N_23343,N_19128,N_18336);
nor U23344 (N_23344,N_18440,N_20937);
nand U23345 (N_23345,N_19059,N_19003);
nor U23346 (N_23346,N_19825,N_20052);
nor U23347 (N_23347,N_18415,N_18377);
xor U23348 (N_23348,N_19155,N_20823);
and U23349 (N_23349,N_18690,N_19940);
or U23350 (N_23350,N_20621,N_18923);
and U23351 (N_23351,N_20699,N_18994);
nand U23352 (N_23352,N_20706,N_20943);
nand U23353 (N_23353,N_18810,N_20852);
nor U23354 (N_23354,N_19373,N_19457);
nand U23355 (N_23355,N_19866,N_19659);
nor U23356 (N_23356,N_18214,N_20439);
or U23357 (N_23357,N_19162,N_18769);
and U23358 (N_23358,N_18864,N_20779);
and U23359 (N_23359,N_18670,N_18217);
nand U23360 (N_23360,N_19636,N_20856);
or U23361 (N_23361,N_18371,N_19421);
and U23362 (N_23362,N_18798,N_18227);
xor U23363 (N_23363,N_20888,N_20651);
xnor U23364 (N_23364,N_19319,N_19379);
nand U23365 (N_23365,N_18404,N_20163);
nand U23366 (N_23366,N_18224,N_20692);
and U23367 (N_23367,N_20712,N_18010);
nand U23368 (N_23368,N_19943,N_18548);
nand U23369 (N_23369,N_20710,N_18310);
nor U23370 (N_23370,N_19049,N_20688);
or U23371 (N_23371,N_19555,N_19286);
or U23372 (N_23372,N_20408,N_19131);
nand U23373 (N_23373,N_18784,N_18833);
and U23374 (N_23374,N_18249,N_18575);
nand U23375 (N_23375,N_19968,N_19979);
xnor U23376 (N_23376,N_19130,N_20565);
nand U23377 (N_23377,N_18096,N_19623);
or U23378 (N_23378,N_20919,N_19682);
nand U23379 (N_23379,N_19882,N_18106);
or U23380 (N_23380,N_18601,N_20149);
nand U23381 (N_23381,N_18862,N_20039);
nor U23382 (N_23382,N_18439,N_19889);
nand U23383 (N_23383,N_18790,N_20766);
nand U23384 (N_23384,N_20835,N_20073);
and U23385 (N_23385,N_18420,N_18377);
and U23386 (N_23386,N_18472,N_20987);
nor U23387 (N_23387,N_18115,N_20826);
and U23388 (N_23388,N_18370,N_20807);
nand U23389 (N_23389,N_18969,N_19514);
or U23390 (N_23390,N_18665,N_19809);
or U23391 (N_23391,N_19274,N_20763);
nor U23392 (N_23392,N_18056,N_18778);
or U23393 (N_23393,N_19971,N_19287);
nor U23394 (N_23394,N_19074,N_18023);
nor U23395 (N_23395,N_18229,N_18027);
xor U23396 (N_23396,N_19946,N_19511);
or U23397 (N_23397,N_18292,N_19707);
or U23398 (N_23398,N_18489,N_20039);
nand U23399 (N_23399,N_19537,N_20555);
or U23400 (N_23400,N_20710,N_18250);
nand U23401 (N_23401,N_20125,N_18190);
nand U23402 (N_23402,N_19347,N_19436);
and U23403 (N_23403,N_18352,N_19823);
nor U23404 (N_23404,N_20542,N_19951);
nor U23405 (N_23405,N_20080,N_18917);
nor U23406 (N_23406,N_18453,N_20854);
xor U23407 (N_23407,N_18560,N_20189);
or U23408 (N_23408,N_20452,N_18803);
or U23409 (N_23409,N_19732,N_19531);
nand U23410 (N_23410,N_18713,N_19282);
xor U23411 (N_23411,N_18355,N_20699);
xnor U23412 (N_23412,N_18706,N_19263);
nor U23413 (N_23413,N_20311,N_20259);
and U23414 (N_23414,N_19537,N_18181);
nand U23415 (N_23415,N_18211,N_18711);
nand U23416 (N_23416,N_19307,N_19510);
xor U23417 (N_23417,N_18683,N_19645);
nor U23418 (N_23418,N_19894,N_19780);
nand U23419 (N_23419,N_18608,N_20949);
xnor U23420 (N_23420,N_20640,N_19373);
and U23421 (N_23421,N_20404,N_19754);
or U23422 (N_23422,N_20118,N_18206);
or U23423 (N_23423,N_18494,N_18211);
nor U23424 (N_23424,N_20447,N_18748);
nand U23425 (N_23425,N_19639,N_18310);
and U23426 (N_23426,N_20517,N_20842);
nor U23427 (N_23427,N_19752,N_20491);
and U23428 (N_23428,N_19045,N_19667);
nor U23429 (N_23429,N_18311,N_18859);
xnor U23430 (N_23430,N_19756,N_20872);
xor U23431 (N_23431,N_18076,N_19608);
nand U23432 (N_23432,N_20160,N_20005);
nor U23433 (N_23433,N_20161,N_19492);
nand U23434 (N_23434,N_18028,N_19040);
nor U23435 (N_23435,N_18106,N_19034);
and U23436 (N_23436,N_18227,N_19690);
nor U23437 (N_23437,N_19756,N_19650);
or U23438 (N_23438,N_18373,N_19229);
or U23439 (N_23439,N_19333,N_18812);
and U23440 (N_23440,N_19962,N_18241);
nor U23441 (N_23441,N_19993,N_19489);
and U23442 (N_23442,N_18567,N_18327);
nand U23443 (N_23443,N_19107,N_19572);
and U23444 (N_23444,N_18449,N_19699);
nand U23445 (N_23445,N_20117,N_19382);
xnor U23446 (N_23446,N_19067,N_20021);
nand U23447 (N_23447,N_20984,N_20171);
or U23448 (N_23448,N_20062,N_18648);
or U23449 (N_23449,N_20446,N_20878);
nor U23450 (N_23450,N_18029,N_20305);
or U23451 (N_23451,N_20057,N_18935);
nand U23452 (N_23452,N_19760,N_20404);
xor U23453 (N_23453,N_19528,N_18769);
or U23454 (N_23454,N_20955,N_20599);
nor U23455 (N_23455,N_20541,N_18356);
or U23456 (N_23456,N_20237,N_18859);
nor U23457 (N_23457,N_19113,N_19428);
and U23458 (N_23458,N_20690,N_19144);
and U23459 (N_23459,N_18281,N_18747);
nor U23460 (N_23460,N_20299,N_18896);
and U23461 (N_23461,N_18544,N_20386);
nand U23462 (N_23462,N_19301,N_19349);
or U23463 (N_23463,N_19032,N_20717);
and U23464 (N_23464,N_18861,N_18601);
nor U23465 (N_23465,N_18376,N_18916);
and U23466 (N_23466,N_20616,N_18654);
and U23467 (N_23467,N_20742,N_18099);
and U23468 (N_23468,N_19681,N_18955);
or U23469 (N_23469,N_18500,N_18489);
xor U23470 (N_23470,N_19999,N_19993);
nand U23471 (N_23471,N_19935,N_18406);
or U23472 (N_23472,N_20405,N_19970);
or U23473 (N_23473,N_18363,N_20337);
nand U23474 (N_23474,N_18504,N_19342);
or U23475 (N_23475,N_19153,N_20001);
or U23476 (N_23476,N_19841,N_18346);
xnor U23477 (N_23477,N_18526,N_20088);
or U23478 (N_23478,N_20226,N_20917);
or U23479 (N_23479,N_18499,N_19419);
and U23480 (N_23480,N_19489,N_18528);
and U23481 (N_23481,N_18422,N_18138);
nand U23482 (N_23482,N_20675,N_19632);
and U23483 (N_23483,N_18717,N_20528);
nor U23484 (N_23484,N_20338,N_18387);
and U23485 (N_23485,N_20426,N_18129);
nand U23486 (N_23486,N_18673,N_18067);
nor U23487 (N_23487,N_19095,N_18812);
nand U23488 (N_23488,N_20673,N_20444);
nand U23489 (N_23489,N_18594,N_18935);
or U23490 (N_23490,N_19825,N_18826);
xnor U23491 (N_23491,N_18492,N_19603);
and U23492 (N_23492,N_18847,N_18257);
or U23493 (N_23493,N_20165,N_18253);
nor U23494 (N_23494,N_18033,N_18402);
and U23495 (N_23495,N_18128,N_19625);
nor U23496 (N_23496,N_19131,N_18825);
and U23497 (N_23497,N_18720,N_18290);
nand U23498 (N_23498,N_20826,N_18169);
or U23499 (N_23499,N_19965,N_18417);
nand U23500 (N_23500,N_19752,N_18314);
nand U23501 (N_23501,N_19397,N_19967);
and U23502 (N_23502,N_18339,N_20838);
nor U23503 (N_23503,N_19461,N_18168);
or U23504 (N_23504,N_18595,N_18865);
nand U23505 (N_23505,N_18623,N_18002);
nand U23506 (N_23506,N_19550,N_18062);
nand U23507 (N_23507,N_18364,N_18629);
nand U23508 (N_23508,N_18482,N_20128);
nand U23509 (N_23509,N_18494,N_18002);
nand U23510 (N_23510,N_20112,N_20828);
nor U23511 (N_23511,N_20656,N_19598);
nor U23512 (N_23512,N_19508,N_18832);
xnor U23513 (N_23513,N_20682,N_18650);
or U23514 (N_23514,N_18973,N_19142);
and U23515 (N_23515,N_19293,N_19121);
nand U23516 (N_23516,N_19280,N_18100);
or U23517 (N_23517,N_18351,N_18383);
xor U23518 (N_23518,N_19561,N_20758);
and U23519 (N_23519,N_18394,N_18785);
xor U23520 (N_23520,N_19969,N_18978);
and U23521 (N_23521,N_18052,N_20119);
and U23522 (N_23522,N_19136,N_20690);
and U23523 (N_23523,N_19786,N_18800);
and U23524 (N_23524,N_20449,N_20370);
and U23525 (N_23525,N_19832,N_20594);
nor U23526 (N_23526,N_20015,N_20068);
and U23527 (N_23527,N_18556,N_20257);
or U23528 (N_23528,N_18438,N_19435);
or U23529 (N_23529,N_18599,N_20401);
nand U23530 (N_23530,N_20102,N_18820);
nand U23531 (N_23531,N_20941,N_19499);
xor U23532 (N_23532,N_18440,N_20159);
and U23533 (N_23533,N_18176,N_19064);
or U23534 (N_23534,N_20884,N_19309);
or U23535 (N_23535,N_18591,N_20426);
xor U23536 (N_23536,N_19950,N_19900);
nor U23537 (N_23537,N_18366,N_18182);
and U23538 (N_23538,N_20743,N_19831);
and U23539 (N_23539,N_19562,N_19770);
nor U23540 (N_23540,N_18333,N_18540);
or U23541 (N_23541,N_19623,N_18740);
nor U23542 (N_23542,N_20080,N_20551);
nor U23543 (N_23543,N_20127,N_18373);
or U23544 (N_23544,N_20697,N_19386);
or U23545 (N_23545,N_19854,N_19373);
and U23546 (N_23546,N_20689,N_19990);
xnor U23547 (N_23547,N_20455,N_18076);
nand U23548 (N_23548,N_20736,N_20389);
nand U23549 (N_23549,N_18307,N_20809);
and U23550 (N_23550,N_19241,N_19812);
or U23551 (N_23551,N_19077,N_18057);
or U23552 (N_23552,N_20125,N_20142);
or U23553 (N_23553,N_19156,N_20610);
nand U23554 (N_23554,N_18473,N_19914);
nand U23555 (N_23555,N_18361,N_18243);
nor U23556 (N_23556,N_18247,N_19118);
or U23557 (N_23557,N_20771,N_20919);
xnor U23558 (N_23558,N_20870,N_20546);
and U23559 (N_23559,N_20166,N_19958);
or U23560 (N_23560,N_19455,N_19775);
nor U23561 (N_23561,N_19814,N_19628);
and U23562 (N_23562,N_19940,N_19863);
nand U23563 (N_23563,N_19346,N_20479);
xnor U23564 (N_23564,N_18397,N_19537);
and U23565 (N_23565,N_19279,N_18071);
xor U23566 (N_23566,N_18356,N_18533);
or U23567 (N_23567,N_19175,N_18714);
and U23568 (N_23568,N_18127,N_18218);
nand U23569 (N_23569,N_20949,N_20451);
or U23570 (N_23570,N_20333,N_20245);
and U23571 (N_23571,N_18027,N_19853);
or U23572 (N_23572,N_18749,N_20292);
and U23573 (N_23573,N_19392,N_19922);
nand U23574 (N_23574,N_18824,N_20619);
and U23575 (N_23575,N_20976,N_20622);
nor U23576 (N_23576,N_18941,N_20844);
nand U23577 (N_23577,N_19876,N_18131);
nand U23578 (N_23578,N_20743,N_19309);
nand U23579 (N_23579,N_18643,N_20638);
nor U23580 (N_23580,N_18986,N_18802);
nand U23581 (N_23581,N_19160,N_18395);
nor U23582 (N_23582,N_20295,N_20604);
xor U23583 (N_23583,N_20520,N_19605);
nand U23584 (N_23584,N_20849,N_20184);
nor U23585 (N_23585,N_18967,N_19203);
or U23586 (N_23586,N_19685,N_19205);
nand U23587 (N_23587,N_20879,N_18229);
or U23588 (N_23588,N_18773,N_20061);
nor U23589 (N_23589,N_19059,N_18275);
xor U23590 (N_23590,N_18570,N_19077);
nor U23591 (N_23591,N_19727,N_20781);
or U23592 (N_23592,N_19123,N_19328);
nand U23593 (N_23593,N_19939,N_20068);
nand U23594 (N_23594,N_18742,N_20338);
nand U23595 (N_23595,N_20592,N_18253);
and U23596 (N_23596,N_20550,N_18448);
or U23597 (N_23597,N_18552,N_19924);
xnor U23598 (N_23598,N_18061,N_18402);
nor U23599 (N_23599,N_20864,N_18740);
xnor U23600 (N_23600,N_18242,N_18512);
or U23601 (N_23601,N_19357,N_19576);
nand U23602 (N_23602,N_19844,N_19795);
and U23603 (N_23603,N_19807,N_19376);
xnor U23604 (N_23604,N_19345,N_18076);
and U23605 (N_23605,N_18390,N_18622);
nand U23606 (N_23606,N_19468,N_19638);
or U23607 (N_23607,N_19802,N_20101);
nor U23608 (N_23608,N_20495,N_19932);
or U23609 (N_23609,N_20152,N_19340);
and U23610 (N_23610,N_19515,N_18709);
and U23611 (N_23611,N_18488,N_20049);
or U23612 (N_23612,N_18562,N_20210);
nor U23613 (N_23613,N_19583,N_19521);
and U23614 (N_23614,N_19606,N_19993);
or U23615 (N_23615,N_18277,N_19494);
and U23616 (N_23616,N_19824,N_19962);
or U23617 (N_23617,N_18069,N_18884);
or U23618 (N_23618,N_20139,N_19083);
nand U23619 (N_23619,N_19759,N_19061);
and U23620 (N_23620,N_18139,N_18627);
nand U23621 (N_23621,N_18902,N_18372);
or U23622 (N_23622,N_19307,N_19969);
and U23623 (N_23623,N_18385,N_20392);
xnor U23624 (N_23624,N_19895,N_19067);
or U23625 (N_23625,N_19244,N_20674);
nor U23626 (N_23626,N_19005,N_20942);
and U23627 (N_23627,N_19176,N_18482);
and U23628 (N_23628,N_19747,N_19790);
xnor U23629 (N_23629,N_18616,N_18884);
or U23630 (N_23630,N_18164,N_19305);
and U23631 (N_23631,N_19282,N_18005);
nand U23632 (N_23632,N_20251,N_18046);
and U23633 (N_23633,N_20711,N_18932);
nor U23634 (N_23634,N_19422,N_20527);
nand U23635 (N_23635,N_18941,N_18235);
nor U23636 (N_23636,N_19863,N_19011);
or U23637 (N_23637,N_20948,N_18525);
or U23638 (N_23638,N_20059,N_19908);
and U23639 (N_23639,N_19256,N_18561);
nor U23640 (N_23640,N_18407,N_18092);
nor U23641 (N_23641,N_19140,N_20777);
nand U23642 (N_23642,N_20058,N_18623);
nor U23643 (N_23643,N_18608,N_18351);
xnor U23644 (N_23644,N_18025,N_20040);
nor U23645 (N_23645,N_20362,N_18134);
nand U23646 (N_23646,N_19827,N_18390);
nand U23647 (N_23647,N_19879,N_19589);
nor U23648 (N_23648,N_19117,N_20225);
or U23649 (N_23649,N_20226,N_18016);
nand U23650 (N_23650,N_20584,N_19035);
nor U23651 (N_23651,N_18694,N_20843);
nand U23652 (N_23652,N_19383,N_20615);
and U23653 (N_23653,N_20889,N_20757);
or U23654 (N_23654,N_18817,N_20170);
xnor U23655 (N_23655,N_18706,N_20702);
nor U23656 (N_23656,N_19487,N_19978);
nor U23657 (N_23657,N_19181,N_18680);
xor U23658 (N_23658,N_19486,N_20060);
and U23659 (N_23659,N_18611,N_19272);
xor U23660 (N_23660,N_20440,N_18292);
or U23661 (N_23661,N_20203,N_19725);
and U23662 (N_23662,N_20559,N_20639);
nor U23663 (N_23663,N_19994,N_20703);
and U23664 (N_23664,N_18249,N_19495);
nor U23665 (N_23665,N_19284,N_19808);
and U23666 (N_23666,N_20868,N_18745);
nor U23667 (N_23667,N_18346,N_19857);
or U23668 (N_23668,N_20620,N_19924);
xnor U23669 (N_23669,N_20270,N_19862);
or U23670 (N_23670,N_20258,N_20410);
nor U23671 (N_23671,N_20680,N_20783);
nand U23672 (N_23672,N_19796,N_19419);
nor U23673 (N_23673,N_18811,N_18903);
nor U23674 (N_23674,N_18067,N_18186);
nand U23675 (N_23675,N_19164,N_20529);
and U23676 (N_23676,N_20855,N_20724);
or U23677 (N_23677,N_19580,N_18781);
and U23678 (N_23678,N_18005,N_18227);
or U23679 (N_23679,N_20908,N_20693);
and U23680 (N_23680,N_20344,N_20633);
nor U23681 (N_23681,N_18905,N_20982);
nor U23682 (N_23682,N_19171,N_19899);
and U23683 (N_23683,N_18411,N_18441);
nand U23684 (N_23684,N_20709,N_19590);
and U23685 (N_23685,N_19524,N_18812);
nor U23686 (N_23686,N_19882,N_19904);
and U23687 (N_23687,N_19248,N_19346);
or U23688 (N_23688,N_18309,N_19086);
and U23689 (N_23689,N_19536,N_19544);
or U23690 (N_23690,N_19778,N_18910);
nor U23691 (N_23691,N_20086,N_19933);
and U23692 (N_23692,N_18742,N_20914);
and U23693 (N_23693,N_19516,N_19307);
and U23694 (N_23694,N_18947,N_18244);
and U23695 (N_23695,N_19889,N_18888);
or U23696 (N_23696,N_20747,N_20908);
or U23697 (N_23697,N_18217,N_20498);
nand U23698 (N_23698,N_20051,N_18715);
and U23699 (N_23699,N_20809,N_20019);
or U23700 (N_23700,N_20972,N_18188);
nor U23701 (N_23701,N_18947,N_18288);
or U23702 (N_23702,N_18543,N_19535);
and U23703 (N_23703,N_19283,N_19060);
nand U23704 (N_23704,N_18671,N_18254);
xnor U23705 (N_23705,N_19895,N_19040);
and U23706 (N_23706,N_18703,N_18427);
nor U23707 (N_23707,N_19157,N_20943);
and U23708 (N_23708,N_20312,N_18509);
nand U23709 (N_23709,N_19569,N_19004);
nor U23710 (N_23710,N_20014,N_18789);
nand U23711 (N_23711,N_18178,N_18273);
and U23712 (N_23712,N_19676,N_18584);
and U23713 (N_23713,N_19769,N_18047);
or U23714 (N_23714,N_20788,N_19019);
nor U23715 (N_23715,N_18227,N_20554);
nand U23716 (N_23716,N_20530,N_19809);
or U23717 (N_23717,N_18730,N_20719);
nor U23718 (N_23718,N_19922,N_19952);
nor U23719 (N_23719,N_18819,N_19784);
xnor U23720 (N_23720,N_18284,N_20097);
and U23721 (N_23721,N_20926,N_20555);
nand U23722 (N_23722,N_18138,N_20546);
and U23723 (N_23723,N_20942,N_18009);
and U23724 (N_23724,N_20876,N_18024);
nor U23725 (N_23725,N_19125,N_20811);
and U23726 (N_23726,N_19214,N_20931);
and U23727 (N_23727,N_19849,N_18200);
and U23728 (N_23728,N_19014,N_20363);
or U23729 (N_23729,N_20719,N_20157);
nor U23730 (N_23730,N_20223,N_18580);
or U23731 (N_23731,N_19795,N_18285);
or U23732 (N_23732,N_19502,N_18898);
and U23733 (N_23733,N_19993,N_19634);
and U23734 (N_23734,N_18102,N_20711);
nand U23735 (N_23735,N_18923,N_18247);
nand U23736 (N_23736,N_20698,N_19088);
or U23737 (N_23737,N_20620,N_18181);
xnor U23738 (N_23738,N_19998,N_18697);
nand U23739 (N_23739,N_20361,N_19302);
or U23740 (N_23740,N_18168,N_18898);
nor U23741 (N_23741,N_18438,N_19817);
nand U23742 (N_23742,N_20391,N_18412);
nor U23743 (N_23743,N_19394,N_19608);
and U23744 (N_23744,N_18730,N_19480);
nand U23745 (N_23745,N_18982,N_19296);
nand U23746 (N_23746,N_19739,N_20867);
nor U23747 (N_23747,N_18618,N_18552);
or U23748 (N_23748,N_19005,N_18171);
nand U23749 (N_23749,N_18380,N_18454);
nor U23750 (N_23750,N_19596,N_19014);
nand U23751 (N_23751,N_18406,N_19257);
nor U23752 (N_23752,N_20776,N_18306);
nand U23753 (N_23753,N_18338,N_19972);
nand U23754 (N_23754,N_18340,N_19228);
nor U23755 (N_23755,N_20249,N_18538);
nand U23756 (N_23756,N_20368,N_19536);
nor U23757 (N_23757,N_20861,N_19118);
nor U23758 (N_23758,N_20202,N_19860);
or U23759 (N_23759,N_20168,N_20166);
nand U23760 (N_23760,N_19048,N_20650);
xnor U23761 (N_23761,N_20303,N_20659);
nor U23762 (N_23762,N_20651,N_18600);
nor U23763 (N_23763,N_19640,N_20137);
or U23764 (N_23764,N_19074,N_19365);
or U23765 (N_23765,N_18988,N_20949);
nand U23766 (N_23766,N_19116,N_20952);
or U23767 (N_23767,N_19683,N_19860);
nand U23768 (N_23768,N_20393,N_20897);
xnor U23769 (N_23769,N_18052,N_19634);
nor U23770 (N_23770,N_19288,N_20122);
or U23771 (N_23771,N_18817,N_20461);
nand U23772 (N_23772,N_20688,N_20433);
and U23773 (N_23773,N_18692,N_18015);
and U23774 (N_23774,N_20589,N_18087);
nand U23775 (N_23775,N_19544,N_20639);
nor U23776 (N_23776,N_19509,N_18479);
nor U23777 (N_23777,N_18653,N_19735);
and U23778 (N_23778,N_19632,N_18468);
nand U23779 (N_23779,N_20004,N_20184);
and U23780 (N_23780,N_19198,N_20226);
and U23781 (N_23781,N_20394,N_20914);
xor U23782 (N_23782,N_19741,N_20186);
nand U23783 (N_23783,N_18348,N_18479);
and U23784 (N_23784,N_19587,N_19651);
and U23785 (N_23785,N_18754,N_19787);
and U23786 (N_23786,N_18983,N_19195);
or U23787 (N_23787,N_18736,N_19408);
nor U23788 (N_23788,N_18861,N_18965);
nor U23789 (N_23789,N_19132,N_18535);
or U23790 (N_23790,N_19838,N_20597);
and U23791 (N_23791,N_18451,N_20111);
and U23792 (N_23792,N_18778,N_19708);
or U23793 (N_23793,N_19768,N_18341);
and U23794 (N_23794,N_20160,N_18184);
or U23795 (N_23795,N_19151,N_20915);
and U23796 (N_23796,N_19711,N_20181);
nor U23797 (N_23797,N_19229,N_18091);
nor U23798 (N_23798,N_20200,N_20587);
and U23799 (N_23799,N_20427,N_18047);
and U23800 (N_23800,N_19787,N_18904);
nand U23801 (N_23801,N_18247,N_19799);
nor U23802 (N_23802,N_19416,N_18652);
nand U23803 (N_23803,N_19478,N_19198);
xnor U23804 (N_23804,N_20050,N_19577);
xor U23805 (N_23805,N_19745,N_20501);
xor U23806 (N_23806,N_18449,N_20901);
xor U23807 (N_23807,N_20821,N_18504);
nand U23808 (N_23808,N_18653,N_18698);
and U23809 (N_23809,N_18845,N_18106);
nand U23810 (N_23810,N_19948,N_18383);
or U23811 (N_23811,N_18370,N_20880);
or U23812 (N_23812,N_20435,N_19928);
nand U23813 (N_23813,N_19353,N_18198);
and U23814 (N_23814,N_20539,N_18295);
nor U23815 (N_23815,N_20557,N_18654);
nor U23816 (N_23816,N_20817,N_18322);
nand U23817 (N_23817,N_18016,N_18251);
xor U23818 (N_23818,N_18712,N_18910);
or U23819 (N_23819,N_18698,N_18234);
xnor U23820 (N_23820,N_19396,N_18457);
and U23821 (N_23821,N_20689,N_18090);
and U23822 (N_23822,N_19001,N_18816);
or U23823 (N_23823,N_20979,N_19693);
and U23824 (N_23824,N_18207,N_20081);
nor U23825 (N_23825,N_20223,N_18256);
and U23826 (N_23826,N_19316,N_18026);
nand U23827 (N_23827,N_18855,N_19149);
nand U23828 (N_23828,N_18146,N_18141);
and U23829 (N_23829,N_19902,N_20238);
nor U23830 (N_23830,N_19059,N_20529);
and U23831 (N_23831,N_19055,N_20382);
nor U23832 (N_23832,N_20287,N_20699);
nor U23833 (N_23833,N_19605,N_18714);
nand U23834 (N_23834,N_19314,N_19371);
or U23835 (N_23835,N_20647,N_18074);
or U23836 (N_23836,N_20176,N_19302);
and U23837 (N_23837,N_20388,N_20826);
and U23838 (N_23838,N_19769,N_19596);
xnor U23839 (N_23839,N_20000,N_18369);
and U23840 (N_23840,N_20893,N_20591);
or U23841 (N_23841,N_20375,N_19673);
or U23842 (N_23842,N_18730,N_18770);
nor U23843 (N_23843,N_19136,N_19316);
or U23844 (N_23844,N_19718,N_18821);
or U23845 (N_23845,N_19259,N_18125);
nor U23846 (N_23846,N_20170,N_19020);
xnor U23847 (N_23847,N_19955,N_20322);
or U23848 (N_23848,N_18492,N_18033);
or U23849 (N_23849,N_19525,N_19625);
xnor U23850 (N_23850,N_18865,N_18681);
and U23851 (N_23851,N_20012,N_19586);
nand U23852 (N_23852,N_18133,N_19778);
nor U23853 (N_23853,N_18655,N_20550);
nor U23854 (N_23854,N_19007,N_19866);
and U23855 (N_23855,N_18249,N_19259);
nand U23856 (N_23856,N_20048,N_19871);
nand U23857 (N_23857,N_18481,N_20239);
or U23858 (N_23858,N_18250,N_18819);
and U23859 (N_23859,N_19289,N_18441);
or U23860 (N_23860,N_19131,N_20172);
and U23861 (N_23861,N_20295,N_19757);
nor U23862 (N_23862,N_19830,N_19053);
nand U23863 (N_23863,N_20496,N_19335);
nor U23864 (N_23864,N_18495,N_19326);
or U23865 (N_23865,N_18865,N_20817);
nand U23866 (N_23866,N_20741,N_18262);
and U23867 (N_23867,N_18599,N_19783);
nor U23868 (N_23868,N_18829,N_18129);
or U23869 (N_23869,N_19977,N_20686);
or U23870 (N_23870,N_18331,N_19747);
nor U23871 (N_23871,N_20576,N_19206);
or U23872 (N_23872,N_20322,N_18705);
xnor U23873 (N_23873,N_18891,N_18696);
and U23874 (N_23874,N_18416,N_19436);
nand U23875 (N_23875,N_20405,N_19242);
nand U23876 (N_23876,N_20014,N_20412);
and U23877 (N_23877,N_18540,N_19193);
nand U23878 (N_23878,N_18818,N_20305);
nand U23879 (N_23879,N_19179,N_19857);
nand U23880 (N_23880,N_18794,N_18556);
or U23881 (N_23881,N_20115,N_19681);
and U23882 (N_23882,N_20531,N_20038);
nand U23883 (N_23883,N_18402,N_19429);
nor U23884 (N_23884,N_19651,N_18207);
nand U23885 (N_23885,N_20408,N_18845);
or U23886 (N_23886,N_19075,N_19356);
xor U23887 (N_23887,N_19296,N_19640);
and U23888 (N_23888,N_18612,N_19582);
nor U23889 (N_23889,N_20953,N_18267);
nor U23890 (N_23890,N_19602,N_20881);
and U23891 (N_23891,N_20058,N_19526);
xnor U23892 (N_23892,N_19322,N_19962);
or U23893 (N_23893,N_19502,N_18355);
nor U23894 (N_23894,N_20298,N_20708);
nand U23895 (N_23895,N_20849,N_20258);
or U23896 (N_23896,N_18203,N_20896);
and U23897 (N_23897,N_18758,N_19419);
nand U23898 (N_23898,N_19635,N_19050);
and U23899 (N_23899,N_20941,N_20625);
and U23900 (N_23900,N_20596,N_18378);
nand U23901 (N_23901,N_18808,N_18362);
nand U23902 (N_23902,N_20486,N_18117);
and U23903 (N_23903,N_20517,N_19991);
and U23904 (N_23904,N_19517,N_18240);
nor U23905 (N_23905,N_18027,N_19901);
nand U23906 (N_23906,N_20695,N_20933);
nand U23907 (N_23907,N_19201,N_18037);
xor U23908 (N_23908,N_19611,N_20658);
or U23909 (N_23909,N_19829,N_18012);
and U23910 (N_23910,N_18237,N_18943);
or U23911 (N_23911,N_19285,N_18552);
nor U23912 (N_23912,N_19828,N_20070);
and U23913 (N_23913,N_20095,N_20977);
or U23914 (N_23914,N_18793,N_18531);
or U23915 (N_23915,N_18292,N_20190);
and U23916 (N_23916,N_20201,N_18229);
xor U23917 (N_23917,N_20340,N_18145);
and U23918 (N_23918,N_20501,N_18639);
xor U23919 (N_23919,N_18987,N_20790);
or U23920 (N_23920,N_20914,N_19055);
or U23921 (N_23921,N_18155,N_20545);
and U23922 (N_23922,N_20806,N_20601);
and U23923 (N_23923,N_19212,N_19959);
and U23924 (N_23924,N_20553,N_18103);
nor U23925 (N_23925,N_19835,N_18895);
and U23926 (N_23926,N_19789,N_18732);
nand U23927 (N_23927,N_18492,N_20135);
or U23928 (N_23928,N_18245,N_19826);
or U23929 (N_23929,N_20823,N_19134);
or U23930 (N_23930,N_19791,N_20870);
nor U23931 (N_23931,N_19301,N_18680);
nor U23932 (N_23932,N_20881,N_20162);
nor U23933 (N_23933,N_20412,N_20366);
nor U23934 (N_23934,N_19562,N_19749);
and U23935 (N_23935,N_18926,N_18141);
and U23936 (N_23936,N_20612,N_18965);
or U23937 (N_23937,N_18859,N_19185);
xor U23938 (N_23938,N_20656,N_20755);
and U23939 (N_23939,N_18554,N_20031);
and U23940 (N_23940,N_18092,N_20776);
nor U23941 (N_23941,N_19219,N_19351);
nor U23942 (N_23942,N_20292,N_19455);
nand U23943 (N_23943,N_20356,N_18566);
nor U23944 (N_23944,N_18461,N_19470);
or U23945 (N_23945,N_19392,N_19086);
nor U23946 (N_23946,N_19683,N_18285);
nand U23947 (N_23947,N_20964,N_20278);
nor U23948 (N_23948,N_18290,N_18398);
nor U23949 (N_23949,N_20358,N_18513);
nor U23950 (N_23950,N_19698,N_18654);
nand U23951 (N_23951,N_18705,N_18813);
nand U23952 (N_23952,N_20710,N_20876);
xor U23953 (N_23953,N_18332,N_19107);
and U23954 (N_23954,N_18290,N_18942);
xor U23955 (N_23955,N_20077,N_19603);
nand U23956 (N_23956,N_18239,N_18979);
or U23957 (N_23957,N_18397,N_20491);
nor U23958 (N_23958,N_20438,N_18770);
and U23959 (N_23959,N_18452,N_20363);
xnor U23960 (N_23960,N_18436,N_19419);
or U23961 (N_23961,N_19932,N_20838);
nand U23962 (N_23962,N_19843,N_19512);
nor U23963 (N_23963,N_19500,N_18716);
and U23964 (N_23964,N_18950,N_20983);
and U23965 (N_23965,N_20820,N_18719);
xnor U23966 (N_23966,N_18096,N_19959);
nand U23967 (N_23967,N_18869,N_20371);
or U23968 (N_23968,N_20572,N_20085);
nand U23969 (N_23969,N_20004,N_19118);
nand U23970 (N_23970,N_20984,N_19777);
or U23971 (N_23971,N_19370,N_19332);
or U23972 (N_23972,N_20252,N_20232);
or U23973 (N_23973,N_19198,N_20302);
xor U23974 (N_23974,N_19505,N_20622);
and U23975 (N_23975,N_19062,N_20133);
and U23976 (N_23976,N_19799,N_20125);
nand U23977 (N_23977,N_19149,N_20791);
nor U23978 (N_23978,N_19995,N_20252);
and U23979 (N_23979,N_18743,N_20664);
and U23980 (N_23980,N_18426,N_19632);
nor U23981 (N_23981,N_19751,N_19802);
nand U23982 (N_23982,N_18831,N_19874);
and U23983 (N_23983,N_18832,N_20146);
or U23984 (N_23984,N_20591,N_18365);
and U23985 (N_23985,N_18309,N_18683);
or U23986 (N_23986,N_20447,N_20048);
nor U23987 (N_23987,N_20008,N_20296);
or U23988 (N_23988,N_19793,N_20669);
and U23989 (N_23989,N_19173,N_19725);
nand U23990 (N_23990,N_20954,N_18729);
nor U23991 (N_23991,N_19438,N_19154);
or U23992 (N_23992,N_20840,N_20429);
and U23993 (N_23993,N_19335,N_18674);
or U23994 (N_23994,N_19587,N_18197);
nand U23995 (N_23995,N_19676,N_18876);
nor U23996 (N_23996,N_19634,N_20426);
or U23997 (N_23997,N_19624,N_18584);
and U23998 (N_23998,N_20938,N_18181);
and U23999 (N_23999,N_19394,N_19809);
or U24000 (N_24000,N_21725,N_21292);
or U24001 (N_24001,N_21823,N_22954);
nor U24002 (N_24002,N_21594,N_22124);
nor U24003 (N_24003,N_22877,N_21205);
xnor U24004 (N_24004,N_23936,N_22974);
or U24005 (N_24005,N_21991,N_22140);
or U24006 (N_24006,N_22719,N_21952);
and U24007 (N_24007,N_22761,N_21568);
nor U24008 (N_24008,N_22293,N_21282);
and U24009 (N_24009,N_21073,N_22408);
or U24010 (N_24010,N_21069,N_21114);
nor U24011 (N_24011,N_21459,N_22378);
nor U24012 (N_24012,N_22928,N_23118);
and U24013 (N_24013,N_21553,N_21284);
and U24014 (N_24014,N_22272,N_21634);
or U24015 (N_24015,N_21920,N_21390);
and U24016 (N_24016,N_21656,N_23937);
xor U24017 (N_24017,N_22855,N_21542);
or U24018 (N_24018,N_21515,N_21224);
xnor U24019 (N_24019,N_23970,N_22969);
nand U24020 (N_24020,N_23402,N_21331);
and U24021 (N_24021,N_22944,N_22031);
nor U24022 (N_24022,N_21572,N_23516);
or U24023 (N_24023,N_22423,N_23761);
and U24024 (N_24024,N_23600,N_23742);
nor U24025 (N_24025,N_23286,N_22906);
or U24026 (N_24026,N_22973,N_23120);
or U24027 (N_24027,N_22304,N_22320);
nand U24028 (N_24028,N_23032,N_21995);
nand U24029 (N_24029,N_23792,N_21537);
nor U24030 (N_24030,N_23218,N_21843);
nand U24031 (N_24031,N_22554,N_23269);
or U24032 (N_24032,N_22352,N_23755);
or U24033 (N_24033,N_21888,N_23663);
and U24034 (N_24034,N_23374,N_23444);
nand U24035 (N_24035,N_23955,N_23851);
and U24036 (N_24036,N_22844,N_23896);
or U24037 (N_24037,N_23299,N_23406);
xor U24038 (N_24038,N_21177,N_23775);
nand U24039 (N_24039,N_21646,N_23573);
nand U24040 (N_24040,N_23505,N_23447);
and U24041 (N_24041,N_22924,N_23488);
xor U24042 (N_24042,N_23574,N_23809);
nor U24043 (N_24043,N_21152,N_23123);
nor U24044 (N_24044,N_23750,N_22672);
or U24045 (N_24045,N_22407,N_23508);
or U24046 (N_24046,N_22958,N_23143);
nand U24047 (N_24047,N_22083,N_22778);
nand U24048 (N_24048,N_23025,N_23588);
nor U24049 (N_24049,N_23031,N_21853);
nand U24050 (N_24050,N_22206,N_23883);
or U24051 (N_24051,N_21321,N_23728);
or U24052 (N_24052,N_22702,N_22120);
and U24053 (N_24053,N_23021,N_23814);
or U24054 (N_24054,N_23745,N_22709);
nor U24055 (N_24055,N_23916,N_22533);
nor U24056 (N_24056,N_22575,N_23939);
nand U24057 (N_24057,N_23502,N_23008);
xor U24058 (N_24058,N_22870,N_22680);
nor U24059 (N_24059,N_23862,N_22972);
nor U24060 (N_24060,N_21828,N_21750);
nor U24061 (N_24061,N_23039,N_23456);
or U24062 (N_24062,N_23966,N_21779);
or U24063 (N_24063,N_23066,N_21000);
and U24064 (N_24064,N_23213,N_21720);
nand U24065 (N_24065,N_21157,N_21852);
or U24066 (N_24066,N_22905,N_21047);
and U24067 (N_24067,N_22627,N_21265);
nand U24068 (N_24068,N_23723,N_21567);
and U24069 (N_24069,N_21729,N_23919);
and U24070 (N_24070,N_21834,N_22400);
and U24071 (N_24071,N_23145,N_22223);
or U24072 (N_24072,N_23906,N_22332);
and U24073 (N_24073,N_23571,N_22292);
nand U24074 (N_24074,N_23355,N_21496);
nor U24075 (N_24075,N_22091,N_23304);
xnor U24076 (N_24076,N_23981,N_22325);
nor U24077 (N_24077,N_22699,N_23210);
nor U24078 (N_24078,N_22899,N_23378);
nor U24079 (N_24079,N_23385,N_23033);
nand U24080 (N_24080,N_23984,N_21717);
and U24081 (N_24081,N_23551,N_22619);
nor U24082 (N_24082,N_22570,N_23368);
and U24083 (N_24083,N_22115,N_22489);
nand U24084 (N_24084,N_23320,N_22035);
nor U24085 (N_24085,N_22903,N_23699);
nand U24086 (N_24086,N_23130,N_23389);
nor U24087 (N_24087,N_22455,N_23191);
and U24088 (N_24088,N_22321,N_22137);
nor U24089 (N_24089,N_22085,N_22545);
and U24090 (N_24090,N_21037,N_21557);
or U24091 (N_24091,N_23894,N_22664);
or U24092 (N_24092,N_21017,N_21765);
xor U24093 (N_24093,N_23659,N_23418);
and U24094 (N_24094,N_21870,N_21733);
nor U24095 (N_24095,N_22056,N_22708);
or U24096 (N_24096,N_22226,N_22801);
and U24097 (N_24097,N_22923,N_22937);
or U24098 (N_24098,N_21923,N_21156);
nor U24099 (N_24099,N_23560,N_23760);
or U24100 (N_24100,N_21016,N_22388);
or U24101 (N_24101,N_22333,N_23810);
or U24102 (N_24102,N_22825,N_23117);
nor U24103 (N_24103,N_21829,N_23382);
nand U24104 (N_24104,N_22979,N_22370);
or U24105 (N_24105,N_22481,N_22516);
nand U24106 (N_24106,N_22858,N_23094);
nor U24107 (N_24107,N_22948,N_21752);
nor U24108 (N_24108,N_23411,N_22757);
nor U24109 (N_24109,N_23122,N_23017);
or U24110 (N_24110,N_23057,N_21879);
and U24111 (N_24111,N_23969,N_21031);
nor U24112 (N_24112,N_23002,N_21874);
and U24113 (N_24113,N_21745,N_23434);
or U24114 (N_24114,N_22249,N_21289);
xnor U24115 (N_24115,N_23314,N_22326);
nand U24116 (N_24116,N_21743,N_23341);
and U24117 (N_24117,N_21094,N_22396);
or U24118 (N_24118,N_23869,N_23221);
nand U24119 (N_24119,N_23649,N_23759);
nor U24120 (N_24120,N_23071,N_22182);
and U24121 (N_24121,N_21066,N_22535);
or U24122 (N_24122,N_23973,N_23178);
nor U24123 (N_24123,N_23043,N_21238);
nand U24124 (N_24124,N_21245,N_22492);
nand U24125 (N_24125,N_22389,N_23662);
nand U24126 (N_24126,N_22945,N_23749);
nor U24127 (N_24127,N_22542,N_21294);
nand U24128 (N_24128,N_23954,N_23983);
nand U24129 (N_24129,N_21800,N_22376);
nor U24130 (N_24130,N_21820,N_23091);
nand U24131 (N_24131,N_21977,N_22068);
or U24132 (N_24132,N_22947,N_23487);
nor U24133 (N_24133,N_22071,N_22084);
nor U24134 (N_24134,N_23391,N_23591);
nor U24135 (N_24135,N_23978,N_22601);
or U24136 (N_24136,N_23914,N_22179);
nand U24137 (N_24137,N_22893,N_21077);
nand U24138 (N_24138,N_21970,N_23089);
nand U24139 (N_24139,N_21010,N_23373);
xnor U24140 (N_24140,N_23696,N_22706);
nor U24141 (N_24141,N_23986,N_21146);
and U24142 (N_24142,N_22902,N_23371);
nand U24143 (N_24143,N_22387,N_21526);
nand U24144 (N_24144,N_22172,N_21796);
or U24145 (N_24145,N_22777,N_22641);
and U24146 (N_24146,N_22462,N_23680);
or U24147 (N_24147,N_23791,N_21814);
nand U24148 (N_24148,N_21540,N_21285);
and U24149 (N_24149,N_21884,N_23853);
and U24150 (N_24150,N_23921,N_23482);
or U24151 (N_24151,N_21081,N_23764);
and U24152 (N_24152,N_22592,N_21601);
nand U24153 (N_24153,N_22475,N_23584);
or U24154 (N_24154,N_22136,N_21428);
nor U24155 (N_24155,N_21742,N_22534);
nor U24156 (N_24156,N_21639,N_23155);
or U24157 (N_24157,N_23525,N_21115);
and U24158 (N_24158,N_22269,N_22668);
or U24159 (N_24159,N_22631,N_23290);
or U24160 (N_24160,N_21642,N_23062);
nor U24161 (N_24161,N_21958,N_22162);
nor U24162 (N_24162,N_23518,N_21383);
or U24163 (N_24163,N_21830,N_23037);
or U24164 (N_24164,N_21994,N_23323);
nor U24165 (N_24165,N_23386,N_21242);
or U24166 (N_24166,N_21948,N_21666);
nand U24167 (N_24167,N_22341,N_23944);
and U24168 (N_24168,N_21524,N_23711);
nor U24169 (N_24169,N_21824,N_23042);
or U24170 (N_24170,N_21423,N_22322);
or U24171 (N_24171,N_23744,N_22665);
and U24172 (N_24172,N_21248,N_21438);
and U24173 (N_24173,N_22879,N_21297);
or U24174 (N_24174,N_23801,N_23654);
or U24175 (N_24175,N_21773,N_21314);
nand U24176 (N_24176,N_23892,N_23151);
nand U24177 (N_24177,N_21614,N_21174);
or U24178 (N_24178,N_21396,N_22482);
xor U24179 (N_24179,N_21237,N_23875);
xor U24180 (N_24180,N_21516,N_23284);
and U24181 (N_24181,N_21484,N_21334);
and U24182 (N_24182,N_21928,N_22549);
xor U24183 (N_24183,N_21650,N_22317);
nand U24184 (N_24184,N_22998,N_22814);
nor U24185 (N_24185,N_23412,N_21556);
nand U24186 (N_24186,N_22161,N_23367);
nand U24187 (N_24187,N_22291,N_23154);
xor U24188 (N_24188,N_22517,N_23507);
nand U24189 (N_24189,N_21789,N_23319);
xor U24190 (N_24190,N_21089,N_23835);
nor U24191 (N_24191,N_22415,N_21988);
nand U24192 (N_24192,N_22251,N_21147);
nor U24193 (N_24193,N_23459,N_23491);
nand U24194 (N_24194,N_23915,N_22882);
or U24195 (N_24195,N_22329,N_23825);
or U24196 (N_24196,N_21858,N_23509);
nor U24197 (N_24197,N_23471,N_21046);
nor U24198 (N_24198,N_22824,N_22051);
nor U24199 (N_24199,N_23831,N_23540);
or U24200 (N_24200,N_22017,N_22457);
and U24201 (N_24201,N_23627,N_21916);
or U24202 (N_24202,N_23812,N_21855);
nand U24203 (N_24203,N_23302,N_23683);
xor U24204 (N_24204,N_22960,N_21402);
xor U24205 (N_24205,N_23622,N_22817);
or U24206 (N_24206,N_22474,N_22577);
or U24207 (N_24207,N_22096,N_21451);
nand U24208 (N_24208,N_21838,N_21458);
nand U24209 (N_24209,N_21398,N_21757);
xor U24210 (N_24210,N_22134,N_23082);
nand U24211 (N_24211,N_23333,N_23099);
nor U24212 (N_24212,N_21783,N_21770);
or U24213 (N_24213,N_23454,N_23793);
nor U24214 (N_24214,N_22160,N_22839);
nand U24215 (N_24215,N_23283,N_22722);
or U24216 (N_24216,N_23818,N_22465);
xnor U24217 (N_24217,N_21809,N_23296);
or U24218 (N_24218,N_22561,N_22646);
nor U24219 (N_24219,N_22397,N_21586);
nand U24220 (N_24220,N_23643,N_23700);
or U24221 (N_24221,N_21247,N_22343);
xor U24222 (N_24222,N_23841,N_21637);
nor U24223 (N_24223,N_21761,N_22621);
nor U24224 (N_24224,N_23186,N_21731);
nor U24225 (N_24225,N_23826,N_21202);
and U24226 (N_24226,N_23293,N_22915);
and U24227 (N_24227,N_23055,N_23451);
nor U24228 (N_24228,N_22831,N_21219);
and U24229 (N_24229,N_23923,N_22956);
nor U24230 (N_24230,N_22738,N_22900);
xor U24231 (N_24231,N_21370,N_21145);
nand U24232 (N_24232,N_21984,N_21722);
nor U24233 (N_24233,N_22088,N_21564);
xnor U24234 (N_24234,N_23597,N_23716);
and U24235 (N_24235,N_22277,N_23985);
nand U24236 (N_24236,N_22864,N_22787);
xor U24237 (N_24237,N_21934,N_23542);
or U24238 (N_24238,N_23767,N_21148);
nand U24239 (N_24239,N_22530,N_22166);
nor U24240 (N_24240,N_22574,N_21444);
nand U24241 (N_24241,N_22185,N_22080);
and U24242 (N_24242,N_21025,N_23880);
and U24243 (N_24243,N_23946,N_21022);
or U24244 (N_24244,N_21559,N_21529);
and U24245 (N_24245,N_21118,N_22776);
nor U24246 (N_24246,N_22502,N_21096);
nand U24247 (N_24247,N_21036,N_22057);
nand U24248 (N_24248,N_22737,N_21348);
or U24249 (N_24249,N_22859,N_21661);
and U24250 (N_24250,N_22107,N_23442);
or U24251 (N_24251,N_23013,N_22135);
and U24252 (N_24252,N_22705,N_21042);
xor U24253 (N_24253,N_21619,N_22404);
and U24254 (N_24254,N_23429,N_23606);
and U24255 (N_24255,N_21197,N_23732);
or U24256 (N_24256,N_22605,N_21741);
and U24257 (N_24257,N_21710,N_22986);
nand U24258 (N_24258,N_22678,N_21771);
xnor U24259 (N_24259,N_21463,N_22469);
or U24260 (N_24260,N_21927,N_23504);
nor U24261 (N_24261,N_23100,N_21088);
nand U24262 (N_24262,N_21364,N_23840);
nor U24263 (N_24263,N_21123,N_23078);
nor U24264 (N_24264,N_22758,N_21164);
nand U24265 (N_24265,N_22072,N_23064);
and U24266 (N_24266,N_22361,N_21756);
and U24267 (N_24267,N_22532,N_22856);
xnor U24268 (N_24268,N_22132,N_22955);
xor U24269 (N_24269,N_22584,N_22997);
or U24270 (N_24270,N_23134,N_21502);
nor U24271 (N_24271,N_23431,N_21320);
and U24272 (N_24272,N_23462,N_23865);
nand U24273 (N_24273,N_22433,N_22466);
or U24274 (N_24274,N_22442,N_21277);
nor U24275 (N_24275,N_21176,N_23215);
or U24276 (N_24276,N_23537,N_21467);
nand U24277 (N_24277,N_23619,N_21850);
and U24278 (N_24278,N_22024,N_21167);
xor U24279 (N_24279,N_23205,N_23772);
nand U24280 (N_24280,N_23305,N_22496);
nor U24281 (N_24281,N_22186,N_23665);
nand U24282 (N_24282,N_22267,N_22591);
or U24283 (N_24283,N_23589,N_21687);
nand U24284 (N_24284,N_21659,N_22886);
or U24285 (N_24285,N_21454,N_21832);
xor U24286 (N_24286,N_23724,N_22984);
and U24287 (N_24287,N_21495,N_23223);
nand U24288 (N_24288,N_22794,N_22454);
nand U24289 (N_24289,N_21701,N_23149);
nor U24290 (N_24290,N_23138,N_21195);
and U24291 (N_24291,N_21813,N_23754);
nor U24292 (N_24292,N_22971,N_21091);
or U24293 (N_24293,N_21845,N_23125);
nand U24294 (N_24294,N_23131,N_22593);
and U24295 (N_24295,N_23212,N_22981);
and U24296 (N_24296,N_23763,N_21827);
nor U24297 (N_24297,N_22772,N_21272);
nand U24298 (N_24298,N_22345,N_21775);
and U24299 (N_24299,N_23365,N_22555);
xor U24300 (N_24300,N_21018,N_22036);
nor U24301 (N_24301,N_23332,N_23988);
or U24302 (N_24302,N_22044,N_23611);
nor U24303 (N_24303,N_22934,N_23357);
nand U24304 (N_24304,N_23360,N_22478);
and U24305 (N_24305,N_22418,N_21403);
nor U24306 (N_24306,N_23783,N_21474);
xnor U24307 (N_24307,N_23010,N_23563);
and U24308 (N_24308,N_21406,N_21216);
or U24309 (N_24309,N_21229,N_22047);
nor U24310 (N_24310,N_21239,N_23280);
or U24311 (N_24311,N_23244,N_21938);
or U24312 (N_24312,N_22774,N_22689);
nand U24313 (N_24313,N_21264,N_23706);
and U24314 (N_24314,N_22257,N_23852);
nand U24315 (N_24315,N_21552,N_21243);
or U24316 (N_24316,N_23803,N_21120);
nor U24317 (N_24317,N_23640,N_23762);
and U24318 (N_24318,N_23908,N_21440);
and U24319 (N_24319,N_21903,N_23498);
and U24320 (N_24320,N_23111,N_23593);
nand U24321 (N_24321,N_21732,N_23725);
nand U24322 (N_24322,N_23383,N_22355);
and U24323 (N_24323,N_21144,N_23048);
nor U24324 (N_24324,N_22691,N_22800);
or U24325 (N_24325,N_22909,N_23068);
nor U24326 (N_24326,N_22896,N_22806);
or U24327 (N_24327,N_23150,N_21449);
or U24328 (N_24328,N_23268,N_23115);
xnor U24329 (N_24329,N_22450,N_23583);
or U24330 (N_24330,N_22655,N_22965);
and U24331 (N_24331,N_22994,N_22437);
nor U24332 (N_24332,N_23576,N_23024);
or U24333 (N_24333,N_23888,N_23870);
nor U24334 (N_24334,N_22263,N_23463);
nand U24335 (N_24335,N_23347,N_21891);
nand U24336 (N_24336,N_21919,N_21034);
xor U24337 (N_24337,N_22007,N_21689);
nor U24338 (N_24338,N_23262,N_22495);
or U24339 (N_24339,N_22414,N_23233);
or U24340 (N_24340,N_21504,N_21186);
nor U24341 (N_24341,N_21367,N_21254);
or U24342 (N_24342,N_22180,N_21906);
or U24343 (N_24343,N_21924,N_21510);
nand U24344 (N_24344,N_22289,N_21108);
and U24345 (N_24345,N_22276,N_23848);
or U24346 (N_24346,N_23996,N_23168);
nor U24347 (N_24347,N_23179,N_23335);
or U24348 (N_24348,N_21393,N_21131);
or U24349 (N_24349,N_21468,N_21020);
and U24350 (N_24350,N_23227,N_22402);
and U24351 (N_24351,N_23208,N_22874);
and U24352 (N_24352,N_22792,N_22082);
nor U24353 (N_24353,N_23965,N_23077);
nand U24354 (N_24354,N_21751,N_23353);
nor U24355 (N_24355,N_22055,N_22254);
or U24356 (N_24356,N_23639,N_22541);
and U24357 (N_24357,N_23443,N_21992);
and U24358 (N_24358,N_21511,N_23421);
xnor U24359 (N_24359,N_21849,N_22034);
nand U24360 (N_24360,N_23202,N_21487);
nor U24361 (N_24361,N_21491,N_23833);
and U24362 (N_24362,N_23850,N_22919);
and U24363 (N_24363,N_23866,N_22459);
and U24364 (N_24364,N_23163,N_21269);
or U24365 (N_24365,N_23426,N_22330);
nor U24366 (N_24366,N_21226,N_23035);
or U24367 (N_24367,N_22014,N_21676);
nand U24368 (N_24368,N_23994,N_21006);
nand U24369 (N_24369,N_22013,N_23860);
nand U24370 (N_24370,N_21339,N_21868);
nor U24371 (N_24371,N_22148,N_23000);
and U24372 (N_24372,N_21442,N_21133);
or U24373 (N_24373,N_22360,N_21035);
or U24374 (N_24374,N_23925,N_22434);
xnor U24375 (N_24375,N_23050,N_21041);
or U24376 (N_24376,N_22287,N_23156);
nand U24377 (N_24377,N_23541,N_22790);
or U24378 (N_24378,N_23080,N_22191);
nand U24379 (N_24379,N_21966,N_21012);
or U24380 (N_24380,N_22500,N_22358);
nand U24381 (N_24381,N_21395,N_21525);
nor U24382 (N_24382,N_21143,N_21949);
and U24383 (N_24383,N_22901,N_21963);
nor U24384 (N_24384,N_22898,N_22959);
xnor U24385 (N_24385,N_23260,N_23846);
xor U24386 (N_24386,N_23387,N_21673);
or U24387 (N_24387,N_22209,N_22990);
xnor U24388 (N_24388,N_23673,N_23450);
or U24389 (N_24389,N_21441,N_23604);
xnor U24390 (N_24390,N_21972,N_21794);
and U24391 (N_24391,N_22066,N_22509);
nor U24392 (N_24392,N_22599,N_21471);
xor U24393 (N_24393,N_22610,N_22704);
nand U24394 (N_24394,N_22092,N_23348);
nor U24395 (N_24395,N_22229,N_23354);
nor U24396 (N_24396,N_21737,N_23631);
nand U24397 (N_24397,N_21158,N_21554);
or U24398 (N_24398,N_21962,N_23821);
or U24399 (N_24399,N_23295,N_22623);
nor U24400 (N_24400,N_23009,N_22413);
and U24401 (N_24401,N_21976,N_22061);
and U24402 (N_24402,N_21786,N_23110);
xor U24403 (N_24403,N_22883,N_23692);
xnor U24404 (N_24404,N_21132,N_23076);
and U24405 (N_24405,N_22198,N_22662);
nor U24406 (N_24406,N_23177,N_21384);
nor U24407 (N_24407,N_21935,N_23494);
nand U24408 (N_24408,N_21753,N_21578);
or U24409 (N_24409,N_23958,N_22027);
and U24410 (N_24410,N_21766,N_23250);
nand U24411 (N_24411,N_22525,N_22743);
or U24412 (N_24412,N_23952,N_21658);
nand U24413 (N_24413,N_22252,N_22245);
or U24414 (N_24414,N_22712,N_22580);
nand U24415 (N_24415,N_21846,N_21230);
xnor U24416 (N_24416,N_21355,N_22957);
and U24417 (N_24417,N_22319,N_21941);
nand U24418 (N_24418,N_21816,N_23172);
or U24419 (N_24419,N_23058,N_23396);
or U24420 (N_24420,N_22356,N_21549);
nand U24421 (N_24421,N_21647,N_22037);
or U24422 (N_24422,N_23489,N_22340);
nand U24423 (N_24423,N_22398,N_23404);
and U24424 (N_24424,N_22242,N_21283);
nand U24425 (N_24425,N_23379,N_21376);
or U24426 (N_24426,N_22836,N_21298);
nor U24427 (N_24427,N_21600,N_22529);
and U24428 (N_24428,N_22045,N_23838);
nor U24429 (N_24429,N_21806,N_23146);
xor U24430 (N_24430,N_21340,N_21629);
or U24431 (N_24431,N_21538,N_21173);
nor U24432 (N_24432,N_23514,N_22274);
nand U24433 (N_24433,N_22519,N_23207);
nor U24434 (N_24434,N_21175,N_21310);
or U24435 (N_24435,N_23733,N_22222);
nor U24436 (N_24436,N_23278,N_21327);
or U24437 (N_24437,N_21086,N_21956);
nor U24438 (N_24438,N_22552,N_21489);
and U24439 (N_24439,N_22985,N_22526);
nor U24440 (N_24440,N_22645,N_21545);
or U24441 (N_24441,N_23475,N_23562);
and U24442 (N_24442,N_23298,N_22564);
and U24443 (N_24443,N_23559,N_21214);
nand U24444 (N_24444,N_21119,N_22147);
nor U24445 (N_24445,N_22250,N_23940);
or U24446 (N_24446,N_21929,N_22150);
xor U24447 (N_24447,N_22904,N_21306);
nand U24448 (N_24448,N_23535,N_23049);
nor U24449 (N_24449,N_21772,N_22951);
or U24450 (N_24450,N_23633,N_22187);
nor U24451 (N_24451,N_22711,N_23521);
nor U24452 (N_24452,N_21712,N_23730);
nand U24453 (N_24453,N_21251,N_22246);
and U24454 (N_24454,N_23872,N_22867);
nor U24455 (N_24455,N_22038,N_21363);
nor U24456 (N_24456,N_22970,N_23625);
or U24457 (N_24457,N_21436,N_21985);
and U24458 (N_24458,N_21307,N_23439);
xor U24459 (N_24459,N_22108,N_22197);
nand U24460 (N_24460,N_21223,N_21345);
nand U24461 (N_24461,N_23085,N_21819);
or U24462 (N_24462,N_22681,N_21207);
or U24463 (N_24463,N_23811,N_21236);
nand U24464 (N_24464,N_23132,N_22062);
xor U24465 (N_24465,N_22950,N_22913);
and U24466 (N_24466,N_21790,N_23088);
nor U24467 (N_24467,N_21950,N_21975);
and U24468 (N_24468,N_21573,N_23081);
or U24469 (N_24469,N_22773,N_21836);
or U24470 (N_24470,N_23530,N_21953);
or U24471 (N_24471,N_23941,N_22546);
and U24472 (N_24472,N_22569,N_22829);
nand U24473 (N_24473,N_22916,N_22079);
and U24474 (N_24474,N_23710,N_21835);
nor U24475 (N_24475,N_21810,N_22324);
and U24476 (N_24476,N_21002,N_21099);
and U24477 (N_24477,N_23231,N_23199);
xor U24478 (N_24478,N_22003,N_21462);
and U24479 (N_24479,N_23859,N_21678);
nor U24480 (N_24480,N_21486,N_23637);
or U24481 (N_24481,N_23282,N_21437);
xnor U24482 (N_24482,N_22169,N_23300);
or U24483 (N_24483,N_21574,N_21873);
nand U24484 (N_24484,N_23737,N_21569);
and U24485 (N_24485,N_23339,N_22302);
nand U24486 (N_24486,N_22406,N_21445);
or U24487 (N_24487,N_23877,N_22953);
or U24488 (N_24488,N_23030,N_23479);
and U24489 (N_24489,N_21851,N_22102);
or U24490 (N_24490,N_21268,N_21802);
or U24491 (N_24491,N_22690,N_22821);
or U24492 (N_24492,N_21135,N_22365);
xnor U24493 (N_24493,N_23170,N_22931);
nand U24494 (N_24494,N_21004,N_22327);
nor U24495 (N_24495,N_23175,N_22967);
and U24496 (N_24496,N_23666,N_23336);
and U24497 (N_24497,N_23552,N_22010);
or U24498 (N_24498,N_21630,N_22349);
or U24499 (N_24499,N_23097,N_21409);
or U24500 (N_24500,N_21369,N_21703);
nand U24501 (N_24501,N_21699,N_22305);
xnor U24502 (N_24502,N_21982,N_23768);
nand U24503 (N_24503,N_22299,N_21183);
or U24504 (N_24504,N_21580,N_23963);
nor U24505 (N_24505,N_21841,N_23093);
nand U24506 (N_24506,N_22271,N_23703);
nor U24507 (N_24507,N_23770,N_23734);
nand U24508 (N_24508,N_23458,N_23328);
and U24509 (N_24509,N_22168,N_21253);
nor U24510 (N_24510,N_21260,N_22968);
and U24511 (N_24511,N_21330,N_21220);
nor U24512 (N_24512,N_22121,N_21215);
xnor U24513 (N_24513,N_23349,N_23797);
and U24514 (N_24514,N_23321,N_22551);
and U24515 (N_24515,N_22025,N_23027);
or U24516 (N_24516,N_22008,N_23599);
nor U24517 (N_24517,N_23748,N_23236);
and U24518 (N_24518,N_23307,N_22946);
and U24519 (N_24519,N_21324,N_23422);
and U24520 (N_24520,N_22259,N_23691);
nand U24521 (N_24521,N_23989,N_23026);
nand U24522 (N_24522,N_23854,N_23529);
nor U24523 (N_24523,N_22089,N_21782);
xor U24524 (N_24524,N_22171,N_21329);
and U24525 (N_24525,N_22049,N_21375);
nor U24526 (N_24526,N_21029,N_22461);
and U24527 (N_24527,N_23844,N_23695);
or U24528 (N_24528,N_21755,N_23272);
or U24529 (N_24529,N_21608,N_21493);
and U24530 (N_24530,N_23229,N_23785);
and U24531 (N_24531,N_22346,N_23964);
and U24532 (N_24532,N_22427,N_21170);
nor U24533 (N_24533,N_22224,N_22211);
xnor U24534 (N_24534,N_23044,N_22921);
or U24535 (N_24535,N_21312,N_23746);
or U24536 (N_24536,N_22366,N_21381);
nand U24537 (N_24537,N_23594,N_23618);
or U24538 (N_24538,N_23648,N_21107);
and U24539 (N_24539,N_22926,N_22654);
or U24540 (N_24540,N_23455,N_23384);
xor U24541 (N_24541,N_22395,N_21696);
nor U24542 (N_24542,N_23598,N_21316);
nor U24543 (N_24543,N_23430,N_23322);
nand U24544 (N_24544,N_22789,N_23263);
and U24545 (N_24545,N_22748,N_23101);
and U24546 (N_24546,N_21617,N_22939);
nor U24547 (N_24547,N_22660,N_23834);
and U24548 (N_24548,N_22572,N_23288);
xor U24549 (N_24549,N_21681,N_21051);
nor U24550 (N_24550,N_21185,N_23040);
and U24551 (N_24551,N_22780,N_22501);
nor U24552 (N_24552,N_23897,N_21013);
nor U24553 (N_24553,N_23795,N_21738);
or U24554 (N_24554,N_21860,N_22510);
nor U24555 (N_24555,N_22908,N_22571);
nor U24556 (N_24556,N_23779,N_21618);
nor U24557 (N_24557,N_21683,N_21943);
xnor U24558 (N_24558,N_21300,N_21512);
and U24559 (N_24559,N_21418,N_22524);
nand U24560 (N_24560,N_22189,N_21648);
nand U24561 (N_24561,N_22671,N_23124);
and U24562 (N_24562,N_22663,N_22538);
and U24563 (N_24563,N_21886,N_21613);
or U24564 (N_24564,N_22608,N_21704);
and U24565 (N_24565,N_23056,N_22002);
and U24566 (N_24566,N_22235,N_23796);
nor U24567 (N_24567,N_23714,N_23148);
xnor U24568 (N_24568,N_23016,N_22458);
nand U24569 (N_24569,N_22157,N_23629);
and U24570 (N_24570,N_22261,N_21453);
or U24571 (N_24571,N_23159,N_22840);
or U24572 (N_24572,N_22557,N_21893);
or U24573 (N_24573,N_21728,N_23338);
nor U24574 (N_24574,N_22688,N_21680);
or U24575 (N_24575,N_23636,N_22728);
nand U24576 (N_24576,N_21825,N_22042);
and U24577 (N_24577,N_21344,N_22219);
nor U24578 (N_24578,N_23316,N_22734);
nand U24579 (N_24579,N_21795,N_21582);
nand U24580 (N_24580,N_21392,N_21599);
or U24581 (N_24581,N_23189,N_21913);
and U24582 (N_24582,N_23949,N_21690);
nand U24583 (N_24583,N_22897,N_21263);
and U24584 (N_24584,N_21273,N_23863);
nand U24585 (N_24585,N_23438,N_21909);
nor U24586 (N_24586,N_21632,N_22726);
nand U24587 (N_24587,N_21106,N_22809);
and U24588 (N_24588,N_23704,N_22520);
or U24589 (N_24589,N_23476,N_23873);
nand U24590 (N_24590,N_21566,N_22280);
nand U24591 (N_24591,N_21204,N_23239);
nor U24592 (N_24592,N_21596,N_23982);
nor U24593 (N_24593,N_21551,N_22767);
nand U24594 (N_24594,N_23603,N_23822);
xnor U24595 (N_24595,N_21414,N_23621);
xor U24596 (N_24596,N_21480,N_22295);
nand U24597 (N_24597,N_22786,N_22075);
nand U24598 (N_24598,N_22138,N_21397);
and U24599 (N_24599,N_21439,N_23513);
nor U24600 (N_24600,N_22383,N_23358);
nand U24601 (N_24601,N_21058,N_23503);
nor U24602 (N_24602,N_22912,N_23142);
or U24603 (N_24603,N_23998,N_22178);
or U24604 (N_24604,N_23567,N_22371);
or U24605 (N_24605,N_21657,N_21033);
nor U24606 (N_24606,N_23976,N_22009);
or U24607 (N_24607,N_22314,N_23904);
and U24608 (N_24608,N_21092,N_23898);
or U24609 (N_24609,N_21308,N_22298);
and U24610 (N_24610,N_22446,N_23528);
nand U24611 (N_24611,N_21374,N_21946);
nand U24612 (N_24612,N_21082,N_23790);
and U24613 (N_24613,N_21071,N_21662);
xnor U24614 (N_24614,N_22692,N_22658);
nor U24615 (N_24615,N_23905,N_22754);
nand U24616 (N_24616,N_22445,N_21922);
nand U24617 (N_24617,N_22798,N_23924);
nor U24618 (N_24618,N_21048,N_22296);
nor U24619 (N_24619,N_23638,N_22228);
xor U24620 (N_24620,N_22464,N_21080);
xnor U24621 (N_24621,N_21981,N_22659);
xor U24622 (N_24622,N_23596,N_22468);
and U24623 (N_24623,N_21513,N_21129);
or U24624 (N_24624,N_22472,N_22723);
nand U24625 (N_24625,N_22724,N_22005);
and U24626 (N_24626,N_22386,N_21258);
nand U24627 (N_24627,N_21389,N_22335);
nor U24628 (N_24628,N_21558,N_22620);
or U24629 (N_24629,N_21754,N_22203);
or U24630 (N_24630,N_22588,N_23756);
nor U24631 (N_24631,N_22648,N_22128);
and U24632 (N_24632,N_23820,N_21964);
nor U24633 (N_24633,N_22710,N_22788);
and U24634 (N_24634,N_23918,N_21457);
xnor U24635 (N_24635,N_22626,N_23885);
nand U24636 (N_24636,N_21481,N_23635);
or U24637 (N_24637,N_21603,N_22258);
nand U24638 (N_24638,N_22674,N_23121);
and U24639 (N_24639,N_23417,N_21461);
xnor U24640 (N_24640,N_21342,N_21067);
nor U24641 (N_24641,N_22233,N_21555);
nand U24642 (N_24642,N_21387,N_23330);
or U24643 (N_24643,N_21328,N_23169);
or U24644 (N_24644,N_21052,N_23277);
nor U24645 (N_24645,N_21562,N_23815);
and U24646 (N_24646,N_23847,N_21848);
and U24647 (N_24647,N_22067,N_23423);
nor U24648 (N_24648,N_23592,N_23579);
or U24649 (N_24649,N_23098,N_23839);
xor U24650 (N_24650,N_23356,N_23201);
xnor U24651 (N_24651,N_21833,N_21075);
nor U24652 (N_24652,N_21032,N_23303);
nand U24653 (N_24653,N_22118,N_22539);
xor U24654 (N_24654,N_23400,N_23095);
and U24655 (N_24655,N_22012,N_22212);
and U24656 (N_24656,N_22852,N_22558);
nand U24657 (N_24657,N_21965,N_23980);
nand U24658 (N_24658,N_23497,N_22987);
xor U24659 (N_24659,N_21179,N_22126);
nand U24660 (N_24660,N_22412,N_21378);
nor U24661 (N_24661,N_22815,N_21138);
xnor U24662 (N_24662,N_22175,N_23517);
or U24663 (N_24663,N_23194,N_21450);
xnor U24664 (N_24664,N_22927,N_21746);
or U24665 (N_24665,N_22409,N_22826);
nor U24666 (N_24666,N_21631,N_23901);
nor U24667 (N_24667,N_22795,N_21577);
and U24668 (N_24668,N_21959,N_22511);
and U24669 (N_24669,N_22232,N_23329);
or U24670 (N_24670,N_21533,N_21498);
nand U24671 (N_24671,N_22028,N_21719);
and U24672 (N_24672,N_21350,N_22687);
or U24673 (N_24673,N_23331,N_21762);
and U24674 (N_24674,N_23808,N_23436);
or U24675 (N_24675,N_21861,N_21854);
nor U24676 (N_24676,N_21876,N_23752);
nand U24677 (N_24677,N_22210,N_21672);
or U24678 (N_24678,N_22751,N_23769);
nand U24679 (N_24679,N_23060,N_22385);
or U24680 (N_24680,N_22497,N_23219);
or U24681 (N_24681,N_23224,N_21180);
or U24682 (N_24682,N_21061,N_23432);
nand U24683 (N_24683,N_21113,N_22811);
nand U24684 (N_24684,N_23003,N_21056);
or U24685 (N_24685,N_22881,N_22230);
nand U24686 (N_24686,N_23740,N_21595);
nand U24687 (N_24687,N_21379,N_23197);
and U24688 (N_24688,N_23246,N_22275);
and U24689 (N_24689,N_21060,N_22207);
nor U24690 (N_24690,N_22675,N_23656);
xor U24691 (N_24691,N_21804,N_22982);
xnor U24692 (N_24692,N_21628,N_23712);
nand U24693 (N_24693,N_23550,N_22639);
nand U24694 (N_24694,N_23069,N_23317);
nor U24695 (N_24695,N_22431,N_22890);
or U24696 (N_24696,N_23586,N_22104);
nand U24697 (N_24697,N_22043,N_22093);
nand U24698 (N_24698,N_23230,N_21235);
nand U24699 (N_24699,N_23782,N_22240);
or U24700 (N_24700,N_23271,N_22419);
and U24701 (N_24701,N_23566,N_21063);
or U24702 (N_24702,N_23344,N_21799);
nor U24703 (N_24703,N_22594,N_22155);
nor U24704 (N_24704,N_22490,N_21209);
xor U24705 (N_24705,N_23876,N_21290);
and U24706 (N_24706,N_22380,N_22508);
nand U24707 (N_24707,N_22869,N_22760);
and U24708 (N_24708,N_21353,N_22399);
xor U24709 (N_24709,N_22315,N_21644);
xnor U24710 (N_24710,N_22281,N_23465);
xor U24711 (N_24711,N_21839,N_22838);
nand U24712 (N_24712,N_21024,N_22992);
nand U24713 (N_24713,N_23819,N_21759);
or U24714 (N_24714,N_22544,N_22215);
and U24715 (N_24715,N_22656,N_22065);
or U24716 (N_24716,N_23318,N_23448);
and U24717 (N_24717,N_22441,N_21611);
nand U24718 (N_24718,N_22606,N_22918);
xnor U24719 (N_24719,N_23135,N_21926);
or U24720 (N_24720,N_21885,N_21896);
nor U24721 (N_24721,N_23158,N_22438);
xor U24722 (N_24722,N_22717,N_22192);
nand U24723 (N_24723,N_21074,N_21279);
or U24724 (N_24724,N_22830,N_22106);
xnor U24725 (N_24725,N_22793,N_22686);
or U24726 (N_24726,N_21875,N_23868);
or U24727 (N_24727,N_22629,N_21707);
xnor U24728 (N_24728,N_21373,N_23405);
or U24729 (N_24729,N_23842,N_21930);
nand U24730 (N_24730,N_23615,N_22683);
nor U24731 (N_24731,N_23470,N_22742);
nand U24732 (N_24732,N_21171,N_21983);
or U24733 (N_24733,N_23614,N_21539);
and U24734 (N_24734,N_21968,N_22518);
xor U24735 (N_24735,N_23047,N_23128);
and U24736 (N_24736,N_23948,N_21083);
nand U24737 (N_24737,N_21665,N_22653);
or U24738 (N_24738,N_21162,N_21702);
nand U24739 (N_24739,N_23190,N_23453);
nand U24740 (N_24740,N_21610,N_21579);
or U24741 (N_24741,N_21521,N_22585);
and U24742 (N_24742,N_22768,N_21093);
nor U24743 (N_24743,N_23655,N_21231);
or U24744 (N_24744,N_22485,N_21009);
xnor U24745 (N_24745,N_23780,N_22943);
nor U24746 (N_24746,N_21677,N_22217);
nor U24747 (N_24747,N_23063,N_23200);
nand U24748 (N_24748,N_21831,N_22609);
or U24749 (N_24749,N_22615,N_21412);
and U24750 (N_24750,N_22195,N_21295);
nor U24751 (N_24751,N_21408,N_22925);
or U24752 (N_24752,N_21864,N_22602);
nor U24753 (N_24753,N_22123,N_22456);
and U24754 (N_24754,N_23106,N_21615);
and U24755 (N_24755,N_21523,N_22347);
nand U24756 (N_24756,N_22344,N_21256);
nor U24757 (N_24757,N_21246,N_22611);
or U24758 (N_24758,N_23226,N_23682);
nor U24759 (N_24759,N_22473,N_23671);
xnor U24760 (N_24760,N_23917,N_23828);
or U24761 (N_24761,N_23727,N_21776);
and U24762 (N_24762,N_21989,N_21110);
nor U24763 (N_24763,N_21413,N_21166);
or U24764 (N_24764,N_23140,N_23327);
nand U24765 (N_24765,N_22750,N_23968);
and U24766 (N_24766,N_22145,N_23974);
nand U24767 (N_24767,N_21410,N_21261);
and U24768 (N_24768,N_21688,N_22208);
or U24769 (N_24769,N_21464,N_23572);
and U24770 (N_24770,N_22070,N_23827);
and U24771 (N_24771,N_23161,N_22995);
nand U24772 (N_24772,N_22090,N_21589);
and U24773 (N_24773,N_22810,N_22194);
nor U24774 (N_24774,N_22253,N_23957);
nor U24775 (N_24775,N_23895,N_21252);
or U24776 (N_24776,N_23837,N_22499);
nor U24777 (N_24777,N_22550,N_21937);
and U24778 (N_24778,N_23256,N_23861);
or U24779 (N_24779,N_23690,N_23926);
xnor U24780 (N_24780,N_21366,N_22736);
and U24781 (N_24781,N_22889,N_21435);
and U24782 (N_24782,N_22624,N_23595);
nor U24783 (N_24783,N_23499,N_22578);
and U24784 (N_24784,N_21587,N_23083);
or U24785 (N_24785,N_23549,N_22781);
or U24786 (N_24786,N_21165,N_21064);
nand U24787 (N_24787,N_23777,N_21456);
nor U24788 (N_24788,N_22756,N_22424);
and U24789 (N_24789,N_22527,N_23658);
nor U24790 (N_24790,N_23247,N_22833);
nor U24791 (N_24791,N_23721,N_23160);
nand U24792 (N_24792,N_22613,N_22447);
nand U24793 (N_24793,N_23800,N_21299);
nand U24794 (N_24794,N_22537,N_23679);
or U24795 (N_24795,N_21917,N_22449);
or U24796 (N_24796,N_23129,N_23209);
nor U24797 (N_24797,N_22785,N_21939);
and U24798 (N_24798,N_22421,N_23004);
nand U24799 (N_24799,N_22476,N_22752);
or U24800 (N_24800,N_22828,N_21940);
or U24801 (N_24801,N_22372,N_23977);
xor U24802 (N_24802,N_22804,N_21954);
nor U24803 (N_24803,N_23620,N_22030);
xnor U24804 (N_24804,N_22862,N_22282);
or U24805 (N_24805,N_21921,N_21225);
or U24806 (N_24806,N_23778,N_23676);
and U24807 (N_24807,N_22220,N_23342);
and U24808 (N_24808,N_21377,N_23943);
nand U24809 (N_24809,N_23441,N_21652);
nand U24810 (N_24810,N_22563,N_22568);
nand U24811 (N_24811,N_21419,N_21336);
nand U24812 (N_24812,N_21193,N_22679);
nand U24813 (N_24813,N_23587,N_22377);
nand U24814 (N_24814,N_22018,N_22628);
nand U24815 (N_24815,N_23393,N_21686);
or U24816 (N_24816,N_22700,N_23281);
and U24817 (N_24817,N_22142,N_23617);
xnor U24818 (N_24818,N_22846,N_21391);
nor U24819 (N_24819,N_21354,N_23312);
and U24820 (N_24820,N_21200,N_22364);
nor U24821 (N_24821,N_21111,N_22410);
or U24822 (N_24822,N_22213,N_21726);
and U24823 (N_24823,N_21999,N_23685);
nor U24824 (N_24824,N_22820,N_22715);
or U24825 (N_24825,N_23261,N_23653);
nand U24826 (N_24826,N_22837,N_21372);
nand U24827 (N_24827,N_21871,N_22779);
or U24828 (N_24828,N_23195,N_21315);
or U24829 (N_24829,N_23991,N_21724);
nor U24830 (N_24830,N_21536,N_21671);
nand U24831 (N_24831,N_21361,N_21059);
nand U24832 (N_24832,N_22735,N_21249);
xor U24833 (N_24833,N_22303,N_22504);
and U24834 (N_24834,N_21137,N_21996);
and U24835 (N_24835,N_21638,N_22638);
and U24836 (N_24836,N_22962,N_23018);
or U24837 (N_24837,N_22884,N_22975);
xor U24838 (N_24838,N_22001,N_22216);
nand U24839 (N_24839,N_23029,N_23484);
xnor U24840 (N_24840,N_22740,N_23717);
and U24841 (N_24841,N_21201,N_21581);
nor U24842 (N_24842,N_23564,N_23927);
or U24843 (N_24843,N_21643,N_22316);
nor U24844 (N_24844,N_22218,N_21900);
or U24845 (N_24845,N_21189,N_23787);
nor U24846 (N_24846,N_22894,N_21607);
nor U24847 (N_24847,N_23242,N_21918);
nand U24848 (N_24848,N_22807,N_21030);
and U24849 (N_24849,N_21747,N_21117);
nand U24850 (N_24850,N_23879,N_23799);
and U24851 (N_24851,N_23582,N_21655);
nor U24852 (N_24852,N_23642,N_21054);
nor U24853 (N_24853,N_21043,N_23771);
xnor U24854 (N_24854,N_23575,N_23127);
nand U24855 (N_24855,N_21213,N_21343);
and U24856 (N_24856,N_22988,N_22131);
nand U24857 (N_24857,N_22351,N_23997);
nand U24858 (N_24858,N_22848,N_23802);
and U24859 (N_24859,N_23446,N_23351);
nor U24860 (N_24860,N_22600,N_22081);
nand U24861 (N_24861,N_21715,N_22307);
nor U24862 (N_24862,N_22514,N_23363);
or U24863 (N_24863,N_22165,N_21425);
and U24864 (N_24864,N_22141,N_23776);
nand U24865 (N_24865,N_23252,N_21869);
and U24866 (N_24866,N_22069,N_23510);
nor U24867 (N_24867,N_21155,N_21910);
and U24868 (N_24868,N_22586,N_22670);
or U24869 (N_24869,N_23019,N_23440);
xor U24870 (N_24870,N_22579,N_21130);
nand U24871 (N_24871,N_23911,N_23394);
and U24872 (N_24872,N_22506,N_23466);
xnor U24873 (N_24873,N_21192,N_23647);
and U24874 (N_24874,N_23698,N_23686);
or U24875 (N_24875,N_22255,N_21027);
and U24876 (N_24876,N_21281,N_21288);
and U24877 (N_24877,N_22871,N_21360);
and U24878 (N_24878,N_22227,N_22630);
nand U24879 (N_24879,N_23945,N_22393);
or U24880 (N_24880,N_21427,N_23255);
nor U24881 (N_24881,N_21401,N_23942);
or U24882 (N_24882,N_22048,N_23912);
xor U24883 (N_24883,N_23136,N_22938);
and U24884 (N_24884,N_22154,N_22435);
xnor U24885 (N_24885,N_23992,N_23774);
and U24886 (N_24886,N_21803,N_22573);
nand U24887 (N_24887,N_23483,N_21460);
and U24888 (N_24888,N_22357,N_23511);
xnor U24889 (N_24889,N_21276,N_23104);
nor U24890 (N_24890,N_23956,N_23693);
and U24891 (N_24891,N_21206,N_23086);
and U24892 (N_24892,N_23501,N_21169);
and U24893 (N_24893,N_22078,N_23109);
nand U24894 (N_24894,N_23678,N_23697);
nand U24895 (N_24895,N_21530,N_22097);
and U24896 (N_24896,N_22060,N_23232);
nor U24897 (N_24897,N_23817,N_23108);
or U24898 (N_24898,N_21011,N_21062);
nand U24899 (N_24899,N_21716,N_21912);
nand U24900 (N_24900,N_22650,N_21228);
nand U24901 (N_24901,N_23308,N_23238);
and U24902 (N_24902,N_23899,N_22707);
nor U24903 (N_24903,N_22268,N_22963);
or U24904 (N_24904,N_23315,N_21416);
nor U24905 (N_24905,N_23581,N_23185);
or U24906 (N_24906,N_22480,N_22854);
and U24907 (N_24907,N_23623,N_23881);
or U24908 (N_24908,N_22566,N_21744);
and U24909 (N_24909,N_23289,N_21151);
nor U24910 (N_24910,N_21807,N_22312);
and U24911 (N_24911,N_21199,N_23556);
nand U24912 (N_24912,N_21184,N_23531);
and U24913 (N_24913,N_22231,N_21604);
nor U24914 (N_24914,N_23397,N_21792);
nor U24915 (N_24915,N_22290,N_22940);
nand U24916 (N_24916,N_21190,N_22288);
nand U24917 (N_24917,N_23610,N_22644);
xnor U24918 (N_24918,N_21055,N_21933);
and U24919 (N_24919,N_23481,N_21492);
and U24920 (N_24920,N_22635,N_22467);
or U24921 (N_24921,N_21023,N_21635);
nand U24922 (N_24922,N_21883,N_21478);
nand U24923 (N_24923,N_23105,N_21944);
or U24924 (N_24924,N_21623,N_22842);
and U24925 (N_24925,N_22966,N_22109);
nand U24926 (N_24926,N_23381,N_21627);
or U24927 (N_24927,N_22993,N_21388);
and U24928 (N_24928,N_21040,N_21560);
nor U24929 (N_24929,N_23652,N_23137);
nand U24930 (N_24930,N_23630,N_23211);
nand U24931 (N_24931,N_23874,N_22243);
xnor U24932 (N_24932,N_21730,N_23377);
and U24933 (N_24933,N_21774,N_23326);
and U24934 (N_24934,N_23410,N_21709);
and U24935 (N_24935,N_21448,N_23419);
and U24936 (N_24936,N_22323,N_23275);
nor U24937 (N_24937,N_22382,N_23496);
and U24938 (N_24938,N_21748,N_23641);
and U24939 (N_24939,N_21911,N_23362);
nor U24940 (N_24940,N_21575,N_23102);
or U24941 (N_24941,N_21386,N_23766);
and U24942 (N_24942,N_22716,N_22636);
or U24943 (N_24943,N_21469,N_23449);
nand U24944 (N_24944,N_23520,N_21508);
nor U24945 (N_24945,N_22094,N_21057);
and U24946 (N_24946,N_21997,N_21482);
and U24947 (N_24947,N_22843,N_22595);
or U24948 (N_24948,N_21805,N_21633);
nor U24949 (N_24949,N_21098,N_23887);
nand U24950 (N_24950,N_22379,N_21161);
nand U24951 (N_24951,N_23460,N_21664);
and U24952 (N_24952,N_21740,N_22749);
or U24953 (N_24953,N_23173,N_22167);
and U24954 (N_24954,N_22697,N_21505);
nand U24955 (N_24955,N_23096,N_21028);
and U24956 (N_24956,N_21641,N_23054);
nand U24957 (N_24957,N_23741,N_21812);
nand U24958 (N_24958,N_23547,N_22247);
nor U24959 (N_24959,N_21104,N_23477);
nand U24960 (N_24960,N_21124,N_22164);
nand U24961 (N_24961,N_23555,N_22417);
nand U24962 (N_24962,N_21501,N_23669);
and U24963 (N_24963,N_23959,N_22453);
or U24964 (N_24964,N_23407,N_22439);
nor U24965 (N_24965,N_22796,N_23807);
and U24966 (N_24966,N_21430,N_21960);
nor U24967 (N_24967,N_22313,N_23126);
nor U24968 (N_24968,N_22214,N_22193);
nor U24969 (N_24969,N_21857,N_21793);
nor U24970 (N_24970,N_22769,N_23285);
nand U24971 (N_24971,N_23660,N_23938);
nor U24972 (N_24972,N_22507,N_22452);
nand U24973 (N_24973,N_21932,N_22122);
or U24974 (N_24974,N_23399,N_23046);
xnor U24975 (N_24975,N_23794,N_22721);
and U24976 (N_24976,N_21085,N_22932);
and U24977 (N_24977,N_21739,N_23612);
nand U24978 (N_24978,N_21163,N_23270);
and U24979 (N_24979,N_22875,N_21234);
or U24980 (N_24980,N_21466,N_21532);
or U24981 (N_24981,N_23931,N_22589);
nor U24982 (N_24982,N_23871,N_21420);
nand U24983 (N_24983,N_21194,N_22976);
or U24984 (N_24984,N_22058,N_23929);
and U24985 (N_24985,N_23569,N_21514);
nor U24986 (N_24986,N_22050,N_22562);
nor U24987 (N_24987,N_21880,N_22753);
and U24988 (N_24988,N_21866,N_21842);
nor U24989 (N_24989,N_23254,N_23012);
and U24990 (N_24990,N_21128,N_22394);
nor U24991 (N_24991,N_22059,N_21974);
nand U24992 (N_24992,N_21259,N_21708);
and U24993 (N_24993,N_21443,N_23087);
or U24994 (N_24994,N_22116,N_23390);
and U24995 (N_24995,N_22156,N_22486);
xor U24996 (N_24996,N_22375,N_21895);
nand U24997 (N_24997,N_21380,N_21477);
and U24998 (N_24998,N_22633,N_21682);
xor U24999 (N_24999,N_23052,N_22318);
or U25000 (N_25000,N_21198,N_21045);
nand U25001 (N_25001,N_22819,N_22170);
nor U25002 (N_25002,N_22657,N_21801);
nand U25003 (N_25003,N_22543,N_21337);
nor U25004 (N_25004,N_23380,N_21097);
nor U25005 (N_25005,N_21087,N_21112);
xor U25006 (N_25006,N_21341,N_21544);
nor U25007 (N_25007,N_22930,N_23103);
and U25008 (N_25008,N_23689,N_23738);
or U25009 (N_25009,N_21149,N_23180);
nor U25010 (N_25010,N_21780,N_21670);
and U25011 (N_25011,N_21723,N_21908);
xor U25012 (N_25012,N_23473,N_21222);
or U25013 (N_25013,N_21785,N_22052);
or U25014 (N_25014,N_21426,N_22270);
nand U25015 (N_25015,N_21811,N_22505);
xor U25016 (N_25016,N_22204,N_22835);
and U25017 (N_25017,N_21969,N_21763);
or U25018 (N_25018,N_21227,N_22746);
or U25019 (N_25019,N_22053,N_21313);
xor U25020 (N_25020,N_23075,N_23364);
nor U25021 (N_25021,N_21332,N_22590);
nand U25022 (N_25022,N_21287,N_21266);
or U25023 (N_25023,N_22054,N_22086);
nor U25024 (N_25024,N_21591,N_21967);
nor U25025 (N_25025,N_22262,N_23266);
and U25026 (N_25026,N_21221,N_23258);
nor U25027 (N_25027,N_23235,N_22999);
nand U25028 (N_25028,N_21588,N_21188);
or U25029 (N_25029,N_22851,N_23687);
or U25030 (N_25030,N_22015,N_21769);
nand U25031 (N_25031,N_21139,N_22339);
or U25032 (N_25032,N_22850,N_23084);
nor U25033 (N_25033,N_22110,N_21706);
and U25034 (N_25034,N_23798,N_21257);
or U25035 (N_25035,N_23265,N_22153);
or U25036 (N_25036,N_23306,N_23829);
nor U25037 (N_25037,N_22016,N_21936);
and U25038 (N_25038,N_22390,N_23961);
nor U25039 (N_25039,N_23878,N_21837);
or U25040 (N_25040,N_23788,N_22483);
nand U25041 (N_25041,N_23824,N_21768);
nor U25042 (N_25042,N_21667,N_21547);
and U25043 (N_25043,N_22512,N_22565);
nand U25044 (N_25044,N_23561,N_22063);
nand U25045 (N_25045,N_21196,N_21405);
and U25046 (N_25046,N_23867,N_23113);
nor U25047 (N_25047,N_21044,N_23403);
nor U25048 (N_25048,N_22384,N_21065);
and U25049 (N_25049,N_21584,N_22105);
nor U25050 (N_25050,N_22603,N_23182);
or U25051 (N_25051,N_21697,N_22783);
or U25052 (N_25052,N_23670,N_23823);
and U25053 (N_25053,N_22745,N_22642);
and U25054 (N_25054,N_22374,N_21267);
nand U25055 (N_25055,N_22432,N_22813);
nand U25056 (N_25056,N_22873,N_22763);
or U25057 (N_25057,N_22237,N_22676);
or U25058 (N_25058,N_21358,N_23468);
or U25059 (N_25059,N_23478,N_22463);
nor U25060 (N_25060,N_22941,N_21727);
nand U25061 (N_25061,N_23739,N_23157);
or U25062 (N_25062,N_21262,N_23753);
nor U25063 (N_25063,N_23345,N_21333);
nor U25064 (N_25064,N_22694,N_22720);
nand U25065 (N_25065,N_22019,N_22184);
nand U25066 (N_25066,N_23166,N_22618);
xor U25067 (N_25067,N_22342,N_22556);
and U25068 (N_25068,N_21291,N_21500);
nand U25069 (N_25069,N_23184,N_23751);
xnor U25070 (N_25070,N_22354,N_23907);
and U25071 (N_25071,N_21178,N_22983);
and U25072 (N_25072,N_23910,N_22849);
nand U25073 (N_25073,N_21240,N_23164);
or U25074 (N_25074,N_23577,N_21434);
nor U25075 (N_25075,N_21278,N_21303);
nor U25076 (N_25076,N_23554,N_21597);
nand U25077 (N_25077,N_21735,N_21563);
or U25078 (N_25078,N_21365,N_23428);
xor U25079 (N_25079,N_21210,N_23427);
nor U25080 (N_25080,N_22732,N_22113);
or U25081 (N_25081,N_23903,N_23506);
or U25082 (N_25082,N_23972,N_22284);
nor U25083 (N_25083,N_23607,N_21338);
nand U25084 (N_25084,N_22977,N_23684);
and U25085 (N_25085,N_23398,N_23294);
nor U25086 (N_25086,N_23979,N_23605);
nand U25087 (N_25087,N_21421,N_21250);
or U25088 (N_25088,N_22868,N_22283);
or U25089 (N_25089,N_21003,N_23065);
or U25090 (N_25090,N_21534,N_22771);
and U25091 (N_25091,N_22391,N_23548);
nor U25092 (N_25092,N_22308,N_22727);
or U25093 (N_25093,N_23051,N_21931);
xnor U25094 (N_25094,N_21126,N_21598);
or U25095 (N_25095,N_22964,N_21822);
and U25096 (N_25096,N_21490,N_22130);
and U25097 (N_25097,N_21892,N_21499);
nand U25098 (N_25098,N_21784,N_21008);
or U25099 (N_25099,N_22479,N_21168);
or U25100 (N_25100,N_21961,N_23141);
nand U25101 (N_25101,N_21781,N_23616);
nor U25102 (N_25102,N_21422,N_23590);
nand U25103 (N_25103,N_23457,N_21764);
and U25104 (N_25104,N_21136,N_23074);
xor U25105 (N_25105,N_23651,N_21522);
nand U25106 (N_25106,N_22337,N_21417);
nand U25107 (N_25107,N_23836,N_22797);
or U25108 (N_25108,N_22367,N_21385);
and U25109 (N_25109,N_21570,N_22536);
nand U25110 (N_25110,N_23366,N_22241);
nand U25111 (N_25111,N_22428,N_22188);
nor U25112 (N_25112,N_21038,N_23276);
and U25113 (N_25113,N_21415,N_23248);
xnor U25114 (N_25114,N_21079,N_22698);
or U25115 (N_25115,N_21309,N_22443);
and U25116 (N_25116,N_21674,N_23602);
and U25117 (N_25117,N_22331,N_23414);
xor U25118 (N_25118,N_23524,N_22095);
nor U25119 (N_25119,N_21621,N_22895);
nor U25120 (N_25120,N_22949,N_22802);
or U25121 (N_25121,N_23519,N_23452);
and U25122 (N_25122,N_23107,N_21583);
nand U25123 (N_25123,N_22205,N_22440);
and U25124 (N_25124,N_21322,N_23165);
nand U25125 (N_25125,N_21636,N_22129);
and U25126 (N_25126,N_21095,N_22117);
nand U25127 (N_25127,N_22265,N_23006);
or U25128 (N_25128,N_21668,N_22818);
nor U25129 (N_25129,N_23987,N_21105);
nand U25130 (N_25130,N_21382,N_22373);
and U25131 (N_25131,N_23805,N_21475);
nor U25132 (N_25132,N_22841,N_21116);
or U25133 (N_25133,N_23526,N_21863);
nor U25134 (N_25134,N_21899,N_23461);
nand U25135 (N_25135,N_21103,N_22163);
and U25136 (N_25136,N_21473,N_21847);
and U25137 (N_25137,N_22643,N_21711);
nand U25138 (N_25138,N_22125,N_21543);
nand U25139 (N_25139,N_23928,N_22493);
nor U25140 (N_25140,N_22832,N_21479);
nor U25141 (N_25141,N_23609,N_23843);
and U25142 (N_25142,N_23558,N_21590);
nand U25143 (N_25143,N_21535,N_22139);
nor U25144 (N_25144,N_22684,N_23539);
or U25145 (N_25145,N_22152,N_23490);
nor U25146 (N_25146,N_22766,N_23688);
nand U25147 (N_25147,N_21808,N_23613);
nand U25148 (N_25148,N_22791,N_21400);
xnor U25149 (N_25149,N_23067,N_22669);
or U25150 (N_25150,N_22133,N_22310);
nor U25151 (N_25151,N_23061,N_21541);
or U25152 (N_25152,N_21957,N_23204);
xnor U25153 (N_25153,N_21986,N_21411);
xnor U25154 (N_25154,N_22991,N_23702);
and U25155 (N_25155,N_22041,N_21527);
and U25156 (N_25156,N_23532,N_22741);
nor U25157 (N_25157,N_23222,N_23645);
and U25158 (N_25158,N_23192,N_22952);
nand U25159 (N_25159,N_21049,N_21494);
nor U25160 (N_25160,N_21528,N_23857);
and U25161 (N_25161,N_23694,N_23784);
nor U25162 (N_25162,N_23005,N_21877);
nand U25163 (N_25163,N_22531,N_21624);
nor U25164 (N_25164,N_22256,N_21232);
nand U25165 (N_25165,N_22405,N_21404);
and U25166 (N_25166,N_22032,N_22425);
nor U25167 (N_25167,N_21109,N_21172);
nor U25168 (N_25168,N_23474,N_22392);
or U25169 (N_25169,N_23070,N_23889);
nor U25170 (N_25170,N_21019,N_22350);
or U25171 (N_25171,N_21447,N_22744);
nor U25172 (N_25172,N_23352,N_21767);
or U25173 (N_25173,N_23297,N_21980);
nand U25174 (N_25174,N_23932,N_23534);
nor U25175 (N_25175,N_23495,N_23626);
nand U25176 (N_25176,N_21531,N_23628);
or U25177 (N_25177,N_23139,N_22739);
or U25178 (N_25178,N_22560,N_22907);
or U25179 (N_25179,N_22583,N_23372);
or U25180 (N_25180,N_23890,N_22816);
or U25181 (N_25181,N_21914,N_22278);
or U25182 (N_25182,N_23990,N_22860);
nor U25183 (N_25183,N_21685,N_23472);
or U25184 (N_25184,N_23203,N_22922);
and U25185 (N_25185,N_21211,N_21998);
and U25186 (N_25186,N_23922,N_21187);
nor U25187 (N_25187,N_21548,N_22730);
xor U25188 (N_25188,N_21159,N_23020);
nor U25189 (N_25189,N_22596,N_23947);
and U25190 (N_25190,N_22604,N_22144);
nand U25191 (N_25191,N_23781,N_22929);
nand U25192 (N_25192,N_22451,N_21894);
xnor U25193 (N_25193,N_21881,N_23090);
and U25194 (N_25194,N_23176,N_23580);
xor U25195 (N_25195,N_21244,N_22119);
and U25196 (N_25196,N_22567,N_23930);
and U25197 (N_25197,N_22103,N_21694);
nand U25198 (N_25198,N_22029,N_23757);
nand U25199 (N_25199,N_23668,N_23171);
nand U25200 (N_25200,N_22149,N_23726);
or U25201 (N_25201,N_21005,N_21497);
nand U25202 (N_25202,N_22101,N_22866);
nand U25203 (N_25203,N_22920,N_23736);
nand U25204 (N_25204,N_23480,N_21684);
or U25205 (N_25205,N_21736,N_22368);
nor U25206 (N_25206,N_23437,N_22640);
or U25207 (N_25207,N_22548,N_21304);
nor U25208 (N_25208,N_22637,N_21955);
or U25209 (N_25209,N_22799,N_21878);
and U25210 (N_25210,N_22422,N_23162);
nand U25211 (N_25211,N_21817,N_22498);
or U25212 (N_25212,N_21296,N_23570);
or U25213 (N_25213,N_23340,N_23674);
nor U25214 (N_25214,N_23073,N_21718);
nor U25215 (N_25215,N_23291,N_22731);
nor U25216 (N_25216,N_22803,N_22876);
nor U25217 (N_25217,N_23713,N_23350);
nand U25218 (N_25218,N_22935,N_23310);
nand U25219 (N_25219,N_21821,N_21905);
and U25220 (N_25220,N_21217,N_23858);
or U25221 (N_25221,N_21844,N_22725);
or U25222 (N_25222,N_22782,N_23538);
and U25223 (N_25223,N_21663,N_23334);
or U25224 (N_25224,N_23485,N_22614);
and U25225 (N_25225,N_22865,N_23079);
nand U25226 (N_25226,N_22023,N_21470);
nor U25227 (N_25227,N_21550,N_23960);
nand U25228 (N_25228,N_21517,N_22297);
and U25229 (N_25229,N_23188,N_22812);
nor U25230 (N_25230,N_22978,N_22695);
nand U25231 (N_25231,N_23038,N_23773);
nand U25232 (N_25232,N_21218,N_23311);
and U25233 (N_25233,N_22667,N_23913);
or U25234 (N_25234,N_23664,N_23337);
or U25235 (N_25235,N_23112,N_22622);
nor U25236 (N_25236,N_23216,N_23845);
nor U25237 (N_25237,N_22980,N_22522);
and U25238 (N_25238,N_22755,N_23369);
nor U25239 (N_25239,N_21326,N_23144);
nand U25240 (N_25240,N_23251,N_22416);
nor U25241 (N_25241,N_23718,N_21788);
and U25242 (N_25242,N_23523,N_22306);
nor U25243 (N_25243,N_21140,N_22348);
or U25244 (N_25244,N_21714,N_21286);
or U25245 (N_25245,N_23119,N_23729);
or U25246 (N_25246,N_22775,N_22765);
xor U25247 (N_25247,N_21978,N_23469);
or U25248 (N_25248,N_21640,N_23361);
nor U25249 (N_25249,N_21150,N_21311);
or U25250 (N_25250,N_22559,N_22336);
or U25251 (N_25251,N_23167,N_23245);
and U25252 (N_25252,N_21749,N_21993);
or U25253 (N_25253,N_22891,N_21902);
and U25254 (N_25254,N_22099,N_21101);
nand U25255 (N_25255,N_21362,N_22183);
xnor U25256 (N_25256,N_21520,N_22582);
nor U25257 (N_25257,N_23962,N_22917);
or U25258 (N_25258,N_23715,N_21675);
nand U25259 (N_25259,N_21693,N_22369);
nand U25260 (N_25260,N_21212,N_21787);
xnor U25261 (N_25261,N_22523,N_23028);
xnor U25262 (N_25262,N_22471,N_23152);
or U25263 (N_25263,N_21431,N_21654);
and U25264 (N_25264,N_21897,N_21507);
nor U25265 (N_25265,N_21271,N_21121);
and U25266 (N_25266,N_22022,N_21084);
xor U25267 (N_25267,N_21270,N_23522);
or U25268 (N_25268,N_21007,N_23343);
nand U25269 (N_25269,N_22151,N_21476);
or U25270 (N_25270,N_22328,N_21691);
nand U25271 (N_25271,N_21695,N_21305);
or U25272 (N_25272,N_21368,N_23971);
nand U25273 (N_25273,N_23072,N_23243);
and U25274 (N_25274,N_23891,N_23804);
nand U25275 (N_25275,N_22607,N_22666);
or U25276 (N_25276,N_22064,N_23565);
nand U25277 (N_25277,N_23415,N_23909);
and U25278 (N_25278,N_21280,N_22301);
nand U25279 (N_25279,N_23259,N_23545);
nand U25280 (N_25280,N_22888,N_21593);
and U25281 (N_25281,N_21371,N_23416);
or U25282 (N_25282,N_23273,N_23092);
or U25283 (N_25283,N_22190,N_22111);
nor U25284 (N_25284,N_23934,N_21001);
nand U25285 (N_25285,N_22363,N_21394);
nand U25286 (N_25286,N_22933,N_21862);
xnor U25287 (N_25287,N_22020,N_21890);
and U25288 (N_25288,N_23392,N_22127);
xor U25289 (N_25289,N_22885,N_21072);
nand U25290 (N_25290,N_23388,N_22260);
nor U25291 (N_25291,N_22264,N_21592);
nor U25292 (N_25292,N_23492,N_22625);
nand U25293 (N_25293,N_22477,N_21700);
nand U25294 (N_25294,N_21758,N_21859);
nand U25295 (N_25295,N_22238,N_22770);
or U25296 (N_25296,N_23174,N_22234);
nor U25297 (N_25297,N_23313,N_22762);
nor U25298 (N_25298,N_21488,N_21777);
nor U25299 (N_25299,N_22176,N_22158);
nand U25300 (N_25300,N_21255,N_23264);
nor U25301 (N_25301,N_23585,N_23601);
xnor U25302 (N_25302,N_21889,N_23249);
nor U25303 (N_25303,N_21335,N_23325);
nor U25304 (N_25304,N_23301,N_22834);
and U25305 (N_25305,N_21182,N_22853);
nor U25306 (N_25306,N_22448,N_21506);
or U25307 (N_25307,N_22805,N_23830);
and U25308 (N_25308,N_21503,N_22279);
and U25309 (N_25309,N_22353,N_21653);
and U25310 (N_25310,N_22632,N_22114);
nor U25311 (N_25311,N_22528,N_23893);
or U25312 (N_25312,N_21323,N_23376);
nand U25313 (N_25313,N_22649,N_21616);
or U25314 (N_25314,N_23001,N_22286);
and U25315 (N_25315,N_23225,N_22021);
xnor U25316 (N_25316,N_21865,N_21942);
or U25317 (N_25317,N_22401,N_22914);
nand U25318 (N_25318,N_21798,N_23234);
nor U25319 (N_25319,N_21713,N_21947);
and U25320 (N_25320,N_23920,N_23993);
nor U25321 (N_25321,N_22491,N_22598);
and U25322 (N_25322,N_21472,N_22470);
nand U25323 (N_25323,N_21585,N_21945);
and U25324 (N_25324,N_23014,N_21692);
or U25325 (N_25325,N_22718,N_23720);
nor U25326 (N_25326,N_23933,N_23370);
nand U25327 (N_25327,N_23856,N_23198);
or U25328 (N_25328,N_22673,N_22196);
xor U25329 (N_25329,N_21791,N_23701);
and U25330 (N_25330,N_22634,N_22540);
nor U25331 (N_25331,N_23543,N_23153);
and U25332 (N_25332,N_23240,N_21319);
nand U25333 (N_25333,N_22300,N_22100);
and U25334 (N_25334,N_22521,N_22266);
and U25335 (N_25335,N_23675,N_22338);
nor U25336 (N_25336,N_21026,N_22733);
nand U25337 (N_25337,N_22677,N_23011);
nand U25338 (N_25338,N_22961,N_22857);
and U25339 (N_25339,N_23116,N_21602);
and U25340 (N_25340,N_22200,N_22430);
or U25341 (N_25341,N_22936,N_21233);
nor U25342 (N_25342,N_23816,N_21669);
nor U25343 (N_25343,N_21973,N_21561);
nand U25344 (N_25344,N_23045,N_23309);
nor U25345 (N_25345,N_21014,N_22000);
or U25346 (N_25346,N_23533,N_22202);
and U25347 (N_25347,N_22703,N_23677);
nand U25348 (N_25348,N_21078,N_23967);
nand U25349 (N_25349,N_22647,N_22159);
nand U25350 (N_25350,N_23193,N_22729);
nand U25351 (N_25351,N_23886,N_22827);
and U25352 (N_25352,N_22845,N_22616);
or U25353 (N_25353,N_21160,N_21760);
or U25354 (N_25354,N_23041,N_22911);
or U25355 (N_25355,N_22547,N_22073);
xnor U25356 (N_25356,N_22989,N_23424);
xnor U25357 (N_25357,N_21721,N_21359);
nor U25358 (N_25358,N_21882,N_22074);
nand U25359 (N_25359,N_23661,N_22652);
xor U25360 (N_25360,N_22311,N_22617);
nand U25361 (N_25361,N_23634,N_23789);
or U25362 (N_25362,N_21102,N_22011);
and U25363 (N_25363,N_23999,N_21660);
nor U25364 (N_25364,N_23667,N_23220);
and U25365 (N_25365,N_21826,N_23053);
and U25366 (N_25366,N_23196,N_22026);
or U25367 (N_25367,N_21649,N_21203);
and U25368 (N_25368,N_22294,N_23747);
xor U25369 (N_25369,N_23735,N_21609);
nand U25370 (N_25370,N_21301,N_21679);
and U25371 (N_25371,N_21125,N_21979);
or U25372 (N_25372,N_21433,N_22597);
nand U25373 (N_25373,N_21241,N_21100);
nor U25374 (N_25374,N_22239,N_21622);
nand U25375 (N_25375,N_21407,N_21275);
and U25376 (N_25376,N_23036,N_23553);
nand U25377 (N_25377,N_21645,N_21734);
nor U25378 (N_25378,N_22087,N_22173);
or U25379 (N_25379,N_23832,N_21068);
and U25380 (N_25380,N_23346,N_23059);
nor U25381 (N_25381,N_21625,N_23034);
xor U25382 (N_25382,N_21191,N_21356);
or U25383 (N_25383,N_21519,N_22863);
nand U25384 (N_25384,N_23536,N_22713);
or U25385 (N_25385,N_23708,N_23650);
and U25386 (N_25386,N_22177,N_22221);
xor U25387 (N_25387,N_22411,N_21898);
nor U25388 (N_25388,N_22494,N_23806);
and U25389 (N_25389,N_23884,N_21293);
nor U25390 (N_25390,N_21429,N_22685);
nor U25391 (N_25391,N_22273,N_22429);
xnor U25392 (N_25392,N_22146,N_22942);
nor U25393 (N_25393,N_23375,N_23408);
and U25394 (N_25394,N_22513,N_21925);
nand U25395 (N_25395,N_21815,N_23217);
or U25396 (N_25396,N_22362,N_23401);
nand U25397 (N_25397,N_23935,N_23743);
nor U25398 (N_25398,N_21127,N_21901);
nor U25399 (N_25399,N_22759,N_21302);
nor U25400 (N_25400,N_23719,N_21446);
xnor U25401 (N_25401,N_21485,N_23849);
or U25402 (N_25402,N_23486,N_21455);
nor U25403 (N_25403,N_22822,N_22784);
and U25404 (N_25404,N_22887,N_21325);
nand U25405 (N_25405,N_23007,N_21349);
nand U25406 (N_25406,N_21452,N_21698);
nor U25407 (N_25407,N_21546,N_23420);
nor U25408 (N_25408,N_23707,N_22006);
and U25409 (N_25409,N_22823,N_23900);
and U25410 (N_25410,N_23722,N_23435);
nor U25411 (N_25411,N_23951,N_22174);
or U25412 (N_25412,N_22309,N_22612);
xor U25413 (N_25413,N_23493,N_23413);
and U25414 (N_25414,N_23632,N_23409);
nand U25415 (N_25415,N_21840,N_23544);
xor U25416 (N_25416,N_21015,N_22878);
nand U25417 (N_25417,N_23214,N_23758);
and U25418 (N_25418,N_23644,N_21465);
nand U25419 (N_25419,N_22701,N_23206);
or U25420 (N_25420,N_21571,N_23657);
and U25421 (N_25421,N_22046,N_23950);
nand U25422 (N_25422,N_22076,N_23855);
or U25423 (N_25423,N_21021,N_23765);
nor U25424 (N_25424,N_23253,N_22039);
nand U25425 (N_25425,N_22892,N_21357);
nand U25426 (N_25426,N_21797,N_22747);
and U25427 (N_25427,N_21887,N_21915);
nand U25428 (N_25428,N_21904,N_23527);
nand U25429 (N_25429,N_22143,N_21352);
nor U25430 (N_25430,N_21483,N_21039);
and U25431 (N_25431,N_23015,N_22426);
nor U25432 (N_25432,N_23731,N_21141);
nand U25433 (N_25433,N_23813,N_23022);
nor U25434 (N_25434,N_23395,N_21620);
nor U25435 (N_25435,N_22872,N_22420);
and U25436 (N_25436,N_22682,N_23292);
and U25437 (N_25437,N_21432,N_23709);
and U25438 (N_25438,N_21347,N_23425);
or U25439 (N_25439,N_22181,N_23237);
nand U25440 (N_25440,N_21318,N_22714);
xnor U25441 (N_25441,N_21154,N_23786);
nand U25442 (N_25442,N_21208,N_22244);
nand U25443 (N_25443,N_21565,N_23546);
nor U25444 (N_25444,N_21050,N_23187);
or U25445 (N_25445,N_23183,N_22515);
nand U25446 (N_25446,N_23705,N_23228);
or U25447 (N_25447,N_22861,N_22444);
or U25448 (N_25448,N_23133,N_23995);
and U25449 (N_25449,N_21867,N_22077);
nor U25450 (N_25450,N_21076,N_22225);
nand U25451 (N_25451,N_22436,N_22359);
nor U25452 (N_25452,N_23267,N_23646);
nor U25453 (N_25453,N_23624,N_23578);
or U25454 (N_25454,N_22764,N_21778);
nor U25455 (N_25455,N_21951,N_22004);
and U25456 (N_25456,N_22651,N_22201);
nor U25457 (N_25457,N_22503,N_21907);
nand U25458 (N_25458,N_23023,N_21605);
and U25459 (N_25459,N_21090,N_23500);
and U25460 (N_25460,N_23568,N_21181);
nand U25461 (N_25461,N_21612,N_23433);
nor U25462 (N_25462,N_21070,N_21399);
nand U25463 (N_25463,N_23324,N_23287);
and U25464 (N_25464,N_21509,N_21518);
and U25465 (N_25465,N_21987,N_22033);
nor U25466 (N_25466,N_22236,N_22661);
nor U25467 (N_25467,N_21346,N_22910);
xor U25468 (N_25468,N_22098,N_21818);
nor U25469 (N_25469,N_21990,N_21274);
and U25470 (N_25470,N_22460,N_21351);
or U25471 (N_25471,N_23464,N_22576);
nand U25472 (N_25472,N_23274,N_22484);
nand U25473 (N_25473,N_23181,N_22587);
nand U25474 (N_25474,N_21576,N_22581);
or U25475 (N_25475,N_21317,N_23864);
or U25476 (N_25476,N_23241,N_22847);
or U25477 (N_25477,N_21606,N_22553);
nand U25478 (N_25478,N_23359,N_22403);
nor U25479 (N_25479,N_21424,N_21122);
or U25480 (N_25480,N_21705,N_22040);
or U25481 (N_25481,N_23975,N_21651);
and U25482 (N_25482,N_23681,N_22488);
or U25483 (N_25483,N_22696,N_22381);
nor U25484 (N_25484,N_23147,N_21134);
xnor U25485 (N_25485,N_23608,N_22199);
and U25486 (N_25486,N_21872,N_23672);
or U25487 (N_25487,N_23279,N_23257);
nor U25488 (N_25488,N_22996,N_21856);
or U25489 (N_25489,N_23467,N_21153);
nor U25490 (N_25490,N_23114,N_23515);
and U25491 (N_25491,N_22248,N_23512);
or U25492 (N_25492,N_23557,N_22334);
nand U25493 (N_25493,N_21971,N_21142);
xor U25494 (N_25494,N_22808,N_22693);
nor U25495 (N_25495,N_22285,N_22112);
nand U25496 (N_25496,N_23882,N_21053);
nand U25497 (N_25497,N_23445,N_23902);
or U25498 (N_25498,N_22880,N_21626);
nor U25499 (N_25499,N_23953,N_22487);
or U25500 (N_25500,N_21876,N_22571);
nand U25501 (N_25501,N_22464,N_22437);
and U25502 (N_25502,N_23481,N_21502);
nor U25503 (N_25503,N_22388,N_22219);
nor U25504 (N_25504,N_21393,N_21932);
or U25505 (N_25505,N_21819,N_22497);
nor U25506 (N_25506,N_21796,N_22886);
xor U25507 (N_25507,N_23104,N_21331);
or U25508 (N_25508,N_23365,N_22285);
or U25509 (N_25509,N_22945,N_23400);
xor U25510 (N_25510,N_23522,N_23617);
nand U25511 (N_25511,N_22732,N_23718);
nor U25512 (N_25512,N_23639,N_22377);
nor U25513 (N_25513,N_21127,N_21532);
and U25514 (N_25514,N_21819,N_21478);
nand U25515 (N_25515,N_22868,N_21664);
and U25516 (N_25516,N_21706,N_21064);
or U25517 (N_25517,N_23501,N_21625);
or U25518 (N_25518,N_22054,N_22608);
nor U25519 (N_25519,N_21368,N_22088);
nor U25520 (N_25520,N_22565,N_21170);
or U25521 (N_25521,N_21042,N_22103);
nor U25522 (N_25522,N_23452,N_23796);
nor U25523 (N_25523,N_22189,N_22780);
or U25524 (N_25524,N_22420,N_22422);
nand U25525 (N_25525,N_21211,N_23031);
or U25526 (N_25526,N_21851,N_22446);
or U25527 (N_25527,N_21417,N_21323);
or U25528 (N_25528,N_21343,N_22627);
or U25529 (N_25529,N_23931,N_21659);
nand U25530 (N_25530,N_22059,N_23126);
nor U25531 (N_25531,N_21603,N_21448);
xor U25532 (N_25532,N_22351,N_23490);
nor U25533 (N_25533,N_21699,N_21359);
or U25534 (N_25534,N_23719,N_23685);
nand U25535 (N_25535,N_23580,N_22080);
and U25536 (N_25536,N_22499,N_21609);
xnor U25537 (N_25537,N_21265,N_22720);
nand U25538 (N_25538,N_22693,N_23900);
and U25539 (N_25539,N_22558,N_23613);
or U25540 (N_25540,N_21162,N_22603);
xnor U25541 (N_25541,N_22969,N_23819);
or U25542 (N_25542,N_21629,N_21170);
and U25543 (N_25543,N_22421,N_22775);
xor U25544 (N_25544,N_22089,N_22512);
and U25545 (N_25545,N_21300,N_22963);
nand U25546 (N_25546,N_21294,N_22832);
and U25547 (N_25547,N_23339,N_22754);
or U25548 (N_25548,N_21068,N_22637);
nor U25549 (N_25549,N_23697,N_23198);
and U25550 (N_25550,N_23635,N_22142);
and U25551 (N_25551,N_21196,N_23812);
and U25552 (N_25552,N_21860,N_22606);
nand U25553 (N_25553,N_22189,N_23102);
xor U25554 (N_25554,N_23184,N_22486);
or U25555 (N_25555,N_23763,N_23949);
and U25556 (N_25556,N_23174,N_23270);
nand U25557 (N_25557,N_22212,N_21834);
nand U25558 (N_25558,N_23872,N_22299);
nor U25559 (N_25559,N_22972,N_23441);
nand U25560 (N_25560,N_23079,N_22694);
xor U25561 (N_25561,N_21694,N_21980);
or U25562 (N_25562,N_23226,N_21596);
nand U25563 (N_25563,N_23242,N_21724);
nand U25564 (N_25564,N_21425,N_23591);
nor U25565 (N_25565,N_23698,N_21648);
or U25566 (N_25566,N_23404,N_23622);
nand U25567 (N_25567,N_23726,N_22561);
or U25568 (N_25568,N_21495,N_21809);
or U25569 (N_25569,N_23389,N_22796);
and U25570 (N_25570,N_23354,N_22480);
nand U25571 (N_25571,N_23251,N_23242);
nor U25572 (N_25572,N_23280,N_21997);
and U25573 (N_25573,N_21682,N_23269);
nand U25574 (N_25574,N_23295,N_23195);
nand U25575 (N_25575,N_21210,N_21885);
nor U25576 (N_25576,N_23009,N_23144);
or U25577 (N_25577,N_23853,N_21502);
nor U25578 (N_25578,N_23471,N_21730);
nand U25579 (N_25579,N_22786,N_22747);
or U25580 (N_25580,N_23646,N_23201);
and U25581 (N_25581,N_22114,N_21203);
and U25582 (N_25582,N_23368,N_22596);
and U25583 (N_25583,N_22648,N_22088);
nor U25584 (N_25584,N_21213,N_23034);
and U25585 (N_25585,N_21600,N_22803);
or U25586 (N_25586,N_21772,N_22009);
nor U25587 (N_25587,N_21362,N_23210);
and U25588 (N_25588,N_21105,N_21608);
xor U25589 (N_25589,N_22475,N_21628);
nand U25590 (N_25590,N_22500,N_23890);
and U25591 (N_25591,N_22988,N_22094);
and U25592 (N_25592,N_21997,N_23647);
or U25593 (N_25593,N_23230,N_22757);
or U25594 (N_25594,N_22449,N_23839);
nand U25595 (N_25595,N_22851,N_23274);
or U25596 (N_25596,N_21915,N_21033);
and U25597 (N_25597,N_21905,N_21668);
nand U25598 (N_25598,N_23143,N_23931);
nor U25599 (N_25599,N_23377,N_22796);
xnor U25600 (N_25600,N_23665,N_23618);
nor U25601 (N_25601,N_22373,N_21483);
xnor U25602 (N_25602,N_23034,N_22900);
nor U25603 (N_25603,N_22416,N_21787);
or U25604 (N_25604,N_23387,N_23072);
nand U25605 (N_25605,N_23943,N_23613);
and U25606 (N_25606,N_21020,N_22240);
nand U25607 (N_25607,N_22122,N_23906);
or U25608 (N_25608,N_21641,N_22349);
or U25609 (N_25609,N_21289,N_21780);
nor U25610 (N_25610,N_23374,N_23556);
nand U25611 (N_25611,N_21218,N_22372);
nand U25612 (N_25612,N_22298,N_22565);
or U25613 (N_25613,N_21644,N_23770);
or U25614 (N_25614,N_21133,N_21324);
nor U25615 (N_25615,N_21331,N_22497);
or U25616 (N_25616,N_23717,N_22774);
and U25617 (N_25617,N_23008,N_23481);
and U25618 (N_25618,N_23104,N_21105);
nand U25619 (N_25619,N_22307,N_21619);
and U25620 (N_25620,N_23729,N_22898);
nand U25621 (N_25621,N_21073,N_23455);
and U25622 (N_25622,N_21213,N_22383);
nor U25623 (N_25623,N_23752,N_21332);
or U25624 (N_25624,N_21760,N_23772);
nor U25625 (N_25625,N_23899,N_21441);
xor U25626 (N_25626,N_21803,N_22222);
xnor U25627 (N_25627,N_22410,N_22552);
or U25628 (N_25628,N_22625,N_21534);
nand U25629 (N_25629,N_21062,N_21304);
nor U25630 (N_25630,N_22035,N_22582);
or U25631 (N_25631,N_22317,N_22516);
nand U25632 (N_25632,N_21499,N_23717);
and U25633 (N_25633,N_21258,N_22781);
or U25634 (N_25634,N_21845,N_21370);
nand U25635 (N_25635,N_21154,N_22007);
nor U25636 (N_25636,N_23364,N_22347);
nor U25637 (N_25637,N_22247,N_21371);
nand U25638 (N_25638,N_23697,N_21467);
or U25639 (N_25639,N_22855,N_21337);
or U25640 (N_25640,N_23555,N_23998);
nand U25641 (N_25641,N_23939,N_23749);
nor U25642 (N_25642,N_22825,N_22705);
or U25643 (N_25643,N_23945,N_21041);
nand U25644 (N_25644,N_22462,N_21088);
and U25645 (N_25645,N_22340,N_22028);
or U25646 (N_25646,N_22986,N_22252);
and U25647 (N_25647,N_23760,N_23317);
nand U25648 (N_25648,N_21751,N_22332);
nor U25649 (N_25649,N_21821,N_22757);
nand U25650 (N_25650,N_21945,N_22204);
nand U25651 (N_25651,N_21148,N_21785);
xor U25652 (N_25652,N_22247,N_21397);
nor U25653 (N_25653,N_22259,N_22861);
nor U25654 (N_25654,N_21259,N_23591);
nor U25655 (N_25655,N_23613,N_21330);
or U25656 (N_25656,N_23750,N_21543);
or U25657 (N_25657,N_22245,N_23107);
and U25658 (N_25658,N_22528,N_22601);
nand U25659 (N_25659,N_21005,N_21053);
and U25660 (N_25660,N_22379,N_23303);
nand U25661 (N_25661,N_21237,N_21521);
nor U25662 (N_25662,N_23296,N_22033);
nor U25663 (N_25663,N_21161,N_21615);
nand U25664 (N_25664,N_22857,N_23214);
and U25665 (N_25665,N_21131,N_21277);
nor U25666 (N_25666,N_21553,N_23316);
xor U25667 (N_25667,N_23328,N_21470);
and U25668 (N_25668,N_22078,N_22634);
nand U25669 (N_25669,N_22645,N_23253);
xor U25670 (N_25670,N_23370,N_21461);
nor U25671 (N_25671,N_23000,N_21823);
nand U25672 (N_25672,N_22610,N_22080);
and U25673 (N_25673,N_22291,N_21215);
nand U25674 (N_25674,N_21876,N_23554);
or U25675 (N_25675,N_23018,N_23272);
or U25676 (N_25676,N_21723,N_23436);
nand U25677 (N_25677,N_21904,N_21148);
nor U25678 (N_25678,N_23345,N_23789);
and U25679 (N_25679,N_22656,N_23215);
nor U25680 (N_25680,N_23683,N_22836);
nand U25681 (N_25681,N_23796,N_21880);
nor U25682 (N_25682,N_23204,N_21927);
nand U25683 (N_25683,N_23603,N_22337);
or U25684 (N_25684,N_23324,N_22401);
and U25685 (N_25685,N_21426,N_22450);
and U25686 (N_25686,N_21204,N_22629);
nand U25687 (N_25687,N_21603,N_21322);
and U25688 (N_25688,N_23054,N_22443);
xnor U25689 (N_25689,N_23407,N_23694);
nor U25690 (N_25690,N_21758,N_23360);
and U25691 (N_25691,N_22746,N_23568);
and U25692 (N_25692,N_21508,N_21167);
nor U25693 (N_25693,N_23844,N_22257);
or U25694 (N_25694,N_22455,N_21154);
nand U25695 (N_25695,N_22538,N_23597);
xnor U25696 (N_25696,N_22717,N_22146);
xor U25697 (N_25697,N_23957,N_21421);
or U25698 (N_25698,N_23247,N_23218);
nand U25699 (N_25699,N_21413,N_21168);
or U25700 (N_25700,N_22903,N_23533);
or U25701 (N_25701,N_21683,N_21828);
and U25702 (N_25702,N_21602,N_23904);
or U25703 (N_25703,N_22261,N_22773);
nor U25704 (N_25704,N_23673,N_23277);
xnor U25705 (N_25705,N_22331,N_23876);
nor U25706 (N_25706,N_21701,N_21669);
nor U25707 (N_25707,N_21409,N_22214);
nand U25708 (N_25708,N_23751,N_22955);
and U25709 (N_25709,N_23275,N_22871);
xnor U25710 (N_25710,N_22358,N_21804);
and U25711 (N_25711,N_23463,N_21940);
nor U25712 (N_25712,N_22727,N_21635);
nor U25713 (N_25713,N_22104,N_21142);
and U25714 (N_25714,N_21876,N_22423);
or U25715 (N_25715,N_22527,N_21396);
xnor U25716 (N_25716,N_23669,N_23049);
nor U25717 (N_25717,N_23000,N_22039);
nand U25718 (N_25718,N_22737,N_22929);
nor U25719 (N_25719,N_22950,N_21561);
nor U25720 (N_25720,N_21639,N_23733);
xnor U25721 (N_25721,N_22977,N_21596);
and U25722 (N_25722,N_21175,N_23778);
or U25723 (N_25723,N_22079,N_22986);
or U25724 (N_25724,N_23776,N_23571);
xor U25725 (N_25725,N_23677,N_22862);
xnor U25726 (N_25726,N_23094,N_23502);
and U25727 (N_25727,N_23013,N_22031);
nand U25728 (N_25728,N_22888,N_23506);
nand U25729 (N_25729,N_23499,N_21755);
or U25730 (N_25730,N_23278,N_23465);
nand U25731 (N_25731,N_21177,N_21487);
and U25732 (N_25732,N_23820,N_22693);
and U25733 (N_25733,N_23986,N_22914);
nand U25734 (N_25734,N_22660,N_22888);
or U25735 (N_25735,N_21581,N_21481);
or U25736 (N_25736,N_23821,N_22097);
or U25737 (N_25737,N_21234,N_21757);
nor U25738 (N_25738,N_21122,N_23910);
xnor U25739 (N_25739,N_21405,N_23266);
or U25740 (N_25740,N_23518,N_23921);
and U25741 (N_25741,N_23110,N_22583);
or U25742 (N_25742,N_22737,N_23168);
nor U25743 (N_25743,N_22800,N_23676);
nor U25744 (N_25744,N_22945,N_22793);
nand U25745 (N_25745,N_22944,N_21005);
nor U25746 (N_25746,N_21773,N_22502);
or U25747 (N_25747,N_23569,N_23529);
nand U25748 (N_25748,N_22507,N_21551);
nor U25749 (N_25749,N_23886,N_22464);
nand U25750 (N_25750,N_22115,N_22909);
and U25751 (N_25751,N_23097,N_23887);
nor U25752 (N_25752,N_23283,N_22744);
nand U25753 (N_25753,N_22419,N_22161);
nand U25754 (N_25754,N_23381,N_23126);
or U25755 (N_25755,N_23851,N_21675);
nand U25756 (N_25756,N_23679,N_21060);
or U25757 (N_25757,N_23507,N_22712);
nand U25758 (N_25758,N_23842,N_23308);
and U25759 (N_25759,N_23366,N_23192);
or U25760 (N_25760,N_22948,N_21939);
and U25761 (N_25761,N_21532,N_23576);
and U25762 (N_25762,N_21338,N_21476);
nor U25763 (N_25763,N_23607,N_21245);
xnor U25764 (N_25764,N_23525,N_21319);
nand U25765 (N_25765,N_21503,N_22330);
or U25766 (N_25766,N_21696,N_23186);
and U25767 (N_25767,N_21615,N_21155);
nor U25768 (N_25768,N_23577,N_21794);
or U25769 (N_25769,N_23088,N_22819);
and U25770 (N_25770,N_21843,N_22219);
nor U25771 (N_25771,N_22477,N_23402);
nand U25772 (N_25772,N_23677,N_21355);
nand U25773 (N_25773,N_23767,N_21586);
xnor U25774 (N_25774,N_22280,N_22081);
and U25775 (N_25775,N_21780,N_21513);
nand U25776 (N_25776,N_22448,N_21156);
nor U25777 (N_25777,N_23473,N_23952);
nand U25778 (N_25778,N_22148,N_21031);
nand U25779 (N_25779,N_23785,N_23083);
nand U25780 (N_25780,N_23212,N_23928);
nand U25781 (N_25781,N_22277,N_23107);
or U25782 (N_25782,N_21842,N_22970);
nand U25783 (N_25783,N_22313,N_22315);
nand U25784 (N_25784,N_23385,N_22775);
nor U25785 (N_25785,N_21336,N_22126);
or U25786 (N_25786,N_21687,N_21994);
and U25787 (N_25787,N_21298,N_22720);
and U25788 (N_25788,N_21718,N_23144);
nor U25789 (N_25789,N_21334,N_23484);
or U25790 (N_25790,N_21649,N_21068);
xnor U25791 (N_25791,N_21172,N_23656);
nor U25792 (N_25792,N_23836,N_23023);
nor U25793 (N_25793,N_22433,N_21639);
nand U25794 (N_25794,N_21081,N_22629);
nor U25795 (N_25795,N_23490,N_21232);
or U25796 (N_25796,N_22889,N_22464);
nand U25797 (N_25797,N_23557,N_23449);
nand U25798 (N_25798,N_22285,N_22338);
nand U25799 (N_25799,N_22816,N_23743);
and U25800 (N_25800,N_22358,N_23764);
xnor U25801 (N_25801,N_22227,N_23221);
nor U25802 (N_25802,N_21001,N_22220);
nor U25803 (N_25803,N_22183,N_23430);
or U25804 (N_25804,N_23215,N_22597);
xnor U25805 (N_25805,N_22877,N_21283);
xnor U25806 (N_25806,N_21398,N_22735);
xnor U25807 (N_25807,N_23606,N_21813);
and U25808 (N_25808,N_21970,N_23759);
and U25809 (N_25809,N_22368,N_22796);
xor U25810 (N_25810,N_22823,N_21839);
and U25811 (N_25811,N_22992,N_21230);
or U25812 (N_25812,N_21434,N_23390);
and U25813 (N_25813,N_21278,N_21463);
or U25814 (N_25814,N_23500,N_22783);
or U25815 (N_25815,N_22411,N_23154);
and U25816 (N_25816,N_22830,N_22047);
nor U25817 (N_25817,N_23762,N_22368);
or U25818 (N_25818,N_21548,N_23920);
nor U25819 (N_25819,N_21711,N_22821);
nand U25820 (N_25820,N_22858,N_23573);
and U25821 (N_25821,N_23680,N_22575);
or U25822 (N_25822,N_21530,N_23425);
and U25823 (N_25823,N_22514,N_21537);
nand U25824 (N_25824,N_23374,N_21639);
and U25825 (N_25825,N_22834,N_22919);
or U25826 (N_25826,N_21261,N_23576);
nor U25827 (N_25827,N_23699,N_23416);
or U25828 (N_25828,N_23987,N_23815);
nand U25829 (N_25829,N_21776,N_21681);
and U25830 (N_25830,N_23650,N_21572);
nor U25831 (N_25831,N_23097,N_21488);
or U25832 (N_25832,N_21404,N_22173);
nand U25833 (N_25833,N_21481,N_21810);
and U25834 (N_25834,N_23045,N_23091);
nor U25835 (N_25835,N_23805,N_23285);
nor U25836 (N_25836,N_22968,N_22802);
xnor U25837 (N_25837,N_22198,N_21052);
nor U25838 (N_25838,N_21869,N_21871);
xnor U25839 (N_25839,N_23033,N_22750);
and U25840 (N_25840,N_23236,N_21273);
nand U25841 (N_25841,N_22657,N_21891);
nand U25842 (N_25842,N_23853,N_22723);
nor U25843 (N_25843,N_21815,N_21985);
and U25844 (N_25844,N_21861,N_21692);
and U25845 (N_25845,N_23949,N_21458);
nand U25846 (N_25846,N_23059,N_22981);
nand U25847 (N_25847,N_21849,N_22653);
nand U25848 (N_25848,N_22986,N_22239);
nand U25849 (N_25849,N_23930,N_22579);
nor U25850 (N_25850,N_23496,N_23534);
nand U25851 (N_25851,N_21656,N_23558);
xnor U25852 (N_25852,N_22428,N_23048);
or U25853 (N_25853,N_23155,N_21992);
or U25854 (N_25854,N_22342,N_22855);
and U25855 (N_25855,N_22733,N_23382);
nand U25856 (N_25856,N_23978,N_22267);
xor U25857 (N_25857,N_23719,N_22880);
and U25858 (N_25858,N_22567,N_23798);
xor U25859 (N_25859,N_23039,N_21072);
nand U25860 (N_25860,N_23109,N_22665);
nand U25861 (N_25861,N_22709,N_22150);
nand U25862 (N_25862,N_23448,N_23923);
and U25863 (N_25863,N_23112,N_22487);
nand U25864 (N_25864,N_22072,N_23280);
nor U25865 (N_25865,N_22790,N_22960);
nor U25866 (N_25866,N_23374,N_22494);
and U25867 (N_25867,N_22020,N_23250);
nor U25868 (N_25868,N_23634,N_23706);
or U25869 (N_25869,N_23034,N_21802);
and U25870 (N_25870,N_23514,N_23453);
nor U25871 (N_25871,N_22765,N_21599);
nor U25872 (N_25872,N_21836,N_23866);
nor U25873 (N_25873,N_23788,N_23171);
nor U25874 (N_25874,N_21553,N_23253);
or U25875 (N_25875,N_23800,N_23033);
xor U25876 (N_25876,N_23658,N_22903);
nor U25877 (N_25877,N_21778,N_23085);
or U25878 (N_25878,N_23970,N_21461);
or U25879 (N_25879,N_22310,N_23516);
nand U25880 (N_25880,N_21356,N_23177);
and U25881 (N_25881,N_23913,N_21953);
or U25882 (N_25882,N_21576,N_22878);
or U25883 (N_25883,N_21937,N_23188);
or U25884 (N_25884,N_21865,N_23738);
or U25885 (N_25885,N_22410,N_22350);
nor U25886 (N_25886,N_21436,N_23438);
or U25887 (N_25887,N_22496,N_23352);
or U25888 (N_25888,N_22605,N_23016);
and U25889 (N_25889,N_22028,N_22899);
and U25890 (N_25890,N_23759,N_22153);
nand U25891 (N_25891,N_23952,N_22647);
or U25892 (N_25892,N_21692,N_23204);
nor U25893 (N_25893,N_23621,N_23065);
or U25894 (N_25894,N_22741,N_21560);
nor U25895 (N_25895,N_21789,N_22080);
nand U25896 (N_25896,N_22381,N_23160);
nand U25897 (N_25897,N_21626,N_23672);
nand U25898 (N_25898,N_23736,N_21791);
and U25899 (N_25899,N_22910,N_21176);
and U25900 (N_25900,N_21798,N_21108);
and U25901 (N_25901,N_22309,N_23621);
or U25902 (N_25902,N_22727,N_23314);
nand U25903 (N_25903,N_23163,N_23909);
xor U25904 (N_25904,N_21828,N_23686);
nand U25905 (N_25905,N_21356,N_22102);
and U25906 (N_25906,N_23572,N_21214);
nand U25907 (N_25907,N_23456,N_21514);
nor U25908 (N_25908,N_22337,N_22539);
nor U25909 (N_25909,N_22913,N_21122);
nor U25910 (N_25910,N_23140,N_22572);
nand U25911 (N_25911,N_21037,N_21834);
nand U25912 (N_25912,N_21688,N_21053);
xnor U25913 (N_25913,N_21406,N_22414);
nand U25914 (N_25914,N_22365,N_21241);
and U25915 (N_25915,N_22282,N_21251);
nor U25916 (N_25916,N_21391,N_22399);
or U25917 (N_25917,N_22304,N_22867);
xnor U25918 (N_25918,N_21504,N_22974);
nor U25919 (N_25919,N_22472,N_21528);
or U25920 (N_25920,N_21046,N_23592);
nor U25921 (N_25921,N_22475,N_22541);
nor U25922 (N_25922,N_21176,N_21599);
and U25923 (N_25923,N_22124,N_22411);
nand U25924 (N_25924,N_23810,N_22038);
nor U25925 (N_25925,N_21201,N_22307);
nor U25926 (N_25926,N_23011,N_22411);
nor U25927 (N_25927,N_22401,N_22463);
or U25928 (N_25928,N_23384,N_22298);
nor U25929 (N_25929,N_23451,N_23385);
xnor U25930 (N_25930,N_21110,N_23916);
nand U25931 (N_25931,N_21588,N_21401);
or U25932 (N_25932,N_21198,N_21695);
nor U25933 (N_25933,N_23111,N_22973);
and U25934 (N_25934,N_23884,N_22209);
nand U25935 (N_25935,N_21474,N_23553);
nor U25936 (N_25936,N_23943,N_21556);
or U25937 (N_25937,N_23665,N_21967);
nand U25938 (N_25938,N_21865,N_21922);
nand U25939 (N_25939,N_21767,N_22999);
xor U25940 (N_25940,N_21657,N_22126);
and U25941 (N_25941,N_23060,N_22305);
xor U25942 (N_25942,N_21876,N_21979);
nor U25943 (N_25943,N_23276,N_22856);
nand U25944 (N_25944,N_23794,N_22584);
nor U25945 (N_25945,N_21811,N_21196);
or U25946 (N_25946,N_21456,N_21911);
and U25947 (N_25947,N_21144,N_23694);
nor U25948 (N_25948,N_21217,N_23170);
nor U25949 (N_25949,N_22945,N_21291);
and U25950 (N_25950,N_23970,N_22117);
and U25951 (N_25951,N_22002,N_23075);
or U25952 (N_25952,N_21305,N_23431);
or U25953 (N_25953,N_22999,N_22231);
or U25954 (N_25954,N_21084,N_21108);
or U25955 (N_25955,N_22893,N_21293);
and U25956 (N_25956,N_22186,N_22936);
nand U25957 (N_25957,N_23541,N_23351);
or U25958 (N_25958,N_22937,N_23555);
xor U25959 (N_25959,N_21978,N_21926);
nor U25960 (N_25960,N_23978,N_23571);
nor U25961 (N_25961,N_21451,N_22358);
nor U25962 (N_25962,N_22764,N_21618);
nand U25963 (N_25963,N_21714,N_22005);
or U25964 (N_25964,N_22921,N_21936);
nand U25965 (N_25965,N_21863,N_22951);
and U25966 (N_25966,N_21350,N_23038);
nand U25967 (N_25967,N_22598,N_23471);
nand U25968 (N_25968,N_22203,N_22047);
or U25969 (N_25969,N_22631,N_21328);
nor U25970 (N_25970,N_23053,N_23971);
nor U25971 (N_25971,N_23530,N_22129);
nand U25972 (N_25972,N_22381,N_22981);
nand U25973 (N_25973,N_23539,N_23337);
and U25974 (N_25974,N_23821,N_22709);
nor U25975 (N_25975,N_23973,N_21586);
and U25976 (N_25976,N_22868,N_23892);
nand U25977 (N_25977,N_22081,N_23304);
or U25978 (N_25978,N_21303,N_22928);
nor U25979 (N_25979,N_23480,N_22460);
nor U25980 (N_25980,N_21953,N_22266);
xnor U25981 (N_25981,N_21646,N_22770);
xor U25982 (N_25982,N_23528,N_21308);
or U25983 (N_25983,N_23502,N_23950);
nand U25984 (N_25984,N_21691,N_21786);
or U25985 (N_25985,N_22984,N_22961);
or U25986 (N_25986,N_21656,N_21893);
and U25987 (N_25987,N_23309,N_21681);
xnor U25988 (N_25988,N_21705,N_21906);
nand U25989 (N_25989,N_23300,N_22996);
xnor U25990 (N_25990,N_22159,N_23637);
nor U25991 (N_25991,N_21402,N_22755);
and U25992 (N_25992,N_21754,N_22250);
or U25993 (N_25993,N_22641,N_22941);
or U25994 (N_25994,N_22636,N_21918);
or U25995 (N_25995,N_22395,N_22398);
nor U25996 (N_25996,N_23095,N_21402);
and U25997 (N_25997,N_23170,N_22390);
and U25998 (N_25998,N_23051,N_21851);
and U25999 (N_25999,N_21403,N_22865);
nand U26000 (N_26000,N_23892,N_23675);
or U26001 (N_26001,N_22595,N_22176);
nor U26002 (N_26002,N_21184,N_23107);
and U26003 (N_26003,N_21507,N_21310);
and U26004 (N_26004,N_23216,N_22872);
xnor U26005 (N_26005,N_21594,N_23867);
or U26006 (N_26006,N_22400,N_23711);
nor U26007 (N_26007,N_23508,N_21749);
and U26008 (N_26008,N_21503,N_23128);
xor U26009 (N_26009,N_23327,N_21043);
nand U26010 (N_26010,N_23540,N_23592);
nand U26011 (N_26011,N_22341,N_21796);
or U26012 (N_26012,N_21791,N_23857);
nand U26013 (N_26013,N_22808,N_23279);
nand U26014 (N_26014,N_21785,N_22818);
xnor U26015 (N_26015,N_21846,N_21732);
and U26016 (N_26016,N_21473,N_23107);
nor U26017 (N_26017,N_23916,N_22020);
and U26018 (N_26018,N_22842,N_23193);
and U26019 (N_26019,N_22194,N_22148);
or U26020 (N_26020,N_21149,N_22297);
nor U26021 (N_26021,N_22465,N_22421);
nand U26022 (N_26022,N_21921,N_23452);
and U26023 (N_26023,N_21211,N_21777);
nor U26024 (N_26024,N_21540,N_21050);
or U26025 (N_26025,N_23252,N_23329);
nor U26026 (N_26026,N_23273,N_21378);
or U26027 (N_26027,N_23885,N_23490);
and U26028 (N_26028,N_21615,N_21042);
or U26029 (N_26029,N_21242,N_23631);
nor U26030 (N_26030,N_21674,N_23520);
or U26031 (N_26031,N_21027,N_22399);
nor U26032 (N_26032,N_22232,N_23058);
and U26033 (N_26033,N_23975,N_23993);
nor U26034 (N_26034,N_21729,N_23606);
nand U26035 (N_26035,N_21350,N_23216);
nand U26036 (N_26036,N_23230,N_22963);
nor U26037 (N_26037,N_23613,N_21133);
and U26038 (N_26038,N_21701,N_23497);
nand U26039 (N_26039,N_23848,N_21420);
nor U26040 (N_26040,N_21051,N_22141);
or U26041 (N_26041,N_21388,N_22476);
nand U26042 (N_26042,N_21183,N_21320);
nor U26043 (N_26043,N_23519,N_23120);
and U26044 (N_26044,N_21064,N_23325);
nor U26045 (N_26045,N_22598,N_22917);
nor U26046 (N_26046,N_21055,N_23741);
and U26047 (N_26047,N_21922,N_21853);
and U26048 (N_26048,N_22412,N_21174);
or U26049 (N_26049,N_22254,N_22062);
or U26050 (N_26050,N_23260,N_21726);
and U26051 (N_26051,N_23650,N_21593);
nor U26052 (N_26052,N_23957,N_23091);
nor U26053 (N_26053,N_23084,N_22232);
nor U26054 (N_26054,N_23651,N_22511);
nand U26055 (N_26055,N_22111,N_22360);
nor U26056 (N_26056,N_22023,N_22552);
or U26057 (N_26057,N_22050,N_23855);
xor U26058 (N_26058,N_21554,N_22295);
nor U26059 (N_26059,N_21869,N_22918);
nand U26060 (N_26060,N_22696,N_22502);
nor U26061 (N_26061,N_23865,N_21869);
xnor U26062 (N_26062,N_22262,N_23677);
xor U26063 (N_26063,N_23786,N_21928);
and U26064 (N_26064,N_22509,N_21019);
nor U26065 (N_26065,N_23853,N_22114);
and U26066 (N_26066,N_23260,N_23358);
and U26067 (N_26067,N_21569,N_22790);
nand U26068 (N_26068,N_22474,N_23585);
nand U26069 (N_26069,N_22656,N_23843);
xnor U26070 (N_26070,N_22741,N_22661);
and U26071 (N_26071,N_22644,N_21418);
xor U26072 (N_26072,N_23890,N_23623);
xnor U26073 (N_26073,N_21223,N_21726);
or U26074 (N_26074,N_21871,N_23285);
nand U26075 (N_26075,N_22084,N_22763);
and U26076 (N_26076,N_21089,N_21513);
and U26077 (N_26077,N_23317,N_22098);
or U26078 (N_26078,N_22325,N_22399);
nand U26079 (N_26079,N_23430,N_22474);
nand U26080 (N_26080,N_21150,N_22328);
nand U26081 (N_26081,N_21636,N_23930);
xor U26082 (N_26082,N_21825,N_22123);
nand U26083 (N_26083,N_21076,N_21260);
nand U26084 (N_26084,N_22140,N_23880);
nand U26085 (N_26085,N_22344,N_21172);
and U26086 (N_26086,N_21732,N_23812);
nor U26087 (N_26087,N_23277,N_21145);
nor U26088 (N_26088,N_21736,N_22387);
xor U26089 (N_26089,N_21100,N_22265);
or U26090 (N_26090,N_22200,N_23181);
and U26091 (N_26091,N_22603,N_22345);
nand U26092 (N_26092,N_22204,N_23064);
or U26093 (N_26093,N_21914,N_22907);
nand U26094 (N_26094,N_22599,N_21474);
or U26095 (N_26095,N_23586,N_23724);
nor U26096 (N_26096,N_21166,N_21953);
or U26097 (N_26097,N_22286,N_22517);
nand U26098 (N_26098,N_21720,N_21620);
or U26099 (N_26099,N_21324,N_22030);
or U26100 (N_26100,N_23671,N_22553);
nor U26101 (N_26101,N_22768,N_23883);
and U26102 (N_26102,N_21894,N_21921);
xnor U26103 (N_26103,N_22728,N_22100);
nor U26104 (N_26104,N_22790,N_23942);
nand U26105 (N_26105,N_21962,N_23118);
xor U26106 (N_26106,N_22293,N_23488);
nand U26107 (N_26107,N_22641,N_21880);
nand U26108 (N_26108,N_21424,N_21749);
and U26109 (N_26109,N_23194,N_22567);
or U26110 (N_26110,N_22199,N_21007);
or U26111 (N_26111,N_21037,N_21237);
nor U26112 (N_26112,N_22948,N_23902);
nor U26113 (N_26113,N_22208,N_21009);
or U26114 (N_26114,N_22843,N_22045);
or U26115 (N_26115,N_22451,N_23658);
xor U26116 (N_26116,N_21456,N_21727);
nand U26117 (N_26117,N_23486,N_21047);
nand U26118 (N_26118,N_23152,N_22018);
nand U26119 (N_26119,N_21427,N_22687);
nor U26120 (N_26120,N_23558,N_21548);
nor U26121 (N_26121,N_22975,N_23425);
and U26122 (N_26122,N_22235,N_22663);
xor U26123 (N_26123,N_21632,N_23326);
or U26124 (N_26124,N_23663,N_22457);
nor U26125 (N_26125,N_22098,N_21259);
xnor U26126 (N_26126,N_23563,N_21358);
or U26127 (N_26127,N_23593,N_21148);
and U26128 (N_26128,N_23201,N_23941);
or U26129 (N_26129,N_22843,N_23073);
nand U26130 (N_26130,N_22067,N_22417);
nand U26131 (N_26131,N_21400,N_21025);
or U26132 (N_26132,N_23017,N_21219);
xor U26133 (N_26133,N_23714,N_23197);
nand U26134 (N_26134,N_23571,N_21183);
and U26135 (N_26135,N_21922,N_22136);
and U26136 (N_26136,N_21388,N_21396);
and U26137 (N_26137,N_21893,N_23614);
nand U26138 (N_26138,N_21271,N_21894);
nor U26139 (N_26139,N_23976,N_21902);
and U26140 (N_26140,N_21278,N_22896);
nand U26141 (N_26141,N_21264,N_22821);
and U26142 (N_26142,N_23443,N_22928);
nand U26143 (N_26143,N_22095,N_23070);
and U26144 (N_26144,N_22862,N_23168);
xor U26145 (N_26145,N_21622,N_22063);
nor U26146 (N_26146,N_23771,N_23218);
or U26147 (N_26147,N_22423,N_22191);
nand U26148 (N_26148,N_22326,N_22937);
nand U26149 (N_26149,N_23371,N_21222);
xnor U26150 (N_26150,N_22206,N_22842);
and U26151 (N_26151,N_23106,N_23507);
or U26152 (N_26152,N_21561,N_21934);
and U26153 (N_26153,N_22977,N_21595);
nand U26154 (N_26154,N_22297,N_23286);
nand U26155 (N_26155,N_21306,N_22668);
and U26156 (N_26156,N_22035,N_22079);
and U26157 (N_26157,N_21744,N_23667);
nor U26158 (N_26158,N_22887,N_22784);
nand U26159 (N_26159,N_22044,N_22944);
nor U26160 (N_26160,N_22695,N_21076);
or U26161 (N_26161,N_22756,N_22282);
nand U26162 (N_26162,N_23093,N_21915);
nor U26163 (N_26163,N_22071,N_23309);
nand U26164 (N_26164,N_21908,N_23111);
or U26165 (N_26165,N_22051,N_21235);
or U26166 (N_26166,N_23281,N_23235);
nand U26167 (N_26167,N_22556,N_22256);
and U26168 (N_26168,N_22162,N_23640);
and U26169 (N_26169,N_23599,N_22955);
nand U26170 (N_26170,N_21955,N_22876);
or U26171 (N_26171,N_22971,N_21903);
or U26172 (N_26172,N_22015,N_22949);
nand U26173 (N_26173,N_23610,N_22722);
and U26174 (N_26174,N_22692,N_22200);
and U26175 (N_26175,N_23244,N_21516);
nand U26176 (N_26176,N_21098,N_21367);
nor U26177 (N_26177,N_22128,N_23008);
nor U26178 (N_26178,N_22071,N_22905);
or U26179 (N_26179,N_23617,N_21496);
or U26180 (N_26180,N_22924,N_22991);
xnor U26181 (N_26181,N_21007,N_23181);
and U26182 (N_26182,N_23054,N_23976);
nor U26183 (N_26183,N_22664,N_21464);
nor U26184 (N_26184,N_23597,N_22031);
nand U26185 (N_26185,N_22262,N_23175);
nor U26186 (N_26186,N_23998,N_23240);
nor U26187 (N_26187,N_23651,N_22261);
and U26188 (N_26188,N_23968,N_23534);
or U26189 (N_26189,N_21390,N_22081);
or U26190 (N_26190,N_23051,N_21774);
and U26191 (N_26191,N_22053,N_21172);
or U26192 (N_26192,N_23424,N_21109);
nand U26193 (N_26193,N_23269,N_21965);
nor U26194 (N_26194,N_23395,N_23782);
and U26195 (N_26195,N_21112,N_22238);
or U26196 (N_26196,N_23287,N_23216);
nand U26197 (N_26197,N_23348,N_21377);
and U26198 (N_26198,N_22545,N_21456);
nand U26199 (N_26199,N_23439,N_21367);
nor U26200 (N_26200,N_22844,N_22312);
nand U26201 (N_26201,N_21019,N_23758);
or U26202 (N_26202,N_22201,N_21495);
nor U26203 (N_26203,N_23168,N_23842);
and U26204 (N_26204,N_22464,N_22345);
nand U26205 (N_26205,N_21323,N_23176);
nor U26206 (N_26206,N_22831,N_21495);
xor U26207 (N_26207,N_23307,N_22796);
nand U26208 (N_26208,N_21878,N_23930);
and U26209 (N_26209,N_21168,N_21994);
and U26210 (N_26210,N_23873,N_21481);
and U26211 (N_26211,N_23139,N_23205);
xor U26212 (N_26212,N_21784,N_21599);
and U26213 (N_26213,N_22172,N_21838);
nand U26214 (N_26214,N_21208,N_21525);
and U26215 (N_26215,N_21760,N_23464);
and U26216 (N_26216,N_23038,N_22132);
or U26217 (N_26217,N_22488,N_23334);
or U26218 (N_26218,N_23820,N_22044);
or U26219 (N_26219,N_21225,N_21849);
nand U26220 (N_26220,N_21092,N_22593);
nor U26221 (N_26221,N_23822,N_23798);
nand U26222 (N_26222,N_21646,N_23165);
and U26223 (N_26223,N_21523,N_23238);
nor U26224 (N_26224,N_22230,N_22808);
and U26225 (N_26225,N_22276,N_22123);
xnor U26226 (N_26226,N_21498,N_22516);
nor U26227 (N_26227,N_23999,N_23384);
nor U26228 (N_26228,N_23082,N_21851);
nor U26229 (N_26229,N_21465,N_21956);
nand U26230 (N_26230,N_21833,N_21408);
nand U26231 (N_26231,N_22452,N_23522);
xor U26232 (N_26232,N_23122,N_21097);
nor U26233 (N_26233,N_23877,N_23726);
xor U26234 (N_26234,N_21548,N_23116);
nor U26235 (N_26235,N_21593,N_23413);
nor U26236 (N_26236,N_23689,N_22615);
or U26237 (N_26237,N_21583,N_21244);
xnor U26238 (N_26238,N_22283,N_22976);
xnor U26239 (N_26239,N_22359,N_23769);
or U26240 (N_26240,N_23899,N_22381);
nor U26241 (N_26241,N_23480,N_21569);
and U26242 (N_26242,N_22715,N_21228);
nor U26243 (N_26243,N_22881,N_22381);
nand U26244 (N_26244,N_21039,N_21495);
and U26245 (N_26245,N_21779,N_21057);
nor U26246 (N_26246,N_23418,N_23231);
nand U26247 (N_26247,N_22357,N_23582);
or U26248 (N_26248,N_22839,N_22481);
and U26249 (N_26249,N_21808,N_22437);
or U26250 (N_26250,N_22359,N_21567);
nor U26251 (N_26251,N_22736,N_21108);
and U26252 (N_26252,N_22751,N_21014);
nor U26253 (N_26253,N_23466,N_23255);
and U26254 (N_26254,N_21871,N_23886);
nand U26255 (N_26255,N_21041,N_22536);
nand U26256 (N_26256,N_21701,N_23600);
nor U26257 (N_26257,N_22676,N_22218);
xnor U26258 (N_26258,N_21332,N_21621);
or U26259 (N_26259,N_23699,N_22982);
nand U26260 (N_26260,N_23482,N_21657);
and U26261 (N_26261,N_22522,N_23326);
and U26262 (N_26262,N_22551,N_22983);
and U26263 (N_26263,N_22018,N_21203);
nand U26264 (N_26264,N_21726,N_22113);
nor U26265 (N_26265,N_22696,N_21750);
or U26266 (N_26266,N_22397,N_21233);
nor U26267 (N_26267,N_21558,N_22611);
xor U26268 (N_26268,N_21207,N_21339);
nor U26269 (N_26269,N_23985,N_22658);
or U26270 (N_26270,N_23413,N_22037);
or U26271 (N_26271,N_21187,N_23997);
xnor U26272 (N_26272,N_22077,N_22259);
nor U26273 (N_26273,N_21676,N_21997);
or U26274 (N_26274,N_22062,N_22733);
and U26275 (N_26275,N_22155,N_21156);
nand U26276 (N_26276,N_23153,N_23148);
and U26277 (N_26277,N_23873,N_21470);
and U26278 (N_26278,N_23612,N_21285);
nor U26279 (N_26279,N_21022,N_23230);
xor U26280 (N_26280,N_21667,N_22240);
and U26281 (N_26281,N_21959,N_22735);
or U26282 (N_26282,N_23152,N_23293);
nor U26283 (N_26283,N_23465,N_22350);
and U26284 (N_26284,N_22218,N_23018);
and U26285 (N_26285,N_21267,N_21917);
xor U26286 (N_26286,N_21231,N_22298);
nand U26287 (N_26287,N_22412,N_23659);
xnor U26288 (N_26288,N_23652,N_21391);
nor U26289 (N_26289,N_23116,N_22057);
and U26290 (N_26290,N_22493,N_22036);
or U26291 (N_26291,N_21126,N_23894);
nand U26292 (N_26292,N_23976,N_23750);
nand U26293 (N_26293,N_21495,N_21992);
nand U26294 (N_26294,N_22427,N_23227);
or U26295 (N_26295,N_21032,N_23504);
or U26296 (N_26296,N_23080,N_22832);
and U26297 (N_26297,N_21591,N_21381);
nand U26298 (N_26298,N_23750,N_23626);
or U26299 (N_26299,N_23996,N_22898);
and U26300 (N_26300,N_23997,N_23858);
and U26301 (N_26301,N_21416,N_22416);
nand U26302 (N_26302,N_22033,N_21050);
nand U26303 (N_26303,N_23204,N_23561);
or U26304 (N_26304,N_22640,N_22326);
nor U26305 (N_26305,N_21270,N_23605);
or U26306 (N_26306,N_22008,N_21476);
or U26307 (N_26307,N_23318,N_21636);
nand U26308 (N_26308,N_23675,N_21017);
xnor U26309 (N_26309,N_21610,N_22234);
nand U26310 (N_26310,N_21499,N_22481);
nand U26311 (N_26311,N_23980,N_23842);
nor U26312 (N_26312,N_22440,N_23795);
nor U26313 (N_26313,N_23679,N_23696);
and U26314 (N_26314,N_21911,N_22427);
nor U26315 (N_26315,N_23270,N_23451);
nor U26316 (N_26316,N_22094,N_22790);
nor U26317 (N_26317,N_21969,N_22712);
and U26318 (N_26318,N_23860,N_21158);
xor U26319 (N_26319,N_23387,N_22849);
nor U26320 (N_26320,N_22019,N_22148);
nand U26321 (N_26321,N_23505,N_22866);
and U26322 (N_26322,N_23671,N_23605);
and U26323 (N_26323,N_23199,N_21851);
nand U26324 (N_26324,N_23773,N_21276);
nand U26325 (N_26325,N_22680,N_21411);
and U26326 (N_26326,N_21679,N_22897);
nor U26327 (N_26327,N_23630,N_21142);
and U26328 (N_26328,N_23906,N_23776);
nand U26329 (N_26329,N_22426,N_23232);
nand U26330 (N_26330,N_23181,N_21942);
xnor U26331 (N_26331,N_22336,N_23182);
nand U26332 (N_26332,N_23502,N_21838);
or U26333 (N_26333,N_22474,N_23600);
and U26334 (N_26334,N_21558,N_21047);
or U26335 (N_26335,N_23932,N_23848);
xnor U26336 (N_26336,N_22502,N_23370);
and U26337 (N_26337,N_22944,N_22589);
or U26338 (N_26338,N_23901,N_22258);
nand U26339 (N_26339,N_23769,N_22848);
and U26340 (N_26340,N_21647,N_23476);
and U26341 (N_26341,N_23880,N_23933);
nor U26342 (N_26342,N_22684,N_22773);
and U26343 (N_26343,N_21463,N_21521);
nand U26344 (N_26344,N_22863,N_22920);
nand U26345 (N_26345,N_21348,N_21453);
and U26346 (N_26346,N_21658,N_23242);
nand U26347 (N_26347,N_21243,N_23320);
xnor U26348 (N_26348,N_21275,N_21453);
or U26349 (N_26349,N_22282,N_23875);
or U26350 (N_26350,N_21036,N_21292);
nor U26351 (N_26351,N_23756,N_22301);
nand U26352 (N_26352,N_23323,N_22917);
nor U26353 (N_26353,N_22762,N_22644);
or U26354 (N_26354,N_22570,N_21853);
and U26355 (N_26355,N_22650,N_21038);
nor U26356 (N_26356,N_21090,N_22756);
or U26357 (N_26357,N_22669,N_22431);
or U26358 (N_26358,N_23138,N_21285);
and U26359 (N_26359,N_22166,N_21799);
and U26360 (N_26360,N_21310,N_22475);
nor U26361 (N_26361,N_21307,N_23074);
and U26362 (N_26362,N_21393,N_22945);
or U26363 (N_26363,N_21509,N_22771);
or U26364 (N_26364,N_23679,N_23118);
nand U26365 (N_26365,N_21502,N_23262);
and U26366 (N_26366,N_22003,N_22335);
or U26367 (N_26367,N_22898,N_22088);
nor U26368 (N_26368,N_22973,N_23816);
nand U26369 (N_26369,N_23635,N_22348);
and U26370 (N_26370,N_23794,N_21298);
nand U26371 (N_26371,N_23647,N_23991);
nand U26372 (N_26372,N_22951,N_21158);
xnor U26373 (N_26373,N_21439,N_23289);
nand U26374 (N_26374,N_21315,N_22223);
xnor U26375 (N_26375,N_22694,N_23265);
nor U26376 (N_26376,N_22422,N_23220);
nor U26377 (N_26377,N_22298,N_23752);
nor U26378 (N_26378,N_21871,N_23768);
or U26379 (N_26379,N_22848,N_21039);
and U26380 (N_26380,N_23304,N_21299);
and U26381 (N_26381,N_23885,N_21360);
nand U26382 (N_26382,N_23707,N_23027);
xnor U26383 (N_26383,N_23500,N_23127);
or U26384 (N_26384,N_23592,N_23909);
nand U26385 (N_26385,N_21260,N_21244);
or U26386 (N_26386,N_21932,N_22682);
nand U26387 (N_26387,N_23490,N_22233);
and U26388 (N_26388,N_22804,N_22121);
and U26389 (N_26389,N_21494,N_23258);
xnor U26390 (N_26390,N_21034,N_22828);
nand U26391 (N_26391,N_21406,N_23934);
and U26392 (N_26392,N_23197,N_23060);
xnor U26393 (N_26393,N_23231,N_23355);
or U26394 (N_26394,N_21471,N_23623);
xnor U26395 (N_26395,N_21131,N_23433);
and U26396 (N_26396,N_22630,N_22813);
and U26397 (N_26397,N_22152,N_21202);
nor U26398 (N_26398,N_23798,N_21009);
nand U26399 (N_26399,N_21256,N_21852);
nand U26400 (N_26400,N_23530,N_22783);
or U26401 (N_26401,N_23029,N_21648);
or U26402 (N_26402,N_22390,N_23463);
or U26403 (N_26403,N_23177,N_22475);
or U26404 (N_26404,N_22868,N_21790);
nor U26405 (N_26405,N_23143,N_22239);
nor U26406 (N_26406,N_21767,N_22163);
or U26407 (N_26407,N_23652,N_21432);
and U26408 (N_26408,N_22666,N_22077);
or U26409 (N_26409,N_21625,N_23569);
nor U26410 (N_26410,N_23522,N_22338);
nand U26411 (N_26411,N_21462,N_21590);
and U26412 (N_26412,N_22674,N_23966);
or U26413 (N_26413,N_21348,N_22201);
or U26414 (N_26414,N_22026,N_22225);
or U26415 (N_26415,N_22170,N_22427);
xnor U26416 (N_26416,N_22385,N_21082);
nor U26417 (N_26417,N_23761,N_22992);
nor U26418 (N_26418,N_23371,N_21354);
or U26419 (N_26419,N_23700,N_23333);
nand U26420 (N_26420,N_22232,N_21195);
and U26421 (N_26421,N_23236,N_21893);
and U26422 (N_26422,N_23303,N_23405);
nor U26423 (N_26423,N_21898,N_22497);
or U26424 (N_26424,N_21734,N_23159);
and U26425 (N_26425,N_23135,N_21599);
xor U26426 (N_26426,N_21383,N_21740);
xnor U26427 (N_26427,N_23439,N_21708);
and U26428 (N_26428,N_21491,N_23526);
nor U26429 (N_26429,N_23492,N_23521);
nor U26430 (N_26430,N_23918,N_21810);
or U26431 (N_26431,N_22085,N_21157);
nand U26432 (N_26432,N_23869,N_22003);
or U26433 (N_26433,N_22133,N_22289);
or U26434 (N_26434,N_21231,N_23299);
nand U26435 (N_26435,N_23318,N_23514);
xor U26436 (N_26436,N_22772,N_21240);
and U26437 (N_26437,N_22076,N_22934);
nand U26438 (N_26438,N_23800,N_22516);
and U26439 (N_26439,N_22076,N_22154);
nor U26440 (N_26440,N_21008,N_21947);
or U26441 (N_26441,N_22129,N_21654);
nand U26442 (N_26442,N_23733,N_22378);
and U26443 (N_26443,N_21674,N_22736);
and U26444 (N_26444,N_22951,N_22832);
or U26445 (N_26445,N_21476,N_22470);
and U26446 (N_26446,N_21555,N_21176);
and U26447 (N_26447,N_21526,N_22855);
and U26448 (N_26448,N_23722,N_21904);
or U26449 (N_26449,N_22525,N_22415);
and U26450 (N_26450,N_21263,N_22080);
nand U26451 (N_26451,N_22423,N_22915);
and U26452 (N_26452,N_23247,N_23889);
and U26453 (N_26453,N_23684,N_23878);
nor U26454 (N_26454,N_22071,N_23645);
and U26455 (N_26455,N_23175,N_22016);
nand U26456 (N_26456,N_21321,N_22649);
nor U26457 (N_26457,N_22575,N_22972);
and U26458 (N_26458,N_22370,N_23092);
and U26459 (N_26459,N_21108,N_22909);
nand U26460 (N_26460,N_21812,N_23393);
nand U26461 (N_26461,N_23717,N_21645);
or U26462 (N_26462,N_21235,N_21143);
or U26463 (N_26463,N_23357,N_21645);
nor U26464 (N_26464,N_23894,N_21507);
nand U26465 (N_26465,N_22847,N_22110);
or U26466 (N_26466,N_22471,N_22765);
or U26467 (N_26467,N_21608,N_22588);
nand U26468 (N_26468,N_22867,N_21182);
nor U26469 (N_26469,N_21076,N_23050);
or U26470 (N_26470,N_21579,N_22637);
xor U26471 (N_26471,N_22124,N_23157);
or U26472 (N_26472,N_23444,N_21587);
or U26473 (N_26473,N_23557,N_23917);
nor U26474 (N_26474,N_21951,N_21484);
nand U26475 (N_26475,N_21974,N_23704);
nand U26476 (N_26476,N_23291,N_23685);
or U26477 (N_26477,N_22912,N_23825);
nor U26478 (N_26478,N_21656,N_23783);
or U26479 (N_26479,N_21933,N_23268);
and U26480 (N_26480,N_22284,N_21953);
or U26481 (N_26481,N_21364,N_21207);
nor U26482 (N_26482,N_22169,N_22681);
nand U26483 (N_26483,N_23646,N_23527);
nor U26484 (N_26484,N_21436,N_23114);
or U26485 (N_26485,N_22203,N_23269);
nor U26486 (N_26486,N_22591,N_21586);
and U26487 (N_26487,N_21018,N_23230);
and U26488 (N_26488,N_23936,N_23396);
or U26489 (N_26489,N_21688,N_22916);
nand U26490 (N_26490,N_23619,N_23041);
or U26491 (N_26491,N_21882,N_23252);
and U26492 (N_26492,N_22188,N_23431);
nand U26493 (N_26493,N_21345,N_22008);
and U26494 (N_26494,N_21473,N_22592);
nand U26495 (N_26495,N_21089,N_21020);
nor U26496 (N_26496,N_21672,N_22987);
xnor U26497 (N_26497,N_21747,N_23176);
nor U26498 (N_26498,N_23783,N_23186);
nand U26499 (N_26499,N_23446,N_22964);
or U26500 (N_26500,N_22115,N_21175);
and U26501 (N_26501,N_21533,N_23843);
xor U26502 (N_26502,N_21473,N_21830);
nor U26503 (N_26503,N_21312,N_22112);
xor U26504 (N_26504,N_23874,N_23533);
and U26505 (N_26505,N_21992,N_22547);
xor U26506 (N_26506,N_23431,N_23565);
nand U26507 (N_26507,N_23946,N_22976);
nand U26508 (N_26508,N_22450,N_21559);
or U26509 (N_26509,N_21763,N_22322);
nor U26510 (N_26510,N_22947,N_23324);
or U26511 (N_26511,N_23945,N_21835);
xnor U26512 (N_26512,N_21327,N_23280);
nand U26513 (N_26513,N_21748,N_22865);
nand U26514 (N_26514,N_21467,N_21413);
and U26515 (N_26515,N_22533,N_22908);
nand U26516 (N_26516,N_21891,N_23127);
and U26517 (N_26517,N_21853,N_21196);
nand U26518 (N_26518,N_21050,N_21063);
or U26519 (N_26519,N_22468,N_22202);
nand U26520 (N_26520,N_23476,N_22877);
or U26521 (N_26521,N_23296,N_23918);
and U26522 (N_26522,N_21691,N_22178);
nand U26523 (N_26523,N_21521,N_21982);
or U26524 (N_26524,N_21143,N_23888);
nor U26525 (N_26525,N_21904,N_23062);
nor U26526 (N_26526,N_23618,N_21948);
and U26527 (N_26527,N_23063,N_23712);
xnor U26528 (N_26528,N_23190,N_22509);
or U26529 (N_26529,N_21788,N_23775);
or U26530 (N_26530,N_21536,N_21300);
and U26531 (N_26531,N_21486,N_21887);
nand U26532 (N_26532,N_23571,N_22821);
or U26533 (N_26533,N_21388,N_22002);
and U26534 (N_26534,N_23728,N_23755);
and U26535 (N_26535,N_22407,N_22320);
nor U26536 (N_26536,N_21306,N_23371);
nor U26537 (N_26537,N_22939,N_23905);
or U26538 (N_26538,N_23079,N_23916);
nand U26539 (N_26539,N_21385,N_22258);
nor U26540 (N_26540,N_22037,N_21276);
or U26541 (N_26541,N_21906,N_21503);
xnor U26542 (N_26542,N_22578,N_21999);
nor U26543 (N_26543,N_22528,N_22691);
nor U26544 (N_26544,N_21247,N_23092);
or U26545 (N_26545,N_21869,N_21330);
nand U26546 (N_26546,N_23005,N_23711);
nand U26547 (N_26547,N_23950,N_21834);
and U26548 (N_26548,N_21534,N_21673);
or U26549 (N_26549,N_22170,N_21094);
nand U26550 (N_26550,N_22550,N_23161);
and U26551 (N_26551,N_22278,N_21034);
nor U26552 (N_26552,N_23700,N_23615);
or U26553 (N_26553,N_23989,N_21268);
nor U26554 (N_26554,N_21404,N_23295);
or U26555 (N_26555,N_21612,N_22076);
and U26556 (N_26556,N_22487,N_23623);
xor U26557 (N_26557,N_23782,N_22719);
nor U26558 (N_26558,N_23130,N_23267);
nand U26559 (N_26559,N_23542,N_23513);
or U26560 (N_26560,N_23279,N_21269);
nor U26561 (N_26561,N_22046,N_23327);
nand U26562 (N_26562,N_21074,N_23778);
or U26563 (N_26563,N_22387,N_22232);
or U26564 (N_26564,N_21456,N_21353);
xnor U26565 (N_26565,N_23082,N_21626);
nand U26566 (N_26566,N_23548,N_21957);
xor U26567 (N_26567,N_21673,N_22599);
nor U26568 (N_26568,N_22258,N_22104);
nand U26569 (N_26569,N_22462,N_21538);
and U26570 (N_26570,N_23619,N_22579);
nor U26571 (N_26571,N_22795,N_22285);
and U26572 (N_26572,N_21679,N_21653);
or U26573 (N_26573,N_21145,N_21640);
and U26574 (N_26574,N_22683,N_22052);
or U26575 (N_26575,N_23983,N_23577);
xnor U26576 (N_26576,N_23800,N_23494);
nand U26577 (N_26577,N_23324,N_23793);
nand U26578 (N_26578,N_22059,N_23221);
nand U26579 (N_26579,N_23222,N_21525);
and U26580 (N_26580,N_22256,N_22185);
or U26581 (N_26581,N_23996,N_22480);
and U26582 (N_26582,N_22870,N_23970);
nor U26583 (N_26583,N_23466,N_21625);
nand U26584 (N_26584,N_21013,N_21660);
or U26585 (N_26585,N_21464,N_21227);
nor U26586 (N_26586,N_22627,N_21465);
or U26587 (N_26587,N_23796,N_22376);
or U26588 (N_26588,N_22750,N_22320);
and U26589 (N_26589,N_21660,N_21292);
and U26590 (N_26590,N_23170,N_22912);
xor U26591 (N_26591,N_23643,N_23092);
or U26592 (N_26592,N_23721,N_22351);
nor U26593 (N_26593,N_22969,N_21339);
or U26594 (N_26594,N_21437,N_23330);
nand U26595 (N_26595,N_23692,N_21974);
and U26596 (N_26596,N_23399,N_22770);
or U26597 (N_26597,N_21611,N_21103);
and U26598 (N_26598,N_21967,N_22273);
xnor U26599 (N_26599,N_21349,N_21348);
nor U26600 (N_26600,N_22251,N_23530);
or U26601 (N_26601,N_21785,N_23516);
nand U26602 (N_26602,N_22769,N_21175);
nand U26603 (N_26603,N_22429,N_22407);
nor U26604 (N_26604,N_22657,N_22545);
or U26605 (N_26605,N_23876,N_22931);
or U26606 (N_26606,N_22580,N_22436);
xnor U26607 (N_26607,N_21154,N_22965);
or U26608 (N_26608,N_22447,N_23220);
and U26609 (N_26609,N_22566,N_21550);
xnor U26610 (N_26610,N_22941,N_21601);
nor U26611 (N_26611,N_22488,N_23502);
and U26612 (N_26612,N_22152,N_22353);
or U26613 (N_26613,N_21187,N_23357);
nor U26614 (N_26614,N_22760,N_22222);
nand U26615 (N_26615,N_23518,N_21656);
nor U26616 (N_26616,N_21495,N_23366);
nor U26617 (N_26617,N_21551,N_23251);
nor U26618 (N_26618,N_21176,N_21467);
xnor U26619 (N_26619,N_23655,N_23493);
nor U26620 (N_26620,N_21362,N_21690);
nor U26621 (N_26621,N_22364,N_21555);
or U26622 (N_26622,N_22420,N_21065);
or U26623 (N_26623,N_23506,N_22337);
or U26624 (N_26624,N_23465,N_23032);
nand U26625 (N_26625,N_22235,N_23264);
nand U26626 (N_26626,N_22557,N_23853);
nand U26627 (N_26627,N_23096,N_21295);
nand U26628 (N_26628,N_22702,N_22672);
nor U26629 (N_26629,N_22600,N_21085);
and U26630 (N_26630,N_23051,N_23890);
and U26631 (N_26631,N_21120,N_22832);
or U26632 (N_26632,N_23541,N_23434);
nand U26633 (N_26633,N_22870,N_22110);
nand U26634 (N_26634,N_21847,N_23380);
and U26635 (N_26635,N_21380,N_23637);
or U26636 (N_26636,N_21954,N_21791);
xnor U26637 (N_26637,N_21859,N_23776);
nor U26638 (N_26638,N_23751,N_23623);
or U26639 (N_26639,N_21667,N_21367);
nand U26640 (N_26640,N_21206,N_23615);
and U26641 (N_26641,N_23965,N_21451);
or U26642 (N_26642,N_23344,N_23699);
nor U26643 (N_26643,N_23418,N_23273);
and U26644 (N_26644,N_22486,N_21775);
or U26645 (N_26645,N_23482,N_22394);
and U26646 (N_26646,N_22736,N_22829);
and U26647 (N_26647,N_22825,N_23991);
and U26648 (N_26648,N_23158,N_21363);
and U26649 (N_26649,N_22086,N_21830);
nand U26650 (N_26650,N_22907,N_22610);
or U26651 (N_26651,N_22697,N_23739);
nand U26652 (N_26652,N_21480,N_23004);
nor U26653 (N_26653,N_21666,N_22736);
nor U26654 (N_26654,N_22823,N_23048);
or U26655 (N_26655,N_23876,N_22075);
and U26656 (N_26656,N_22570,N_22435);
nor U26657 (N_26657,N_21752,N_22048);
nor U26658 (N_26658,N_23023,N_23183);
nor U26659 (N_26659,N_21947,N_21663);
nor U26660 (N_26660,N_23041,N_23753);
or U26661 (N_26661,N_23371,N_21634);
and U26662 (N_26662,N_22297,N_21091);
nand U26663 (N_26663,N_21744,N_23722);
nor U26664 (N_26664,N_23412,N_23871);
nor U26665 (N_26665,N_21265,N_22830);
nor U26666 (N_26666,N_22072,N_23734);
and U26667 (N_26667,N_21665,N_21673);
and U26668 (N_26668,N_22509,N_22051);
or U26669 (N_26669,N_23089,N_23277);
nor U26670 (N_26670,N_23672,N_22997);
nor U26671 (N_26671,N_22977,N_22784);
nor U26672 (N_26672,N_23818,N_21323);
or U26673 (N_26673,N_23232,N_22031);
xor U26674 (N_26674,N_23973,N_21315);
nor U26675 (N_26675,N_21226,N_23989);
nand U26676 (N_26676,N_22487,N_21314);
nor U26677 (N_26677,N_21197,N_23212);
and U26678 (N_26678,N_21184,N_22093);
or U26679 (N_26679,N_21663,N_23584);
nand U26680 (N_26680,N_21059,N_23428);
or U26681 (N_26681,N_23292,N_22208);
and U26682 (N_26682,N_22395,N_22572);
nor U26683 (N_26683,N_22927,N_23476);
nand U26684 (N_26684,N_21815,N_21002);
or U26685 (N_26685,N_21775,N_23713);
or U26686 (N_26686,N_22713,N_23656);
xor U26687 (N_26687,N_22435,N_22957);
or U26688 (N_26688,N_22966,N_23342);
or U26689 (N_26689,N_23472,N_23923);
or U26690 (N_26690,N_23747,N_22376);
nor U26691 (N_26691,N_22866,N_23478);
or U26692 (N_26692,N_22387,N_23032);
xor U26693 (N_26693,N_22646,N_23033);
xnor U26694 (N_26694,N_23004,N_21364);
nor U26695 (N_26695,N_23633,N_22167);
and U26696 (N_26696,N_22095,N_23386);
nand U26697 (N_26697,N_22861,N_23805);
xnor U26698 (N_26698,N_22569,N_22842);
and U26699 (N_26699,N_23709,N_21196);
or U26700 (N_26700,N_23241,N_21974);
nor U26701 (N_26701,N_23277,N_21051);
nor U26702 (N_26702,N_21459,N_23988);
nor U26703 (N_26703,N_22610,N_22852);
nand U26704 (N_26704,N_21830,N_22627);
and U26705 (N_26705,N_23771,N_21808);
and U26706 (N_26706,N_21434,N_21822);
nor U26707 (N_26707,N_23441,N_22802);
nor U26708 (N_26708,N_23904,N_22283);
nand U26709 (N_26709,N_21034,N_21706);
nand U26710 (N_26710,N_21068,N_22759);
xor U26711 (N_26711,N_22527,N_22785);
nor U26712 (N_26712,N_23191,N_23314);
or U26713 (N_26713,N_22558,N_21152);
or U26714 (N_26714,N_22998,N_21898);
nor U26715 (N_26715,N_21730,N_23342);
nand U26716 (N_26716,N_21824,N_23552);
or U26717 (N_26717,N_21992,N_21431);
or U26718 (N_26718,N_22961,N_21308);
nand U26719 (N_26719,N_22425,N_22647);
and U26720 (N_26720,N_22006,N_22939);
and U26721 (N_26721,N_22921,N_23442);
or U26722 (N_26722,N_22795,N_21582);
or U26723 (N_26723,N_23693,N_22855);
nor U26724 (N_26724,N_21684,N_22226);
nand U26725 (N_26725,N_22804,N_21242);
nand U26726 (N_26726,N_23552,N_21440);
nor U26727 (N_26727,N_23015,N_23148);
and U26728 (N_26728,N_23893,N_22832);
nand U26729 (N_26729,N_22243,N_21752);
and U26730 (N_26730,N_22012,N_22242);
nor U26731 (N_26731,N_22385,N_22795);
nor U26732 (N_26732,N_22928,N_23690);
nor U26733 (N_26733,N_21408,N_21088);
xor U26734 (N_26734,N_23512,N_23474);
nor U26735 (N_26735,N_23880,N_21888);
nand U26736 (N_26736,N_21257,N_23518);
nand U26737 (N_26737,N_23010,N_21072);
and U26738 (N_26738,N_23357,N_23226);
or U26739 (N_26739,N_21626,N_23766);
nor U26740 (N_26740,N_21146,N_22358);
nor U26741 (N_26741,N_22618,N_23777);
nor U26742 (N_26742,N_21457,N_21669);
nor U26743 (N_26743,N_23810,N_23428);
nand U26744 (N_26744,N_22387,N_22867);
nor U26745 (N_26745,N_22119,N_23494);
nor U26746 (N_26746,N_22207,N_21175);
and U26747 (N_26747,N_23551,N_22174);
xnor U26748 (N_26748,N_21392,N_21296);
xnor U26749 (N_26749,N_21243,N_23354);
and U26750 (N_26750,N_23397,N_22985);
or U26751 (N_26751,N_22208,N_23255);
and U26752 (N_26752,N_22401,N_22495);
or U26753 (N_26753,N_22766,N_22145);
and U26754 (N_26754,N_22168,N_22418);
or U26755 (N_26755,N_23884,N_21764);
or U26756 (N_26756,N_22969,N_21996);
and U26757 (N_26757,N_22467,N_21592);
xor U26758 (N_26758,N_23217,N_23112);
nand U26759 (N_26759,N_21594,N_22182);
and U26760 (N_26760,N_22071,N_23141);
or U26761 (N_26761,N_21412,N_22584);
and U26762 (N_26762,N_23145,N_23448);
or U26763 (N_26763,N_22992,N_22386);
nor U26764 (N_26764,N_23935,N_23995);
nor U26765 (N_26765,N_22844,N_21595);
or U26766 (N_26766,N_22365,N_22534);
nor U26767 (N_26767,N_23680,N_22924);
and U26768 (N_26768,N_23965,N_23510);
nor U26769 (N_26769,N_21779,N_21241);
nor U26770 (N_26770,N_21306,N_23211);
nand U26771 (N_26771,N_23068,N_22445);
nand U26772 (N_26772,N_23220,N_21318);
nand U26773 (N_26773,N_23526,N_21214);
nor U26774 (N_26774,N_23890,N_21599);
nand U26775 (N_26775,N_22694,N_21082);
nand U26776 (N_26776,N_22723,N_22601);
nor U26777 (N_26777,N_21712,N_21044);
or U26778 (N_26778,N_23250,N_21750);
and U26779 (N_26779,N_22404,N_22289);
nor U26780 (N_26780,N_22622,N_23436);
and U26781 (N_26781,N_21346,N_22968);
xor U26782 (N_26782,N_21199,N_23148);
nor U26783 (N_26783,N_22037,N_23750);
nor U26784 (N_26784,N_21809,N_22643);
nand U26785 (N_26785,N_22050,N_22601);
nand U26786 (N_26786,N_23273,N_21221);
nand U26787 (N_26787,N_22749,N_21192);
nand U26788 (N_26788,N_23931,N_23895);
nand U26789 (N_26789,N_23578,N_22127);
xor U26790 (N_26790,N_21163,N_23509);
and U26791 (N_26791,N_23369,N_22018);
or U26792 (N_26792,N_23633,N_22431);
nor U26793 (N_26793,N_21674,N_22834);
nor U26794 (N_26794,N_21316,N_22237);
and U26795 (N_26795,N_23748,N_22231);
or U26796 (N_26796,N_23896,N_23842);
nand U26797 (N_26797,N_21060,N_21988);
and U26798 (N_26798,N_23354,N_23630);
nor U26799 (N_26799,N_23215,N_22623);
or U26800 (N_26800,N_22796,N_22730);
xor U26801 (N_26801,N_23308,N_23008);
and U26802 (N_26802,N_22084,N_23528);
xnor U26803 (N_26803,N_21832,N_21754);
or U26804 (N_26804,N_23641,N_21004);
or U26805 (N_26805,N_22332,N_23991);
and U26806 (N_26806,N_21054,N_21041);
or U26807 (N_26807,N_23677,N_21349);
nor U26808 (N_26808,N_22900,N_23330);
and U26809 (N_26809,N_21262,N_22248);
or U26810 (N_26810,N_23574,N_21361);
nor U26811 (N_26811,N_21514,N_21645);
xor U26812 (N_26812,N_22563,N_23829);
xnor U26813 (N_26813,N_22794,N_23150);
nor U26814 (N_26814,N_23651,N_21904);
nand U26815 (N_26815,N_21541,N_21692);
nor U26816 (N_26816,N_23407,N_21909);
nand U26817 (N_26817,N_22204,N_21262);
and U26818 (N_26818,N_23981,N_21158);
nor U26819 (N_26819,N_23049,N_23432);
nand U26820 (N_26820,N_21172,N_22727);
nand U26821 (N_26821,N_21980,N_21566);
or U26822 (N_26822,N_23707,N_21631);
nand U26823 (N_26823,N_22330,N_23576);
and U26824 (N_26824,N_23802,N_22368);
nand U26825 (N_26825,N_22558,N_23386);
xor U26826 (N_26826,N_23168,N_21873);
xor U26827 (N_26827,N_22106,N_21521);
xor U26828 (N_26828,N_21498,N_23051);
xnor U26829 (N_26829,N_22325,N_21579);
nand U26830 (N_26830,N_22195,N_21481);
and U26831 (N_26831,N_21393,N_22135);
nor U26832 (N_26832,N_22171,N_23947);
and U26833 (N_26833,N_22460,N_23286);
or U26834 (N_26834,N_21032,N_23032);
nor U26835 (N_26835,N_23260,N_22675);
and U26836 (N_26836,N_23449,N_22386);
and U26837 (N_26837,N_21982,N_23518);
nand U26838 (N_26838,N_21662,N_22885);
xor U26839 (N_26839,N_22881,N_22676);
xor U26840 (N_26840,N_21076,N_23305);
nor U26841 (N_26841,N_22158,N_22927);
and U26842 (N_26842,N_23571,N_22697);
or U26843 (N_26843,N_22806,N_23057);
and U26844 (N_26844,N_21031,N_21404);
or U26845 (N_26845,N_22773,N_21547);
or U26846 (N_26846,N_23602,N_22186);
or U26847 (N_26847,N_22278,N_23655);
nor U26848 (N_26848,N_22615,N_22650);
nand U26849 (N_26849,N_22824,N_23959);
or U26850 (N_26850,N_22306,N_22720);
nor U26851 (N_26851,N_23441,N_23109);
or U26852 (N_26852,N_23272,N_22770);
and U26853 (N_26853,N_22199,N_21788);
nor U26854 (N_26854,N_22885,N_21282);
and U26855 (N_26855,N_22995,N_22955);
or U26856 (N_26856,N_23409,N_22427);
or U26857 (N_26857,N_22787,N_22881);
or U26858 (N_26858,N_22182,N_22289);
xor U26859 (N_26859,N_22220,N_23385);
and U26860 (N_26860,N_22952,N_23382);
nor U26861 (N_26861,N_21369,N_22032);
nor U26862 (N_26862,N_22826,N_21979);
nor U26863 (N_26863,N_22844,N_21474);
and U26864 (N_26864,N_21234,N_21058);
or U26865 (N_26865,N_22599,N_21236);
or U26866 (N_26866,N_22342,N_23769);
and U26867 (N_26867,N_21336,N_21227);
or U26868 (N_26868,N_21662,N_21129);
or U26869 (N_26869,N_23385,N_23664);
nand U26870 (N_26870,N_22320,N_21653);
or U26871 (N_26871,N_21416,N_23849);
xnor U26872 (N_26872,N_21817,N_23976);
nor U26873 (N_26873,N_23610,N_21065);
nor U26874 (N_26874,N_22310,N_23883);
or U26875 (N_26875,N_22997,N_21869);
or U26876 (N_26876,N_23559,N_23575);
or U26877 (N_26877,N_21772,N_21912);
nor U26878 (N_26878,N_22801,N_21451);
and U26879 (N_26879,N_21221,N_22594);
nand U26880 (N_26880,N_22118,N_22533);
nand U26881 (N_26881,N_21051,N_21311);
nor U26882 (N_26882,N_22758,N_23529);
nand U26883 (N_26883,N_22177,N_21154);
or U26884 (N_26884,N_22148,N_23335);
and U26885 (N_26885,N_21398,N_21845);
nand U26886 (N_26886,N_21039,N_23958);
nand U26887 (N_26887,N_21627,N_23735);
or U26888 (N_26888,N_23236,N_21603);
nand U26889 (N_26889,N_21381,N_22393);
nor U26890 (N_26890,N_23695,N_23177);
nor U26891 (N_26891,N_21959,N_22949);
nand U26892 (N_26892,N_21739,N_22896);
or U26893 (N_26893,N_22614,N_22430);
or U26894 (N_26894,N_22055,N_23790);
and U26895 (N_26895,N_22479,N_23088);
xor U26896 (N_26896,N_22436,N_23727);
nand U26897 (N_26897,N_23849,N_21152);
nor U26898 (N_26898,N_23129,N_22738);
nand U26899 (N_26899,N_21528,N_21553);
xor U26900 (N_26900,N_21294,N_22893);
or U26901 (N_26901,N_21609,N_21370);
nor U26902 (N_26902,N_21972,N_23755);
xor U26903 (N_26903,N_21021,N_23590);
and U26904 (N_26904,N_23372,N_21728);
nand U26905 (N_26905,N_21921,N_23733);
nor U26906 (N_26906,N_21528,N_22576);
and U26907 (N_26907,N_23847,N_22385);
or U26908 (N_26908,N_22354,N_21171);
nand U26909 (N_26909,N_22891,N_21823);
nand U26910 (N_26910,N_22231,N_23524);
and U26911 (N_26911,N_21427,N_22925);
or U26912 (N_26912,N_22966,N_23846);
nand U26913 (N_26913,N_22692,N_23808);
nor U26914 (N_26914,N_22480,N_23593);
and U26915 (N_26915,N_23046,N_23027);
and U26916 (N_26916,N_22231,N_22000);
nand U26917 (N_26917,N_22472,N_23686);
and U26918 (N_26918,N_21483,N_21741);
nor U26919 (N_26919,N_23542,N_21638);
and U26920 (N_26920,N_21273,N_22653);
nand U26921 (N_26921,N_21242,N_22829);
nand U26922 (N_26922,N_21906,N_22590);
nand U26923 (N_26923,N_23337,N_22215);
xnor U26924 (N_26924,N_21972,N_22159);
nor U26925 (N_26925,N_22470,N_22901);
or U26926 (N_26926,N_23714,N_22345);
nor U26927 (N_26927,N_21022,N_22460);
nor U26928 (N_26928,N_22883,N_22286);
and U26929 (N_26929,N_23395,N_23445);
and U26930 (N_26930,N_21685,N_21011);
or U26931 (N_26931,N_21144,N_22310);
and U26932 (N_26932,N_23745,N_23251);
nor U26933 (N_26933,N_23795,N_21920);
nor U26934 (N_26934,N_22814,N_21184);
and U26935 (N_26935,N_21196,N_23363);
nor U26936 (N_26936,N_23830,N_23335);
and U26937 (N_26937,N_23167,N_23362);
xor U26938 (N_26938,N_23252,N_21146);
or U26939 (N_26939,N_21963,N_21881);
nand U26940 (N_26940,N_23537,N_21452);
nor U26941 (N_26941,N_22059,N_21450);
or U26942 (N_26942,N_23245,N_22930);
xnor U26943 (N_26943,N_23681,N_21692);
nor U26944 (N_26944,N_22180,N_22623);
and U26945 (N_26945,N_21523,N_23423);
nand U26946 (N_26946,N_23803,N_22612);
and U26947 (N_26947,N_23707,N_21589);
nor U26948 (N_26948,N_21612,N_23292);
xor U26949 (N_26949,N_23230,N_23425);
or U26950 (N_26950,N_21827,N_22117);
xnor U26951 (N_26951,N_23546,N_22453);
nor U26952 (N_26952,N_22417,N_22344);
or U26953 (N_26953,N_21909,N_23717);
nand U26954 (N_26954,N_22055,N_22732);
and U26955 (N_26955,N_21786,N_22774);
nor U26956 (N_26956,N_22353,N_22068);
and U26957 (N_26957,N_22885,N_23807);
nor U26958 (N_26958,N_23602,N_22253);
and U26959 (N_26959,N_22243,N_23852);
nor U26960 (N_26960,N_22006,N_21726);
or U26961 (N_26961,N_21711,N_23244);
nand U26962 (N_26962,N_22372,N_23221);
and U26963 (N_26963,N_21049,N_23738);
nor U26964 (N_26964,N_23137,N_21691);
nand U26965 (N_26965,N_23250,N_22247);
or U26966 (N_26966,N_22694,N_22998);
and U26967 (N_26967,N_21669,N_22174);
and U26968 (N_26968,N_22348,N_21848);
and U26969 (N_26969,N_22442,N_23958);
nor U26970 (N_26970,N_21276,N_22062);
nand U26971 (N_26971,N_22000,N_23548);
xor U26972 (N_26972,N_21780,N_22433);
nand U26973 (N_26973,N_23746,N_23768);
xnor U26974 (N_26974,N_21803,N_22087);
nand U26975 (N_26975,N_21198,N_22711);
and U26976 (N_26976,N_23323,N_23801);
nor U26977 (N_26977,N_23101,N_21172);
or U26978 (N_26978,N_21902,N_22609);
and U26979 (N_26979,N_21350,N_21933);
nor U26980 (N_26980,N_21789,N_21062);
nand U26981 (N_26981,N_21608,N_23179);
nor U26982 (N_26982,N_21120,N_23422);
and U26983 (N_26983,N_21976,N_23553);
and U26984 (N_26984,N_21699,N_22387);
nor U26985 (N_26985,N_23198,N_21586);
nor U26986 (N_26986,N_22299,N_21986);
and U26987 (N_26987,N_22336,N_22418);
or U26988 (N_26988,N_21694,N_22383);
nand U26989 (N_26989,N_22370,N_21117);
nand U26990 (N_26990,N_23182,N_22308);
xor U26991 (N_26991,N_21622,N_23518);
and U26992 (N_26992,N_23168,N_21426);
xor U26993 (N_26993,N_22696,N_22001);
or U26994 (N_26994,N_22917,N_22097);
nand U26995 (N_26995,N_22933,N_21135);
or U26996 (N_26996,N_21210,N_22196);
or U26997 (N_26997,N_22937,N_23766);
or U26998 (N_26998,N_22164,N_22134);
and U26999 (N_26999,N_22995,N_23707);
nand U27000 (N_27000,N_24504,N_25584);
nor U27001 (N_27001,N_24732,N_25146);
nand U27002 (N_27002,N_25736,N_26186);
nor U27003 (N_27003,N_26866,N_26678);
and U27004 (N_27004,N_26403,N_25130);
or U27005 (N_27005,N_25538,N_26728);
xor U27006 (N_27006,N_26995,N_26843);
nand U27007 (N_27007,N_25669,N_25479);
or U27008 (N_27008,N_24740,N_26423);
and U27009 (N_27009,N_25650,N_25104);
nor U27010 (N_27010,N_24897,N_25340);
or U27011 (N_27011,N_25115,N_25370);
or U27012 (N_27012,N_25872,N_24491);
or U27013 (N_27013,N_26558,N_25785);
nor U27014 (N_27014,N_24852,N_24091);
or U27015 (N_27015,N_24139,N_24649);
xor U27016 (N_27016,N_25621,N_24945);
nor U27017 (N_27017,N_26431,N_24238);
nand U27018 (N_27018,N_24900,N_26551);
and U27019 (N_27019,N_26677,N_26424);
and U27020 (N_27020,N_24735,N_25038);
nand U27021 (N_27021,N_26791,N_26545);
or U27022 (N_27022,N_24212,N_25577);
nor U27023 (N_27023,N_25176,N_26386);
nor U27024 (N_27024,N_24145,N_25218);
or U27025 (N_27025,N_25452,N_24709);
or U27026 (N_27026,N_26406,N_25599);
nor U27027 (N_27027,N_26065,N_26364);
xnor U27028 (N_27028,N_25738,N_24357);
nor U27029 (N_27029,N_26407,N_25786);
nor U27030 (N_27030,N_24921,N_25014);
and U27031 (N_27031,N_24330,N_24194);
xnor U27032 (N_27032,N_26648,N_25744);
or U27033 (N_27033,N_24669,N_24997);
nand U27034 (N_27034,N_25983,N_24154);
xor U27035 (N_27035,N_24049,N_25398);
and U27036 (N_27036,N_25093,N_25583);
nor U27037 (N_27037,N_25234,N_26183);
and U27038 (N_27038,N_26654,N_26565);
or U27039 (N_27039,N_25002,N_24213);
nand U27040 (N_27040,N_25391,N_25593);
and U27041 (N_27041,N_24152,N_26026);
nand U27042 (N_27042,N_24946,N_24097);
nand U27043 (N_27043,N_25450,N_25019);
nand U27044 (N_27044,N_24363,N_26979);
or U27045 (N_27045,N_25823,N_25609);
nor U27046 (N_27046,N_25148,N_25498);
nor U27047 (N_27047,N_25525,N_24959);
or U27048 (N_27048,N_24260,N_25890);
and U27049 (N_27049,N_26753,N_26780);
or U27050 (N_27050,N_24231,N_24808);
nor U27051 (N_27051,N_26361,N_24624);
xor U27052 (N_27052,N_26328,N_25341);
nor U27053 (N_27053,N_26923,N_25062);
xnor U27054 (N_27054,N_24784,N_26211);
nor U27055 (N_27055,N_25974,N_25631);
or U27056 (N_27056,N_25371,N_25718);
nand U27057 (N_27057,N_26299,N_25368);
or U27058 (N_27058,N_24632,N_26835);
nor U27059 (N_27059,N_25421,N_25702);
nor U27060 (N_27060,N_24009,N_24613);
nor U27061 (N_27061,N_25161,N_25318);
and U27062 (N_27062,N_25681,N_26850);
xnor U27063 (N_27063,N_25292,N_26461);
and U27064 (N_27064,N_25249,N_24289);
nor U27065 (N_27065,N_26176,N_24577);
nand U27066 (N_27066,N_25505,N_25187);
and U27067 (N_27067,N_24058,N_25815);
xor U27068 (N_27068,N_24418,N_25261);
nand U27069 (N_27069,N_25534,N_25747);
nand U27070 (N_27070,N_25385,N_25544);
and U27071 (N_27071,N_24114,N_26153);
nand U27072 (N_27072,N_24383,N_24739);
nand U27073 (N_27073,N_24439,N_24667);
or U27074 (N_27074,N_25833,N_25588);
nand U27075 (N_27075,N_26974,N_26944);
and U27076 (N_27076,N_25199,N_26067);
and U27077 (N_27077,N_24606,N_26968);
or U27078 (N_27078,N_25539,N_26707);
and U27079 (N_27079,N_25745,N_24720);
nand U27080 (N_27080,N_24377,N_25485);
nor U27081 (N_27081,N_25826,N_24521);
nand U27082 (N_27082,N_24636,N_24074);
nand U27083 (N_27083,N_26945,N_24053);
or U27084 (N_27084,N_26370,N_25726);
nand U27085 (N_27085,N_24863,N_24711);
or U27086 (N_27086,N_25020,N_25016);
nor U27087 (N_27087,N_25004,N_25540);
or U27088 (N_27088,N_25694,N_24722);
nand U27089 (N_27089,N_24648,N_25478);
and U27090 (N_27090,N_24218,N_25152);
or U27091 (N_27091,N_26720,N_25467);
and U27092 (N_27092,N_26468,N_24036);
nor U27093 (N_27093,N_26820,N_24562);
or U27094 (N_27094,N_25862,N_26520);
or U27095 (N_27095,N_26323,N_25801);
nand U27096 (N_27096,N_26773,N_25388);
nand U27097 (N_27097,N_24136,N_26643);
and U27098 (N_27098,N_25784,N_24535);
or U27099 (N_27099,N_24005,N_24542);
nand U27100 (N_27100,N_24887,N_25873);
nor U27101 (N_27101,N_25759,N_24858);
nand U27102 (N_27102,N_26957,N_24890);
nor U27103 (N_27103,N_24021,N_26268);
nor U27104 (N_27104,N_25437,N_26693);
nand U27105 (N_27105,N_24666,N_25289);
and U27106 (N_27106,N_25773,N_24634);
nor U27107 (N_27107,N_26870,N_26795);
nor U27108 (N_27108,N_25290,N_24083);
nand U27109 (N_27109,N_25231,N_26589);
nand U27110 (N_27110,N_26725,N_25931);
nor U27111 (N_27111,N_25838,N_25326);
or U27112 (N_27112,N_25765,N_24790);
nor U27113 (N_27113,N_26683,N_26803);
nand U27114 (N_27114,N_24826,N_26929);
or U27115 (N_27115,N_26642,N_26527);
nand U27116 (N_27116,N_26383,N_24864);
and U27117 (N_27117,N_24293,N_25095);
or U27118 (N_27118,N_24037,N_26477);
nand U27119 (N_27119,N_25915,N_25114);
xnor U27120 (N_27120,N_24108,N_25822);
nor U27121 (N_27121,N_26482,N_26878);
xor U27122 (N_27122,N_24251,N_26288);
nor U27123 (N_27123,N_25851,N_25715);
or U27124 (N_27124,N_25676,N_26395);
xor U27125 (N_27125,N_24656,N_25783);
and U27126 (N_27126,N_24814,N_24555);
xnor U27127 (N_27127,N_25521,N_26263);
and U27128 (N_27128,N_24726,N_25174);
or U27129 (N_27129,N_26077,N_25628);
and U27130 (N_27130,N_25888,N_26155);
nand U27131 (N_27131,N_25712,N_26733);
nand U27132 (N_27132,N_24170,N_25163);
or U27133 (N_27133,N_25256,N_24873);
or U27134 (N_27134,N_25466,N_24967);
nand U27135 (N_27135,N_25597,N_26682);
and U27136 (N_27136,N_25527,N_24811);
and U27137 (N_27137,N_24962,N_26718);
nand U27138 (N_27138,N_26048,N_26248);
and U27139 (N_27139,N_25419,N_24318);
xor U27140 (N_27140,N_26647,N_25052);
and U27141 (N_27141,N_24322,N_25659);
and U27142 (N_27142,N_25899,N_24423);
nand U27143 (N_27143,N_25168,N_24684);
nand U27144 (N_27144,N_25557,N_26412);
nor U27145 (N_27145,N_25345,N_24766);
nand U27146 (N_27146,N_26189,N_26053);
nor U27147 (N_27147,N_26123,N_24248);
nand U27148 (N_27148,N_26651,N_26840);
nor U27149 (N_27149,N_26076,N_26083);
xor U27150 (N_27150,N_24929,N_26131);
nand U27151 (N_27151,N_26745,N_24940);
nand U27152 (N_27152,N_25253,N_25924);
nand U27153 (N_27153,N_24909,N_25991);
nand U27154 (N_27154,N_26941,N_26860);
and U27155 (N_27155,N_24072,N_24980);
nor U27156 (N_27156,N_24177,N_24285);
and U27157 (N_27157,N_25259,N_24874);
or U27158 (N_27158,N_25435,N_25606);
nor U27159 (N_27159,N_26821,N_25463);
nor U27160 (N_27160,N_26485,N_25275);
nand U27161 (N_27161,N_25845,N_26761);
nand U27162 (N_27162,N_26710,N_25749);
nand U27163 (N_27163,N_24261,N_25528);
xor U27164 (N_27164,N_25775,N_25229);
nor U27165 (N_27165,N_25036,N_25761);
xor U27166 (N_27166,N_26425,N_26830);
or U27167 (N_27167,N_24147,N_25379);
nor U27168 (N_27168,N_25175,N_26627);
xnor U27169 (N_27169,N_25482,N_25280);
or U27170 (N_27170,N_25953,N_26632);
nor U27171 (N_27171,N_26854,N_26798);
and U27172 (N_27172,N_26614,N_24460);
nand U27173 (N_27173,N_24288,N_25999);
nand U27174 (N_27174,N_26719,N_25039);
and U27175 (N_27175,N_24801,N_26254);
xor U27176 (N_27176,N_25150,N_24806);
or U27177 (N_27177,N_24331,N_24111);
nand U27178 (N_27178,N_24938,N_24388);
and U27179 (N_27179,N_25821,N_25415);
or U27180 (N_27180,N_26169,N_24870);
or U27181 (N_27181,N_24197,N_24239);
and U27182 (N_27182,N_25212,N_26980);
nand U27183 (N_27183,N_26797,N_24845);
nand U27184 (N_27184,N_26224,N_24465);
and U27185 (N_27185,N_26991,N_24519);
and U27186 (N_27186,N_25067,N_25751);
xnor U27187 (N_27187,N_24839,N_26448);
and U27188 (N_27188,N_24373,N_24672);
nor U27189 (N_27189,N_24000,N_26905);
nor U27190 (N_27190,N_26063,N_25877);
and U27191 (N_27191,N_26846,N_24633);
and U27192 (N_27192,N_25490,N_26027);
nand U27193 (N_27193,N_24158,N_24923);
and U27194 (N_27194,N_24934,N_25041);
nand U27195 (N_27195,N_24280,N_25118);
nor U27196 (N_27196,N_24242,N_26039);
nor U27197 (N_27197,N_24565,N_24048);
nand U27198 (N_27198,N_26593,N_26289);
nor U27199 (N_27199,N_24983,N_25220);
xor U27200 (N_27200,N_24107,N_26316);
and U27201 (N_27201,N_25687,N_25449);
or U27202 (N_27202,N_25686,N_26368);
nor U27203 (N_27203,N_25812,N_24469);
xor U27204 (N_27204,N_26935,N_24544);
or U27205 (N_27205,N_26298,N_26989);
or U27206 (N_27206,N_26279,N_24159);
nand U27207 (N_27207,N_24155,N_26812);
or U27208 (N_27208,N_26338,N_24570);
or U27209 (N_27209,N_26899,N_25875);
or U27210 (N_27210,N_25003,N_26727);
and U27211 (N_27211,N_24494,N_25278);
xnor U27212 (N_27212,N_24586,N_24226);
and U27213 (N_27213,N_26709,N_24339);
nor U27214 (N_27214,N_24458,N_24384);
and U27215 (N_27215,N_24531,N_25917);
and U27216 (N_27216,N_26774,N_25767);
or U27217 (N_27217,N_26217,N_24138);
xnor U27218 (N_27218,N_24172,N_24440);
nor U27219 (N_27219,N_24392,N_26213);
or U27220 (N_27220,N_25887,N_24654);
nand U27221 (N_27221,N_26985,N_24530);
xnor U27222 (N_27222,N_25075,N_25670);
or U27223 (N_27223,N_24203,N_26743);
or U27224 (N_27224,N_24605,N_24710);
nor U27225 (N_27225,N_26483,N_26195);
nor U27226 (N_27226,N_24413,N_25938);
nand U27227 (N_27227,N_26529,N_26351);
or U27228 (N_27228,N_25630,N_25852);
nand U27229 (N_27229,N_26952,N_25012);
xor U27230 (N_27230,N_24270,N_25087);
nor U27231 (N_27231,N_25354,N_25362);
or U27232 (N_27232,N_26225,N_24335);
nor U27233 (N_27233,N_26926,N_24085);
and U27234 (N_27234,N_24856,N_24575);
nand U27235 (N_27235,N_25835,N_26629);
and U27236 (N_27236,N_25460,N_26928);
or U27237 (N_27237,N_26162,N_26602);
or U27238 (N_27238,N_24210,N_26241);
and U27239 (N_27239,N_25470,N_24976);
nor U27240 (N_27240,N_26635,N_26239);
xnor U27241 (N_27241,N_24034,N_24830);
or U27242 (N_27242,N_25192,N_25941);
nand U27243 (N_27243,N_24958,N_26401);
or U27244 (N_27244,N_25904,N_25017);
and U27245 (N_27245,N_26624,N_24682);
xor U27246 (N_27246,N_26555,N_26817);
or U27247 (N_27247,N_26816,N_24110);
and U27248 (N_27248,N_24217,N_25186);
nor U27249 (N_27249,N_26964,N_25119);
and U27250 (N_27250,N_24611,N_25853);
or U27251 (N_27251,N_26092,N_24397);
nand U27252 (N_27252,N_25181,N_24041);
nand U27253 (N_27253,N_25171,N_26575);
xor U27254 (N_27254,N_25214,N_25423);
and U27255 (N_27255,N_26003,N_25222);
and U27256 (N_27256,N_24370,N_26055);
xnor U27257 (N_27257,N_26937,N_24786);
xnor U27258 (N_27258,N_25572,N_25806);
and U27259 (N_27259,N_25026,N_26746);
or U27260 (N_27260,N_24355,N_26863);
nand U27261 (N_27261,N_26327,N_24961);
and U27262 (N_27262,N_25366,N_25856);
nor U27263 (N_27263,N_26324,N_25475);
or U27264 (N_27264,N_24326,N_25081);
or U27265 (N_27265,N_25264,N_24499);
or U27266 (N_27266,N_26507,N_26531);
nand U27267 (N_27267,N_25982,N_26885);
xnor U27268 (N_27268,N_26621,N_25328);
nor U27269 (N_27269,N_25590,N_25160);
nand U27270 (N_27270,N_25509,N_25978);
nor U27271 (N_27271,N_26024,N_26455);
nor U27272 (N_27272,N_26286,N_25042);
nand U27273 (N_27273,N_26013,N_26559);
nand U27274 (N_27274,N_24733,N_26564);
and U27275 (N_27275,N_26486,N_25934);
nand U27276 (N_27276,N_26690,N_24467);
or U27277 (N_27277,N_24479,N_25740);
nor U27278 (N_27278,N_25513,N_26956);
or U27279 (N_27279,N_26818,N_26842);
nand U27280 (N_27280,N_26523,N_24972);
or U27281 (N_27281,N_24222,N_25811);
xor U27282 (N_27282,N_24804,N_24866);
nand U27283 (N_27283,N_24886,N_26182);
and U27284 (N_27284,N_24680,N_25204);
and U27285 (N_27285,N_26924,N_26269);
nand U27286 (N_27286,N_24595,N_25569);
nor U27287 (N_27287,N_26016,N_24604);
nand U27288 (N_27288,N_26524,N_26150);
nand U27289 (N_27289,N_25595,N_26184);
nor U27290 (N_27290,N_25344,N_24825);
nor U27291 (N_27291,N_25741,N_25357);
nor U27292 (N_27292,N_24442,N_25541);
nand U27293 (N_27293,N_25356,N_25307);
nand U27294 (N_27294,N_26100,N_24968);
or U27295 (N_27295,N_26047,N_24300);
xnor U27296 (N_27296,N_25517,N_24878);
or U27297 (N_27297,N_24496,N_25276);
nand U27298 (N_27298,N_26976,N_26344);
or U27299 (N_27299,N_26156,N_24650);
xor U27300 (N_27300,N_25703,N_24130);
and U27301 (N_27301,N_25350,N_24497);
xor U27302 (N_27302,N_25529,N_24812);
and U27303 (N_27303,N_24396,N_26366);
and U27304 (N_27304,N_25651,N_24779);
or U27305 (N_27305,N_24471,N_25300);
nand U27306 (N_27306,N_24073,N_24411);
nand U27307 (N_27307,N_24834,N_26729);
nor U27308 (N_27308,N_24781,N_24548);
nor U27309 (N_27309,N_26768,N_25589);
and U27310 (N_27310,N_25027,N_26825);
nor U27311 (N_27311,N_25400,N_26416);
and U27312 (N_27312,N_26157,N_25921);
nand U27313 (N_27313,N_26538,N_24061);
nor U27314 (N_27314,N_26634,N_25469);
nor U27315 (N_27315,N_25869,N_26751);
or U27316 (N_27316,N_25837,N_24325);
or U27317 (N_27317,N_24516,N_24892);
and U27318 (N_27318,N_25660,N_24931);
nand U27319 (N_27319,N_26235,N_24895);
or U27320 (N_27320,N_26265,N_25262);
xor U27321 (N_27321,N_26561,N_25916);
or U27322 (N_27322,N_24902,N_26574);
nor U27323 (N_27323,N_24459,N_25946);
xor U27324 (N_27324,N_26392,N_25602);
or U27325 (N_27325,N_25442,N_26367);
xor U27326 (N_27326,N_25009,N_26847);
nor U27327 (N_27327,N_24725,N_26017);
nor U27328 (N_27328,N_24894,N_26603);
and U27329 (N_27329,N_26726,N_25136);
or U27330 (N_27330,N_25793,N_25549);
nor U27331 (N_27331,N_26947,N_26560);
and U27332 (N_27332,N_25241,N_24615);
and U27333 (N_27333,N_24679,N_24428);
nor U27334 (N_27334,N_24328,N_24303);
nor U27335 (N_27335,N_25263,N_25349);
xor U27336 (N_27336,N_26916,N_25070);
or U27337 (N_27337,N_24712,N_26303);
nand U27338 (N_27338,N_25827,N_25361);
xor U27339 (N_27339,N_24284,N_25184);
and U27340 (N_27340,N_24332,N_25975);
nand U27341 (N_27341,N_25179,N_26029);
nor U27342 (N_27342,N_24059,N_26948);
nand U27343 (N_27343,N_26072,N_26623);
and U27344 (N_27344,N_26390,N_25792);
nor U27345 (N_27345,N_26573,N_24584);
xnor U27346 (N_27346,N_26925,N_24556);
or U27347 (N_27347,N_24143,N_24872);
and U27348 (N_27348,N_26539,N_24118);
nand U27349 (N_27349,N_24574,N_26806);
xnor U27350 (N_27350,N_26496,N_25834);
nand U27351 (N_27351,N_25059,N_26626);
nand U27352 (N_27352,N_24693,N_26480);
or U27353 (N_27353,N_26236,N_24241);
and U27354 (N_27354,N_24175,N_25386);
nand U27355 (N_27355,N_25126,N_25024);
nor U27356 (N_27356,N_25867,N_26345);
xnor U27357 (N_27357,N_25447,N_26692);
or U27358 (N_27358,N_24778,N_26095);
and U27359 (N_27359,N_25291,N_26737);
or U27360 (N_27360,N_25560,N_24630);
xor U27361 (N_27361,N_24823,N_25501);
nand U27362 (N_27362,N_24445,N_25173);
or U27363 (N_27363,N_25418,N_24743);
or U27364 (N_27364,N_25188,N_24153);
and U27365 (N_27365,N_26101,N_26240);
or U27366 (N_27366,N_25518,N_26414);
and U27367 (N_27367,N_26877,N_24977);
and U27368 (N_27368,N_24951,N_24865);
nand U27369 (N_27369,N_25891,N_26904);
nor U27370 (N_27370,N_25170,N_25496);
nor U27371 (N_27371,N_25769,N_25486);
nor U27372 (N_27372,N_25295,N_24879);
and U27373 (N_27373,N_26919,N_26384);
nand U27374 (N_27374,N_25566,N_25780);
nand U27375 (N_27375,N_24686,N_26554);
and U27376 (N_27376,N_25607,N_26584);
nand U27377 (N_27377,N_26911,N_26158);
and U27378 (N_27378,N_25074,N_24821);
and U27379 (N_27379,N_24244,N_26967);
or U27380 (N_27380,N_24131,N_24358);
and U27381 (N_27381,N_24532,N_25582);
nor U27382 (N_27382,N_24398,N_25010);
and U27383 (N_27383,N_25255,N_26571);
xnor U27384 (N_27384,N_26826,N_24974);
nor U27385 (N_27385,N_26867,N_24279);
or U27386 (N_27386,N_26108,N_24514);
nand U27387 (N_27387,N_26848,N_24768);
nand U27388 (N_27388,N_26417,N_25436);
nand U27389 (N_27389,N_26159,N_26884);
and U27390 (N_27390,N_25299,N_24117);
and U27391 (N_27391,N_25412,N_26580);
nor U27392 (N_27392,N_26618,N_25704);
nor U27393 (N_27393,N_25491,N_26596);
or U27394 (N_27394,N_26740,N_25454);
or U27395 (N_27395,N_24321,N_24035);
nand U27396 (N_27396,N_25992,N_24381);
nor U27397 (N_27397,N_25816,N_24472);
xor U27398 (N_27398,N_24783,N_24193);
nand U27399 (N_27399,N_24068,N_24166);
nor U27400 (N_27400,N_24142,N_25409);
xnor U27401 (N_27401,N_24849,N_25661);
and U27402 (N_27402,N_24290,N_26936);
and U27403 (N_27403,N_24375,N_24291);
or U27404 (N_27404,N_26106,N_25481);
and U27405 (N_27405,N_26413,N_24190);
and U27406 (N_27406,N_26232,N_25193);
and U27407 (N_27407,N_24387,N_26231);
xnor U27408 (N_27408,N_25839,N_26702);
nand U27409 (N_27409,N_24071,N_25579);
nor U27410 (N_27410,N_24718,N_25427);
and U27411 (N_27411,N_25266,N_24016);
or U27412 (N_27412,N_26018,N_25313);
xor U27413 (N_27413,N_25734,N_26649);
nor U27414 (N_27414,N_26715,N_24207);
nor U27415 (N_27415,N_26285,N_26191);
or U27416 (N_27416,N_26234,N_24956);
and U27417 (N_27417,N_26363,N_25503);
and U27418 (N_27418,N_26051,N_25764);
nand U27419 (N_27419,N_25526,N_26205);
nor U27420 (N_27420,N_25376,N_24341);
and U27421 (N_27421,N_24753,N_26317);
nand U27422 (N_27422,N_25265,N_24343);
nand U27423 (N_27423,N_26148,N_25476);
nand U27424 (N_27424,N_25757,N_24463);
and U27425 (N_27425,N_24716,N_26282);
and U27426 (N_27426,N_26958,N_26275);
nand U27427 (N_27427,N_26022,N_24127);
or U27428 (N_27428,N_26291,N_24581);
nor U27429 (N_27429,N_24827,N_26853);
nor U27430 (N_27430,N_26177,N_24196);
xnor U27431 (N_27431,N_24729,N_25157);
or U27432 (N_27432,N_25406,N_24706);
nor U27433 (N_27433,N_26732,N_24149);
nor U27434 (N_27434,N_26829,N_25322);
nor U27435 (N_27435,N_24018,N_24017);
nor U27436 (N_27436,N_26909,N_24908);
and U27437 (N_27437,N_24425,N_26515);
and U27438 (N_27438,N_26165,N_25373);
or U27439 (N_27439,N_25656,N_24451);
nand U27440 (N_27440,N_26152,N_25183);
xor U27441 (N_27441,N_26784,N_24764);
xnor U27442 (N_27442,N_25558,N_26297);
and U27443 (N_27443,N_24174,N_26378);
xor U27444 (N_27444,N_26717,N_25201);
nand U27445 (N_27445,N_24757,N_25401);
and U27446 (N_27446,N_26498,N_25208);
and U27447 (N_27447,N_25940,N_26404);
nor U27448 (N_27448,N_25304,N_25381);
nor U27449 (N_27449,N_26942,N_26792);
nand U27450 (N_27450,N_24794,N_24868);
and U27451 (N_27451,N_26971,N_25779);
xnor U27452 (N_27452,N_24354,N_24299);
xnor U27453 (N_27453,N_24903,N_26664);
or U27454 (N_27454,N_25760,N_24657);
nor U27455 (N_27455,N_24309,N_26434);
or U27456 (N_27456,N_25968,N_24861);
nor U27457 (N_27457,N_24533,N_24637);
or U27458 (N_27458,N_26568,N_24340);
nor U27459 (N_27459,N_25717,N_25287);
xnor U27460 (N_27460,N_24558,N_24181);
nor U27461 (N_27461,N_25018,N_24503);
xor U27462 (N_27462,N_26075,N_24004);
nand U27463 (N_27463,N_24797,N_24102);
xor U27464 (N_27464,N_26836,N_25546);
and U27465 (N_27465,N_24677,N_24919);
and U27466 (N_27466,N_26548,N_25239);
and U27467 (N_27467,N_24717,N_25441);
nand U27468 (N_27468,N_26606,N_25374);
and U27469 (N_27469,N_25622,N_26781);
nand U27470 (N_27470,N_25570,N_25535);
nor U27471 (N_27471,N_25825,N_25013);
or U27472 (N_27472,N_25798,N_26517);
or U27473 (N_27473,N_25605,N_24250);
nor U27474 (N_27474,N_26526,N_26997);
nor U27475 (N_27475,N_24543,N_24663);
and U27476 (N_27476,N_26495,N_24055);
nand U27477 (N_27477,N_26469,N_25858);
or U27478 (N_27478,N_25337,N_25001);
nand U27479 (N_27479,N_26969,N_25556);
nand U27480 (N_27480,N_24295,N_25099);
and U27481 (N_27481,N_26880,N_24043);
nor U27482 (N_27482,N_25166,N_25653);
or U27483 (N_27483,N_25665,N_26959);
or U27484 (N_27484,N_26744,N_24084);
nor U27485 (N_27485,N_26783,N_26547);
nor U27486 (N_27486,N_24828,N_24982);
nand U27487 (N_27487,N_26822,N_25443);
nor U27488 (N_27488,N_24006,N_24067);
or U27489 (N_27489,N_26750,N_25683);
nand U27490 (N_27490,N_25190,N_24529);
nand U27491 (N_27491,N_26509,N_26419);
nand U27492 (N_27492,N_25925,N_24406);
or U27493 (N_27493,N_25302,N_26879);
and U27494 (N_27494,N_25855,N_26389);
nor U27495 (N_27495,N_24349,N_25217);
nor U27496 (N_27496,N_24728,N_25652);
and U27497 (N_27497,N_25440,N_26349);
and U27498 (N_27498,N_24368,N_24167);
nand U27499 (N_27499,N_24013,N_24096);
and U27500 (N_27500,N_25121,N_26805);
nor U27501 (N_27501,N_24401,N_25483);
or U27502 (N_27502,N_24875,N_24393);
nand U27503 (N_27503,N_24587,N_26178);
nor U27504 (N_27504,N_25962,N_25531);
nor U27505 (N_27505,N_25484,N_24582);
and U27506 (N_27506,N_24296,N_24436);
or U27507 (N_27507,N_24090,N_25248);
nand U27508 (N_27508,N_25565,N_26839);
xor U27509 (N_27509,N_26973,N_25250);
xnor U27510 (N_27510,N_26569,N_26210);
nor U27511 (N_27511,N_26049,N_24612);
nor U27512 (N_27512,N_26811,N_24378);
or U27513 (N_27513,N_24835,N_24776);
nor U27514 (N_27514,N_24692,N_24178);
nor U27515 (N_27515,N_24583,N_25850);
or U27516 (N_27516,N_26940,N_24180);
nor U27517 (N_27517,N_24947,N_25271);
nor U27518 (N_27518,N_26309,N_25296);
xnor U27519 (N_27519,N_26109,N_25473);
nand U27520 (N_27520,N_26827,N_24386);
nand U27521 (N_27521,N_26244,N_26492);
nand U27522 (N_27522,N_26563,N_25841);
or U27523 (N_27523,N_25389,N_26124);
xnor U27524 (N_27524,N_25151,N_25935);
nand U27525 (N_27525,N_25444,N_24025);
nand U27526 (N_27526,N_24113,N_24225);
nand U27527 (N_27527,N_24763,N_25189);
or U27528 (N_27528,N_26463,N_25111);
or U27529 (N_27529,N_26661,N_26620);
xnor U27530 (N_27530,N_25548,N_24473);
nand U27531 (N_27531,N_24115,N_26410);
nor U27532 (N_27532,N_24410,N_25878);
xnor U27533 (N_27533,N_25301,N_26684);
nand U27534 (N_27534,N_24598,N_25408);
or U27535 (N_27535,N_25939,N_24485);
nor U27536 (N_27536,N_26411,N_24829);
nand U27537 (N_27537,N_26397,N_26978);
nor U27538 (N_27538,N_26314,N_24374);
nand U27539 (N_27539,N_24855,N_26775);
nor U27540 (N_27540,N_26954,N_26544);
nand U27541 (N_27541,N_24329,N_26685);
nor U27542 (N_27542,N_24789,N_24506);
or U27543 (N_27543,N_26009,N_25487);
nand U27544 (N_27544,N_24457,N_24342);
nand U27545 (N_27545,N_26097,N_24880);
nand U27546 (N_27546,N_24668,N_25781);
and U27547 (N_27547,N_24168,N_26594);
nand U27548 (N_27548,N_26864,N_25141);
and U27549 (N_27549,N_26474,N_25021);
nand U27550 (N_27550,N_24696,N_25963);
nand U27551 (N_27551,N_26278,N_26464);
nor U27552 (N_27552,N_25674,N_24256);
nand U27553 (N_27553,N_26704,N_24105);
and U27554 (N_27554,N_24122,N_25108);
or U27555 (N_27555,N_26889,N_24209);
nand U27556 (N_27556,N_26915,N_24367);
and U27557 (N_27557,N_24511,N_25918);
nor U27558 (N_27558,N_25365,N_26387);
nand U27559 (N_27559,N_25794,N_24585);
nand U27560 (N_27560,N_25955,N_24204);
or U27561 (N_27561,N_26179,N_24077);
and U27562 (N_27562,N_26907,N_24515);
and U27563 (N_27563,N_25334,N_26587);
nor U27564 (N_27564,N_24844,N_24490);
nand U27565 (N_27565,N_25537,N_24925);
or U27566 (N_27566,N_25094,N_25031);
nor U27567 (N_27567,N_25865,N_25147);
nand U27568 (N_27568,N_25451,N_26331);
xnor U27569 (N_27569,N_24052,N_25644);
xnor U27570 (N_27570,N_25227,N_26516);
nand U27571 (N_27571,N_24936,N_26350);
or U27572 (N_27572,N_25497,N_26491);
or U27573 (N_27573,N_24229,N_26385);
nor U27574 (N_27574,N_25554,N_26875);
nand U27575 (N_27575,N_25034,N_25284);
nor U27576 (N_27576,N_25461,N_26922);
or U27577 (N_27577,N_24086,N_25124);
or U27578 (N_27578,N_24913,N_24123);
and U27579 (N_27579,N_26375,N_26576);
nor U27580 (N_27580,N_26188,N_25859);
nor U27581 (N_27581,N_24963,N_24702);
or U27582 (N_27582,N_25820,N_25297);
or U27583 (N_27583,N_26214,N_24910);
nor U27584 (N_27584,N_25729,N_25843);
and U27585 (N_27585,N_24010,N_26341);
nor U27586 (N_27586,N_26566,N_25677);
nor U27587 (N_27587,N_24271,N_24389);
and U27588 (N_27588,N_25453,N_26807);
nand U27589 (N_27589,N_24930,N_25197);
xor U27590 (N_27590,N_24437,N_24089);
or U27591 (N_27591,N_26247,N_24227);
nand U27592 (N_27592,N_24022,N_24953);
and U27593 (N_27593,N_26168,N_26352);
and U27594 (N_27594,N_25646,N_26394);
nand U27595 (N_27595,N_26963,N_25567);
nand U27596 (N_27596,N_26982,N_26611);
or U27597 (N_27597,N_25106,N_26204);
nand U27598 (N_27598,N_24885,N_25053);
or U27599 (N_27599,N_26758,N_25763);
or U27600 (N_27600,N_24211,N_26012);
nor U27601 (N_27601,N_25688,N_24165);
and U27602 (N_27602,N_26723,N_24552);
or U27603 (N_27603,N_24427,N_26200);
nand U27604 (N_27604,N_26020,N_24815);
and U27605 (N_27605,N_24477,N_26591);
or U27606 (N_27606,N_26070,N_26794);
and U27607 (N_27607,N_25011,N_26308);
or U27608 (N_27608,N_26061,N_25267);
and U27609 (N_27609,N_24602,N_26660);
nor U27610 (N_27610,N_26831,N_24944);
xor U27611 (N_27611,N_24380,N_25079);
and U27612 (N_27612,N_24438,N_25624);
xor U27613 (N_27613,N_26776,N_24750);
nand U27614 (N_27614,N_25545,N_24434);
or U27615 (N_27615,N_24561,N_24435);
and U27616 (N_27616,N_26994,N_25654);
or U27617 (N_27617,N_25682,N_26943);
or U27618 (N_27618,N_26851,N_26307);
or U27619 (N_27619,N_26586,N_26030);
nor U27620 (N_27620,N_25854,N_26376);
and U27621 (N_27621,N_24361,N_25105);
nand U27622 (N_27622,N_26804,N_24989);
or U27623 (N_27623,N_25343,N_26598);
or U27624 (N_27624,N_26694,N_26164);
and U27625 (N_27625,N_26510,N_26334);
or U27626 (N_27626,N_25399,N_26245);
and U27627 (N_27627,N_25323,N_24474);
or U27628 (N_27628,N_24660,N_26296);
xnor U27629 (N_27629,N_25731,N_25977);
nand U27630 (N_27630,N_24986,N_24971);
nor U27631 (N_27631,N_24069,N_25701);
or U27632 (N_27632,N_24590,N_26052);
or U27633 (N_27633,N_25489,N_25308);
nor U27634 (N_27634,N_25626,N_24263);
nand U27635 (N_27635,N_26823,N_25260);
or U27636 (N_27636,N_26522,N_25571);
nand U27637 (N_27637,N_24027,N_26104);
and U27638 (N_27638,N_24802,N_24220);
nor U27639 (N_27639,N_25807,N_24399);
nand U27640 (N_27640,N_25756,N_24714);
or U27641 (N_27641,N_24744,N_25056);
nand U27642 (N_27642,N_24747,N_24002);
and U27643 (N_27643,N_26320,N_24352);
and U27644 (N_27644,N_26362,N_24362);
and U27645 (N_27645,N_25233,N_24629);
nand U27646 (N_27646,N_24780,N_24822);
and U27647 (N_27647,N_26144,N_24681);
nor U27648 (N_27648,N_24889,N_24287);
nor U27649 (N_27649,N_24658,N_25647);
nor U27650 (N_27650,N_25563,N_24896);
and U27651 (N_27651,N_26223,N_25164);
nor U27652 (N_27652,N_25494,N_25885);
nand U27653 (N_27653,N_24156,N_24112);
nand U27654 (N_27654,N_25294,N_25506);
nand U27655 (N_27655,N_26295,N_26686);
or U27656 (N_27656,N_26699,N_24871);
xor U27657 (N_27657,N_25937,N_24893);
xor U27658 (N_27658,N_24215,N_25732);
nand U27659 (N_27659,N_26069,N_24782);
nor U27660 (N_27660,N_25959,N_26824);
nand U27661 (N_27661,N_25237,N_25303);
nor U27662 (N_27662,N_25247,N_26405);
xnor U27663 (N_27663,N_26960,N_24076);
and U27664 (N_27664,N_24545,N_26542);
and U27665 (N_27665,N_25254,N_24973);
or U27666 (N_27666,N_25426,N_24432);
or U27667 (N_27667,N_26292,N_25216);
or U27668 (N_27668,N_25901,N_26767);
and U27669 (N_27669,N_26930,N_26032);
nor U27670 (N_27670,N_26306,N_24001);
nand U27671 (N_27671,N_26462,N_26277);
nor U27672 (N_27672,N_24949,N_26086);
nand U27673 (N_27673,N_26470,N_26519);
nor U27674 (N_27674,N_25319,N_24670);
nand U27675 (N_27675,N_26137,N_26190);
nand U27676 (N_27676,N_24255,N_26050);
nor U27677 (N_27677,N_26613,N_25936);
or U27678 (N_27678,N_24501,N_25985);
nand U27679 (N_27679,N_25377,N_24164);
nor U27680 (N_27680,N_24843,N_26736);
xnor U27681 (N_27681,N_26479,N_26121);
nand U27682 (N_27682,N_24307,N_26484);
nor U27683 (N_27683,N_25321,N_24737);
or U27684 (N_27684,N_25634,N_24426);
and U27685 (N_27685,N_24282,N_24645);
and U27686 (N_27686,N_25905,N_25564);
nor U27687 (N_27687,N_24915,N_24727);
and U27688 (N_27688,N_25876,N_25082);
nor U27689 (N_27689,N_25914,N_25714);
nor U27690 (N_27690,N_25964,N_26442);
nand U27691 (N_27691,N_26513,N_25456);
or U27692 (N_27692,N_26062,N_26253);
or U27693 (N_27693,N_26192,N_26382);
nor U27694 (N_27694,N_24994,N_25530);
xnor U27695 (N_27695,N_24767,N_24975);
nand U27696 (N_27696,N_24394,N_25508);
and U27697 (N_27697,N_24752,N_24274);
nand U27698 (N_27698,N_25817,N_24988);
nor U27699 (N_27699,N_26229,N_26756);
or U27700 (N_27700,N_25643,N_25552);
nand U27701 (N_27701,N_25615,N_24032);
nor U27702 (N_27702,N_26002,N_25668);
and U27703 (N_27703,N_25520,N_24955);
and U27704 (N_27704,N_24623,N_25007);
nand U27705 (N_27705,N_25252,N_26134);
or U27706 (N_27706,N_24553,N_24415);
and U27707 (N_27707,N_25050,N_26681);
and U27708 (N_27708,N_26934,N_24746);
nor U27709 (N_27709,N_26505,N_26336);
or U27710 (N_27710,N_25127,N_25950);
nor U27711 (N_27711,N_26914,N_25730);
or U27712 (N_27712,N_25397,N_26762);
nor U27713 (N_27713,N_25547,N_25603);
nor U27714 (N_27714,N_25191,N_25156);
and U27715 (N_27715,N_25971,N_24539);
nand U27716 (N_27716,N_26537,N_25355);
and U27717 (N_27717,N_25629,N_25719);
nand U27718 (N_27718,N_24011,N_26708);
and U27719 (N_27719,N_24526,N_26233);
or U27720 (N_27720,N_25984,N_24653);
and U27721 (N_27721,N_25112,N_24347);
and U27722 (N_27722,N_26196,N_25874);
or U27723 (N_27723,N_25351,N_24954);
and U27724 (N_27724,N_24749,N_25684);
nand U27725 (N_27725,N_24901,N_24818);
or U27726 (N_27726,N_24799,N_24995);
nand U27727 (N_27727,N_26099,N_26110);
nor U27728 (N_27728,N_24444,N_25960);
nand U27729 (N_27729,N_26644,N_25455);
nor U27730 (N_27730,N_24234,N_26379);
nand U27731 (N_27731,N_25948,N_24964);
and U27732 (N_27732,N_24563,N_26193);
nor U27733 (N_27733,N_24012,N_24121);
or U27734 (N_27734,N_25840,N_26841);
nand U27735 (N_27735,N_26933,N_24468);
and U27736 (N_27736,N_25332,N_26894);
or U27737 (N_27737,N_25084,N_26060);
and U27738 (N_27738,N_25808,N_25459);
nor U27739 (N_27739,N_24643,N_24433);
and U27740 (N_27740,N_25819,N_25543);
nor U27741 (N_27741,N_24524,N_26102);
nand U27742 (N_27742,N_24775,N_24456);
or U27743 (N_27743,N_26837,N_26357);
or U27744 (N_27744,N_24985,N_24860);
xnor U27745 (N_27745,N_24182,N_26260);
nor U27746 (N_27746,N_24761,N_25107);
and U27747 (N_27747,N_26655,N_26588);
xor U27748 (N_27748,N_26872,N_26631);
nand U27749 (N_27749,N_24128,N_25857);
or U27750 (N_27750,N_25068,N_24267);
and U27751 (N_27751,N_24316,N_25158);
nand U27752 (N_27752,N_26763,N_26090);
or U27753 (N_27753,N_24655,N_25033);
and U27754 (N_27754,N_24219,N_25433);
and U27755 (N_27755,N_26962,N_24928);
nor U27756 (N_27756,N_24031,N_26494);
xor U27757 (N_27757,N_24614,N_25619);
nand U27758 (N_27758,N_25213,N_26601);
nor U27759 (N_27759,N_25932,N_24608);
and U27760 (N_27760,N_25089,N_26226);
and U27761 (N_27761,N_26266,N_26865);
nand U27762 (N_27762,N_26691,N_24695);
nor U27763 (N_27763,N_24979,N_26712);
nand U27764 (N_27764,N_24509,N_26730);
nand U27765 (N_27765,N_26813,N_26581);
nor U27766 (N_27766,N_24308,N_24466);
and U27767 (N_27767,N_26869,N_26284);
nand U27768 (N_27768,N_26873,N_24200);
or U27769 (N_27769,N_25410,N_25980);
nor U27770 (N_27770,N_25169,N_26354);
nand U27771 (N_27771,N_24809,N_25000);
and U27772 (N_27772,N_25006,N_26374);
xnor U27773 (N_27773,N_24920,N_25586);
nand U27774 (N_27774,N_24232,N_25311);
and U27775 (N_27775,N_26742,N_25005);
nand U27776 (N_27776,N_26501,N_26508);
nand U27777 (N_27777,N_24850,N_24935);
or U27778 (N_27778,N_24571,N_26778);
and U27779 (N_27779,N_26000,N_25618);
nor U27780 (N_27780,N_26466,N_24907);
xnor U27781 (N_27781,N_25055,N_26111);
nand U27782 (N_27782,N_24772,N_24421);
nand U27783 (N_27783,N_24541,N_26001);
or U27784 (N_27784,N_26999,N_24774);
xnor U27785 (N_27785,N_24424,N_26011);
and U27786 (N_27786,N_24707,N_24987);
nand U27787 (N_27787,N_26222,N_25125);
and U27788 (N_27788,N_24745,N_25329);
nor U27789 (N_27789,N_25438,N_24119);
and U27790 (N_27790,N_24042,N_26833);
or U27791 (N_27791,N_26315,N_24652);
or U27792 (N_27792,N_24481,N_24592);
or U27793 (N_27793,N_25090,N_26619);
or U27794 (N_27794,N_25696,N_26656);
nor U27795 (N_27795,N_26975,N_24453);
or U27796 (N_27796,N_24877,N_24952);
and U27797 (N_27797,N_25883,N_26696);
nand U27798 (N_27798,N_24698,N_25232);
and U27799 (N_27799,N_24576,N_25743);
or U27800 (N_27800,N_24236,N_26992);
nand U27801 (N_27801,N_25672,N_26421);
nand U27802 (N_27802,N_26897,N_26858);
or U27803 (N_27803,N_25325,N_24705);
and U27804 (N_27804,N_25040,N_25988);
or U27805 (N_27805,N_26785,N_24116);
and U27806 (N_27806,N_25128,N_25210);
nor U27807 (N_27807,N_24721,N_25847);
xor U27808 (N_27808,N_24618,N_25054);
nor U27809 (N_27809,N_26452,N_26703);
and U27810 (N_27810,N_24547,N_25117);
xnor U27811 (N_27811,N_25309,N_25774);
and U27812 (N_27812,N_26711,N_25109);
and U27813 (N_27813,N_26161,N_25097);
or U27814 (N_27814,N_26175,N_24933);
and U27815 (N_27815,N_24588,N_26369);
nand U27816 (N_27816,N_24292,N_26347);
nor U27817 (N_27817,N_25353,N_24252);
nor U27818 (N_27818,N_24346,N_24638);
and U27819 (N_27819,N_24276,N_24254);
and U27820 (N_27820,N_26949,N_26749);
nand U27821 (N_27821,N_24044,N_26673);
xor U27822 (N_27822,N_24651,N_24817);
nand U27823 (N_27823,N_26122,N_26731);
nor U27824 (N_27824,N_24911,N_25071);
or U27825 (N_27825,N_26465,N_24120);
or U27826 (N_27826,N_26243,N_25532);
and U27827 (N_27827,N_26140,N_24412);
nor U27828 (N_27828,N_24498,N_26902);
nor U27829 (N_27829,N_26305,N_26662);
or U27830 (N_27830,N_25086,N_24441);
xor U27831 (N_27831,N_25698,N_26698);
nor U27832 (N_27832,N_26360,N_26171);
nand U27833 (N_27833,N_25211,N_26310);
and U27834 (N_27834,N_24315,N_26680);
nor U27835 (N_27835,N_25331,N_25954);
nor U27836 (N_27836,N_24785,N_26085);
nand U27837 (N_27837,N_26876,N_26636);
nor U27838 (N_27838,N_25462,N_24452);
nor U27839 (N_27839,N_24833,N_24080);
nand U27840 (N_27840,N_24603,N_26887);
nor U27841 (N_27841,N_25632,N_25768);
or U27842 (N_27842,N_24301,N_24187);
and U27843 (N_27843,N_26530,N_25305);
and U27844 (N_27844,N_25414,N_24162);
nor U27845 (N_27845,N_25973,N_24047);
nand U27846 (N_27846,N_26256,N_24408);
nor U27847 (N_27847,N_26610,N_24891);
nand U27848 (N_27848,N_25405,N_26340);
and U27849 (N_27849,N_24500,N_25986);
or U27850 (N_27850,N_24518,N_24057);
and U27851 (N_27851,N_24573,N_25346);
nor U27852 (N_27852,N_25568,N_26739);
and U27853 (N_27853,N_24273,N_26136);
and U27854 (N_27854,N_26422,N_26359);
or U27855 (N_27855,N_26891,N_24505);
nor U27856 (N_27856,N_25866,N_25134);
or U27857 (N_27857,N_25848,N_26272);
nand U27858 (N_27858,N_25384,N_26553);
and U27859 (N_27859,N_24851,N_26185);
nand U27860 (N_27860,N_24414,N_25244);
or U27861 (N_27861,N_24066,N_24619);
nand U27862 (N_27862,N_25347,N_26716);
and U27863 (N_27863,N_25739,N_24566);
and U27864 (N_27864,N_24673,N_24859);
xor U27865 (N_27865,N_25279,N_24694);
nand U27866 (N_27866,N_26646,N_25043);
or U27867 (N_27867,N_25209,N_24125);
and U27868 (N_27868,N_25735,N_24171);
xnor U27869 (N_27869,N_24836,N_25306);
nand U27870 (N_27870,N_26302,N_26667);
or U27871 (N_27871,N_26373,N_25268);
and U27872 (N_27872,N_26146,N_25091);
nand U27873 (N_27873,N_24070,N_25085);
and U27874 (N_27874,N_25789,N_24950);
and U27875 (N_27875,N_25861,N_25207);
nand U27876 (N_27876,N_26255,N_26105);
and U27877 (N_27877,N_24050,N_24353);
nor U27878 (N_27878,N_26868,N_24008);
xnor U27879 (N_27879,N_24486,N_24337);
nor U27880 (N_27880,N_24447,N_25142);
or U27881 (N_27881,N_25956,N_24416);
nor U27882 (N_27882,N_26450,N_25522);
and U27883 (N_27883,N_26326,N_25240);
nor U27884 (N_27884,N_26637,N_26687);
and U27885 (N_27885,N_25600,N_26058);
nor U27886 (N_27886,N_25777,N_26766);
nand U27887 (N_27887,N_24186,N_25065);
nor U27888 (N_27888,N_26458,N_26579);
nand U27889 (N_27889,N_26093,N_25981);
nor U27890 (N_27890,N_25748,N_24371);
nand U27891 (N_27891,N_26628,N_25912);
nand U27892 (N_27892,N_26800,N_24476);
nand U27893 (N_27893,N_24205,N_24993);
nand U27894 (N_27894,N_26057,N_26721);
and U27895 (N_27895,N_25339,N_24482);
or U27896 (N_27896,N_24098,N_25927);
or U27897 (N_27897,N_26600,N_26986);
or U27898 (N_27898,N_25516,N_26330);
and U27899 (N_27899,N_25242,N_25957);
xnor U27900 (N_27900,N_26116,N_25638);
nor U27901 (N_27901,N_26788,N_24446);
nand U27902 (N_27902,N_24578,N_24140);
nor U27903 (N_27903,N_26427,N_26215);
nor U27904 (N_27904,N_26951,N_25895);
xor U27905 (N_27905,N_25809,N_24832);
nand U27906 (N_27906,N_24831,N_24151);
nor U27907 (N_27907,N_25771,N_25472);
and U27908 (N_27908,N_24554,N_26657);
nand U27909 (N_27909,N_25396,N_24601);
nand U27910 (N_27910,N_24610,N_25995);
xnor U27911 (N_27911,N_25695,N_24422);
and U27912 (N_27912,N_24443,N_26203);
nor U27913 (N_27913,N_25420,N_24664);
nand U27914 (N_27914,N_24713,N_26037);
nand U27915 (N_27915,N_25246,N_25824);
or U27916 (N_27916,N_25131,N_24157);
nand U27917 (N_27917,N_25047,N_24905);
or U27918 (N_27918,N_25635,N_26230);
nor U27919 (N_27919,N_26449,N_26227);
nor U27920 (N_27920,N_24419,N_24771);
or U27921 (N_27921,N_24365,N_25692);
and U27922 (N_27922,N_24246,N_26525);
and U27923 (N_27923,N_25182,N_24134);
xor U27924 (N_27924,N_24146,N_26700);
nand U27925 (N_27925,N_25555,N_26771);
nand U27926 (N_27926,N_24723,N_25363);
nor U27927 (N_27927,N_25996,N_26356);
nand U27928 (N_27928,N_26892,N_25502);
nand U27929 (N_27929,N_26886,N_24689);
or U27930 (N_27930,N_25269,N_26570);
or U27931 (N_27931,N_25430,N_24334);
nand U27932 (N_27932,N_24063,N_25429);
nor U27933 (N_27933,N_26113,N_26160);
nor U27934 (N_27934,N_26665,N_24480);
xnor U27935 (N_27935,N_26920,N_25512);
xor U27936 (N_27936,N_25610,N_25818);
nor U27937 (N_27937,N_26276,N_25800);
nor U27938 (N_27938,N_24003,N_25581);
nor U27939 (N_27939,N_24758,N_24943);
xor U27940 (N_27940,N_24641,N_24088);
and U27941 (N_27941,N_26054,N_25314);
and U27942 (N_27942,N_24742,N_26197);
xnor U27943 (N_27943,N_26760,N_26514);
xnor U27944 (N_27944,N_24064,N_26481);
nor U27945 (N_27945,N_24228,N_25342);
nor U27946 (N_27946,N_24773,N_26301);
and U27947 (N_27947,N_25614,N_25092);
nor U27948 (N_27948,N_25049,N_25465);
or U27949 (N_27949,N_25274,N_26497);
and U27950 (N_27950,N_25257,N_24247);
or U27951 (N_27951,N_25286,N_24259);
nand U27952 (N_27952,N_26772,N_26433);
xnor U27953 (N_27953,N_26493,N_25762);
nand U27954 (N_27954,N_25432,N_25911);
xor U27955 (N_27955,N_26046,N_25145);
nand U27956 (N_27956,N_25662,N_24283);
or U27957 (N_27957,N_26274,N_26034);
nor U27958 (N_27958,N_25445,N_25697);
or U27959 (N_27959,N_25898,N_26759);
or U27960 (N_27960,N_26908,N_24275);
nor U27961 (N_27961,N_24559,N_25333);
or U27962 (N_27962,N_26490,N_24991);
nand U27963 (N_27963,N_24028,N_26676);
or U27964 (N_27964,N_24258,N_25710);
and U27965 (N_27965,N_25392,N_25471);
and U27966 (N_27966,N_26511,N_26251);
and U27967 (N_27967,N_24224,N_25413);
xor U27968 (N_27968,N_24350,N_24508);
and U27969 (N_27969,N_26149,N_26283);
or U27970 (N_27970,N_26770,N_25575);
or U27971 (N_27971,N_25680,N_26910);
and U27972 (N_27972,N_25057,N_25312);
nand U27973 (N_27973,N_24277,N_24922);
nand U27974 (N_27974,N_24837,N_24917);
or U27975 (N_27975,N_24599,N_26988);
or U27976 (N_27976,N_25372,N_25515);
and U27977 (N_27977,N_24087,N_24765);
or U27978 (N_27978,N_24665,N_25790);
and U27979 (N_27979,N_26151,N_24338);
nand U27980 (N_27980,N_26023,N_25069);
nand U27981 (N_27981,N_26089,N_24867);
nor U27982 (N_27982,N_24674,N_25495);
and U27983 (N_27983,N_24372,N_25952);
or U27984 (N_27984,N_24161,N_24600);
nor U27985 (N_27985,N_24715,N_26607);
xor U27986 (N_27986,N_26004,N_24513);
or U27987 (N_27987,N_26080,N_24007);
or U27988 (N_27988,N_24819,N_26638);
xnor U27989 (N_27989,N_25641,N_26572);
nand U27990 (N_27990,N_26556,N_26180);
xor U27991 (N_27991,N_25524,N_25283);
nand U27992 (N_27992,N_25037,N_26040);
nor U27993 (N_27993,N_24591,N_26506);
or U27994 (N_27994,N_25649,N_24525);
and U27995 (N_27995,N_26318,N_25499);
nor U27996 (N_27996,N_26755,N_26166);
and U27997 (N_27997,N_24992,N_24360);
and U27998 (N_27998,N_25320,N_24884);
nor U27999 (N_27999,N_26998,N_25997);
nand U28000 (N_28000,N_24314,N_25382);
nand U28001 (N_28001,N_26881,N_24607);
xnor U28002 (N_28002,N_24488,N_24286);
and U28003 (N_28003,N_25666,N_24628);
nand U28004 (N_28004,N_25903,N_24594);
xnor U28005 (N_28005,N_25805,N_26237);
nor U28006 (N_28006,N_25863,N_25913);
and U28007 (N_28007,N_24914,N_26453);
xnor U28008 (N_28008,N_24323,N_24173);
nor U28009 (N_28009,N_25587,N_25906);
nand U28010 (N_28010,N_25245,N_24183);
and U28011 (N_28011,N_26552,N_26896);
nand U28012 (N_28012,N_24023,N_24937);
nor U28013 (N_28013,N_25022,N_25434);
nand U28014 (N_28014,N_25023,N_24400);
nand U28015 (N_28015,N_26578,N_25965);
nor U28016 (N_28016,N_25709,N_24557);
or U28017 (N_28017,N_26849,N_26145);
and U28018 (N_28018,N_25892,N_25636);
nor U28019 (N_28019,N_24201,N_25120);
and U28020 (N_28020,N_25958,N_25132);
nor U28021 (N_28021,N_25700,N_24311);
nand U28022 (N_28022,N_26567,N_26983);
nand U28023 (N_28023,N_26087,N_26834);
nand U28024 (N_28024,N_25842,N_25073);
xnor U28025 (N_28025,N_26258,N_26447);
nand U28026 (N_28026,N_24095,N_24567);
or U28027 (N_28027,N_25711,N_25766);
and U28028 (N_28028,N_24420,N_26819);
nor U28029 (N_28029,N_25135,N_25723);
xnor U28030 (N_28030,N_25612,N_25076);
nand U28031 (N_28031,N_24065,N_26782);
or U28032 (N_28032,N_24208,N_26064);
nand U28033 (N_28033,N_26500,N_25153);
and U28034 (N_28034,N_24390,N_26293);
nor U28035 (N_28035,N_26467,N_26582);
nor U28036 (N_28036,N_26893,N_26939);
and U28037 (N_28037,N_25533,N_26126);
nor U28038 (N_28038,N_25078,N_24690);
or U28039 (N_28039,N_24770,N_25116);
nor U28040 (N_28040,N_24015,N_25015);
or U28041 (N_28041,N_24492,N_24464);
or U28042 (N_28042,N_24688,N_25281);
or U28043 (N_28043,N_25542,N_25951);
xnor U28044 (N_28044,N_25689,N_26754);
and U28045 (N_28045,N_26088,N_26640);
and U28046 (N_28046,N_25202,N_25492);
and U28047 (N_28047,N_25464,N_26187);
nor U28048 (N_28048,N_25474,N_24687);
and U28049 (N_28049,N_26201,N_24759);
xor U28050 (N_28050,N_24449,N_26769);
nand U28051 (N_28051,N_25802,N_25282);
xnor U28052 (N_28052,N_24704,N_25795);
nand U28053 (N_28053,N_25889,N_24106);
and U28054 (N_28054,N_26512,N_25226);
nor U28055 (N_28055,N_26005,N_25025);
or U28056 (N_28056,N_24272,N_24793);
or U28057 (N_28057,N_25870,N_26617);
and U28058 (N_28058,N_25831,N_25510);
nor U28059 (N_28059,N_26946,N_26459);
nand U28060 (N_28060,N_25029,N_26457);
and U28061 (N_28061,N_26446,N_26015);
and U28062 (N_28062,N_24404,N_24510);
nor U28063 (N_28063,N_24527,N_25721);
and U28064 (N_28064,N_25272,N_25782);
nor U28065 (N_28065,N_24853,N_26918);
nand U28066 (N_28066,N_26882,N_26358);
nand U28067 (N_28067,N_26981,N_26312);
nand U28068 (N_28068,N_24489,N_26532);
and U28069 (N_28069,N_24431,N_26701);
nand U28070 (N_28070,N_26021,N_26198);
or U28071 (N_28071,N_26371,N_26130);
or U28072 (N_28072,N_26734,N_25667);
nor U28073 (N_28073,N_25755,N_25395);
nand U28074 (N_28074,N_25077,N_24319);
or U28075 (N_28075,N_26096,N_24609);
nor U28076 (N_28076,N_25616,N_26199);
xor U28077 (N_28077,N_26420,N_26663);
nor U28078 (N_28078,N_25750,N_26035);
nand U28079 (N_28079,N_26838,N_25884);
xnor U28080 (N_28080,N_25514,N_24417);
nand U28081 (N_28081,N_25846,N_25909);
xor U28082 (N_28082,N_24268,N_26445);
or U28083 (N_28083,N_26748,N_26735);
nand U28084 (N_28084,N_24269,N_25411);
or U28085 (N_28085,N_25724,N_24345);
nor U28086 (N_28086,N_25737,N_26333);
nand U28087 (N_28087,N_26036,N_24927);
nor U28088 (N_28088,N_24391,N_24109);
nand U28089 (N_28089,N_26488,N_26534);
or U28090 (N_28090,N_25797,N_24748);
nand U28091 (N_28091,N_26521,N_24642);
and U28092 (N_28092,N_26429,N_26078);
nand U28093 (N_28093,N_24625,N_25691);
or U28094 (N_28094,N_26845,N_26906);
xor U28095 (N_28095,N_25979,N_24912);
nor U28096 (N_28096,N_25221,N_24056);
xnor U28097 (N_28097,N_26612,N_25129);
and U28098 (N_28098,N_26871,N_25713);
nand U28099 (N_28099,N_25390,N_24033);
and U28100 (N_28100,N_24195,N_26353);
nor U28101 (N_28101,N_25424,N_24788);
or U28102 (N_28102,N_24046,N_24214);
nand U28103 (N_28103,N_26221,N_26163);
xor U28104 (N_28104,N_26112,N_26802);
xor U28105 (N_28105,N_24163,N_25072);
nor U28106 (N_28106,N_25149,N_25477);
nor U28107 (N_28107,N_26679,N_26118);
and U28108 (N_28108,N_24685,N_24838);
nand U28109 (N_28109,N_26844,N_24470);
nand U28110 (N_28110,N_24235,N_25639);
or U28111 (N_28111,N_25671,N_24932);
nand U28112 (N_28112,N_26697,N_26503);
and U28113 (N_28113,N_25369,N_25998);
nor U28114 (N_28114,N_24144,N_25562);
nand U28115 (N_28115,N_26828,N_25428);
nor U28116 (N_28116,N_24523,N_24978);
or U28117 (N_28117,N_25367,N_25673);
and U28118 (N_28118,N_25844,N_26987);
and U28119 (N_28119,N_25693,N_26972);
nor U28120 (N_28120,N_26418,N_25536);
or U28121 (N_28121,N_24313,N_25664);
nand U28122 (N_28122,N_26900,N_26861);
or U28123 (N_28123,N_25458,N_26659);
nor U28124 (N_28124,N_24395,N_26066);
and U28125 (N_28125,N_25277,N_26476);
or U28126 (N_28126,N_24137,N_24454);
nand U28127 (N_28127,N_26966,N_24324);
or U28128 (N_28128,N_25138,N_26890);
and U28129 (N_28129,N_25690,N_24662);
nand U28130 (N_28130,N_25648,N_24382);
nand U28131 (N_28131,N_25407,N_25550);
nand U28132 (N_28132,N_24310,N_25625);
nor U28133 (N_28133,N_25679,N_24848);
and U28134 (N_28134,N_24741,N_24126);
and U28135 (N_28135,N_24675,N_24593);
and U28136 (N_28136,N_24569,N_26098);
and U28137 (N_28137,N_26355,N_26451);
nor U28138 (N_28138,N_24560,N_24661);
xor U28139 (N_28139,N_25404,N_25500);
xor U28140 (N_28140,N_24093,N_25422);
and U28141 (N_28141,N_24265,N_26901);
nor U28142 (N_28142,N_25088,N_25733);
or U28143 (N_28143,N_24820,N_24876);
or U28144 (N_28144,N_25722,N_26174);
and U28145 (N_28145,N_24430,N_24621);
nand U28146 (N_28146,N_26670,N_25330);
and U28147 (N_28147,N_24169,N_25642);
nor U28148 (N_28148,N_24206,N_24029);
and U28149 (N_28149,N_24079,N_25637);
and U28150 (N_28150,N_25896,N_25967);
nand U28151 (N_28151,N_25480,N_24192);
nand U28152 (N_28152,N_26460,N_24676);
xor U28153 (N_28153,N_25860,N_24580);
xnor U28154 (N_28154,N_25378,N_25993);
nand U28155 (N_28155,N_26348,N_24483);
xor U28156 (N_28156,N_25008,N_24882);
xor U28157 (N_28157,N_24230,N_26007);
nor U28158 (N_28158,N_26809,N_26597);
nor U28159 (N_28159,N_26608,N_25200);
nor U28160 (N_28160,N_26456,N_26440);
and U28161 (N_28161,N_25776,N_26862);
and U28162 (N_28162,N_24941,N_26181);
and U28163 (N_28163,N_25140,N_26220);
nand U28164 (N_28164,N_24719,N_24327);
nor U28165 (N_28165,N_24810,N_26489);
nand U28166 (N_28166,N_24787,N_26028);
nand U28167 (N_28167,N_26068,N_26622);
and U28168 (N_28168,N_24407,N_25504);
nor U28169 (N_28169,N_25989,N_25969);
nand U28170 (N_28170,N_24188,N_25836);
nor U28171 (N_28171,N_24429,N_24730);
nor U28172 (N_28172,N_25273,N_24369);
or U28173 (N_28173,N_25907,N_26810);
and U28174 (N_28174,N_26262,N_26409);
nand U28175 (N_28175,N_24351,N_26172);
nor U28176 (N_28176,N_24462,N_26133);
nand U28177 (N_28177,N_25046,N_26249);
nand U28178 (N_28178,N_26970,N_25045);
and U28179 (N_28179,N_26444,N_26883);
or U28180 (N_28180,N_26815,N_25926);
nor U28181 (N_28181,N_25154,N_25058);
or U28182 (N_28182,N_26073,N_25559);
nor U28183 (N_28183,N_25394,N_26808);
or U28184 (N_28184,N_26135,N_24475);
or U28185 (N_28185,N_24199,N_26304);
nor U28186 (N_28186,N_26400,N_24708);
or U28187 (N_28187,N_26921,N_26321);
and U28188 (N_28188,N_24233,N_25943);
xor U28189 (N_28189,N_26019,N_25645);
and U28190 (N_28190,N_24862,N_24176);
and U28191 (N_28191,N_24703,N_26322);
nor U28192 (N_28192,N_25592,N_26536);
and U28193 (N_28193,N_24092,N_25617);
nand U28194 (N_28194,N_26045,N_24448);
or U28195 (N_28195,N_24402,N_26504);
or U28196 (N_28196,N_24262,N_24635);
xnor U28197 (N_28197,N_26472,N_24366);
or U28198 (N_28198,N_25338,N_24100);
or U28199 (N_28199,N_26977,N_25596);
nand U28200 (N_28200,N_24045,N_26706);
nand U28201 (N_28201,N_24179,N_26747);
and U28202 (N_28202,N_24409,N_24969);
or U28203 (N_28203,N_26346,N_24631);
or U28204 (N_28204,N_26319,N_26856);
and U28205 (N_28205,N_24644,N_25336);
and U28206 (N_28206,N_24237,N_25604);
and U28207 (N_28207,N_25591,N_25352);
or U28208 (N_28208,N_26329,N_24150);
nor U28209 (N_28209,N_26641,N_25044);
or U28210 (N_28210,N_25990,N_24769);
or U28211 (N_28211,N_26984,N_24926);
nor U28212 (N_28212,N_24996,N_26025);
nand U28213 (N_28213,N_24731,N_26041);
nand U28214 (N_28214,N_26094,N_26129);
nand U28215 (N_28215,N_25194,N_25439);
nor U28216 (N_28216,N_25699,N_24700);
nor U28217 (N_28217,N_25961,N_25813);
nor U28218 (N_28218,N_25655,N_25972);
and U28219 (N_28219,N_25923,N_25387);
xnor U28220 (N_28220,N_24736,N_24356);
and U28221 (N_28221,N_26543,N_26398);
nand U28222 (N_28222,N_25324,N_24738);
nor U28223 (N_28223,N_24132,N_26562);
or U28224 (N_28224,N_24579,N_25716);
nor U28225 (N_28225,N_26938,N_26590);
or U28226 (N_28226,N_24795,N_25380);
nand U28227 (N_28227,N_25110,N_26107);
and U28228 (N_28228,N_26888,N_24191);
nor U28229 (N_28229,N_25360,N_26927);
and U28230 (N_28230,N_25335,N_25137);
and U28231 (N_28231,N_24939,N_25235);
or U28232 (N_28232,N_26343,N_26793);
nand U28233 (N_28233,N_24534,N_25375);
nand U28234 (N_28234,N_26132,N_24540);
nand U28235 (N_28235,N_24455,N_24189);
xor U28236 (N_28236,N_25810,N_26014);
and U28237 (N_28237,N_24792,N_25315);
nand U28238 (N_28238,N_26439,N_25293);
or U28239 (N_28239,N_26741,N_26895);
nand U28240 (N_28240,N_26605,N_26857);
and U28241 (N_28241,N_25758,N_24484);
and U28242 (N_28242,N_26955,N_25573);
nor U28243 (N_28243,N_26206,N_24385);
nor U28244 (N_28244,N_24755,N_26008);
nor U28245 (N_28245,N_26859,N_24376);
and U28246 (N_28246,N_25970,N_24124);
nor U28247 (N_28247,N_26079,N_25594);
and U28248 (N_28248,N_24141,N_24842);
or U28249 (N_28249,N_26688,N_26625);
and U28250 (N_28250,N_24364,N_26372);
and U28251 (N_28251,N_24751,N_25947);
nor U28252 (N_28252,N_25928,N_26300);
nand U28253 (N_28253,N_25753,N_24626);
and U28254 (N_28254,N_24671,N_24678);
and U28255 (N_28255,N_24359,N_24699);
or U28256 (N_28256,N_26038,N_24942);
nand U28257 (N_28257,N_24627,N_25728);
nand U28258 (N_28258,N_25167,N_25416);
nand U28259 (N_28259,N_24981,N_26246);
nor U28260 (N_28260,N_24014,N_26218);
nor U28261 (N_28261,N_25886,N_24800);
nand U28262 (N_28262,N_25223,N_25705);
nor U28263 (N_28263,N_25159,N_26261);
nand U28264 (N_28264,N_24094,N_25675);
xor U28265 (N_28265,N_24502,N_26082);
and U28266 (N_28266,N_25185,N_26426);
nand U28267 (N_28267,N_25113,N_26402);
xor U28268 (N_28268,N_24639,N_24312);
nor U28269 (N_28269,N_24344,N_25706);
nor U28270 (N_28270,N_26814,N_24701);
or U28271 (N_28271,N_24507,N_25879);
nand U28272 (N_28272,N_24075,N_25754);
nor U28273 (N_28273,N_25383,N_26208);
nor U28274 (N_28274,N_26669,N_26281);
nand U28275 (N_28275,N_25402,N_26674);
and U28276 (N_28276,N_24294,N_24724);
or U28277 (N_28277,N_25894,N_26294);
or U28278 (N_28278,N_26695,N_24754);
and U28279 (N_28279,N_26950,N_25364);
and U28280 (N_28280,N_26119,N_24683);
xor U28281 (N_28281,N_26996,N_25804);
and U28282 (N_28282,N_24266,N_26675);
or U28283 (N_28283,N_26787,N_25103);
or U28284 (N_28284,N_25133,N_24082);
nor U28285 (N_28285,N_26432,N_26633);
or U28286 (N_28286,N_25788,N_25796);
nand U28287 (N_28287,N_26499,N_24906);
or U28288 (N_28288,N_25030,N_26393);
or U28289 (N_28289,N_26238,N_25348);
or U28290 (N_28290,N_25035,N_24333);
nor U28291 (N_28291,N_25298,N_24019);
or U28292 (N_28292,N_26777,N_24918);
nand U28293 (N_28293,N_24133,N_25206);
or U28294 (N_28294,N_24791,N_24589);
xor U28295 (N_28295,N_26609,N_24965);
and U28296 (N_28296,N_25511,N_24984);
nand U28297 (N_28297,N_24305,N_25060);
and U28298 (N_28298,N_25578,N_26722);
or U28299 (N_28299,N_25457,N_25258);
nor U28300 (N_28300,N_26595,N_25488);
nor U28301 (N_28301,N_24104,N_24051);
nor U28302 (N_28302,N_26033,N_26441);
nor U28303 (N_28303,N_25251,N_24807);
and U28304 (N_28304,N_25032,N_26965);
and U28305 (N_28305,N_25551,N_24841);
and U28306 (N_28306,N_26264,N_26961);
nor U28307 (N_28307,N_26653,N_26388);
nor U28308 (N_28308,N_24135,N_25966);
nor U28309 (N_28309,N_25707,N_26202);
or U28310 (N_28310,N_26990,N_25627);
and U28311 (N_28311,N_26313,N_25224);
and U28312 (N_28312,N_25585,N_25598);
nand U28313 (N_28313,N_26031,N_26381);
nand U28314 (N_28314,N_26714,N_24040);
or U28315 (N_28315,N_25064,N_25752);
nand U28316 (N_28316,N_26339,N_26242);
and U28317 (N_28317,N_25663,N_24026);
nor U28318 (N_28318,N_24549,N_24336);
or U28319 (N_28319,N_25864,N_24302);
and U28320 (N_28320,N_24306,N_24517);
nor U28321 (N_28321,N_26091,N_25561);
nor U28322 (N_28322,N_26454,N_26228);
or U28323 (N_28323,N_25920,N_25393);
and U28324 (N_28324,N_26332,N_25613);
xnor U28325 (N_28325,N_25908,N_24081);
nor U28326 (N_28326,N_25803,N_24243);
nand U28327 (N_28327,N_26399,N_26652);
and U28328 (N_28328,N_25236,N_26337);
nand U28329 (N_28329,N_24253,N_24522);
or U28330 (N_28330,N_24062,N_25746);
or U28331 (N_28331,N_24216,N_26391);
or U28332 (N_28332,N_24990,N_26380);
and U28333 (N_28333,N_25061,N_25468);
or U28334 (N_28334,N_26757,N_25238);
or U28335 (N_28335,N_25868,N_26786);
and U28336 (N_28336,N_25897,N_24551);
nor U28337 (N_28337,N_26430,N_24257);
nor U28338 (N_28338,N_25640,N_24478);
and U28339 (N_28339,N_25945,N_25881);
xor U28340 (N_28340,N_24883,N_26672);
or U28341 (N_28341,N_26084,N_26898);
nand U28342 (N_28342,N_26533,N_24240);
nand U28343 (N_28343,N_25219,N_25143);
and U28344 (N_28344,N_26658,N_25243);
or U28345 (N_28345,N_24320,N_26528);
and U28346 (N_28346,N_25215,N_26127);
nor U28347 (N_28347,N_26074,N_26115);
or U28348 (N_28348,N_26056,N_24129);
and U28349 (N_28349,N_26103,N_26365);
xor U28350 (N_28350,N_25976,N_26290);
nor U28351 (N_28351,N_24078,N_24805);
and U28352 (N_28352,N_24756,N_25576);
and U28353 (N_28353,N_24024,N_24403);
xnor U28354 (N_28354,N_25123,N_25900);
nor U28355 (N_28355,N_26535,N_26852);
or U28356 (N_28356,N_24185,N_25608);
nand U28357 (N_28357,N_25431,N_25949);
or U28358 (N_28358,N_24060,N_24537);
nor U28359 (N_28359,N_26705,N_26671);
xor U28360 (N_28360,N_24278,N_26855);
or U28361 (N_28361,N_26173,N_25658);
nor U28362 (N_28362,N_25708,N_26689);
nor U28363 (N_28363,N_26724,N_26142);
and U28364 (N_28364,N_24568,N_25098);
nand U28365 (N_28365,N_26585,N_25063);
xnor U28366 (N_28366,N_25799,N_24854);
nand U28367 (N_28367,N_26147,N_25922);
nand U28368 (N_28368,N_25910,N_24813);
xnor U28369 (N_28369,N_25316,N_26931);
and U28370 (N_28370,N_24461,N_25523);
or U28371 (N_28371,N_24546,N_24904);
and U28372 (N_28372,N_26668,N_24198);
nand U28373 (N_28373,N_25177,N_24512);
nand U28374 (N_28374,N_26903,N_26443);
nand U28375 (N_28375,N_26396,N_26779);
and U28376 (N_28376,N_26799,N_25317);
nand U28377 (N_28377,N_26832,N_25611);
or U28378 (N_28378,N_26342,N_26209);
or U28379 (N_28379,N_25230,N_24221);
and U28380 (N_28380,N_25574,N_25080);
and U28381 (N_28381,N_24538,N_24857);
or U28382 (N_28382,N_25657,N_24762);
nor U28383 (N_28383,N_26993,N_25725);
nand U28384 (N_28384,N_24520,N_24054);
nand U28385 (N_28385,N_26273,N_24881);
and U28386 (N_28386,N_26765,N_26874);
xnor U28387 (N_28387,N_24184,N_25678);
nor U28388 (N_28388,N_25228,N_24596);
nor U28389 (N_28389,N_26415,N_26645);
or U28390 (N_28390,N_26311,N_26271);
nand U28391 (N_28391,N_26796,N_26081);
nor U28392 (N_28392,N_26437,N_24487);
nand U28393 (N_28393,N_25225,N_26280);
and U28394 (N_28394,N_25285,N_26764);
or U28395 (N_28395,N_25507,N_26639);
nand U28396 (N_28396,N_24038,N_26071);
or U28397 (N_28397,N_26043,N_25100);
nor U28398 (N_28398,N_26557,N_24796);
xor U28399 (N_28399,N_26592,N_24099);
and U28400 (N_28400,N_24297,N_25102);
or U28401 (N_28401,N_26917,N_24899);
nor U28402 (N_28402,N_26139,N_26615);
nor U28403 (N_28403,N_26287,N_25028);
or U28404 (N_28404,N_26170,N_24202);
nand U28405 (N_28405,N_26577,N_25832);
and U28406 (N_28406,N_25929,N_26325);
nor U28407 (N_28407,N_24148,N_24999);
and U28408 (N_28408,N_24304,N_25205);
nor U28409 (N_28409,N_25493,N_25791);
nand U28410 (N_28410,N_26250,N_25994);
or U28411 (N_28411,N_24298,N_25620);
or U28412 (N_28412,N_25720,N_24550);
and U28413 (N_28413,N_26207,N_25358);
or U28414 (N_28414,N_24970,N_25987);
nand U28415 (N_28415,N_24030,N_24160);
and U28416 (N_28416,N_24528,N_25829);
and U28417 (N_28417,N_24245,N_26599);
nor U28418 (N_28418,N_25849,N_26167);
nor U28419 (N_28419,N_25310,N_25155);
nand U28420 (N_28420,N_25519,N_24617);
nand U28421 (N_28421,N_26216,N_25580);
nor U28422 (N_28422,N_26502,N_25902);
or U28423 (N_28423,N_24966,N_26471);
or U28424 (N_28424,N_24846,N_26790);
nand U28425 (N_28425,N_26478,N_24847);
and U28426 (N_28426,N_24281,N_26650);
or U28427 (N_28427,N_25882,N_25051);
nand U28428 (N_28428,N_25553,N_24957);
or U28429 (N_28429,N_24998,N_24249);
or U28430 (N_28430,N_24622,N_26546);
or U28431 (N_28431,N_24734,N_24898);
or U28432 (N_28432,N_26257,N_25814);
or U28433 (N_28433,N_26377,N_25162);
nand U28434 (N_28434,N_24869,N_26125);
or U28435 (N_28435,N_24803,N_25417);
or U28436 (N_28436,N_25871,N_24924);
nand U28437 (N_28437,N_25403,N_26932);
or U28438 (N_28438,N_26752,N_25165);
nor U28439 (N_28439,N_25180,N_26408);
nor U28440 (N_28440,N_26666,N_25083);
or U28441 (N_28441,N_25828,N_25930);
nor U28442 (N_28442,N_26270,N_26335);
nand U28443 (N_28443,N_25172,N_26138);
xnor U28444 (N_28444,N_26042,N_25919);
and U28445 (N_28445,N_25778,N_25066);
nor U28446 (N_28446,N_25203,N_24493);
nor U28447 (N_28447,N_26117,N_26259);
nand U28448 (N_28448,N_26473,N_26436);
or U28449 (N_28449,N_26252,N_24405);
and U28450 (N_28450,N_26435,N_24691);
nand U28451 (N_28451,N_26114,N_24101);
or U28452 (N_28452,N_26604,N_26912);
and U28453 (N_28453,N_24798,N_26475);
or U28454 (N_28454,N_26630,N_25359);
and U28455 (N_28455,N_26438,N_24640);
and U28456 (N_28456,N_26487,N_26518);
and U28457 (N_28457,N_25685,N_26128);
nand U28458 (N_28458,N_26616,N_25101);
and U28459 (N_28459,N_25096,N_26549);
nand U28460 (N_28460,N_25880,N_26801);
and U28461 (N_28461,N_24450,N_25139);
nor U28462 (N_28462,N_25623,N_26154);
or U28463 (N_28463,N_24616,N_25048);
xor U28464 (N_28464,N_24760,N_25446);
nand U28465 (N_28465,N_25195,N_24264);
nor U28466 (N_28466,N_24646,N_24777);
nor U28467 (N_28467,N_25830,N_26713);
xor U28468 (N_28468,N_25633,N_24948);
nand U28469 (N_28469,N_26141,N_24223);
nand U28470 (N_28470,N_24495,N_24697);
and U28471 (N_28471,N_26059,N_24564);
nand U28472 (N_28472,N_26044,N_24103);
nor U28473 (N_28473,N_25944,N_26212);
nand U28474 (N_28474,N_25893,N_26006);
nand U28475 (N_28475,N_26120,N_24916);
or U28476 (N_28476,N_24379,N_26541);
nand U28477 (N_28477,N_26194,N_24824);
and U28478 (N_28478,N_24572,N_26219);
nor U28479 (N_28479,N_26738,N_24348);
nor U28480 (N_28480,N_26143,N_25933);
nand U28481 (N_28481,N_24536,N_25270);
and U28482 (N_28482,N_26428,N_24647);
nor U28483 (N_28483,N_25942,N_24888);
and U28484 (N_28484,N_26583,N_25122);
nand U28485 (N_28485,N_24039,N_24620);
xor U28486 (N_28486,N_24840,N_24960);
or U28487 (N_28487,N_25425,N_24020);
or U28488 (N_28488,N_25196,N_24317);
nand U28489 (N_28489,N_24659,N_25288);
and U28490 (N_28490,N_26789,N_25448);
or U28491 (N_28491,N_26953,N_26267);
xor U28492 (N_28492,N_25198,N_25770);
or U28493 (N_28493,N_24597,N_26550);
and U28494 (N_28494,N_25601,N_25772);
and U28495 (N_28495,N_25742,N_25327);
nand U28496 (N_28496,N_26913,N_25144);
nand U28497 (N_28497,N_26540,N_25178);
or U28498 (N_28498,N_25787,N_25727);
and U28499 (N_28499,N_24816,N_26010);
and U28500 (N_28500,N_26037,N_24152);
nand U28501 (N_28501,N_24809,N_26083);
or U28502 (N_28502,N_26841,N_24544);
or U28503 (N_28503,N_24220,N_26329);
nand U28504 (N_28504,N_26363,N_24884);
nor U28505 (N_28505,N_24287,N_26498);
nand U28506 (N_28506,N_26157,N_24261);
and U28507 (N_28507,N_26776,N_24147);
nor U28508 (N_28508,N_24700,N_26974);
xor U28509 (N_28509,N_24856,N_25664);
nand U28510 (N_28510,N_24841,N_24689);
nor U28511 (N_28511,N_25692,N_24519);
nor U28512 (N_28512,N_26250,N_24787);
nor U28513 (N_28513,N_24491,N_24672);
or U28514 (N_28514,N_24036,N_25148);
nand U28515 (N_28515,N_24563,N_26915);
or U28516 (N_28516,N_24151,N_26821);
or U28517 (N_28517,N_25357,N_25211);
and U28518 (N_28518,N_26618,N_24449);
nand U28519 (N_28519,N_25226,N_24337);
nor U28520 (N_28520,N_25729,N_26551);
xor U28521 (N_28521,N_26214,N_25984);
or U28522 (N_28522,N_25987,N_24684);
nor U28523 (N_28523,N_25066,N_26708);
or U28524 (N_28524,N_25082,N_25972);
nand U28525 (N_28525,N_24278,N_26470);
nand U28526 (N_28526,N_26440,N_24191);
nand U28527 (N_28527,N_25619,N_25575);
nand U28528 (N_28528,N_24139,N_24935);
nand U28529 (N_28529,N_24468,N_25304);
nor U28530 (N_28530,N_24382,N_26514);
and U28531 (N_28531,N_24632,N_26067);
or U28532 (N_28532,N_24428,N_25733);
nand U28533 (N_28533,N_25319,N_25199);
and U28534 (N_28534,N_24171,N_24872);
and U28535 (N_28535,N_24516,N_25531);
nand U28536 (N_28536,N_24928,N_25804);
and U28537 (N_28537,N_26842,N_25728);
xnor U28538 (N_28538,N_24815,N_25413);
xnor U28539 (N_28539,N_26397,N_25928);
nor U28540 (N_28540,N_26683,N_24881);
nand U28541 (N_28541,N_24043,N_26258);
xor U28542 (N_28542,N_24670,N_26616);
or U28543 (N_28543,N_26794,N_24981);
nor U28544 (N_28544,N_25409,N_26337);
and U28545 (N_28545,N_25377,N_24115);
nand U28546 (N_28546,N_24407,N_25966);
and U28547 (N_28547,N_26307,N_24050);
or U28548 (N_28548,N_25965,N_26509);
nor U28549 (N_28549,N_25996,N_24653);
xnor U28550 (N_28550,N_26584,N_26469);
xor U28551 (N_28551,N_26908,N_26705);
or U28552 (N_28552,N_26095,N_26085);
nand U28553 (N_28553,N_24976,N_26603);
nor U28554 (N_28554,N_25477,N_24114);
nor U28555 (N_28555,N_26259,N_24156);
nand U28556 (N_28556,N_24193,N_25032);
xor U28557 (N_28557,N_26320,N_25964);
nor U28558 (N_28558,N_24719,N_26904);
or U28559 (N_28559,N_25392,N_26666);
or U28560 (N_28560,N_25037,N_26864);
nor U28561 (N_28561,N_25455,N_25949);
and U28562 (N_28562,N_24542,N_25362);
nor U28563 (N_28563,N_26661,N_26104);
nand U28564 (N_28564,N_26128,N_26141);
and U28565 (N_28565,N_26140,N_26652);
nor U28566 (N_28566,N_26841,N_26199);
nand U28567 (N_28567,N_24679,N_25786);
or U28568 (N_28568,N_24517,N_25376);
or U28569 (N_28569,N_24562,N_26024);
or U28570 (N_28570,N_25042,N_25383);
nand U28571 (N_28571,N_25052,N_25384);
nor U28572 (N_28572,N_24047,N_26321);
nand U28573 (N_28573,N_24680,N_25535);
or U28574 (N_28574,N_26105,N_25324);
nor U28575 (N_28575,N_24869,N_26898);
and U28576 (N_28576,N_26511,N_26654);
xor U28577 (N_28577,N_25756,N_25818);
xnor U28578 (N_28578,N_25893,N_24404);
nor U28579 (N_28579,N_25195,N_24120);
and U28580 (N_28580,N_24548,N_25038);
and U28581 (N_28581,N_25741,N_26925);
or U28582 (N_28582,N_25388,N_26311);
or U28583 (N_28583,N_24475,N_25429);
nor U28584 (N_28584,N_25740,N_26676);
and U28585 (N_28585,N_26615,N_24145);
nand U28586 (N_28586,N_26581,N_26218);
nor U28587 (N_28587,N_26850,N_26635);
nand U28588 (N_28588,N_25457,N_25892);
and U28589 (N_28589,N_24142,N_24428);
or U28590 (N_28590,N_24815,N_26403);
and U28591 (N_28591,N_26612,N_26644);
nand U28592 (N_28592,N_25579,N_24588);
nor U28593 (N_28593,N_26546,N_26816);
or U28594 (N_28594,N_25838,N_24350);
nor U28595 (N_28595,N_26131,N_24955);
nor U28596 (N_28596,N_25492,N_25188);
nand U28597 (N_28597,N_25681,N_24354);
and U28598 (N_28598,N_25020,N_25248);
nor U28599 (N_28599,N_25062,N_25288);
xor U28600 (N_28600,N_26259,N_26082);
nand U28601 (N_28601,N_26871,N_24216);
or U28602 (N_28602,N_26124,N_26664);
nor U28603 (N_28603,N_24007,N_26394);
or U28604 (N_28604,N_24722,N_25078);
nand U28605 (N_28605,N_25375,N_24325);
nor U28606 (N_28606,N_24858,N_25166);
and U28607 (N_28607,N_24106,N_26960);
nand U28608 (N_28608,N_24231,N_25460);
and U28609 (N_28609,N_24347,N_24050);
nand U28610 (N_28610,N_25072,N_24138);
or U28611 (N_28611,N_26267,N_24099);
nor U28612 (N_28612,N_25713,N_26085);
or U28613 (N_28613,N_26635,N_25921);
and U28614 (N_28614,N_24731,N_26028);
and U28615 (N_28615,N_24580,N_26799);
nand U28616 (N_28616,N_26719,N_24863);
and U28617 (N_28617,N_25370,N_24946);
nand U28618 (N_28618,N_24452,N_25199);
nand U28619 (N_28619,N_26741,N_26712);
nand U28620 (N_28620,N_25977,N_24846);
nand U28621 (N_28621,N_25423,N_24201);
nand U28622 (N_28622,N_24619,N_24929);
nand U28623 (N_28623,N_25753,N_26734);
nor U28624 (N_28624,N_24052,N_26639);
or U28625 (N_28625,N_24444,N_25988);
xor U28626 (N_28626,N_26971,N_26433);
nor U28627 (N_28627,N_25437,N_25921);
nor U28628 (N_28628,N_26214,N_25743);
nand U28629 (N_28629,N_25814,N_25655);
or U28630 (N_28630,N_26400,N_24264);
and U28631 (N_28631,N_25532,N_24463);
or U28632 (N_28632,N_25189,N_26713);
or U28633 (N_28633,N_24718,N_24904);
and U28634 (N_28634,N_26425,N_25902);
xnor U28635 (N_28635,N_25858,N_24445);
and U28636 (N_28636,N_24775,N_26196);
xor U28637 (N_28637,N_24919,N_26697);
or U28638 (N_28638,N_25814,N_24907);
nand U28639 (N_28639,N_24700,N_24214);
nand U28640 (N_28640,N_25659,N_25370);
nor U28641 (N_28641,N_26785,N_24072);
nor U28642 (N_28642,N_25216,N_24393);
nand U28643 (N_28643,N_25878,N_24850);
or U28644 (N_28644,N_25081,N_24293);
and U28645 (N_28645,N_24622,N_24940);
and U28646 (N_28646,N_25566,N_26544);
xnor U28647 (N_28647,N_26912,N_25527);
and U28648 (N_28648,N_25996,N_26816);
or U28649 (N_28649,N_26947,N_26206);
or U28650 (N_28650,N_26828,N_24930);
nor U28651 (N_28651,N_26635,N_26038);
or U28652 (N_28652,N_26956,N_26295);
xnor U28653 (N_28653,N_26351,N_24141);
and U28654 (N_28654,N_24624,N_26503);
or U28655 (N_28655,N_25049,N_24848);
nor U28656 (N_28656,N_25564,N_26661);
nor U28657 (N_28657,N_26871,N_26810);
nand U28658 (N_28658,N_26290,N_26224);
or U28659 (N_28659,N_26358,N_25787);
and U28660 (N_28660,N_24496,N_25825);
and U28661 (N_28661,N_25877,N_26008);
nand U28662 (N_28662,N_25850,N_24271);
and U28663 (N_28663,N_25882,N_26115);
and U28664 (N_28664,N_24285,N_25232);
nand U28665 (N_28665,N_25192,N_24203);
or U28666 (N_28666,N_24045,N_25543);
nand U28667 (N_28667,N_26854,N_24385);
nor U28668 (N_28668,N_24275,N_24092);
and U28669 (N_28669,N_26256,N_24132);
and U28670 (N_28670,N_24890,N_25801);
nor U28671 (N_28671,N_25072,N_25015);
nand U28672 (N_28672,N_24697,N_25836);
nor U28673 (N_28673,N_25017,N_26887);
and U28674 (N_28674,N_26408,N_24976);
and U28675 (N_28675,N_25439,N_25106);
and U28676 (N_28676,N_25608,N_26141);
nand U28677 (N_28677,N_24779,N_26706);
or U28678 (N_28678,N_25448,N_26970);
and U28679 (N_28679,N_26031,N_26130);
nand U28680 (N_28680,N_26934,N_25823);
nor U28681 (N_28681,N_24884,N_25024);
and U28682 (N_28682,N_25641,N_25685);
or U28683 (N_28683,N_26753,N_24803);
xor U28684 (N_28684,N_24188,N_25347);
nand U28685 (N_28685,N_24776,N_24659);
or U28686 (N_28686,N_26272,N_26820);
nor U28687 (N_28687,N_24678,N_26722);
nand U28688 (N_28688,N_25414,N_26538);
nor U28689 (N_28689,N_24126,N_24716);
and U28690 (N_28690,N_25416,N_25017);
xnor U28691 (N_28691,N_26637,N_26414);
and U28692 (N_28692,N_26444,N_26734);
or U28693 (N_28693,N_24254,N_26547);
nor U28694 (N_28694,N_25125,N_26593);
or U28695 (N_28695,N_25844,N_24505);
nor U28696 (N_28696,N_24852,N_26892);
nor U28697 (N_28697,N_25297,N_25435);
nor U28698 (N_28698,N_26453,N_24672);
and U28699 (N_28699,N_25669,N_26395);
or U28700 (N_28700,N_25563,N_25994);
or U28701 (N_28701,N_24400,N_26013);
nand U28702 (N_28702,N_26959,N_25878);
nor U28703 (N_28703,N_24453,N_25688);
nor U28704 (N_28704,N_24447,N_24708);
nor U28705 (N_28705,N_25953,N_24979);
or U28706 (N_28706,N_26759,N_24382);
nand U28707 (N_28707,N_26159,N_24612);
xnor U28708 (N_28708,N_26121,N_26767);
nor U28709 (N_28709,N_24651,N_25141);
nand U28710 (N_28710,N_24869,N_26621);
xor U28711 (N_28711,N_25821,N_25893);
nor U28712 (N_28712,N_26319,N_25469);
and U28713 (N_28713,N_26022,N_26119);
nor U28714 (N_28714,N_26689,N_24587);
nand U28715 (N_28715,N_25096,N_24968);
nand U28716 (N_28716,N_25433,N_24715);
nor U28717 (N_28717,N_26754,N_25638);
nand U28718 (N_28718,N_25047,N_24719);
nand U28719 (N_28719,N_24539,N_26787);
and U28720 (N_28720,N_26518,N_24728);
nand U28721 (N_28721,N_24804,N_26698);
or U28722 (N_28722,N_26299,N_26494);
nand U28723 (N_28723,N_26572,N_25607);
xnor U28724 (N_28724,N_25641,N_26523);
nand U28725 (N_28725,N_25605,N_25190);
and U28726 (N_28726,N_24577,N_25633);
and U28727 (N_28727,N_25517,N_24383);
and U28728 (N_28728,N_26360,N_25737);
and U28729 (N_28729,N_24499,N_26293);
nand U28730 (N_28730,N_26024,N_26809);
nand U28731 (N_28731,N_24420,N_25497);
and U28732 (N_28732,N_24982,N_24858);
or U28733 (N_28733,N_24699,N_25602);
and U28734 (N_28734,N_25672,N_25728);
nand U28735 (N_28735,N_26675,N_26802);
nor U28736 (N_28736,N_25068,N_26917);
or U28737 (N_28737,N_25175,N_26489);
xnor U28738 (N_28738,N_24309,N_24509);
or U28739 (N_28739,N_26438,N_24068);
and U28740 (N_28740,N_24709,N_24216);
or U28741 (N_28741,N_25391,N_26554);
and U28742 (N_28742,N_26695,N_24756);
nand U28743 (N_28743,N_26758,N_24657);
nor U28744 (N_28744,N_25998,N_25705);
or U28745 (N_28745,N_25077,N_26365);
and U28746 (N_28746,N_26885,N_26166);
nor U28747 (N_28747,N_26158,N_26627);
nand U28748 (N_28748,N_26492,N_26908);
and U28749 (N_28749,N_25188,N_26945);
nand U28750 (N_28750,N_26995,N_25062);
and U28751 (N_28751,N_26187,N_24826);
and U28752 (N_28752,N_24629,N_24816);
nand U28753 (N_28753,N_26851,N_24335);
nand U28754 (N_28754,N_25914,N_25869);
nand U28755 (N_28755,N_26002,N_24416);
nand U28756 (N_28756,N_26876,N_24796);
nor U28757 (N_28757,N_26048,N_24210);
nor U28758 (N_28758,N_24238,N_24914);
and U28759 (N_28759,N_24791,N_24781);
or U28760 (N_28760,N_25623,N_25911);
or U28761 (N_28761,N_25647,N_25411);
or U28762 (N_28762,N_26845,N_25289);
nor U28763 (N_28763,N_24409,N_25712);
and U28764 (N_28764,N_25790,N_26143);
nand U28765 (N_28765,N_25716,N_25355);
nand U28766 (N_28766,N_25388,N_26530);
or U28767 (N_28767,N_24934,N_26390);
nor U28768 (N_28768,N_26283,N_25829);
and U28769 (N_28769,N_24600,N_24395);
and U28770 (N_28770,N_25377,N_24287);
xnor U28771 (N_28771,N_25511,N_26257);
nand U28772 (N_28772,N_24002,N_24485);
and U28773 (N_28773,N_25096,N_25963);
xnor U28774 (N_28774,N_26325,N_26524);
nor U28775 (N_28775,N_24434,N_24672);
and U28776 (N_28776,N_25701,N_26735);
xnor U28777 (N_28777,N_25811,N_26903);
nand U28778 (N_28778,N_25352,N_25162);
and U28779 (N_28779,N_26557,N_25050);
nand U28780 (N_28780,N_26833,N_26907);
nor U28781 (N_28781,N_25483,N_25949);
or U28782 (N_28782,N_26110,N_26997);
nor U28783 (N_28783,N_24884,N_26911);
or U28784 (N_28784,N_26389,N_24364);
nor U28785 (N_28785,N_26404,N_25213);
and U28786 (N_28786,N_24315,N_25737);
nand U28787 (N_28787,N_26771,N_26305);
nand U28788 (N_28788,N_24178,N_25127);
nand U28789 (N_28789,N_25920,N_24470);
and U28790 (N_28790,N_25747,N_25694);
nand U28791 (N_28791,N_24116,N_25469);
nor U28792 (N_28792,N_24049,N_26465);
and U28793 (N_28793,N_26147,N_26842);
nor U28794 (N_28794,N_24467,N_25150);
nor U28795 (N_28795,N_24529,N_24092);
xnor U28796 (N_28796,N_24990,N_24628);
nor U28797 (N_28797,N_24285,N_24031);
or U28798 (N_28798,N_24617,N_24552);
or U28799 (N_28799,N_24890,N_25488);
or U28800 (N_28800,N_25700,N_26917);
nand U28801 (N_28801,N_24376,N_25073);
nand U28802 (N_28802,N_26612,N_26563);
nor U28803 (N_28803,N_26850,N_26489);
nand U28804 (N_28804,N_26366,N_26990);
nor U28805 (N_28805,N_25349,N_25825);
nand U28806 (N_28806,N_26112,N_26927);
nand U28807 (N_28807,N_26038,N_24232);
xnor U28808 (N_28808,N_24829,N_25436);
nor U28809 (N_28809,N_24277,N_25905);
nor U28810 (N_28810,N_25180,N_26365);
nand U28811 (N_28811,N_25281,N_24140);
nand U28812 (N_28812,N_25062,N_24789);
nand U28813 (N_28813,N_24934,N_25934);
or U28814 (N_28814,N_24687,N_24861);
and U28815 (N_28815,N_24002,N_24858);
nor U28816 (N_28816,N_26735,N_24876);
xor U28817 (N_28817,N_26299,N_26610);
and U28818 (N_28818,N_25102,N_25668);
nor U28819 (N_28819,N_24095,N_26297);
or U28820 (N_28820,N_25749,N_25589);
or U28821 (N_28821,N_25609,N_26409);
nand U28822 (N_28822,N_25960,N_25663);
nor U28823 (N_28823,N_25634,N_25857);
xnor U28824 (N_28824,N_25993,N_24595);
nand U28825 (N_28825,N_26111,N_25833);
nor U28826 (N_28826,N_25312,N_24408);
or U28827 (N_28827,N_26315,N_24325);
nor U28828 (N_28828,N_26946,N_25460);
or U28829 (N_28829,N_25154,N_24288);
nor U28830 (N_28830,N_25312,N_24569);
nand U28831 (N_28831,N_26078,N_24700);
xor U28832 (N_28832,N_26409,N_26010);
and U28833 (N_28833,N_24010,N_26413);
and U28834 (N_28834,N_25272,N_25791);
nand U28835 (N_28835,N_26993,N_26795);
and U28836 (N_28836,N_25014,N_26171);
or U28837 (N_28837,N_25637,N_24454);
and U28838 (N_28838,N_26349,N_26917);
xor U28839 (N_28839,N_25862,N_26368);
nor U28840 (N_28840,N_25543,N_25830);
nor U28841 (N_28841,N_26432,N_24153);
nand U28842 (N_28842,N_26386,N_24172);
and U28843 (N_28843,N_25762,N_26586);
or U28844 (N_28844,N_26171,N_25844);
and U28845 (N_28845,N_26379,N_26345);
or U28846 (N_28846,N_26824,N_24320);
xor U28847 (N_28847,N_26696,N_25467);
and U28848 (N_28848,N_26287,N_24208);
nand U28849 (N_28849,N_24853,N_25931);
and U28850 (N_28850,N_24960,N_24788);
and U28851 (N_28851,N_24187,N_26085);
and U28852 (N_28852,N_26946,N_26887);
nor U28853 (N_28853,N_24907,N_24690);
or U28854 (N_28854,N_24104,N_24951);
and U28855 (N_28855,N_25068,N_26648);
xor U28856 (N_28856,N_25642,N_26272);
nand U28857 (N_28857,N_24404,N_25314);
nor U28858 (N_28858,N_25763,N_26210);
nand U28859 (N_28859,N_26184,N_26015);
or U28860 (N_28860,N_24140,N_25710);
nand U28861 (N_28861,N_26693,N_24496);
nand U28862 (N_28862,N_25469,N_25983);
nand U28863 (N_28863,N_26005,N_25332);
or U28864 (N_28864,N_24463,N_26929);
or U28865 (N_28865,N_24037,N_25932);
or U28866 (N_28866,N_26772,N_26585);
and U28867 (N_28867,N_26112,N_26948);
nand U28868 (N_28868,N_25631,N_25007);
or U28869 (N_28869,N_24620,N_26221);
and U28870 (N_28870,N_25335,N_25153);
nand U28871 (N_28871,N_26131,N_25309);
nor U28872 (N_28872,N_25859,N_26132);
or U28873 (N_28873,N_26255,N_26328);
and U28874 (N_28874,N_26109,N_25143);
nor U28875 (N_28875,N_24059,N_26922);
or U28876 (N_28876,N_25528,N_26018);
xor U28877 (N_28877,N_26319,N_25048);
xnor U28878 (N_28878,N_26119,N_26577);
nor U28879 (N_28879,N_26742,N_25837);
nor U28880 (N_28880,N_24311,N_24262);
nand U28881 (N_28881,N_25905,N_26466);
or U28882 (N_28882,N_24385,N_24441);
and U28883 (N_28883,N_24867,N_26969);
nand U28884 (N_28884,N_26438,N_26752);
nor U28885 (N_28885,N_26909,N_26899);
xor U28886 (N_28886,N_26055,N_25586);
and U28887 (N_28887,N_25210,N_26165);
nor U28888 (N_28888,N_25073,N_26957);
nand U28889 (N_28889,N_26968,N_24491);
and U28890 (N_28890,N_25850,N_24705);
xor U28891 (N_28891,N_26258,N_25811);
or U28892 (N_28892,N_24566,N_25516);
or U28893 (N_28893,N_24586,N_26786);
and U28894 (N_28894,N_25884,N_26384);
and U28895 (N_28895,N_25385,N_25806);
nand U28896 (N_28896,N_26151,N_24006);
nor U28897 (N_28897,N_25934,N_25621);
nor U28898 (N_28898,N_25401,N_26388);
nand U28899 (N_28899,N_26234,N_25413);
xnor U28900 (N_28900,N_24093,N_26797);
nor U28901 (N_28901,N_26663,N_25569);
and U28902 (N_28902,N_24608,N_24046);
nor U28903 (N_28903,N_24958,N_25349);
nor U28904 (N_28904,N_25310,N_26971);
and U28905 (N_28905,N_24640,N_26202);
nand U28906 (N_28906,N_26092,N_25216);
and U28907 (N_28907,N_24153,N_24579);
nand U28908 (N_28908,N_26219,N_24113);
nor U28909 (N_28909,N_26390,N_24564);
and U28910 (N_28910,N_24850,N_24678);
and U28911 (N_28911,N_26941,N_25427);
or U28912 (N_28912,N_24332,N_24298);
nor U28913 (N_28913,N_25653,N_26132);
nor U28914 (N_28914,N_25084,N_25901);
nor U28915 (N_28915,N_24889,N_24847);
or U28916 (N_28916,N_24509,N_26574);
nand U28917 (N_28917,N_25434,N_25785);
or U28918 (N_28918,N_25369,N_25644);
nand U28919 (N_28919,N_26667,N_24009);
and U28920 (N_28920,N_26365,N_25335);
nor U28921 (N_28921,N_26420,N_24100);
nor U28922 (N_28922,N_24769,N_25044);
and U28923 (N_28923,N_24905,N_25781);
nor U28924 (N_28924,N_24998,N_26459);
and U28925 (N_28925,N_25221,N_24243);
nor U28926 (N_28926,N_26711,N_26135);
xnor U28927 (N_28927,N_26720,N_25668);
and U28928 (N_28928,N_26062,N_25538);
xor U28929 (N_28929,N_25712,N_26325);
nand U28930 (N_28930,N_24135,N_24801);
and U28931 (N_28931,N_25502,N_24652);
and U28932 (N_28932,N_25099,N_26020);
nor U28933 (N_28933,N_25472,N_25030);
or U28934 (N_28934,N_26268,N_24788);
or U28935 (N_28935,N_24652,N_24162);
and U28936 (N_28936,N_25162,N_26428);
nor U28937 (N_28937,N_24857,N_26940);
and U28938 (N_28938,N_24683,N_24047);
and U28939 (N_28939,N_26317,N_25619);
nor U28940 (N_28940,N_24863,N_25781);
or U28941 (N_28941,N_24808,N_25969);
nand U28942 (N_28942,N_24063,N_26336);
nor U28943 (N_28943,N_26934,N_24604);
and U28944 (N_28944,N_26194,N_25033);
and U28945 (N_28945,N_26647,N_26315);
or U28946 (N_28946,N_25542,N_24090);
or U28947 (N_28947,N_24412,N_24298);
or U28948 (N_28948,N_24843,N_24683);
nor U28949 (N_28949,N_25946,N_24970);
and U28950 (N_28950,N_26079,N_24952);
nand U28951 (N_28951,N_24704,N_26726);
or U28952 (N_28952,N_25586,N_24845);
and U28953 (N_28953,N_24429,N_26484);
nor U28954 (N_28954,N_26974,N_25872);
or U28955 (N_28955,N_26234,N_24190);
or U28956 (N_28956,N_25590,N_26428);
nor U28957 (N_28957,N_26891,N_25892);
nand U28958 (N_28958,N_25651,N_24611);
nor U28959 (N_28959,N_24286,N_25208);
nor U28960 (N_28960,N_24176,N_24681);
xnor U28961 (N_28961,N_24070,N_24603);
nand U28962 (N_28962,N_24072,N_25454);
nand U28963 (N_28963,N_26509,N_24894);
and U28964 (N_28964,N_25845,N_25681);
nor U28965 (N_28965,N_26529,N_25383);
nand U28966 (N_28966,N_25545,N_25701);
or U28967 (N_28967,N_24912,N_24995);
nand U28968 (N_28968,N_24856,N_26609);
or U28969 (N_28969,N_24160,N_26998);
and U28970 (N_28970,N_26485,N_25873);
nor U28971 (N_28971,N_25477,N_24919);
nand U28972 (N_28972,N_26609,N_25987);
nand U28973 (N_28973,N_24891,N_25739);
nor U28974 (N_28974,N_26618,N_24392);
xor U28975 (N_28975,N_26616,N_25478);
and U28976 (N_28976,N_25573,N_25205);
nor U28977 (N_28977,N_26547,N_24072);
or U28978 (N_28978,N_26532,N_25477);
and U28979 (N_28979,N_26603,N_26737);
or U28980 (N_28980,N_25741,N_26832);
nand U28981 (N_28981,N_24261,N_26814);
or U28982 (N_28982,N_26705,N_24505);
nor U28983 (N_28983,N_26112,N_26457);
and U28984 (N_28984,N_26887,N_25540);
or U28985 (N_28985,N_25774,N_26853);
and U28986 (N_28986,N_24181,N_24404);
or U28987 (N_28987,N_24563,N_24890);
xor U28988 (N_28988,N_24918,N_26185);
and U28989 (N_28989,N_26707,N_24231);
nand U28990 (N_28990,N_24888,N_26864);
nand U28991 (N_28991,N_24448,N_24879);
and U28992 (N_28992,N_26668,N_24199);
nor U28993 (N_28993,N_24193,N_26642);
and U28994 (N_28994,N_25886,N_26230);
or U28995 (N_28995,N_25971,N_24898);
or U28996 (N_28996,N_26186,N_25605);
nor U28997 (N_28997,N_26985,N_25866);
or U28998 (N_28998,N_26626,N_26077);
and U28999 (N_28999,N_25782,N_25188);
nor U29000 (N_29000,N_25358,N_25418);
nand U29001 (N_29001,N_24403,N_26433);
nand U29002 (N_29002,N_24382,N_26972);
or U29003 (N_29003,N_24742,N_25034);
nor U29004 (N_29004,N_24998,N_25505);
nor U29005 (N_29005,N_24520,N_25817);
xnor U29006 (N_29006,N_25699,N_26618);
or U29007 (N_29007,N_26002,N_24771);
or U29008 (N_29008,N_25297,N_25888);
or U29009 (N_29009,N_24132,N_25751);
or U29010 (N_29010,N_25786,N_24960);
nand U29011 (N_29011,N_25388,N_26070);
xnor U29012 (N_29012,N_25770,N_25420);
nor U29013 (N_29013,N_25954,N_26295);
xnor U29014 (N_29014,N_26858,N_24563);
and U29015 (N_29015,N_26280,N_25666);
xnor U29016 (N_29016,N_26751,N_24030);
xnor U29017 (N_29017,N_25214,N_24840);
or U29018 (N_29018,N_25124,N_24926);
xnor U29019 (N_29019,N_24829,N_24125);
xor U29020 (N_29020,N_25973,N_26689);
nand U29021 (N_29021,N_26603,N_26457);
or U29022 (N_29022,N_25455,N_24542);
nor U29023 (N_29023,N_25871,N_24077);
xor U29024 (N_29024,N_25326,N_25308);
nor U29025 (N_29025,N_25941,N_25535);
nor U29026 (N_29026,N_26245,N_26354);
nand U29027 (N_29027,N_26435,N_26891);
nor U29028 (N_29028,N_26337,N_25833);
xor U29029 (N_29029,N_25021,N_24094);
or U29030 (N_29030,N_24809,N_25442);
xor U29031 (N_29031,N_26585,N_24305);
xnor U29032 (N_29032,N_26702,N_24416);
and U29033 (N_29033,N_24056,N_24847);
and U29034 (N_29034,N_25745,N_24131);
nand U29035 (N_29035,N_24836,N_26232);
nand U29036 (N_29036,N_25980,N_24997);
and U29037 (N_29037,N_24861,N_24013);
nand U29038 (N_29038,N_26200,N_24476);
xor U29039 (N_29039,N_24891,N_25305);
nor U29040 (N_29040,N_24847,N_25826);
nor U29041 (N_29041,N_25156,N_25531);
nor U29042 (N_29042,N_25997,N_24370);
nand U29043 (N_29043,N_25232,N_25604);
xor U29044 (N_29044,N_26371,N_26253);
or U29045 (N_29045,N_24772,N_25442);
xnor U29046 (N_29046,N_26929,N_26938);
xor U29047 (N_29047,N_24275,N_25436);
nand U29048 (N_29048,N_24016,N_24447);
xnor U29049 (N_29049,N_26076,N_26864);
nor U29050 (N_29050,N_26353,N_26693);
xor U29051 (N_29051,N_24380,N_24465);
and U29052 (N_29052,N_25166,N_26877);
xor U29053 (N_29053,N_24512,N_24380);
or U29054 (N_29054,N_26900,N_24194);
or U29055 (N_29055,N_26088,N_24632);
nor U29056 (N_29056,N_24749,N_25176);
nand U29057 (N_29057,N_25613,N_26731);
nor U29058 (N_29058,N_25947,N_24239);
nand U29059 (N_29059,N_24447,N_26445);
nor U29060 (N_29060,N_24165,N_24251);
or U29061 (N_29061,N_26533,N_25951);
and U29062 (N_29062,N_26532,N_25378);
and U29063 (N_29063,N_26104,N_26285);
nand U29064 (N_29064,N_24849,N_24827);
or U29065 (N_29065,N_25474,N_25697);
nor U29066 (N_29066,N_26717,N_26269);
or U29067 (N_29067,N_24257,N_24020);
nand U29068 (N_29068,N_26180,N_24218);
nand U29069 (N_29069,N_24193,N_25968);
and U29070 (N_29070,N_26822,N_25385);
nand U29071 (N_29071,N_25884,N_24856);
nor U29072 (N_29072,N_26921,N_25084);
nor U29073 (N_29073,N_24662,N_26781);
and U29074 (N_29074,N_26041,N_26218);
and U29075 (N_29075,N_24183,N_24215);
xnor U29076 (N_29076,N_25426,N_26128);
nand U29077 (N_29077,N_26202,N_25059);
nand U29078 (N_29078,N_25977,N_25236);
or U29079 (N_29079,N_26782,N_24739);
and U29080 (N_29080,N_25326,N_26931);
nor U29081 (N_29081,N_24702,N_25474);
and U29082 (N_29082,N_24844,N_26701);
nor U29083 (N_29083,N_24535,N_25187);
or U29084 (N_29084,N_25911,N_24220);
or U29085 (N_29085,N_24739,N_26236);
nand U29086 (N_29086,N_24355,N_25522);
nand U29087 (N_29087,N_26933,N_26336);
nand U29088 (N_29088,N_26916,N_25939);
or U29089 (N_29089,N_26699,N_25411);
and U29090 (N_29090,N_25313,N_24132);
nor U29091 (N_29091,N_26211,N_26374);
nand U29092 (N_29092,N_24689,N_26927);
or U29093 (N_29093,N_26481,N_25917);
nand U29094 (N_29094,N_24984,N_25723);
nand U29095 (N_29095,N_26750,N_24399);
or U29096 (N_29096,N_26195,N_24065);
or U29097 (N_29097,N_26780,N_26910);
nand U29098 (N_29098,N_24387,N_24869);
nor U29099 (N_29099,N_24196,N_26642);
and U29100 (N_29100,N_24091,N_26544);
and U29101 (N_29101,N_24447,N_26762);
or U29102 (N_29102,N_24617,N_26625);
or U29103 (N_29103,N_24919,N_26434);
or U29104 (N_29104,N_26226,N_26590);
and U29105 (N_29105,N_25689,N_24197);
and U29106 (N_29106,N_24499,N_25463);
or U29107 (N_29107,N_24921,N_24575);
and U29108 (N_29108,N_25717,N_25134);
or U29109 (N_29109,N_26152,N_25166);
or U29110 (N_29110,N_24132,N_26633);
nor U29111 (N_29111,N_26073,N_26050);
or U29112 (N_29112,N_26562,N_25903);
nor U29113 (N_29113,N_24414,N_24807);
and U29114 (N_29114,N_25295,N_24958);
nand U29115 (N_29115,N_24098,N_26364);
and U29116 (N_29116,N_25484,N_24711);
nor U29117 (N_29117,N_26789,N_26550);
or U29118 (N_29118,N_25115,N_25913);
nand U29119 (N_29119,N_26203,N_26028);
and U29120 (N_29120,N_25413,N_26261);
nor U29121 (N_29121,N_24193,N_24212);
nand U29122 (N_29122,N_25384,N_25004);
nand U29123 (N_29123,N_26113,N_26990);
or U29124 (N_29124,N_24729,N_24132);
or U29125 (N_29125,N_25657,N_24847);
nand U29126 (N_29126,N_26068,N_24389);
and U29127 (N_29127,N_25060,N_24108);
xor U29128 (N_29128,N_24071,N_25802);
nor U29129 (N_29129,N_26077,N_25512);
and U29130 (N_29130,N_26802,N_26084);
xor U29131 (N_29131,N_25580,N_26533);
and U29132 (N_29132,N_25180,N_25152);
nand U29133 (N_29133,N_26930,N_24097);
xor U29134 (N_29134,N_26453,N_24340);
nor U29135 (N_29135,N_26572,N_25205);
nand U29136 (N_29136,N_24969,N_24654);
or U29137 (N_29137,N_26816,N_25253);
nand U29138 (N_29138,N_24656,N_24850);
nor U29139 (N_29139,N_25313,N_24240);
nand U29140 (N_29140,N_25489,N_26943);
nand U29141 (N_29141,N_25284,N_26959);
xor U29142 (N_29142,N_24678,N_24698);
nor U29143 (N_29143,N_26606,N_25909);
or U29144 (N_29144,N_25850,N_26601);
nor U29145 (N_29145,N_25012,N_24869);
nor U29146 (N_29146,N_24074,N_25807);
nor U29147 (N_29147,N_24577,N_24756);
nand U29148 (N_29148,N_24237,N_24060);
nand U29149 (N_29149,N_24273,N_25690);
nand U29150 (N_29150,N_26885,N_26494);
and U29151 (N_29151,N_24772,N_24185);
nor U29152 (N_29152,N_26615,N_26178);
nor U29153 (N_29153,N_25904,N_26977);
nand U29154 (N_29154,N_24713,N_26202);
or U29155 (N_29155,N_26688,N_25487);
nand U29156 (N_29156,N_26298,N_26506);
xor U29157 (N_29157,N_25260,N_26070);
or U29158 (N_29158,N_26303,N_26393);
or U29159 (N_29159,N_24462,N_24045);
and U29160 (N_29160,N_24954,N_26558);
nand U29161 (N_29161,N_24407,N_26612);
or U29162 (N_29162,N_26749,N_26111);
nand U29163 (N_29163,N_25025,N_26374);
or U29164 (N_29164,N_25579,N_24768);
or U29165 (N_29165,N_24394,N_24041);
and U29166 (N_29166,N_24954,N_26914);
or U29167 (N_29167,N_25648,N_26527);
nor U29168 (N_29168,N_24379,N_25517);
nor U29169 (N_29169,N_25398,N_25138);
and U29170 (N_29170,N_25041,N_24409);
nor U29171 (N_29171,N_24678,N_26035);
nand U29172 (N_29172,N_25972,N_25367);
or U29173 (N_29173,N_24857,N_24601);
and U29174 (N_29174,N_25327,N_25858);
or U29175 (N_29175,N_25536,N_25379);
or U29176 (N_29176,N_25857,N_24641);
nor U29177 (N_29177,N_25945,N_26833);
nor U29178 (N_29178,N_24947,N_24491);
nand U29179 (N_29179,N_26791,N_26604);
nand U29180 (N_29180,N_24233,N_24249);
nand U29181 (N_29181,N_24163,N_24682);
and U29182 (N_29182,N_25603,N_26517);
nor U29183 (N_29183,N_24160,N_26183);
or U29184 (N_29184,N_26105,N_26392);
or U29185 (N_29185,N_25324,N_26634);
nor U29186 (N_29186,N_26720,N_26041);
nor U29187 (N_29187,N_24743,N_24879);
nor U29188 (N_29188,N_25132,N_25063);
or U29189 (N_29189,N_24005,N_26310);
nor U29190 (N_29190,N_25141,N_24015);
nor U29191 (N_29191,N_25815,N_24887);
and U29192 (N_29192,N_24864,N_25337);
or U29193 (N_29193,N_26186,N_24168);
nand U29194 (N_29194,N_24682,N_25849);
nand U29195 (N_29195,N_26229,N_24735);
or U29196 (N_29196,N_26458,N_26908);
or U29197 (N_29197,N_24139,N_24491);
nor U29198 (N_29198,N_24705,N_25096);
and U29199 (N_29199,N_25350,N_24264);
and U29200 (N_29200,N_26218,N_25617);
nor U29201 (N_29201,N_25776,N_24102);
and U29202 (N_29202,N_25517,N_25816);
and U29203 (N_29203,N_24491,N_26277);
nand U29204 (N_29204,N_24992,N_24024);
xor U29205 (N_29205,N_24602,N_25320);
nand U29206 (N_29206,N_25498,N_24269);
xor U29207 (N_29207,N_26292,N_24653);
and U29208 (N_29208,N_26405,N_25228);
and U29209 (N_29209,N_26656,N_25638);
or U29210 (N_29210,N_24115,N_25156);
or U29211 (N_29211,N_25905,N_25143);
and U29212 (N_29212,N_26535,N_26577);
xnor U29213 (N_29213,N_25181,N_24187);
xor U29214 (N_29214,N_26286,N_25068);
nor U29215 (N_29215,N_25862,N_24173);
nand U29216 (N_29216,N_25917,N_25519);
nor U29217 (N_29217,N_26445,N_24603);
nand U29218 (N_29218,N_24701,N_24268);
nor U29219 (N_29219,N_25644,N_26143);
or U29220 (N_29220,N_24520,N_24424);
or U29221 (N_29221,N_25279,N_24133);
nand U29222 (N_29222,N_25681,N_25601);
or U29223 (N_29223,N_24926,N_25649);
or U29224 (N_29224,N_24123,N_24142);
nor U29225 (N_29225,N_25098,N_25570);
and U29226 (N_29226,N_24109,N_24772);
and U29227 (N_29227,N_24351,N_24320);
or U29228 (N_29228,N_25690,N_25116);
xor U29229 (N_29229,N_25552,N_25754);
or U29230 (N_29230,N_25360,N_25635);
nand U29231 (N_29231,N_24520,N_26648);
nand U29232 (N_29232,N_24665,N_25989);
or U29233 (N_29233,N_24631,N_24949);
nor U29234 (N_29234,N_26791,N_24559);
xnor U29235 (N_29235,N_24879,N_26902);
or U29236 (N_29236,N_25840,N_25542);
or U29237 (N_29237,N_25824,N_25316);
and U29238 (N_29238,N_24930,N_25706);
nor U29239 (N_29239,N_24240,N_26640);
or U29240 (N_29240,N_26222,N_24268);
nor U29241 (N_29241,N_26967,N_26409);
or U29242 (N_29242,N_24530,N_26180);
and U29243 (N_29243,N_25560,N_26536);
or U29244 (N_29244,N_26700,N_25314);
nor U29245 (N_29245,N_24054,N_24254);
nor U29246 (N_29246,N_24491,N_24808);
nor U29247 (N_29247,N_26235,N_25678);
nor U29248 (N_29248,N_26951,N_24854);
nor U29249 (N_29249,N_24943,N_24245);
nand U29250 (N_29250,N_24866,N_25736);
nor U29251 (N_29251,N_24506,N_26264);
and U29252 (N_29252,N_24131,N_26436);
nand U29253 (N_29253,N_24773,N_26428);
or U29254 (N_29254,N_25172,N_26959);
and U29255 (N_29255,N_25411,N_25614);
nand U29256 (N_29256,N_25849,N_24063);
nor U29257 (N_29257,N_26950,N_24407);
nor U29258 (N_29258,N_25986,N_24128);
nand U29259 (N_29259,N_25496,N_24980);
and U29260 (N_29260,N_25179,N_26937);
or U29261 (N_29261,N_25269,N_24438);
or U29262 (N_29262,N_25169,N_25533);
nor U29263 (N_29263,N_26857,N_24269);
nand U29264 (N_29264,N_25969,N_25520);
or U29265 (N_29265,N_24431,N_26394);
nand U29266 (N_29266,N_24705,N_24134);
and U29267 (N_29267,N_24086,N_26785);
nand U29268 (N_29268,N_26218,N_26521);
and U29269 (N_29269,N_24185,N_25618);
and U29270 (N_29270,N_25469,N_26509);
nor U29271 (N_29271,N_24416,N_25469);
xor U29272 (N_29272,N_25791,N_26044);
nand U29273 (N_29273,N_24531,N_26754);
and U29274 (N_29274,N_26044,N_25085);
and U29275 (N_29275,N_26322,N_25327);
nor U29276 (N_29276,N_24249,N_24323);
nand U29277 (N_29277,N_24044,N_26341);
nand U29278 (N_29278,N_24703,N_25038);
nand U29279 (N_29279,N_25888,N_26213);
nand U29280 (N_29280,N_25555,N_26789);
nand U29281 (N_29281,N_26165,N_25033);
and U29282 (N_29282,N_25875,N_25518);
nor U29283 (N_29283,N_24935,N_24246);
or U29284 (N_29284,N_25133,N_25649);
and U29285 (N_29285,N_24676,N_24505);
nand U29286 (N_29286,N_25099,N_25754);
and U29287 (N_29287,N_25349,N_24577);
xnor U29288 (N_29288,N_24884,N_24138);
xnor U29289 (N_29289,N_26402,N_26287);
nor U29290 (N_29290,N_25891,N_24895);
xnor U29291 (N_29291,N_26736,N_24188);
xor U29292 (N_29292,N_24535,N_25550);
nor U29293 (N_29293,N_26128,N_25185);
or U29294 (N_29294,N_24099,N_24041);
and U29295 (N_29295,N_26020,N_24530);
nor U29296 (N_29296,N_26015,N_26461);
nand U29297 (N_29297,N_24653,N_24835);
or U29298 (N_29298,N_24369,N_24573);
or U29299 (N_29299,N_26450,N_26842);
xnor U29300 (N_29300,N_25458,N_24751);
nand U29301 (N_29301,N_26809,N_26472);
or U29302 (N_29302,N_24996,N_24199);
or U29303 (N_29303,N_25358,N_25115);
nor U29304 (N_29304,N_26813,N_24315);
or U29305 (N_29305,N_25374,N_25591);
and U29306 (N_29306,N_24571,N_24622);
or U29307 (N_29307,N_24586,N_24233);
or U29308 (N_29308,N_24865,N_24646);
and U29309 (N_29309,N_25351,N_24779);
nor U29310 (N_29310,N_25864,N_24676);
or U29311 (N_29311,N_26528,N_24080);
nand U29312 (N_29312,N_24080,N_26397);
and U29313 (N_29313,N_25247,N_26499);
or U29314 (N_29314,N_25751,N_24978);
nand U29315 (N_29315,N_24827,N_24670);
nor U29316 (N_29316,N_25609,N_24852);
or U29317 (N_29317,N_24137,N_24595);
nor U29318 (N_29318,N_26454,N_26981);
or U29319 (N_29319,N_24006,N_26702);
nor U29320 (N_29320,N_25435,N_25819);
and U29321 (N_29321,N_25849,N_24393);
nor U29322 (N_29322,N_26829,N_26809);
nor U29323 (N_29323,N_26175,N_26578);
and U29324 (N_29324,N_26914,N_26130);
xnor U29325 (N_29325,N_26688,N_24017);
nor U29326 (N_29326,N_25327,N_25721);
and U29327 (N_29327,N_25819,N_26637);
nand U29328 (N_29328,N_25292,N_26901);
xnor U29329 (N_29329,N_26779,N_26906);
and U29330 (N_29330,N_25414,N_25991);
nand U29331 (N_29331,N_24893,N_26465);
nand U29332 (N_29332,N_25466,N_24214);
and U29333 (N_29333,N_24365,N_24614);
nor U29334 (N_29334,N_24976,N_24458);
xor U29335 (N_29335,N_26156,N_26032);
nor U29336 (N_29336,N_25353,N_25193);
nor U29337 (N_29337,N_26779,N_24750);
xor U29338 (N_29338,N_26471,N_26010);
nor U29339 (N_29339,N_26524,N_26292);
nor U29340 (N_29340,N_24067,N_24845);
nor U29341 (N_29341,N_25203,N_25355);
nor U29342 (N_29342,N_25053,N_25643);
or U29343 (N_29343,N_26967,N_26676);
xnor U29344 (N_29344,N_26426,N_26774);
and U29345 (N_29345,N_25611,N_25918);
nand U29346 (N_29346,N_24859,N_26917);
or U29347 (N_29347,N_24392,N_25319);
or U29348 (N_29348,N_26565,N_25225);
and U29349 (N_29349,N_24381,N_26950);
nand U29350 (N_29350,N_24447,N_25739);
nand U29351 (N_29351,N_24127,N_26660);
nand U29352 (N_29352,N_26874,N_26738);
or U29353 (N_29353,N_25087,N_25423);
nand U29354 (N_29354,N_25510,N_26320);
and U29355 (N_29355,N_26345,N_26370);
nand U29356 (N_29356,N_26243,N_26764);
nor U29357 (N_29357,N_24959,N_25061);
and U29358 (N_29358,N_24814,N_25128);
and U29359 (N_29359,N_24791,N_26647);
xor U29360 (N_29360,N_25619,N_26933);
or U29361 (N_29361,N_26023,N_24734);
nand U29362 (N_29362,N_26955,N_25511);
and U29363 (N_29363,N_24255,N_25665);
or U29364 (N_29364,N_26664,N_25743);
or U29365 (N_29365,N_25792,N_25037);
and U29366 (N_29366,N_25037,N_25449);
nand U29367 (N_29367,N_25890,N_26080);
nor U29368 (N_29368,N_26508,N_25670);
or U29369 (N_29369,N_26081,N_24778);
and U29370 (N_29370,N_24142,N_25613);
nor U29371 (N_29371,N_24232,N_25834);
or U29372 (N_29372,N_26110,N_25150);
nand U29373 (N_29373,N_26824,N_25534);
nand U29374 (N_29374,N_24921,N_24992);
nor U29375 (N_29375,N_26033,N_24183);
or U29376 (N_29376,N_24150,N_26830);
nand U29377 (N_29377,N_24346,N_24343);
xnor U29378 (N_29378,N_25868,N_24954);
xor U29379 (N_29379,N_24368,N_26359);
or U29380 (N_29380,N_24973,N_24012);
or U29381 (N_29381,N_26958,N_25164);
or U29382 (N_29382,N_24274,N_26222);
nand U29383 (N_29383,N_24227,N_25250);
nor U29384 (N_29384,N_25204,N_26489);
nor U29385 (N_29385,N_25252,N_26013);
and U29386 (N_29386,N_25482,N_26765);
nand U29387 (N_29387,N_26826,N_24073);
and U29388 (N_29388,N_26524,N_24754);
nand U29389 (N_29389,N_24990,N_26956);
and U29390 (N_29390,N_24550,N_24348);
or U29391 (N_29391,N_24105,N_26895);
nor U29392 (N_29392,N_24328,N_25921);
nor U29393 (N_29393,N_25215,N_25799);
nand U29394 (N_29394,N_26314,N_25620);
or U29395 (N_29395,N_25459,N_26532);
nand U29396 (N_29396,N_25465,N_26618);
nor U29397 (N_29397,N_25570,N_24168);
nor U29398 (N_29398,N_26090,N_26707);
nand U29399 (N_29399,N_24298,N_24163);
nand U29400 (N_29400,N_26163,N_24854);
xor U29401 (N_29401,N_26262,N_24024);
xnor U29402 (N_29402,N_25698,N_26368);
and U29403 (N_29403,N_25478,N_24666);
or U29404 (N_29404,N_25971,N_26315);
nor U29405 (N_29405,N_24664,N_24352);
and U29406 (N_29406,N_24310,N_24735);
and U29407 (N_29407,N_26688,N_24970);
nor U29408 (N_29408,N_25595,N_24613);
and U29409 (N_29409,N_26285,N_25910);
nor U29410 (N_29410,N_25686,N_24340);
and U29411 (N_29411,N_24725,N_25657);
nand U29412 (N_29412,N_24371,N_25130);
and U29413 (N_29413,N_26696,N_26121);
nor U29414 (N_29414,N_25782,N_25238);
and U29415 (N_29415,N_24703,N_24564);
nor U29416 (N_29416,N_24495,N_25408);
or U29417 (N_29417,N_26162,N_24787);
or U29418 (N_29418,N_24111,N_25319);
and U29419 (N_29419,N_24706,N_26221);
and U29420 (N_29420,N_26537,N_24245);
or U29421 (N_29421,N_26230,N_26827);
nor U29422 (N_29422,N_25045,N_26383);
xor U29423 (N_29423,N_24462,N_26118);
and U29424 (N_29424,N_26962,N_25028);
nor U29425 (N_29425,N_25630,N_26927);
xor U29426 (N_29426,N_25357,N_26464);
and U29427 (N_29427,N_25040,N_24141);
nand U29428 (N_29428,N_24197,N_25947);
or U29429 (N_29429,N_25070,N_25030);
nor U29430 (N_29430,N_25539,N_26525);
nor U29431 (N_29431,N_26529,N_26349);
and U29432 (N_29432,N_24339,N_24318);
and U29433 (N_29433,N_25523,N_24151);
nor U29434 (N_29434,N_26869,N_25953);
nand U29435 (N_29435,N_26545,N_26444);
or U29436 (N_29436,N_25612,N_24088);
xnor U29437 (N_29437,N_25305,N_24183);
and U29438 (N_29438,N_24815,N_26030);
nor U29439 (N_29439,N_25496,N_26486);
or U29440 (N_29440,N_24711,N_26582);
nor U29441 (N_29441,N_24792,N_25053);
and U29442 (N_29442,N_26546,N_24390);
xor U29443 (N_29443,N_26398,N_26518);
or U29444 (N_29444,N_25966,N_24895);
or U29445 (N_29445,N_25393,N_24447);
or U29446 (N_29446,N_24347,N_26559);
nand U29447 (N_29447,N_24945,N_26715);
nor U29448 (N_29448,N_25844,N_25665);
and U29449 (N_29449,N_26089,N_26191);
or U29450 (N_29450,N_24931,N_25915);
nor U29451 (N_29451,N_25778,N_25652);
and U29452 (N_29452,N_25316,N_24950);
nor U29453 (N_29453,N_25453,N_24194);
and U29454 (N_29454,N_25521,N_26675);
xnor U29455 (N_29455,N_26532,N_25568);
or U29456 (N_29456,N_26370,N_26338);
xor U29457 (N_29457,N_25185,N_26509);
nand U29458 (N_29458,N_24599,N_25224);
xnor U29459 (N_29459,N_25996,N_24438);
and U29460 (N_29460,N_26724,N_24158);
xnor U29461 (N_29461,N_25953,N_25718);
and U29462 (N_29462,N_26870,N_26604);
xnor U29463 (N_29463,N_25805,N_24247);
or U29464 (N_29464,N_24397,N_25426);
nor U29465 (N_29465,N_25375,N_25392);
nor U29466 (N_29466,N_25485,N_24184);
nand U29467 (N_29467,N_24113,N_25135);
and U29468 (N_29468,N_25010,N_24445);
or U29469 (N_29469,N_26118,N_26803);
nand U29470 (N_29470,N_25537,N_24508);
or U29471 (N_29471,N_25271,N_24623);
or U29472 (N_29472,N_24828,N_26739);
nor U29473 (N_29473,N_24236,N_25331);
nand U29474 (N_29474,N_26835,N_25989);
nor U29475 (N_29475,N_26684,N_24568);
nand U29476 (N_29476,N_25705,N_24379);
and U29477 (N_29477,N_26676,N_25058);
or U29478 (N_29478,N_24947,N_25681);
and U29479 (N_29479,N_25303,N_24517);
nand U29480 (N_29480,N_26451,N_26406);
nor U29481 (N_29481,N_26448,N_25901);
nor U29482 (N_29482,N_25007,N_25024);
xnor U29483 (N_29483,N_26252,N_26815);
nor U29484 (N_29484,N_26213,N_26132);
nand U29485 (N_29485,N_26977,N_24442);
and U29486 (N_29486,N_26483,N_24740);
nor U29487 (N_29487,N_24730,N_24763);
and U29488 (N_29488,N_24674,N_24661);
or U29489 (N_29489,N_26595,N_26607);
xor U29490 (N_29490,N_26295,N_25513);
nor U29491 (N_29491,N_26376,N_26406);
or U29492 (N_29492,N_26826,N_24980);
nand U29493 (N_29493,N_25334,N_25078);
or U29494 (N_29494,N_25035,N_26875);
xnor U29495 (N_29495,N_26511,N_24604);
or U29496 (N_29496,N_26514,N_26226);
nand U29497 (N_29497,N_24761,N_26674);
and U29498 (N_29498,N_24207,N_24719);
nand U29499 (N_29499,N_26267,N_26312);
or U29500 (N_29500,N_25082,N_25805);
nand U29501 (N_29501,N_25506,N_26658);
nand U29502 (N_29502,N_24389,N_24606);
nor U29503 (N_29503,N_25781,N_26594);
or U29504 (N_29504,N_24256,N_25470);
or U29505 (N_29505,N_24907,N_25054);
nand U29506 (N_29506,N_24068,N_24498);
and U29507 (N_29507,N_25403,N_26279);
nor U29508 (N_29508,N_24557,N_24945);
and U29509 (N_29509,N_25145,N_25434);
nand U29510 (N_29510,N_26174,N_24671);
or U29511 (N_29511,N_25259,N_25387);
and U29512 (N_29512,N_26728,N_24051);
nand U29513 (N_29513,N_24637,N_24902);
and U29514 (N_29514,N_26801,N_26571);
or U29515 (N_29515,N_25682,N_25525);
nor U29516 (N_29516,N_26098,N_24584);
nor U29517 (N_29517,N_24094,N_25173);
nor U29518 (N_29518,N_25477,N_26741);
nor U29519 (N_29519,N_24581,N_24357);
nor U29520 (N_29520,N_26324,N_26051);
or U29521 (N_29521,N_25461,N_24458);
and U29522 (N_29522,N_25961,N_25906);
and U29523 (N_29523,N_24643,N_24815);
and U29524 (N_29524,N_25629,N_25916);
nor U29525 (N_29525,N_26221,N_25855);
nand U29526 (N_29526,N_25316,N_26129);
nor U29527 (N_29527,N_24397,N_24279);
xor U29528 (N_29528,N_26747,N_24905);
or U29529 (N_29529,N_24075,N_26807);
or U29530 (N_29530,N_26192,N_26662);
nor U29531 (N_29531,N_25588,N_25098);
xnor U29532 (N_29532,N_26130,N_24229);
or U29533 (N_29533,N_24673,N_25008);
nand U29534 (N_29534,N_24740,N_24686);
nand U29535 (N_29535,N_25534,N_26592);
and U29536 (N_29536,N_26888,N_26184);
nor U29537 (N_29537,N_24208,N_24659);
nor U29538 (N_29538,N_24128,N_26119);
nor U29539 (N_29539,N_25142,N_24507);
nand U29540 (N_29540,N_24420,N_24251);
nand U29541 (N_29541,N_25883,N_24705);
nor U29542 (N_29542,N_25295,N_26932);
or U29543 (N_29543,N_24565,N_25153);
nand U29544 (N_29544,N_24278,N_24522);
or U29545 (N_29545,N_26553,N_26028);
or U29546 (N_29546,N_24775,N_26537);
or U29547 (N_29547,N_25726,N_26803);
nand U29548 (N_29548,N_24514,N_24119);
nand U29549 (N_29549,N_24133,N_25268);
xnor U29550 (N_29550,N_25209,N_25754);
nor U29551 (N_29551,N_25875,N_24916);
nand U29552 (N_29552,N_24195,N_25355);
or U29553 (N_29553,N_25646,N_25816);
or U29554 (N_29554,N_25644,N_24332);
nand U29555 (N_29555,N_26634,N_24875);
nand U29556 (N_29556,N_25775,N_25363);
and U29557 (N_29557,N_26073,N_25087);
or U29558 (N_29558,N_26419,N_24552);
nor U29559 (N_29559,N_25943,N_24409);
nand U29560 (N_29560,N_24517,N_25146);
or U29561 (N_29561,N_26068,N_24611);
nor U29562 (N_29562,N_25658,N_26258);
nor U29563 (N_29563,N_24413,N_24158);
xor U29564 (N_29564,N_26370,N_24748);
nor U29565 (N_29565,N_25180,N_25760);
and U29566 (N_29566,N_26736,N_24276);
and U29567 (N_29567,N_26178,N_26502);
and U29568 (N_29568,N_25618,N_25511);
or U29569 (N_29569,N_26731,N_24826);
xor U29570 (N_29570,N_25821,N_26269);
nor U29571 (N_29571,N_24672,N_25802);
nor U29572 (N_29572,N_24320,N_24099);
xor U29573 (N_29573,N_25596,N_24164);
nand U29574 (N_29574,N_25126,N_26080);
nor U29575 (N_29575,N_26859,N_25182);
and U29576 (N_29576,N_25474,N_24673);
nor U29577 (N_29577,N_26587,N_25296);
and U29578 (N_29578,N_25501,N_25687);
nor U29579 (N_29579,N_25048,N_24712);
nor U29580 (N_29580,N_26041,N_24126);
xor U29581 (N_29581,N_24620,N_25698);
nor U29582 (N_29582,N_25725,N_24411);
and U29583 (N_29583,N_24931,N_24364);
nand U29584 (N_29584,N_25212,N_24196);
nor U29585 (N_29585,N_24721,N_24785);
nand U29586 (N_29586,N_24398,N_24014);
nor U29587 (N_29587,N_25091,N_24009);
nand U29588 (N_29588,N_25212,N_24157);
and U29589 (N_29589,N_24234,N_24457);
and U29590 (N_29590,N_26961,N_25685);
or U29591 (N_29591,N_24705,N_25831);
and U29592 (N_29592,N_26130,N_24047);
and U29593 (N_29593,N_24496,N_24352);
nor U29594 (N_29594,N_26704,N_25121);
xnor U29595 (N_29595,N_25908,N_24701);
nor U29596 (N_29596,N_24573,N_24750);
nand U29597 (N_29597,N_24212,N_26018);
and U29598 (N_29598,N_24578,N_24833);
xnor U29599 (N_29599,N_26013,N_25556);
xor U29600 (N_29600,N_25850,N_24593);
nand U29601 (N_29601,N_24655,N_26171);
and U29602 (N_29602,N_24249,N_26109);
and U29603 (N_29603,N_26701,N_26089);
and U29604 (N_29604,N_25297,N_24757);
nand U29605 (N_29605,N_24327,N_26957);
nor U29606 (N_29606,N_25464,N_26451);
nand U29607 (N_29607,N_26937,N_25850);
nor U29608 (N_29608,N_24839,N_24946);
or U29609 (N_29609,N_26823,N_24147);
or U29610 (N_29610,N_24367,N_25257);
or U29611 (N_29611,N_24400,N_26091);
and U29612 (N_29612,N_26802,N_24576);
xnor U29613 (N_29613,N_25367,N_26638);
or U29614 (N_29614,N_26380,N_26525);
nor U29615 (N_29615,N_25966,N_25394);
nor U29616 (N_29616,N_25897,N_26784);
or U29617 (N_29617,N_24340,N_26110);
and U29618 (N_29618,N_24198,N_26843);
or U29619 (N_29619,N_26593,N_24552);
nor U29620 (N_29620,N_26290,N_26745);
nor U29621 (N_29621,N_25150,N_26353);
or U29622 (N_29622,N_24115,N_26587);
xor U29623 (N_29623,N_25897,N_25880);
nor U29624 (N_29624,N_26753,N_24856);
nand U29625 (N_29625,N_25087,N_24153);
and U29626 (N_29626,N_24551,N_24222);
nor U29627 (N_29627,N_24791,N_24409);
and U29628 (N_29628,N_26486,N_26585);
nor U29629 (N_29629,N_26875,N_25493);
or U29630 (N_29630,N_24918,N_26998);
nand U29631 (N_29631,N_26443,N_24611);
or U29632 (N_29632,N_26439,N_26142);
and U29633 (N_29633,N_26117,N_25686);
and U29634 (N_29634,N_25623,N_25537);
nand U29635 (N_29635,N_26326,N_26368);
nor U29636 (N_29636,N_24679,N_25606);
or U29637 (N_29637,N_24254,N_26097);
nor U29638 (N_29638,N_25321,N_26695);
and U29639 (N_29639,N_24456,N_25536);
nor U29640 (N_29640,N_26000,N_26904);
xor U29641 (N_29641,N_24883,N_24190);
nor U29642 (N_29642,N_24287,N_26150);
or U29643 (N_29643,N_26924,N_24064);
or U29644 (N_29644,N_24589,N_24448);
nor U29645 (N_29645,N_26006,N_26580);
or U29646 (N_29646,N_24607,N_26986);
and U29647 (N_29647,N_26005,N_26150);
nor U29648 (N_29648,N_25508,N_24784);
or U29649 (N_29649,N_25933,N_25742);
or U29650 (N_29650,N_24193,N_25046);
nor U29651 (N_29651,N_24867,N_26449);
or U29652 (N_29652,N_25700,N_24911);
xor U29653 (N_29653,N_25745,N_25355);
nand U29654 (N_29654,N_24953,N_26871);
xnor U29655 (N_29655,N_24027,N_25009);
nor U29656 (N_29656,N_25148,N_26084);
nand U29657 (N_29657,N_25252,N_26437);
nand U29658 (N_29658,N_26215,N_26372);
and U29659 (N_29659,N_24735,N_25411);
or U29660 (N_29660,N_25420,N_26571);
and U29661 (N_29661,N_24927,N_26449);
or U29662 (N_29662,N_24866,N_25261);
nand U29663 (N_29663,N_24467,N_24199);
or U29664 (N_29664,N_25238,N_25237);
xor U29665 (N_29665,N_25714,N_24802);
or U29666 (N_29666,N_24846,N_24163);
nand U29667 (N_29667,N_24959,N_25850);
and U29668 (N_29668,N_24237,N_25222);
nand U29669 (N_29669,N_26993,N_24648);
and U29670 (N_29670,N_25615,N_24023);
nand U29671 (N_29671,N_26481,N_26559);
nand U29672 (N_29672,N_26549,N_26631);
and U29673 (N_29673,N_24756,N_26521);
and U29674 (N_29674,N_26037,N_26156);
or U29675 (N_29675,N_26827,N_24757);
nand U29676 (N_29676,N_24609,N_26187);
nand U29677 (N_29677,N_24873,N_25347);
nor U29678 (N_29678,N_24700,N_26970);
nor U29679 (N_29679,N_26616,N_25739);
nand U29680 (N_29680,N_25774,N_24027);
xnor U29681 (N_29681,N_25267,N_24182);
and U29682 (N_29682,N_25814,N_25874);
nand U29683 (N_29683,N_25167,N_24327);
and U29684 (N_29684,N_24288,N_24526);
or U29685 (N_29685,N_25035,N_24960);
nand U29686 (N_29686,N_25811,N_24342);
or U29687 (N_29687,N_26148,N_26374);
and U29688 (N_29688,N_24805,N_26946);
and U29689 (N_29689,N_24229,N_25854);
nand U29690 (N_29690,N_26080,N_25345);
nor U29691 (N_29691,N_24082,N_25951);
xor U29692 (N_29692,N_24347,N_24171);
nor U29693 (N_29693,N_26608,N_26611);
xnor U29694 (N_29694,N_24859,N_25745);
and U29695 (N_29695,N_25590,N_24071);
nand U29696 (N_29696,N_25682,N_25213);
nor U29697 (N_29697,N_24878,N_26802);
or U29698 (N_29698,N_25436,N_25741);
and U29699 (N_29699,N_26252,N_26634);
and U29700 (N_29700,N_24838,N_26722);
nand U29701 (N_29701,N_25771,N_26068);
and U29702 (N_29702,N_24828,N_24736);
nand U29703 (N_29703,N_26577,N_24988);
xor U29704 (N_29704,N_26659,N_25862);
or U29705 (N_29705,N_24419,N_26119);
nor U29706 (N_29706,N_24152,N_25292);
or U29707 (N_29707,N_25056,N_26302);
nor U29708 (N_29708,N_24512,N_24716);
nor U29709 (N_29709,N_26079,N_25508);
nand U29710 (N_29710,N_25613,N_26983);
nor U29711 (N_29711,N_25081,N_26530);
and U29712 (N_29712,N_24360,N_24323);
and U29713 (N_29713,N_26422,N_24834);
or U29714 (N_29714,N_25096,N_24270);
or U29715 (N_29715,N_24985,N_24952);
and U29716 (N_29716,N_25039,N_25564);
and U29717 (N_29717,N_24634,N_26042);
nand U29718 (N_29718,N_25175,N_26456);
nand U29719 (N_29719,N_25216,N_24614);
and U29720 (N_29720,N_24674,N_24182);
nor U29721 (N_29721,N_25367,N_24606);
and U29722 (N_29722,N_25397,N_25794);
or U29723 (N_29723,N_26913,N_24543);
xnor U29724 (N_29724,N_25113,N_25819);
or U29725 (N_29725,N_26384,N_25949);
nand U29726 (N_29726,N_24340,N_24090);
and U29727 (N_29727,N_26058,N_24671);
nor U29728 (N_29728,N_25102,N_25391);
and U29729 (N_29729,N_26847,N_26497);
or U29730 (N_29730,N_26258,N_25555);
nand U29731 (N_29731,N_26433,N_25952);
xnor U29732 (N_29732,N_25629,N_25934);
nor U29733 (N_29733,N_24753,N_24631);
nor U29734 (N_29734,N_24718,N_24950);
or U29735 (N_29735,N_26268,N_25682);
and U29736 (N_29736,N_26136,N_26986);
or U29737 (N_29737,N_26402,N_26742);
or U29738 (N_29738,N_24836,N_26484);
nand U29739 (N_29739,N_26350,N_25315);
nand U29740 (N_29740,N_25740,N_25778);
nand U29741 (N_29741,N_24572,N_24433);
or U29742 (N_29742,N_26620,N_26162);
or U29743 (N_29743,N_25756,N_26745);
xor U29744 (N_29744,N_24964,N_25937);
and U29745 (N_29745,N_24192,N_25927);
nand U29746 (N_29746,N_25477,N_24482);
nand U29747 (N_29747,N_25936,N_26934);
xnor U29748 (N_29748,N_24278,N_26130);
and U29749 (N_29749,N_26919,N_26826);
and U29750 (N_29750,N_25078,N_25149);
nor U29751 (N_29751,N_24266,N_26408);
and U29752 (N_29752,N_26902,N_26522);
nand U29753 (N_29753,N_24073,N_25594);
and U29754 (N_29754,N_25751,N_26760);
nor U29755 (N_29755,N_24459,N_26017);
or U29756 (N_29756,N_25916,N_24667);
nand U29757 (N_29757,N_24596,N_24225);
and U29758 (N_29758,N_25727,N_26992);
and U29759 (N_29759,N_26074,N_25810);
nand U29760 (N_29760,N_24569,N_26801);
and U29761 (N_29761,N_24902,N_26578);
or U29762 (N_29762,N_26960,N_24051);
and U29763 (N_29763,N_24067,N_25248);
nand U29764 (N_29764,N_26760,N_25567);
or U29765 (N_29765,N_25566,N_24552);
or U29766 (N_29766,N_24888,N_26033);
and U29767 (N_29767,N_24934,N_24742);
or U29768 (N_29768,N_24567,N_26836);
xnor U29769 (N_29769,N_25977,N_24350);
nand U29770 (N_29770,N_26037,N_26640);
xor U29771 (N_29771,N_24833,N_26906);
nor U29772 (N_29772,N_26042,N_25011);
nand U29773 (N_29773,N_24237,N_24309);
or U29774 (N_29774,N_26926,N_26427);
nand U29775 (N_29775,N_25378,N_26891);
nand U29776 (N_29776,N_26355,N_25503);
nand U29777 (N_29777,N_26354,N_26530);
nand U29778 (N_29778,N_25487,N_26296);
nand U29779 (N_29779,N_26544,N_24449);
nand U29780 (N_29780,N_25341,N_25905);
nand U29781 (N_29781,N_24596,N_24683);
and U29782 (N_29782,N_25333,N_26005);
nor U29783 (N_29783,N_24428,N_25597);
nor U29784 (N_29784,N_24751,N_25301);
nand U29785 (N_29785,N_25250,N_25807);
and U29786 (N_29786,N_25109,N_25010);
or U29787 (N_29787,N_24059,N_24758);
and U29788 (N_29788,N_26204,N_26804);
nand U29789 (N_29789,N_24090,N_25372);
nor U29790 (N_29790,N_24628,N_26957);
nor U29791 (N_29791,N_25586,N_24083);
and U29792 (N_29792,N_24652,N_25037);
nor U29793 (N_29793,N_26098,N_25522);
nand U29794 (N_29794,N_26196,N_24319);
nand U29795 (N_29795,N_24350,N_26396);
and U29796 (N_29796,N_24716,N_25656);
and U29797 (N_29797,N_24335,N_24637);
or U29798 (N_29798,N_25001,N_26479);
nor U29799 (N_29799,N_25041,N_26637);
nand U29800 (N_29800,N_24713,N_25084);
xnor U29801 (N_29801,N_26245,N_24332);
nand U29802 (N_29802,N_25118,N_24598);
and U29803 (N_29803,N_24777,N_25040);
nor U29804 (N_29804,N_24925,N_25519);
nor U29805 (N_29805,N_26391,N_26651);
nor U29806 (N_29806,N_26680,N_26740);
nor U29807 (N_29807,N_25023,N_26251);
or U29808 (N_29808,N_25182,N_24444);
or U29809 (N_29809,N_25234,N_24077);
and U29810 (N_29810,N_26436,N_25076);
nor U29811 (N_29811,N_26748,N_25998);
nor U29812 (N_29812,N_24195,N_26069);
nor U29813 (N_29813,N_26570,N_26475);
nand U29814 (N_29814,N_26356,N_25277);
nand U29815 (N_29815,N_26171,N_26441);
nor U29816 (N_29816,N_25313,N_26649);
nor U29817 (N_29817,N_26804,N_26892);
and U29818 (N_29818,N_24867,N_26571);
and U29819 (N_29819,N_25266,N_24863);
and U29820 (N_29820,N_25401,N_24849);
or U29821 (N_29821,N_25075,N_24606);
xnor U29822 (N_29822,N_25346,N_24970);
nand U29823 (N_29823,N_25937,N_24167);
xnor U29824 (N_29824,N_26477,N_26280);
nand U29825 (N_29825,N_26007,N_26038);
nand U29826 (N_29826,N_25212,N_24999);
nor U29827 (N_29827,N_26581,N_26802);
nor U29828 (N_29828,N_25321,N_26627);
and U29829 (N_29829,N_24491,N_26773);
nor U29830 (N_29830,N_24160,N_26780);
nor U29831 (N_29831,N_26786,N_24161);
nor U29832 (N_29832,N_25498,N_26722);
or U29833 (N_29833,N_26289,N_25411);
and U29834 (N_29834,N_26335,N_24066);
nand U29835 (N_29835,N_24731,N_26530);
nand U29836 (N_29836,N_26226,N_24550);
nand U29837 (N_29837,N_24783,N_24936);
and U29838 (N_29838,N_26470,N_24500);
xor U29839 (N_29839,N_25280,N_25766);
or U29840 (N_29840,N_25919,N_26355);
and U29841 (N_29841,N_26756,N_25659);
or U29842 (N_29842,N_26147,N_25527);
xnor U29843 (N_29843,N_26027,N_26539);
nor U29844 (N_29844,N_24449,N_25694);
nor U29845 (N_29845,N_25060,N_25102);
and U29846 (N_29846,N_26710,N_25918);
or U29847 (N_29847,N_24281,N_24894);
xnor U29848 (N_29848,N_24427,N_25673);
nor U29849 (N_29849,N_24687,N_25525);
nand U29850 (N_29850,N_26395,N_25726);
and U29851 (N_29851,N_25490,N_25161);
nor U29852 (N_29852,N_26288,N_25793);
xor U29853 (N_29853,N_26427,N_25549);
and U29854 (N_29854,N_24597,N_26659);
xnor U29855 (N_29855,N_25224,N_25545);
nand U29856 (N_29856,N_25688,N_24109);
or U29857 (N_29857,N_25460,N_25944);
or U29858 (N_29858,N_25853,N_26116);
nand U29859 (N_29859,N_25824,N_25140);
and U29860 (N_29860,N_24305,N_26612);
or U29861 (N_29861,N_25046,N_25502);
xnor U29862 (N_29862,N_24110,N_24273);
xor U29863 (N_29863,N_25053,N_25314);
nor U29864 (N_29864,N_24941,N_24563);
or U29865 (N_29865,N_24537,N_26090);
nor U29866 (N_29866,N_24357,N_24512);
nand U29867 (N_29867,N_26804,N_24602);
nor U29868 (N_29868,N_24136,N_26564);
and U29869 (N_29869,N_26465,N_24906);
nor U29870 (N_29870,N_26723,N_26972);
and U29871 (N_29871,N_26692,N_24025);
or U29872 (N_29872,N_25546,N_24964);
nor U29873 (N_29873,N_25650,N_25603);
nand U29874 (N_29874,N_26624,N_26588);
nor U29875 (N_29875,N_26478,N_26838);
or U29876 (N_29876,N_26317,N_25864);
and U29877 (N_29877,N_24406,N_26686);
or U29878 (N_29878,N_26020,N_26412);
or U29879 (N_29879,N_26434,N_25160);
nand U29880 (N_29880,N_24083,N_25821);
and U29881 (N_29881,N_26544,N_24035);
nor U29882 (N_29882,N_24346,N_26763);
or U29883 (N_29883,N_26065,N_24980);
and U29884 (N_29884,N_26346,N_24606);
and U29885 (N_29885,N_25342,N_25154);
nand U29886 (N_29886,N_24466,N_26655);
and U29887 (N_29887,N_24403,N_26210);
and U29888 (N_29888,N_25647,N_26592);
xor U29889 (N_29889,N_26766,N_26027);
or U29890 (N_29890,N_25941,N_24160);
nor U29891 (N_29891,N_24919,N_24580);
nand U29892 (N_29892,N_26108,N_25450);
nand U29893 (N_29893,N_24199,N_25880);
nand U29894 (N_29894,N_24486,N_26539);
and U29895 (N_29895,N_26301,N_24107);
nor U29896 (N_29896,N_24659,N_26674);
and U29897 (N_29897,N_26594,N_24174);
nand U29898 (N_29898,N_26099,N_26013);
and U29899 (N_29899,N_24941,N_25058);
nor U29900 (N_29900,N_24894,N_24988);
nor U29901 (N_29901,N_26338,N_24413);
nor U29902 (N_29902,N_26991,N_26573);
nand U29903 (N_29903,N_24415,N_25907);
and U29904 (N_29904,N_26357,N_25923);
xor U29905 (N_29905,N_26796,N_25830);
or U29906 (N_29906,N_24795,N_25253);
or U29907 (N_29907,N_26462,N_25090);
nand U29908 (N_29908,N_24973,N_24717);
and U29909 (N_29909,N_25552,N_26840);
nand U29910 (N_29910,N_26112,N_25430);
nor U29911 (N_29911,N_25991,N_24389);
nand U29912 (N_29912,N_25243,N_26467);
xnor U29913 (N_29913,N_26765,N_24130);
and U29914 (N_29914,N_25195,N_26171);
or U29915 (N_29915,N_25920,N_26713);
nand U29916 (N_29916,N_25982,N_25302);
nand U29917 (N_29917,N_25676,N_26728);
nand U29918 (N_29918,N_25491,N_25949);
nor U29919 (N_29919,N_25239,N_24548);
nor U29920 (N_29920,N_25919,N_25382);
nand U29921 (N_29921,N_26215,N_24372);
or U29922 (N_29922,N_26205,N_26811);
or U29923 (N_29923,N_25678,N_26624);
or U29924 (N_29924,N_25891,N_26949);
or U29925 (N_29925,N_26972,N_24788);
nor U29926 (N_29926,N_24980,N_24327);
nor U29927 (N_29927,N_25038,N_24689);
nor U29928 (N_29928,N_26705,N_25752);
or U29929 (N_29929,N_25696,N_24509);
xnor U29930 (N_29930,N_24724,N_26634);
or U29931 (N_29931,N_26488,N_25652);
xor U29932 (N_29932,N_25475,N_24810);
and U29933 (N_29933,N_25180,N_26808);
nand U29934 (N_29934,N_25534,N_26366);
and U29935 (N_29935,N_26099,N_24772);
or U29936 (N_29936,N_24773,N_25718);
or U29937 (N_29937,N_25628,N_25352);
or U29938 (N_29938,N_26597,N_25008);
and U29939 (N_29939,N_24664,N_26834);
and U29940 (N_29940,N_26708,N_26682);
xnor U29941 (N_29941,N_25468,N_26391);
nor U29942 (N_29942,N_25393,N_24056);
xnor U29943 (N_29943,N_25743,N_24327);
and U29944 (N_29944,N_26608,N_25298);
or U29945 (N_29945,N_25084,N_25285);
nor U29946 (N_29946,N_24413,N_26333);
nand U29947 (N_29947,N_25506,N_26732);
or U29948 (N_29948,N_24975,N_25912);
xnor U29949 (N_29949,N_25903,N_25734);
or U29950 (N_29950,N_24433,N_24560);
and U29951 (N_29951,N_26302,N_26732);
and U29952 (N_29952,N_25032,N_25200);
or U29953 (N_29953,N_26358,N_26487);
and U29954 (N_29954,N_26710,N_25323);
or U29955 (N_29955,N_25852,N_26571);
xnor U29956 (N_29956,N_24318,N_25218);
or U29957 (N_29957,N_25121,N_26388);
or U29958 (N_29958,N_26936,N_25262);
xor U29959 (N_29959,N_26965,N_25342);
xnor U29960 (N_29960,N_25745,N_25845);
nand U29961 (N_29961,N_25185,N_25434);
or U29962 (N_29962,N_25052,N_24544);
or U29963 (N_29963,N_26876,N_24798);
and U29964 (N_29964,N_24359,N_25680);
nand U29965 (N_29965,N_25692,N_25653);
xor U29966 (N_29966,N_24487,N_26295);
and U29967 (N_29967,N_26450,N_24769);
and U29968 (N_29968,N_25697,N_25520);
nand U29969 (N_29969,N_24342,N_26205);
and U29970 (N_29970,N_26567,N_25607);
nor U29971 (N_29971,N_25084,N_24340);
nand U29972 (N_29972,N_24369,N_26362);
or U29973 (N_29973,N_24127,N_25181);
nor U29974 (N_29974,N_25581,N_24541);
or U29975 (N_29975,N_25098,N_25941);
xor U29976 (N_29976,N_26815,N_26013);
nand U29977 (N_29977,N_25888,N_24175);
nor U29978 (N_29978,N_26173,N_26392);
and U29979 (N_29979,N_24289,N_24043);
nand U29980 (N_29980,N_24990,N_25491);
nand U29981 (N_29981,N_26751,N_26166);
xnor U29982 (N_29982,N_24682,N_25097);
xnor U29983 (N_29983,N_25232,N_25052);
nand U29984 (N_29984,N_24807,N_26849);
or U29985 (N_29985,N_26744,N_26684);
and U29986 (N_29986,N_25299,N_25783);
nand U29987 (N_29987,N_26440,N_25411);
or U29988 (N_29988,N_26771,N_25360);
or U29989 (N_29989,N_24363,N_25793);
and U29990 (N_29990,N_24190,N_26154);
nand U29991 (N_29991,N_24605,N_24981);
or U29992 (N_29992,N_24226,N_26727);
nand U29993 (N_29993,N_25158,N_24994);
or U29994 (N_29994,N_25255,N_26752);
and U29995 (N_29995,N_24574,N_25910);
nor U29996 (N_29996,N_25642,N_24638);
nor U29997 (N_29997,N_24906,N_25353);
or U29998 (N_29998,N_26241,N_26416);
nor U29999 (N_29999,N_25932,N_24219);
xnor UO_0 (O_0,N_28713,N_29463);
nor UO_1 (O_1,N_28609,N_28159);
nand UO_2 (O_2,N_28197,N_29793);
xor UO_3 (O_3,N_28525,N_27538);
xor UO_4 (O_4,N_29116,N_27818);
nor UO_5 (O_5,N_28783,N_29470);
nand UO_6 (O_6,N_29440,N_29069);
or UO_7 (O_7,N_28594,N_28590);
nor UO_8 (O_8,N_27147,N_27105);
nor UO_9 (O_9,N_29500,N_27264);
xnor UO_10 (O_10,N_29811,N_29998);
nand UO_11 (O_11,N_28807,N_27155);
or UO_12 (O_12,N_27111,N_27323);
or UO_13 (O_13,N_29645,N_29469);
nor UO_14 (O_14,N_29297,N_29676);
nand UO_15 (O_15,N_29745,N_27258);
or UO_16 (O_16,N_29573,N_27179);
or UO_17 (O_17,N_29859,N_29395);
nand UO_18 (O_18,N_28795,N_27228);
nor UO_19 (O_19,N_29136,N_29090);
or UO_20 (O_20,N_27613,N_29327);
nor UO_21 (O_21,N_27029,N_29046);
and UO_22 (O_22,N_29163,N_28800);
and UO_23 (O_23,N_29402,N_28926);
nor UO_24 (O_24,N_28799,N_29738);
nand UO_25 (O_25,N_27471,N_29442);
or UO_26 (O_26,N_29369,N_28942);
or UO_27 (O_27,N_29564,N_29436);
or UO_28 (O_28,N_28318,N_27922);
or UO_29 (O_29,N_29729,N_27187);
nor UO_30 (O_30,N_27243,N_28112);
or UO_31 (O_31,N_29814,N_27259);
and UO_32 (O_32,N_27807,N_29822);
and UO_33 (O_33,N_29887,N_29340);
nand UO_34 (O_34,N_27221,N_27123);
nand UO_35 (O_35,N_28405,N_28516);
or UO_36 (O_36,N_28764,N_29108);
nand UO_37 (O_37,N_29909,N_29051);
xnor UO_38 (O_38,N_28135,N_28975);
nor UO_39 (O_39,N_28346,N_28538);
and UO_40 (O_40,N_27495,N_27732);
or UO_41 (O_41,N_27663,N_27509);
or UO_42 (O_42,N_27767,N_27245);
nor UO_43 (O_43,N_27063,N_27300);
nand UO_44 (O_44,N_27059,N_27974);
nand UO_45 (O_45,N_27257,N_29653);
and UO_46 (O_46,N_27330,N_29431);
nor UO_47 (O_47,N_27594,N_27354);
nand UO_48 (O_48,N_29558,N_27592);
nor UO_49 (O_49,N_27771,N_27142);
nand UO_50 (O_50,N_29200,N_28787);
nand UO_51 (O_51,N_27931,N_28261);
and UO_52 (O_52,N_29040,N_29259);
nor UO_53 (O_53,N_29888,N_28130);
xor UO_54 (O_54,N_28736,N_27557);
nand UO_55 (O_55,N_29199,N_28856);
xor UO_56 (O_56,N_28341,N_28133);
and UO_57 (O_57,N_27737,N_27086);
and UO_58 (O_58,N_27348,N_28234);
or UO_59 (O_59,N_28671,N_29527);
nor UO_60 (O_60,N_29902,N_27353);
and UO_61 (O_61,N_27313,N_29457);
and UO_62 (O_62,N_27854,N_29192);
and UO_63 (O_63,N_28232,N_29838);
nand UO_64 (O_64,N_28083,N_29915);
nor UO_65 (O_65,N_29741,N_29430);
xnor UO_66 (O_66,N_29922,N_28064);
nor UO_67 (O_67,N_29854,N_27904);
nand UO_68 (O_68,N_29810,N_27181);
nor UO_69 (O_69,N_28715,N_28763);
or UO_70 (O_70,N_27791,N_29841);
nand UO_71 (O_71,N_28936,N_29740);
xor UO_72 (O_72,N_28499,N_27892);
nand UO_73 (O_73,N_29139,N_29452);
xnor UO_74 (O_74,N_27046,N_28305);
and UO_75 (O_75,N_27388,N_27579);
and UO_76 (O_76,N_27661,N_27335);
nor UO_77 (O_77,N_29592,N_28427);
or UO_78 (O_78,N_28390,N_28802);
xor UO_79 (O_79,N_28769,N_27716);
or UO_80 (O_80,N_29635,N_29026);
or UO_81 (O_81,N_28356,N_29298);
and UO_82 (O_82,N_27829,N_29744);
nand UO_83 (O_83,N_29076,N_27101);
and UO_84 (O_84,N_28729,N_29984);
and UO_85 (O_85,N_28418,N_28812);
or UO_86 (O_86,N_28482,N_27017);
nand UO_87 (O_87,N_27654,N_27697);
nor UO_88 (O_88,N_29765,N_28436);
or UO_89 (O_89,N_29906,N_29794);
nand UO_90 (O_90,N_27902,N_29596);
nor UO_91 (O_91,N_27834,N_29017);
and UO_92 (O_92,N_27433,N_28309);
and UO_93 (O_93,N_29828,N_28208);
nor UO_94 (O_94,N_29386,N_28943);
nor UO_95 (O_95,N_29060,N_29677);
or UO_96 (O_96,N_27048,N_28424);
xnor UO_97 (O_97,N_27239,N_29089);
nand UO_98 (O_98,N_27996,N_27503);
nor UO_99 (O_99,N_27479,N_28473);
or UO_100 (O_100,N_28015,N_29043);
nand UO_101 (O_101,N_28563,N_29987);
or UO_102 (O_102,N_28735,N_29972);
and UO_103 (O_103,N_27207,N_27368);
xnor UO_104 (O_104,N_28697,N_29183);
or UO_105 (O_105,N_27961,N_29346);
or UO_106 (O_106,N_29176,N_29349);
or UO_107 (O_107,N_29388,N_28552);
nor UO_108 (O_108,N_29979,N_28278);
nor UO_109 (O_109,N_28182,N_29003);
nand UO_110 (O_110,N_29492,N_27830);
nand UO_111 (O_111,N_27790,N_29770);
or UO_112 (O_112,N_29570,N_28251);
nor UO_113 (O_113,N_27997,N_27696);
nor UO_114 (O_114,N_28411,N_27513);
and UO_115 (O_115,N_29066,N_27753);
nor UO_116 (O_116,N_27315,N_28878);
nand UO_117 (O_117,N_27943,N_27061);
or UO_118 (O_118,N_29561,N_27911);
and UO_119 (O_119,N_28838,N_29256);
and UO_120 (O_120,N_28545,N_28329);
nand UO_121 (O_121,N_29864,N_27201);
nand UO_122 (O_122,N_28727,N_28958);
and UO_123 (O_123,N_27066,N_29569);
and UO_124 (O_124,N_28254,N_29265);
nand UO_125 (O_125,N_29840,N_28292);
nor UO_126 (O_126,N_28378,N_28521);
nand UO_127 (O_127,N_28326,N_29119);
nand UO_128 (O_128,N_29542,N_28851);
xnor UO_129 (O_129,N_28056,N_28136);
xnor UO_130 (O_130,N_28307,N_27988);
nand UO_131 (O_131,N_28149,N_27390);
and UO_132 (O_132,N_28751,N_28435);
nand UO_133 (O_133,N_27333,N_27395);
nor UO_134 (O_134,N_28080,N_28123);
xor UO_135 (O_135,N_28887,N_29456);
and UO_136 (O_136,N_27377,N_29622);
and UO_137 (O_137,N_27140,N_29184);
xnor UO_138 (O_138,N_28164,N_28191);
nand UO_139 (O_139,N_27777,N_29152);
or UO_140 (O_140,N_29866,N_27837);
nand UO_141 (O_141,N_28919,N_29719);
nor UO_142 (O_142,N_27669,N_27692);
xnor UO_143 (O_143,N_28823,N_29245);
nand UO_144 (O_144,N_28223,N_29555);
or UO_145 (O_145,N_27549,N_27569);
or UO_146 (O_146,N_29524,N_28263);
and UO_147 (O_147,N_28479,N_27003);
xnor UO_148 (O_148,N_29768,N_28820);
or UO_149 (O_149,N_27383,N_29935);
and UO_150 (O_150,N_27516,N_28465);
or UO_151 (O_151,N_28540,N_29389);
xnor UO_152 (O_152,N_29264,N_28839);
or UO_153 (O_153,N_27277,N_27435);
or UO_154 (O_154,N_29313,N_29001);
nor UO_155 (O_155,N_29604,N_28095);
nand UO_156 (O_156,N_29952,N_27720);
nor UO_157 (O_157,N_29280,N_27519);
or UO_158 (O_158,N_28970,N_29113);
and UO_159 (O_159,N_28954,N_28102);
nor UO_160 (O_160,N_28454,N_28432);
and UO_161 (O_161,N_27452,N_29825);
or UO_162 (O_162,N_29379,N_29960);
nand UO_163 (O_163,N_29112,N_27415);
and UO_164 (O_164,N_27189,N_28766);
or UO_165 (O_165,N_29600,N_27560);
or UO_166 (O_166,N_29534,N_29632);
nand UO_167 (O_167,N_27328,N_28833);
nand UO_168 (O_168,N_27664,N_29285);
and UO_169 (O_169,N_28216,N_27907);
nor UO_170 (O_170,N_28573,N_29231);
nand UO_171 (O_171,N_27849,N_29853);
and UO_172 (O_172,N_29048,N_28646);
or UO_173 (O_173,N_27242,N_28669);
and UO_174 (O_174,N_29938,N_27916);
nor UO_175 (O_175,N_28829,N_27143);
nand UO_176 (O_176,N_29077,N_29597);
nand UO_177 (O_177,N_29688,N_27180);
nor UO_178 (O_178,N_28923,N_29757);
nand UO_179 (O_179,N_29631,N_27256);
nand UO_180 (O_180,N_28199,N_29743);
or UO_181 (O_181,N_27392,N_27989);
or UO_182 (O_182,N_27506,N_28925);
and UO_183 (O_183,N_27404,N_27969);
and UO_184 (O_184,N_27623,N_29024);
nand UO_185 (O_185,N_29267,N_27526);
nor UO_186 (O_186,N_27889,N_28630);
nor UO_187 (O_187,N_29144,N_28407);
xnor UO_188 (O_188,N_29595,N_27158);
nand UO_189 (O_189,N_27420,N_29962);
nand UO_190 (O_190,N_29959,N_29512);
or UO_191 (O_191,N_28379,N_28698);
nor UO_192 (O_192,N_27204,N_28895);
or UO_193 (O_193,N_27018,N_28652);
or UO_194 (O_194,N_28181,N_27825);
nor UO_195 (O_195,N_28090,N_27548);
or UO_196 (O_196,N_28816,N_27803);
nand UO_197 (O_197,N_27119,N_27662);
xnor UO_198 (O_198,N_28265,N_29750);
nand UO_199 (O_199,N_29494,N_29879);
nor UO_200 (O_200,N_28998,N_28046);
nor UO_201 (O_201,N_28592,N_27114);
nand UO_202 (O_202,N_28439,N_27026);
nor UO_203 (O_203,N_28018,N_27596);
nand UO_204 (O_204,N_29391,N_27776);
and UO_205 (O_205,N_29449,N_28549);
nor UO_206 (O_206,N_28255,N_27843);
and UO_207 (O_207,N_27608,N_29507);
or UO_208 (O_208,N_27038,N_27067);
or UO_209 (O_209,N_28349,N_28298);
nor UO_210 (O_210,N_29191,N_27770);
nor UO_211 (O_211,N_28249,N_29050);
nand UO_212 (O_212,N_28272,N_28685);
xnor UO_213 (O_213,N_27741,N_28534);
xnor UO_214 (O_214,N_27443,N_28333);
nand UO_215 (O_215,N_28979,N_28917);
or UO_216 (O_216,N_27115,N_27149);
and UO_217 (O_217,N_27480,N_27617);
nor UO_218 (O_218,N_27271,N_27231);
and UO_219 (O_219,N_27612,N_28988);
nor UO_220 (O_220,N_29680,N_29733);
nor UO_221 (O_221,N_27681,N_29846);
and UO_222 (O_222,N_29437,N_27251);
xor UO_223 (O_223,N_29913,N_28423);
and UO_224 (O_224,N_28959,N_27075);
or UO_225 (O_225,N_28012,N_28717);
and UO_226 (O_226,N_28931,N_29746);
nor UO_227 (O_227,N_27319,N_29813);
nand UO_228 (O_228,N_28137,N_27401);
and UO_229 (O_229,N_29889,N_29292);
and UO_230 (O_230,N_28585,N_29704);
nand UO_231 (O_231,N_29455,N_29477);
nand UO_232 (O_232,N_29146,N_28239);
xnor UO_233 (O_233,N_29934,N_29362);
xor UO_234 (O_234,N_28877,N_28648);
and UO_235 (O_235,N_27021,N_29488);
and UO_236 (O_236,N_29637,N_27108);
or UO_237 (O_237,N_29010,N_28033);
nor UO_238 (O_238,N_27650,N_29783);
nor UO_239 (O_239,N_28962,N_29240);
nand UO_240 (O_240,N_29400,N_28148);
and UO_241 (O_241,N_29869,N_27937);
or UO_242 (O_242,N_28376,N_28395);
and UO_243 (O_243,N_28704,N_28675);
nor UO_244 (O_244,N_29634,N_27196);
nand UO_245 (O_245,N_28176,N_29105);
or UO_246 (O_246,N_29749,N_28964);
nand UO_247 (O_247,N_28950,N_28422);
and UO_248 (O_248,N_27938,N_28172);
nand UO_249 (O_249,N_28971,N_29401);
nor UO_250 (O_250,N_27533,N_29279);
or UO_251 (O_251,N_29971,N_28955);
nand UO_252 (O_252,N_27117,N_27894);
or UO_253 (O_253,N_29905,N_27883);
or UO_254 (O_254,N_28062,N_29111);
and UO_255 (O_255,N_28830,N_27651);
nor UO_256 (O_256,N_28093,N_27094);
or UO_257 (O_257,N_28299,N_29826);
or UO_258 (O_258,N_29381,N_27260);
and UO_259 (O_259,N_28290,N_27879);
nand UO_260 (O_260,N_29848,N_27578);
xor UO_261 (O_261,N_27322,N_29304);
nor UO_262 (O_262,N_27727,N_28639);
and UO_263 (O_263,N_28126,N_28242);
nor UO_264 (O_264,N_28616,N_29383);
nor UO_265 (O_265,N_29792,N_29357);
and UO_266 (O_266,N_28118,N_28775);
and UO_267 (O_267,N_28668,N_29608);
or UO_268 (O_268,N_29390,N_28387);
or UO_269 (O_269,N_28899,N_27614);
or UO_270 (O_270,N_27817,N_29038);
or UO_271 (O_271,N_29602,N_27811);
nor UO_272 (O_272,N_29013,N_27908);
nor UO_273 (O_273,N_29617,N_29588);
and UO_274 (O_274,N_28173,N_28900);
and UO_275 (O_275,N_29158,N_27762);
xnor UO_276 (O_276,N_28007,N_29693);
or UO_277 (O_277,N_27972,N_29643);
and UO_278 (O_278,N_28791,N_27287);
nor UO_279 (O_279,N_28940,N_27559);
nand UO_280 (O_280,N_28233,N_29774);
and UO_281 (O_281,N_27097,N_29165);
and UO_282 (O_282,N_27083,N_29258);
nand UO_283 (O_283,N_27006,N_27622);
and UO_284 (O_284,N_27970,N_27437);
nand UO_285 (O_285,N_27919,N_29319);
nand UO_286 (O_286,N_29443,N_29651);
nand UO_287 (O_287,N_27289,N_29718);
and UO_288 (O_288,N_29658,N_27051);
or UO_289 (O_289,N_28099,N_28916);
nand UO_290 (O_290,N_29249,N_29843);
xnor UO_291 (O_291,N_28328,N_29928);
nor UO_292 (O_292,N_29428,N_29343);
nor UO_293 (O_293,N_28313,N_28868);
nand UO_294 (O_294,N_28687,N_29097);
nand UO_295 (O_295,N_29504,N_27504);
or UO_296 (O_296,N_27855,N_28773);
nor UO_297 (O_297,N_29802,N_29659);
nor UO_298 (O_298,N_29098,N_28282);
xor UO_299 (O_299,N_28653,N_28359);
nor UO_300 (O_300,N_29930,N_29877);
nand UO_301 (O_301,N_27358,N_29329);
xnor UO_302 (O_302,N_28588,N_28896);
and UO_303 (O_303,N_29503,N_28336);
nand UO_304 (O_304,N_27165,N_28711);
and UO_305 (O_305,N_28276,N_27840);
nor UO_306 (O_306,N_28984,N_28957);
nand UO_307 (O_307,N_29851,N_29664);
or UO_308 (O_308,N_27831,N_28296);
or UO_309 (O_309,N_27899,N_28973);
nand UO_310 (O_310,N_29065,N_27124);
and UO_311 (O_311,N_27331,N_27652);
nand UO_312 (O_312,N_28300,N_28651);
and UO_313 (O_313,N_28695,N_29241);
and UO_314 (O_314,N_28902,N_28315);
or UO_315 (O_315,N_27958,N_29257);
and UO_316 (O_316,N_27011,N_29876);
and UO_317 (O_317,N_27898,N_29781);
xnor UO_318 (O_318,N_28548,N_27413);
xnor UO_319 (O_319,N_27810,N_28048);
nor UO_320 (O_320,N_27213,N_29845);
and UO_321 (O_321,N_27699,N_28470);
nor UO_322 (O_322,N_28060,N_29506);
and UO_323 (O_323,N_29818,N_29904);
and UO_324 (O_324,N_29226,N_28170);
xor UO_325 (O_325,N_27144,N_28863);
nand UO_326 (O_326,N_29014,N_28391);
xnor UO_327 (O_327,N_29737,N_27601);
and UO_328 (O_328,N_28714,N_27792);
nand UO_329 (O_329,N_29281,N_27477);
or UO_330 (O_330,N_28890,N_29047);
nor UO_331 (O_331,N_27556,N_27379);
nor UO_332 (O_332,N_28385,N_29875);
nor UO_333 (O_333,N_28221,N_29131);
and UO_334 (O_334,N_29263,N_29919);
nor UO_335 (O_335,N_29961,N_27173);
nor UO_336 (O_336,N_27933,N_27303);
or UO_337 (O_337,N_28228,N_27900);
nor UO_338 (O_338,N_29893,N_29762);
or UO_339 (O_339,N_27041,N_29705);
nand UO_340 (O_340,N_28710,N_27740);
xor UO_341 (O_341,N_29018,N_28835);
or UO_342 (O_342,N_27500,N_29352);
nor UO_343 (O_343,N_29006,N_27798);
nand UO_344 (O_344,N_28344,N_29100);
nor UO_345 (O_345,N_29490,N_28758);
and UO_346 (O_346,N_28617,N_27019);
nand UO_347 (O_347,N_28235,N_29661);
or UO_348 (O_348,N_28343,N_28266);
nor UO_349 (O_349,N_29342,N_28415);
and UO_350 (O_350,N_29977,N_27054);
nand UO_351 (O_351,N_28319,N_29268);
and UO_352 (O_352,N_28138,N_27724);
nor UO_353 (O_353,N_28051,N_28458);
nand UO_354 (O_354,N_29434,N_27233);
or UO_355 (O_355,N_29035,N_28485);
or UO_356 (O_356,N_27024,N_29412);
or UO_357 (O_357,N_27921,N_28712);
or UO_358 (O_358,N_29538,N_28096);
nor UO_359 (O_359,N_28495,N_27963);
and UO_360 (O_360,N_27278,N_28103);
xnor UO_361 (O_361,N_27736,N_29374);
xnor UO_362 (O_362,N_28610,N_29880);
xor UO_363 (O_363,N_27658,N_27483);
nand UO_364 (O_364,N_28380,N_29337);
nor UO_365 (O_365,N_27307,N_28157);
nand UO_366 (O_366,N_27215,N_28022);
and UO_367 (O_367,N_27424,N_27926);
and UO_368 (O_368,N_27139,N_29535);
xor UO_369 (O_369,N_29414,N_27308);
nor UO_370 (O_370,N_28185,N_28279);
xor UO_371 (O_371,N_28151,N_28915);
or UO_372 (O_372,N_29416,N_29439);
nand UO_373 (O_373,N_27641,N_28416);
and UO_374 (O_374,N_27905,N_29471);
or UO_375 (O_375,N_27028,N_27229);
nor UO_376 (O_376,N_27530,N_29795);
or UO_377 (O_377,N_27253,N_27202);
or UO_378 (O_378,N_27070,N_29734);
and UO_379 (O_379,N_28969,N_29168);
xor UO_380 (O_380,N_27610,N_27694);
xnor UO_381 (O_381,N_28854,N_28226);
nand UO_382 (O_382,N_27357,N_28094);
nor UO_383 (O_383,N_27248,N_28768);
or UO_384 (O_384,N_28857,N_27138);
xnor UO_385 (O_385,N_28815,N_27891);
nand UO_386 (O_386,N_29916,N_28792);
or UO_387 (O_387,N_29423,N_27396);
nor UO_388 (O_388,N_29944,N_29238);
or UO_389 (O_389,N_27188,N_27940);
xnor UO_390 (O_390,N_29147,N_28660);
xor UO_391 (O_391,N_27064,N_27025);
nand UO_392 (O_392,N_29034,N_29620);
or UO_393 (O_393,N_27567,N_27295);
nor UO_394 (O_394,N_29284,N_27965);
and UO_395 (O_395,N_27174,N_27800);
nand UO_396 (O_396,N_29732,N_27291);
xor UO_397 (O_397,N_29489,N_28035);
or UO_398 (O_398,N_28044,N_29212);
nor UO_399 (O_399,N_28743,N_29206);
or UO_400 (O_400,N_29751,N_27962);
and UO_401 (O_401,N_29260,N_28143);
nor UO_402 (O_402,N_27045,N_27216);
and UO_403 (O_403,N_28338,N_29261);
or UO_404 (O_404,N_27742,N_29326);
or UO_405 (O_405,N_27707,N_29511);
nor UO_406 (O_406,N_27624,N_29912);
or UO_407 (O_407,N_27570,N_29759);
and UO_408 (O_408,N_28734,N_28358);
nor UO_409 (O_409,N_27723,N_29673);
nor UO_410 (O_410,N_29198,N_27555);
nor UO_411 (O_411,N_29126,N_28752);
and UO_412 (O_412,N_27678,N_28201);
nand UO_413 (O_413,N_27448,N_27957);
or UO_414 (O_414,N_29609,N_27869);
nand UO_415 (O_415,N_27376,N_28209);
xor UO_416 (O_416,N_27351,N_29910);
nor UO_417 (O_417,N_29679,N_29099);
xnor UO_418 (O_418,N_29269,N_28446);
nand UO_419 (O_419,N_29755,N_28933);
xor UO_420 (O_420,N_27507,N_29925);
or UO_421 (O_421,N_27850,N_29545);
nand UO_422 (O_422,N_27876,N_28043);
nor UO_423 (O_423,N_28113,N_27620);
and UO_424 (O_424,N_28977,N_29985);
nand UO_425 (O_425,N_29957,N_28566);
or UO_426 (O_426,N_27593,N_28141);
and UO_427 (O_427,N_28991,N_28528);
and UO_428 (O_428,N_27375,N_27721);
nand UO_429 (O_429,N_28939,N_27113);
and UO_430 (O_430,N_29173,N_27468);
or UO_431 (O_431,N_28865,N_29160);
nor UO_432 (O_432,N_27252,N_29418);
nand UO_433 (O_433,N_27691,N_29054);
or UO_434 (O_434,N_29537,N_29502);
and UO_435 (O_435,N_28375,N_27451);
or UO_436 (O_436,N_29501,N_28274);
and UO_437 (O_437,N_28562,N_27730);
and UO_438 (O_438,N_29782,N_28961);
and UO_439 (O_439,N_29235,N_29482);
xnor UO_440 (O_440,N_28597,N_28611);
and UO_441 (O_441,N_28690,N_28809);
or UO_442 (O_442,N_27566,N_29937);
nor UO_443 (O_443,N_29016,N_27896);
nand UO_444 (O_444,N_29367,N_28894);
xnor UO_445 (O_445,N_28072,N_27544);
and UO_446 (O_446,N_27481,N_27217);
or UO_447 (O_447,N_27005,N_28124);
or UO_448 (O_448,N_27668,N_27527);
xor UO_449 (O_449,N_29523,N_27558);
nand UO_450 (O_450,N_29574,N_28455);
nand UO_451 (O_451,N_27634,N_29188);
and UO_452 (O_452,N_29104,N_29368);
nand UO_453 (O_453,N_28230,N_28845);
nand UO_454 (O_454,N_29921,N_29530);
and UO_455 (O_455,N_29899,N_27056);
and UO_456 (O_456,N_27980,N_28819);
nand UO_457 (O_457,N_28510,N_28577);
xnor UO_458 (O_458,N_27112,N_27665);
nor UO_459 (O_459,N_28347,N_29092);
nor UO_460 (O_460,N_29873,N_27102);
xor UO_461 (O_461,N_27604,N_27884);
or UO_462 (O_462,N_29467,N_28881);
nand UO_463 (O_463,N_29674,N_29669);
nor UO_464 (O_464,N_29012,N_27877);
nor UO_465 (O_465,N_27655,N_29638);
nor UO_466 (O_466,N_29178,N_28508);
or UO_467 (O_467,N_28122,N_27214);
and UO_468 (O_468,N_28640,N_28161);
xor UO_469 (O_469,N_28440,N_27983);
or UO_470 (O_470,N_29946,N_27738);
nor UO_471 (O_471,N_29137,N_28335);
and UO_472 (O_472,N_28457,N_28146);
nor UO_473 (O_473,N_27341,N_27247);
nand UO_474 (O_474,N_27946,N_29565);
nand UO_475 (O_475,N_28505,N_28397);
nor UO_476 (O_476,N_29621,N_29509);
and UO_477 (O_477,N_29788,N_28903);
nor UO_478 (O_478,N_29236,N_27903);
nor UO_479 (O_479,N_28175,N_28303);
xnor UO_480 (O_480,N_27960,N_27674);
and UO_481 (O_481,N_27764,N_27979);
nand UO_482 (O_482,N_28659,N_28127);
nor UO_483 (O_483,N_28023,N_29756);
xor UO_484 (O_484,N_29115,N_28901);
nor UO_485 (O_485,N_29692,N_27012);
or UO_486 (O_486,N_29917,N_29195);
nand UO_487 (O_487,N_28091,N_28636);
and UO_488 (O_488,N_27326,N_28568);
nor UO_489 (O_489,N_28488,N_27848);
nor UO_490 (O_490,N_29219,N_27490);
or UO_491 (O_491,N_28623,N_27708);
nor UO_492 (O_492,N_29886,N_29372);
or UO_493 (O_493,N_29308,N_29208);
or UO_494 (O_494,N_29106,N_27999);
or UO_495 (O_495,N_28889,N_29128);
or UO_496 (O_496,N_29626,N_27316);
and UO_497 (O_497,N_29218,N_29143);
or UO_498 (O_498,N_27890,N_27409);
nand UO_499 (O_499,N_29495,N_27702);
or UO_500 (O_500,N_28997,N_27191);
xor UO_501 (O_501,N_28417,N_29836);
nand UO_502 (O_502,N_29358,N_29145);
or UO_503 (O_503,N_28109,N_29045);
or UO_504 (O_504,N_28077,N_28428);
and UO_505 (O_505,N_29769,N_28810);
nand UO_506 (O_506,N_28702,N_29963);
xnor UO_507 (O_507,N_27844,N_28377);
and UO_508 (O_508,N_28657,N_29255);
nor UO_509 (O_509,N_28104,N_27676);
nor UO_510 (O_510,N_27587,N_27643);
and UO_511 (O_511,N_29725,N_29586);
nor UO_512 (O_512,N_28382,N_29712);
or UO_513 (O_513,N_29328,N_29177);
nand UO_514 (O_514,N_29812,N_29064);
xor UO_515 (O_515,N_28321,N_28363);
xnor UO_516 (O_516,N_28403,N_27164);
xor UO_517 (O_517,N_28804,N_29196);
xnor UO_518 (O_518,N_27089,N_28999);
or UO_519 (O_519,N_28207,N_27531);
or UO_520 (O_520,N_29625,N_29323);
or UO_521 (O_521,N_28183,N_28361);
xor UO_522 (O_522,N_28231,N_27129);
or UO_523 (O_523,N_27071,N_27687);
and UO_524 (O_524,N_28317,N_27606);
and UO_525 (O_525,N_29295,N_29666);
nand UO_526 (O_526,N_28345,N_28448);
or UO_527 (O_527,N_28569,N_27910);
or UO_528 (O_528,N_28121,N_28430);
or UO_529 (O_529,N_27363,N_28559);
xnor UO_530 (O_530,N_27126,N_29594);
xnor UO_531 (O_531,N_27182,N_29299);
nand UO_532 (O_532,N_29384,N_27082);
nand UO_533 (O_533,N_29125,N_28813);
and UO_534 (O_534,N_29075,N_28551);
or UO_535 (O_535,N_28425,N_28667);
and UO_536 (O_536,N_28978,N_28946);
and UO_537 (O_537,N_27981,N_27486);
nor UO_538 (O_538,N_28576,N_27246);
nand UO_539 (O_539,N_27915,N_28767);
nor UO_540 (O_540,N_27583,N_27282);
and UO_541 (O_541,N_27197,N_29974);
and UO_542 (O_542,N_28491,N_29239);
nor UO_543 (O_543,N_27301,N_27093);
or UO_544 (O_544,N_29832,N_27867);
nand UO_545 (O_545,N_29403,N_29228);
and UO_546 (O_546,N_29325,N_27540);
and UO_547 (O_547,N_29522,N_28858);
and UO_548 (O_548,N_29011,N_29205);
or UO_549 (O_549,N_28968,N_29052);
nor UO_550 (O_550,N_29084,N_28876);
and UO_551 (O_551,N_28029,N_27534);
or UO_552 (O_552,N_29900,N_27194);
or UO_553 (O_553,N_29031,N_27107);
nand UO_554 (O_554,N_29964,N_28537);
and UO_555 (O_555,N_28184,N_28441);
nand UO_556 (O_556,N_27203,N_29947);
nand UO_557 (O_557,N_28402,N_28213);
nor UO_558 (O_558,N_27380,N_29380);
and UO_559 (O_559,N_28281,N_29275);
nand UO_560 (O_560,N_27865,N_28575);
nand UO_561 (O_561,N_29148,N_29189);
nand UO_562 (O_562,N_29335,N_27945);
nand UO_563 (O_563,N_27552,N_28331);
and UO_564 (O_564,N_27757,N_27036);
nand UO_565 (O_565,N_29703,N_29767);
or UO_566 (O_566,N_27636,N_28108);
xnor UO_567 (O_567,N_27014,N_28620);
xnor UO_568 (O_568,N_28332,N_29465);
or UO_569 (O_569,N_29672,N_28277);
or UO_570 (O_570,N_28088,N_29780);
nand UO_571 (O_571,N_29114,N_27092);
nor UO_572 (O_572,N_27971,N_29800);
or UO_573 (O_573,N_29682,N_28880);
and UO_574 (O_574,N_28987,N_27788);
and UO_575 (O_575,N_27266,N_29531);
or UO_576 (O_576,N_28312,N_28860);
or UO_577 (O_577,N_27190,N_29955);
and UO_578 (O_578,N_27459,N_28066);
and UO_579 (O_579,N_29305,N_29454);
or UO_580 (O_580,N_27756,N_28467);
or UO_581 (O_581,N_29914,N_27484);
and UO_582 (O_582,N_27550,N_29073);
nand UO_583 (O_583,N_27227,N_28512);
nor UO_584 (O_584,N_28747,N_28938);
nand UO_585 (O_585,N_28178,N_29382);
or UO_586 (O_586,N_27947,N_29655);
and UO_587 (O_587,N_29373,N_27386);
and UO_588 (O_588,N_29307,N_28111);
or UO_589 (O_589,N_29486,N_27780);
nand UO_590 (O_590,N_29398,N_29159);
or UO_591 (O_591,N_27514,N_27993);
nor UO_592 (O_592,N_29656,N_28098);
nand UO_593 (O_593,N_28294,N_27049);
nand UO_594 (O_594,N_28392,N_27302);
and UO_595 (O_595,N_27332,N_27603);
or UO_596 (O_596,N_28935,N_27009);
nand UO_597 (O_597,N_29222,N_27185);
nand UO_598 (O_598,N_27501,N_27299);
and UO_599 (O_599,N_28542,N_29243);
nand UO_600 (O_600,N_29493,N_27037);
nand UO_601 (O_601,N_28280,N_29020);
and UO_602 (O_602,N_27078,N_29883);
nor UO_603 (O_603,N_28179,N_27739);
or UO_604 (O_604,N_27728,N_27934);
xnor UO_605 (O_605,N_29994,N_29803);
or UO_606 (O_606,N_27935,N_28606);
nor UO_607 (O_607,N_28250,N_27499);
and UO_608 (O_608,N_28911,N_29474);
nand UO_609 (O_609,N_29197,N_28259);
xnor UO_610 (O_610,N_29533,N_28794);
nand UO_611 (O_611,N_27088,N_27541);
or UO_612 (O_612,N_28709,N_27745);
nand UO_613 (O_613,N_29706,N_28907);
or UO_614 (O_614,N_29577,N_28119);
and UO_615 (O_615,N_27529,N_27498);
or UO_616 (O_616,N_28608,N_29683);
nand UO_617 (O_617,N_29763,N_28666);
or UO_618 (O_618,N_27927,N_27478);
or UO_619 (O_619,N_29487,N_27199);
or UO_620 (O_620,N_27023,N_29172);
nor UO_621 (O_621,N_28401,N_29742);
nand UO_622 (O_622,N_27735,N_27485);
xor UO_623 (O_623,N_29897,N_27536);
or UO_624 (O_624,N_28167,N_27518);
nor UO_625 (O_625,N_29544,N_29378);
nor UO_626 (O_626,N_28069,N_27132);
or UO_627 (O_627,N_28314,N_29234);
nand UO_628 (O_628,N_29923,N_28355);
nand UO_629 (O_629,N_28558,N_28205);
and UO_630 (O_630,N_28850,N_27878);
nor UO_631 (O_631,N_27445,N_29053);
xnor UO_632 (O_632,N_27441,N_27584);
or UO_633 (O_633,N_27367,N_28981);
xor UO_634 (O_634,N_27033,N_27822);
and UO_635 (O_635,N_29995,N_28746);
or UO_636 (O_636,N_28644,N_28982);
nand UO_637 (O_637,N_29435,N_29294);
or UO_638 (O_638,N_27690,N_27421);
xnor UO_639 (O_639,N_29691,N_29778);
nand UO_640 (O_640,N_29083,N_29223);
or UO_641 (O_641,N_27494,N_27492);
nor UO_642 (O_642,N_29220,N_29130);
xor UO_643 (O_643,N_28028,N_28543);
xnor UO_644 (O_644,N_27824,N_27648);
nand UO_645 (O_645,N_28368,N_28774);
xor UO_646 (O_646,N_29546,N_27466);
nand UO_647 (O_647,N_27611,N_27096);
or UO_648 (O_648,N_28909,N_27719);
nand UO_649 (O_649,N_27489,N_28871);
nand UO_650 (O_650,N_27966,N_29697);
nor UO_651 (O_651,N_27659,N_27267);
nand UO_652 (O_652,N_29970,N_27422);
nor UO_653 (O_653,N_29039,N_27660);
nand UO_654 (O_654,N_28930,N_27360);
or UO_655 (O_655,N_29301,N_27975);
nand UO_656 (O_656,N_29118,N_27779);
and UO_657 (O_657,N_28514,N_27647);
xor UO_658 (O_658,N_28948,N_29175);
nand UO_659 (O_659,N_28934,N_29156);
and UO_660 (O_660,N_27475,N_27868);
nor UO_661 (O_661,N_29933,N_28638);
and UO_662 (O_662,N_28914,N_28438);
or UO_663 (O_663,N_27031,N_27842);
nand UO_664 (O_664,N_27637,N_28010);
nand UO_665 (O_665,N_27436,N_29356);
and UO_666 (O_666,N_28744,N_29953);
and UO_667 (O_667,N_27821,N_28381);
nor UO_668 (O_668,N_28092,N_28034);
and UO_669 (O_669,N_29376,N_29607);
and UO_670 (O_670,N_28976,N_28475);
or UO_671 (O_671,N_28990,N_28229);
nand UO_672 (O_672,N_27618,N_29649);
or UO_673 (O_673,N_29686,N_29950);
and UO_674 (O_674,N_27684,N_28486);
nand UO_675 (O_675,N_27909,N_28513);
and UO_676 (O_676,N_27121,N_27683);
or UO_677 (O_677,N_29480,N_29429);
nand UO_678 (O_678,N_28506,N_28031);
or UO_679 (O_679,N_29711,N_27670);
nor UO_680 (O_680,N_28803,N_27688);
and UO_681 (O_681,N_28607,N_29521);
nor UO_682 (O_682,N_28853,N_28445);
nor UO_683 (O_683,N_29041,N_27440);
or UO_684 (O_684,N_27789,N_28582);
and UO_685 (O_685,N_29419,N_29306);
nor UO_686 (O_686,N_27572,N_28536);
nand UO_687 (O_687,N_27772,N_27949);
nor UO_688 (O_688,N_29539,N_27091);
or UO_689 (O_689,N_28586,N_28886);
or UO_690 (O_690,N_29739,N_27802);
nor UO_691 (O_691,N_29107,N_27532);
nor UO_692 (O_692,N_28673,N_28680);
nor UO_693 (O_693,N_28306,N_28596);
nand UO_694 (O_694,N_27973,N_29421);
and UO_695 (O_695,N_27134,N_27157);
and UO_696 (O_696,N_28866,N_27835);
and UO_697 (O_697,N_27152,N_28196);
nor UO_698 (O_698,N_28295,N_29833);
and UO_699 (O_699,N_27359,N_28052);
nand UO_700 (O_700,N_27679,N_29408);
nor UO_701 (O_701,N_27146,N_29473);
xnor UO_702 (O_702,N_27491,N_28760);
nand UO_703 (O_703,N_27077,N_28716);
or UO_704 (O_704,N_28252,N_29807);
and UO_705 (O_705,N_28081,N_28643);
or UO_706 (O_706,N_27167,N_28225);
nor UO_707 (O_707,N_27220,N_27356);
or UO_708 (O_708,N_27978,N_27598);
xnor UO_709 (O_709,N_27939,N_29771);
or UO_710 (O_710,N_27930,N_27766);
nor UO_711 (O_711,N_27057,N_29580);
or UO_712 (O_712,N_27116,N_27497);
and UO_713 (O_713,N_28664,N_29078);
and UO_714 (O_714,N_29815,N_27682);
nor UO_715 (O_715,N_27912,N_29820);
xnor UO_716 (O_716,N_29796,N_27956);
and UO_717 (O_717,N_27044,N_28019);
and UO_718 (O_718,N_28471,N_27310);
nor UO_719 (O_719,N_28656,N_27763);
nor UO_720 (O_720,N_28214,N_29215);
nor UO_721 (O_721,N_29339,N_29566);
and UO_722 (O_722,N_29606,N_28190);
or UO_723 (O_723,N_28904,N_27434);
xnor UO_724 (O_724,N_28433,N_28145);
and UO_725 (O_725,N_29747,N_29290);
or UO_726 (O_726,N_27255,N_28257);
nor UO_727 (O_727,N_27016,N_29568);
nor UO_728 (O_728,N_29056,N_27685);
nand UO_729 (O_729,N_27873,N_28701);
and UO_730 (O_730,N_29484,N_27553);
and UO_731 (O_731,N_27545,N_28187);
or UO_732 (O_732,N_29321,N_28362);
nand UO_733 (O_733,N_28808,N_27212);
nor UO_734 (O_734,N_28614,N_29681);
or UO_735 (O_735,N_27060,N_27465);
or UO_736 (O_736,N_28264,N_27482);
or UO_737 (O_737,N_28826,N_27222);
nand UO_738 (O_738,N_28509,N_28837);
xor UO_739 (O_739,N_29816,N_28604);
or UO_740 (O_740,N_28555,N_27711);
and UO_741 (O_741,N_29660,N_28311);
nor UO_742 (O_742,N_28168,N_29361);
or UO_743 (O_743,N_29274,N_29748);
and UO_744 (O_744,N_29857,N_29248);
nor UO_745 (O_745,N_28101,N_27427);
or UO_746 (O_746,N_28676,N_29969);
nor UO_747 (O_747,N_28945,N_28017);
nand UO_748 (O_748,N_27977,N_29870);
nor UO_749 (O_749,N_27275,N_28393);
xor UO_750 (O_750,N_29121,N_28078);
or UO_751 (O_751,N_29445,N_27917);
and UO_752 (O_752,N_29898,N_27206);
or UO_753 (O_753,N_28539,N_28700);
xor UO_754 (O_754,N_28409,N_28186);
xor UO_755 (O_755,N_29556,N_27773);
nor UO_756 (O_756,N_28322,N_28262);
or UO_757 (O_757,N_27656,N_27680);
and UO_758 (O_758,N_27262,N_28831);
or UO_759 (O_759,N_29855,N_28677);
nor UO_760 (O_760,N_28843,N_27344);
nor UO_761 (O_761,N_27350,N_27369);
nor UO_762 (O_762,N_27847,N_29464);
and UO_763 (O_763,N_27431,N_27671);
nand UO_764 (O_764,N_28632,N_28824);
nor UO_765 (O_765,N_29187,N_29551);
nor UO_766 (O_766,N_28761,N_28983);
or UO_767 (O_767,N_27397,N_29978);
and UO_768 (O_768,N_28785,N_29458);
nand UO_769 (O_769,N_29980,N_27200);
nand UO_770 (O_770,N_28500,N_27796);
nand UO_771 (O_771,N_27525,N_29093);
xor UO_772 (O_772,N_28260,N_29540);
nor UO_773 (O_773,N_27428,N_28348);
nand UO_774 (O_774,N_28692,N_27968);
xor UO_775 (O_775,N_28460,N_29593);
or UO_776 (O_776,N_28699,N_27286);
and UO_777 (O_777,N_28600,N_29668);
nor UO_778 (O_778,N_29310,N_29049);
and UO_779 (O_779,N_27995,N_29976);
nor UO_780 (O_780,N_28166,N_27133);
and UO_781 (O_781,N_28398,N_28507);
xnor UO_782 (O_782,N_27642,N_28974);
nor UO_783 (O_783,N_29140,N_29370);
nor UO_784 (O_784,N_28778,N_29345);
or UO_785 (O_785,N_27469,N_29009);
xor UO_786 (O_786,N_27254,N_29613);
or UO_787 (O_787,N_28053,N_29790);
or UO_788 (O_788,N_29827,N_28086);
nor UO_789 (O_789,N_29646,N_28762);
or UO_790 (O_790,N_27626,N_27370);
nor UO_791 (O_791,N_27321,N_28818);
or UO_792 (O_792,N_27042,N_29572);
nand UO_793 (O_793,N_27474,N_28517);
nor UO_794 (O_794,N_28570,N_27677);
or UO_795 (O_795,N_29409,N_27951);
or UO_796 (O_796,N_27412,N_29232);
nor UO_797 (O_797,N_29117,N_27106);
nor UO_798 (O_798,N_28832,N_28003);
nand UO_799 (O_799,N_27705,N_28463);
nand UO_800 (O_800,N_27460,N_27888);
xor UO_801 (O_801,N_27901,N_27597);
and UO_802 (O_802,N_27885,N_29528);
nand UO_803 (O_803,N_28776,N_28944);
xnor UO_804 (O_804,N_27602,N_29037);
or UO_805 (O_805,N_28797,N_28780);
nand UO_806 (O_806,N_28518,N_27502);
xor UO_807 (O_807,N_27856,N_27959);
nand UO_808 (O_808,N_28068,N_29871);
xnor UO_809 (O_809,N_28089,N_28110);
nand UO_810 (O_810,N_27524,N_28844);
nand UO_811 (O_811,N_27022,N_29966);
nor UO_812 (O_812,N_27419,N_28655);
or UO_813 (O_813,N_28189,N_27585);
nand UO_814 (O_814,N_29541,N_29721);
nand UO_815 (O_815,N_27166,N_27733);
xnor UO_816 (O_816,N_28770,N_27568);
nand UO_817 (O_817,N_29155,N_29169);
nor UO_818 (O_818,N_28030,N_27327);
xor UO_819 (O_819,N_28076,N_27193);
or UO_820 (O_820,N_28248,N_29929);
or UO_821 (O_821,N_28271,N_27081);
nor UO_822 (O_822,N_27932,N_27575);
nor UO_823 (O_823,N_27382,N_28827);
and UO_824 (O_824,N_28293,N_28892);
nor UO_825 (O_825,N_29213,N_29891);
or UO_826 (O_826,N_28932,N_29623);
nand UO_827 (O_827,N_28786,N_28288);
or UO_828 (O_828,N_29324,N_28006);
xnor UO_829 (O_829,N_28725,N_28330);
nor UO_830 (O_830,N_29519,N_29615);
and UO_831 (O_831,N_28073,N_27871);
nand UO_832 (O_832,N_29858,N_29862);
or UO_833 (O_833,N_27058,N_27586);
xnor UO_834 (O_834,N_27457,N_28560);
nor UO_835 (O_835,N_29071,N_28749);
xnor UO_836 (O_836,N_28115,N_28884);
nand UO_837 (O_837,N_28882,N_27364);
nor UO_838 (O_838,N_28000,N_28572);
nor UO_839 (O_839,N_29153,N_27689);
or UO_840 (O_840,N_29699,N_28649);
xor UO_841 (O_841,N_27250,N_27627);
or UO_842 (O_842,N_29791,N_27274);
nand UO_843 (O_843,N_28451,N_29366);
nand UO_844 (O_844,N_28374,N_29941);
or UO_845 (O_845,N_28243,N_29070);
or UO_846 (O_846,N_29134,N_27467);
nor UO_847 (O_847,N_28334,N_28864);
nor UO_848 (O_848,N_29983,N_29293);
and UO_849 (O_849,N_27862,N_29392);
and UO_850 (O_850,N_27628,N_27365);
nand UO_851 (O_851,N_28523,N_29311);
and UO_852 (O_852,N_29135,N_29868);
nand UO_853 (O_853,N_29127,N_28049);
xnor UO_854 (O_854,N_29975,N_29808);
nand UO_855 (O_855,N_29644,N_27456);
nor UO_856 (O_856,N_27758,N_28502);
nor UO_857 (O_857,N_28481,N_27759);
and UO_858 (O_858,N_27942,N_27423);
and UO_859 (O_859,N_27002,N_28434);
or UO_860 (O_860,N_29225,N_29648);
xnor UO_861 (O_861,N_28579,N_28503);
nor UO_862 (O_862,N_27095,N_27893);
nand UO_863 (O_863,N_28765,N_29110);
nand UO_864 (O_864,N_29201,N_28921);
or UO_865 (O_865,N_27007,N_28472);
and UO_866 (O_866,N_28834,N_27393);
or UO_867 (O_867,N_27389,N_29920);
and UO_868 (O_868,N_27405,N_27210);
or UO_869 (O_869,N_29532,N_27551);
and UO_870 (O_870,N_29427,N_29926);
or UO_871 (O_871,N_27408,N_28952);
and UO_872 (O_872,N_27750,N_29927);
nand UO_873 (O_873,N_27128,N_29476);
xor UO_874 (O_874,N_27340,N_28245);
and UO_875 (O_875,N_27136,N_28805);
xnor UO_876 (O_876,N_29731,N_27595);
or UO_877 (O_877,N_29460,N_28841);
nand UO_878 (O_878,N_29852,N_28873);
and UO_879 (O_879,N_28989,N_29027);
nor UO_880 (O_880,N_29518,N_29211);
xor UO_881 (O_881,N_29174,N_29943);
nor UO_882 (O_882,N_28595,N_27131);
nor UO_883 (O_883,N_29417,N_29939);
or UO_884 (O_884,N_29334,N_27281);
nor UO_885 (O_885,N_29185,N_28360);
and UO_886 (O_886,N_27649,N_27381);
nand UO_887 (O_887,N_28163,N_27032);
and UO_888 (O_888,N_29958,N_29360);
nor UO_889 (O_889,N_27985,N_28922);
or UO_890 (O_890,N_28493,N_29954);
nor UO_891 (O_891,N_29582,N_28897);
or UO_892 (O_892,N_28039,N_29717);
nand UO_893 (O_893,N_27845,N_29831);
nor UO_894 (O_894,N_29948,N_29513);
nor UO_895 (O_895,N_29872,N_27591);
or UO_896 (O_896,N_29799,N_28703);
xnor UO_897 (O_897,N_28450,N_27852);
or UO_898 (O_898,N_27887,N_28147);
nand UO_899 (O_899,N_28928,N_28742);
and UO_900 (O_900,N_29730,N_27269);
nand UO_901 (O_901,N_27241,N_27290);
nand UO_902 (O_902,N_27571,N_27135);
and UO_903 (O_903,N_27561,N_28386);
and UO_904 (O_904,N_28840,N_29583);
or UO_905 (O_905,N_28372,N_27069);
and UO_906 (O_906,N_28061,N_27374);
and UO_907 (O_907,N_28951,N_29775);
or UO_908 (O_908,N_28215,N_29124);
nor UO_909 (O_909,N_29193,N_27704);
or UO_910 (O_910,N_29895,N_27053);
or UO_911 (O_911,N_28461,N_29314);
or UO_912 (O_912,N_27874,N_27653);
nor UO_913 (O_913,N_28683,N_27838);
or UO_914 (O_914,N_28162,N_29882);
xor UO_915 (O_915,N_29404,N_27812);
nor UO_916 (O_916,N_29496,N_28211);
or UO_917 (O_917,N_29999,N_28324);
or UO_918 (O_918,N_29315,N_29433);
nand UO_919 (O_919,N_28708,N_28872);
nor UO_920 (O_920,N_27765,N_28100);
nand UO_921 (O_921,N_27755,N_29896);
nor UO_922 (O_922,N_28218,N_27339);
xor UO_923 (O_923,N_29554,N_27870);
and UO_924 (O_924,N_28634,N_28057);
or UO_925 (O_925,N_29590,N_27573);
nand UO_926 (O_926,N_27832,N_28153);
or UO_927 (O_927,N_27463,N_28339);
and UO_928 (O_928,N_27398,N_28637);
nand UO_929 (O_929,N_29141,N_28836);
xnor UO_930 (O_930,N_29186,N_27547);
or UO_931 (O_931,N_27293,N_29685);
and UO_932 (O_932,N_27294,N_27752);
and UO_933 (O_933,N_27564,N_29639);
or UO_934 (O_934,N_29251,N_29413);
and UO_935 (O_935,N_29589,N_29167);
or UO_936 (O_936,N_29365,N_27027);
nor UO_937 (O_937,N_28420,N_29505);
and UO_938 (O_938,N_29426,N_27841);
nand UO_939 (O_939,N_28615,N_29951);
nand UO_940 (O_940,N_27297,N_29063);
nand UO_941 (O_941,N_28670,N_27145);
or UO_942 (O_942,N_27355,N_27314);
xnor UO_943 (O_943,N_27881,N_27387);
and UO_944 (O_944,N_28825,N_29250);
and UO_945 (O_945,N_27998,N_27775);
nor UO_946 (O_946,N_28437,N_28796);
or UO_947 (O_947,N_27864,N_28426);
and UO_948 (O_948,N_27923,N_28273);
nor UO_949 (O_949,N_28464,N_29761);
nor UO_950 (O_950,N_27402,N_27941);
and UO_951 (O_951,N_29085,N_29394);
and UO_952 (O_952,N_28980,N_29931);
and UO_953 (O_953,N_28285,N_28679);
nand UO_954 (O_954,N_28301,N_28009);
or UO_955 (O_955,N_29067,N_29940);
nor UO_956 (O_956,N_29475,N_27455);
nor UO_957 (O_957,N_27230,N_28396);
or UO_958 (O_958,N_28898,N_29667);
nor UO_959 (O_959,N_27161,N_28546);
nand UO_960 (O_960,N_29377,N_29008);
or UO_961 (O_961,N_27192,N_27219);
nor UO_962 (O_962,N_28619,N_29425);
nand UO_963 (O_963,N_29986,N_28532);
nand UO_964 (O_964,N_27808,N_28139);
and UO_965 (O_965,N_28287,N_27713);
and UO_966 (O_966,N_28754,N_28665);
or UO_967 (O_967,N_27866,N_29202);
or UO_968 (O_968,N_28021,N_29459);
nor UO_969 (O_969,N_29591,N_28564);
or UO_970 (O_970,N_27347,N_28414);
and UO_971 (O_971,N_28079,N_28730);
and UO_972 (O_972,N_29997,N_28626);
or UO_973 (O_973,N_28036,N_28489);
nand UO_974 (O_974,N_27714,N_28661);
nand UO_975 (O_975,N_28477,N_29630);
or UO_976 (O_976,N_27337,N_28304);
or UO_977 (O_977,N_27543,N_28227);
and UO_978 (O_978,N_28696,N_28447);
or UO_979 (O_979,N_28027,N_29350);
or UO_980 (O_980,N_28748,N_28498);
nor UO_981 (O_981,N_27235,N_27168);
nor UO_982 (O_982,N_27853,N_28444);
nor UO_983 (O_983,N_29233,N_28553);
and UO_984 (O_984,N_29096,N_28497);
nand UO_985 (O_985,N_27693,N_29341);
xnor UO_986 (O_986,N_28867,N_27342);
nor UO_987 (O_987,N_28781,N_29300);
nor UO_988 (O_988,N_29088,N_27169);
or UO_989 (O_989,N_29081,N_28212);
nand UO_990 (O_990,N_29936,N_29776);
nor UO_991 (O_991,N_29441,N_27546);
xnor UO_992 (O_992,N_27639,N_28504);
and UO_993 (O_993,N_27487,N_29585);
nor UO_994 (O_994,N_27052,N_27918);
nor UO_995 (O_995,N_27698,N_27633);
or UO_996 (O_996,N_27992,N_27913);
nand UO_997 (O_997,N_28759,N_27099);
or UO_998 (O_998,N_29654,N_29633);
or UO_999 (O_999,N_28453,N_29722);
nor UO_1000 (O_1000,N_27391,N_29736);
xor UO_1001 (O_1001,N_27814,N_27700);
or UO_1002 (O_1002,N_27748,N_28645);
xor UO_1003 (O_1003,N_28004,N_28801);
or UO_1004 (O_1004,N_29628,N_28756);
or UO_1005 (O_1005,N_29863,N_29204);
and UO_1006 (O_1006,N_27488,N_29061);
or UO_1007 (O_1007,N_29694,N_28530);
and UO_1008 (O_1008,N_29120,N_27517);
or UO_1009 (O_1009,N_27731,N_29918);
nor UO_1010 (O_1010,N_28733,N_27880);
xnor UO_1011 (O_1011,N_27806,N_27747);
xnor UO_1012 (O_1012,N_29989,N_27872);
nand UO_1013 (O_1013,N_27863,N_27882);
nor UO_1014 (O_1014,N_29805,N_28480);
xnor UO_1015 (O_1015,N_28177,N_29723);
nand UO_1016 (O_1016,N_29945,N_27774);
or UO_1017 (O_1017,N_29221,N_29844);
and UO_1018 (O_1018,N_27013,N_27065);
nand UO_1019 (O_1019,N_28862,N_28599);
nand UO_1020 (O_1020,N_28155,N_29835);
and UO_1021 (O_1021,N_29161,N_28547);
nor UO_1022 (O_1022,N_27406,N_28419);
and UO_1023 (O_1023,N_28745,N_28814);
nor UO_1024 (O_1024,N_27084,N_27444);
nor UO_1025 (O_1025,N_28366,N_29082);
or UO_1026 (O_1026,N_27156,N_29801);
nor UO_1027 (O_1027,N_28237,N_28128);
nand UO_1028 (O_1028,N_27461,N_29839);
and UO_1029 (O_1029,N_27644,N_29773);
or UO_1030 (O_1030,N_29619,N_28494);
nand UO_1031 (O_1031,N_29652,N_27118);
nand UO_1032 (O_1032,N_29216,N_27580);
nor UO_1033 (O_1033,N_27325,N_28247);
nor UO_1034 (O_1034,N_29695,N_27588);
or UO_1035 (O_1035,N_28220,N_27346);
or UO_1036 (O_1036,N_28684,N_27991);
or UO_1037 (O_1037,N_27263,N_28750);
xnor UO_1038 (O_1038,N_28399,N_29446);
and UO_1039 (O_1039,N_29059,N_29624);
nand UO_1040 (O_1040,N_29303,N_28487);
nor UO_1041 (O_1041,N_27362,N_27125);
nand UO_1042 (O_1042,N_27343,N_29214);
nand UO_1043 (O_1043,N_28621,N_28050);
or UO_1044 (O_1044,N_27819,N_29272);
xor UO_1045 (O_1045,N_28678,N_29080);
and UO_1046 (O_1046,N_29150,N_28996);
xnor UO_1047 (O_1047,N_27528,N_28140);
or UO_1048 (O_1048,N_29779,N_29266);
nor UO_1049 (O_1049,N_28847,N_27240);
nor UO_1050 (O_1050,N_29347,N_29567);
nand UO_1051 (O_1051,N_29354,N_27635);
nor UO_1052 (O_1052,N_28258,N_27760);
nor UO_1053 (O_1053,N_29702,N_27725);
xor UO_1054 (O_1054,N_27860,N_28065);
or UO_1055 (O_1055,N_27280,N_28650);
nand UO_1056 (O_1056,N_27781,N_27283);
and UO_1057 (O_1057,N_28412,N_27666);
or UO_1058 (O_1058,N_28584,N_29129);
nor UO_1059 (O_1059,N_29453,N_29371);
xnor UO_1060 (O_1060,N_29363,N_28811);
nor UO_1061 (O_1061,N_29415,N_29696);
or UO_1062 (O_1062,N_28688,N_29499);
nor UO_1063 (O_1063,N_27110,N_29277);
nand UO_1064 (O_1064,N_27417,N_27607);
and UO_1065 (O_1065,N_29847,N_27520);
nand UO_1066 (O_1066,N_29698,N_29033);
nor UO_1067 (O_1067,N_29510,N_27329);
nand UO_1068 (O_1068,N_28674,N_29684);
nand UO_1069 (O_1069,N_28132,N_27630);
nor UO_1070 (O_1070,N_27616,N_29406);
and UO_1071 (O_1071,N_27349,N_29021);
and UO_1072 (O_1072,N_27265,N_27447);
xnor UO_1073 (O_1073,N_27726,N_28026);
xnor UO_1074 (O_1074,N_28152,N_29576);
nor UO_1075 (O_1075,N_28323,N_28635);
nand UO_1076 (O_1076,N_28353,N_29498);
and UO_1077 (O_1077,N_28483,N_28589);
and UO_1078 (O_1078,N_27249,N_28720);
nor UO_1079 (O_1079,N_29675,N_27450);
xor UO_1080 (O_1080,N_28995,N_27268);
or UO_1081 (O_1081,N_29091,N_27195);
or UO_1082 (O_1082,N_29605,N_28384);
and UO_1083 (O_1083,N_29320,N_28097);
nor UO_1084 (O_1084,N_28757,N_27505);
nand UO_1085 (O_1085,N_29466,N_27787);
and UO_1086 (O_1086,N_27120,N_27914);
and UO_1087 (O_1087,N_28662,N_27673);
or UO_1088 (O_1088,N_29316,N_27924);
and UO_1089 (O_1089,N_28910,N_28370);
nor UO_1090 (O_1090,N_29993,N_29094);
nand UO_1091 (O_1091,N_28256,N_28556);
or UO_1092 (O_1092,N_28055,N_28144);
or UO_1093 (O_1093,N_29559,N_28924);
or UO_1094 (O_1094,N_27218,N_27015);
and UO_1095 (O_1095,N_29516,N_28642);
and UO_1096 (O_1096,N_28920,N_29547);
and UO_1097 (O_1097,N_27846,N_27234);
nand UO_1098 (O_1098,N_28874,N_27906);
or UO_1099 (O_1099,N_29557,N_27170);
or UO_1100 (O_1100,N_27743,N_28478);
nand UO_1101 (O_1101,N_28937,N_28107);
and UO_1102 (O_1102,N_29806,N_29701);
xnor UO_1103 (O_1103,N_28654,N_27799);
and UO_1104 (O_1104,N_28106,N_28120);
nand UO_1105 (O_1105,N_28024,N_28268);
xor UO_1106 (O_1106,N_29000,N_27508);
nor UO_1107 (O_1107,N_27055,N_27833);
nor UO_1108 (O_1108,N_29525,N_27010);
and UO_1109 (O_1109,N_27712,N_27619);
nand UO_1110 (O_1110,N_28531,N_28005);
nor UO_1111 (O_1111,N_28949,N_27839);
and UO_1112 (O_1112,N_28721,N_27537);
nand UO_1113 (O_1113,N_29375,N_29996);
nor UO_1114 (O_1114,N_29562,N_29662);
nor UO_1115 (O_1115,N_29636,N_28413);
or UO_1116 (O_1116,N_27122,N_28732);
or UO_1117 (O_1117,N_27625,N_27305);
xnor UO_1118 (O_1118,N_28722,N_27950);
or UO_1119 (O_1119,N_29042,N_28484);
or UO_1120 (O_1120,N_29690,N_27542);
nor UO_1121 (O_1121,N_27826,N_29028);
nor UO_1122 (O_1122,N_29834,N_29397);
nand UO_1123 (O_1123,N_28219,N_28966);
and UO_1124 (O_1124,N_28798,N_28842);
nor UO_1125 (O_1125,N_28682,N_29407);
nor UO_1126 (O_1126,N_27172,N_27279);
or UO_1127 (O_1127,N_29764,N_28142);
nand UO_1128 (O_1128,N_29317,N_29276);
or UO_1129 (O_1129,N_28535,N_28574);
and UO_1130 (O_1130,N_27198,N_29149);
and UO_1131 (O_1131,N_27224,N_27072);
nand UO_1132 (O_1132,N_29728,N_29973);
and UO_1133 (O_1133,N_27801,N_28156);
nand UO_1134 (O_1134,N_28171,N_28116);
nor UO_1135 (O_1135,N_28658,N_28204);
nand UO_1136 (O_1136,N_28605,N_29289);
nor UO_1137 (O_1137,N_27418,N_27886);
or UO_1138 (O_1138,N_27778,N_28501);
or UO_1139 (O_1139,N_29309,N_27675);
nand UO_1140 (O_1140,N_27897,N_29162);
or UO_1141 (O_1141,N_27967,N_27554);
or UO_1142 (O_1142,N_28105,N_28206);
and UO_1143 (O_1143,N_28821,N_27394);
and UO_1144 (O_1144,N_28075,N_29678);
or UO_1145 (O_1145,N_29968,N_28476);
and UO_1146 (O_1146,N_28627,N_28001);
xnor UO_1147 (O_1147,N_28160,N_28628);
nor UO_1148 (O_1148,N_29603,N_27836);
nor UO_1149 (O_1149,N_29179,N_28963);
and UO_1150 (O_1150,N_27384,N_27709);
xnor UO_1151 (O_1151,N_28406,N_28601);
nand UO_1152 (O_1152,N_27288,N_28550);
nand UO_1153 (O_1153,N_29288,N_27521);
xor UO_1154 (O_1154,N_29629,N_29019);
or UO_1155 (O_1155,N_27646,N_27074);
nand UO_1156 (O_1156,N_28325,N_28443);
nor UO_1157 (O_1157,N_28195,N_27425);
nand UO_1158 (O_1158,N_29157,N_27209);
and UO_1159 (O_1159,N_29478,N_28337);
and UO_1160 (O_1160,N_27920,N_28625);
nor UO_1161 (O_1161,N_27030,N_28404);
nor UO_1162 (O_1162,N_29612,N_27470);
and UO_1163 (O_1163,N_29715,N_27851);
nor UO_1164 (O_1164,N_27827,N_28992);
xor UO_1165 (O_1165,N_27309,N_28849);
nand UO_1166 (O_1166,N_29550,N_27523);
and UO_1167 (O_1167,N_29727,N_29282);
nor UO_1168 (O_1168,N_27510,N_29351);
or UO_1169 (O_1169,N_29752,N_29894);
nand UO_1170 (O_1170,N_28275,N_29967);
and UO_1171 (O_1171,N_28011,N_28738);
and UO_1172 (O_1172,N_27710,N_29312);
xnor UO_1173 (O_1173,N_29584,N_28002);
nor UO_1174 (O_1174,N_27784,N_28777);
and UO_1175 (O_1175,N_29514,N_28782);
and UO_1176 (O_1176,N_29344,N_27324);
or UO_1177 (O_1177,N_29641,N_27177);
or UO_1178 (O_1178,N_27040,N_28373);
nand UO_1179 (O_1179,N_27338,N_27320);
and UO_1180 (O_1180,N_27087,N_28354);
and UO_1181 (O_1181,N_27925,N_28117);
or UO_1182 (O_1182,N_29903,N_29244);
xor UO_1183 (O_1183,N_29708,N_28071);
or UO_1184 (O_1184,N_27104,N_28918);
nor UO_1185 (O_1185,N_29472,N_28883);
or UO_1186 (O_1186,N_28352,N_27782);
nand UO_1187 (O_1187,N_28554,N_29348);
xor UO_1188 (O_1188,N_27414,N_27273);
nand UO_1189 (O_1189,N_29004,N_28074);
or UO_1190 (O_1190,N_27432,N_28705);
and UO_1191 (O_1191,N_29025,N_27043);
nand UO_1192 (O_1192,N_29181,N_29142);
xnor UO_1193 (O_1193,N_28037,N_28134);
nor UO_1194 (O_1194,N_29599,N_27211);
nand UO_1195 (O_1195,N_28452,N_29444);
or UO_1196 (O_1196,N_29491,N_28519);
and UO_1197 (O_1197,N_29022,N_29787);
xnor UO_1198 (O_1198,N_28681,N_28193);
nand UO_1199 (O_1199,N_28286,N_27047);
nand UO_1200 (O_1200,N_28192,N_27020);
nor UO_1201 (O_1201,N_27987,N_29670);
or UO_1202 (O_1202,N_29029,N_27236);
and UO_1203 (O_1203,N_27645,N_29884);
nand UO_1204 (O_1204,N_27148,N_28875);
or UO_1205 (O_1205,N_27859,N_27621);
nor UO_1206 (O_1206,N_27449,N_27496);
and UO_1207 (O_1207,N_27318,N_29055);
xnor UO_1208 (O_1208,N_28772,N_29821);
xor UO_1209 (O_1209,N_27751,N_28041);
nand UO_1210 (O_1210,N_28994,N_29058);
nor UO_1211 (O_1211,N_29789,N_28686);
nand UO_1212 (O_1212,N_27238,N_29229);
nor UO_1213 (O_1213,N_28316,N_29336);
or UO_1214 (O_1214,N_27098,N_28158);
nand UO_1215 (O_1215,N_29246,N_29296);
xnor UO_1216 (O_1216,N_29552,N_27631);
nand UO_1217 (O_1217,N_29447,N_27577);
nand UO_1218 (O_1218,N_29515,N_27100);
or UO_1219 (O_1219,N_29908,N_29860);
nor UO_1220 (O_1220,N_29901,N_28131);
nand UO_1221 (O_1221,N_29536,N_29411);
or UO_1222 (O_1222,N_29581,N_27244);
nand UO_1223 (O_1223,N_29057,N_28310);
and UO_1224 (O_1224,N_29209,N_29422);
xnor UO_1225 (O_1225,N_27372,N_28217);
or UO_1226 (O_1226,N_27403,N_28731);
nor UO_1227 (O_1227,N_27718,N_28200);
and UO_1228 (O_1228,N_29663,N_29074);
or UO_1229 (O_1229,N_29647,N_29874);
and UO_1230 (O_1230,N_27823,N_27539);
xnor UO_1231 (O_1231,N_27261,N_28828);
and UO_1232 (O_1232,N_27729,N_27336);
nand UO_1233 (O_1233,N_28706,N_27439);
nor UO_1234 (O_1234,N_27184,N_27276);
or UO_1235 (O_1235,N_29758,N_29079);
or UO_1236 (O_1236,N_29990,N_28612);
or UO_1237 (O_1237,N_27473,N_29575);
or UO_1238 (O_1238,N_27034,N_29735);
or UO_1239 (O_1239,N_29353,N_27462);
nor UO_1240 (O_1240,N_29032,N_29123);
nor UO_1241 (O_1241,N_28522,N_29164);
and UO_1242 (O_1242,N_29405,N_27183);
and UO_1243 (O_1243,N_29151,N_27783);
nor UO_1244 (O_1244,N_28408,N_29270);
or UO_1245 (O_1245,N_27001,N_29036);
and UO_1246 (O_1246,N_27695,N_28456);
or UO_1247 (O_1247,N_29777,N_27004);
nand UO_1248 (O_1248,N_29956,N_29044);
or UO_1249 (O_1249,N_28779,N_27430);
nand UO_1250 (O_1250,N_28269,N_27141);
or UO_1251 (O_1251,N_28741,N_29109);
nand UO_1252 (O_1252,N_27109,N_28598);
or UO_1253 (O_1253,N_27150,N_29007);
nand UO_1254 (O_1254,N_29689,N_28474);
nor UO_1255 (O_1255,N_28388,N_29424);
or UO_1256 (O_1256,N_28965,N_29154);
or UO_1257 (O_1257,N_28580,N_28082);
nor UO_1258 (O_1258,N_27175,N_27599);
nor UO_1259 (O_1259,N_28449,N_28350);
nor UO_1260 (O_1260,N_27954,N_29571);
xor UO_1261 (O_1261,N_27162,N_28042);
nand UO_1262 (O_1262,N_28986,N_28855);
nand UO_1263 (O_1263,N_28793,N_28085);
xor UO_1264 (O_1264,N_29210,N_27600);
and UO_1265 (O_1265,N_28369,N_29687);
and UO_1266 (O_1266,N_27226,N_29062);
or UO_1267 (O_1267,N_29396,N_27638);
or UO_1268 (O_1268,N_27493,N_27312);
nand UO_1269 (O_1269,N_27990,N_27875);
nand UO_1270 (O_1270,N_29924,N_27062);
and UO_1271 (O_1271,N_28410,N_27426);
and UO_1272 (O_1272,N_28340,N_28879);
nand UO_1273 (O_1273,N_27127,N_29578);
nor UO_1274 (O_1274,N_27232,N_27944);
nor UO_1275 (O_1275,N_27964,N_29322);
or UO_1276 (O_1276,N_27385,N_29122);
or UO_1277 (O_1277,N_29287,N_27154);
xnor UO_1278 (O_1278,N_28059,N_29804);
nor UO_1279 (O_1279,N_28308,N_29330);
nand UO_1280 (O_1280,N_28527,N_27039);
and UO_1281 (O_1281,N_29760,N_28070);
nand UO_1282 (O_1282,N_28067,N_27178);
nand UO_1283 (O_1283,N_29942,N_27797);
or UO_1284 (O_1284,N_28342,N_29483);
xor UO_1285 (O_1285,N_29023,N_28737);
xor UO_1286 (O_1286,N_29230,N_28240);
nor UO_1287 (O_1287,N_29823,N_27512);
or UO_1288 (O_1288,N_29171,N_27657);
and UO_1289 (O_1289,N_29965,N_28581);
nor UO_1290 (O_1290,N_27458,N_29549);
nor UO_1291 (O_1291,N_29797,N_27749);
xnor UO_1292 (O_1292,N_27769,N_29911);
xnor UO_1293 (O_1293,N_28270,N_27090);
and UO_1294 (O_1294,N_28544,N_28693);
and UO_1295 (O_1295,N_27085,N_28058);
or UO_1296 (O_1296,N_29461,N_28253);
and UO_1297 (O_1297,N_27785,N_27137);
nor UO_1298 (O_1298,N_27955,N_27590);
or UO_1299 (O_1299,N_28492,N_27399);
and UO_1300 (O_1300,N_27813,N_29224);
nor UO_1301 (O_1301,N_28008,N_27130);
or UO_1302 (O_1302,N_27296,N_28587);
and UO_1303 (O_1303,N_28613,N_28913);
or UO_1304 (O_1304,N_27317,N_28817);
nand UO_1305 (O_1305,N_29949,N_28755);
nand UO_1306 (O_1306,N_29798,N_28154);
and UO_1307 (O_1307,N_28174,N_29850);
or UO_1308 (O_1308,N_27828,N_29720);
nand UO_1309 (O_1309,N_28846,N_27407);
and UO_1310 (O_1310,N_29611,N_29587);
and UO_1311 (O_1311,N_29772,N_27565);
and UO_1312 (O_1312,N_29448,N_29650);
nor UO_1313 (O_1313,N_29332,N_29291);
nor UO_1314 (O_1314,N_27816,N_28941);
and UO_1315 (O_1315,N_27411,N_27976);
nor UO_1316 (O_1316,N_27416,N_29410);
and UO_1317 (O_1317,N_28602,N_29166);
xnor UO_1318 (O_1318,N_27366,N_28165);
and UO_1319 (O_1319,N_27171,N_29207);
nand UO_1320 (O_1320,N_28267,N_29817);
and UO_1321 (O_1321,N_27272,N_29203);
nor UO_1322 (O_1322,N_29982,N_27073);
nand UO_1323 (O_1323,N_29992,N_28020);
and UO_1324 (O_1324,N_27667,N_28947);
nor UO_1325 (O_1325,N_29627,N_28180);
and UO_1326 (O_1326,N_29830,N_28956);
nor UO_1327 (O_1327,N_29553,N_28806);
and UO_1328 (O_1328,N_28014,N_28515);
xnor UO_1329 (O_1329,N_27511,N_29724);
and UO_1330 (O_1330,N_27080,N_28631);
and UO_1331 (O_1331,N_28431,N_27223);
and UO_1332 (O_1332,N_29138,N_28740);
nand UO_1333 (O_1333,N_27270,N_27361);
nand UO_1334 (O_1334,N_28198,N_29359);
nand UO_1335 (O_1335,N_27744,N_29420);
or UO_1336 (O_1336,N_29247,N_27858);
nand UO_1337 (O_1337,N_28869,N_29861);
nand UO_1338 (O_1338,N_29087,N_29331);
and UO_1339 (O_1339,N_28953,N_28520);
nand UO_1340 (O_1340,N_27581,N_27163);
nor UO_1341 (O_1341,N_29601,N_29753);
nor UO_1342 (O_1342,N_27334,N_29981);
or UO_1343 (O_1343,N_29842,N_28084);
nor UO_1344 (O_1344,N_27672,N_27754);
nand UO_1345 (O_1345,N_28054,N_28726);
and UO_1346 (O_1346,N_28583,N_28442);
nor UO_1347 (O_1347,N_27795,N_27982);
or UO_1348 (O_1348,N_27371,N_27050);
and UO_1349 (O_1349,N_27562,N_29640);
and UO_1350 (O_1350,N_27345,N_29133);
nand UO_1351 (O_1351,N_28371,N_29526);
or UO_1352 (O_1352,N_28169,N_29355);
or UO_1353 (O_1353,N_28985,N_27563);
and UO_1354 (O_1354,N_29278,N_29182);
nor UO_1355 (O_1355,N_29338,N_28429);
or UO_1356 (O_1356,N_27454,N_27820);
or UO_1357 (O_1357,N_29809,N_28906);
xor UO_1358 (O_1358,N_29399,N_28327);
nor UO_1359 (O_1359,N_29318,N_29892);
or UO_1360 (O_1360,N_27442,N_28960);
or UO_1361 (O_1361,N_29766,N_29103);
nor UO_1362 (O_1362,N_28789,N_28578);
and UO_1363 (O_1363,N_29227,N_29302);
and UO_1364 (O_1364,N_29438,N_29068);
nand UO_1365 (O_1365,N_27574,N_29462);
xnor UO_1366 (O_1366,N_28462,N_29543);
or UO_1367 (O_1367,N_28557,N_27160);
nor UO_1368 (O_1368,N_27632,N_28222);
or UO_1369 (O_1369,N_28241,N_29907);
xnor UO_1370 (O_1370,N_27589,N_28210);
or UO_1371 (O_1371,N_28529,N_28739);
nor UO_1372 (O_1372,N_28469,N_27640);
and UO_1373 (O_1373,N_28790,N_29878);
and UO_1374 (O_1374,N_28784,N_28238);
or UO_1375 (O_1375,N_28045,N_28567);
xnor UO_1376 (O_1376,N_28289,N_28848);
or UO_1377 (O_1377,N_28905,N_27515);
or UO_1378 (O_1378,N_28150,N_28244);
xnor UO_1379 (O_1379,N_27809,N_28365);
nand UO_1380 (O_1380,N_29785,N_28490);
or UO_1381 (O_1381,N_27068,N_27429);
nor UO_1382 (O_1382,N_29286,N_28561);
nor UO_1383 (O_1383,N_29132,N_27629);
nand UO_1384 (O_1384,N_29824,N_28753);
nand UO_1385 (O_1385,N_28893,N_28929);
nand UO_1386 (O_1386,N_29642,N_28694);
or UO_1387 (O_1387,N_29598,N_27186);
nor UO_1388 (O_1388,N_29217,N_29579);
xor UO_1389 (O_1389,N_27734,N_27576);
and UO_1390 (O_1390,N_28302,N_27535);
and UO_1391 (O_1391,N_29194,N_28624);
and UO_1392 (O_1392,N_27076,N_29101);
nand UO_1393 (O_1393,N_28524,N_27008);
nor UO_1394 (O_1394,N_29849,N_27000);
and UO_1395 (O_1395,N_28389,N_28641);
nor UO_1396 (O_1396,N_28633,N_28723);
or UO_1397 (O_1397,N_29754,N_28511);
nand UO_1398 (O_1398,N_29710,N_28291);
and UO_1399 (O_1399,N_28888,N_28047);
and UO_1400 (O_1400,N_27715,N_27298);
xnor UO_1401 (O_1401,N_27176,N_28040);
or UO_1402 (O_1402,N_27857,N_27928);
or UO_1403 (O_1403,N_28663,N_29497);
nor UO_1404 (O_1404,N_28861,N_28852);
nor UO_1405 (O_1405,N_28728,N_29508);
or UO_1406 (O_1406,N_28013,N_27952);
and UO_1407 (O_1407,N_27035,N_29726);
or UO_1408 (O_1408,N_29700,N_29015);
and UO_1409 (O_1409,N_28114,N_29005);
nand UO_1410 (O_1410,N_28591,N_29784);
xor UO_1411 (O_1411,N_27410,N_28236);
nand UO_1412 (O_1412,N_27717,N_28647);
nand UO_1413 (O_1413,N_28284,N_27476);
nand UO_1414 (O_1414,N_27805,N_28032);
xnor UO_1415 (O_1415,N_28533,N_29881);
and UO_1416 (O_1416,N_29387,N_29273);
or UO_1417 (O_1417,N_28367,N_28565);
nor UO_1418 (O_1418,N_27861,N_29856);
nand UO_1419 (O_1419,N_28038,N_28459);
nor UO_1420 (O_1420,N_28870,N_29610);
or UO_1421 (O_1421,N_27103,N_29829);
nand UO_1422 (O_1422,N_28788,N_27786);
xnor UO_1423 (O_1423,N_29529,N_27582);
and UO_1424 (O_1424,N_27208,N_27615);
nand UO_1425 (O_1425,N_27400,N_29548);
nor UO_1426 (O_1426,N_28087,N_28025);
and UO_1427 (O_1427,N_29242,N_29560);
and UO_1428 (O_1428,N_28885,N_28394);
xor UO_1429 (O_1429,N_29252,N_27761);
or UO_1430 (O_1430,N_27609,N_27986);
nand UO_1431 (O_1431,N_29885,N_29671);
and UO_1432 (O_1432,N_29707,N_28859);
and UO_1433 (O_1433,N_27722,N_28891);
or UO_1434 (O_1434,N_29614,N_28283);
or UO_1435 (O_1435,N_29385,N_28629);
or UO_1436 (O_1436,N_29451,N_29709);
xnor UO_1437 (O_1437,N_28541,N_28689);
and UO_1438 (O_1438,N_29716,N_29237);
nand UO_1439 (O_1439,N_28618,N_27205);
or UO_1440 (O_1440,N_28912,N_28972);
and UO_1441 (O_1441,N_27936,N_29481);
and UO_1442 (O_1442,N_28822,N_29714);
and UO_1443 (O_1443,N_27815,N_28718);
nor UO_1444 (O_1444,N_28129,N_27793);
nand UO_1445 (O_1445,N_27794,N_29253);
or UO_1446 (O_1446,N_28707,N_27284);
and UO_1447 (O_1447,N_29520,N_29988);
and UO_1448 (O_1448,N_28593,N_29190);
nor UO_1449 (O_1449,N_28691,N_27306);
xor UO_1450 (O_1450,N_29517,N_29865);
and UO_1451 (O_1451,N_29271,N_27746);
or UO_1452 (O_1452,N_27311,N_28202);
nand UO_1453 (O_1453,N_29819,N_27706);
nor UO_1454 (O_1454,N_27453,N_28421);
or UO_1455 (O_1455,N_27472,N_28603);
or UO_1456 (O_1456,N_28383,N_28400);
or UO_1457 (O_1457,N_28246,N_29468);
nor UO_1458 (O_1458,N_27446,N_27352);
or UO_1459 (O_1459,N_29095,N_28719);
and UO_1460 (O_1460,N_29283,N_29563);
nor UO_1461 (O_1461,N_27522,N_28468);
nand UO_1462 (O_1462,N_28297,N_28993);
nor UO_1463 (O_1463,N_27378,N_29072);
nor UO_1464 (O_1464,N_29890,N_28016);
nand UO_1465 (O_1465,N_28357,N_27237);
and UO_1466 (O_1466,N_27153,N_28194);
and UO_1467 (O_1467,N_27159,N_28351);
nor UO_1468 (O_1468,N_27701,N_28224);
or UO_1469 (O_1469,N_27605,N_29102);
nor UO_1470 (O_1470,N_27703,N_29932);
nor UO_1471 (O_1471,N_28724,N_29485);
and UO_1472 (O_1472,N_29479,N_28672);
or UO_1473 (O_1473,N_29030,N_27292);
and UO_1474 (O_1474,N_28125,N_27895);
nand UO_1475 (O_1475,N_29450,N_29254);
nor UO_1476 (O_1476,N_27768,N_28526);
nand UO_1477 (O_1477,N_27984,N_29867);
and UO_1478 (O_1478,N_29713,N_29665);
nand UO_1479 (O_1479,N_29086,N_28622);
and UO_1480 (O_1480,N_28908,N_29364);
nor UO_1481 (O_1481,N_27225,N_29333);
nor UO_1482 (O_1482,N_27438,N_27373);
nor UO_1483 (O_1483,N_27804,N_28063);
and UO_1484 (O_1484,N_29657,N_27285);
and UO_1485 (O_1485,N_28967,N_29170);
xor UO_1486 (O_1486,N_28771,N_29393);
xnor UO_1487 (O_1487,N_27994,N_29262);
and UO_1488 (O_1488,N_28927,N_27079);
nor UO_1489 (O_1489,N_27953,N_28203);
and UO_1490 (O_1490,N_27948,N_29786);
nor UO_1491 (O_1491,N_27151,N_29180);
nor UO_1492 (O_1492,N_28188,N_29618);
nand UO_1493 (O_1493,N_29837,N_29991);
and UO_1494 (O_1494,N_27686,N_27929);
or UO_1495 (O_1495,N_29616,N_28496);
and UO_1496 (O_1496,N_28571,N_29002);
nor UO_1497 (O_1497,N_28364,N_28320);
nor UO_1498 (O_1498,N_29432,N_27464);
xor UO_1499 (O_1499,N_28466,N_27304);
nand UO_1500 (O_1500,N_28167,N_28281);
nor UO_1501 (O_1501,N_29557,N_27304);
or UO_1502 (O_1502,N_27541,N_27018);
nand UO_1503 (O_1503,N_28377,N_28787);
nor UO_1504 (O_1504,N_29415,N_29896);
or UO_1505 (O_1505,N_27009,N_27055);
nand UO_1506 (O_1506,N_27364,N_29923);
or UO_1507 (O_1507,N_28973,N_27627);
and UO_1508 (O_1508,N_27132,N_28407);
nor UO_1509 (O_1509,N_29058,N_28689);
nand UO_1510 (O_1510,N_27822,N_27009);
or UO_1511 (O_1511,N_28890,N_28170);
nor UO_1512 (O_1512,N_27059,N_29258);
nor UO_1513 (O_1513,N_28874,N_28186);
nand UO_1514 (O_1514,N_29145,N_28281);
xnor UO_1515 (O_1515,N_27193,N_28243);
and UO_1516 (O_1516,N_29976,N_27517);
nor UO_1517 (O_1517,N_29816,N_27117);
and UO_1518 (O_1518,N_28208,N_28974);
and UO_1519 (O_1519,N_29869,N_27400);
nor UO_1520 (O_1520,N_29329,N_29113);
or UO_1521 (O_1521,N_28842,N_29555);
nor UO_1522 (O_1522,N_27450,N_29017);
or UO_1523 (O_1523,N_27800,N_28689);
nor UO_1524 (O_1524,N_29637,N_29302);
or UO_1525 (O_1525,N_29324,N_28843);
and UO_1526 (O_1526,N_28688,N_29103);
nand UO_1527 (O_1527,N_28767,N_27224);
nor UO_1528 (O_1528,N_28565,N_28911);
nor UO_1529 (O_1529,N_27194,N_27703);
and UO_1530 (O_1530,N_28759,N_28961);
nor UO_1531 (O_1531,N_29692,N_29162);
xnor UO_1532 (O_1532,N_27179,N_28757);
or UO_1533 (O_1533,N_28872,N_27570);
or UO_1534 (O_1534,N_29262,N_28004);
nand UO_1535 (O_1535,N_29935,N_27807);
or UO_1536 (O_1536,N_28944,N_27484);
nand UO_1537 (O_1537,N_28172,N_29789);
and UO_1538 (O_1538,N_27623,N_27352);
nand UO_1539 (O_1539,N_28142,N_28544);
or UO_1540 (O_1540,N_27092,N_29794);
nand UO_1541 (O_1541,N_28161,N_29079);
nor UO_1542 (O_1542,N_29569,N_29476);
nor UO_1543 (O_1543,N_28356,N_29671);
and UO_1544 (O_1544,N_27497,N_27928);
nor UO_1545 (O_1545,N_29428,N_28102);
and UO_1546 (O_1546,N_27183,N_27128);
nor UO_1547 (O_1547,N_29127,N_29316);
and UO_1548 (O_1548,N_29149,N_28601);
and UO_1549 (O_1549,N_28086,N_28927);
and UO_1550 (O_1550,N_28983,N_29545);
nor UO_1551 (O_1551,N_28800,N_28642);
nand UO_1552 (O_1552,N_27594,N_29241);
and UO_1553 (O_1553,N_27971,N_29873);
and UO_1554 (O_1554,N_27856,N_27401);
nand UO_1555 (O_1555,N_29021,N_28698);
nor UO_1556 (O_1556,N_28918,N_28422);
or UO_1557 (O_1557,N_28457,N_29130);
and UO_1558 (O_1558,N_28514,N_28342);
nand UO_1559 (O_1559,N_28059,N_29628);
xnor UO_1560 (O_1560,N_29964,N_28062);
and UO_1561 (O_1561,N_28665,N_28450);
nand UO_1562 (O_1562,N_29347,N_29284);
nand UO_1563 (O_1563,N_27540,N_27534);
xnor UO_1564 (O_1564,N_28211,N_28245);
and UO_1565 (O_1565,N_28695,N_29003);
and UO_1566 (O_1566,N_27956,N_28842);
nand UO_1567 (O_1567,N_28322,N_28392);
nand UO_1568 (O_1568,N_28092,N_28864);
nand UO_1569 (O_1569,N_28909,N_27515);
xor UO_1570 (O_1570,N_28305,N_29801);
nand UO_1571 (O_1571,N_28417,N_29324);
or UO_1572 (O_1572,N_29713,N_28950);
nand UO_1573 (O_1573,N_28015,N_28558);
and UO_1574 (O_1574,N_28740,N_27860);
nand UO_1575 (O_1575,N_27980,N_28429);
nor UO_1576 (O_1576,N_27883,N_29637);
xor UO_1577 (O_1577,N_29916,N_29579);
nor UO_1578 (O_1578,N_29360,N_27210);
nand UO_1579 (O_1579,N_27861,N_28352);
nor UO_1580 (O_1580,N_27951,N_27300);
or UO_1581 (O_1581,N_28420,N_28383);
xor UO_1582 (O_1582,N_29053,N_29601);
and UO_1583 (O_1583,N_28660,N_28820);
or UO_1584 (O_1584,N_27565,N_29685);
or UO_1585 (O_1585,N_29078,N_28933);
nor UO_1586 (O_1586,N_28967,N_29150);
nand UO_1587 (O_1587,N_28196,N_28468);
and UO_1588 (O_1588,N_28632,N_27329);
and UO_1589 (O_1589,N_27341,N_29821);
or UO_1590 (O_1590,N_28566,N_29994);
or UO_1591 (O_1591,N_27149,N_28389);
xnor UO_1592 (O_1592,N_29142,N_28086);
nand UO_1593 (O_1593,N_28166,N_29573);
nor UO_1594 (O_1594,N_29958,N_28579);
and UO_1595 (O_1595,N_28911,N_27447);
or UO_1596 (O_1596,N_28225,N_29537);
nor UO_1597 (O_1597,N_29232,N_27058);
or UO_1598 (O_1598,N_28493,N_27486);
nand UO_1599 (O_1599,N_27192,N_28002);
and UO_1600 (O_1600,N_28930,N_29792);
xnor UO_1601 (O_1601,N_27381,N_28941);
nor UO_1602 (O_1602,N_29641,N_27214);
and UO_1603 (O_1603,N_27832,N_29090);
nor UO_1604 (O_1604,N_29413,N_27995);
or UO_1605 (O_1605,N_29090,N_28834);
and UO_1606 (O_1606,N_28355,N_29152);
and UO_1607 (O_1607,N_29092,N_27943);
or UO_1608 (O_1608,N_27911,N_29207);
and UO_1609 (O_1609,N_28072,N_28998);
and UO_1610 (O_1610,N_28103,N_28514);
nor UO_1611 (O_1611,N_29755,N_28017);
nand UO_1612 (O_1612,N_29405,N_27036);
nand UO_1613 (O_1613,N_27727,N_28708);
nor UO_1614 (O_1614,N_29762,N_28407);
xor UO_1615 (O_1615,N_29341,N_28360);
nand UO_1616 (O_1616,N_28849,N_27113);
nor UO_1617 (O_1617,N_29745,N_29948);
and UO_1618 (O_1618,N_27136,N_27138);
or UO_1619 (O_1619,N_27091,N_27124);
nor UO_1620 (O_1620,N_27735,N_27070);
and UO_1621 (O_1621,N_28751,N_29493);
xor UO_1622 (O_1622,N_27309,N_28518);
or UO_1623 (O_1623,N_29855,N_29275);
nand UO_1624 (O_1624,N_28629,N_27161);
and UO_1625 (O_1625,N_28790,N_27996);
or UO_1626 (O_1626,N_28059,N_27861);
nand UO_1627 (O_1627,N_29612,N_27332);
nor UO_1628 (O_1628,N_27825,N_28942);
nor UO_1629 (O_1629,N_27350,N_27079);
nand UO_1630 (O_1630,N_28219,N_27056);
nor UO_1631 (O_1631,N_29886,N_28197);
or UO_1632 (O_1632,N_28772,N_27007);
xnor UO_1633 (O_1633,N_27690,N_27408);
nor UO_1634 (O_1634,N_28771,N_29197);
and UO_1635 (O_1635,N_29523,N_28440);
or UO_1636 (O_1636,N_28518,N_27473);
nor UO_1637 (O_1637,N_28405,N_27515);
and UO_1638 (O_1638,N_29055,N_28170);
nor UO_1639 (O_1639,N_29302,N_27217);
or UO_1640 (O_1640,N_28646,N_28311);
nor UO_1641 (O_1641,N_28162,N_27004);
or UO_1642 (O_1642,N_28779,N_29748);
and UO_1643 (O_1643,N_27525,N_29291);
or UO_1644 (O_1644,N_28790,N_29715);
and UO_1645 (O_1645,N_29232,N_28153);
or UO_1646 (O_1646,N_27403,N_28177);
or UO_1647 (O_1647,N_29063,N_27766);
nor UO_1648 (O_1648,N_29205,N_27946);
nand UO_1649 (O_1649,N_27817,N_29355);
nand UO_1650 (O_1650,N_29982,N_27735);
nand UO_1651 (O_1651,N_29625,N_29858);
nand UO_1652 (O_1652,N_29143,N_27576);
or UO_1653 (O_1653,N_29249,N_29817);
nor UO_1654 (O_1654,N_29167,N_28968);
nor UO_1655 (O_1655,N_28426,N_29101);
xor UO_1656 (O_1656,N_28553,N_28897);
nand UO_1657 (O_1657,N_27823,N_29158);
nor UO_1658 (O_1658,N_28580,N_29828);
and UO_1659 (O_1659,N_29154,N_29368);
or UO_1660 (O_1660,N_27101,N_29560);
and UO_1661 (O_1661,N_29402,N_27205);
or UO_1662 (O_1662,N_28866,N_27109);
and UO_1663 (O_1663,N_27992,N_27625);
nand UO_1664 (O_1664,N_27515,N_27355);
nor UO_1665 (O_1665,N_28969,N_29462);
or UO_1666 (O_1666,N_27144,N_29084);
nand UO_1667 (O_1667,N_27741,N_28996);
nand UO_1668 (O_1668,N_27305,N_27863);
and UO_1669 (O_1669,N_27916,N_27641);
xor UO_1670 (O_1670,N_29265,N_28234);
nor UO_1671 (O_1671,N_28044,N_28271);
nand UO_1672 (O_1672,N_28382,N_28652);
and UO_1673 (O_1673,N_29947,N_28484);
or UO_1674 (O_1674,N_29826,N_28579);
and UO_1675 (O_1675,N_28696,N_29439);
and UO_1676 (O_1676,N_28619,N_28393);
xnor UO_1677 (O_1677,N_27999,N_27851);
or UO_1678 (O_1678,N_28883,N_28639);
nor UO_1679 (O_1679,N_29275,N_28492);
or UO_1680 (O_1680,N_29889,N_29865);
nand UO_1681 (O_1681,N_27051,N_27927);
or UO_1682 (O_1682,N_28615,N_28752);
xor UO_1683 (O_1683,N_29584,N_28174);
and UO_1684 (O_1684,N_28430,N_29176);
xor UO_1685 (O_1685,N_29114,N_28811);
nand UO_1686 (O_1686,N_27197,N_28218);
nand UO_1687 (O_1687,N_28197,N_28668);
and UO_1688 (O_1688,N_28169,N_28597);
or UO_1689 (O_1689,N_29082,N_29739);
or UO_1690 (O_1690,N_28461,N_28466);
nand UO_1691 (O_1691,N_29166,N_28348);
or UO_1692 (O_1692,N_29895,N_27308);
nand UO_1693 (O_1693,N_27665,N_27163);
nand UO_1694 (O_1694,N_28459,N_28191);
or UO_1695 (O_1695,N_29364,N_28268);
nor UO_1696 (O_1696,N_27334,N_29950);
nand UO_1697 (O_1697,N_28821,N_28593);
xnor UO_1698 (O_1698,N_29384,N_29194);
nand UO_1699 (O_1699,N_29076,N_29140);
and UO_1700 (O_1700,N_28060,N_29209);
and UO_1701 (O_1701,N_27743,N_29183);
nor UO_1702 (O_1702,N_27775,N_28580);
nor UO_1703 (O_1703,N_29169,N_27535);
and UO_1704 (O_1704,N_27691,N_28626);
nor UO_1705 (O_1705,N_27456,N_27290);
nand UO_1706 (O_1706,N_27858,N_27992);
and UO_1707 (O_1707,N_28351,N_28849);
nor UO_1708 (O_1708,N_29787,N_27227);
nor UO_1709 (O_1709,N_29236,N_29365);
or UO_1710 (O_1710,N_29262,N_28539);
xnor UO_1711 (O_1711,N_27670,N_27303);
nor UO_1712 (O_1712,N_28588,N_28052);
xnor UO_1713 (O_1713,N_29098,N_29253);
and UO_1714 (O_1714,N_28564,N_29720);
and UO_1715 (O_1715,N_29625,N_29525);
xor UO_1716 (O_1716,N_28051,N_29793);
nor UO_1717 (O_1717,N_29712,N_28683);
or UO_1718 (O_1718,N_27628,N_28338);
or UO_1719 (O_1719,N_28345,N_28867);
or UO_1720 (O_1720,N_28344,N_28355);
xor UO_1721 (O_1721,N_28598,N_29095);
nand UO_1722 (O_1722,N_27708,N_29467);
nand UO_1723 (O_1723,N_28553,N_27642);
nand UO_1724 (O_1724,N_29903,N_29715);
nand UO_1725 (O_1725,N_29674,N_29722);
and UO_1726 (O_1726,N_27065,N_28933);
nand UO_1727 (O_1727,N_29009,N_29603);
and UO_1728 (O_1728,N_27334,N_29130);
nand UO_1729 (O_1729,N_28896,N_29262);
or UO_1730 (O_1730,N_27769,N_28958);
nand UO_1731 (O_1731,N_28159,N_27140);
or UO_1732 (O_1732,N_27621,N_27181);
or UO_1733 (O_1733,N_28725,N_28556);
nor UO_1734 (O_1734,N_29126,N_27784);
nand UO_1735 (O_1735,N_27313,N_28336);
nor UO_1736 (O_1736,N_27388,N_29332);
and UO_1737 (O_1737,N_27671,N_27969);
or UO_1738 (O_1738,N_29620,N_29087);
and UO_1739 (O_1739,N_27460,N_27383);
or UO_1740 (O_1740,N_29036,N_27378);
xor UO_1741 (O_1741,N_27942,N_29655);
and UO_1742 (O_1742,N_27041,N_27237);
or UO_1743 (O_1743,N_29170,N_27397);
and UO_1744 (O_1744,N_27332,N_29525);
or UO_1745 (O_1745,N_29666,N_27935);
and UO_1746 (O_1746,N_29413,N_29526);
or UO_1747 (O_1747,N_28060,N_29707);
nor UO_1748 (O_1748,N_28100,N_28428);
nand UO_1749 (O_1749,N_28709,N_29763);
nor UO_1750 (O_1750,N_29375,N_28216);
nand UO_1751 (O_1751,N_27138,N_27731);
or UO_1752 (O_1752,N_28794,N_29100);
nand UO_1753 (O_1753,N_27169,N_29472);
nand UO_1754 (O_1754,N_28677,N_29610);
nand UO_1755 (O_1755,N_29180,N_27749);
and UO_1756 (O_1756,N_29322,N_29541);
or UO_1757 (O_1757,N_28745,N_27127);
or UO_1758 (O_1758,N_29300,N_27470);
or UO_1759 (O_1759,N_27390,N_29219);
nor UO_1760 (O_1760,N_27609,N_27249);
xor UO_1761 (O_1761,N_29466,N_29157);
nand UO_1762 (O_1762,N_27922,N_27306);
and UO_1763 (O_1763,N_28401,N_28784);
nand UO_1764 (O_1764,N_27824,N_29319);
and UO_1765 (O_1765,N_29839,N_29047);
and UO_1766 (O_1766,N_28031,N_28859);
and UO_1767 (O_1767,N_29713,N_29542);
nand UO_1768 (O_1768,N_27837,N_29255);
and UO_1769 (O_1769,N_27313,N_27634);
or UO_1770 (O_1770,N_29410,N_27342);
or UO_1771 (O_1771,N_28293,N_28830);
and UO_1772 (O_1772,N_27257,N_28756);
and UO_1773 (O_1773,N_29786,N_29935);
nand UO_1774 (O_1774,N_28699,N_27519);
xnor UO_1775 (O_1775,N_28784,N_27475);
and UO_1776 (O_1776,N_28518,N_27914);
or UO_1777 (O_1777,N_28487,N_29819);
xnor UO_1778 (O_1778,N_28258,N_28755);
and UO_1779 (O_1779,N_28072,N_27453);
and UO_1780 (O_1780,N_28023,N_29054);
or UO_1781 (O_1781,N_29272,N_27909);
xnor UO_1782 (O_1782,N_27904,N_29052);
nor UO_1783 (O_1783,N_27321,N_27150);
nor UO_1784 (O_1784,N_27151,N_29219);
xnor UO_1785 (O_1785,N_27570,N_28947);
and UO_1786 (O_1786,N_29607,N_29222);
or UO_1787 (O_1787,N_29481,N_28855);
or UO_1788 (O_1788,N_29853,N_28881);
or UO_1789 (O_1789,N_27010,N_28870);
or UO_1790 (O_1790,N_27879,N_27692);
nor UO_1791 (O_1791,N_27855,N_29591);
nand UO_1792 (O_1792,N_28962,N_29832);
and UO_1793 (O_1793,N_28941,N_27736);
nand UO_1794 (O_1794,N_28197,N_27804);
or UO_1795 (O_1795,N_29019,N_28431);
nor UO_1796 (O_1796,N_28567,N_27760);
nand UO_1797 (O_1797,N_27495,N_29214);
nor UO_1798 (O_1798,N_27239,N_28216);
and UO_1799 (O_1799,N_28110,N_28725);
nand UO_1800 (O_1800,N_28607,N_29822);
and UO_1801 (O_1801,N_28366,N_27127);
and UO_1802 (O_1802,N_28171,N_27889);
and UO_1803 (O_1803,N_27035,N_29281);
nor UO_1804 (O_1804,N_29266,N_28355);
nor UO_1805 (O_1805,N_28580,N_27834);
nor UO_1806 (O_1806,N_28487,N_28746);
nand UO_1807 (O_1807,N_29684,N_28257);
or UO_1808 (O_1808,N_27985,N_28501);
nand UO_1809 (O_1809,N_29668,N_29959);
or UO_1810 (O_1810,N_29910,N_28091);
and UO_1811 (O_1811,N_29103,N_27133);
xor UO_1812 (O_1812,N_28521,N_27444);
nor UO_1813 (O_1813,N_29963,N_28742);
nand UO_1814 (O_1814,N_27204,N_27895);
nand UO_1815 (O_1815,N_27464,N_29567);
nor UO_1816 (O_1816,N_28550,N_29117);
nand UO_1817 (O_1817,N_28914,N_29934);
and UO_1818 (O_1818,N_28889,N_28430);
nand UO_1819 (O_1819,N_29653,N_29316);
and UO_1820 (O_1820,N_28811,N_27266);
nand UO_1821 (O_1821,N_29892,N_28719);
or UO_1822 (O_1822,N_29729,N_29789);
or UO_1823 (O_1823,N_28324,N_28648);
nand UO_1824 (O_1824,N_27507,N_29232);
or UO_1825 (O_1825,N_29541,N_28970);
nand UO_1826 (O_1826,N_29256,N_29297);
nor UO_1827 (O_1827,N_27672,N_29124);
xor UO_1828 (O_1828,N_27992,N_28379);
nand UO_1829 (O_1829,N_27391,N_29418);
nor UO_1830 (O_1830,N_29572,N_29676);
nand UO_1831 (O_1831,N_27986,N_29745);
xor UO_1832 (O_1832,N_29418,N_27138);
and UO_1833 (O_1833,N_27015,N_29530);
and UO_1834 (O_1834,N_28125,N_28139);
or UO_1835 (O_1835,N_29700,N_28684);
and UO_1836 (O_1836,N_28783,N_29605);
nor UO_1837 (O_1837,N_28629,N_29207);
or UO_1838 (O_1838,N_29346,N_27848);
nand UO_1839 (O_1839,N_28648,N_29339);
and UO_1840 (O_1840,N_28305,N_29489);
and UO_1841 (O_1841,N_29076,N_29787);
nor UO_1842 (O_1842,N_28836,N_29481);
xor UO_1843 (O_1843,N_27192,N_29722);
or UO_1844 (O_1844,N_29337,N_29237);
nand UO_1845 (O_1845,N_27843,N_27026);
nand UO_1846 (O_1846,N_27128,N_27524);
nand UO_1847 (O_1847,N_29679,N_28656);
nand UO_1848 (O_1848,N_29816,N_27412);
nor UO_1849 (O_1849,N_28322,N_27782);
or UO_1850 (O_1850,N_28116,N_29902);
nand UO_1851 (O_1851,N_27664,N_28998);
and UO_1852 (O_1852,N_28781,N_29970);
nand UO_1853 (O_1853,N_28977,N_29777);
nor UO_1854 (O_1854,N_28716,N_27738);
nand UO_1855 (O_1855,N_28161,N_27597);
or UO_1856 (O_1856,N_29446,N_28494);
nor UO_1857 (O_1857,N_29778,N_27799);
xor UO_1858 (O_1858,N_29787,N_28281);
nor UO_1859 (O_1859,N_28355,N_27834);
xnor UO_1860 (O_1860,N_27056,N_29994);
nand UO_1861 (O_1861,N_27347,N_28641);
or UO_1862 (O_1862,N_29732,N_28137);
nor UO_1863 (O_1863,N_28725,N_29444);
or UO_1864 (O_1864,N_28248,N_27917);
and UO_1865 (O_1865,N_28799,N_29585);
or UO_1866 (O_1866,N_27558,N_29285);
nand UO_1867 (O_1867,N_29622,N_28340);
or UO_1868 (O_1868,N_29867,N_29086);
nand UO_1869 (O_1869,N_28740,N_29854);
nor UO_1870 (O_1870,N_28223,N_29932);
and UO_1871 (O_1871,N_28387,N_29273);
or UO_1872 (O_1872,N_27148,N_27662);
nand UO_1873 (O_1873,N_29068,N_29995);
nand UO_1874 (O_1874,N_27700,N_28231);
nor UO_1875 (O_1875,N_28067,N_27847);
nand UO_1876 (O_1876,N_28525,N_27343);
or UO_1877 (O_1877,N_29884,N_27007);
and UO_1878 (O_1878,N_28064,N_29815);
and UO_1879 (O_1879,N_28108,N_28187);
and UO_1880 (O_1880,N_28366,N_28424);
or UO_1881 (O_1881,N_28305,N_29707);
and UO_1882 (O_1882,N_29141,N_27863);
xnor UO_1883 (O_1883,N_27383,N_28639);
and UO_1884 (O_1884,N_29073,N_29999);
nand UO_1885 (O_1885,N_27060,N_27258);
nand UO_1886 (O_1886,N_27244,N_27895);
or UO_1887 (O_1887,N_27475,N_27404);
and UO_1888 (O_1888,N_27336,N_27558);
or UO_1889 (O_1889,N_27392,N_29552);
nor UO_1890 (O_1890,N_27207,N_29128);
and UO_1891 (O_1891,N_29737,N_28883);
or UO_1892 (O_1892,N_27199,N_29212);
nor UO_1893 (O_1893,N_28724,N_29440);
nand UO_1894 (O_1894,N_28493,N_27614);
and UO_1895 (O_1895,N_29670,N_28856);
nand UO_1896 (O_1896,N_29865,N_28041);
xor UO_1897 (O_1897,N_27588,N_27680);
or UO_1898 (O_1898,N_28856,N_29242);
nor UO_1899 (O_1899,N_29171,N_28976);
nor UO_1900 (O_1900,N_28325,N_27706);
nor UO_1901 (O_1901,N_29193,N_28123);
and UO_1902 (O_1902,N_27227,N_29391);
or UO_1903 (O_1903,N_27093,N_28760);
nor UO_1904 (O_1904,N_27704,N_28525);
or UO_1905 (O_1905,N_27124,N_29848);
or UO_1906 (O_1906,N_29041,N_29880);
nand UO_1907 (O_1907,N_28250,N_27520);
nor UO_1908 (O_1908,N_27297,N_29564);
nand UO_1909 (O_1909,N_27370,N_29950);
nand UO_1910 (O_1910,N_28584,N_29537);
and UO_1911 (O_1911,N_28144,N_29449);
nand UO_1912 (O_1912,N_27062,N_28956);
nor UO_1913 (O_1913,N_27532,N_29206);
nand UO_1914 (O_1914,N_28167,N_27991);
nand UO_1915 (O_1915,N_29791,N_29889);
or UO_1916 (O_1916,N_29657,N_27827);
or UO_1917 (O_1917,N_27883,N_28075);
or UO_1918 (O_1918,N_27135,N_29746);
nand UO_1919 (O_1919,N_27838,N_29731);
xnor UO_1920 (O_1920,N_27905,N_28540);
nor UO_1921 (O_1921,N_28360,N_29211);
nand UO_1922 (O_1922,N_27274,N_28376);
and UO_1923 (O_1923,N_29187,N_28703);
nor UO_1924 (O_1924,N_27143,N_28594);
nor UO_1925 (O_1925,N_29073,N_29223);
or UO_1926 (O_1926,N_29415,N_29215);
nand UO_1927 (O_1927,N_27312,N_27100);
nand UO_1928 (O_1928,N_29536,N_29565);
or UO_1929 (O_1929,N_27625,N_29162);
nand UO_1930 (O_1930,N_28346,N_28292);
nor UO_1931 (O_1931,N_27494,N_28365);
xnor UO_1932 (O_1932,N_29333,N_27823);
nor UO_1933 (O_1933,N_29986,N_27658);
and UO_1934 (O_1934,N_28536,N_29758);
and UO_1935 (O_1935,N_29855,N_29414);
or UO_1936 (O_1936,N_27113,N_27852);
nand UO_1937 (O_1937,N_27954,N_28260);
nor UO_1938 (O_1938,N_27779,N_28435);
nor UO_1939 (O_1939,N_27840,N_28443);
nand UO_1940 (O_1940,N_28539,N_28264);
nand UO_1941 (O_1941,N_27553,N_29787);
nand UO_1942 (O_1942,N_27922,N_28498);
nor UO_1943 (O_1943,N_27191,N_28371);
nor UO_1944 (O_1944,N_29106,N_27339);
xor UO_1945 (O_1945,N_28899,N_29286);
and UO_1946 (O_1946,N_28071,N_29720);
nor UO_1947 (O_1947,N_27478,N_28430);
nand UO_1948 (O_1948,N_28698,N_29584);
xnor UO_1949 (O_1949,N_28361,N_28168);
or UO_1950 (O_1950,N_27346,N_29792);
or UO_1951 (O_1951,N_28491,N_29827);
nor UO_1952 (O_1952,N_27721,N_28969);
xnor UO_1953 (O_1953,N_27999,N_29188);
or UO_1954 (O_1954,N_28115,N_28593);
and UO_1955 (O_1955,N_29329,N_27993);
or UO_1956 (O_1956,N_29625,N_27447);
or UO_1957 (O_1957,N_27136,N_27691);
or UO_1958 (O_1958,N_29888,N_29646);
nand UO_1959 (O_1959,N_29953,N_28906);
or UO_1960 (O_1960,N_28257,N_29575);
nor UO_1961 (O_1961,N_28796,N_29886);
nand UO_1962 (O_1962,N_28072,N_27616);
nand UO_1963 (O_1963,N_28570,N_28548);
nor UO_1964 (O_1964,N_28804,N_29308);
and UO_1965 (O_1965,N_28804,N_29970);
or UO_1966 (O_1966,N_29957,N_29387);
or UO_1967 (O_1967,N_28973,N_27886);
nand UO_1968 (O_1968,N_28485,N_28250);
nor UO_1969 (O_1969,N_27852,N_29291);
and UO_1970 (O_1970,N_28755,N_27202);
nor UO_1971 (O_1971,N_28153,N_27985);
and UO_1972 (O_1972,N_28966,N_28063);
nor UO_1973 (O_1973,N_29383,N_28977);
and UO_1974 (O_1974,N_28720,N_29300);
nand UO_1975 (O_1975,N_27681,N_27346);
nand UO_1976 (O_1976,N_28185,N_27794);
or UO_1977 (O_1977,N_29202,N_27740);
nand UO_1978 (O_1978,N_29700,N_29867);
nand UO_1979 (O_1979,N_29969,N_29306);
and UO_1980 (O_1980,N_27262,N_28719);
or UO_1981 (O_1981,N_27485,N_27391);
and UO_1982 (O_1982,N_28884,N_27846);
nor UO_1983 (O_1983,N_29279,N_29124);
or UO_1984 (O_1984,N_29703,N_27710);
nor UO_1985 (O_1985,N_28401,N_27163);
or UO_1986 (O_1986,N_27120,N_29729);
nand UO_1987 (O_1987,N_27359,N_27312);
nor UO_1988 (O_1988,N_27113,N_28474);
nor UO_1989 (O_1989,N_29892,N_27417);
or UO_1990 (O_1990,N_27103,N_27429);
nor UO_1991 (O_1991,N_29676,N_29437);
or UO_1992 (O_1992,N_28813,N_28188);
and UO_1993 (O_1993,N_29765,N_27017);
or UO_1994 (O_1994,N_27954,N_27293);
and UO_1995 (O_1995,N_27386,N_29999);
nor UO_1996 (O_1996,N_29022,N_27795);
nor UO_1997 (O_1997,N_29705,N_27895);
or UO_1998 (O_1998,N_27930,N_27716);
or UO_1999 (O_1999,N_27102,N_27509);
and UO_2000 (O_2000,N_28787,N_28873);
nand UO_2001 (O_2001,N_28253,N_27726);
nor UO_2002 (O_2002,N_27694,N_27732);
and UO_2003 (O_2003,N_29447,N_28933);
nor UO_2004 (O_2004,N_28895,N_29223);
and UO_2005 (O_2005,N_27897,N_29924);
nor UO_2006 (O_2006,N_28723,N_28609);
nor UO_2007 (O_2007,N_28173,N_29215);
xnor UO_2008 (O_2008,N_29385,N_28443);
nand UO_2009 (O_2009,N_29266,N_28631);
and UO_2010 (O_2010,N_27628,N_29256);
or UO_2011 (O_2011,N_28412,N_29599);
and UO_2012 (O_2012,N_28471,N_27967);
xnor UO_2013 (O_2013,N_27129,N_28255);
nand UO_2014 (O_2014,N_28049,N_29818);
nand UO_2015 (O_2015,N_29872,N_28881);
nand UO_2016 (O_2016,N_27663,N_29168);
nand UO_2017 (O_2017,N_28737,N_29189);
or UO_2018 (O_2018,N_29268,N_29589);
nand UO_2019 (O_2019,N_29347,N_27257);
or UO_2020 (O_2020,N_28048,N_29653);
or UO_2021 (O_2021,N_29945,N_28241);
nor UO_2022 (O_2022,N_27240,N_28097);
xnor UO_2023 (O_2023,N_29740,N_29021);
or UO_2024 (O_2024,N_29420,N_28410);
nand UO_2025 (O_2025,N_27948,N_28719);
and UO_2026 (O_2026,N_27463,N_29653);
nand UO_2027 (O_2027,N_28943,N_27057);
nor UO_2028 (O_2028,N_28339,N_27078);
nand UO_2029 (O_2029,N_27369,N_29762);
nand UO_2030 (O_2030,N_27831,N_27074);
nand UO_2031 (O_2031,N_29970,N_27024);
nor UO_2032 (O_2032,N_27560,N_28289);
xnor UO_2033 (O_2033,N_29566,N_29211);
and UO_2034 (O_2034,N_29760,N_28003);
and UO_2035 (O_2035,N_27159,N_28680);
and UO_2036 (O_2036,N_27728,N_28603);
or UO_2037 (O_2037,N_27767,N_29689);
nand UO_2038 (O_2038,N_29391,N_28330);
nor UO_2039 (O_2039,N_29747,N_29774);
nand UO_2040 (O_2040,N_28082,N_28230);
nand UO_2041 (O_2041,N_28797,N_28188);
nand UO_2042 (O_2042,N_27615,N_28047);
nor UO_2043 (O_2043,N_28500,N_28577);
and UO_2044 (O_2044,N_29045,N_29221);
or UO_2045 (O_2045,N_27597,N_27553);
nand UO_2046 (O_2046,N_27935,N_28273);
and UO_2047 (O_2047,N_27378,N_29502);
nor UO_2048 (O_2048,N_29021,N_29843);
and UO_2049 (O_2049,N_28475,N_28031);
nor UO_2050 (O_2050,N_28128,N_28780);
and UO_2051 (O_2051,N_29321,N_27025);
and UO_2052 (O_2052,N_28079,N_29442);
and UO_2053 (O_2053,N_27116,N_27765);
and UO_2054 (O_2054,N_29986,N_28320);
xor UO_2055 (O_2055,N_29703,N_27610);
nand UO_2056 (O_2056,N_29070,N_28678);
nor UO_2057 (O_2057,N_27745,N_28118);
or UO_2058 (O_2058,N_28010,N_28173);
and UO_2059 (O_2059,N_29927,N_28125);
and UO_2060 (O_2060,N_27128,N_29038);
xnor UO_2061 (O_2061,N_28329,N_28597);
nor UO_2062 (O_2062,N_28389,N_29477);
nor UO_2063 (O_2063,N_29423,N_27720);
xnor UO_2064 (O_2064,N_29986,N_29339);
and UO_2065 (O_2065,N_28756,N_27952);
nor UO_2066 (O_2066,N_29773,N_27736);
nor UO_2067 (O_2067,N_28801,N_27790);
nor UO_2068 (O_2068,N_29777,N_28719);
or UO_2069 (O_2069,N_29494,N_29340);
nor UO_2070 (O_2070,N_29799,N_29498);
or UO_2071 (O_2071,N_28146,N_27871);
nand UO_2072 (O_2072,N_28955,N_28717);
or UO_2073 (O_2073,N_27670,N_28484);
and UO_2074 (O_2074,N_29806,N_28100);
nand UO_2075 (O_2075,N_29755,N_27628);
xor UO_2076 (O_2076,N_29117,N_27568);
nor UO_2077 (O_2077,N_27097,N_29579);
nand UO_2078 (O_2078,N_28136,N_28976);
nand UO_2079 (O_2079,N_27202,N_28340);
and UO_2080 (O_2080,N_28282,N_27512);
nor UO_2081 (O_2081,N_28019,N_27636);
nand UO_2082 (O_2082,N_28371,N_27638);
and UO_2083 (O_2083,N_28789,N_28974);
or UO_2084 (O_2084,N_28163,N_28364);
nor UO_2085 (O_2085,N_27642,N_28418);
nand UO_2086 (O_2086,N_27415,N_29021);
nor UO_2087 (O_2087,N_29758,N_27716);
or UO_2088 (O_2088,N_28816,N_28036);
xnor UO_2089 (O_2089,N_29110,N_27695);
nand UO_2090 (O_2090,N_29275,N_28617);
nand UO_2091 (O_2091,N_28905,N_28040);
and UO_2092 (O_2092,N_29975,N_27984);
nor UO_2093 (O_2093,N_28713,N_29224);
or UO_2094 (O_2094,N_27391,N_28976);
or UO_2095 (O_2095,N_29870,N_27310);
or UO_2096 (O_2096,N_29386,N_27373);
nor UO_2097 (O_2097,N_28753,N_29393);
and UO_2098 (O_2098,N_27415,N_27248);
nor UO_2099 (O_2099,N_29359,N_27541);
nand UO_2100 (O_2100,N_28623,N_29857);
nand UO_2101 (O_2101,N_28056,N_27558);
and UO_2102 (O_2102,N_28766,N_29527);
nor UO_2103 (O_2103,N_29505,N_29763);
and UO_2104 (O_2104,N_27502,N_29216);
nor UO_2105 (O_2105,N_29940,N_28301);
and UO_2106 (O_2106,N_29250,N_28238);
nand UO_2107 (O_2107,N_27391,N_29968);
or UO_2108 (O_2108,N_28299,N_28198);
and UO_2109 (O_2109,N_29904,N_27852);
and UO_2110 (O_2110,N_29388,N_28645);
and UO_2111 (O_2111,N_29659,N_28808);
and UO_2112 (O_2112,N_27778,N_29579);
and UO_2113 (O_2113,N_29659,N_27323);
xnor UO_2114 (O_2114,N_28996,N_29669);
and UO_2115 (O_2115,N_29999,N_29851);
and UO_2116 (O_2116,N_28447,N_27150);
or UO_2117 (O_2117,N_28401,N_27770);
nor UO_2118 (O_2118,N_29346,N_27992);
nor UO_2119 (O_2119,N_28728,N_28898);
or UO_2120 (O_2120,N_28172,N_28901);
nand UO_2121 (O_2121,N_28066,N_27220);
and UO_2122 (O_2122,N_28288,N_28054);
nor UO_2123 (O_2123,N_28073,N_28941);
nand UO_2124 (O_2124,N_28831,N_28160);
nor UO_2125 (O_2125,N_27561,N_28900);
and UO_2126 (O_2126,N_29935,N_29607);
nor UO_2127 (O_2127,N_29254,N_28518);
nor UO_2128 (O_2128,N_27324,N_28980);
nor UO_2129 (O_2129,N_28315,N_28846);
or UO_2130 (O_2130,N_28710,N_29247);
xnor UO_2131 (O_2131,N_27063,N_28145);
nor UO_2132 (O_2132,N_27782,N_29698);
xnor UO_2133 (O_2133,N_27046,N_29690);
xnor UO_2134 (O_2134,N_27917,N_27394);
xnor UO_2135 (O_2135,N_28095,N_27824);
or UO_2136 (O_2136,N_29903,N_29340);
nand UO_2137 (O_2137,N_28496,N_28010);
or UO_2138 (O_2138,N_27387,N_27343);
nor UO_2139 (O_2139,N_27717,N_27981);
nor UO_2140 (O_2140,N_28999,N_29395);
nor UO_2141 (O_2141,N_29958,N_28513);
xnor UO_2142 (O_2142,N_29193,N_28288);
xnor UO_2143 (O_2143,N_29153,N_28173);
and UO_2144 (O_2144,N_28562,N_27461);
nor UO_2145 (O_2145,N_27647,N_27068);
or UO_2146 (O_2146,N_28740,N_28735);
or UO_2147 (O_2147,N_29248,N_27924);
xor UO_2148 (O_2148,N_27647,N_27262);
or UO_2149 (O_2149,N_28027,N_28870);
and UO_2150 (O_2150,N_29914,N_29644);
and UO_2151 (O_2151,N_28878,N_28068);
or UO_2152 (O_2152,N_28248,N_27507);
and UO_2153 (O_2153,N_29857,N_27520);
nor UO_2154 (O_2154,N_28914,N_29435);
and UO_2155 (O_2155,N_28555,N_29074);
nand UO_2156 (O_2156,N_29896,N_28762);
nor UO_2157 (O_2157,N_28302,N_29690);
nand UO_2158 (O_2158,N_29939,N_29519);
nand UO_2159 (O_2159,N_28792,N_28779);
or UO_2160 (O_2160,N_29891,N_27349);
or UO_2161 (O_2161,N_28253,N_29272);
xor UO_2162 (O_2162,N_29244,N_27013);
and UO_2163 (O_2163,N_29034,N_28375);
nand UO_2164 (O_2164,N_29950,N_28068);
nand UO_2165 (O_2165,N_28836,N_27630);
nand UO_2166 (O_2166,N_29347,N_28197);
xnor UO_2167 (O_2167,N_28954,N_27911);
xor UO_2168 (O_2168,N_29469,N_28675);
and UO_2169 (O_2169,N_27941,N_28576);
xor UO_2170 (O_2170,N_27309,N_27728);
and UO_2171 (O_2171,N_28918,N_28023);
xnor UO_2172 (O_2172,N_27289,N_27822);
nor UO_2173 (O_2173,N_27527,N_28462);
or UO_2174 (O_2174,N_29367,N_28600);
nand UO_2175 (O_2175,N_28436,N_28640);
and UO_2176 (O_2176,N_27753,N_27078);
and UO_2177 (O_2177,N_27386,N_28004);
xor UO_2178 (O_2178,N_29021,N_29197);
and UO_2179 (O_2179,N_28938,N_29071);
or UO_2180 (O_2180,N_28068,N_27234);
or UO_2181 (O_2181,N_27278,N_28042);
xor UO_2182 (O_2182,N_28623,N_29876);
xor UO_2183 (O_2183,N_27363,N_28852);
nor UO_2184 (O_2184,N_29731,N_29412);
and UO_2185 (O_2185,N_27338,N_27930);
and UO_2186 (O_2186,N_29144,N_29243);
or UO_2187 (O_2187,N_29548,N_28480);
nor UO_2188 (O_2188,N_29165,N_29508);
nor UO_2189 (O_2189,N_29707,N_28335);
or UO_2190 (O_2190,N_27793,N_28728);
and UO_2191 (O_2191,N_28832,N_29160);
and UO_2192 (O_2192,N_28474,N_27412);
xnor UO_2193 (O_2193,N_29592,N_28324);
nor UO_2194 (O_2194,N_27990,N_28982);
nor UO_2195 (O_2195,N_28677,N_28597);
nand UO_2196 (O_2196,N_29124,N_27193);
nand UO_2197 (O_2197,N_28290,N_29878);
and UO_2198 (O_2198,N_29248,N_29324);
nand UO_2199 (O_2199,N_28905,N_27107);
nor UO_2200 (O_2200,N_29474,N_29173);
or UO_2201 (O_2201,N_29175,N_27039);
nor UO_2202 (O_2202,N_29795,N_27900);
nor UO_2203 (O_2203,N_27307,N_28730);
nand UO_2204 (O_2204,N_29788,N_29992);
nand UO_2205 (O_2205,N_28125,N_27928);
nor UO_2206 (O_2206,N_28247,N_29986);
nand UO_2207 (O_2207,N_29517,N_28655);
nor UO_2208 (O_2208,N_27850,N_27042);
nand UO_2209 (O_2209,N_27611,N_28639);
nand UO_2210 (O_2210,N_27830,N_27233);
xnor UO_2211 (O_2211,N_27099,N_29661);
nor UO_2212 (O_2212,N_28410,N_27370);
and UO_2213 (O_2213,N_29800,N_28404);
nand UO_2214 (O_2214,N_28983,N_28727);
and UO_2215 (O_2215,N_29944,N_27961);
and UO_2216 (O_2216,N_27248,N_27874);
and UO_2217 (O_2217,N_28798,N_27035);
nand UO_2218 (O_2218,N_27538,N_29949);
and UO_2219 (O_2219,N_27009,N_29147);
and UO_2220 (O_2220,N_27529,N_28516);
nand UO_2221 (O_2221,N_29024,N_28911);
or UO_2222 (O_2222,N_29732,N_27567);
and UO_2223 (O_2223,N_27866,N_29198);
and UO_2224 (O_2224,N_29559,N_29034);
nor UO_2225 (O_2225,N_29731,N_28040);
nand UO_2226 (O_2226,N_29703,N_29109);
nand UO_2227 (O_2227,N_29139,N_29538);
and UO_2228 (O_2228,N_28329,N_28762);
and UO_2229 (O_2229,N_28628,N_27050);
xnor UO_2230 (O_2230,N_27530,N_29207);
or UO_2231 (O_2231,N_29620,N_29333);
nor UO_2232 (O_2232,N_29318,N_27386);
or UO_2233 (O_2233,N_29988,N_27578);
and UO_2234 (O_2234,N_29538,N_27205);
nand UO_2235 (O_2235,N_27421,N_29126);
nor UO_2236 (O_2236,N_28491,N_27158);
nor UO_2237 (O_2237,N_29751,N_29571);
xor UO_2238 (O_2238,N_28643,N_29001);
nor UO_2239 (O_2239,N_28021,N_28817);
nand UO_2240 (O_2240,N_27065,N_29050);
nand UO_2241 (O_2241,N_29078,N_29370);
nand UO_2242 (O_2242,N_28668,N_27527);
or UO_2243 (O_2243,N_28612,N_28133);
xor UO_2244 (O_2244,N_29862,N_28448);
xnor UO_2245 (O_2245,N_27240,N_28633);
and UO_2246 (O_2246,N_28060,N_27686);
nand UO_2247 (O_2247,N_28658,N_28180);
nor UO_2248 (O_2248,N_29119,N_27681);
xor UO_2249 (O_2249,N_29105,N_29980);
nor UO_2250 (O_2250,N_29743,N_28125);
and UO_2251 (O_2251,N_29259,N_28182);
and UO_2252 (O_2252,N_27964,N_29284);
or UO_2253 (O_2253,N_29455,N_29524);
and UO_2254 (O_2254,N_28769,N_29289);
nand UO_2255 (O_2255,N_27580,N_29251);
nand UO_2256 (O_2256,N_28720,N_27692);
or UO_2257 (O_2257,N_27750,N_29370);
or UO_2258 (O_2258,N_28079,N_28292);
nor UO_2259 (O_2259,N_29622,N_27733);
and UO_2260 (O_2260,N_29004,N_29664);
xor UO_2261 (O_2261,N_29755,N_28797);
nor UO_2262 (O_2262,N_27208,N_28140);
or UO_2263 (O_2263,N_28492,N_28803);
nor UO_2264 (O_2264,N_27298,N_27852);
nor UO_2265 (O_2265,N_29900,N_27383);
xor UO_2266 (O_2266,N_27969,N_29303);
and UO_2267 (O_2267,N_27405,N_28106);
nand UO_2268 (O_2268,N_29785,N_27269);
nor UO_2269 (O_2269,N_29906,N_28823);
xor UO_2270 (O_2270,N_28533,N_28041);
nor UO_2271 (O_2271,N_28654,N_27631);
or UO_2272 (O_2272,N_27501,N_27385);
nand UO_2273 (O_2273,N_28689,N_29940);
and UO_2274 (O_2274,N_28799,N_29139);
or UO_2275 (O_2275,N_29903,N_28642);
xor UO_2276 (O_2276,N_29925,N_27146);
xor UO_2277 (O_2277,N_28704,N_27707);
xor UO_2278 (O_2278,N_27279,N_29622);
nor UO_2279 (O_2279,N_27698,N_27442);
and UO_2280 (O_2280,N_29242,N_29911);
and UO_2281 (O_2281,N_27682,N_27144);
or UO_2282 (O_2282,N_29737,N_29800);
nor UO_2283 (O_2283,N_29770,N_28912);
nand UO_2284 (O_2284,N_28030,N_29820);
nand UO_2285 (O_2285,N_27089,N_27396);
or UO_2286 (O_2286,N_29244,N_29784);
xnor UO_2287 (O_2287,N_27211,N_28016);
or UO_2288 (O_2288,N_29434,N_27901);
or UO_2289 (O_2289,N_29373,N_29386);
and UO_2290 (O_2290,N_29336,N_29905);
nand UO_2291 (O_2291,N_28850,N_29058);
or UO_2292 (O_2292,N_27859,N_29057);
or UO_2293 (O_2293,N_27194,N_27076);
nor UO_2294 (O_2294,N_29542,N_27148);
nor UO_2295 (O_2295,N_29110,N_29694);
nor UO_2296 (O_2296,N_29594,N_28641);
and UO_2297 (O_2297,N_29296,N_28818);
and UO_2298 (O_2298,N_29959,N_27287);
and UO_2299 (O_2299,N_28345,N_29763);
nor UO_2300 (O_2300,N_29785,N_27277);
or UO_2301 (O_2301,N_29525,N_27328);
nor UO_2302 (O_2302,N_29465,N_29468);
nor UO_2303 (O_2303,N_29620,N_29193);
nor UO_2304 (O_2304,N_28373,N_27020);
and UO_2305 (O_2305,N_27213,N_28827);
or UO_2306 (O_2306,N_27219,N_27026);
nand UO_2307 (O_2307,N_28804,N_29557);
and UO_2308 (O_2308,N_28551,N_29502);
nand UO_2309 (O_2309,N_27889,N_27894);
xnor UO_2310 (O_2310,N_27306,N_27971);
or UO_2311 (O_2311,N_27958,N_29561);
nor UO_2312 (O_2312,N_28630,N_29769);
or UO_2313 (O_2313,N_27702,N_27456);
xor UO_2314 (O_2314,N_27171,N_28010);
xnor UO_2315 (O_2315,N_28141,N_29656);
xnor UO_2316 (O_2316,N_28062,N_28980);
or UO_2317 (O_2317,N_27740,N_29910);
xnor UO_2318 (O_2318,N_28544,N_28724);
and UO_2319 (O_2319,N_27225,N_29196);
nand UO_2320 (O_2320,N_29240,N_29691);
nand UO_2321 (O_2321,N_27898,N_29552);
nand UO_2322 (O_2322,N_27063,N_29610);
nor UO_2323 (O_2323,N_28575,N_27862);
nor UO_2324 (O_2324,N_28770,N_28691);
nor UO_2325 (O_2325,N_27084,N_28393);
nand UO_2326 (O_2326,N_28737,N_28619);
and UO_2327 (O_2327,N_29955,N_29614);
or UO_2328 (O_2328,N_29749,N_29874);
nor UO_2329 (O_2329,N_27152,N_28137);
nor UO_2330 (O_2330,N_28178,N_27359);
or UO_2331 (O_2331,N_27690,N_27560);
or UO_2332 (O_2332,N_29568,N_28777);
xor UO_2333 (O_2333,N_28191,N_28320);
nand UO_2334 (O_2334,N_29044,N_29343);
and UO_2335 (O_2335,N_29618,N_28631);
nand UO_2336 (O_2336,N_27046,N_28089);
nand UO_2337 (O_2337,N_27718,N_29070);
nand UO_2338 (O_2338,N_27556,N_29633);
nor UO_2339 (O_2339,N_27162,N_27418);
or UO_2340 (O_2340,N_29166,N_29209);
or UO_2341 (O_2341,N_29343,N_28897);
nor UO_2342 (O_2342,N_28091,N_28728);
or UO_2343 (O_2343,N_29567,N_29225);
nor UO_2344 (O_2344,N_29963,N_27999);
or UO_2345 (O_2345,N_28512,N_29538);
and UO_2346 (O_2346,N_28530,N_28542);
and UO_2347 (O_2347,N_29942,N_29966);
and UO_2348 (O_2348,N_27185,N_28403);
or UO_2349 (O_2349,N_27539,N_27805);
nor UO_2350 (O_2350,N_29922,N_28275);
nor UO_2351 (O_2351,N_28423,N_27729);
and UO_2352 (O_2352,N_29946,N_28204);
and UO_2353 (O_2353,N_28909,N_28194);
or UO_2354 (O_2354,N_27480,N_27836);
nand UO_2355 (O_2355,N_28567,N_28746);
and UO_2356 (O_2356,N_28538,N_27061);
or UO_2357 (O_2357,N_29083,N_29887);
or UO_2358 (O_2358,N_29097,N_28893);
or UO_2359 (O_2359,N_29090,N_29946);
and UO_2360 (O_2360,N_28475,N_29630);
nor UO_2361 (O_2361,N_29525,N_28454);
nor UO_2362 (O_2362,N_27606,N_28643);
nand UO_2363 (O_2363,N_28429,N_28790);
nand UO_2364 (O_2364,N_28121,N_27927);
or UO_2365 (O_2365,N_28275,N_28072);
nand UO_2366 (O_2366,N_27112,N_27908);
or UO_2367 (O_2367,N_27411,N_28683);
xnor UO_2368 (O_2368,N_29921,N_29538);
or UO_2369 (O_2369,N_29180,N_28309);
and UO_2370 (O_2370,N_28586,N_28964);
nor UO_2371 (O_2371,N_29205,N_28112);
or UO_2372 (O_2372,N_27028,N_27985);
and UO_2373 (O_2373,N_29121,N_29429);
or UO_2374 (O_2374,N_29109,N_29555);
nor UO_2375 (O_2375,N_27051,N_28893);
nand UO_2376 (O_2376,N_27019,N_28458);
nor UO_2377 (O_2377,N_27656,N_27920);
and UO_2378 (O_2378,N_29817,N_27363);
nand UO_2379 (O_2379,N_29599,N_29919);
or UO_2380 (O_2380,N_29178,N_27029);
nor UO_2381 (O_2381,N_27498,N_29413);
nor UO_2382 (O_2382,N_28902,N_28746);
nand UO_2383 (O_2383,N_29783,N_29437);
xnor UO_2384 (O_2384,N_28483,N_28041);
and UO_2385 (O_2385,N_29496,N_27561);
or UO_2386 (O_2386,N_29871,N_29861);
or UO_2387 (O_2387,N_27672,N_29198);
nand UO_2388 (O_2388,N_28233,N_28611);
or UO_2389 (O_2389,N_27023,N_29708);
or UO_2390 (O_2390,N_29141,N_27085);
and UO_2391 (O_2391,N_27037,N_28021);
or UO_2392 (O_2392,N_29403,N_29312);
nor UO_2393 (O_2393,N_29909,N_29076);
nand UO_2394 (O_2394,N_27717,N_29763);
and UO_2395 (O_2395,N_27139,N_28728);
or UO_2396 (O_2396,N_27213,N_29204);
and UO_2397 (O_2397,N_27546,N_27766);
or UO_2398 (O_2398,N_29773,N_28143);
nand UO_2399 (O_2399,N_27342,N_27185);
nand UO_2400 (O_2400,N_28173,N_27965);
nor UO_2401 (O_2401,N_27176,N_29205);
or UO_2402 (O_2402,N_27591,N_29238);
and UO_2403 (O_2403,N_29245,N_27285);
or UO_2404 (O_2404,N_27437,N_29801);
xnor UO_2405 (O_2405,N_29321,N_28178);
nand UO_2406 (O_2406,N_28385,N_29203);
and UO_2407 (O_2407,N_27095,N_28601);
nand UO_2408 (O_2408,N_28870,N_28883);
nand UO_2409 (O_2409,N_29633,N_29696);
nor UO_2410 (O_2410,N_27192,N_28683);
or UO_2411 (O_2411,N_28312,N_28962);
xor UO_2412 (O_2412,N_28310,N_27163);
nor UO_2413 (O_2413,N_28687,N_29265);
nand UO_2414 (O_2414,N_29276,N_27041);
and UO_2415 (O_2415,N_27810,N_29946);
nor UO_2416 (O_2416,N_29099,N_29393);
or UO_2417 (O_2417,N_29472,N_27247);
and UO_2418 (O_2418,N_28643,N_29778);
xnor UO_2419 (O_2419,N_27459,N_28241);
nor UO_2420 (O_2420,N_27178,N_29406);
xor UO_2421 (O_2421,N_29361,N_28461);
and UO_2422 (O_2422,N_28387,N_27210);
nor UO_2423 (O_2423,N_28006,N_27787);
nand UO_2424 (O_2424,N_29816,N_28964);
or UO_2425 (O_2425,N_28196,N_28740);
or UO_2426 (O_2426,N_28492,N_28888);
and UO_2427 (O_2427,N_28015,N_28108);
nand UO_2428 (O_2428,N_27527,N_28415);
and UO_2429 (O_2429,N_27321,N_29762);
nor UO_2430 (O_2430,N_29457,N_28134);
nor UO_2431 (O_2431,N_28536,N_27917);
and UO_2432 (O_2432,N_28883,N_28483);
and UO_2433 (O_2433,N_29293,N_29417);
nand UO_2434 (O_2434,N_27279,N_29061);
or UO_2435 (O_2435,N_28952,N_28708);
nor UO_2436 (O_2436,N_27781,N_29302);
nand UO_2437 (O_2437,N_29299,N_29542);
or UO_2438 (O_2438,N_28290,N_28764);
xnor UO_2439 (O_2439,N_28424,N_27674);
nand UO_2440 (O_2440,N_29288,N_28501);
nand UO_2441 (O_2441,N_28352,N_28846);
nor UO_2442 (O_2442,N_29922,N_27912);
nand UO_2443 (O_2443,N_29851,N_29413);
or UO_2444 (O_2444,N_27486,N_28325);
or UO_2445 (O_2445,N_29137,N_29149);
nand UO_2446 (O_2446,N_29161,N_28784);
nor UO_2447 (O_2447,N_29552,N_27917);
xor UO_2448 (O_2448,N_29005,N_28026);
or UO_2449 (O_2449,N_28025,N_27225);
nor UO_2450 (O_2450,N_29202,N_27718);
nand UO_2451 (O_2451,N_29925,N_27742);
and UO_2452 (O_2452,N_27062,N_29353);
nand UO_2453 (O_2453,N_27908,N_27757);
nand UO_2454 (O_2454,N_28151,N_29918);
nor UO_2455 (O_2455,N_28578,N_28523);
or UO_2456 (O_2456,N_29273,N_29106);
nand UO_2457 (O_2457,N_29921,N_28926);
or UO_2458 (O_2458,N_27745,N_28661);
and UO_2459 (O_2459,N_27743,N_29539);
or UO_2460 (O_2460,N_27071,N_29467);
xnor UO_2461 (O_2461,N_28701,N_27899);
or UO_2462 (O_2462,N_28133,N_27782);
nor UO_2463 (O_2463,N_28031,N_27400);
or UO_2464 (O_2464,N_27403,N_29871);
nor UO_2465 (O_2465,N_27306,N_28324);
nor UO_2466 (O_2466,N_29766,N_28622);
or UO_2467 (O_2467,N_28879,N_27138);
and UO_2468 (O_2468,N_27124,N_28554);
and UO_2469 (O_2469,N_28773,N_27854);
xor UO_2470 (O_2470,N_29618,N_29714);
xor UO_2471 (O_2471,N_27884,N_27788);
nor UO_2472 (O_2472,N_28219,N_27218);
nor UO_2473 (O_2473,N_28390,N_27718);
nand UO_2474 (O_2474,N_28330,N_27109);
and UO_2475 (O_2475,N_28576,N_28686);
and UO_2476 (O_2476,N_27793,N_27376);
nor UO_2477 (O_2477,N_29132,N_27533);
or UO_2478 (O_2478,N_28953,N_28882);
nor UO_2479 (O_2479,N_27344,N_27589);
and UO_2480 (O_2480,N_27598,N_27830);
and UO_2481 (O_2481,N_28104,N_27731);
and UO_2482 (O_2482,N_28053,N_28912);
nor UO_2483 (O_2483,N_28126,N_29938);
or UO_2484 (O_2484,N_28517,N_28132);
and UO_2485 (O_2485,N_29972,N_29956);
nor UO_2486 (O_2486,N_28277,N_27081);
nand UO_2487 (O_2487,N_27279,N_28756);
nand UO_2488 (O_2488,N_27071,N_29967);
and UO_2489 (O_2489,N_29230,N_27132);
nor UO_2490 (O_2490,N_28929,N_28111);
and UO_2491 (O_2491,N_27734,N_28690);
nand UO_2492 (O_2492,N_29408,N_28364);
and UO_2493 (O_2493,N_27591,N_28618);
xor UO_2494 (O_2494,N_29372,N_27395);
nand UO_2495 (O_2495,N_28835,N_27823);
and UO_2496 (O_2496,N_28490,N_28959);
xor UO_2497 (O_2497,N_29582,N_28693);
nand UO_2498 (O_2498,N_27173,N_27912);
and UO_2499 (O_2499,N_27312,N_28283);
nor UO_2500 (O_2500,N_28973,N_29751);
nor UO_2501 (O_2501,N_27000,N_29627);
nand UO_2502 (O_2502,N_27150,N_27703);
nor UO_2503 (O_2503,N_27533,N_27988);
nand UO_2504 (O_2504,N_27871,N_27392);
xnor UO_2505 (O_2505,N_27048,N_28689);
nand UO_2506 (O_2506,N_28615,N_27838);
nand UO_2507 (O_2507,N_29627,N_28479);
nand UO_2508 (O_2508,N_29099,N_29566);
xor UO_2509 (O_2509,N_28690,N_29335);
nor UO_2510 (O_2510,N_27682,N_28802);
and UO_2511 (O_2511,N_28033,N_27340);
or UO_2512 (O_2512,N_27281,N_27449);
xnor UO_2513 (O_2513,N_27529,N_28821);
and UO_2514 (O_2514,N_27084,N_27349);
nor UO_2515 (O_2515,N_29817,N_28027);
or UO_2516 (O_2516,N_29665,N_27114);
nor UO_2517 (O_2517,N_29539,N_27884);
and UO_2518 (O_2518,N_28785,N_28739);
nand UO_2519 (O_2519,N_28121,N_27280);
and UO_2520 (O_2520,N_29073,N_29080);
nor UO_2521 (O_2521,N_28224,N_29553);
nand UO_2522 (O_2522,N_29468,N_29090);
nand UO_2523 (O_2523,N_28703,N_29953);
nand UO_2524 (O_2524,N_28433,N_28509);
nand UO_2525 (O_2525,N_27817,N_28002);
nor UO_2526 (O_2526,N_28498,N_27413);
nand UO_2527 (O_2527,N_27956,N_29714);
nor UO_2528 (O_2528,N_27990,N_29822);
nor UO_2529 (O_2529,N_28589,N_29278);
xor UO_2530 (O_2530,N_29900,N_28038);
and UO_2531 (O_2531,N_29240,N_29061);
nor UO_2532 (O_2532,N_28181,N_28639);
nand UO_2533 (O_2533,N_27978,N_29904);
or UO_2534 (O_2534,N_28867,N_29674);
nor UO_2535 (O_2535,N_29637,N_28774);
nand UO_2536 (O_2536,N_27690,N_27143);
nand UO_2537 (O_2537,N_28178,N_27176);
or UO_2538 (O_2538,N_29339,N_27596);
nor UO_2539 (O_2539,N_29265,N_27160);
nor UO_2540 (O_2540,N_29353,N_28958);
and UO_2541 (O_2541,N_27354,N_28490);
nor UO_2542 (O_2542,N_28091,N_27697);
and UO_2543 (O_2543,N_29701,N_28424);
nor UO_2544 (O_2544,N_28364,N_27248);
or UO_2545 (O_2545,N_28867,N_29888);
and UO_2546 (O_2546,N_27564,N_29842);
xnor UO_2547 (O_2547,N_29150,N_27695);
and UO_2548 (O_2548,N_29959,N_27323);
nand UO_2549 (O_2549,N_29231,N_27897);
nor UO_2550 (O_2550,N_28121,N_29034);
xnor UO_2551 (O_2551,N_29749,N_29625);
nand UO_2552 (O_2552,N_27189,N_29203);
and UO_2553 (O_2553,N_27589,N_28233);
xor UO_2554 (O_2554,N_27256,N_27787);
or UO_2555 (O_2555,N_28468,N_29829);
or UO_2556 (O_2556,N_27636,N_27251);
nand UO_2557 (O_2557,N_29668,N_29178);
or UO_2558 (O_2558,N_27466,N_27217);
nor UO_2559 (O_2559,N_29369,N_28451);
xor UO_2560 (O_2560,N_29388,N_29848);
nand UO_2561 (O_2561,N_27985,N_27277);
or UO_2562 (O_2562,N_27857,N_27025);
nand UO_2563 (O_2563,N_29402,N_27014);
or UO_2564 (O_2564,N_27343,N_27995);
nor UO_2565 (O_2565,N_29269,N_28625);
or UO_2566 (O_2566,N_29315,N_29057);
and UO_2567 (O_2567,N_28016,N_27994);
nand UO_2568 (O_2568,N_29278,N_28507);
nor UO_2569 (O_2569,N_28593,N_29675);
nor UO_2570 (O_2570,N_27199,N_27520);
xnor UO_2571 (O_2571,N_28206,N_27661);
nand UO_2572 (O_2572,N_27941,N_28419);
or UO_2573 (O_2573,N_29804,N_27568);
nor UO_2574 (O_2574,N_27504,N_27743);
and UO_2575 (O_2575,N_27259,N_27907);
and UO_2576 (O_2576,N_28245,N_27374);
nor UO_2577 (O_2577,N_29107,N_29353);
nand UO_2578 (O_2578,N_29597,N_29002);
and UO_2579 (O_2579,N_29604,N_28444);
nand UO_2580 (O_2580,N_28675,N_29175);
xnor UO_2581 (O_2581,N_27480,N_27328);
xor UO_2582 (O_2582,N_27011,N_28742);
or UO_2583 (O_2583,N_28750,N_29767);
and UO_2584 (O_2584,N_29759,N_27482);
xor UO_2585 (O_2585,N_29285,N_28233);
or UO_2586 (O_2586,N_29158,N_27175);
and UO_2587 (O_2587,N_27015,N_27589);
or UO_2588 (O_2588,N_28141,N_29585);
nor UO_2589 (O_2589,N_27657,N_28583);
nor UO_2590 (O_2590,N_28680,N_28876);
nor UO_2591 (O_2591,N_28500,N_28276);
xor UO_2592 (O_2592,N_29204,N_27804);
nand UO_2593 (O_2593,N_27556,N_27180);
or UO_2594 (O_2594,N_27106,N_29424);
or UO_2595 (O_2595,N_28748,N_29708);
nand UO_2596 (O_2596,N_29183,N_28830);
nand UO_2597 (O_2597,N_27528,N_29501);
nor UO_2598 (O_2598,N_27127,N_29174);
nand UO_2599 (O_2599,N_29742,N_27134);
nor UO_2600 (O_2600,N_27189,N_28755);
xnor UO_2601 (O_2601,N_28257,N_29231);
and UO_2602 (O_2602,N_28345,N_27673);
nor UO_2603 (O_2603,N_27479,N_28747);
and UO_2604 (O_2604,N_27770,N_27576);
or UO_2605 (O_2605,N_27365,N_27487);
and UO_2606 (O_2606,N_29106,N_27309);
nor UO_2607 (O_2607,N_28283,N_28263);
nand UO_2608 (O_2608,N_29484,N_29086);
and UO_2609 (O_2609,N_27909,N_29063);
nand UO_2610 (O_2610,N_27804,N_29805);
xnor UO_2611 (O_2611,N_27560,N_27257);
nand UO_2612 (O_2612,N_27855,N_27102);
nor UO_2613 (O_2613,N_29923,N_27155);
nand UO_2614 (O_2614,N_27676,N_29242);
xor UO_2615 (O_2615,N_28612,N_29867);
nand UO_2616 (O_2616,N_27519,N_27516);
nor UO_2617 (O_2617,N_29690,N_27142);
nand UO_2618 (O_2618,N_27713,N_27027);
and UO_2619 (O_2619,N_27817,N_27190);
or UO_2620 (O_2620,N_27272,N_27269);
or UO_2621 (O_2621,N_29403,N_28476);
nand UO_2622 (O_2622,N_27159,N_28794);
nor UO_2623 (O_2623,N_28449,N_28852);
xnor UO_2624 (O_2624,N_29727,N_28192);
and UO_2625 (O_2625,N_28200,N_29160);
nor UO_2626 (O_2626,N_27342,N_29120);
nor UO_2627 (O_2627,N_29079,N_27829);
or UO_2628 (O_2628,N_29604,N_29434);
and UO_2629 (O_2629,N_28934,N_28049);
nor UO_2630 (O_2630,N_27863,N_27161);
xnor UO_2631 (O_2631,N_27558,N_29505);
nand UO_2632 (O_2632,N_28053,N_28087);
and UO_2633 (O_2633,N_27615,N_28077);
nor UO_2634 (O_2634,N_28488,N_29229);
or UO_2635 (O_2635,N_27018,N_29947);
or UO_2636 (O_2636,N_28987,N_28719);
and UO_2637 (O_2637,N_27520,N_27912);
and UO_2638 (O_2638,N_27238,N_29306);
nor UO_2639 (O_2639,N_28177,N_29812);
and UO_2640 (O_2640,N_27147,N_29452);
nor UO_2641 (O_2641,N_29796,N_28877);
nor UO_2642 (O_2642,N_27497,N_28725);
nor UO_2643 (O_2643,N_28758,N_28205);
nor UO_2644 (O_2644,N_27663,N_27806);
or UO_2645 (O_2645,N_28591,N_29700);
xnor UO_2646 (O_2646,N_28770,N_29945);
nand UO_2647 (O_2647,N_29721,N_27110);
and UO_2648 (O_2648,N_27719,N_29815);
nor UO_2649 (O_2649,N_28751,N_27910);
nand UO_2650 (O_2650,N_28564,N_27184);
nand UO_2651 (O_2651,N_28568,N_29093);
nor UO_2652 (O_2652,N_28339,N_28294);
nor UO_2653 (O_2653,N_28385,N_28238);
or UO_2654 (O_2654,N_29692,N_28825);
nand UO_2655 (O_2655,N_27726,N_27112);
nand UO_2656 (O_2656,N_27532,N_29578);
nor UO_2657 (O_2657,N_27409,N_27384);
or UO_2658 (O_2658,N_27698,N_28615);
nand UO_2659 (O_2659,N_28163,N_29077);
nand UO_2660 (O_2660,N_29456,N_27979);
xor UO_2661 (O_2661,N_27082,N_27089);
and UO_2662 (O_2662,N_27155,N_27005);
and UO_2663 (O_2663,N_27017,N_28086);
and UO_2664 (O_2664,N_29162,N_28065);
nor UO_2665 (O_2665,N_29074,N_29318);
and UO_2666 (O_2666,N_27097,N_28463);
nand UO_2667 (O_2667,N_29226,N_27901);
nor UO_2668 (O_2668,N_27090,N_29756);
nor UO_2669 (O_2669,N_27957,N_27154);
xor UO_2670 (O_2670,N_29502,N_28837);
xor UO_2671 (O_2671,N_29017,N_27447);
and UO_2672 (O_2672,N_29742,N_27045);
nand UO_2673 (O_2673,N_28256,N_27460);
or UO_2674 (O_2674,N_29548,N_28324);
nand UO_2675 (O_2675,N_28469,N_27898);
nor UO_2676 (O_2676,N_29853,N_27382);
nor UO_2677 (O_2677,N_29867,N_28079);
and UO_2678 (O_2678,N_27005,N_29411);
or UO_2679 (O_2679,N_29804,N_27583);
and UO_2680 (O_2680,N_28057,N_28914);
or UO_2681 (O_2681,N_28155,N_28338);
nand UO_2682 (O_2682,N_29353,N_28155);
and UO_2683 (O_2683,N_29716,N_27268);
nor UO_2684 (O_2684,N_28914,N_29510);
nand UO_2685 (O_2685,N_28772,N_29389);
nor UO_2686 (O_2686,N_27035,N_27629);
and UO_2687 (O_2687,N_27162,N_28701);
xor UO_2688 (O_2688,N_28092,N_27031);
nand UO_2689 (O_2689,N_27009,N_28283);
or UO_2690 (O_2690,N_28029,N_28761);
nand UO_2691 (O_2691,N_27720,N_27031);
nand UO_2692 (O_2692,N_29583,N_29750);
and UO_2693 (O_2693,N_28807,N_27189);
nand UO_2694 (O_2694,N_27706,N_27752);
or UO_2695 (O_2695,N_27349,N_27649);
and UO_2696 (O_2696,N_28673,N_29064);
xor UO_2697 (O_2697,N_29055,N_29319);
and UO_2698 (O_2698,N_27585,N_28704);
nor UO_2699 (O_2699,N_28372,N_28564);
and UO_2700 (O_2700,N_28316,N_27152);
and UO_2701 (O_2701,N_27844,N_28579);
and UO_2702 (O_2702,N_27673,N_29832);
or UO_2703 (O_2703,N_28157,N_27817);
nand UO_2704 (O_2704,N_28360,N_29505);
or UO_2705 (O_2705,N_28941,N_27045);
and UO_2706 (O_2706,N_27324,N_28681);
or UO_2707 (O_2707,N_27513,N_28185);
and UO_2708 (O_2708,N_29126,N_29889);
xor UO_2709 (O_2709,N_29789,N_29462);
nand UO_2710 (O_2710,N_27919,N_28781);
nand UO_2711 (O_2711,N_27101,N_28616);
nand UO_2712 (O_2712,N_28005,N_27986);
or UO_2713 (O_2713,N_28296,N_28597);
and UO_2714 (O_2714,N_27153,N_29900);
or UO_2715 (O_2715,N_29005,N_27207);
and UO_2716 (O_2716,N_27170,N_27723);
and UO_2717 (O_2717,N_29219,N_27654);
nor UO_2718 (O_2718,N_28372,N_27848);
nor UO_2719 (O_2719,N_29203,N_27360);
and UO_2720 (O_2720,N_29223,N_27327);
nor UO_2721 (O_2721,N_27335,N_29194);
nor UO_2722 (O_2722,N_28693,N_29431);
nand UO_2723 (O_2723,N_27722,N_29062);
nand UO_2724 (O_2724,N_27277,N_28215);
nor UO_2725 (O_2725,N_28201,N_27985);
or UO_2726 (O_2726,N_29568,N_29560);
nor UO_2727 (O_2727,N_28289,N_29594);
nor UO_2728 (O_2728,N_27583,N_27122);
nand UO_2729 (O_2729,N_29109,N_27774);
nor UO_2730 (O_2730,N_27927,N_29806);
and UO_2731 (O_2731,N_28127,N_27574);
or UO_2732 (O_2732,N_27066,N_29231);
or UO_2733 (O_2733,N_27033,N_27345);
and UO_2734 (O_2734,N_29611,N_27023);
xnor UO_2735 (O_2735,N_29585,N_29950);
or UO_2736 (O_2736,N_27179,N_27321);
or UO_2737 (O_2737,N_28682,N_29334);
and UO_2738 (O_2738,N_28647,N_29950);
nand UO_2739 (O_2739,N_28360,N_27503);
or UO_2740 (O_2740,N_27940,N_28590);
nand UO_2741 (O_2741,N_28262,N_28786);
or UO_2742 (O_2742,N_28709,N_28281);
nand UO_2743 (O_2743,N_27198,N_29895);
or UO_2744 (O_2744,N_28591,N_27392);
nand UO_2745 (O_2745,N_27462,N_27294);
nand UO_2746 (O_2746,N_27755,N_28531);
nand UO_2747 (O_2747,N_29978,N_28780);
nand UO_2748 (O_2748,N_28227,N_28238);
nor UO_2749 (O_2749,N_28630,N_29812);
or UO_2750 (O_2750,N_29478,N_29396);
or UO_2751 (O_2751,N_27354,N_28487);
nor UO_2752 (O_2752,N_27314,N_27324);
or UO_2753 (O_2753,N_28951,N_28314);
xnor UO_2754 (O_2754,N_29975,N_29278);
and UO_2755 (O_2755,N_28472,N_28697);
and UO_2756 (O_2756,N_29932,N_28792);
nand UO_2757 (O_2757,N_28846,N_28865);
nand UO_2758 (O_2758,N_28270,N_27700);
and UO_2759 (O_2759,N_28092,N_28220);
and UO_2760 (O_2760,N_27253,N_29872);
nand UO_2761 (O_2761,N_27256,N_28149);
nand UO_2762 (O_2762,N_27119,N_27835);
nor UO_2763 (O_2763,N_29631,N_29590);
or UO_2764 (O_2764,N_27373,N_28370);
or UO_2765 (O_2765,N_28186,N_29667);
nor UO_2766 (O_2766,N_29339,N_27373);
or UO_2767 (O_2767,N_29608,N_28233);
or UO_2768 (O_2768,N_29821,N_28168);
and UO_2769 (O_2769,N_27408,N_27118);
nand UO_2770 (O_2770,N_27343,N_29478);
nand UO_2771 (O_2771,N_27895,N_27488);
nor UO_2772 (O_2772,N_28471,N_29345);
nor UO_2773 (O_2773,N_28121,N_29859);
xor UO_2774 (O_2774,N_27009,N_27568);
nor UO_2775 (O_2775,N_29844,N_27778);
and UO_2776 (O_2776,N_29395,N_27196);
nand UO_2777 (O_2777,N_27524,N_28271);
xor UO_2778 (O_2778,N_27001,N_28045);
or UO_2779 (O_2779,N_28711,N_28961);
nor UO_2780 (O_2780,N_27548,N_29752);
xnor UO_2781 (O_2781,N_28437,N_29506);
nand UO_2782 (O_2782,N_27135,N_27684);
nand UO_2783 (O_2783,N_29204,N_28837);
nand UO_2784 (O_2784,N_27006,N_27347);
or UO_2785 (O_2785,N_29175,N_29806);
nand UO_2786 (O_2786,N_29056,N_28755);
or UO_2787 (O_2787,N_27622,N_29789);
nor UO_2788 (O_2788,N_27969,N_27726);
and UO_2789 (O_2789,N_27870,N_28686);
nor UO_2790 (O_2790,N_27811,N_28105);
or UO_2791 (O_2791,N_28644,N_28439);
nand UO_2792 (O_2792,N_29435,N_28521);
and UO_2793 (O_2793,N_29047,N_28447);
nand UO_2794 (O_2794,N_29819,N_28199);
and UO_2795 (O_2795,N_28458,N_29171);
nor UO_2796 (O_2796,N_29139,N_29219);
or UO_2797 (O_2797,N_27260,N_27198);
or UO_2798 (O_2798,N_28786,N_29824);
nor UO_2799 (O_2799,N_28586,N_29708);
nand UO_2800 (O_2800,N_28636,N_29585);
nor UO_2801 (O_2801,N_29358,N_28184);
xnor UO_2802 (O_2802,N_28733,N_27400);
xnor UO_2803 (O_2803,N_28018,N_27370);
nand UO_2804 (O_2804,N_28709,N_28796);
nor UO_2805 (O_2805,N_29312,N_28018);
xnor UO_2806 (O_2806,N_27681,N_28646);
nand UO_2807 (O_2807,N_28619,N_28296);
nand UO_2808 (O_2808,N_29373,N_28399);
nand UO_2809 (O_2809,N_29811,N_27229);
nor UO_2810 (O_2810,N_28114,N_29561);
or UO_2811 (O_2811,N_28055,N_27579);
or UO_2812 (O_2812,N_29095,N_28884);
nor UO_2813 (O_2813,N_27432,N_27410);
or UO_2814 (O_2814,N_28767,N_28261);
and UO_2815 (O_2815,N_27190,N_28228);
or UO_2816 (O_2816,N_29311,N_28344);
nor UO_2817 (O_2817,N_27570,N_28032);
nor UO_2818 (O_2818,N_27097,N_28982);
nor UO_2819 (O_2819,N_28924,N_29057);
nand UO_2820 (O_2820,N_28244,N_27617);
nand UO_2821 (O_2821,N_27197,N_27094);
xor UO_2822 (O_2822,N_27486,N_29931);
or UO_2823 (O_2823,N_28452,N_28026);
or UO_2824 (O_2824,N_28505,N_29354);
and UO_2825 (O_2825,N_27469,N_29439);
nand UO_2826 (O_2826,N_29775,N_29559);
nand UO_2827 (O_2827,N_28426,N_27764);
or UO_2828 (O_2828,N_28731,N_27412);
nor UO_2829 (O_2829,N_29100,N_28697);
and UO_2830 (O_2830,N_28068,N_28597);
nand UO_2831 (O_2831,N_29088,N_29746);
nand UO_2832 (O_2832,N_29888,N_27603);
nor UO_2833 (O_2833,N_29983,N_29676);
nor UO_2834 (O_2834,N_27752,N_29076);
nand UO_2835 (O_2835,N_28745,N_28884);
xor UO_2836 (O_2836,N_27337,N_28235);
or UO_2837 (O_2837,N_28131,N_28648);
nand UO_2838 (O_2838,N_27057,N_28781);
or UO_2839 (O_2839,N_28672,N_28851);
nand UO_2840 (O_2840,N_27520,N_29385);
nor UO_2841 (O_2841,N_28602,N_29975);
and UO_2842 (O_2842,N_27532,N_29900);
or UO_2843 (O_2843,N_28317,N_28215);
nor UO_2844 (O_2844,N_28611,N_28170);
nor UO_2845 (O_2845,N_29568,N_27467);
and UO_2846 (O_2846,N_29592,N_28945);
nand UO_2847 (O_2847,N_27403,N_27274);
and UO_2848 (O_2848,N_29273,N_28148);
nand UO_2849 (O_2849,N_27219,N_27412);
or UO_2850 (O_2850,N_27873,N_27710);
or UO_2851 (O_2851,N_28954,N_29112);
nor UO_2852 (O_2852,N_28389,N_27924);
xnor UO_2853 (O_2853,N_29556,N_28328);
or UO_2854 (O_2854,N_29165,N_28174);
nand UO_2855 (O_2855,N_28951,N_28519);
nand UO_2856 (O_2856,N_27805,N_29537);
nor UO_2857 (O_2857,N_29930,N_27441);
nor UO_2858 (O_2858,N_27336,N_28296);
nor UO_2859 (O_2859,N_28945,N_27424);
nand UO_2860 (O_2860,N_28018,N_27657);
or UO_2861 (O_2861,N_28212,N_27191);
or UO_2862 (O_2862,N_27280,N_28100);
and UO_2863 (O_2863,N_29148,N_27744);
and UO_2864 (O_2864,N_29055,N_28336);
nand UO_2865 (O_2865,N_28958,N_28432);
and UO_2866 (O_2866,N_27923,N_29940);
nor UO_2867 (O_2867,N_27132,N_28858);
nor UO_2868 (O_2868,N_28460,N_29104);
xor UO_2869 (O_2869,N_27457,N_28287);
nor UO_2870 (O_2870,N_29783,N_27261);
nand UO_2871 (O_2871,N_29007,N_29604);
nor UO_2872 (O_2872,N_27357,N_29761);
nor UO_2873 (O_2873,N_28880,N_28055);
nor UO_2874 (O_2874,N_29183,N_29195);
or UO_2875 (O_2875,N_29048,N_28052);
nor UO_2876 (O_2876,N_27884,N_28852);
or UO_2877 (O_2877,N_29997,N_29517);
xnor UO_2878 (O_2878,N_29743,N_28908);
nand UO_2879 (O_2879,N_27704,N_28301);
nor UO_2880 (O_2880,N_28217,N_28345);
and UO_2881 (O_2881,N_27013,N_27227);
and UO_2882 (O_2882,N_28976,N_27983);
or UO_2883 (O_2883,N_27635,N_27563);
nand UO_2884 (O_2884,N_29411,N_29772);
nand UO_2885 (O_2885,N_29262,N_27825);
nand UO_2886 (O_2886,N_27414,N_27655);
or UO_2887 (O_2887,N_29702,N_28951);
and UO_2888 (O_2888,N_28789,N_29322);
or UO_2889 (O_2889,N_29978,N_28279);
or UO_2890 (O_2890,N_29622,N_28207);
nand UO_2891 (O_2891,N_27656,N_27723);
nand UO_2892 (O_2892,N_28588,N_29168);
nor UO_2893 (O_2893,N_28285,N_29427);
or UO_2894 (O_2894,N_27483,N_28364);
nor UO_2895 (O_2895,N_29550,N_29741);
nor UO_2896 (O_2896,N_29206,N_28675);
or UO_2897 (O_2897,N_29028,N_29204);
or UO_2898 (O_2898,N_27287,N_29266);
or UO_2899 (O_2899,N_28420,N_27779);
nor UO_2900 (O_2900,N_29682,N_29799);
nand UO_2901 (O_2901,N_28782,N_28677);
nor UO_2902 (O_2902,N_28851,N_28111);
or UO_2903 (O_2903,N_29672,N_28124);
nand UO_2904 (O_2904,N_28372,N_29294);
and UO_2905 (O_2905,N_28920,N_29562);
xnor UO_2906 (O_2906,N_29349,N_28558);
nand UO_2907 (O_2907,N_28322,N_29072);
nor UO_2908 (O_2908,N_29363,N_28655);
nor UO_2909 (O_2909,N_28847,N_27972);
xnor UO_2910 (O_2910,N_29814,N_27126);
nor UO_2911 (O_2911,N_29702,N_28017);
nor UO_2912 (O_2912,N_28349,N_29978);
or UO_2913 (O_2913,N_29656,N_28415);
nor UO_2914 (O_2914,N_27446,N_29821);
nor UO_2915 (O_2915,N_29996,N_28403);
or UO_2916 (O_2916,N_27158,N_27787);
nor UO_2917 (O_2917,N_29196,N_29497);
or UO_2918 (O_2918,N_27755,N_29131);
nor UO_2919 (O_2919,N_28436,N_27931);
and UO_2920 (O_2920,N_27235,N_28910);
or UO_2921 (O_2921,N_28888,N_28977);
nor UO_2922 (O_2922,N_28832,N_27416);
nand UO_2923 (O_2923,N_29190,N_27182);
or UO_2924 (O_2924,N_27610,N_28237);
xnor UO_2925 (O_2925,N_28705,N_27465);
and UO_2926 (O_2926,N_29646,N_27406);
nor UO_2927 (O_2927,N_27393,N_29364);
or UO_2928 (O_2928,N_29427,N_29314);
and UO_2929 (O_2929,N_27680,N_29704);
and UO_2930 (O_2930,N_27106,N_29532);
and UO_2931 (O_2931,N_27409,N_28478);
xnor UO_2932 (O_2932,N_29251,N_29137);
nand UO_2933 (O_2933,N_28331,N_27800);
nor UO_2934 (O_2934,N_27504,N_27273);
nand UO_2935 (O_2935,N_28200,N_29037);
nor UO_2936 (O_2936,N_28399,N_29849);
nor UO_2937 (O_2937,N_29426,N_27941);
and UO_2938 (O_2938,N_28908,N_29458);
or UO_2939 (O_2939,N_27119,N_27990);
and UO_2940 (O_2940,N_29329,N_27643);
nand UO_2941 (O_2941,N_29072,N_28019);
or UO_2942 (O_2942,N_28593,N_27919);
or UO_2943 (O_2943,N_29556,N_29984);
nand UO_2944 (O_2944,N_28052,N_29396);
nor UO_2945 (O_2945,N_27931,N_28243);
and UO_2946 (O_2946,N_29256,N_29226);
and UO_2947 (O_2947,N_28081,N_27034);
or UO_2948 (O_2948,N_29214,N_28982);
nand UO_2949 (O_2949,N_28764,N_29470);
or UO_2950 (O_2950,N_29607,N_29983);
nand UO_2951 (O_2951,N_27201,N_27221);
or UO_2952 (O_2952,N_27192,N_29676);
or UO_2953 (O_2953,N_29414,N_28696);
nand UO_2954 (O_2954,N_29953,N_27673);
nand UO_2955 (O_2955,N_27539,N_29168);
nor UO_2956 (O_2956,N_28241,N_28777);
xnor UO_2957 (O_2957,N_28650,N_27331);
and UO_2958 (O_2958,N_29158,N_27676);
and UO_2959 (O_2959,N_27771,N_29580);
nor UO_2960 (O_2960,N_27680,N_29166);
nor UO_2961 (O_2961,N_27555,N_29114);
nor UO_2962 (O_2962,N_27664,N_27197);
xnor UO_2963 (O_2963,N_28221,N_29164);
or UO_2964 (O_2964,N_27349,N_29188);
or UO_2965 (O_2965,N_27841,N_28992);
xnor UO_2966 (O_2966,N_27293,N_29250);
and UO_2967 (O_2967,N_27091,N_28568);
nand UO_2968 (O_2968,N_28218,N_28087);
nor UO_2969 (O_2969,N_27412,N_29019);
nor UO_2970 (O_2970,N_29195,N_28357);
nor UO_2971 (O_2971,N_28431,N_27732);
nor UO_2972 (O_2972,N_28939,N_27353);
or UO_2973 (O_2973,N_28838,N_29284);
nor UO_2974 (O_2974,N_29959,N_27861);
nand UO_2975 (O_2975,N_28578,N_27913);
nand UO_2976 (O_2976,N_28524,N_27685);
and UO_2977 (O_2977,N_28959,N_28844);
nand UO_2978 (O_2978,N_27536,N_29973);
nand UO_2979 (O_2979,N_27825,N_28535);
nand UO_2980 (O_2980,N_27116,N_28877);
nand UO_2981 (O_2981,N_28057,N_28990);
xnor UO_2982 (O_2982,N_29170,N_28941);
nor UO_2983 (O_2983,N_27258,N_27379);
and UO_2984 (O_2984,N_27922,N_29532);
nor UO_2985 (O_2985,N_27488,N_28421);
nor UO_2986 (O_2986,N_29292,N_28827);
nand UO_2987 (O_2987,N_28304,N_27616);
and UO_2988 (O_2988,N_28417,N_27589);
and UO_2989 (O_2989,N_28315,N_27682);
nand UO_2990 (O_2990,N_28089,N_27364);
nor UO_2991 (O_2991,N_28676,N_28608);
nand UO_2992 (O_2992,N_28935,N_29065);
nor UO_2993 (O_2993,N_28425,N_27469);
or UO_2994 (O_2994,N_27943,N_28550);
xnor UO_2995 (O_2995,N_27400,N_27222);
or UO_2996 (O_2996,N_27094,N_28506);
or UO_2997 (O_2997,N_27453,N_29779);
or UO_2998 (O_2998,N_27515,N_28597);
and UO_2999 (O_2999,N_28736,N_27948);
nor UO_3000 (O_3000,N_27028,N_27434);
or UO_3001 (O_3001,N_27811,N_29936);
nand UO_3002 (O_3002,N_27633,N_27832);
nand UO_3003 (O_3003,N_29001,N_28202);
or UO_3004 (O_3004,N_29890,N_29504);
nor UO_3005 (O_3005,N_29964,N_29723);
nor UO_3006 (O_3006,N_29120,N_27046);
or UO_3007 (O_3007,N_28693,N_28477);
or UO_3008 (O_3008,N_28115,N_27954);
xnor UO_3009 (O_3009,N_29821,N_28496);
nand UO_3010 (O_3010,N_28334,N_29572);
nand UO_3011 (O_3011,N_27972,N_29005);
or UO_3012 (O_3012,N_28173,N_29752);
xnor UO_3013 (O_3013,N_28555,N_28933);
xor UO_3014 (O_3014,N_29063,N_28872);
nand UO_3015 (O_3015,N_29697,N_28424);
nand UO_3016 (O_3016,N_27371,N_28998);
nand UO_3017 (O_3017,N_29578,N_29527);
or UO_3018 (O_3018,N_29062,N_28380);
nor UO_3019 (O_3019,N_28609,N_29517);
or UO_3020 (O_3020,N_27283,N_28382);
or UO_3021 (O_3021,N_29003,N_27947);
or UO_3022 (O_3022,N_27397,N_28281);
and UO_3023 (O_3023,N_27073,N_29811);
nor UO_3024 (O_3024,N_29605,N_27128);
nor UO_3025 (O_3025,N_28077,N_28637);
and UO_3026 (O_3026,N_27592,N_28867);
or UO_3027 (O_3027,N_28697,N_28274);
or UO_3028 (O_3028,N_27743,N_28259);
and UO_3029 (O_3029,N_27429,N_28257);
or UO_3030 (O_3030,N_27240,N_29317);
nor UO_3031 (O_3031,N_28495,N_28691);
or UO_3032 (O_3032,N_29005,N_27395);
nand UO_3033 (O_3033,N_27594,N_27615);
xor UO_3034 (O_3034,N_29405,N_27543);
xnor UO_3035 (O_3035,N_27341,N_28465);
nand UO_3036 (O_3036,N_28418,N_27632);
nor UO_3037 (O_3037,N_28712,N_29026);
xor UO_3038 (O_3038,N_28510,N_29092);
and UO_3039 (O_3039,N_28481,N_28382);
or UO_3040 (O_3040,N_28052,N_28746);
nor UO_3041 (O_3041,N_27316,N_27980);
nor UO_3042 (O_3042,N_27520,N_28409);
nand UO_3043 (O_3043,N_27664,N_29993);
nor UO_3044 (O_3044,N_28362,N_27686);
nand UO_3045 (O_3045,N_29006,N_29794);
xnor UO_3046 (O_3046,N_29734,N_27591);
and UO_3047 (O_3047,N_28927,N_29527);
nand UO_3048 (O_3048,N_28404,N_27269);
nor UO_3049 (O_3049,N_28380,N_29384);
and UO_3050 (O_3050,N_28982,N_29354);
or UO_3051 (O_3051,N_27201,N_28204);
or UO_3052 (O_3052,N_28067,N_28528);
nand UO_3053 (O_3053,N_29056,N_27850);
nand UO_3054 (O_3054,N_27641,N_28872);
nor UO_3055 (O_3055,N_28197,N_28533);
nand UO_3056 (O_3056,N_29234,N_28114);
and UO_3057 (O_3057,N_28030,N_28197);
nand UO_3058 (O_3058,N_27321,N_27270);
and UO_3059 (O_3059,N_29820,N_27378);
nand UO_3060 (O_3060,N_29396,N_27283);
xor UO_3061 (O_3061,N_27570,N_27436);
or UO_3062 (O_3062,N_28668,N_27422);
nand UO_3063 (O_3063,N_27646,N_29284);
and UO_3064 (O_3064,N_29704,N_28151);
nor UO_3065 (O_3065,N_27642,N_29025);
or UO_3066 (O_3066,N_29643,N_29521);
or UO_3067 (O_3067,N_28583,N_28585);
nand UO_3068 (O_3068,N_28193,N_27634);
nor UO_3069 (O_3069,N_28953,N_29970);
or UO_3070 (O_3070,N_27281,N_29084);
or UO_3071 (O_3071,N_27874,N_29592);
xnor UO_3072 (O_3072,N_28474,N_27337);
nand UO_3073 (O_3073,N_27229,N_28292);
nand UO_3074 (O_3074,N_27816,N_29044);
nor UO_3075 (O_3075,N_29001,N_28855);
or UO_3076 (O_3076,N_29977,N_29513);
nor UO_3077 (O_3077,N_28468,N_28285);
nor UO_3078 (O_3078,N_27599,N_29464);
xor UO_3079 (O_3079,N_27249,N_27425);
nand UO_3080 (O_3080,N_28136,N_29898);
or UO_3081 (O_3081,N_29279,N_28106);
nand UO_3082 (O_3082,N_29831,N_27073);
nor UO_3083 (O_3083,N_28819,N_27368);
or UO_3084 (O_3084,N_28779,N_28686);
or UO_3085 (O_3085,N_29918,N_27450);
nand UO_3086 (O_3086,N_29221,N_28181);
nor UO_3087 (O_3087,N_27260,N_29847);
or UO_3088 (O_3088,N_29481,N_29852);
nor UO_3089 (O_3089,N_27371,N_29587);
nor UO_3090 (O_3090,N_29141,N_27721);
and UO_3091 (O_3091,N_29089,N_28128);
or UO_3092 (O_3092,N_27552,N_28150);
and UO_3093 (O_3093,N_27380,N_28624);
nand UO_3094 (O_3094,N_27521,N_29276);
nor UO_3095 (O_3095,N_28855,N_28112);
and UO_3096 (O_3096,N_28903,N_27639);
xnor UO_3097 (O_3097,N_28802,N_29547);
and UO_3098 (O_3098,N_29265,N_29088);
nand UO_3099 (O_3099,N_27149,N_27883);
nor UO_3100 (O_3100,N_28611,N_29954);
and UO_3101 (O_3101,N_28628,N_27663);
nor UO_3102 (O_3102,N_27381,N_28704);
or UO_3103 (O_3103,N_27895,N_27690);
xnor UO_3104 (O_3104,N_28935,N_27667);
nand UO_3105 (O_3105,N_29869,N_27072);
nand UO_3106 (O_3106,N_28974,N_27035);
nand UO_3107 (O_3107,N_28139,N_29664);
xor UO_3108 (O_3108,N_28988,N_27380);
nand UO_3109 (O_3109,N_28262,N_27727);
nor UO_3110 (O_3110,N_27128,N_29289);
nor UO_3111 (O_3111,N_28827,N_28988);
or UO_3112 (O_3112,N_28464,N_27167);
nor UO_3113 (O_3113,N_29654,N_27360);
and UO_3114 (O_3114,N_29215,N_27264);
nor UO_3115 (O_3115,N_29716,N_27114);
nor UO_3116 (O_3116,N_28233,N_29090);
nor UO_3117 (O_3117,N_28448,N_28222);
or UO_3118 (O_3118,N_28635,N_27550);
xor UO_3119 (O_3119,N_27953,N_29777);
or UO_3120 (O_3120,N_28514,N_28634);
nor UO_3121 (O_3121,N_29673,N_28721);
nor UO_3122 (O_3122,N_28801,N_27344);
nor UO_3123 (O_3123,N_29938,N_29799);
and UO_3124 (O_3124,N_27001,N_27329);
nand UO_3125 (O_3125,N_29545,N_27883);
nor UO_3126 (O_3126,N_28453,N_27644);
nand UO_3127 (O_3127,N_27940,N_27622);
and UO_3128 (O_3128,N_27109,N_29344);
or UO_3129 (O_3129,N_27641,N_27333);
nand UO_3130 (O_3130,N_27862,N_29917);
nor UO_3131 (O_3131,N_28742,N_28797);
and UO_3132 (O_3132,N_27324,N_28010);
or UO_3133 (O_3133,N_27701,N_28504);
or UO_3134 (O_3134,N_28098,N_28408);
and UO_3135 (O_3135,N_27786,N_27795);
nand UO_3136 (O_3136,N_27472,N_27070);
nand UO_3137 (O_3137,N_27813,N_29677);
nand UO_3138 (O_3138,N_27205,N_27734);
nand UO_3139 (O_3139,N_28091,N_27710);
nand UO_3140 (O_3140,N_29083,N_28187);
or UO_3141 (O_3141,N_28623,N_28376);
xor UO_3142 (O_3142,N_28499,N_27178);
nand UO_3143 (O_3143,N_28105,N_29209);
or UO_3144 (O_3144,N_28087,N_29790);
and UO_3145 (O_3145,N_28449,N_27823);
or UO_3146 (O_3146,N_29493,N_28373);
and UO_3147 (O_3147,N_28099,N_29690);
or UO_3148 (O_3148,N_29266,N_27537);
and UO_3149 (O_3149,N_28494,N_27501);
xor UO_3150 (O_3150,N_28971,N_28756);
xnor UO_3151 (O_3151,N_27343,N_27805);
and UO_3152 (O_3152,N_28068,N_29603);
nor UO_3153 (O_3153,N_29278,N_29227);
or UO_3154 (O_3154,N_27140,N_27995);
and UO_3155 (O_3155,N_29753,N_28437);
nand UO_3156 (O_3156,N_29958,N_28838);
nand UO_3157 (O_3157,N_28869,N_29337);
or UO_3158 (O_3158,N_29754,N_28571);
xnor UO_3159 (O_3159,N_27735,N_28990);
nand UO_3160 (O_3160,N_27146,N_29988);
and UO_3161 (O_3161,N_28485,N_27228);
and UO_3162 (O_3162,N_29837,N_28871);
and UO_3163 (O_3163,N_29148,N_28753);
nor UO_3164 (O_3164,N_27037,N_28714);
or UO_3165 (O_3165,N_27819,N_27075);
nand UO_3166 (O_3166,N_28432,N_28003);
and UO_3167 (O_3167,N_28809,N_27848);
nor UO_3168 (O_3168,N_29215,N_29568);
nor UO_3169 (O_3169,N_27752,N_29604);
or UO_3170 (O_3170,N_29571,N_29730);
xor UO_3171 (O_3171,N_28081,N_27516);
and UO_3172 (O_3172,N_28464,N_27529);
nand UO_3173 (O_3173,N_28809,N_28515);
nand UO_3174 (O_3174,N_29888,N_28170);
nand UO_3175 (O_3175,N_28425,N_29048);
or UO_3176 (O_3176,N_27523,N_28078);
or UO_3177 (O_3177,N_28961,N_27796);
and UO_3178 (O_3178,N_29137,N_29891);
and UO_3179 (O_3179,N_27742,N_27226);
xnor UO_3180 (O_3180,N_29869,N_29595);
or UO_3181 (O_3181,N_29272,N_28997);
nor UO_3182 (O_3182,N_27439,N_29313);
nor UO_3183 (O_3183,N_27033,N_28677);
nor UO_3184 (O_3184,N_28945,N_29760);
nand UO_3185 (O_3185,N_27779,N_29883);
and UO_3186 (O_3186,N_29602,N_28649);
nor UO_3187 (O_3187,N_27138,N_29688);
and UO_3188 (O_3188,N_29011,N_28162);
and UO_3189 (O_3189,N_28006,N_27542);
nor UO_3190 (O_3190,N_29297,N_29169);
nor UO_3191 (O_3191,N_29851,N_28806);
and UO_3192 (O_3192,N_27274,N_28669);
nand UO_3193 (O_3193,N_27156,N_29368);
and UO_3194 (O_3194,N_29207,N_27047);
and UO_3195 (O_3195,N_27939,N_28863);
nor UO_3196 (O_3196,N_27253,N_27348);
or UO_3197 (O_3197,N_27590,N_28439);
or UO_3198 (O_3198,N_28862,N_27593);
nand UO_3199 (O_3199,N_29826,N_27358);
and UO_3200 (O_3200,N_29075,N_27604);
nand UO_3201 (O_3201,N_29375,N_27073);
and UO_3202 (O_3202,N_27397,N_27077);
or UO_3203 (O_3203,N_28489,N_29618);
and UO_3204 (O_3204,N_28206,N_28024);
or UO_3205 (O_3205,N_28403,N_28237);
and UO_3206 (O_3206,N_28721,N_29955);
and UO_3207 (O_3207,N_27146,N_29128);
or UO_3208 (O_3208,N_29074,N_27284);
nand UO_3209 (O_3209,N_28781,N_28423);
and UO_3210 (O_3210,N_29393,N_28888);
or UO_3211 (O_3211,N_28264,N_29379);
nand UO_3212 (O_3212,N_28910,N_27581);
xor UO_3213 (O_3213,N_29908,N_29540);
xor UO_3214 (O_3214,N_29073,N_28723);
and UO_3215 (O_3215,N_27960,N_28503);
nor UO_3216 (O_3216,N_27712,N_27686);
nand UO_3217 (O_3217,N_27445,N_28535);
nand UO_3218 (O_3218,N_27391,N_27277);
and UO_3219 (O_3219,N_29188,N_27442);
nor UO_3220 (O_3220,N_29814,N_27244);
xnor UO_3221 (O_3221,N_29092,N_29503);
nand UO_3222 (O_3222,N_29984,N_27408);
nor UO_3223 (O_3223,N_29571,N_27432);
xor UO_3224 (O_3224,N_29754,N_27289);
nor UO_3225 (O_3225,N_27227,N_28673);
nor UO_3226 (O_3226,N_29880,N_27318);
nor UO_3227 (O_3227,N_28228,N_29211);
nand UO_3228 (O_3228,N_28379,N_28358);
or UO_3229 (O_3229,N_27874,N_28029);
nor UO_3230 (O_3230,N_28243,N_28706);
nor UO_3231 (O_3231,N_29558,N_27880);
and UO_3232 (O_3232,N_29290,N_28861);
and UO_3233 (O_3233,N_29113,N_27361);
or UO_3234 (O_3234,N_27948,N_28542);
or UO_3235 (O_3235,N_27949,N_27134);
nor UO_3236 (O_3236,N_27400,N_27253);
nand UO_3237 (O_3237,N_27657,N_28078);
xor UO_3238 (O_3238,N_28262,N_27914);
or UO_3239 (O_3239,N_28907,N_29430);
and UO_3240 (O_3240,N_27714,N_29547);
and UO_3241 (O_3241,N_28804,N_29329);
and UO_3242 (O_3242,N_27000,N_29801);
nor UO_3243 (O_3243,N_27643,N_28054);
nand UO_3244 (O_3244,N_27545,N_28644);
xnor UO_3245 (O_3245,N_29510,N_28435);
or UO_3246 (O_3246,N_27161,N_28305);
nor UO_3247 (O_3247,N_28575,N_27133);
nor UO_3248 (O_3248,N_29598,N_27758);
xor UO_3249 (O_3249,N_28362,N_27496);
or UO_3250 (O_3250,N_27873,N_29189);
nor UO_3251 (O_3251,N_27062,N_28589);
or UO_3252 (O_3252,N_29613,N_28463);
xnor UO_3253 (O_3253,N_29638,N_28745);
or UO_3254 (O_3254,N_29073,N_27521);
nand UO_3255 (O_3255,N_27167,N_27114);
and UO_3256 (O_3256,N_27082,N_27629);
and UO_3257 (O_3257,N_28157,N_29097);
nor UO_3258 (O_3258,N_28612,N_28414);
nor UO_3259 (O_3259,N_27450,N_29181);
and UO_3260 (O_3260,N_27134,N_28546);
or UO_3261 (O_3261,N_27567,N_27444);
nor UO_3262 (O_3262,N_27933,N_28639);
or UO_3263 (O_3263,N_27950,N_28173);
or UO_3264 (O_3264,N_29451,N_28873);
xnor UO_3265 (O_3265,N_29294,N_27875);
and UO_3266 (O_3266,N_29373,N_29158);
nor UO_3267 (O_3267,N_27090,N_28932);
or UO_3268 (O_3268,N_29961,N_29097);
nor UO_3269 (O_3269,N_28367,N_29110);
or UO_3270 (O_3270,N_28531,N_28652);
nor UO_3271 (O_3271,N_29402,N_27791);
nand UO_3272 (O_3272,N_28873,N_28478);
and UO_3273 (O_3273,N_27011,N_28536);
or UO_3274 (O_3274,N_27162,N_28930);
nor UO_3275 (O_3275,N_28080,N_28025);
and UO_3276 (O_3276,N_28527,N_28649);
and UO_3277 (O_3277,N_27862,N_29181);
xnor UO_3278 (O_3278,N_27097,N_28720);
or UO_3279 (O_3279,N_29353,N_28667);
or UO_3280 (O_3280,N_29856,N_27648);
and UO_3281 (O_3281,N_29083,N_28288);
xnor UO_3282 (O_3282,N_27608,N_28460);
nand UO_3283 (O_3283,N_29346,N_29285);
nand UO_3284 (O_3284,N_28697,N_27781);
nand UO_3285 (O_3285,N_27967,N_29408);
or UO_3286 (O_3286,N_29524,N_27997);
nand UO_3287 (O_3287,N_27839,N_28738);
or UO_3288 (O_3288,N_29130,N_28701);
nor UO_3289 (O_3289,N_29543,N_29289);
and UO_3290 (O_3290,N_28807,N_27331);
nor UO_3291 (O_3291,N_28923,N_27539);
or UO_3292 (O_3292,N_28924,N_29215);
and UO_3293 (O_3293,N_27508,N_28894);
nand UO_3294 (O_3294,N_28561,N_28663);
and UO_3295 (O_3295,N_29997,N_29856);
nor UO_3296 (O_3296,N_28133,N_29964);
and UO_3297 (O_3297,N_27633,N_27672);
xnor UO_3298 (O_3298,N_29823,N_27011);
nor UO_3299 (O_3299,N_28279,N_27592);
and UO_3300 (O_3300,N_29695,N_27523);
and UO_3301 (O_3301,N_27604,N_28958);
or UO_3302 (O_3302,N_27608,N_28674);
nor UO_3303 (O_3303,N_29981,N_28793);
xnor UO_3304 (O_3304,N_29644,N_28352);
nand UO_3305 (O_3305,N_28379,N_28633);
and UO_3306 (O_3306,N_29811,N_29439);
nor UO_3307 (O_3307,N_27292,N_28414);
and UO_3308 (O_3308,N_28433,N_27418);
or UO_3309 (O_3309,N_29900,N_28977);
xnor UO_3310 (O_3310,N_28555,N_29194);
and UO_3311 (O_3311,N_27781,N_29097);
and UO_3312 (O_3312,N_27722,N_29896);
and UO_3313 (O_3313,N_29831,N_27365);
and UO_3314 (O_3314,N_29048,N_29244);
nand UO_3315 (O_3315,N_29033,N_28705);
and UO_3316 (O_3316,N_29552,N_27280);
and UO_3317 (O_3317,N_27155,N_27966);
or UO_3318 (O_3318,N_29158,N_27574);
nor UO_3319 (O_3319,N_28219,N_29833);
nand UO_3320 (O_3320,N_29196,N_27595);
nor UO_3321 (O_3321,N_29158,N_29971);
or UO_3322 (O_3322,N_27388,N_29863);
xor UO_3323 (O_3323,N_29722,N_27715);
or UO_3324 (O_3324,N_28236,N_29462);
nor UO_3325 (O_3325,N_27538,N_28679);
or UO_3326 (O_3326,N_29778,N_28131);
nand UO_3327 (O_3327,N_29703,N_29820);
nor UO_3328 (O_3328,N_28693,N_27147);
and UO_3329 (O_3329,N_27167,N_28087);
and UO_3330 (O_3330,N_28186,N_29483);
nor UO_3331 (O_3331,N_29493,N_29583);
nor UO_3332 (O_3332,N_27438,N_29112);
nand UO_3333 (O_3333,N_27509,N_29907);
nor UO_3334 (O_3334,N_29346,N_28202);
nand UO_3335 (O_3335,N_28519,N_28182);
xor UO_3336 (O_3336,N_27283,N_29399);
and UO_3337 (O_3337,N_29284,N_28434);
nor UO_3338 (O_3338,N_29656,N_28769);
nand UO_3339 (O_3339,N_28922,N_28165);
or UO_3340 (O_3340,N_29460,N_27378);
and UO_3341 (O_3341,N_29375,N_28572);
nor UO_3342 (O_3342,N_27294,N_29182);
or UO_3343 (O_3343,N_29226,N_27967);
nor UO_3344 (O_3344,N_29127,N_29014);
nor UO_3345 (O_3345,N_28578,N_29715);
and UO_3346 (O_3346,N_28867,N_28929);
and UO_3347 (O_3347,N_29143,N_29908);
nand UO_3348 (O_3348,N_29483,N_28135);
and UO_3349 (O_3349,N_29512,N_29111);
or UO_3350 (O_3350,N_29866,N_28379);
and UO_3351 (O_3351,N_29846,N_28949);
xnor UO_3352 (O_3352,N_27402,N_29137);
and UO_3353 (O_3353,N_27062,N_27588);
nor UO_3354 (O_3354,N_28525,N_27611);
and UO_3355 (O_3355,N_28736,N_28651);
nor UO_3356 (O_3356,N_28780,N_28833);
nor UO_3357 (O_3357,N_27982,N_27856);
or UO_3358 (O_3358,N_28621,N_28829);
nor UO_3359 (O_3359,N_27276,N_28911);
or UO_3360 (O_3360,N_28305,N_29211);
xnor UO_3361 (O_3361,N_29697,N_28560);
nor UO_3362 (O_3362,N_27456,N_28523);
or UO_3363 (O_3363,N_29457,N_28306);
and UO_3364 (O_3364,N_29502,N_29644);
and UO_3365 (O_3365,N_27559,N_28037);
and UO_3366 (O_3366,N_28633,N_28821);
nand UO_3367 (O_3367,N_28811,N_28279);
and UO_3368 (O_3368,N_27677,N_28288);
xor UO_3369 (O_3369,N_27918,N_27074);
nand UO_3370 (O_3370,N_28851,N_29291);
nand UO_3371 (O_3371,N_29559,N_28093);
or UO_3372 (O_3372,N_29256,N_28235);
nand UO_3373 (O_3373,N_27161,N_29949);
xor UO_3374 (O_3374,N_28890,N_27496);
nor UO_3375 (O_3375,N_28429,N_29565);
nand UO_3376 (O_3376,N_28891,N_29357);
nor UO_3377 (O_3377,N_27674,N_29046);
nand UO_3378 (O_3378,N_27015,N_28162);
and UO_3379 (O_3379,N_29721,N_28402);
nand UO_3380 (O_3380,N_27090,N_29702);
or UO_3381 (O_3381,N_29934,N_28657);
nand UO_3382 (O_3382,N_28443,N_28856);
and UO_3383 (O_3383,N_27093,N_27702);
or UO_3384 (O_3384,N_29934,N_27335);
and UO_3385 (O_3385,N_29137,N_27250);
or UO_3386 (O_3386,N_29792,N_29549);
nand UO_3387 (O_3387,N_28229,N_28611);
or UO_3388 (O_3388,N_27656,N_28651);
nor UO_3389 (O_3389,N_27320,N_29315);
and UO_3390 (O_3390,N_28608,N_29890);
or UO_3391 (O_3391,N_28762,N_27267);
nor UO_3392 (O_3392,N_28911,N_27230);
and UO_3393 (O_3393,N_28768,N_28288);
and UO_3394 (O_3394,N_28644,N_28035);
nand UO_3395 (O_3395,N_27029,N_29262);
nor UO_3396 (O_3396,N_27755,N_28360);
or UO_3397 (O_3397,N_27852,N_28520);
and UO_3398 (O_3398,N_27284,N_27695);
nor UO_3399 (O_3399,N_28543,N_27462);
and UO_3400 (O_3400,N_28611,N_28855);
and UO_3401 (O_3401,N_29138,N_29456);
or UO_3402 (O_3402,N_29457,N_29622);
nand UO_3403 (O_3403,N_27379,N_29997);
and UO_3404 (O_3404,N_27448,N_29206);
nand UO_3405 (O_3405,N_29137,N_27422);
nor UO_3406 (O_3406,N_27002,N_28694);
nor UO_3407 (O_3407,N_28067,N_27550);
nor UO_3408 (O_3408,N_27864,N_27083);
nand UO_3409 (O_3409,N_28606,N_28401);
nor UO_3410 (O_3410,N_27255,N_28283);
and UO_3411 (O_3411,N_28972,N_29865);
and UO_3412 (O_3412,N_28022,N_27877);
and UO_3413 (O_3413,N_27564,N_28116);
nand UO_3414 (O_3414,N_27363,N_27132);
and UO_3415 (O_3415,N_28757,N_28499);
or UO_3416 (O_3416,N_27274,N_29566);
or UO_3417 (O_3417,N_29322,N_28020);
nor UO_3418 (O_3418,N_28891,N_29662);
xor UO_3419 (O_3419,N_29603,N_28558);
or UO_3420 (O_3420,N_27347,N_27082);
and UO_3421 (O_3421,N_29487,N_27109);
and UO_3422 (O_3422,N_27373,N_29366);
nor UO_3423 (O_3423,N_27932,N_27931);
nor UO_3424 (O_3424,N_27110,N_29492);
nand UO_3425 (O_3425,N_28218,N_29632);
xnor UO_3426 (O_3426,N_27723,N_27647);
or UO_3427 (O_3427,N_29664,N_28668);
and UO_3428 (O_3428,N_28451,N_29958);
nand UO_3429 (O_3429,N_27154,N_29199);
nor UO_3430 (O_3430,N_29123,N_29622);
and UO_3431 (O_3431,N_27054,N_28811);
and UO_3432 (O_3432,N_28500,N_28840);
xnor UO_3433 (O_3433,N_29751,N_27011);
nand UO_3434 (O_3434,N_28816,N_27595);
and UO_3435 (O_3435,N_29425,N_28644);
xor UO_3436 (O_3436,N_29114,N_27159);
and UO_3437 (O_3437,N_29635,N_29138);
xnor UO_3438 (O_3438,N_29436,N_27565);
nor UO_3439 (O_3439,N_27793,N_27198);
or UO_3440 (O_3440,N_29715,N_29349);
nand UO_3441 (O_3441,N_28770,N_28833);
xnor UO_3442 (O_3442,N_27182,N_27694);
nor UO_3443 (O_3443,N_29594,N_29086);
nand UO_3444 (O_3444,N_29182,N_27305);
nand UO_3445 (O_3445,N_28474,N_27983);
nor UO_3446 (O_3446,N_27601,N_29713);
or UO_3447 (O_3447,N_28688,N_29357);
nand UO_3448 (O_3448,N_28089,N_27214);
or UO_3449 (O_3449,N_28552,N_27842);
nand UO_3450 (O_3450,N_27784,N_28978);
nor UO_3451 (O_3451,N_27128,N_27487);
or UO_3452 (O_3452,N_28039,N_27676);
xor UO_3453 (O_3453,N_28658,N_28831);
nor UO_3454 (O_3454,N_27074,N_27961);
or UO_3455 (O_3455,N_29062,N_29365);
and UO_3456 (O_3456,N_28115,N_29873);
and UO_3457 (O_3457,N_28137,N_27802);
or UO_3458 (O_3458,N_27776,N_29106);
or UO_3459 (O_3459,N_28606,N_28182);
and UO_3460 (O_3460,N_28136,N_28827);
xor UO_3461 (O_3461,N_27432,N_28626);
and UO_3462 (O_3462,N_28869,N_29400);
nand UO_3463 (O_3463,N_29473,N_27841);
xnor UO_3464 (O_3464,N_27280,N_28421);
or UO_3465 (O_3465,N_27507,N_28159);
and UO_3466 (O_3466,N_29983,N_28893);
or UO_3467 (O_3467,N_27848,N_27893);
nor UO_3468 (O_3468,N_29794,N_29675);
and UO_3469 (O_3469,N_27977,N_29048);
xor UO_3470 (O_3470,N_28490,N_29186);
and UO_3471 (O_3471,N_29609,N_28727);
or UO_3472 (O_3472,N_27807,N_29349);
and UO_3473 (O_3473,N_28323,N_29248);
xnor UO_3474 (O_3474,N_27393,N_29707);
xor UO_3475 (O_3475,N_28741,N_29628);
and UO_3476 (O_3476,N_29287,N_28477);
and UO_3477 (O_3477,N_27905,N_29133);
and UO_3478 (O_3478,N_28560,N_27634);
nand UO_3479 (O_3479,N_29925,N_28564);
and UO_3480 (O_3480,N_28170,N_28445);
or UO_3481 (O_3481,N_29149,N_28503);
nor UO_3482 (O_3482,N_27677,N_28879);
or UO_3483 (O_3483,N_28888,N_29752);
and UO_3484 (O_3484,N_28942,N_29259);
and UO_3485 (O_3485,N_27402,N_28397);
xnor UO_3486 (O_3486,N_28012,N_29019);
xor UO_3487 (O_3487,N_29487,N_29739);
and UO_3488 (O_3488,N_28562,N_29858);
nand UO_3489 (O_3489,N_27355,N_29462);
or UO_3490 (O_3490,N_29246,N_28937);
nand UO_3491 (O_3491,N_28538,N_29481);
nor UO_3492 (O_3492,N_27115,N_29119);
nand UO_3493 (O_3493,N_27686,N_29079);
xor UO_3494 (O_3494,N_29984,N_27247);
or UO_3495 (O_3495,N_29395,N_28318);
nor UO_3496 (O_3496,N_29804,N_27339);
nand UO_3497 (O_3497,N_28279,N_27497);
and UO_3498 (O_3498,N_29689,N_28099);
and UO_3499 (O_3499,N_29227,N_28097);
endmodule