module basic_1000_10000_1500_5_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_360,In_721);
nor U1 (N_1,In_694,In_455);
or U2 (N_2,In_90,In_792);
nor U3 (N_3,In_927,In_991);
or U4 (N_4,In_590,In_936);
nor U5 (N_5,In_237,In_881);
or U6 (N_6,In_28,In_373);
and U7 (N_7,In_942,In_262);
nand U8 (N_8,In_492,In_950);
or U9 (N_9,In_122,In_918);
and U10 (N_10,In_720,In_634);
nor U11 (N_11,In_645,In_862);
and U12 (N_12,In_248,In_3);
nor U13 (N_13,In_616,In_632);
nand U14 (N_14,In_808,In_739);
nor U15 (N_15,In_929,In_718);
nand U16 (N_16,In_615,In_199);
nand U17 (N_17,In_993,In_368);
or U18 (N_18,In_555,In_635);
or U19 (N_19,In_217,In_656);
and U20 (N_20,In_556,In_323);
nand U21 (N_21,In_767,In_218);
nor U22 (N_22,In_160,In_740);
and U23 (N_23,In_290,In_200);
and U24 (N_24,In_416,In_981);
nor U25 (N_25,In_866,In_236);
nand U26 (N_26,In_195,In_975);
nand U27 (N_27,In_855,In_267);
and U28 (N_28,In_971,In_994);
or U29 (N_29,In_435,In_520);
or U30 (N_30,In_388,In_321);
or U31 (N_31,In_679,In_289);
or U32 (N_32,In_507,In_148);
and U33 (N_33,In_513,In_329);
nand U34 (N_34,In_370,In_81);
and U35 (N_35,In_36,In_6);
nor U36 (N_36,In_755,In_444);
nor U37 (N_37,In_749,In_146);
xor U38 (N_38,In_805,In_654);
nand U39 (N_39,In_559,In_502);
or U40 (N_40,In_371,In_608);
nor U41 (N_41,In_754,In_491);
or U42 (N_42,In_191,In_98);
nand U43 (N_43,In_980,In_358);
or U44 (N_44,In_79,In_563);
or U45 (N_45,In_147,In_274);
nor U46 (N_46,In_481,In_397);
or U47 (N_47,In_834,In_110);
and U48 (N_48,In_383,In_134);
and U49 (N_49,In_87,In_51);
nand U50 (N_50,In_803,In_607);
and U51 (N_51,In_965,In_489);
and U52 (N_52,In_457,In_16);
or U53 (N_53,In_220,In_858);
xor U54 (N_54,In_784,In_103);
and U55 (N_55,In_104,In_505);
or U56 (N_56,In_546,In_63);
or U57 (N_57,In_888,In_677);
xor U58 (N_58,In_377,In_156);
or U59 (N_59,In_990,In_265);
and U60 (N_60,In_209,In_791);
nor U61 (N_61,In_390,In_964);
nor U62 (N_62,In_339,In_931);
nand U63 (N_63,In_818,In_72);
xnor U64 (N_64,In_362,In_509);
and U65 (N_65,In_182,In_292);
or U66 (N_66,In_838,In_252);
nand U67 (N_67,In_700,In_954);
and U68 (N_68,In_437,In_347);
and U69 (N_69,In_259,In_982);
and U70 (N_70,In_37,In_427);
nor U71 (N_71,In_447,In_899);
nand U72 (N_72,In_144,In_807);
nor U73 (N_73,In_42,In_526);
nand U74 (N_74,In_958,In_553);
and U75 (N_75,In_610,In_790);
nand U76 (N_76,In_298,In_760);
xor U77 (N_77,In_583,In_568);
nor U78 (N_78,In_744,In_227);
nor U79 (N_79,In_500,In_585);
or U80 (N_80,In_295,In_841);
nand U81 (N_81,In_810,In_666);
or U82 (N_82,In_955,In_598);
nand U83 (N_83,In_158,In_973);
nand U84 (N_84,In_935,In_466);
and U85 (N_85,In_470,In_854);
or U86 (N_86,In_892,In_743);
nand U87 (N_87,In_839,In_727);
nand U88 (N_88,In_562,In_83);
nand U89 (N_89,In_450,In_787);
nor U90 (N_90,In_917,In_658);
nor U91 (N_91,In_281,In_877);
nand U92 (N_92,In_864,In_401);
nor U93 (N_93,In_573,In_452);
nand U94 (N_94,In_746,In_748);
nor U95 (N_95,In_602,In_552);
and U96 (N_96,In_359,In_436);
nand U97 (N_97,In_208,In_531);
nor U98 (N_98,In_843,In_233);
or U99 (N_99,In_959,In_712);
nor U100 (N_100,In_123,In_575);
nor U101 (N_101,In_27,In_883);
nor U102 (N_102,In_86,In_245);
nor U103 (N_103,In_693,In_8);
or U104 (N_104,In_827,In_326);
and U105 (N_105,In_972,In_882);
nor U106 (N_106,In_223,In_544);
xnor U107 (N_107,In_714,In_938);
and U108 (N_108,In_558,In_974);
and U109 (N_109,In_212,In_17);
and U110 (N_110,In_317,In_617);
or U111 (N_111,In_196,In_78);
and U112 (N_112,In_89,In_340);
nor U113 (N_113,In_478,In_823);
nor U114 (N_114,In_33,In_282);
nor U115 (N_115,In_893,In_957);
and U116 (N_116,In_0,In_538);
nor U117 (N_117,In_372,In_438);
or U118 (N_118,In_557,In_922);
nand U119 (N_119,In_809,In_53);
or U120 (N_120,In_723,In_742);
nand U121 (N_121,In_701,In_511);
and U122 (N_122,In_462,In_93);
or U123 (N_123,In_382,In_345);
and U124 (N_124,In_667,In_247);
and U125 (N_125,In_570,In_409);
or U126 (N_126,In_706,In_73);
and U127 (N_127,In_924,In_327);
or U128 (N_128,In_225,In_226);
nor U129 (N_129,In_2,In_750);
xor U130 (N_130,In_205,In_966);
nand U131 (N_131,In_756,In_782);
nand U132 (N_132,In_9,In_822);
or U133 (N_133,In_312,In_198);
nand U134 (N_134,In_774,In_770);
nand U135 (N_135,In_149,In_571);
nand U136 (N_136,In_905,In_771);
nor U137 (N_137,In_629,In_386);
or U138 (N_138,In_947,In_896);
or U139 (N_139,In_670,In_643);
nor U140 (N_140,In_765,In_514);
nor U141 (N_141,In_745,In_357);
nand U142 (N_142,In_167,In_525);
nand U143 (N_143,In_288,In_441);
nand U144 (N_144,In_92,In_941);
and U145 (N_145,In_126,In_630);
or U146 (N_146,In_296,In_496);
nand U147 (N_147,In_460,In_330);
xor U148 (N_148,In_547,In_343);
nand U149 (N_149,In_389,In_829);
nand U150 (N_150,In_423,In_846);
nor U151 (N_151,In_474,In_676);
and U152 (N_152,In_836,In_703);
or U153 (N_153,In_94,In_952);
xor U154 (N_154,In_828,In_678);
and U155 (N_155,In_166,In_400);
xor U156 (N_156,In_130,In_406);
or U157 (N_157,In_203,In_914);
and U158 (N_158,In_934,In_946);
nor U159 (N_159,In_453,In_251);
or U160 (N_160,In_367,In_915);
and U161 (N_161,In_550,In_683);
and U162 (N_162,In_5,In_324);
nand U163 (N_163,In_420,In_532);
or U164 (N_164,In_270,In_354);
or U165 (N_165,In_80,In_66);
and U166 (N_166,In_395,In_876);
or U167 (N_167,In_219,In_417);
and U168 (N_168,In_257,In_762);
or U169 (N_169,In_54,In_169);
or U170 (N_170,In_878,In_434);
nand U171 (N_171,In_926,In_495);
nand U172 (N_172,In_768,In_242);
or U173 (N_173,In_99,In_897);
and U174 (N_174,In_900,In_937);
and U175 (N_175,In_136,In_908);
and U176 (N_176,In_303,In_535);
nor U177 (N_177,In_232,In_987);
nand U178 (N_178,In_599,In_832);
nand U179 (N_179,In_651,In_962);
and U180 (N_180,In_459,In_685);
or U181 (N_181,In_675,In_164);
nand U182 (N_182,In_341,In_172);
nor U183 (N_183,In_369,In_884);
nor U184 (N_184,In_800,In_471);
nor U185 (N_185,In_439,In_465);
or U186 (N_186,In_43,In_300);
or U187 (N_187,In_185,In_969);
or U188 (N_188,In_680,In_766);
nand U189 (N_189,In_793,In_361);
nor U190 (N_190,In_837,In_688);
or U191 (N_191,In_190,In_34);
or U192 (N_192,In_432,In_414);
nand U193 (N_193,In_68,In_118);
nor U194 (N_194,In_886,In_485);
or U195 (N_195,In_816,In_879);
xnor U196 (N_196,In_636,In_761);
nor U197 (N_197,In_61,In_398);
nor U198 (N_198,In_736,In_596);
nand U199 (N_199,In_111,In_308);
xnor U200 (N_200,In_569,In_258);
nand U201 (N_201,In_549,In_19);
and U202 (N_202,In_426,In_45);
and U203 (N_203,In_25,In_293);
nand U204 (N_204,In_348,In_530);
and U205 (N_205,In_566,In_777);
and U206 (N_206,In_71,In_625);
nor U207 (N_207,In_333,In_729);
and U208 (N_208,In_309,In_527);
nand U209 (N_209,In_261,In_517);
nand U210 (N_210,In_405,In_229);
nand U211 (N_211,In_758,In_819);
nor U212 (N_212,In_631,In_109);
or U213 (N_213,In_673,In_264);
nor U214 (N_214,In_366,In_451);
nor U215 (N_215,In_528,In_804);
nand U216 (N_216,In_814,In_129);
and U217 (N_217,In_699,In_101);
or U218 (N_218,In_415,In_230);
nand U219 (N_219,In_584,In_131);
nand U220 (N_220,In_194,In_88);
and U221 (N_221,In_446,In_458);
nand U222 (N_222,In_375,In_895);
and U223 (N_223,In_722,In_454);
nand U224 (N_224,In_778,In_662);
or U225 (N_225,In_222,In_997);
nor U226 (N_226,In_363,In_320);
nand U227 (N_227,In_968,In_337);
nand U228 (N_228,In_487,In_889);
xnor U229 (N_229,In_404,In_567);
and U230 (N_230,In_425,In_216);
nand U231 (N_231,In_275,In_757);
and U232 (N_232,In_15,In_865);
nand U233 (N_233,In_413,In_91);
nor U234 (N_234,In_859,In_238);
and U235 (N_235,In_40,In_910);
nand U236 (N_236,In_789,In_812);
or U237 (N_237,In_603,In_112);
and U238 (N_238,In_263,In_463);
nand U239 (N_239,In_477,In_518);
and U240 (N_240,In_687,In_875);
or U241 (N_241,In_572,In_84);
or U242 (N_242,In_76,In_387);
nor U243 (N_243,In_243,In_860);
nor U244 (N_244,In_7,In_665);
nor U245 (N_245,In_633,In_543);
nor U246 (N_246,In_898,In_904);
and U247 (N_247,In_923,In_175);
and U248 (N_248,In_763,In_648);
or U249 (N_249,In_336,In_440);
nor U250 (N_250,In_286,In_23);
xor U251 (N_251,In_856,In_783);
nand U252 (N_252,In_788,In_430);
or U253 (N_253,In_254,In_74);
nand U254 (N_254,In_379,In_649);
nor U255 (N_255,In_276,In_197);
or U256 (N_256,In_921,In_508);
and U257 (N_257,In_142,In_154);
nor U258 (N_258,In_284,In_612);
nor U259 (N_259,In_582,In_621);
nand U260 (N_260,In_497,In_140);
nor U261 (N_261,In_671,In_797);
nor U262 (N_262,In_52,In_796);
and U263 (N_263,In_996,In_695);
and U264 (N_264,In_211,In_874);
and U265 (N_265,In_561,In_418);
and U266 (N_266,In_586,In_737);
and U267 (N_267,In_709,In_85);
nand U268 (N_268,In_861,In_589);
nand U269 (N_269,In_183,In_125);
nand U270 (N_270,In_193,In_912);
or U271 (N_271,In_165,In_995);
nand U272 (N_272,In_717,In_565);
nor U273 (N_273,In_798,In_786);
or U274 (N_274,In_202,In_913);
and U275 (N_275,In_189,In_132);
nand U276 (N_276,In_494,In_176);
or U277 (N_277,In_493,In_143);
and U278 (N_278,In_32,In_732);
or U279 (N_279,In_272,In_332);
nand U280 (N_280,In_920,In_127);
nor U281 (N_281,In_448,In_121);
nand U282 (N_282,In_141,In_313);
or U283 (N_283,In_244,In_719);
nor U284 (N_284,In_322,In_38);
nor U285 (N_285,In_747,In_581);
nand U286 (N_286,In_620,In_668);
and U287 (N_287,In_698,In_138);
or U288 (N_288,In_442,In_759);
nor U289 (N_289,In_128,In_869);
and U290 (N_290,In_619,In_419);
nand U291 (N_291,In_515,In_519);
or U292 (N_292,In_639,In_628);
or U293 (N_293,In_403,In_215);
nand U294 (N_294,In_277,In_207);
and U295 (N_295,In_187,In_848);
and U296 (N_296,In_593,In_960);
or U297 (N_297,In_985,In_945);
nor U298 (N_298,In_213,In_657);
nand U299 (N_299,In_464,In_314);
or U300 (N_300,In_510,In_335);
or U301 (N_301,In_342,In_830);
or U302 (N_302,In_351,In_802);
or U303 (N_303,In_940,In_170);
or U304 (N_304,In_186,In_393);
or U305 (N_305,In_20,In_374);
nor U306 (N_306,In_595,In_21);
nor U307 (N_307,In_133,In_894);
or U308 (N_308,In_887,In_60);
and U309 (N_309,In_738,In_609);
nor U310 (N_310,In_157,In_311);
nor U311 (N_311,In_825,In_652);
nand U312 (N_312,In_588,In_663);
or U313 (N_313,In_533,In_710);
nor U314 (N_314,In_986,In_151);
and U315 (N_315,In_529,In_412);
xnor U316 (N_316,In_704,In_820);
or U317 (N_317,In_301,In_906);
nand U318 (N_318,In_772,In_534);
or U319 (N_319,In_429,In_137);
or U320 (N_320,In_192,In_50);
and U321 (N_321,In_953,In_844);
and U322 (N_322,In_482,In_690);
nand U323 (N_323,In_168,In_62);
or U324 (N_324,In_306,In_153);
nor U325 (N_325,In_963,In_806);
or U326 (N_326,In_214,In_95);
or U327 (N_327,In_407,In_831);
nor U328 (N_328,In_411,In_152);
nor U329 (N_329,In_781,In_106);
nand U330 (N_330,In_490,In_39);
nand U331 (N_331,In_541,In_163);
nor U332 (N_332,In_967,In_548);
and U333 (N_333,In_944,In_611);
nand U334 (N_334,In_116,In_70);
nor U335 (N_335,In_653,In_989);
or U336 (N_336,In_642,In_280);
nor U337 (N_337,In_235,In_473);
nor U338 (N_338,In_551,In_716);
and U339 (N_339,In_682,In_82);
or U340 (N_340,In_349,In_824);
and U341 (N_341,In_433,In_385);
nand U342 (N_342,In_711,In_319);
and U343 (N_343,In_847,In_305);
and U344 (N_344,In_872,In_124);
and U345 (N_345,In_424,In_512);
nand U346 (N_346,In_75,In_475);
or U347 (N_347,In_857,In_26);
and U348 (N_348,In_249,In_726);
or U349 (N_349,In_161,In_692);
or U350 (N_350,In_410,In_24);
and U351 (N_351,In_499,In_752);
and U352 (N_352,In_31,In_622);
nand U353 (N_353,In_999,In_600);
or U354 (N_354,In_256,In_145);
and U355 (N_355,In_867,In_638);
and U356 (N_356,In_30,In_472);
nor U357 (N_357,In_880,In_979);
nand U358 (N_358,In_250,In_443);
nand U359 (N_359,In_978,In_449);
nor U360 (N_360,In_117,In_697);
nand U361 (N_361,In_850,In_102);
nor U362 (N_362,In_307,In_291);
nand U363 (N_363,In_948,In_461);
and U364 (N_364,In_554,In_334);
or U365 (N_365,In_811,In_833);
nor U366 (N_366,In_331,In_325);
and U367 (N_367,In_776,In_852);
and U368 (N_368,In_97,In_302);
nand U369 (N_369,In_919,In_399);
nor U370 (N_370,In_346,In_579);
nor U371 (N_371,In_41,In_984);
nand U372 (N_372,In_956,In_328);
nor U373 (N_373,In_916,In_932);
and U374 (N_374,In_577,In_356);
or U375 (N_375,In_206,In_479);
nor U376 (N_376,In_469,In_480);
and U377 (N_377,In_728,In_537);
nand U378 (N_378,In_891,In_64);
nand U379 (N_379,In_815,In_14);
nor U380 (N_380,In_647,In_764);
or U381 (N_381,In_542,In_344);
and U382 (N_382,In_174,In_909);
nand U383 (N_383,In_188,In_951);
and U384 (N_384,In_177,In_105);
or U385 (N_385,In_135,In_863);
nand U386 (N_386,In_396,In_422);
and U387 (N_387,In_624,In_853);
nand U388 (N_388,In_294,In_113);
xnor U389 (N_389,In_162,In_870);
nor U390 (N_390,In_637,In_840);
or U391 (N_391,In_501,In_44);
or U392 (N_392,In_686,In_890);
and U393 (N_393,In_115,In_350);
nor U394 (N_394,In_201,In_659);
or U395 (N_395,In_467,In_939);
nor U396 (N_396,In_601,In_885);
nand U397 (N_397,In_775,In_181);
or U398 (N_398,In_456,In_684);
or U399 (N_399,In_483,In_646);
and U400 (N_400,In_100,In_46);
or U401 (N_401,In_849,In_661);
and U402 (N_402,In_785,In_283);
or U403 (N_403,In_725,In_484);
nand U404 (N_404,In_304,In_655);
and U405 (N_405,In_523,In_983);
nor U406 (N_406,In_623,In_260);
nor U407 (N_407,In_155,In_57);
nor U408 (N_408,In_310,In_735);
nor U409 (N_409,In_681,In_391);
or U410 (N_410,In_943,In_524);
or U411 (N_411,In_315,In_67);
nor U412 (N_412,In_576,In_285);
and U413 (N_413,In_171,In_708);
nand U414 (N_414,In_540,In_907);
nand U415 (N_415,In_817,In_925);
or U416 (N_416,In_614,In_392);
nor U417 (N_417,In_55,In_578);
nor U418 (N_418,In_431,In_378);
and U419 (N_419,In_799,In_241);
and U420 (N_420,In_504,In_992);
and U421 (N_421,In_707,In_835);
and U422 (N_422,In_239,In_564);
nand U423 (N_423,In_901,In_734);
nand U424 (N_424,In_516,In_488);
or U425 (N_425,In_178,In_911);
and U426 (N_426,In_231,In_949);
nor U427 (N_427,In_180,In_715);
and U428 (N_428,In_741,In_873);
nor U429 (N_429,In_228,In_355);
nand U430 (N_430,In_587,In_11);
or U431 (N_431,In_660,In_521);
nand U432 (N_432,In_733,In_753);
nor U433 (N_433,In_376,In_380);
and U434 (N_434,In_664,In_644);
nand U435 (N_435,In_318,In_976);
or U436 (N_436,In_605,In_506);
or U437 (N_437,In_591,In_365);
nand U438 (N_438,In_269,In_316);
nor U439 (N_439,In_107,In_114);
nor U440 (N_440,In_626,In_179);
and U441 (N_441,In_35,In_845);
and U442 (N_442,In_353,In_297);
nand U443 (N_443,In_279,In_545);
or U444 (N_444,In_536,In_618);
and U445 (N_445,In_381,In_29);
or U446 (N_446,In_139,In_650);
nor U447 (N_447,In_696,In_255);
nor U448 (N_448,In_408,In_713);
xnor U449 (N_449,In_780,In_669);
and U450 (N_450,In_539,In_594);
nor U451 (N_451,In_794,In_4);
nor U452 (N_452,In_65,In_560);
nor U453 (N_453,In_119,In_22);
or U454 (N_454,In_18,In_691);
nor U455 (N_455,In_826,In_724);
nand U456 (N_456,In_801,In_266);
nor U457 (N_457,In_580,In_77);
nand U458 (N_458,In_352,In_702);
nand U459 (N_459,In_299,In_338);
nor U460 (N_460,In_730,In_184);
nand U461 (N_461,In_705,In_159);
nor U462 (N_462,In_253,In_173);
or U463 (N_463,In_287,In_58);
or U464 (N_464,In_672,In_476);
or U465 (N_465,In_120,In_604);
and U466 (N_466,In_498,In_240);
nand U467 (N_467,In_278,In_364);
and U468 (N_468,In_970,In_428);
or U469 (N_469,In_674,In_12);
and U470 (N_470,In_868,In_597);
nor U471 (N_471,In_769,In_1);
nand U472 (N_472,In_204,In_779);
nand U473 (N_473,In_468,In_384);
and U474 (N_474,In_402,In_933);
xnor U475 (N_475,In_641,In_821);
or U476 (N_476,In_49,In_627);
nor U477 (N_477,In_903,In_96);
or U478 (N_478,In_47,In_928);
nand U479 (N_479,In_486,In_977);
and U480 (N_480,In_10,In_592);
nor U481 (N_481,In_394,In_871);
and U482 (N_482,In_998,In_842);
or U483 (N_483,In_773,In_13);
nor U484 (N_484,In_606,In_59);
or U485 (N_485,In_574,In_613);
or U486 (N_486,In_988,In_522);
nand U487 (N_487,In_246,In_271);
nand U488 (N_488,In_851,In_48);
nand U489 (N_489,In_421,In_224);
nand U490 (N_490,In_930,In_961);
or U491 (N_491,In_503,In_689);
nor U492 (N_492,In_902,In_795);
nand U493 (N_493,In_221,In_640);
nand U494 (N_494,In_234,In_273);
or U495 (N_495,In_69,In_108);
nor U496 (N_496,In_445,In_731);
and U497 (N_497,In_268,In_210);
or U498 (N_498,In_813,In_150);
and U499 (N_499,In_751,In_56);
or U500 (N_500,In_945,In_117);
or U501 (N_501,In_690,In_568);
nand U502 (N_502,In_650,In_923);
and U503 (N_503,In_735,In_856);
nand U504 (N_504,In_73,In_598);
or U505 (N_505,In_337,In_433);
nand U506 (N_506,In_739,In_145);
nor U507 (N_507,In_620,In_650);
nand U508 (N_508,In_441,In_899);
nand U509 (N_509,In_884,In_86);
and U510 (N_510,In_931,In_308);
nand U511 (N_511,In_40,In_22);
nor U512 (N_512,In_980,In_3);
and U513 (N_513,In_874,In_365);
and U514 (N_514,In_231,In_620);
and U515 (N_515,In_835,In_439);
or U516 (N_516,In_481,In_899);
and U517 (N_517,In_948,In_825);
or U518 (N_518,In_544,In_288);
nand U519 (N_519,In_754,In_386);
and U520 (N_520,In_432,In_31);
and U521 (N_521,In_267,In_271);
nor U522 (N_522,In_17,In_405);
nor U523 (N_523,In_180,In_776);
or U524 (N_524,In_89,In_47);
nor U525 (N_525,In_654,In_533);
nor U526 (N_526,In_718,In_862);
nor U527 (N_527,In_192,In_736);
and U528 (N_528,In_761,In_534);
and U529 (N_529,In_716,In_283);
nand U530 (N_530,In_74,In_284);
and U531 (N_531,In_762,In_213);
xor U532 (N_532,In_623,In_784);
nand U533 (N_533,In_508,In_319);
nor U534 (N_534,In_399,In_808);
nor U535 (N_535,In_637,In_324);
nand U536 (N_536,In_202,In_669);
nand U537 (N_537,In_240,In_316);
and U538 (N_538,In_387,In_708);
xor U539 (N_539,In_749,In_821);
or U540 (N_540,In_360,In_451);
and U541 (N_541,In_756,In_614);
or U542 (N_542,In_568,In_913);
and U543 (N_543,In_622,In_474);
nand U544 (N_544,In_505,In_403);
and U545 (N_545,In_483,In_615);
and U546 (N_546,In_568,In_987);
and U547 (N_547,In_410,In_351);
nor U548 (N_548,In_804,In_109);
or U549 (N_549,In_647,In_238);
and U550 (N_550,In_579,In_928);
nor U551 (N_551,In_137,In_29);
nor U552 (N_552,In_63,In_923);
nor U553 (N_553,In_242,In_478);
nor U554 (N_554,In_244,In_836);
nor U555 (N_555,In_123,In_613);
or U556 (N_556,In_22,In_644);
and U557 (N_557,In_780,In_269);
nor U558 (N_558,In_582,In_744);
nand U559 (N_559,In_82,In_222);
or U560 (N_560,In_414,In_848);
or U561 (N_561,In_780,In_28);
or U562 (N_562,In_435,In_528);
nor U563 (N_563,In_896,In_703);
or U564 (N_564,In_292,In_10);
and U565 (N_565,In_752,In_107);
nand U566 (N_566,In_197,In_105);
nor U567 (N_567,In_883,In_370);
or U568 (N_568,In_724,In_629);
and U569 (N_569,In_909,In_387);
nand U570 (N_570,In_600,In_284);
and U571 (N_571,In_115,In_423);
and U572 (N_572,In_837,In_842);
nor U573 (N_573,In_557,In_826);
nand U574 (N_574,In_218,In_477);
or U575 (N_575,In_792,In_713);
or U576 (N_576,In_724,In_2);
nand U577 (N_577,In_818,In_404);
or U578 (N_578,In_726,In_222);
nor U579 (N_579,In_185,In_346);
or U580 (N_580,In_772,In_73);
or U581 (N_581,In_488,In_81);
or U582 (N_582,In_804,In_955);
and U583 (N_583,In_818,In_3);
nor U584 (N_584,In_319,In_542);
or U585 (N_585,In_859,In_517);
nand U586 (N_586,In_422,In_987);
or U587 (N_587,In_256,In_925);
nor U588 (N_588,In_173,In_499);
and U589 (N_589,In_982,In_948);
nor U590 (N_590,In_12,In_934);
nand U591 (N_591,In_698,In_81);
or U592 (N_592,In_688,In_339);
xor U593 (N_593,In_32,In_715);
nand U594 (N_594,In_920,In_896);
nor U595 (N_595,In_351,In_344);
nand U596 (N_596,In_771,In_629);
nand U597 (N_597,In_336,In_707);
or U598 (N_598,In_378,In_123);
nor U599 (N_599,In_956,In_605);
nor U600 (N_600,In_883,In_343);
nor U601 (N_601,In_651,In_46);
nand U602 (N_602,In_398,In_373);
nor U603 (N_603,In_726,In_255);
or U604 (N_604,In_660,In_753);
nand U605 (N_605,In_556,In_626);
nor U606 (N_606,In_525,In_399);
nor U607 (N_607,In_419,In_92);
nor U608 (N_608,In_388,In_968);
nor U609 (N_609,In_180,In_135);
or U610 (N_610,In_424,In_202);
nor U611 (N_611,In_734,In_381);
nor U612 (N_612,In_16,In_543);
and U613 (N_613,In_699,In_33);
and U614 (N_614,In_946,In_606);
or U615 (N_615,In_995,In_61);
or U616 (N_616,In_735,In_753);
and U617 (N_617,In_353,In_179);
nor U618 (N_618,In_639,In_942);
or U619 (N_619,In_222,In_307);
nor U620 (N_620,In_300,In_28);
nor U621 (N_621,In_596,In_280);
nand U622 (N_622,In_427,In_239);
nor U623 (N_623,In_139,In_590);
nand U624 (N_624,In_260,In_206);
nand U625 (N_625,In_206,In_273);
and U626 (N_626,In_891,In_588);
or U627 (N_627,In_91,In_397);
xor U628 (N_628,In_476,In_164);
nor U629 (N_629,In_224,In_645);
or U630 (N_630,In_262,In_620);
or U631 (N_631,In_794,In_863);
nand U632 (N_632,In_741,In_316);
nand U633 (N_633,In_200,In_534);
or U634 (N_634,In_588,In_413);
nor U635 (N_635,In_347,In_639);
and U636 (N_636,In_595,In_824);
and U637 (N_637,In_271,In_519);
nand U638 (N_638,In_289,In_589);
nand U639 (N_639,In_232,In_585);
nand U640 (N_640,In_77,In_747);
or U641 (N_641,In_9,In_441);
and U642 (N_642,In_624,In_488);
nand U643 (N_643,In_7,In_512);
nor U644 (N_644,In_134,In_671);
or U645 (N_645,In_665,In_853);
nand U646 (N_646,In_582,In_306);
and U647 (N_647,In_24,In_290);
or U648 (N_648,In_241,In_332);
and U649 (N_649,In_66,In_142);
and U650 (N_650,In_180,In_577);
nand U651 (N_651,In_850,In_649);
nand U652 (N_652,In_559,In_983);
or U653 (N_653,In_210,In_890);
or U654 (N_654,In_154,In_576);
or U655 (N_655,In_244,In_17);
nor U656 (N_656,In_5,In_598);
or U657 (N_657,In_936,In_572);
nand U658 (N_658,In_53,In_216);
or U659 (N_659,In_97,In_796);
nor U660 (N_660,In_122,In_906);
and U661 (N_661,In_567,In_484);
nand U662 (N_662,In_988,In_525);
or U663 (N_663,In_618,In_75);
nor U664 (N_664,In_726,In_414);
nor U665 (N_665,In_24,In_892);
nor U666 (N_666,In_149,In_764);
nand U667 (N_667,In_315,In_666);
nor U668 (N_668,In_151,In_94);
nand U669 (N_669,In_611,In_21);
nor U670 (N_670,In_624,In_258);
or U671 (N_671,In_52,In_798);
nor U672 (N_672,In_791,In_738);
or U673 (N_673,In_875,In_757);
or U674 (N_674,In_953,In_268);
nor U675 (N_675,In_63,In_661);
nand U676 (N_676,In_547,In_395);
nor U677 (N_677,In_593,In_659);
xor U678 (N_678,In_1,In_900);
and U679 (N_679,In_141,In_388);
nor U680 (N_680,In_682,In_650);
nand U681 (N_681,In_848,In_562);
xnor U682 (N_682,In_423,In_222);
nand U683 (N_683,In_45,In_365);
and U684 (N_684,In_34,In_600);
and U685 (N_685,In_118,In_220);
and U686 (N_686,In_226,In_889);
or U687 (N_687,In_734,In_104);
nor U688 (N_688,In_472,In_675);
and U689 (N_689,In_592,In_696);
or U690 (N_690,In_474,In_616);
nand U691 (N_691,In_782,In_621);
nor U692 (N_692,In_207,In_790);
nand U693 (N_693,In_845,In_122);
nor U694 (N_694,In_625,In_139);
nor U695 (N_695,In_410,In_632);
or U696 (N_696,In_960,In_432);
and U697 (N_697,In_957,In_688);
and U698 (N_698,In_374,In_300);
or U699 (N_699,In_711,In_446);
or U700 (N_700,In_630,In_85);
and U701 (N_701,In_153,In_402);
nand U702 (N_702,In_253,In_625);
xnor U703 (N_703,In_262,In_165);
nand U704 (N_704,In_459,In_646);
nand U705 (N_705,In_64,In_808);
nor U706 (N_706,In_283,In_870);
or U707 (N_707,In_989,In_632);
and U708 (N_708,In_79,In_455);
and U709 (N_709,In_279,In_58);
and U710 (N_710,In_520,In_614);
nor U711 (N_711,In_572,In_563);
nor U712 (N_712,In_481,In_625);
nor U713 (N_713,In_13,In_948);
nor U714 (N_714,In_169,In_672);
xnor U715 (N_715,In_189,In_51);
or U716 (N_716,In_101,In_137);
nand U717 (N_717,In_49,In_373);
nand U718 (N_718,In_132,In_47);
nand U719 (N_719,In_363,In_777);
or U720 (N_720,In_668,In_570);
nor U721 (N_721,In_787,In_620);
nand U722 (N_722,In_816,In_196);
nand U723 (N_723,In_133,In_41);
and U724 (N_724,In_2,In_198);
nor U725 (N_725,In_594,In_935);
or U726 (N_726,In_377,In_442);
and U727 (N_727,In_862,In_952);
nand U728 (N_728,In_172,In_993);
xor U729 (N_729,In_8,In_824);
or U730 (N_730,In_24,In_336);
or U731 (N_731,In_266,In_292);
nand U732 (N_732,In_326,In_411);
nand U733 (N_733,In_467,In_739);
and U734 (N_734,In_198,In_759);
nor U735 (N_735,In_374,In_814);
and U736 (N_736,In_821,In_257);
or U737 (N_737,In_413,In_535);
nor U738 (N_738,In_57,In_525);
or U739 (N_739,In_955,In_228);
nand U740 (N_740,In_870,In_982);
or U741 (N_741,In_6,In_405);
nand U742 (N_742,In_551,In_152);
nor U743 (N_743,In_986,In_949);
nor U744 (N_744,In_353,In_495);
and U745 (N_745,In_880,In_171);
xor U746 (N_746,In_723,In_361);
and U747 (N_747,In_61,In_103);
nor U748 (N_748,In_100,In_589);
nor U749 (N_749,In_36,In_540);
nor U750 (N_750,In_567,In_776);
and U751 (N_751,In_679,In_731);
and U752 (N_752,In_998,In_580);
and U753 (N_753,In_526,In_239);
nor U754 (N_754,In_777,In_72);
or U755 (N_755,In_638,In_12);
nand U756 (N_756,In_653,In_368);
nand U757 (N_757,In_743,In_795);
nor U758 (N_758,In_762,In_710);
or U759 (N_759,In_364,In_299);
nand U760 (N_760,In_852,In_981);
and U761 (N_761,In_993,In_410);
or U762 (N_762,In_841,In_314);
nand U763 (N_763,In_823,In_638);
or U764 (N_764,In_373,In_163);
or U765 (N_765,In_750,In_469);
and U766 (N_766,In_880,In_992);
nor U767 (N_767,In_468,In_290);
nand U768 (N_768,In_652,In_576);
and U769 (N_769,In_784,In_248);
nand U770 (N_770,In_413,In_985);
nand U771 (N_771,In_660,In_786);
nor U772 (N_772,In_694,In_588);
nor U773 (N_773,In_535,In_730);
nor U774 (N_774,In_295,In_536);
or U775 (N_775,In_444,In_198);
and U776 (N_776,In_744,In_759);
or U777 (N_777,In_963,In_22);
or U778 (N_778,In_900,In_289);
or U779 (N_779,In_386,In_496);
nor U780 (N_780,In_509,In_392);
and U781 (N_781,In_444,In_626);
nor U782 (N_782,In_945,In_793);
nand U783 (N_783,In_29,In_719);
nor U784 (N_784,In_269,In_281);
and U785 (N_785,In_78,In_784);
and U786 (N_786,In_188,In_56);
and U787 (N_787,In_920,In_500);
and U788 (N_788,In_327,In_161);
and U789 (N_789,In_188,In_293);
nand U790 (N_790,In_411,In_288);
and U791 (N_791,In_150,In_28);
and U792 (N_792,In_89,In_883);
nor U793 (N_793,In_373,In_934);
xor U794 (N_794,In_555,In_896);
or U795 (N_795,In_238,In_614);
nor U796 (N_796,In_930,In_327);
nor U797 (N_797,In_421,In_155);
xnor U798 (N_798,In_462,In_420);
nand U799 (N_799,In_219,In_854);
nor U800 (N_800,In_357,In_56);
or U801 (N_801,In_783,In_984);
nand U802 (N_802,In_735,In_87);
or U803 (N_803,In_378,In_249);
or U804 (N_804,In_955,In_741);
or U805 (N_805,In_278,In_799);
nor U806 (N_806,In_230,In_757);
nand U807 (N_807,In_548,In_527);
and U808 (N_808,In_966,In_442);
or U809 (N_809,In_534,In_602);
and U810 (N_810,In_54,In_539);
or U811 (N_811,In_273,In_146);
and U812 (N_812,In_682,In_74);
and U813 (N_813,In_383,In_655);
nor U814 (N_814,In_622,In_517);
or U815 (N_815,In_650,In_242);
nor U816 (N_816,In_272,In_825);
and U817 (N_817,In_997,In_793);
nand U818 (N_818,In_13,In_642);
and U819 (N_819,In_221,In_268);
and U820 (N_820,In_267,In_317);
and U821 (N_821,In_162,In_993);
nor U822 (N_822,In_95,In_453);
nor U823 (N_823,In_154,In_309);
nor U824 (N_824,In_574,In_2);
nor U825 (N_825,In_110,In_988);
and U826 (N_826,In_897,In_744);
nor U827 (N_827,In_185,In_887);
nor U828 (N_828,In_90,In_301);
nor U829 (N_829,In_719,In_610);
or U830 (N_830,In_180,In_424);
or U831 (N_831,In_846,In_448);
nand U832 (N_832,In_606,In_936);
nor U833 (N_833,In_190,In_567);
and U834 (N_834,In_194,In_513);
nand U835 (N_835,In_67,In_620);
nor U836 (N_836,In_560,In_340);
or U837 (N_837,In_611,In_401);
or U838 (N_838,In_647,In_925);
nand U839 (N_839,In_295,In_959);
and U840 (N_840,In_17,In_367);
and U841 (N_841,In_286,In_896);
nand U842 (N_842,In_888,In_965);
nor U843 (N_843,In_649,In_325);
or U844 (N_844,In_483,In_515);
nor U845 (N_845,In_424,In_375);
and U846 (N_846,In_998,In_892);
nor U847 (N_847,In_502,In_65);
or U848 (N_848,In_887,In_528);
nand U849 (N_849,In_290,In_0);
xnor U850 (N_850,In_233,In_188);
and U851 (N_851,In_613,In_771);
nand U852 (N_852,In_684,In_311);
or U853 (N_853,In_667,In_999);
and U854 (N_854,In_15,In_734);
nor U855 (N_855,In_522,In_136);
nor U856 (N_856,In_663,In_724);
or U857 (N_857,In_762,In_857);
nor U858 (N_858,In_449,In_997);
nand U859 (N_859,In_740,In_349);
nand U860 (N_860,In_986,In_295);
nand U861 (N_861,In_627,In_617);
nand U862 (N_862,In_534,In_929);
nor U863 (N_863,In_961,In_391);
and U864 (N_864,In_859,In_525);
nor U865 (N_865,In_241,In_474);
and U866 (N_866,In_935,In_511);
and U867 (N_867,In_326,In_435);
or U868 (N_868,In_354,In_105);
or U869 (N_869,In_168,In_763);
and U870 (N_870,In_980,In_109);
and U871 (N_871,In_536,In_97);
nand U872 (N_872,In_776,In_349);
or U873 (N_873,In_906,In_20);
and U874 (N_874,In_553,In_602);
nor U875 (N_875,In_526,In_582);
or U876 (N_876,In_684,In_860);
xor U877 (N_877,In_75,In_882);
and U878 (N_878,In_197,In_747);
or U879 (N_879,In_408,In_521);
or U880 (N_880,In_575,In_453);
nor U881 (N_881,In_317,In_595);
or U882 (N_882,In_2,In_346);
nor U883 (N_883,In_283,In_78);
xor U884 (N_884,In_476,In_94);
nand U885 (N_885,In_968,In_696);
nor U886 (N_886,In_317,In_955);
or U887 (N_887,In_28,In_433);
or U888 (N_888,In_23,In_9);
nand U889 (N_889,In_336,In_972);
or U890 (N_890,In_843,In_367);
nand U891 (N_891,In_706,In_870);
or U892 (N_892,In_404,In_548);
nand U893 (N_893,In_9,In_624);
and U894 (N_894,In_849,In_955);
and U895 (N_895,In_893,In_523);
nand U896 (N_896,In_505,In_587);
and U897 (N_897,In_579,In_322);
nor U898 (N_898,In_16,In_499);
and U899 (N_899,In_41,In_291);
nor U900 (N_900,In_532,In_901);
or U901 (N_901,In_154,In_47);
nor U902 (N_902,In_618,In_237);
and U903 (N_903,In_933,In_515);
nor U904 (N_904,In_716,In_676);
nand U905 (N_905,In_421,In_321);
and U906 (N_906,In_613,In_558);
nand U907 (N_907,In_569,In_25);
or U908 (N_908,In_56,In_782);
xor U909 (N_909,In_131,In_105);
nand U910 (N_910,In_463,In_436);
and U911 (N_911,In_70,In_295);
nor U912 (N_912,In_469,In_560);
and U913 (N_913,In_578,In_255);
nor U914 (N_914,In_103,In_362);
nor U915 (N_915,In_318,In_346);
nor U916 (N_916,In_543,In_658);
nor U917 (N_917,In_126,In_722);
or U918 (N_918,In_341,In_520);
nand U919 (N_919,In_836,In_39);
and U920 (N_920,In_526,In_481);
and U921 (N_921,In_106,In_815);
or U922 (N_922,In_98,In_156);
nand U923 (N_923,In_385,In_913);
nor U924 (N_924,In_449,In_520);
nor U925 (N_925,In_325,In_25);
or U926 (N_926,In_257,In_761);
nor U927 (N_927,In_984,In_544);
xor U928 (N_928,In_247,In_383);
nand U929 (N_929,In_654,In_777);
nand U930 (N_930,In_450,In_895);
nor U931 (N_931,In_512,In_445);
nor U932 (N_932,In_111,In_82);
and U933 (N_933,In_424,In_518);
xnor U934 (N_934,In_984,In_581);
nor U935 (N_935,In_822,In_197);
nand U936 (N_936,In_783,In_879);
nand U937 (N_937,In_43,In_312);
nand U938 (N_938,In_738,In_342);
nand U939 (N_939,In_193,In_447);
and U940 (N_940,In_756,In_708);
nand U941 (N_941,In_536,In_987);
or U942 (N_942,In_409,In_580);
and U943 (N_943,In_582,In_603);
and U944 (N_944,In_959,In_581);
and U945 (N_945,In_291,In_910);
and U946 (N_946,In_504,In_114);
and U947 (N_947,In_260,In_765);
or U948 (N_948,In_689,In_322);
xnor U949 (N_949,In_700,In_723);
or U950 (N_950,In_205,In_819);
nor U951 (N_951,In_554,In_238);
nand U952 (N_952,In_398,In_500);
and U953 (N_953,In_281,In_698);
and U954 (N_954,In_0,In_895);
nand U955 (N_955,In_754,In_773);
or U956 (N_956,In_809,In_13);
nor U957 (N_957,In_507,In_498);
nor U958 (N_958,In_314,In_836);
or U959 (N_959,In_96,In_80);
and U960 (N_960,In_821,In_908);
and U961 (N_961,In_568,In_85);
and U962 (N_962,In_81,In_604);
and U963 (N_963,In_64,In_10);
or U964 (N_964,In_188,In_326);
nand U965 (N_965,In_460,In_22);
nand U966 (N_966,In_117,In_387);
or U967 (N_967,In_603,In_790);
or U968 (N_968,In_801,In_122);
nand U969 (N_969,In_822,In_592);
nand U970 (N_970,In_875,In_716);
nand U971 (N_971,In_578,In_64);
or U972 (N_972,In_513,In_573);
nand U973 (N_973,In_884,In_961);
xor U974 (N_974,In_900,In_417);
nor U975 (N_975,In_428,In_631);
nor U976 (N_976,In_832,In_732);
or U977 (N_977,In_412,In_532);
nor U978 (N_978,In_888,In_524);
nor U979 (N_979,In_246,In_125);
and U980 (N_980,In_242,In_558);
and U981 (N_981,In_442,In_753);
nor U982 (N_982,In_673,In_499);
and U983 (N_983,In_332,In_148);
and U984 (N_984,In_323,In_176);
and U985 (N_985,In_24,In_924);
or U986 (N_986,In_468,In_723);
or U987 (N_987,In_835,In_280);
and U988 (N_988,In_814,In_633);
and U989 (N_989,In_693,In_812);
nand U990 (N_990,In_473,In_18);
nand U991 (N_991,In_78,In_764);
or U992 (N_992,In_482,In_218);
and U993 (N_993,In_699,In_85);
and U994 (N_994,In_396,In_254);
xnor U995 (N_995,In_721,In_328);
or U996 (N_996,In_802,In_519);
nand U997 (N_997,In_683,In_670);
or U998 (N_998,In_469,In_29);
nor U999 (N_999,In_726,In_253);
or U1000 (N_1000,In_347,In_49);
nand U1001 (N_1001,In_394,In_757);
nor U1002 (N_1002,In_670,In_171);
nor U1003 (N_1003,In_105,In_723);
or U1004 (N_1004,In_479,In_223);
nand U1005 (N_1005,In_585,In_511);
or U1006 (N_1006,In_603,In_919);
nor U1007 (N_1007,In_951,In_16);
xor U1008 (N_1008,In_872,In_264);
nand U1009 (N_1009,In_963,In_481);
nor U1010 (N_1010,In_622,In_349);
nand U1011 (N_1011,In_194,In_790);
nand U1012 (N_1012,In_22,In_994);
or U1013 (N_1013,In_942,In_850);
nand U1014 (N_1014,In_154,In_731);
nand U1015 (N_1015,In_429,In_483);
nor U1016 (N_1016,In_237,In_555);
nand U1017 (N_1017,In_425,In_958);
or U1018 (N_1018,In_867,In_841);
and U1019 (N_1019,In_909,In_210);
nand U1020 (N_1020,In_253,In_773);
nor U1021 (N_1021,In_518,In_15);
nor U1022 (N_1022,In_671,In_414);
nor U1023 (N_1023,In_727,In_369);
nor U1024 (N_1024,In_427,In_774);
nor U1025 (N_1025,In_944,In_440);
nor U1026 (N_1026,In_301,In_883);
nand U1027 (N_1027,In_158,In_371);
and U1028 (N_1028,In_729,In_595);
and U1029 (N_1029,In_593,In_231);
or U1030 (N_1030,In_172,In_461);
nor U1031 (N_1031,In_909,In_960);
nor U1032 (N_1032,In_590,In_759);
nand U1033 (N_1033,In_851,In_279);
nand U1034 (N_1034,In_373,In_795);
nand U1035 (N_1035,In_1,In_206);
or U1036 (N_1036,In_518,In_723);
nand U1037 (N_1037,In_820,In_611);
nor U1038 (N_1038,In_296,In_280);
nand U1039 (N_1039,In_816,In_671);
xor U1040 (N_1040,In_375,In_463);
and U1041 (N_1041,In_337,In_845);
nand U1042 (N_1042,In_653,In_415);
and U1043 (N_1043,In_214,In_796);
or U1044 (N_1044,In_600,In_90);
nor U1045 (N_1045,In_358,In_749);
nand U1046 (N_1046,In_913,In_689);
and U1047 (N_1047,In_999,In_882);
and U1048 (N_1048,In_105,In_890);
or U1049 (N_1049,In_220,In_147);
or U1050 (N_1050,In_292,In_367);
nand U1051 (N_1051,In_910,In_804);
nand U1052 (N_1052,In_609,In_302);
or U1053 (N_1053,In_360,In_291);
or U1054 (N_1054,In_659,In_523);
and U1055 (N_1055,In_229,In_817);
nor U1056 (N_1056,In_602,In_418);
nor U1057 (N_1057,In_94,In_928);
or U1058 (N_1058,In_200,In_508);
nor U1059 (N_1059,In_45,In_991);
or U1060 (N_1060,In_945,In_699);
or U1061 (N_1061,In_450,In_154);
nor U1062 (N_1062,In_923,In_528);
and U1063 (N_1063,In_827,In_221);
nor U1064 (N_1064,In_390,In_617);
or U1065 (N_1065,In_577,In_860);
nand U1066 (N_1066,In_42,In_694);
nand U1067 (N_1067,In_506,In_958);
nor U1068 (N_1068,In_362,In_913);
and U1069 (N_1069,In_243,In_651);
and U1070 (N_1070,In_355,In_152);
nor U1071 (N_1071,In_120,In_32);
nor U1072 (N_1072,In_553,In_975);
nand U1073 (N_1073,In_580,In_397);
xor U1074 (N_1074,In_620,In_60);
or U1075 (N_1075,In_77,In_690);
nor U1076 (N_1076,In_169,In_978);
nand U1077 (N_1077,In_371,In_519);
or U1078 (N_1078,In_483,In_994);
nand U1079 (N_1079,In_506,In_144);
or U1080 (N_1080,In_777,In_47);
xnor U1081 (N_1081,In_842,In_622);
nand U1082 (N_1082,In_469,In_134);
nor U1083 (N_1083,In_919,In_677);
and U1084 (N_1084,In_732,In_987);
and U1085 (N_1085,In_820,In_144);
nor U1086 (N_1086,In_712,In_579);
nor U1087 (N_1087,In_256,In_323);
nor U1088 (N_1088,In_443,In_746);
nand U1089 (N_1089,In_933,In_755);
nand U1090 (N_1090,In_942,In_949);
nand U1091 (N_1091,In_318,In_79);
nand U1092 (N_1092,In_767,In_861);
and U1093 (N_1093,In_596,In_895);
or U1094 (N_1094,In_12,In_327);
nor U1095 (N_1095,In_164,In_14);
or U1096 (N_1096,In_705,In_507);
or U1097 (N_1097,In_770,In_71);
nor U1098 (N_1098,In_341,In_716);
and U1099 (N_1099,In_575,In_680);
or U1100 (N_1100,In_337,In_419);
or U1101 (N_1101,In_482,In_222);
nand U1102 (N_1102,In_285,In_618);
or U1103 (N_1103,In_807,In_780);
nand U1104 (N_1104,In_703,In_435);
nand U1105 (N_1105,In_751,In_511);
or U1106 (N_1106,In_152,In_443);
and U1107 (N_1107,In_438,In_625);
nand U1108 (N_1108,In_586,In_801);
nand U1109 (N_1109,In_6,In_335);
and U1110 (N_1110,In_714,In_430);
nand U1111 (N_1111,In_361,In_473);
and U1112 (N_1112,In_605,In_490);
nor U1113 (N_1113,In_108,In_699);
and U1114 (N_1114,In_151,In_193);
nor U1115 (N_1115,In_13,In_703);
nand U1116 (N_1116,In_399,In_653);
and U1117 (N_1117,In_932,In_74);
xnor U1118 (N_1118,In_18,In_309);
nand U1119 (N_1119,In_44,In_38);
or U1120 (N_1120,In_438,In_415);
and U1121 (N_1121,In_331,In_989);
nand U1122 (N_1122,In_645,In_995);
nand U1123 (N_1123,In_968,In_365);
or U1124 (N_1124,In_128,In_390);
and U1125 (N_1125,In_657,In_740);
and U1126 (N_1126,In_193,In_139);
and U1127 (N_1127,In_733,In_372);
or U1128 (N_1128,In_348,In_24);
nand U1129 (N_1129,In_15,In_402);
nor U1130 (N_1130,In_12,In_76);
nor U1131 (N_1131,In_145,In_133);
xnor U1132 (N_1132,In_374,In_774);
or U1133 (N_1133,In_309,In_588);
nand U1134 (N_1134,In_936,In_742);
nor U1135 (N_1135,In_674,In_444);
or U1136 (N_1136,In_23,In_871);
nand U1137 (N_1137,In_688,In_106);
nand U1138 (N_1138,In_194,In_298);
nand U1139 (N_1139,In_483,In_816);
xor U1140 (N_1140,In_854,In_610);
or U1141 (N_1141,In_132,In_120);
nor U1142 (N_1142,In_578,In_494);
or U1143 (N_1143,In_729,In_31);
nand U1144 (N_1144,In_996,In_175);
or U1145 (N_1145,In_994,In_175);
or U1146 (N_1146,In_904,In_425);
nor U1147 (N_1147,In_644,In_901);
nand U1148 (N_1148,In_532,In_586);
and U1149 (N_1149,In_550,In_205);
or U1150 (N_1150,In_488,In_528);
and U1151 (N_1151,In_223,In_378);
nand U1152 (N_1152,In_928,In_580);
nand U1153 (N_1153,In_447,In_537);
and U1154 (N_1154,In_690,In_650);
nand U1155 (N_1155,In_367,In_854);
or U1156 (N_1156,In_943,In_692);
nand U1157 (N_1157,In_473,In_769);
or U1158 (N_1158,In_555,In_995);
and U1159 (N_1159,In_856,In_575);
xor U1160 (N_1160,In_216,In_710);
nor U1161 (N_1161,In_724,In_410);
nor U1162 (N_1162,In_988,In_47);
and U1163 (N_1163,In_751,In_480);
nor U1164 (N_1164,In_380,In_350);
nor U1165 (N_1165,In_726,In_33);
and U1166 (N_1166,In_55,In_321);
nand U1167 (N_1167,In_620,In_838);
and U1168 (N_1168,In_754,In_964);
nand U1169 (N_1169,In_476,In_358);
and U1170 (N_1170,In_991,In_540);
or U1171 (N_1171,In_93,In_958);
and U1172 (N_1172,In_435,In_494);
nor U1173 (N_1173,In_904,In_508);
and U1174 (N_1174,In_735,In_129);
or U1175 (N_1175,In_951,In_496);
and U1176 (N_1176,In_980,In_750);
nor U1177 (N_1177,In_534,In_746);
and U1178 (N_1178,In_190,In_328);
nand U1179 (N_1179,In_439,In_261);
nor U1180 (N_1180,In_163,In_111);
nand U1181 (N_1181,In_709,In_265);
nor U1182 (N_1182,In_910,In_868);
xor U1183 (N_1183,In_184,In_860);
or U1184 (N_1184,In_409,In_54);
nor U1185 (N_1185,In_55,In_457);
and U1186 (N_1186,In_739,In_821);
nand U1187 (N_1187,In_332,In_931);
nand U1188 (N_1188,In_84,In_727);
nor U1189 (N_1189,In_399,In_108);
or U1190 (N_1190,In_134,In_903);
and U1191 (N_1191,In_279,In_898);
and U1192 (N_1192,In_897,In_235);
nor U1193 (N_1193,In_115,In_486);
and U1194 (N_1194,In_785,In_727);
nor U1195 (N_1195,In_625,In_65);
or U1196 (N_1196,In_531,In_310);
nor U1197 (N_1197,In_294,In_857);
nor U1198 (N_1198,In_415,In_314);
or U1199 (N_1199,In_463,In_296);
nand U1200 (N_1200,In_719,In_142);
nor U1201 (N_1201,In_624,In_158);
nor U1202 (N_1202,In_39,In_782);
nor U1203 (N_1203,In_272,In_919);
or U1204 (N_1204,In_117,In_28);
nand U1205 (N_1205,In_950,In_592);
or U1206 (N_1206,In_35,In_183);
xnor U1207 (N_1207,In_103,In_596);
and U1208 (N_1208,In_557,In_631);
and U1209 (N_1209,In_842,In_957);
and U1210 (N_1210,In_629,In_755);
nor U1211 (N_1211,In_914,In_976);
nor U1212 (N_1212,In_17,In_151);
nor U1213 (N_1213,In_152,In_786);
and U1214 (N_1214,In_788,In_419);
and U1215 (N_1215,In_953,In_524);
nor U1216 (N_1216,In_292,In_933);
or U1217 (N_1217,In_889,In_996);
nor U1218 (N_1218,In_175,In_218);
nor U1219 (N_1219,In_482,In_264);
or U1220 (N_1220,In_366,In_179);
nand U1221 (N_1221,In_394,In_154);
nor U1222 (N_1222,In_887,In_355);
or U1223 (N_1223,In_930,In_393);
or U1224 (N_1224,In_710,In_953);
nand U1225 (N_1225,In_920,In_308);
or U1226 (N_1226,In_647,In_849);
or U1227 (N_1227,In_378,In_305);
and U1228 (N_1228,In_551,In_966);
nand U1229 (N_1229,In_216,In_440);
and U1230 (N_1230,In_904,In_630);
or U1231 (N_1231,In_381,In_801);
and U1232 (N_1232,In_554,In_831);
and U1233 (N_1233,In_146,In_3);
nor U1234 (N_1234,In_944,In_477);
and U1235 (N_1235,In_611,In_26);
nor U1236 (N_1236,In_357,In_364);
or U1237 (N_1237,In_696,In_921);
nor U1238 (N_1238,In_877,In_598);
nor U1239 (N_1239,In_792,In_982);
and U1240 (N_1240,In_64,In_825);
and U1241 (N_1241,In_700,In_610);
or U1242 (N_1242,In_238,In_86);
nand U1243 (N_1243,In_479,In_990);
and U1244 (N_1244,In_741,In_207);
or U1245 (N_1245,In_876,In_964);
nor U1246 (N_1246,In_491,In_536);
and U1247 (N_1247,In_474,In_925);
and U1248 (N_1248,In_508,In_34);
and U1249 (N_1249,In_423,In_373);
and U1250 (N_1250,In_237,In_594);
and U1251 (N_1251,In_571,In_11);
nand U1252 (N_1252,In_554,In_787);
and U1253 (N_1253,In_967,In_152);
nor U1254 (N_1254,In_104,In_668);
nor U1255 (N_1255,In_349,In_581);
or U1256 (N_1256,In_887,In_132);
and U1257 (N_1257,In_2,In_483);
nand U1258 (N_1258,In_727,In_724);
and U1259 (N_1259,In_200,In_481);
or U1260 (N_1260,In_94,In_530);
or U1261 (N_1261,In_64,In_285);
and U1262 (N_1262,In_943,In_438);
or U1263 (N_1263,In_882,In_435);
or U1264 (N_1264,In_970,In_510);
and U1265 (N_1265,In_928,In_842);
and U1266 (N_1266,In_236,In_536);
and U1267 (N_1267,In_181,In_586);
nand U1268 (N_1268,In_609,In_344);
nand U1269 (N_1269,In_15,In_954);
nor U1270 (N_1270,In_596,In_156);
nand U1271 (N_1271,In_915,In_154);
nor U1272 (N_1272,In_51,In_831);
nor U1273 (N_1273,In_717,In_927);
and U1274 (N_1274,In_808,In_26);
or U1275 (N_1275,In_583,In_392);
xor U1276 (N_1276,In_213,In_586);
nor U1277 (N_1277,In_858,In_6);
or U1278 (N_1278,In_823,In_961);
xor U1279 (N_1279,In_617,In_808);
and U1280 (N_1280,In_735,In_508);
nor U1281 (N_1281,In_266,In_333);
or U1282 (N_1282,In_697,In_873);
nand U1283 (N_1283,In_349,In_565);
nand U1284 (N_1284,In_680,In_110);
nor U1285 (N_1285,In_940,In_142);
and U1286 (N_1286,In_767,In_110);
nand U1287 (N_1287,In_525,In_557);
nor U1288 (N_1288,In_895,In_227);
and U1289 (N_1289,In_64,In_946);
nand U1290 (N_1290,In_508,In_412);
or U1291 (N_1291,In_486,In_72);
or U1292 (N_1292,In_427,In_259);
or U1293 (N_1293,In_563,In_731);
nand U1294 (N_1294,In_266,In_843);
or U1295 (N_1295,In_238,In_399);
nand U1296 (N_1296,In_32,In_443);
and U1297 (N_1297,In_361,In_752);
or U1298 (N_1298,In_889,In_477);
nor U1299 (N_1299,In_565,In_446);
nor U1300 (N_1300,In_491,In_713);
nor U1301 (N_1301,In_438,In_584);
nor U1302 (N_1302,In_593,In_826);
or U1303 (N_1303,In_323,In_745);
and U1304 (N_1304,In_963,In_7);
and U1305 (N_1305,In_627,In_792);
and U1306 (N_1306,In_508,In_72);
or U1307 (N_1307,In_977,In_815);
or U1308 (N_1308,In_788,In_873);
nand U1309 (N_1309,In_79,In_828);
nor U1310 (N_1310,In_218,In_542);
or U1311 (N_1311,In_951,In_770);
xor U1312 (N_1312,In_164,In_12);
or U1313 (N_1313,In_763,In_41);
nand U1314 (N_1314,In_979,In_735);
nor U1315 (N_1315,In_181,In_785);
nor U1316 (N_1316,In_99,In_582);
nand U1317 (N_1317,In_232,In_479);
nand U1318 (N_1318,In_459,In_704);
nand U1319 (N_1319,In_959,In_773);
and U1320 (N_1320,In_580,In_658);
or U1321 (N_1321,In_772,In_403);
nand U1322 (N_1322,In_513,In_36);
nor U1323 (N_1323,In_483,In_929);
nand U1324 (N_1324,In_266,In_102);
and U1325 (N_1325,In_46,In_141);
and U1326 (N_1326,In_758,In_401);
or U1327 (N_1327,In_454,In_968);
and U1328 (N_1328,In_864,In_382);
nand U1329 (N_1329,In_572,In_677);
or U1330 (N_1330,In_235,In_44);
nor U1331 (N_1331,In_733,In_771);
nor U1332 (N_1332,In_603,In_931);
nand U1333 (N_1333,In_166,In_970);
or U1334 (N_1334,In_848,In_459);
nor U1335 (N_1335,In_845,In_82);
nor U1336 (N_1336,In_121,In_748);
or U1337 (N_1337,In_513,In_470);
xor U1338 (N_1338,In_355,In_944);
nand U1339 (N_1339,In_232,In_549);
nand U1340 (N_1340,In_76,In_718);
and U1341 (N_1341,In_738,In_597);
xnor U1342 (N_1342,In_514,In_114);
nand U1343 (N_1343,In_808,In_614);
or U1344 (N_1344,In_973,In_541);
nand U1345 (N_1345,In_438,In_941);
or U1346 (N_1346,In_90,In_120);
nand U1347 (N_1347,In_941,In_901);
nor U1348 (N_1348,In_89,In_539);
nand U1349 (N_1349,In_565,In_383);
or U1350 (N_1350,In_534,In_898);
nor U1351 (N_1351,In_546,In_703);
nor U1352 (N_1352,In_899,In_439);
and U1353 (N_1353,In_839,In_122);
nand U1354 (N_1354,In_192,In_814);
nand U1355 (N_1355,In_388,In_734);
or U1356 (N_1356,In_966,In_776);
nor U1357 (N_1357,In_974,In_561);
nor U1358 (N_1358,In_873,In_758);
or U1359 (N_1359,In_110,In_84);
nand U1360 (N_1360,In_979,In_251);
xnor U1361 (N_1361,In_811,In_354);
nand U1362 (N_1362,In_759,In_945);
and U1363 (N_1363,In_799,In_708);
nand U1364 (N_1364,In_436,In_872);
or U1365 (N_1365,In_710,In_590);
or U1366 (N_1366,In_366,In_874);
nand U1367 (N_1367,In_20,In_34);
nor U1368 (N_1368,In_924,In_674);
or U1369 (N_1369,In_998,In_659);
and U1370 (N_1370,In_545,In_536);
and U1371 (N_1371,In_735,In_636);
nor U1372 (N_1372,In_223,In_221);
or U1373 (N_1373,In_817,In_34);
nor U1374 (N_1374,In_601,In_410);
nand U1375 (N_1375,In_796,In_532);
xnor U1376 (N_1376,In_330,In_345);
nand U1377 (N_1377,In_396,In_210);
or U1378 (N_1378,In_938,In_72);
nand U1379 (N_1379,In_326,In_935);
nand U1380 (N_1380,In_205,In_835);
nand U1381 (N_1381,In_111,In_525);
nand U1382 (N_1382,In_999,In_117);
nand U1383 (N_1383,In_386,In_673);
or U1384 (N_1384,In_265,In_530);
xnor U1385 (N_1385,In_426,In_384);
xnor U1386 (N_1386,In_627,In_464);
nor U1387 (N_1387,In_372,In_110);
nor U1388 (N_1388,In_245,In_647);
or U1389 (N_1389,In_464,In_952);
or U1390 (N_1390,In_946,In_792);
and U1391 (N_1391,In_881,In_567);
and U1392 (N_1392,In_609,In_652);
nand U1393 (N_1393,In_975,In_520);
nand U1394 (N_1394,In_940,In_589);
nor U1395 (N_1395,In_581,In_985);
or U1396 (N_1396,In_100,In_431);
nor U1397 (N_1397,In_94,In_659);
or U1398 (N_1398,In_627,In_586);
nand U1399 (N_1399,In_441,In_573);
nor U1400 (N_1400,In_968,In_484);
or U1401 (N_1401,In_227,In_730);
and U1402 (N_1402,In_122,In_206);
nor U1403 (N_1403,In_81,In_689);
nor U1404 (N_1404,In_98,In_204);
nand U1405 (N_1405,In_216,In_142);
or U1406 (N_1406,In_355,In_494);
and U1407 (N_1407,In_902,In_170);
and U1408 (N_1408,In_664,In_528);
or U1409 (N_1409,In_7,In_850);
nor U1410 (N_1410,In_435,In_740);
and U1411 (N_1411,In_860,In_360);
and U1412 (N_1412,In_762,In_77);
and U1413 (N_1413,In_956,In_886);
nand U1414 (N_1414,In_929,In_56);
and U1415 (N_1415,In_219,In_409);
nand U1416 (N_1416,In_405,In_751);
nand U1417 (N_1417,In_836,In_137);
or U1418 (N_1418,In_7,In_379);
nor U1419 (N_1419,In_585,In_336);
nand U1420 (N_1420,In_770,In_683);
nor U1421 (N_1421,In_297,In_933);
nor U1422 (N_1422,In_777,In_231);
nand U1423 (N_1423,In_337,In_637);
nand U1424 (N_1424,In_847,In_714);
nand U1425 (N_1425,In_932,In_251);
or U1426 (N_1426,In_81,In_185);
and U1427 (N_1427,In_320,In_562);
or U1428 (N_1428,In_56,In_659);
nand U1429 (N_1429,In_603,In_366);
or U1430 (N_1430,In_616,In_222);
and U1431 (N_1431,In_819,In_166);
and U1432 (N_1432,In_961,In_852);
nor U1433 (N_1433,In_924,In_369);
nand U1434 (N_1434,In_123,In_169);
or U1435 (N_1435,In_333,In_853);
or U1436 (N_1436,In_116,In_606);
nand U1437 (N_1437,In_3,In_352);
nor U1438 (N_1438,In_987,In_493);
nor U1439 (N_1439,In_439,In_131);
and U1440 (N_1440,In_754,In_650);
or U1441 (N_1441,In_323,In_843);
or U1442 (N_1442,In_586,In_828);
nand U1443 (N_1443,In_83,In_255);
and U1444 (N_1444,In_343,In_827);
or U1445 (N_1445,In_609,In_527);
nor U1446 (N_1446,In_304,In_414);
or U1447 (N_1447,In_28,In_563);
and U1448 (N_1448,In_956,In_690);
nor U1449 (N_1449,In_318,In_746);
nor U1450 (N_1450,In_209,In_972);
nand U1451 (N_1451,In_404,In_199);
nor U1452 (N_1452,In_554,In_22);
nand U1453 (N_1453,In_990,In_575);
nor U1454 (N_1454,In_930,In_771);
and U1455 (N_1455,In_15,In_48);
xor U1456 (N_1456,In_821,In_272);
or U1457 (N_1457,In_13,In_300);
and U1458 (N_1458,In_624,In_966);
and U1459 (N_1459,In_564,In_668);
or U1460 (N_1460,In_935,In_51);
or U1461 (N_1461,In_392,In_185);
nor U1462 (N_1462,In_141,In_877);
nor U1463 (N_1463,In_389,In_328);
and U1464 (N_1464,In_905,In_570);
nand U1465 (N_1465,In_102,In_246);
or U1466 (N_1466,In_111,In_57);
nand U1467 (N_1467,In_317,In_727);
or U1468 (N_1468,In_723,In_629);
xor U1469 (N_1469,In_786,In_144);
nand U1470 (N_1470,In_302,In_240);
nand U1471 (N_1471,In_345,In_349);
and U1472 (N_1472,In_308,In_140);
and U1473 (N_1473,In_440,In_164);
nor U1474 (N_1474,In_427,In_790);
nand U1475 (N_1475,In_114,In_820);
or U1476 (N_1476,In_567,In_301);
nor U1477 (N_1477,In_723,In_857);
or U1478 (N_1478,In_957,In_216);
nor U1479 (N_1479,In_988,In_162);
xor U1480 (N_1480,In_870,In_576);
nor U1481 (N_1481,In_394,In_661);
or U1482 (N_1482,In_912,In_941);
or U1483 (N_1483,In_352,In_686);
nand U1484 (N_1484,In_81,In_335);
and U1485 (N_1485,In_769,In_580);
and U1486 (N_1486,In_111,In_280);
nand U1487 (N_1487,In_648,In_903);
or U1488 (N_1488,In_995,In_999);
nand U1489 (N_1489,In_379,In_933);
nor U1490 (N_1490,In_187,In_571);
xor U1491 (N_1491,In_360,In_899);
or U1492 (N_1492,In_555,In_64);
and U1493 (N_1493,In_368,In_946);
and U1494 (N_1494,In_75,In_795);
and U1495 (N_1495,In_747,In_883);
or U1496 (N_1496,In_890,In_834);
nand U1497 (N_1497,In_335,In_98);
nand U1498 (N_1498,In_37,In_930);
nor U1499 (N_1499,In_300,In_914);
and U1500 (N_1500,In_734,In_516);
and U1501 (N_1501,In_838,In_455);
nand U1502 (N_1502,In_72,In_911);
nor U1503 (N_1503,In_272,In_588);
or U1504 (N_1504,In_287,In_713);
and U1505 (N_1505,In_852,In_205);
and U1506 (N_1506,In_998,In_983);
nor U1507 (N_1507,In_67,In_738);
nand U1508 (N_1508,In_687,In_919);
nor U1509 (N_1509,In_948,In_962);
nand U1510 (N_1510,In_687,In_679);
xor U1511 (N_1511,In_995,In_107);
and U1512 (N_1512,In_798,In_353);
or U1513 (N_1513,In_458,In_464);
and U1514 (N_1514,In_747,In_837);
nor U1515 (N_1515,In_127,In_880);
nand U1516 (N_1516,In_906,In_371);
and U1517 (N_1517,In_634,In_346);
or U1518 (N_1518,In_750,In_661);
or U1519 (N_1519,In_96,In_284);
nor U1520 (N_1520,In_985,In_74);
nand U1521 (N_1521,In_601,In_171);
or U1522 (N_1522,In_869,In_571);
or U1523 (N_1523,In_696,In_243);
and U1524 (N_1524,In_711,In_930);
nor U1525 (N_1525,In_606,In_685);
and U1526 (N_1526,In_669,In_416);
and U1527 (N_1527,In_712,In_719);
nor U1528 (N_1528,In_808,In_609);
nand U1529 (N_1529,In_674,In_220);
or U1530 (N_1530,In_368,In_904);
or U1531 (N_1531,In_872,In_335);
xor U1532 (N_1532,In_100,In_485);
and U1533 (N_1533,In_892,In_604);
nand U1534 (N_1534,In_636,In_887);
or U1535 (N_1535,In_350,In_43);
and U1536 (N_1536,In_137,In_496);
or U1537 (N_1537,In_831,In_211);
or U1538 (N_1538,In_258,In_740);
nor U1539 (N_1539,In_320,In_999);
nand U1540 (N_1540,In_24,In_198);
nor U1541 (N_1541,In_364,In_564);
and U1542 (N_1542,In_87,In_366);
nor U1543 (N_1543,In_695,In_903);
and U1544 (N_1544,In_862,In_280);
and U1545 (N_1545,In_152,In_340);
and U1546 (N_1546,In_89,In_738);
and U1547 (N_1547,In_148,In_985);
nor U1548 (N_1548,In_749,In_259);
nand U1549 (N_1549,In_726,In_723);
nor U1550 (N_1550,In_685,In_895);
xnor U1551 (N_1551,In_890,In_226);
nand U1552 (N_1552,In_878,In_616);
xnor U1553 (N_1553,In_565,In_386);
or U1554 (N_1554,In_899,In_419);
nor U1555 (N_1555,In_140,In_965);
and U1556 (N_1556,In_773,In_642);
and U1557 (N_1557,In_643,In_480);
or U1558 (N_1558,In_900,In_324);
and U1559 (N_1559,In_784,In_378);
xor U1560 (N_1560,In_411,In_836);
nand U1561 (N_1561,In_873,In_75);
nor U1562 (N_1562,In_205,In_173);
nor U1563 (N_1563,In_436,In_979);
or U1564 (N_1564,In_133,In_113);
or U1565 (N_1565,In_155,In_576);
nand U1566 (N_1566,In_881,In_39);
and U1567 (N_1567,In_208,In_897);
or U1568 (N_1568,In_544,In_153);
nand U1569 (N_1569,In_634,In_646);
xor U1570 (N_1570,In_792,In_665);
and U1571 (N_1571,In_637,In_80);
nor U1572 (N_1572,In_830,In_525);
and U1573 (N_1573,In_708,In_622);
nor U1574 (N_1574,In_324,In_212);
and U1575 (N_1575,In_449,In_121);
or U1576 (N_1576,In_443,In_521);
and U1577 (N_1577,In_336,In_705);
and U1578 (N_1578,In_693,In_467);
nor U1579 (N_1579,In_160,In_355);
or U1580 (N_1580,In_677,In_920);
nor U1581 (N_1581,In_4,In_234);
nand U1582 (N_1582,In_892,In_383);
and U1583 (N_1583,In_780,In_11);
nor U1584 (N_1584,In_239,In_30);
nor U1585 (N_1585,In_784,In_370);
nor U1586 (N_1586,In_861,In_883);
and U1587 (N_1587,In_353,In_169);
nand U1588 (N_1588,In_981,In_367);
nor U1589 (N_1589,In_474,In_181);
nand U1590 (N_1590,In_267,In_787);
or U1591 (N_1591,In_592,In_180);
nor U1592 (N_1592,In_632,In_787);
nor U1593 (N_1593,In_105,In_52);
nor U1594 (N_1594,In_564,In_835);
nand U1595 (N_1595,In_833,In_920);
and U1596 (N_1596,In_924,In_30);
or U1597 (N_1597,In_883,In_901);
nor U1598 (N_1598,In_930,In_625);
nand U1599 (N_1599,In_495,In_815);
or U1600 (N_1600,In_435,In_480);
nor U1601 (N_1601,In_614,In_290);
or U1602 (N_1602,In_143,In_328);
nand U1603 (N_1603,In_866,In_647);
or U1604 (N_1604,In_379,In_636);
or U1605 (N_1605,In_949,In_989);
nor U1606 (N_1606,In_701,In_781);
and U1607 (N_1607,In_271,In_244);
and U1608 (N_1608,In_382,In_629);
nand U1609 (N_1609,In_955,In_378);
and U1610 (N_1610,In_971,In_183);
nand U1611 (N_1611,In_456,In_66);
or U1612 (N_1612,In_362,In_250);
nor U1613 (N_1613,In_800,In_933);
nand U1614 (N_1614,In_621,In_580);
nor U1615 (N_1615,In_145,In_710);
or U1616 (N_1616,In_507,In_180);
nor U1617 (N_1617,In_545,In_336);
and U1618 (N_1618,In_698,In_454);
and U1619 (N_1619,In_276,In_2);
nand U1620 (N_1620,In_272,In_75);
nand U1621 (N_1621,In_843,In_273);
nor U1622 (N_1622,In_824,In_531);
nand U1623 (N_1623,In_15,In_307);
nor U1624 (N_1624,In_665,In_329);
or U1625 (N_1625,In_859,In_711);
nand U1626 (N_1626,In_763,In_393);
nand U1627 (N_1627,In_438,In_207);
nor U1628 (N_1628,In_510,In_704);
nor U1629 (N_1629,In_833,In_717);
nor U1630 (N_1630,In_134,In_332);
and U1631 (N_1631,In_578,In_187);
xor U1632 (N_1632,In_695,In_696);
nor U1633 (N_1633,In_497,In_379);
nor U1634 (N_1634,In_348,In_435);
or U1635 (N_1635,In_833,In_778);
xnor U1636 (N_1636,In_217,In_185);
nand U1637 (N_1637,In_314,In_439);
nand U1638 (N_1638,In_904,In_549);
or U1639 (N_1639,In_200,In_493);
and U1640 (N_1640,In_953,In_619);
nand U1641 (N_1641,In_241,In_370);
nor U1642 (N_1642,In_262,In_860);
or U1643 (N_1643,In_490,In_93);
nor U1644 (N_1644,In_916,In_367);
nor U1645 (N_1645,In_697,In_335);
or U1646 (N_1646,In_11,In_286);
and U1647 (N_1647,In_398,In_663);
or U1648 (N_1648,In_297,In_234);
and U1649 (N_1649,In_259,In_870);
nor U1650 (N_1650,In_374,In_575);
nor U1651 (N_1651,In_538,In_372);
nand U1652 (N_1652,In_350,In_267);
nand U1653 (N_1653,In_584,In_92);
nor U1654 (N_1654,In_551,In_757);
and U1655 (N_1655,In_532,In_155);
nor U1656 (N_1656,In_354,In_559);
nor U1657 (N_1657,In_239,In_556);
and U1658 (N_1658,In_577,In_382);
nor U1659 (N_1659,In_185,In_691);
nand U1660 (N_1660,In_846,In_606);
or U1661 (N_1661,In_84,In_782);
or U1662 (N_1662,In_647,In_914);
and U1663 (N_1663,In_133,In_164);
or U1664 (N_1664,In_941,In_952);
and U1665 (N_1665,In_31,In_416);
xor U1666 (N_1666,In_746,In_376);
nand U1667 (N_1667,In_327,In_127);
nor U1668 (N_1668,In_529,In_623);
nor U1669 (N_1669,In_905,In_510);
nor U1670 (N_1670,In_665,In_489);
and U1671 (N_1671,In_515,In_357);
nand U1672 (N_1672,In_545,In_439);
or U1673 (N_1673,In_492,In_845);
nand U1674 (N_1674,In_967,In_16);
nor U1675 (N_1675,In_612,In_241);
or U1676 (N_1676,In_783,In_704);
nand U1677 (N_1677,In_74,In_649);
nor U1678 (N_1678,In_621,In_237);
nor U1679 (N_1679,In_441,In_498);
or U1680 (N_1680,In_297,In_375);
nand U1681 (N_1681,In_994,In_250);
and U1682 (N_1682,In_387,In_409);
nand U1683 (N_1683,In_572,In_584);
or U1684 (N_1684,In_121,In_296);
nor U1685 (N_1685,In_101,In_403);
or U1686 (N_1686,In_965,In_408);
or U1687 (N_1687,In_380,In_566);
or U1688 (N_1688,In_68,In_901);
nand U1689 (N_1689,In_341,In_487);
or U1690 (N_1690,In_556,In_788);
nor U1691 (N_1691,In_297,In_621);
nand U1692 (N_1692,In_297,In_951);
and U1693 (N_1693,In_167,In_38);
nand U1694 (N_1694,In_358,In_827);
nand U1695 (N_1695,In_865,In_719);
nor U1696 (N_1696,In_912,In_1);
or U1697 (N_1697,In_820,In_641);
nor U1698 (N_1698,In_881,In_487);
or U1699 (N_1699,In_886,In_8);
nor U1700 (N_1700,In_495,In_923);
or U1701 (N_1701,In_176,In_682);
and U1702 (N_1702,In_259,In_894);
nor U1703 (N_1703,In_218,In_90);
nand U1704 (N_1704,In_820,In_75);
and U1705 (N_1705,In_378,In_38);
and U1706 (N_1706,In_166,In_5);
and U1707 (N_1707,In_716,In_980);
and U1708 (N_1708,In_521,In_759);
or U1709 (N_1709,In_169,In_290);
or U1710 (N_1710,In_647,In_240);
nand U1711 (N_1711,In_244,In_633);
nor U1712 (N_1712,In_526,In_940);
nand U1713 (N_1713,In_210,In_606);
nand U1714 (N_1714,In_945,In_607);
and U1715 (N_1715,In_393,In_96);
nand U1716 (N_1716,In_317,In_446);
nand U1717 (N_1717,In_579,In_907);
nor U1718 (N_1718,In_384,In_671);
and U1719 (N_1719,In_79,In_615);
and U1720 (N_1720,In_93,In_946);
or U1721 (N_1721,In_79,In_135);
nand U1722 (N_1722,In_272,In_929);
and U1723 (N_1723,In_704,In_24);
or U1724 (N_1724,In_2,In_861);
or U1725 (N_1725,In_515,In_382);
or U1726 (N_1726,In_972,In_824);
or U1727 (N_1727,In_822,In_957);
nor U1728 (N_1728,In_484,In_705);
or U1729 (N_1729,In_100,In_9);
or U1730 (N_1730,In_20,In_589);
and U1731 (N_1731,In_579,In_518);
or U1732 (N_1732,In_396,In_12);
and U1733 (N_1733,In_152,In_796);
and U1734 (N_1734,In_546,In_149);
and U1735 (N_1735,In_947,In_843);
or U1736 (N_1736,In_629,In_466);
or U1737 (N_1737,In_809,In_320);
or U1738 (N_1738,In_61,In_744);
and U1739 (N_1739,In_534,In_15);
or U1740 (N_1740,In_649,In_966);
nor U1741 (N_1741,In_160,In_678);
nand U1742 (N_1742,In_552,In_836);
and U1743 (N_1743,In_299,In_11);
nand U1744 (N_1744,In_15,In_219);
xor U1745 (N_1745,In_626,In_505);
nand U1746 (N_1746,In_453,In_928);
or U1747 (N_1747,In_559,In_853);
or U1748 (N_1748,In_57,In_571);
or U1749 (N_1749,In_681,In_273);
nor U1750 (N_1750,In_601,In_927);
nand U1751 (N_1751,In_280,In_78);
xnor U1752 (N_1752,In_439,In_525);
or U1753 (N_1753,In_210,In_641);
and U1754 (N_1754,In_273,In_480);
and U1755 (N_1755,In_828,In_985);
and U1756 (N_1756,In_461,In_223);
nand U1757 (N_1757,In_297,In_877);
nor U1758 (N_1758,In_391,In_871);
or U1759 (N_1759,In_430,In_62);
nor U1760 (N_1760,In_408,In_852);
and U1761 (N_1761,In_110,In_71);
or U1762 (N_1762,In_8,In_70);
nor U1763 (N_1763,In_97,In_527);
or U1764 (N_1764,In_7,In_459);
and U1765 (N_1765,In_475,In_216);
nand U1766 (N_1766,In_434,In_463);
and U1767 (N_1767,In_944,In_64);
nand U1768 (N_1768,In_212,In_477);
nand U1769 (N_1769,In_749,In_792);
nand U1770 (N_1770,In_446,In_613);
or U1771 (N_1771,In_331,In_181);
nand U1772 (N_1772,In_342,In_351);
nand U1773 (N_1773,In_56,In_880);
and U1774 (N_1774,In_667,In_995);
and U1775 (N_1775,In_73,In_674);
and U1776 (N_1776,In_827,In_334);
nor U1777 (N_1777,In_571,In_215);
or U1778 (N_1778,In_380,In_3);
and U1779 (N_1779,In_266,In_711);
nor U1780 (N_1780,In_241,In_410);
nand U1781 (N_1781,In_185,In_598);
and U1782 (N_1782,In_899,In_452);
or U1783 (N_1783,In_530,In_947);
nand U1784 (N_1784,In_388,In_670);
xnor U1785 (N_1785,In_363,In_543);
and U1786 (N_1786,In_639,In_856);
nor U1787 (N_1787,In_377,In_887);
nor U1788 (N_1788,In_245,In_588);
and U1789 (N_1789,In_247,In_734);
and U1790 (N_1790,In_693,In_353);
nor U1791 (N_1791,In_194,In_129);
nand U1792 (N_1792,In_292,In_818);
or U1793 (N_1793,In_305,In_107);
nor U1794 (N_1794,In_124,In_558);
nor U1795 (N_1795,In_661,In_744);
and U1796 (N_1796,In_579,In_815);
nand U1797 (N_1797,In_655,In_711);
or U1798 (N_1798,In_885,In_593);
and U1799 (N_1799,In_859,In_740);
nor U1800 (N_1800,In_442,In_468);
nor U1801 (N_1801,In_161,In_950);
nand U1802 (N_1802,In_652,In_341);
and U1803 (N_1803,In_875,In_198);
nor U1804 (N_1804,In_81,In_850);
nand U1805 (N_1805,In_334,In_106);
nor U1806 (N_1806,In_572,In_206);
or U1807 (N_1807,In_895,In_291);
nor U1808 (N_1808,In_720,In_650);
nor U1809 (N_1809,In_734,In_679);
or U1810 (N_1810,In_386,In_784);
and U1811 (N_1811,In_118,In_841);
and U1812 (N_1812,In_565,In_311);
or U1813 (N_1813,In_554,In_935);
and U1814 (N_1814,In_284,In_916);
nor U1815 (N_1815,In_640,In_672);
or U1816 (N_1816,In_764,In_626);
and U1817 (N_1817,In_444,In_155);
and U1818 (N_1818,In_3,In_296);
nor U1819 (N_1819,In_166,In_457);
and U1820 (N_1820,In_71,In_969);
nor U1821 (N_1821,In_318,In_998);
and U1822 (N_1822,In_254,In_502);
xor U1823 (N_1823,In_233,In_548);
and U1824 (N_1824,In_461,In_848);
nor U1825 (N_1825,In_265,In_294);
nand U1826 (N_1826,In_993,In_105);
nor U1827 (N_1827,In_390,In_423);
or U1828 (N_1828,In_17,In_235);
or U1829 (N_1829,In_410,In_418);
nor U1830 (N_1830,In_563,In_291);
or U1831 (N_1831,In_972,In_583);
nand U1832 (N_1832,In_540,In_243);
or U1833 (N_1833,In_727,In_172);
and U1834 (N_1834,In_272,In_999);
nand U1835 (N_1835,In_536,In_355);
nor U1836 (N_1836,In_824,In_148);
or U1837 (N_1837,In_971,In_802);
or U1838 (N_1838,In_426,In_174);
and U1839 (N_1839,In_204,In_284);
and U1840 (N_1840,In_397,In_561);
nand U1841 (N_1841,In_648,In_466);
or U1842 (N_1842,In_958,In_340);
nand U1843 (N_1843,In_27,In_159);
nand U1844 (N_1844,In_406,In_316);
nor U1845 (N_1845,In_712,In_450);
or U1846 (N_1846,In_37,In_370);
or U1847 (N_1847,In_721,In_406);
and U1848 (N_1848,In_527,In_907);
and U1849 (N_1849,In_91,In_184);
or U1850 (N_1850,In_390,In_358);
xor U1851 (N_1851,In_771,In_438);
nor U1852 (N_1852,In_106,In_339);
and U1853 (N_1853,In_214,In_249);
nor U1854 (N_1854,In_41,In_58);
nand U1855 (N_1855,In_880,In_932);
or U1856 (N_1856,In_704,In_801);
and U1857 (N_1857,In_939,In_807);
nor U1858 (N_1858,In_532,In_23);
nand U1859 (N_1859,In_619,In_918);
nor U1860 (N_1860,In_736,In_926);
or U1861 (N_1861,In_77,In_141);
nand U1862 (N_1862,In_484,In_880);
nor U1863 (N_1863,In_661,In_943);
nand U1864 (N_1864,In_948,In_503);
nor U1865 (N_1865,In_321,In_711);
nand U1866 (N_1866,In_13,In_855);
nand U1867 (N_1867,In_470,In_733);
or U1868 (N_1868,In_717,In_173);
and U1869 (N_1869,In_236,In_633);
nor U1870 (N_1870,In_896,In_74);
nand U1871 (N_1871,In_560,In_16);
or U1872 (N_1872,In_943,In_830);
and U1873 (N_1873,In_95,In_138);
nor U1874 (N_1874,In_188,In_877);
or U1875 (N_1875,In_65,In_735);
and U1876 (N_1876,In_86,In_641);
nor U1877 (N_1877,In_105,In_777);
nor U1878 (N_1878,In_714,In_510);
nor U1879 (N_1879,In_454,In_689);
nor U1880 (N_1880,In_755,In_124);
nand U1881 (N_1881,In_538,In_105);
or U1882 (N_1882,In_575,In_471);
nor U1883 (N_1883,In_483,In_658);
and U1884 (N_1884,In_992,In_892);
nor U1885 (N_1885,In_257,In_751);
or U1886 (N_1886,In_309,In_424);
and U1887 (N_1887,In_14,In_748);
nor U1888 (N_1888,In_838,In_746);
and U1889 (N_1889,In_770,In_889);
nor U1890 (N_1890,In_601,In_99);
nand U1891 (N_1891,In_771,In_672);
and U1892 (N_1892,In_966,In_368);
nand U1893 (N_1893,In_167,In_125);
nor U1894 (N_1894,In_83,In_468);
and U1895 (N_1895,In_590,In_726);
nand U1896 (N_1896,In_337,In_276);
nand U1897 (N_1897,In_14,In_912);
and U1898 (N_1898,In_248,In_435);
and U1899 (N_1899,In_469,In_586);
and U1900 (N_1900,In_485,In_206);
nand U1901 (N_1901,In_91,In_223);
or U1902 (N_1902,In_919,In_123);
nand U1903 (N_1903,In_419,In_411);
or U1904 (N_1904,In_163,In_399);
and U1905 (N_1905,In_165,In_655);
or U1906 (N_1906,In_973,In_866);
xnor U1907 (N_1907,In_217,In_396);
and U1908 (N_1908,In_364,In_528);
and U1909 (N_1909,In_590,In_724);
or U1910 (N_1910,In_861,In_209);
and U1911 (N_1911,In_832,In_57);
or U1912 (N_1912,In_357,In_181);
nor U1913 (N_1913,In_294,In_252);
nor U1914 (N_1914,In_161,In_652);
or U1915 (N_1915,In_768,In_186);
nor U1916 (N_1916,In_649,In_249);
nand U1917 (N_1917,In_63,In_65);
and U1918 (N_1918,In_887,In_40);
or U1919 (N_1919,In_271,In_546);
or U1920 (N_1920,In_512,In_655);
and U1921 (N_1921,In_870,In_703);
and U1922 (N_1922,In_591,In_717);
and U1923 (N_1923,In_600,In_713);
or U1924 (N_1924,In_193,In_962);
or U1925 (N_1925,In_163,In_79);
and U1926 (N_1926,In_372,In_912);
nor U1927 (N_1927,In_331,In_346);
nand U1928 (N_1928,In_843,In_354);
and U1929 (N_1929,In_615,In_858);
nor U1930 (N_1930,In_363,In_54);
and U1931 (N_1931,In_545,In_151);
or U1932 (N_1932,In_0,In_899);
nor U1933 (N_1933,In_427,In_719);
nor U1934 (N_1934,In_651,In_58);
nor U1935 (N_1935,In_739,In_766);
nor U1936 (N_1936,In_800,In_55);
nor U1937 (N_1937,In_215,In_342);
or U1938 (N_1938,In_64,In_347);
and U1939 (N_1939,In_829,In_652);
nor U1940 (N_1940,In_775,In_942);
xor U1941 (N_1941,In_884,In_999);
nor U1942 (N_1942,In_104,In_301);
or U1943 (N_1943,In_169,In_469);
or U1944 (N_1944,In_503,In_262);
and U1945 (N_1945,In_764,In_211);
or U1946 (N_1946,In_253,In_623);
nand U1947 (N_1947,In_968,In_623);
or U1948 (N_1948,In_757,In_40);
or U1949 (N_1949,In_397,In_591);
or U1950 (N_1950,In_548,In_880);
or U1951 (N_1951,In_680,In_104);
or U1952 (N_1952,In_151,In_885);
and U1953 (N_1953,In_873,In_931);
nand U1954 (N_1954,In_350,In_739);
and U1955 (N_1955,In_791,In_844);
or U1956 (N_1956,In_862,In_957);
nand U1957 (N_1957,In_12,In_119);
nor U1958 (N_1958,In_991,In_832);
and U1959 (N_1959,In_669,In_395);
nor U1960 (N_1960,In_929,In_77);
nor U1961 (N_1961,In_716,In_113);
or U1962 (N_1962,In_812,In_54);
and U1963 (N_1963,In_906,In_745);
nand U1964 (N_1964,In_694,In_383);
nor U1965 (N_1965,In_647,In_949);
nor U1966 (N_1966,In_878,In_448);
nand U1967 (N_1967,In_806,In_704);
nand U1968 (N_1968,In_6,In_260);
nand U1969 (N_1969,In_804,In_298);
nand U1970 (N_1970,In_686,In_19);
nor U1971 (N_1971,In_852,In_600);
and U1972 (N_1972,In_527,In_217);
nor U1973 (N_1973,In_205,In_130);
or U1974 (N_1974,In_642,In_861);
or U1975 (N_1975,In_257,In_752);
or U1976 (N_1976,In_732,In_78);
nand U1977 (N_1977,In_797,In_115);
nand U1978 (N_1978,In_358,In_874);
nor U1979 (N_1979,In_288,In_37);
nand U1980 (N_1980,In_211,In_625);
nor U1981 (N_1981,In_128,In_971);
and U1982 (N_1982,In_242,In_238);
nand U1983 (N_1983,In_984,In_616);
or U1984 (N_1984,In_285,In_167);
or U1985 (N_1985,In_87,In_683);
or U1986 (N_1986,In_670,In_846);
nor U1987 (N_1987,In_413,In_358);
nor U1988 (N_1988,In_317,In_979);
or U1989 (N_1989,In_763,In_815);
nand U1990 (N_1990,In_957,In_909);
nand U1991 (N_1991,In_546,In_333);
nor U1992 (N_1992,In_926,In_179);
and U1993 (N_1993,In_919,In_424);
nand U1994 (N_1994,In_935,In_702);
nor U1995 (N_1995,In_556,In_567);
or U1996 (N_1996,In_158,In_798);
nor U1997 (N_1997,In_652,In_120);
or U1998 (N_1998,In_92,In_755);
or U1999 (N_1999,In_918,In_314);
nand U2000 (N_2000,N_86,N_1944);
and U2001 (N_2001,N_846,N_1274);
and U2002 (N_2002,N_88,N_85);
and U2003 (N_2003,N_417,N_1926);
nand U2004 (N_2004,N_1940,N_840);
or U2005 (N_2005,N_1629,N_1083);
nor U2006 (N_2006,N_47,N_987);
nand U2007 (N_2007,N_956,N_1857);
or U2008 (N_2008,N_1820,N_887);
or U2009 (N_2009,N_786,N_266);
nor U2010 (N_2010,N_842,N_1033);
and U2011 (N_2011,N_1790,N_1863);
nand U2012 (N_2012,N_905,N_863);
nand U2013 (N_2013,N_1414,N_1688);
nand U2014 (N_2014,N_183,N_1171);
or U2015 (N_2015,N_652,N_1600);
or U2016 (N_2016,N_402,N_1040);
or U2017 (N_2017,N_216,N_1708);
nor U2018 (N_2018,N_675,N_495);
or U2019 (N_2019,N_22,N_923);
nand U2020 (N_2020,N_681,N_899);
and U2021 (N_2021,N_1938,N_1750);
nand U2022 (N_2022,N_1272,N_1775);
xnor U2023 (N_2023,N_548,N_1215);
nand U2024 (N_2024,N_725,N_1675);
or U2025 (N_2025,N_166,N_434);
and U2026 (N_2026,N_167,N_184);
and U2027 (N_2027,N_148,N_695);
or U2028 (N_2028,N_1304,N_1713);
and U2029 (N_2029,N_1946,N_1764);
and U2030 (N_2030,N_1167,N_674);
and U2031 (N_2031,N_1170,N_1021);
nand U2032 (N_2032,N_300,N_454);
nor U2033 (N_2033,N_691,N_1140);
or U2034 (N_2034,N_673,N_724);
nor U2035 (N_2035,N_1253,N_1475);
nor U2036 (N_2036,N_506,N_1914);
nand U2037 (N_2037,N_741,N_253);
nand U2038 (N_2038,N_962,N_1486);
or U2039 (N_2039,N_188,N_1130);
nor U2040 (N_2040,N_818,N_731);
nor U2041 (N_2041,N_1206,N_912);
xor U2042 (N_2042,N_12,N_74);
and U2043 (N_2043,N_294,N_38);
xor U2044 (N_2044,N_102,N_1386);
or U2045 (N_2045,N_1590,N_1331);
or U2046 (N_2046,N_589,N_505);
and U2047 (N_2047,N_1730,N_1110);
or U2048 (N_2048,N_20,N_1570);
nand U2049 (N_2049,N_207,N_464);
xnor U2050 (N_2050,N_229,N_1611);
and U2051 (N_2051,N_901,N_221);
and U2052 (N_2052,N_1227,N_1250);
or U2053 (N_2053,N_764,N_1067);
nor U2054 (N_2054,N_1280,N_99);
or U2055 (N_2055,N_1180,N_814);
nand U2056 (N_2056,N_1222,N_432);
or U2057 (N_2057,N_1886,N_1120);
nand U2058 (N_2058,N_1329,N_140);
and U2059 (N_2059,N_306,N_1893);
nand U2060 (N_2060,N_1562,N_1522);
and U2061 (N_2061,N_356,N_778);
nand U2062 (N_2062,N_1044,N_1614);
nand U2063 (N_2063,N_1121,N_664);
xnor U2064 (N_2064,N_1073,N_1768);
nor U2065 (N_2065,N_1723,N_1363);
nor U2066 (N_2066,N_1582,N_896);
and U2067 (N_2067,N_954,N_580);
nand U2068 (N_2068,N_240,N_325);
or U2069 (N_2069,N_1419,N_1450);
nor U2070 (N_2070,N_1126,N_1022);
nand U2071 (N_2071,N_806,N_1341);
and U2072 (N_2072,N_1578,N_256);
and U2073 (N_2073,N_1879,N_1109);
nand U2074 (N_2074,N_133,N_1816);
and U2075 (N_2075,N_1338,N_303);
xor U2076 (N_2076,N_1855,N_555);
nand U2077 (N_2077,N_1667,N_628);
and U2078 (N_2078,N_1279,N_1906);
or U2079 (N_2079,N_359,N_1814);
and U2080 (N_2080,N_271,N_1326);
xnor U2081 (N_2081,N_1057,N_1860);
nand U2082 (N_2082,N_1846,N_1849);
or U2083 (N_2083,N_235,N_1664);
or U2084 (N_2084,N_960,N_1512);
or U2085 (N_2085,N_1469,N_1742);
nor U2086 (N_2086,N_596,N_1544);
nand U2087 (N_2087,N_1618,N_1737);
and U2088 (N_2088,N_1704,N_329);
and U2089 (N_2089,N_53,N_1769);
and U2090 (N_2090,N_1308,N_1869);
nand U2091 (N_2091,N_1878,N_1736);
and U2092 (N_2092,N_576,N_635);
nand U2093 (N_2093,N_1901,N_1592);
or U2094 (N_2094,N_1690,N_1795);
nand U2095 (N_2095,N_1276,N_493);
or U2096 (N_2096,N_791,N_394);
nor U2097 (N_2097,N_1453,N_570);
nand U2098 (N_2098,N_83,N_1984);
nand U2099 (N_2099,N_513,N_261);
and U2100 (N_2100,N_1931,N_1043);
nand U2101 (N_2101,N_976,N_208);
xnor U2102 (N_2102,N_1706,N_1612);
nand U2103 (N_2103,N_526,N_345);
nor U2104 (N_2104,N_350,N_696);
nor U2105 (N_2105,N_699,N_639);
nand U2106 (N_2106,N_683,N_1184);
or U2107 (N_2107,N_593,N_105);
or U2108 (N_2108,N_572,N_1828);
nand U2109 (N_2109,N_1594,N_1373);
or U2110 (N_2110,N_1097,N_1298);
or U2111 (N_2111,N_1151,N_1166);
nand U2112 (N_2112,N_751,N_18);
xnor U2113 (N_2113,N_585,N_997);
nand U2114 (N_2114,N_1301,N_217);
and U2115 (N_2115,N_1413,N_1471);
xor U2116 (N_2116,N_621,N_1316);
or U2117 (N_2117,N_1754,N_1444);
and U2118 (N_2118,N_1609,N_1672);
or U2119 (N_2119,N_1342,N_1064);
and U2120 (N_2120,N_868,N_1965);
or U2121 (N_2121,N_120,N_733);
xnor U2122 (N_2122,N_433,N_162);
or U2123 (N_2123,N_1913,N_799);
or U2124 (N_2124,N_1942,N_150);
nor U2125 (N_2125,N_446,N_693);
nand U2126 (N_2126,N_66,N_128);
nor U2127 (N_2127,N_1104,N_813);
nand U2128 (N_2128,N_1464,N_659);
and U2129 (N_2129,N_1610,N_755);
or U2130 (N_2130,N_1972,N_753);
nor U2131 (N_2131,N_736,N_865);
or U2132 (N_2132,N_1756,N_1840);
or U2133 (N_2133,N_1183,N_514);
or U2134 (N_2134,N_1069,N_784);
and U2135 (N_2135,N_169,N_474);
nand U2136 (N_2136,N_1302,N_1241);
nor U2137 (N_2137,N_1422,N_265);
nor U2138 (N_2138,N_223,N_528);
and U2139 (N_2139,N_599,N_1002);
nand U2140 (N_2140,N_1431,N_415);
nor U2141 (N_2141,N_1597,N_1026);
nand U2142 (N_2142,N_1321,N_1966);
nand U2143 (N_2143,N_1516,N_1988);
nor U2144 (N_2144,N_1583,N_139);
or U2145 (N_2145,N_1251,N_1693);
nor U2146 (N_2146,N_149,N_595);
and U2147 (N_2147,N_1229,N_1613);
and U2148 (N_2148,N_283,N_1446);
nor U2149 (N_2149,N_765,N_1927);
nand U2150 (N_2150,N_663,N_682);
and U2151 (N_2151,N_904,N_92);
nand U2152 (N_2152,N_1156,N_1369);
or U2153 (N_2153,N_1681,N_812);
and U2154 (N_2154,N_1564,N_1237);
or U2155 (N_2155,N_878,N_129);
nor U2156 (N_2156,N_1347,N_1461);
nand U2157 (N_2157,N_930,N_479);
and U2158 (N_2158,N_200,N_214);
nand U2159 (N_2159,N_1786,N_116);
and U2160 (N_2160,N_1105,N_436);
or U2161 (N_2161,N_1416,N_1652);
nor U2162 (N_2162,N_1697,N_951);
nand U2163 (N_2163,N_158,N_131);
or U2164 (N_2164,N_1649,N_24);
nand U2165 (N_2165,N_1725,N_365);
or U2166 (N_2166,N_703,N_145);
nor U2167 (N_2167,N_1314,N_993);
and U2168 (N_2168,N_71,N_62);
or U2169 (N_2169,N_503,N_445);
or U2170 (N_2170,N_112,N_1330);
or U2171 (N_2171,N_1604,N_1454);
and U2172 (N_2172,N_800,N_219);
or U2173 (N_2173,N_369,N_344);
or U2174 (N_2174,N_971,N_701);
nand U2175 (N_2175,N_520,N_134);
and U2176 (N_2176,N_1394,N_1545);
nor U2177 (N_2177,N_1969,N_636);
or U2178 (N_2178,N_141,N_1114);
and U2179 (N_2179,N_1962,N_893);
nand U2180 (N_2180,N_544,N_1729);
or U2181 (N_2181,N_592,N_1970);
nor U2182 (N_2182,N_859,N_1560);
or U2183 (N_2183,N_480,N_1382);
or U2184 (N_2184,N_1565,N_1949);
nor U2185 (N_2185,N_911,N_1325);
nor U2186 (N_2186,N_117,N_114);
xnor U2187 (N_2187,N_364,N_309);
xnor U2188 (N_2188,N_1261,N_298);
and U2189 (N_2189,N_561,N_1967);
or U2190 (N_2190,N_525,N_13);
or U2191 (N_2191,N_1306,N_195);
nor U2192 (N_2192,N_209,N_1839);
nor U2193 (N_2193,N_1287,N_281);
nand U2194 (N_2194,N_1624,N_1157);
nor U2195 (N_2195,N_1749,N_1502);
or U2196 (N_2196,N_1975,N_1835);
nor U2197 (N_2197,N_130,N_1344);
or U2198 (N_2198,N_1062,N_860);
or U2199 (N_2199,N_1936,N_762);
and U2200 (N_2200,N_823,N_1550);
and U2201 (N_2201,N_1520,N_1596);
and U2202 (N_2202,N_850,N_1848);
or U2203 (N_2203,N_1559,N_1717);
and U2204 (N_2204,N_510,N_1054);
and U2205 (N_2205,N_259,N_705);
nor U2206 (N_2206,N_940,N_0);
and U2207 (N_2207,N_648,N_1755);
nand U2208 (N_2208,N_1854,N_552);
nand U2209 (N_2209,N_371,N_1438);
nor U2210 (N_2210,N_1147,N_1143);
or U2211 (N_2211,N_456,N_1493);
and U2212 (N_2212,N_398,N_1925);
and U2213 (N_2213,N_1881,N_460);
nand U2214 (N_2214,N_611,N_407);
and U2215 (N_2215,N_26,N_647);
nor U2216 (N_2216,N_632,N_808);
nand U2217 (N_2217,N_212,N_656);
nand U2218 (N_2218,N_824,N_1960);
nor U2219 (N_2219,N_734,N_1456);
or U2220 (N_2220,N_180,N_1865);
and U2221 (N_2221,N_1117,N_1617);
and U2222 (N_2222,N_154,N_1154);
nor U2223 (N_2223,N_1794,N_605);
or U2224 (N_2224,N_387,N_676);
nand U2225 (N_2225,N_1765,N_1499);
nor U2226 (N_2226,N_989,N_1626);
and U2227 (N_2227,N_1451,N_1716);
or U2228 (N_2228,N_1248,N_629);
nor U2229 (N_2229,N_1116,N_1015);
and U2230 (N_2230,N_1579,N_1265);
nand U2231 (N_2231,N_107,N_759);
nand U2232 (N_2232,N_442,N_1599);
and U2233 (N_2233,N_1483,N_1513);
nor U2234 (N_2234,N_945,N_1952);
and U2235 (N_2235,N_575,N_363);
and U2236 (N_2236,N_462,N_190);
nand U2237 (N_2237,N_1551,N_512);
nand U2238 (N_2238,N_1976,N_1247);
nor U2239 (N_2239,N_773,N_1379);
or U2240 (N_2240,N_54,N_1005);
and U2241 (N_2241,N_1996,N_1286);
or U2242 (N_2242,N_630,N_1296);
or U2243 (N_2243,N_1294,N_143);
nor U2244 (N_2244,N_710,N_1176);
nor U2245 (N_2245,N_518,N_849);
xnor U2246 (N_2246,N_471,N_43);
or U2247 (N_2247,N_553,N_832);
nor U2248 (N_2248,N_1554,N_412);
and U2249 (N_2249,N_1616,N_1809);
or U2250 (N_2250,N_343,N_355);
or U2251 (N_2251,N_1362,N_1683);
and U2252 (N_2252,N_714,N_393);
nor U2253 (N_2253,N_1734,N_368);
nor U2254 (N_2254,N_1397,N_428);
nor U2255 (N_2255,N_98,N_616);
nor U2256 (N_2256,N_702,N_1384);
nand U2257 (N_2257,N_643,N_1941);
and U2258 (N_2258,N_1887,N_1255);
nor U2259 (N_2259,N_1799,N_807);
or U2260 (N_2260,N_1646,N_96);
nand U2261 (N_2261,N_943,N_3);
nor U2262 (N_2262,N_1696,N_280);
nor U2263 (N_2263,N_1220,N_1478);
nor U2264 (N_2264,N_450,N_227);
nor U2265 (N_2265,N_299,N_1415);
and U2266 (N_2266,N_1532,N_1024);
nor U2267 (N_2267,N_941,N_247);
nand U2268 (N_2268,N_587,N_672);
nand U2269 (N_2269,N_583,N_67);
nand U2270 (N_2270,N_1084,N_1213);
and U2271 (N_2271,N_921,N_79);
and U2272 (N_2272,N_1739,N_1139);
or U2273 (N_2273,N_882,N_1779);
and U2274 (N_2274,N_973,N_1694);
or U2275 (N_2275,N_551,N_944);
nand U2276 (N_2276,N_631,N_396);
or U2277 (N_2277,N_401,N_1523);
and U2278 (N_2278,N_1270,N_1071);
or U2279 (N_2279,N_1217,N_1317);
nor U2280 (N_2280,N_1094,N_1871);
and U2281 (N_2281,N_346,N_826);
nor U2282 (N_2282,N_1922,N_1258);
nor U2283 (N_2283,N_178,N_523);
nor U2284 (N_2284,N_1098,N_706);
nand U2285 (N_2285,N_151,N_1907);
and U2286 (N_2286,N_668,N_210);
nor U2287 (N_2287,N_1133,N_524);
nor U2288 (N_2288,N_1636,N_1945);
nand U2289 (N_2289,N_1273,N_408);
and U2290 (N_2290,N_841,N_1702);
or U2291 (N_2291,N_1986,N_392);
or U2292 (N_2292,N_1312,N_658);
xor U2293 (N_2293,N_1254,N_1621);
nand U2294 (N_2294,N_2,N_649);
and U2295 (N_2295,N_1519,N_1541);
nand U2296 (N_2296,N_239,N_925);
nor U2297 (N_2297,N_307,N_521);
nor U2298 (N_2298,N_1197,N_929);
nor U2299 (N_2299,N_830,N_186);
and U2300 (N_2300,N_1465,N_248);
or U2301 (N_2301,N_678,N_1808);
nand U2302 (N_2302,N_1390,N_374);
or U2303 (N_2303,N_995,N_665);
and U2304 (N_2304,N_1086,N_895);
nand U2305 (N_2305,N_1365,N_317);
nand U2306 (N_2306,N_934,N_349);
nand U2307 (N_2307,N_861,N_427);
or U2308 (N_2308,N_1305,N_1676);
or U2309 (N_2309,N_856,N_33);
or U2310 (N_2310,N_890,N_1804);
nor U2311 (N_2311,N_1787,N_65);
nor U2312 (N_2312,N_1123,N_1531);
or U2313 (N_2313,N_1577,N_566);
or U2314 (N_2314,N_1797,N_439);
or U2315 (N_2315,N_1412,N_558);
nor U2316 (N_2316,N_1008,N_836);
or U2317 (N_2317,N_740,N_1684);
or U2318 (N_2318,N_1263,N_745);
or U2319 (N_2319,N_1640,N_625);
xor U2320 (N_2320,N_254,N_1028);
nor U2321 (N_2321,N_827,N_1953);
or U2322 (N_2322,N_1993,N_1818);
and U2323 (N_2323,N_707,N_1266);
nand U2324 (N_2324,N_203,N_782);
nand U2325 (N_2325,N_802,N_1977);
nor U2326 (N_2326,N_1549,N_1175);
or U2327 (N_2327,N_100,N_1371);
or U2328 (N_2328,N_597,N_1671);
nor U2329 (N_2329,N_1426,N_968);
nand U2330 (N_2330,N_1920,N_63);
or U2331 (N_2331,N_179,N_508);
nand U2332 (N_2332,N_1353,N_977);
or U2333 (N_2333,N_1351,N_1858);
or U2334 (N_2334,N_571,N_332);
or U2335 (N_2335,N_1715,N_501);
nor U2336 (N_2336,N_1072,N_378);
nor U2337 (N_2337,N_57,N_1245);
or U2338 (N_2338,N_242,N_756);
nor U2339 (N_2339,N_1627,N_1368);
nand U2340 (N_2340,N_498,N_1246);
nor U2341 (N_2341,N_1595,N_1585);
nor U2342 (N_2342,N_1481,N_637);
nor U2343 (N_2343,N_1070,N_1670);
and U2344 (N_2344,N_386,N_1884);
nand U2345 (N_2345,N_233,N_961);
nand U2346 (N_2346,N_1101,N_384);
nor U2347 (N_2347,N_626,N_704);
and U2348 (N_2348,N_1673,N_1211);
nand U2349 (N_2349,N_1662,N_477);
nor U2350 (N_2350,N_1911,N_153);
and U2351 (N_2351,N_926,N_1603);
and U2352 (N_2352,N_1805,N_924);
nor U2353 (N_2353,N_711,N_979);
nor U2354 (N_2354,N_1574,N_1815);
xnor U2355 (N_2355,N_422,N_1271);
xnor U2356 (N_2356,N_1643,N_48);
and U2357 (N_2357,N_763,N_867);
nand U2358 (N_2358,N_645,N_1692);
nand U2359 (N_2359,N_275,N_1186);
or U2360 (N_2360,N_1556,N_1058);
or U2361 (N_2361,N_601,N_604);
or U2362 (N_2362,N_1555,N_1168);
and U2363 (N_2363,N_1908,N_152);
and U2364 (N_2364,N_1987,N_11);
nand U2365 (N_2365,N_1623,N_302);
or U2366 (N_2366,N_788,N_395);
and U2367 (N_2367,N_52,N_103);
and U2368 (N_2368,N_1743,N_1047);
or U2369 (N_2369,N_602,N_310);
or U2370 (N_2370,N_1909,N_1476);
nand U2371 (N_2371,N_796,N_892);
or U2372 (N_2372,N_404,N_1146);
nand U2373 (N_2373,N_466,N_4);
or U2374 (N_2374,N_328,N_1872);
or U2375 (N_2375,N_746,N_918);
nor U2376 (N_2376,N_1902,N_366);
nor U2377 (N_2377,N_447,N_1081);
nand U2378 (N_2378,N_1727,N_1127);
nand U2379 (N_2379,N_1018,N_568);
nand U2380 (N_2380,N_749,N_1437);
and U2381 (N_2381,N_1686,N_776);
or U2382 (N_2382,N_1598,N_1447);
nand U2383 (N_2383,N_420,N_1772);
nand U2384 (N_2384,N_1877,N_231);
nand U2385 (N_2385,N_949,N_1687);
and U2386 (N_2386,N_321,N_482);
or U2387 (N_2387,N_1359,N_1607);
and U2388 (N_2388,N_1773,N_124);
and U2389 (N_2389,N_1292,N_40);
nor U2390 (N_2390,N_312,N_1158);
or U2391 (N_2391,N_967,N_1788);
nand U2392 (N_2392,N_232,N_487);
nor U2393 (N_2393,N_1882,N_1992);
or U2394 (N_2394,N_1537,N_273);
nor U2395 (N_2395,N_1830,N_1129);
nand U2396 (N_2396,N_998,N_1642);
nand U2397 (N_2397,N_1075,N_258);
or U2398 (N_2398,N_1517,N_1700);
and U2399 (N_2399,N_1731,N_641);
nor U2400 (N_2400,N_192,N_1542);
or U2401 (N_2401,N_488,N_483);
xor U2402 (N_2402,N_72,N_1060);
nor U2403 (N_2403,N_947,N_1710);
and U2404 (N_2404,N_1231,N_29);
nand U2405 (N_2405,N_230,N_1488);
and U2406 (N_2406,N_1457,N_515);
and U2407 (N_2407,N_1034,N_774);
nand U2408 (N_2408,N_457,N_476);
or U2409 (N_2409,N_1495,N_1943);
or U2410 (N_2410,N_1315,N_472);
and U2411 (N_2411,N_975,N_1707);
nand U2412 (N_2412,N_1806,N_1165);
and U2413 (N_2413,N_1289,N_1588);
or U2414 (N_2414,N_1496,N_1866);
nand U2415 (N_2415,N_1290,N_564);
nor U2416 (N_2416,N_339,N_1979);
nor U2417 (N_2417,N_1791,N_1712);
or U2418 (N_2418,N_839,N_1695);
or U2419 (N_2419,N_633,N_252);
nor U2420 (N_2420,N_463,N_623);
nor U2421 (N_2421,N_1540,N_137);
nand U2422 (N_2422,N_1398,N_61);
or U2423 (N_2423,N_958,N_500);
nor U2424 (N_2424,N_7,N_950);
nor U2425 (N_2425,N_1356,N_1239);
nor U2426 (N_2426,N_361,N_1467);
nand U2427 (N_2427,N_1747,N_41);
nor U2428 (N_2428,N_1148,N_399);
nor U2429 (N_2429,N_136,N_1722);
or U2430 (N_2430,N_1999,N_295);
nand U2431 (N_2431,N_787,N_1844);
and U2432 (N_2432,N_1961,N_1510);
or U2433 (N_2433,N_1441,N_160);
nand U2434 (N_2434,N_610,N_453);
or U2435 (N_2435,N_1277,N_142);
nor U2436 (N_2436,N_1548,N_1605);
nand U2437 (N_2437,N_1096,N_390);
nand U2438 (N_2438,N_1163,N_620);
or U2439 (N_2439,N_39,N_517);
nand U2440 (N_2440,N_494,N_1494);
or U2441 (N_2441,N_1930,N_1323);
nand U2442 (N_2442,N_638,N_1763);
nor U2443 (N_2443,N_1430,N_400);
or U2444 (N_2444,N_809,N_1501);
nor U2445 (N_2445,N_1894,N_978);
nor U2446 (N_2446,N_1917,N_694);
nor U2447 (N_2447,N_1401,N_1291);
nor U2448 (N_2448,N_1630,N_411);
and U2449 (N_2449,N_1701,N_1918);
nand U2450 (N_2450,N_1087,N_1448);
or U2451 (N_2451,N_748,N_1219);
nor U2452 (N_2452,N_563,N_449);
or U2453 (N_2453,N_64,N_1826);
and U2454 (N_2454,N_9,N_441);
nand U2455 (N_2455,N_1023,N_1051);
nor U2456 (N_2456,N_1234,N_1784);
and U2457 (N_2457,N_922,N_1421);
nor U2458 (N_2458,N_1631,N_1460);
nor U2459 (N_2459,N_1526,N_196);
and U2460 (N_2460,N_1653,N_222);
nor U2461 (N_2461,N_270,N_970);
and U2462 (N_2462,N_1014,N_475);
nor U2463 (N_2463,N_104,N_1746);
nand U2464 (N_2464,N_1740,N_1758);
and U2465 (N_2465,N_1851,N_1776);
nor U2466 (N_2466,N_497,N_1632);
and U2467 (N_2467,N_1796,N_1395);
and U2468 (N_2468,N_1903,N_1682);
and U2469 (N_2469,N_874,N_851);
nand U2470 (N_2470,N_173,N_218);
nor U2471 (N_2471,N_138,N_1455);
or U2472 (N_2472,N_942,N_1593);
and U2473 (N_2473,N_1714,N_1619);
or U2474 (N_2474,N_268,N_1155);
or U2475 (N_2475,N_1997,N_461);
or U2476 (N_2476,N_1181,N_1487);
nor U2477 (N_2477,N_770,N_1406);
xor U2478 (N_2478,N_224,N_1159);
nand U2479 (N_2479,N_499,N_669);
nor U2480 (N_2480,N_421,N_805);
nor U2481 (N_2481,N_1821,N_397);
xor U2482 (N_2482,N_742,N_304);
nor U2483 (N_2483,N_1678,N_1425);
or U2484 (N_2484,N_972,N_58);
and U2485 (N_2485,N_822,N_1408);
and U2486 (N_2486,N_1659,N_1334);
nor U2487 (N_2487,N_1989,N_56);
nand U2488 (N_2488,N_409,N_334);
and U2489 (N_2489,N_290,N_467);
nand U2490 (N_2490,N_189,N_1337);
nand U2491 (N_2491,N_249,N_341);
and U2492 (N_2492,N_747,N_829);
or U2493 (N_2493,N_1663,N_1571);
or U2494 (N_2494,N_1569,N_1898);
or U2495 (N_2495,N_1521,N_305);
nand U2496 (N_2496,N_790,N_69);
and U2497 (N_2497,N_320,N_594);
nand U2498 (N_2498,N_95,N_654);
or U2499 (N_2499,N_1399,N_185);
nor U2500 (N_2500,N_781,N_1536);
nand U2501 (N_2501,N_110,N_579);
and U2502 (N_2502,N_319,N_1720);
and U2503 (N_2503,N_844,N_1050);
and U2504 (N_2504,N_614,N_1169);
or U2505 (N_2505,N_1751,N_313);
or U2506 (N_2506,N_535,N_1196);
or U2507 (N_2507,N_795,N_36);
nand U2508 (N_2508,N_1738,N_1132);
and U2509 (N_2509,N_1500,N_1873);
nand U2510 (N_2510,N_1557,N_990);
and U2511 (N_2511,N_23,N_1012);
and U2512 (N_2512,N_156,N_1509);
nor U2513 (N_2513,N_1374,N_1506);
or U2514 (N_2514,N_713,N_1240);
or U2515 (N_2515,N_992,N_348);
and U2516 (N_2516,N_1576,N_1124);
or U2517 (N_2517,N_952,N_1392);
nand U2518 (N_2518,N_1134,N_478);
or U2519 (N_2519,N_410,N_1311);
and U2520 (N_2520,N_1400,N_1777);
nand U2521 (N_2521,N_1332,N_1178);
nand U2522 (N_2522,N_144,N_423);
nand U2523 (N_2523,N_871,N_1466);
nand U2524 (N_2524,N_1077,N_855);
nand U2525 (N_2525,N_262,N_490);
nand U2526 (N_2526,N_1119,N_1587);
nor U2527 (N_2527,N_1733,N_82);
or U2528 (N_2528,N_1726,N_607);
xor U2529 (N_2529,N_1568,N_225);
and U2530 (N_2530,N_1709,N_1224);
and U2531 (N_2531,N_991,N_1090);
or U2532 (N_2532,N_168,N_679);
xnor U2533 (N_2533,N_1985,N_889);
or U2534 (N_2534,N_1434,N_123);
nor U2535 (N_2535,N_965,N_1088);
or U2536 (N_2536,N_539,N_980);
and U2537 (N_2537,N_1396,N_838);
or U2538 (N_2538,N_627,N_1971);
nand U2539 (N_2539,N_1093,N_1679);
or U2540 (N_2540,N_202,N_847);
and U2541 (N_2541,N_1393,N_1783);
and U2542 (N_2542,N_1053,N_615);
nand U2543 (N_2543,N_127,N_1812);
nand U2544 (N_2544,N_1209,N_1324);
nor U2545 (N_2545,N_49,N_1378);
nand U2546 (N_2546,N_1061,N_170);
and U2547 (N_2547,N_547,N_1994);
or U2548 (N_2548,N_815,N_1238);
nand U2549 (N_2549,N_640,N_1459);
and U2550 (N_2550,N_1472,N_245);
nor U2551 (N_2551,N_1990,N_1327);
nor U2552 (N_2552,N_1845,N_1982);
and U2553 (N_2553,N_817,N_89);
nor U2554 (N_2554,N_780,N_282);
nand U2555 (N_2555,N_1514,N_16);
or U2556 (N_2556,N_1563,N_709);
nand U2557 (N_2557,N_1748,N_1904);
nor U2558 (N_2558,N_831,N_1160);
nor U2559 (N_2559,N_920,N_985);
and U2560 (N_2560,N_1389,N_1935);
nand U2561 (N_2561,N_879,N_1661);
or U2562 (N_2562,N_1602,N_1364);
nand U2563 (N_2563,N_122,N_1829);
nand U2564 (N_2564,N_1862,N_697);
nand U2565 (N_2565,N_1644,N_1320);
nor U2566 (N_2566,N_1528,N_1198);
and U2567 (N_2567,N_391,N_171);
or U2568 (N_2568,N_1628,N_1089);
or U2569 (N_2569,N_81,N_1402);
nor U2570 (N_2570,N_1256,N_1432);
nand U2571 (N_2571,N_172,N_1766);
nand U2572 (N_2572,N_870,N_1335);
and U2573 (N_2573,N_1003,N_1793);
and U2574 (N_2574,N_541,N_293);
or U2575 (N_2575,N_354,N_999);
or U2576 (N_2576,N_1173,N_21);
or U2577 (N_2577,N_353,N_1868);
nand U2578 (N_2578,N_606,N_612);
and U2579 (N_2579,N_1482,N_296);
nand U2580 (N_2580,N_590,N_1063);
or U2581 (N_2581,N_1191,N_529);
or U2582 (N_2582,N_1037,N_455);
nand U2583 (N_2583,N_1032,N_1009);
nor U2584 (N_2584,N_569,N_1162);
nand U2585 (N_2585,N_1233,N_1439);
nand U2586 (N_2586,N_279,N_175);
nand U2587 (N_2587,N_1638,N_516);
nand U2588 (N_2588,N_1136,N_28);
and U2589 (N_2589,N_1883,N_199);
or U2590 (N_2590,N_1606,N_769);
nor U2591 (N_2591,N_650,N_1954);
nand U2592 (N_2592,N_91,N_737);
nand U2593 (N_2593,N_1719,N_1284);
xor U2594 (N_2594,N_660,N_567);
xnor U2595 (N_2595,N_848,N_1346);
or U2596 (N_2596,N_1436,N_1208);
and U2597 (N_2597,N_726,N_1428);
or U2598 (N_2598,N_468,N_1625);
or U2599 (N_2599,N_284,N_1354);
or U2600 (N_2600,N_932,N_382);
or U2601 (N_2601,N_426,N_1182);
or U2602 (N_2602,N_1435,N_1031);
or U2603 (N_2603,N_1336,N_1349);
or U2604 (N_2604,N_1059,N_886);
and U2605 (N_2605,N_201,N_559);
nand U2606 (N_2606,N_388,N_845);
or U2607 (N_2607,N_1744,N_966);
or U2608 (N_2608,N_819,N_496);
and U2609 (N_2609,N_291,N_732);
and U2610 (N_2610,N_1867,N_1185);
nand U2611 (N_2611,N_549,N_276);
nand U2612 (N_2612,N_519,N_1870);
or U2613 (N_2613,N_260,N_1131);
nand U2614 (N_2614,N_1955,N_1484);
nand U2615 (N_2615,N_1885,N_351);
nor U2616 (N_2616,N_527,N_1891);
nor U2617 (N_2617,N_1677,N_1318);
nand U2618 (N_2618,N_730,N_1202);
nand U2619 (N_2619,N_504,N_1463);
nand U2620 (N_2620,N_1491,N_25);
xnor U2621 (N_2621,N_862,N_228);
or U2622 (N_2622,N_459,N_1216);
and U2623 (N_2623,N_285,N_443);
or U2624 (N_2624,N_161,N_1259);
and U2625 (N_2625,N_768,N_308);
nand U2626 (N_2626,N_1055,N_546);
or U2627 (N_2627,N_1916,N_1691);
or U2628 (N_2628,N_1080,N_352);
nand U2629 (N_2629,N_877,N_1843);
or U2630 (N_2630,N_1888,N_1201);
and U2631 (N_2631,N_1339,N_335);
and U2632 (N_2632,N_73,N_1230);
nand U2633 (N_2633,N_6,N_383);
or U2634 (N_2634,N_1367,N_1900);
and U2635 (N_2635,N_994,N_1300);
nand U2636 (N_2636,N_661,N_1760);
nor U2637 (N_2637,N_452,N_1038);
nor U2638 (N_2638,N_1288,N_872);
nor U2639 (N_2639,N_1001,N_1995);
and U2640 (N_2640,N_1479,N_19);
or U2641 (N_2641,N_1543,N_181);
or U2642 (N_2642,N_1172,N_507);
nor U2643 (N_2643,N_1194,N_1504);
nor U2644 (N_2644,N_758,N_1998);
xnor U2645 (N_2645,N_1910,N_828);
or U2646 (N_2646,N_1823,N_125);
nor U2647 (N_2647,N_1100,N_1832);
nand U2648 (N_2648,N_1118,N_1407);
or U2649 (N_2649,N_716,N_727);
nand U2650 (N_2650,N_1838,N_1534);
or U2651 (N_2651,N_1068,N_1689);
nand U2652 (N_2652,N_667,N_206);
or U2653 (N_2653,N_609,N_577);
and U2654 (N_2654,N_931,N_1388);
xnor U2655 (N_2655,N_1190,N_801);
and U2656 (N_2656,N_1417,N_573);
nand U2657 (N_2657,N_1780,N_1745);
nand U2658 (N_2658,N_157,N_1552);
and U2659 (N_2659,N_1125,N_618);
nor U2660 (N_2660,N_1572,N_919);
or U2661 (N_2661,N_1924,N_1381);
and U2662 (N_2662,N_1852,N_1391);
and U2663 (N_2663,N_94,N_948);
nor U2664 (N_2664,N_1007,N_1409);
or U2665 (N_2665,N_311,N_928);
and U2666 (N_2666,N_600,N_1699);
and U2667 (N_2667,N_1959,N_301);
nor U2668 (N_2668,N_1427,N_581);
and U2669 (N_2669,N_1584,N_486);
and U2670 (N_2670,N_1633,N_634);
and U2671 (N_2671,N_1785,N_543);
nor U2672 (N_2672,N_1620,N_419);
or U2673 (N_2673,N_106,N_885);
nor U2674 (N_2674,N_113,N_1650);
nand U2675 (N_2675,N_1641,N_1187);
nor U2676 (N_2676,N_680,N_389);
and U2677 (N_2677,N_534,N_833);
and U2678 (N_2678,N_1297,N_761);
nor U2679 (N_2679,N_1978,N_984);
nand U2680 (N_2680,N_1669,N_14);
nor U2681 (N_2681,N_121,N_834);
or U2682 (N_2682,N_1375,N_416);
nor U2683 (N_2683,N_1950,N_718);
nor U2684 (N_2684,N_405,N_1242);
or U2685 (N_2685,N_584,N_1876);
and U2686 (N_2686,N_1781,N_241);
nand U2687 (N_2687,N_338,N_565);
and U2688 (N_2688,N_779,N_720);
nor U2689 (N_2689,N_1313,N_530);
and U2690 (N_2690,N_1387,N_689);
nor U2691 (N_2691,N_1199,N_1899);
xnor U2692 (N_2692,N_362,N_1307);
or U2693 (N_2693,N_470,N_622);
or U2694 (N_2694,N_739,N_884);
nand U2695 (N_2695,N_858,N_274);
and U2696 (N_2696,N_93,N_174);
nor U2697 (N_2697,N_1411,N_1929);
or U2698 (N_2698,N_909,N_686);
and U2699 (N_2699,N_852,N_1189);
or U2700 (N_2700,N_1340,N_1892);
and U2701 (N_2701,N_1810,N_1218);
and U2702 (N_2702,N_1933,N_358);
or U2703 (N_2703,N_1462,N_619);
nand U2704 (N_2704,N_1529,N_1905);
and U2705 (N_2705,N_670,N_286);
nor U2706 (N_2706,N_917,N_1964);
or U2707 (N_2707,N_1921,N_1041);
nand U2708 (N_2708,N_97,N_1477);
and U2709 (N_2709,N_719,N_1645);
nand U2710 (N_2710,N_698,N_176);
and U2711 (N_2711,N_700,N_955);
and U2712 (N_2712,N_1759,N_1833);
and U2713 (N_2713,N_1575,N_603);
and U2714 (N_2714,N_1767,N_1405);
and U2715 (N_2715,N_974,N_1092);
and U2716 (N_2716,N_1153,N_76);
and U2717 (N_2717,N_376,N_413);
xor U2718 (N_2718,N_1078,N_1824);
and U2719 (N_2719,N_772,N_1065);
or U2720 (N_2720,N_75,N_1827);
or U2721 (N_2721,N_1912,N_1035);
or U2722 (N_2722,N_37,N_869);
or U2723 (N_2723,N_1380,N_1282);
nor U2724 (N_2724,N_1957,N_915);
nand U2725 (N_2725,N_1226,N_1762);
and U2726 (N_2726,N_226,N_1046);
or U2727 (N_2727,N_1535,N_1214);
or U2728 (N_2728,N_1511,N_1179);
or U2729 (N_2729,N_684,N_78);
or U2730 (N_2730,N_582,N_30);
and U2731 (N_2731,N_316,N_333);
and U2732 (N_2732,N_1525,N_1983);
nor U2733 (N_2733,N_837,N_322);
nor U2734 (N_2734,N_1836,N_1586);
and U2735 (N_2735,N_1801,N_1262);
nand U2736 (N_2736,N_492,N_792);
or U2737 (N_2737,N_789,N_794);
or U2738 (N_2738,N_1267,N_77);
nor U2739 (N_2739,N_1660,N_1842);
and U2740 (N_2740,N_729,N_1951);
or U2741 (N_2741,N_1076,N_743);
or U2742 (N_2742,N_444,N_45);
nor U2743 (N_2743,N_1376,N_1923);
or U2744 (N_2744,N_1006,N_1106);
nor U2745 (N_2745,N_87,N_1637);
or U2746 (N_2746,N_810,N_1027);
nand U2747 (N_2747,N_1385,N_750);
nand U2748 (N_2748,N_377,N_437);
nand U2749 (N_2749,N_372,N_1666);
nand U2750 (N_2750,N_367,N_1711);
and U2751 (N_2751,N_938,N_723);
nand U2752 (N_2752,N_728,N_1647);
nor U2753 (N_2753,N_435,N_898);
and U2754 (N_2754,N_297,N_163);
nor U2755 (N_2755,N_1761,N_511);
and U2756 (N_2756,N_1480,N_1505);
or U2757 (N_2757,N_31,N_1333);
nand U2758 (N_2758,N_1225,N_1048);
and U2759 (N_2759,N_1200,N_1490);
xor U2760 (N_2760,N_1252,N_340);
nand U2761 (N_2761,N_1355,N_1141);
and U2762 (N_2762,N_1771,N_1260);
and U2763 (N_2763,N_1732,N_1703);
and U2764 (N_2764,N_1831,N_1403);
and U2765 (N_2765,N_811,N_900);
nor U2766 (N_2766,N_1580,N_1657);
or U2767 (N_2767,N_357,N_251);
or U2768 (N_2768,N_70,N_1192);
nand U2769 (N_2769,N_908,N_891);
nor U2770 (N_2770,N_722,N_347);
or U2771 (N_2771,N_1896,N_147);
and U2772 (N_2772,N_164,N_757);
nand U2773 (N_2773,N_1825,N_1377);
nor U2774 (N_2774,N_1658,N_988);
nand U2775 (N_2775,N_246,N_1591);
nor U2776 (N_2776,N_1221,N_5);
or U2777 (N_2777,N_653,N_1056);
or U2778 (N_2778,N_1947,N_873);
and U2779 (N_2779,N_211,N_1547);
or U2780 (N_2780,N_375,N_1188);
nand U2781 (N_2781,N_1019,N_288);
or U2782 (N_2782,N_717,N_708);
or U2783 (N_2783,N_1648,N_671);
or U2784 (N_2784,N_1091,N_1728);
nand U2785 (N_2785,N_642,N_370);
or U2786 (N_2786,N_690,N_1856);
or U2787 (N_2787,N_1895,N_937);
or U2788 (N_2788,N_927,N_1654);
or U2789 (N_2789,N_1608,N_798);
nand U2790 (N_2790,N_108,N_1753);
nand U2791 (N_2791,N_1656,N_1473);
or U2792 (N_2792,N_267,N_692);
nor U2793 (N_2793,N_1052,N_1232);
and U2794 (N_2794,N_1474,N_1880);
and U2795 (N_2795,N_1561,N_550);
nor U2796 (N_2796,N_205,N_767);
nand U2797 (N_2797,N_1782,N_381);
and U2798 (N_2798,N_1249,N_1010);
and U2799 (N_2799,N_1889,N_1573);
and U2800 (N_2800,N_820,N_913);
nand U2801 (N_2801,N_458,N_1113);
nand U2802 (N_2802,N_1497,N_1423);
nand U2803 (N_2803,N_10,N_1859);
nor U2804 (N_2804,N_752,N_1309);
nand U2805 (N_2805,N_1974,N_406);
nand U2806 (N_2806,N_1489,N_1128);
xor U2807 (N_2807,N_193,N_1698);
and U2808 (N_2808,N_1834,N_1303);
nor U2809 (N_2809,N_666,N_418);
nand U2810 (N_2810,N_1819,N_1752);
and U2811 (N_2811,N_277,N_1622);
or U2812 (N_2812,N_1207,N_1538);
and U2813 (N_2813,N_644,N_1358);
nand U2814 (N_2814,N_646,N_15);
or U2815 (N_2815,N_1508,N_484);
nor U2816 (N_2816,N_907,N_1195);
and U2817 (N_2817,N_1370,N_1212);
and U2818 (N_2818,N_119,N_473);
nor U2819 (N_2819,N_1085,N_1518);
nor U2820 (N_2820,N_1817,N_1352);
nor U2821 (N_2821,N_481,N_236);
or U2822 (N_2822,N_1470,N_1939);
xnor U2823 (N_2823,N_785,N_588);
and U2824 (N_2824,N_1567,N_843);
nor U2825 (N_2825,N_1980,N_1404);
nand U2826 (N_2826,N_1343,N_996);
nor U2827 (N_2827,N_1236,N_502);
nor U2828 (N_2828,N_1928,N_1800);
or U2829 (N_2829,N_556,N_1164);
nand U2830 (N_2830,N_982,N_981);
xnor U2831 (N_2831,N_1278,N_1348);
nand U2832 (N_2832,N_916,N_243);
or U2833 (N_2833,N_803,N_964);
and U2834 (N_2834,N_1115,N_1066);
or U2835 (N_2835,N_532,N_1458);
nand U2836 (N_2836,N_754,N_330);
or U2837 (N_2837,N_894,N_1674);
nor U2838 (N_2838,N_198,N_939);
or U2839 (N_2839,N_1802,N_557);
and U2840 (N_2840,N_1811,N_531);
or U2841 (N_2841,N_1036,N_1269);
and U2842 (N_2842,N_1932,N_1792);
nand U2843 (N_2843,N_465,N_536);
nand U2844 (N_2844,N_1442,N_1145);
or U2845 (N_2845,N_1937,N_1235);
nor U2846 (N_2846,N_560,N_875);
nor U2847 (N_2847,N_115,N_655);
nand U2848 (N_2848,N_657,N_1443);
nand U2849 (N_2849,N_257,N_1102);
or U2850 (N_2850,N_1122,N_883);
and U2851 (N_2851,N_1082,N_1721);
and U2852 (N_2852,N_1203,N_289);
or U2853 (N_2853,N_1468,N_1360);
nor U2854 (N_2854,N_1948,N_194);
xor U2855 (N_2855,N_1973,N_986);
or U2856 (N_2856,N_1310,N_1524);
and U2857 (N_2857,N_591,N_777);
nor U2858 (N_2858,N_866,N_1357);
nand U2859 (N_2859,N_1553,N_959);
or U2860 (N_2860,N_857,N_292);
and U2861 (N_2861,N_373,N_238);
nor U2862 (N_2862,N_425,N_90);
or U2863 (N_2863,N_1205,N_738);
nand U2864 (N_2864,N_1042,N_331);
or U2865 (N_2865,N_469,N_59);
and U2866 (N_2866,N_963,N_135);
and U2867 (N_2867,N_1045,N_766);
nor U2868 (N_2868,N_1107,N_651);
nand U2869 (N_2869,N_109,N_318);
or U2870 (N_2870,N_1897,N_379);
xor U2871 (N_2871,N_191,N_1099);
or U2872 (N_2872,N_1639,N_342);
and U2873 (N_2873,N_1533,N_430);
nand U2874 (N_2874,N_1013,N_489);
and U2875 (N_2875,N_403,N_1958);
nor U2876 (N_2876,N_1049,N_1345);
nor U2877 (N_2877,N_662,N_1135);
and U2878 (N_2878,N_220,N_1566);
or U2879 (N_2879,N_1498,N_1228);
nor U2880 (N_2880,N_1025,N_1546);
or U2881 (N_2881,N_1204,N_624);
nand U2882 (N_2882,N_111,N_27);
or U2883 (N_2883,N_17,N_578);
and U2884 (N_2884,N_60,N_42);
nand U2885 (N_2885,N_897,N_1705);
and U2886 (N_2886,N_1449,N_1152);
nand U2887 (N_2887,N_1177,N_617);
nand U2888 (N_2888,N_1,N_1527);
nand U2889 (N_2889,N_159,N_237);
nand U2890 (N_2890,N_44,N_1837);
nor U2891 (N_2891,N_1492,N_272);
or U2892 (N_2892,N_126,N_1017);
nand U2893 (N_2893,N_429,N_825);
and U2894 (N_2894,N_775,N_1452);
nand U2895 (N_2895,N_55,N_424);
nand U2896 (N_2896,N_132,N_1850);
or U2897 (N_2897,N_1789,N_1655);
nor U2898 (N_2898,N_215,N_876);
xor U2899 (N_2899,N_1798,N_1956);
or U2900 (N_2900,N_1864,N_197);
nand U2901 (N_2901,N_1112,N_1295);
or U2902 (N_2902,N_1161,N_1651);
nand U2903 (N_2903,N_1420,N_1095);
nand U2904 (N_2904,N_269,N_936);
nor U2905 (N_2905,N_1039,N_1503);
nor U2906 (N_2906,N_1515,N_1016);
xnor U2907 (N_2907,N_1144,N_1718);
nand U2908 (N_2908,N_906,N_1445);
nor U2909 (N_2909,N_101,N_880);
nand U2910 (N_2910,N_32,N_538);
or U2911 (N_2911,N_287,N_1111);
nand U2912 (N_2912,N_1210,N_182);
nor U2913 (N_2913,N_485,N_35);
or U2914 (N_2914,N_1963,N_1813);
nor U2915 (N_2915,N_1429,N_263);
and U2916 (N_2916,N_1665,N_545);
nand U2917 (N_2917,N_969,N_1530);
or U2918 (N_2918,N_677,N_8);
or U2919 (N_2919,N_1275,N_914);
nor U2920 (N_2920,N_760,N_118);
nand U2921 (N_2921,N_360,N_336);
nand U2922 (N_2922,N_853,N_1011);
or U2923 (N_2923,N_155,N_1149);
or U2924 (N_2924,N_68,N_554);
and U2925 (N_2925,N_1322,N_324);
nor U2926 (N_2926,N_1281,N_1934);
and U2927 (N_2927,N_314,N_685);
and U2928 (N_2928,N_1366,N_431);
nand U2929 (N_2929,N_1680,N_1138);
and U2930 (N_2930,N_34,N_1778);
and U2931 (N_2931,N_278,N_1150);
and U2932 (N_2932,N_1074,N_1485);
or U2933 (N_2933,N_204,N_1589);
nor U2934 (N_2934,N_84,N_1724);
or U2935 (N_2935,N_1919,N_1875);
nand U2936 (N_2936,N_327,N_562);
nand U2937 (N_2937,N_1861,N_451);
nand U2938 (N_2938,N_323,N_1103);
or U2939 (N_2939,N_1841,N_234);
or U2940 (N_2940,N_1424,N_213);
nand U2941 (N_2941,N_821,N_783);
xnor U2942 (N_2942,N_953,N_608);
nor U2943 (N_2943,N_1299,N_1601);
nor U2944 (N_2944,N_1264,N_1319);
or U2945 (N_2945,N_1174,N_1383);
nand U2946 (N_2946,N_1822,N_542);
or U2947 (N_2947,N_1968,N_735);
nand U2948 (N_2948,N_1915,N_1774);
and U2949 (N_2949,N_1361,N_933);
and U2950 (N_2950,N_688,N_51);
nor U2951 (N_2951,N_881,N_835);
or U2952 (N_2952,N_1079,N_146);
or U2953 (N_2953,N_797,N_414);
and U2954 (N_2954,N_1635,N_1108);
and U2955 (N_2955,N_1615,N_326);
nand U2956 (N_2956,N_1293,N_1991);
nor U2957 (N_2957,N_1507,N_1741);
nand U2958 (N_2958,N_1142,N_598);
and U2959 (N_2959,N_864,N_491);
nor U2960 (N_2960,N_1328,N_1410);
nand U2961 (N_2961,N_522,N_1685);
nor U2962 (N_2962,N_1668,N_1853);
or U2963 (N_2963,N_804,N_1874);
and U2964 (N_2964,N_1243,N_1803);
and U2965 (N_2965,N_1890,N_902);
nand U2966 (N_2966,N_1581,N_1257);
or U2967 (N_2967,N_448,N_264);
nor U2968 (N_2968,N_1418,N_721);
nor U2969 (N_2969,N_744,N_935);
or U2970 (N_2970,N_1433,N_1350);
and U2971 (N_2971,N_250,N_715);
nor U2972 (N_2972,N_816,N_793);
and U2973 (N_2973,N_385,N_910);
nor U2974 (N_2974,N_80,N_946);
nor U2975 (N_2975,N_1440,N_687);
nor U2976 (N_2976,N_380,N_574);
or U2977 (N_2977,N_165,N_244);
nor U2978 (N_2978,N_1735,N_903);
or U2979 (N_2979,N_1981,N_438);
or U2980 (N_2980,N_1757,N_1539);
nor U2981 (N_2981,N_50,N_187);
or U2982 (N_2982,N_613,N_1372);
nand U2983 (N_2983,N_337,N_1634);
nor U2984 (N_2984,N_1268,N_586);
nor U2985 (N_2985,N_854,N_888);
xnor U2986 (N_2986,N_315,N_771);
nand U2987 (N_2987,N_177,N_255);
or U2988 (N_2988,N_1020,N_1223);
or U2989 (N_2989,N_509,N_46);
or U2990 (N_2990,N_537,N_1770);
nor U2991 (N_2991,N_533,N_440);
and U2992 (N_2992,N_1807,N_712);
or U2993 (N_2993,N_1847,N_1029);
nand U2994 (N_2994,N_1558,N_1030);
nor U2995 (N_2995,N_1000,N_1244);
and U2996 (N_2996,N_540,N_1193);
nand U2997 (N_2997,N_1283,N_1285);
nor U2998 (N_2998,N_1137,N_1004);
nor U2999 (N_2999,N_983,N_957);
nor U3000 (N_3000,N_493,N_3);
and U3001 (N_3001,N_1309,N_1795);
nand U3002 (N_3002,N_1452,N_1703);
xnor U3003 (N_3003,N_366,N_208);
nor U3004 (N_3004,N_674,N_1664);
nand U3005 (N_3005,N_1794,N_1427);
or U3006 (N_3006,N_1136,N_1645);
or U3007 (N_3007,N_669,N_730);
and U3008 (N_3008,N_1795,N_1954);
nand U3009 (N_3009,N_724,N_879);
or U3010 (N_3010,N_1893,N_1478);
nor U3011 (N_3011,N_1902,N_1586);
or U3012 (N_3012,N_163,N_1835);
or U3013 (N_3013,N_1685,N_1532);
nand U3014 (N_3014,N_752,N_1281);
or U3015 (N_3015,N_940,N_1050);
nand U3016 (N_3016,N_1980,N_1122);
nor U3017 (N_3017,N_1015,N_1155);
or U3018 (N_3018,N_1602,N_543);
nor U3019 (N_3019,N_876,N_1856);
nor U3020 (N_3020,N_1151,N_1281);
nor U3021 (N_3021,N_1738,N_1710);
nand U3022 (N_3022,N_1604,N_305);
or U3023 (N_3023,N_1431,N_49);
nor U3024 (N_3024,N_293,N_605);
and U3025 (N_3025,N_698,N_603);
and U3026 (N_3026,N_547,N_683);
nor U3027 (N_3027,N_1427,N_0);
nor U3028 (N_3028,N_796,N_60);
nor U3029 (N_3029,N_1107,N_1500);
or U3030 (N_3030,N_554,N_1217);
nor U3031 (N_3031,N_1330,N_1329);
nor U3032 (N_3032,N_1228,N_776);
and U3033 (N_3033,N_975,N_1010);
or U3034 (N_3034,N_1878,N_829);
nor U3035 (N_3035,N_522,N_972);
and U3036 (N_3036,N_845,N_1416);
and U3037 (N_3037,N_834,N_837);
nand U3038 (N_3038,N_205,N_577);
and U3039 (N_3039,N_1358,N_86);
nor U3040 (N_3040,N_1586,N_300);
nand U3041 (N_3041,N_440,N_841);
nand U3042 (N_3042,N_1860,N_355);
and U3043 (N_3043,N_349,N_1107);
nor U3044 (N_3044,N_1580,N_607);
or U3045 (N_3045,N_92,N_936);
and U3046 (N_3046,N_813,N_1335);
or U3047 (N_3047,N_1913,N_470);
and U3048 (N_3048,N_549,N_365);
or U3049 (N_3049,N_826,N_539);
nand U3050 (N_3050,N_457,N_1701);
or U3051 (N_3051,N_806,N_740);
or U3052 (N_3052,N_1827,N_1748);
or U3053 (N_3053,N_123,N_1969);
nor U3054 (N_3054,N_541,N_99);
nor U3055 (N_3055,N_1127,N_1788);
nand U3056 (N_3056,N_1369,N_728);
nand U3057 (N_3057,N_789,N_1067);
or U3058 (N_3058,N_367,N_1690);
nor U3059 (N_3059,N_479,N_1471);
and U3060 (N_3060,N_1082,N_883);
nand U3061 (N_3061,N_1071,N_1756);
nor U3062 (N_3062,N_1130,N_974);
nand U3063 (N_3063,N_1568,N_551);
and U3064 (N_3064,N_736,N_1966);
nand U3065 (N_3065,N_133,N_1827);
and U3066 (N_3066,N_15,N_937);
and U3067 (N_3067,N_804,N_1368);
nand U3068 (N_3068,N_1401,N_1006);
and U3069 (N_3069,N_651,N_473);
and U3070 (N_3070,N_1558,N_1010);
or U3071 (N_3071,N_951,N_353);
nor U3072 (N_3072,N_1639,N_1988);
nand U3073 (N_3073,N_1298,N_1604);
nor U3074 (N_3074,N_133,N_704);
or U3075 (N_3075,N_1960,N_374);
and U3076 (N_3076,N_669,N_1793);
nor U3077 (N_3077,N_1205,N_1969);
and U3078 (N_3078,N_1480,N_619);
nor U3079 (N_3079,N_1600,N_1077);
or U3080 (N_3080,N_857,N_602);
nor U3081 (N_3081,N_115,N_245);
xnor U3082 (N_3082,N_1220,N_239);
nor U3083 (N_3083,N_664,N_1278);
nor U3084 (N_3084,N_1034,N_557);
nand U3085 (N_3085,N_292,N_1541);
nor U3086 (N_3086,N_875,N_874);
nand U3087 (N_3087,N_862,N_1528);
or U3088 (N_3088,N_1183,N_1627);
nand U3089 (N_3089,N_1226,N_1147);
or U3090 (N_3090,N_1005,N_231);
or U3091 (N_3091,N_1812,N_1507);
nand U3092 (N_3092,N_632,N_295);
nor U3093 (N_3093,N_662,N_82);
nor U3094 (N_3094,N_1778,N_1028);
nor U3095 (N_3095,N_1307,N_1529);
nor U3096 (N_3096,N_693,N_1370);
nor U3097 (N_3097,N_624,N_860);
nor U3098 (N_3098,N_1370,N_1151);
xnor U3099 (N_3099,N_1163,N_474);
and U3100 (N_3100,N_879,N_239);
or U3101 (N_3101,N_1007,N_768);
or U3102 (N_3102,N_1728,N_1160);
and U3103 (N_3103,N_1743,N_315);
and U3104 (N_3104,N_311,N_1859);
nand U3105 (N_3105,N_1124,N_152);
nand U3106 (N_3106,N_1925,N_1613);
and U3107 (N_3107,N_429,N_604);
or U3108 (N_3108,N_1362,N_899);
and U3109 (N_3109,N_1062,N_994);
or U3110 (N_3110,N_1804,N_1949);
or U3111 (N_3111,N_92,N_47);
and U3112 (N_3112,N_1319,N_1395);
nor U3113 (N_3113,N_1396,N_134);
nor U3114 (N_3114,N_7,N_1399);
nand U3115 (N_3115,N_609,N_1649);
and U3116 (N_3116,N_1700,N_187);
and U3117 (N_3117,N_1264,N_879);
nor U3118 (N_3118,N_1760,N_1956);
and U3119 (N_3119,N_1443,N_296);
nor U3120 (N_3120,N_1190,N_610);
or U3121 (N_3121,N_273,N_462);
nor U3122 (N_3122,N_607,N_1063);
nand U3123 (N_3123,N_519,N_1683);
nand U3124 (N_3124,N_571,N_1069);
or U3125 (N_3125,N_799,N_1257);
xnor U3126 (N_3126,N_319,N_1268);
nand U3127 (N_3127,N_1392,N_638);
nand U3128 (N_3128,N_1493,N_705);
and U3129 (N_3129,N_1936,N_32);
nand U3130 (N_3130,N_723,N_337);
xor U3131 (N_3131,N_1570,N_1281);
and U3132 (N_3132,N_621,N_860);
and U3133 (N_3133,N_424,N_1676);
nand U3134 (N_3134,N_1718,N_754);
nor U3135 (N_3135,N_979,N_625);
nand U3136 (N_3136,N_1702,N_562);
nor U3137 (N_3137,N_466,N_399);
or U3138 (N_3138,N_598,N_1488);
nand U3139 (N_3139,N_1254,N_55);
nand U3140 (N_3140,N_329,N_1777);
nand U3141 (N_3141,N_673,N_1092);
nand U3142 (N_3142,N_588,N_736);
and U3143 (N_3143,N_1535,N_1193);
nor U3144 (N_3144,N_1217,N_1593);
nor U3145 (N_3145,N_686,N_1965);
nor U3146 (N_3146,N_1324,N_3);
xnor U3147 (N_3147,N_44,N_465);
and U3148 (N_3148,N_677,N_1099);
nor U3149 (N_3149,N_464,N_583);
nand U3150 (N_3150,N_922,N_443);
or U3151 (N_3151,N_89,N_1760);
nor U3152 (N_3152,N_32,N_722);
nand U3153 (N_3153,N_491,N_655);
and U3154 (N_3154,N_726,N_1972);
nand U3155 (N_3155,N_501,N_1455);
and U3156 (N_3156,N_578,N_1159);
or U3157 (N_3157,N_816,N_1643);
nor U3158 (N_3158,N_667,N_1863);
or U3159 (N_3159,N_216,N_1386);
nand U3160 (N_3160,N_1534,N_1911);
nand U3161 (N_3161,N_1340,N_538);
or U3162 (N_3162,N_476,N_696);
nor U3163 (N_3163,N_1160,N_430);
nor U3164 (N_3164,N_97,N_276);
or U3165 (N_3165,N_1293,N_431);
or U3166 (N_3166,N_669,N_483);
nor U3167 (N_3167,N_434,N_1667);
nand U3168 (N_3168,N_355,N_696);
and U3169 (N_3169,N_229,N_1817);
nor U3170 (N_3170,N_81,N_1757);
xnor U3171 (N_3171,N_1005,N_856);
or U3172 (N_3172,N_1454,N_990);
or U3173 (N_3173,N_1908,N_171);
and U3174 (N_3174,N_467,N_556);
or U3175 (N_3175,N_1725,N_1887);
and U3176 (N_3176,N_791,N_1150);
or U3177 (N_3177,N_1485,N_1165);
nor U3178 (N_3178,N_859,N_831);
or U3179 (N_3179,N_22,N_1824);
nand U3180 (N_3180,N_168,N_1093);
nor U3181 (N_3181,N_41,N_535);
and U3182 (N_3182,N_348,N_871);
nand U3183 (N_3183,N_426,N_209);
nor U3184 (N_3184,N_698,N_1619);
and U3185 (N_3185,N_827,N_1242);
nand U3186 (N_3186,N_840,N_1138);
or U3187 (N_3187,N_1095,N_1096);
nor U3188 (N_3188,N_183,N_330);
nor U3189 (N_3189,N_1088,N_1237);
nand U3190 (N_3190,N_593,N_1965);
nand U3191 (N_3191,N_703,N_403);
or U3192 (N_3192,N_1426,N_721);
and U3193 (N_3193,N_709,N_166);
nor U3194 (N_3194,N_1089,N_1774);
nor U3195 (N_3195,N_453,N_91);
or U3196 (N_3196,N_1099,N_116);
or U3197 (N_3197,N_535,N_757);
or U3198 (N_3198,N_335,N_313);
xnor U3199 (N_3199,N_415,N_675);
and U3200 (N_3200,N_1833,N_1352);
nor U3201 (N_3201,N_1592,N_750);
xnor U3202 (N_3202,N_1545,N_1280);
nor U3203 (N_3203,N_163,N_1130);
nor U3204 (N_3204,N_1173,N_1799);
and U3205 (N_3205,N_1764,N_1075);
and U3206 (N_3206,N_125,N_1318);
nor U3207 (N_3207,N_109,N_730);
nor U3208 (N_3208,N_1301,N_1637);
and U3209 (N_3209,N_884,N_1926);
xor U3210 (N_3210,N_605,N_1201);
nand U3211 (N_3211,N_619,N_424);
and U3212 (N_3212,N_1482,N_1600);
nor U3213 (N_3213,N_174,N_1488);
and U3214 (N_3214,N_1191,N_700);
and U3215 (N_3215,N_1810,N_652);
nor U3216 (N_3216,N_1314,N_1193);
nor U3217 (N_3217,N_1540,N_1196);
or U3218 (N_3218,N_291,N_481);
nor U3219 (N_3219,N_1915,N_1436);
nor U3220 (N_3220,N_175,N_57);
or U3221 (N_3221,N_1157,N_1926);
xor U3222 (N_3222,N_1055,N_905);
nand U3223 (N_3223,N_249,N_1089);
nor U3224 (N_3224,N_324,N_1797);
nor U3225 (N_3225,N_1016,N_702);
nor U3226 (N_3226,N_1175,N_900);
nor U3227 (N_3227,N_1728,N_597);
nand U3228 (N_3228,N_161,N_410);
nand U3229 (N_3229,N_973,N_710);
nand U3230 (N_3230,N_936,N_1496);
and U3231 (N_3231,N_1544,N_444);
nand U3232 (N_3232,N_1562,N_1484);
nor U3233 (N_3233,N_226,N_1382);
or U3234 (N_3234,N_1719,N_1228);
nand U3235 (N_3235,N_202,N_33);
and U3236 (N_3236,N_159,N_320);
and U3237 (N_3237,N_507,N_1418);
nor U3238 (N_3238,N_259,N_890);
nor U3239 (N_3239,N_1560,N_926);
or U3240 (N_3240,N_767,N_1108);
or U3241 (N_3241,N_925,N_69);
nand U3242 (N_3242,N_849,N_1044);
nand U3243 (N_3243,N_1488,N_1648);
or U3244 (N_3244,N_1104,N_1381);
nand U3245 (N_3245,N_712,N_1532);
and U3246 (N_3246,N_1746,N_876);
nand U3247 (N_3247,N_1750,N_1662);
nor U3248 (N_3248,N_1930,N_1876);
and U3249 (N_3249,N_95,N_1324);
nor U3250 (N_3250,N_1971,N_1727);
or U3251 (N_3251,N_215,N_1243);
or U3252 (N_3252,N_403,N_661);
or U3253 (N_3253,N_72,N_360);
nor U3254 (N_3254,N_720,N_1408);
nor U3255 (N_3255,N_912,N_42);
nor U3256 (N_3256,N_823,N_982);
nand U3257 (N_3257,N_1495,N_610);
nor U3258 (N_3258,N_1283,N_1848);
xnor U3259 (N_3259,N_1004,N_370);
or U3260 (N_3260,N_1421,N_1734);
or U3261 (N_3261,N_1,N_1878);
or U3262 (N_3262,N_921,N_1486);
nand U3263 (N_3263,N_1271,N_1979);
nand U3264 (N_3264,N_800,N_1366);
nand U3265 (N_3265,N_528,N_1680);
and U3266 (N_3266,N_70,N_545);
and U3267 (N_3267,N_1186,N_39);
or U3268 (N_3268,N_203,N_1188);
nor U3269 (N_3269,N_1569,N_1906);
nand U3270 (N_3270,N_1205,N_994);
or U3271 (N_3271,N_403,N_821);
nand U3272 (N_3272,N_879,N_1638);
or U3273 (N_3273,N_1763,N_1048);
or U3274 (N_3274,N_1464,N_928);
or U3275 (N_3275,N_242,N_1147);
and U3276 (N_3276,N_176,N_1798);
nand U3277 (N_3277,N_1136,N_860);
nand U3278 (N_3278,N_1851,N_758);
or U3279 (N_3279,N_1558,N_1407);
nand U3280 (N_3280,N_586,N_1114);
and U3281 (N_3281,N_11,N_686);
nor U3282 (N_3282,N_1052,N_1376);
nand U3283 (N_3283,N_458,N_1275);
or U3284 (N_3284,N_1744,N_779);
nand U3285 (N_3285,N_633,N_1085);
nand U3286 (N_3286,N_486,N_539);
or U3287 (N_3287,N_1396,N_927);
or U3288 (N_3288,N_925,N_176);
nor U3289 (N_3289,N_147,N_1208);
nand U3290 (N_3290,N_817,N_1391);
nor U3291 (N_3291,N_1981,N_707);
nor U3292 (N_3292,N_308,N_1785);
or U3293 (N_3293,N_507,N_434);
or U3294 (N_3294,N_1886,N_1925);
xnor U3295 (N_3295,N_1642,N_1732);
and U3296 (N_3296,N_1841,N_1911);
nor U3297 (N_3297,N_491,N_724);
and U3298 (N_3298,N_1698,N_174);
nor U3299 (N_3299,N_1044,N_277);
or U3300 (N_3300,N_1268,N_298);
nor U3301 (N_3301,N_173,N_1298);
and U3302 (N_3302,N_1814,N_1254);
or U3303 (N_3303,N_782,N_1592);
nand U3304 (N_3304,N_156,N_1521);
nand U3305 (N_3305,N_1363,N_1159);
or U3306 (N_3306,N_543,N_270);
nand U3307 (N_3307,N_1599,N_914);
xnor U3308 (N_3308,N_1470,N_1144);
and U3309 (N_3309,N_987,N_942);
and U3310 (N_3310,N_134,N_791);
or U3311 (N_3311,N_564,N_1628);
nand U3312 (N_3312,N_390,N_686);
or U3313 (N_3313,N_433,N_41);
or U3314 (N_3314,N_1299,N_963);
xor U3315 (N_3315,N_618,N_881);
or U3316 (N_3316,N_1803,N_544);
or U3317 (N_3317,N_1139,N_760);
nand U3318 (N_3318,N_504,N_1726);
or U3319 (N_3319,N_641,N_1038);
and U3320 (N_3320,N_254,N_1833);
and U3321 (N_3321,N_1322,N_214);
nand U3322 (N_3322,N_367,N_1235);
nor U3323 (N_3323,N_1985,N_509);
nor U3324 (N_3324,N_1537,N_1021);
nor U3325 (N_3325,N_969,N_1951);
or U3326 (N_3326,N_541,N_91);
and U3327 (N_3327,N_36,N_1870);
or U3328 (N_3328,N_170,N_946);
or U3329 (N_3329,N_1076,N_1432);
or U3330 (N_3330,N_1690,N_691);
nor U3331 (N_3331,N_739,N_1515);
nor U3332 (N_3332,N_1793,N_1108);
xnor U3333 (N_3333,N_1964,N_240);
and U3334 (N_3334,N_907,N_1813);
and U3335 (N_3335,N_80,N_966);
nand U3336 (N_3336,N_1012,N_309);
nand U3337 (N_3337,N_1131,N_993);
xnor U3338 (N_3338,N_1416,N_1267);
nand U3339 (N_3339,N_501,N_1182);
and U3340 (N_3340,N_155,N_652);
or U3341 (N_3341,N_1387,N_279);
nor U3342 (N_3342,N_141,N_1243);
and U3343 (N_3343,N_685,N_539);
and U3344 (N_3344,N_1428,N_811);
or U3345 (N_3345,N_1517,N_1900);
or U3346 (N_3346,N_1886,N_116);
nand U3347 (N_3347,N_1215,N_1138);
and U3348 (N_3348,N_1672,N_182);
or U3349 (N_3349,N_1933,N_1878);
nand U3350 (N_3350,N_554,N_203);
or U3351 (N_3351,N_788,N_568);
and U3352 (N_3352,N_1362,N_897);
nand U3353 (N_3353,N_1775,N_1892);
and U3354 (N_3354,N_1925,N_1884);
nor U3355 (N_3355,N_1896,N_249);
nor U3356 (N_3356,N_476,N_1817);
or U3357 (N_3357,N_1983,N_166);
or U3358 (N_3358,N_819,N_1369);
nand U3359 (N_3359,N_1797,N_943);
or U3360 (N_3360,N_565,N_394);
or U3361 (N_3361,N_676,N_1895);
or U3362 (N_3362,N_355,N_512);
nand U3363 (N_3363,N_437,N_1527);
xnor U3364 (N_3364,N_33,N_623);
or U3365 (N_3365,N_1318,N_587);
nand U3366 (N_3366,N_543,N_47);
nand U3367 (N_3367,N_1972,N_1940);
xnor U3368 (N_3368,N_266,N_1157);
nor U3369 (N_3369,N_1632,N_155);
nor U3370 (N_3370,N_1229,N_1923);
nor U3371 (N_3371,N_1917,N_1913);
nor U3372 (N_3372,N_1958,N_952);
or U3373 (N_3373,N_996,N_786);
and U3374 (N_3374,N_261,N_333);
and U3375 (N_3375,N_1183,N_984);
or U3376 (N_3376,N_1888,N_1364);
and U3377 (N_3377,N_512,N_1534);
or U3378 (N_3378,N_892,N_590);
and U3379 (N_3379,N_405,N_217);
and U3380 (N_3380,N_27,N_675);
nor U3381 (N_3381,N_1125,N_1169);
or U3382 (N_3382,N_1377,N_1944);
nor U3383 (N_3383,N_390,N_844);
and U3384 (N_3384,N_1073,N_1704);
nand U3385 (N_3385,N_1925,N_534);
nor U3386 (N_3386,N_361,N_536);
nand U3387 (N_3387,N_1107,N_1281);
nand U3388 (N_3388,N_18,N_343);
or U3389 (N_3389,N_863,N_738);
or U3390 (N_3390,N_680,N_1614);
nand U3391 (N_3391,N_1462,N_938);
nor U3392 (N_3392,N_763,N_557);
nand U3393 (N_3393,N_1081,N_1454);
nand U3394 (N_3394,N_1798,N_1251);
and U3395 (N_3395,N_703,N_1347);
nand U3396 (N_3396,N_115,N_804);
nand U3397 (N_3397,N_1229,N_1661);
nand U3398 (N_3398,N_1914,N_505);
nor U3399 (N_3399,N_999,N_257);
or U3400 (N_3400,N_1936,N_1375);
and U3401 (N_3401,N_859,N_573);
nor U3402 (N_3402,N_936,N_261);
nand U3403 (N_3403,N_1557,N_690);
and U3404 (N_3404,N_366,N_1748);
and U3405 (N_3405,N_283,N_1695);
nor U3406 (N_3406,N_1693,N_967);
nand U3407 (N_3407,N_897,N_1441);
and U3408 (N_3408,N_1461,N_280);
xnor U3409 (N_3409,N_1230,N_1941);
nand U3410 (N_3410,N_158,N_1458);
nand U3411 (N_3411,N_243,N_17);
or U3412 (N_3412,N_528,N_1277);
or U3413 (N_3413,N_562,N_768);
nor U3414 (N_3414,N_424,N_1071);
nor U3415 (N_3415,N_580,N_1986);
nor U3416 (N_3416,N_1744,N_63);
nand U3417 (N_3417,N_1105,N_1708);
nor U3418 (N_3418,N_43,N_365);
nor U3419 (N_3419,N_1022,N_1550);
nand U3420 (N_3420,N_692,N_1935);
nand U3421 (N_3421,N_1657,N_579);
and U3422 (N_3422,N_1958,N_1700);
and U3423 (N_3423,N_1889,N_1835);
or U3424 (N_3424,N_658,N_494);
or U3425 (N_3425,N_295,N_1100);
nand U3426 (N_3426,N_250,N_509);
nand U3427 (N_3427,N_433,N_1360);
nand U3428 (N_3428,N_224,N_924);
nand U3429 (N_3429,N_956,N_851);
nand U3430 (N_3430,N_1880,N_1253);
or U3431 (N_3431,N_408,N_1548);
and U3432 (N_3432,N_1945,N_1741);
and U3433 (N_3433,N_384,N_496);
and U3434 (N_3434,N_1752,N_1181);
and U3435 (N_3435,N_874,N_1464);
or U3436 (N_3436,N_63,N_1251);
nand U3437 (N_3437,N_513,N_1780);
nand U3438 (N_3438,N_1209,N_453);
and U3439 (N_3439,N_541,N_1987);
nor U3440 (N_3440,N_474,N_489);
and U3441 (N_3441,N_1085,N_1478);
and U3442 (N_3442,N_1958,N_515);
or U3443 (N_3443,N_1919,N_1398);
and U3444 (N_3444,N_1443,N_812);
nand U3445 (N_3445,N_346,N_879);
nand U3446 (N_3446,N_548,N_774);
or U3447 (N_3447,N_1883,N_457);
or U3448 (N_3448,N_315,N_807);
and U3449 (N_3449,N_512,N_1286);
and U3450 (N_3450,N_1319,N_1888);
or U3451 (N_3451,N_261,N_1022);
nand U3452 (N_3452,N_785,N_1608);
or U3453 (N_3453,N_525,N_700);
xnor U3454 (N_3454,N_793,N_790);
xor U3455 (N_3455,N_616,N_1254);
and U3456 (N_3456,N_654,N_844);
and U3457 (N_3457,N_348,N_36);
and U3458 (N_3458,N_1862,N_1331);
and U3459 (N_3459,N_1726,N_1837);
nand U3460 (N_3460,N_1194,N_198);
nor U3461 (N_3461,N_1397,N_388);
and U3462 (N_3462,N_657,N_1618);
nor U3463 (N_3463,N_1955,N_247);
or U3464 (N_3464,N_678,N_533);
nor U3465 (N_3465,N_1632,N_1763);
or U3466 (N_3466,N_1915,N_1872);
nor U3467 (N_3467,N_1735,N_651);
nor U3468 (N_3468,N_1410,N_353);
and U3469 (N_3469,N_1987,N_1595);
and U3470 (N_3470,N_1351,N_607);
nor U3471 (N_3471,N_283,N_1121);
nor U3472 (N_3472,N_1986,N_1948);
nand U3473 (N_3473,N_339,N_1012);
nor U3474 (N_3474,N_703,N_1492);
and U3475 (N_3475,N_846,N_755);
nand U3476 (N_3476,N_1489,N_1075);
nand U3477 (N_3477,N_948,N_1070);
and U3478 (N_3478,N_809,N_1992);
and U3479 (N_3479,N_223,N_1804);
or U3480 (N_3480,N_776,N_1788);
nand U3481 (N_3481,N_490,N_1664);
nand U3482 (N_3482,N_930,N_1959);
nand U3483 (N_3483,N_1337,N_689);
nand U3484 (N_3484,N_266,N_867);
nor U3485 (N_3485,N_1370,N_661);
nand U3486 (N_3486,N_79,N_1032);
or U3487 (N_3487,N_1683,N_1816);
nor U3488 (N_3488,N_1994,N_553);
nor U3489 (N_3489,N_1949,N_1996);
and U3490 (N_3490,N_144,N_1738);
and U3491 (N_3491,N_429,N_813);
nand U3492 (N_3492,N_23,N_410);
nor U3493 (N_3493,N_828,N_1990);
nor U3494 (N_3494,N_925,N_372);
nor U3495 (N_3495,N_1949,N_1948);
nor U3496 (N_3496,N_1442,N_1863);
nor U3497 (N_3497,N_1929,N_1992);
nand U3498 (N_3498,N_175,N_165);
nand U3499 (N_3499,N_1613,N_1234);
nor U3500 (N_3500,N_867,N_1137);
nand U3501 (N_3501,N_1812,N_1782);
and U3502 (N_3502,N_145,N_1704);
and U3503 (N_3503,N_916,N_447);
or U3504 (N_3504,N_1675,N_52);
nor U3505 (N_3505,N_1534,N_162);
nor U3506 (N_3506,N_796,N_802);
or U3507 (N_3507,N_794,N_553);
or U3508 (N_3508,N_1218,N_1927);
or U3509 (N_3509,N_873,N_1316);
nand U3510 (N_3510,N_1402,N_1275);
xnor U3511 (N_3511,N_1879,N_411);
and U3512 (N_3512,N_1462,N_1997);
nand U3513 (N_3513,N_658,N_367);
nor U3514 (N_3514,N_1484,N_1234);
and U3515 (N_3515,N_156,N_1654);
nor U3516 (N_3516,N_1285,N_952);
or U3517 (N_3517,N_1315,N_783);
and U3518 (N_3518,N_1338,N_1469);
nor U3519 (N_3519,N_1088,N_1566);
or U3520 (N_3520,N_1618,N_402);
or U3521 (N_3521,N_648,N_5);
nor U3522 (N_3522,N_1758,N_1995);
nand U3523 (N_3523,N_1045,N_1574);
and U3524 (N_3524,N_1821,N_1363);
or U3525 (N_3525,N_507,N_282);
nor U3526 (N_3526,N_1824,N_1008);
nand U3527 (N_3527,N_673,N_757);
nor U3528 (N_3528,N_1873,N_1458);
and U3529 (N_3529,N_715,N_1760);
xnor U3530 (N_3530,N_537,N_84);
or U3531 (N_3531,N_571,N_1369);
nand U3532 (N_3532,N_180,N_323);
and U3533 (N_3533,N_1143,N_1082);
or U3534 (N_3534,N_275,N_801);
nand U3535 (N_3535,N_1020,N_1487);
and U3536 (N_3536,N_1043,N_354);
nor U3537 (N_3537,N_1227,N_455);
and U3538 (N_3538,N_1489,N_35);
xnor U3539 (N_3539,N_1928,N_1516);
nor U3540 (N_3540,N_1831,N_714);
nand U3541 (N_3541,N_214,N_567);
and U3542 (N_3542,N_312,N_570);
nor U3543 (N_3543,N_195,N_1046);
nor U3544 (N_3544,N_820,N_134);
and U3545 (N_3545,N_1772,N_1190);
and U3546 (N_3546,N_231,N_99);
and U3547 (N_3547,N_1932,N_1612);
nand U3548 (N_3548,N_1085,N_1542);
nor U3549 (N_3549,N_415,N_1057);
and U3550 (N_3550,N_1740,N_297);
or U3551 (N_3551,N_120,N_1194);
and U3552 (N_3552,N_1288,N_914);
and U3553 (N_3553,N_593,N_1469);
and U3554 (N_3554,N_1230,N_989);
nand U3555 (N_3555,N_354,N_1304);
nor U3556 (N_3556,N_1662,N_1887);
or U3557 (N_3557,N_1515,N_1622);
nand U3558 (N_3558,N_1700,N_105);
or U3559 (N_3559,N_610,N_734);
and U3560 (N_3560,N_809,N_973);
nand U3561 (N_3561,N_1789,N_252);
or U3562 (N_3562,N_1447,N_1148);
nor U3563 (N_3563,N_146,N_1706);
or U3564 (N_3564,N_1633,N_523);
nor U3565 (N_3565,N_1047,N_1948);
nand U3566 (N_3566,N_1791,N_1908);
or U3567 (N_3567,N_1385,N_461);
nor U3568 (N_3568,N_1021,N_219);
nor U3569 (N_3569,N_1845,N_1472);
and U3570 (N_3570,N_13,N_397);
nand U3571 (N_3571,N_786,N_619);
nor U3572 (N_3572,N_525,N_1968);
or U3573 (N_3573,N_1390,N_63);
and U3574 (N_3574,N_1540,N_1430);
nor U3575 (N_3575,N_487,N_1732);
or U3576 (N_3576,N_1154,N_1308);
nor U3577 (N_3577,N_666,N_1361);
nand U3578 (N_3578,N_1233,N_301);
nand U3579 (N_3579,N_963,N_1088);
nor U3580 (N_3580,N_247,N_1616);
nor U3581 (N_3581,N_831,N_1243);
nor U3582 (N_3582,N_1012,N_1881);
or U3583 (N_3583,N_1895,N_225);
nor U3584 (N_3584,N_1550,N_1371);
or U3585 (N_3585,N_1684,N_846);
nor U3586 (N_3586,N_1978,N_1813);
or U3587 (N_3587,N_1294,N_1224);
nor U3588 (N_3588,N_723,N_779);
nand U3589 (N_3589,N_1576,N_331);
nand U3590 (N_3590,N_774,N_593);
nand U3591 (N_3591,N_1718,N_266);
or U3592 (N_3592,N_151,N_1437);
nor U3593 (N_3593,N_748,N_1204);
xor U3594 (N_3594,N_653,N_775);
nor U3595 (N_3595,N_190,N_1578);
and U3596 (N_3596,N_1464,N_1636);
and U3597 (N_3597,N_1904,N_1649);
and U3598 (N_3598,N_1822,N_983);
nor U3599 (N_3599,N_449,N_832);
nor U3600 (N_3600,N_1098,N_1557);
nor U3601 (N_3601,N_1301,N_476);
or U3602 (N_3602,N_726,N_364);
or U3603 (N_3603,N_1956,N_767);
nor U3604 (N_3604,N_361,N_1002);
nand U3605 (N_3605,N_944,N_1453);
nor U3606 (N_3606,N_1614,N_1260);
nor U3607 (N_3607,N_445,N_893);
and U3608 (N_3608,N_749,N_459);
xor U3609 (N_3609,N_1759,N_1145);
and U3610 (N_3610,N_991,N_1862);
and U3611 (N_3611,N_153,N_1945);
nand U3612 (N_3612,N_714,N_368);
nor U3613 (N_3613,N_1483,N_856);
nor U3614 (N_3614,N_1312,N_1218);
and U3615 (N_3615,N_1847,N_1727);
or U3616 (N_3616,N_1000,N_1747);
xor U3617 (N_3617,N_257,N_1703);
and U3618 (N_3618,N_1470,N_1473);
or U3619 (N_3619,N_263,N_621);
nand U3620 (N_3620,N_109,N_802);
and U3621 (N_3621,N_1251,N_1621);
nand U3622 (N_3622,N_212,N_786);
nor U3623 (N_3623,N_1165,N_75);
and U3624 (N_3624,N_1520,N_285);
nor U3625 (N_3625,N_1878,N_245);
and U3626 (N_3626,N_1657,N_1568);
or U3627 (N_3627,N_1593,N_32);
nand U3628 (N_3628,N_1490,N_1126);
and U3629 (N_3629,N_1580,N_117);
nand U3630 (N_3630,N_241,N_1430);
nor U3631 (N_3631,N_1051,N_1614);
nand U3632 (N_3632,N_607,N_1114);
nand U3633 (N_3633,N_1188,N_1279);
and U3634 (N_3634,N_1375,N_1408);
nand U3635 (N_3635,N_1122,N_1740);
nand U3636 (N_3636,N_1505,N_726);
and U3637 (N_3637,N_441,N_31);
and U3638 (N_3638,N_118,N_1899);
nor U3639 (N_3639,N_441,N_277);
nand U3640 (N_3640,N_1258,N_114);
or U3641 (N_3641,N_93,N_153);
or U3642 (N_3642,N_848,N_1508);
and U3643 (N_3643,N_195,N_24);
nor U3644 (N_3644,N_1952,N_250);
nand U3645 (N_3645,N_1226,N_1266);
nand U3646 (N_3646,N_1840,N_1231);
or U3647 (N_3647,N_1201,N_526);
and U3648 (N_3648,N_1504,N_1750);
nor U3649 (N_3649,N_1293,N_1103);
and U3650 (N_3650,N_494,N_1722);
nand U3651 (N_3651,N_528,N_577);
or U3652 (N_3652,N_993,N_348);
and U3653 (N_3653,N_1504,N_1437);
or U3654 (N_3654,N_118,N_949);
or U3655 (N_3655,N_955,N_423);
or U3656 (N_3656,N_674,N_954);
and U3657 (N_3657,N_773,N_1494);
and U3658 (N_3658,N_244,N_1518);
nand U3659 (N_3659,N_1942,N_1607);
nand U3660 (N_3660,N_1392,N_725);
nand U3661 (N_3661,N_1757,N_899);
and U3662 (N_3662,N_1243,N_1652);
or U3663 (N_3663,N_1960,N_1942);
nor U3664 (N_3664,N_346,N_1178);
and U3665 (N_3665,N_631,N_1397);
nand U3666 (N_3666,N_669,N_382);
or U3667 (N_3667,N_521,N_699);
or U3668 (N_3668,N_1695,N_725);
or U3669 (N_3669,N_1621,N_714);
nand U3670 (N_3670,N_750,N_693);
or U3671 (N_3671,N_1599,N_903);
nand U3672 (N_3672,N_1463,N_1992);
nor U3673 (N_3673,N_1677,N_860);
or U3674 (N_3674,N_586,N_628);
nand U3675 (N_3675,N_1009,N_1417);
nand U3676 (N_3676,N_642,N_1599);
or U3677 (N_3677,N_1591,N_458);
or U3678 (N_3678,N_1162,N_1589);
or U3679 (N_3679,N_1136,N_725);
and U3680 (N_3680,N_1576,N_1561);
nand U3681 (N_3681,N_896,N_829);
nor U3682 (N_3682,N_546,N_711);
and U3683 (N_3683,N_1775,N_251);
nand U3684 (N_3684,N_46,N_298);
xnor U3685 (N_3685,N_1138,N_780);
nor U3686 (N_3686,N_1748,N_147);
or U3687 (N_3687,N_152,N_1944);
nor U3688 (N_3688,N_156,N_1378);
nand U3689 (N_3689,N_553,N_211);
nand U3690 (N_3690,N_30,N_1613);
and U3691 (N_3691,N_1148,N_1817);
and U3692 (N_3692,N_1216,N_607);
and U3693 (N_3693,N_1805,N_1311);
or U3694 (N_3694,N_1121,N_118);
nand U3695 (N_3695,N_426,N_1688);
or U3696 (N_3696,N_1395,N_326);
nand U3697 (N_3697,N_1491,N_790);
or U3698 (N_3698,N_254,N_1599);
and U3699 (N_3699,N_1273,N_1644);
nor U3700 (N_3700,N_1923,N_19);
and U3701 (N_3701,N_175,N_1654);
or U3702 (N_3702,N_1184,N_1410);
nor U3703 (N_3703,N_37,N_539);
nor U3704 (N_3704,N_169,N_1809);
nor U3705 (N_3705,N_336,N_532);
or U3706 (N_3706,N_282,N_1975);
or U3707 (N_3707,N_1040,N_1632);
and U3708 (N_3708,N_536,N_1579);
nand U3709 (N_3709,N_1657,N_1725);
or U3710 (N_3710,N_1817,N_1957);
nand U3711 (N_3711,N_342,N_1347);
or U3712 (N_3712,N_1497,N_246);
or U3713 (N_3713,N_1920,N_867);
and U3714 (N_3714,N_311,N_1947);
or U3715 (N_3715,N_681,N_72);
nand U3716 (N_3716,N_1172,N_1062);
or U3717 (N_3717,N_1913,N_764);
nand U3718 (N_3718,N_110,N_1390);
or U3719 (N_3719,N_856,N_97);
or U3720 (N_3720,N_579,N_616);
nand U3721 (N_3721,N_570,N_1570);
and U3722 (N_3722,N_813,N_1116);
nor U3723 (N_3723,N_1627,N_1717);
nand U3724 (N_3724,N_1159,N_1798);
nor U3725 (N_3725,N_153,N_1818);
or U3726 (N_3726,N_1632,N_1987);
nor U3727 (N_3727,N_547,N_447);
xor U3728 (N_3728,N_1991,N_1494);
nor U3729 (N_3729,N_1140,N_1302);
nor U3730 (N_3730,N_399,N_1258);
and U3731 (N_3731,N_1464,N_338);
or U3732 (N_3732,N_274,N_623);
nand U3733 (N_3733,N_1514,N_773);
or U3734 (N_3734,N_1227,N_917);
nand U3735 (N_3735,N_67,N_256);
or U3736 (N_3736,N_766,N_757);
nand U3737 (N_3737,N_710,N_854);
and U3738 (N_3738,N_471,N_1517);
nand U3739 (N_3739,N_1336,N_908);
nor U3740 (N_3740,N_246,N_1278);
and U3741 (N_3741,N_899,N_1729);
or U3742 (N_3742,N_1229,N_67);
nand U3743 (N_3743,N_743,N_28);
nor U3744 (N_3744,N_1005,N_1373);
or U3745 (N_3745,N_1031,N_1840);
nand U3746 (N_3746,N_82,N_1843);
or U3747 (N_3747,N_912,N_1239);
nand U3748 (N_3748,N_702,N_819);
nand U3749 (N_3749,N_1371,N_428);
nand U3750 (N_3750,N_99,N_1957);
nand U3751 (N_3751,N_185,N_853);
nor U3752 (N_3752,N_1482,N_1131);
nor U3753 (N_3753,N_1394,N_1761);
or U3754 (N_3754,N_606,N_735);
and U3755 (N_3755,N_342,N_205);
nor U3756 (N_3756,N_1979,N_717);
or U3757 (N_3757,N_599,N_1898);
or U3758 (N_3758,N_1636,N_735);
and U3759 (N_3759,N_678,N_1584);
and U3760 (N_3760,N_310,N_1016);
or U3761 (N_3761,N_1466,N_1461);
nor U3762 (N_3762,N_1383,N_690);
or U3763 (N_3763,N_1361,N_1717);
or U3764 (N_3764,N_887,N_1691);
or U3765 (N_3765,N_721,N_1421);
nor U3766 (N_3766,N_418,N_1134);
and U3767 (N_3767,N_1727,N_1319);
or U3768 (N_3768,N_473,N_470);
nor U3769 (N_3769,N_739,N_1643);
and U3770 (N_3770,N_1611,N_1025);
nor U3771 (N_3771,N_254,N_0);
and U3772 (N_3772,N_651,N_1039);
nor U3773 (N_3773,N_1529,N_478);
nand U3774 (N_3774,N_732,N_371);
or U3775 (N_3775,N_234,N_1915);
or U3776 (N_3776,N_1485,N_1111);
nor U3777 (N_3777,N_1441,N_1520);
nand U3778 (N_3778,N_1551,N_1614);
nor U3779 (N_3779,N_674,N_1592);
nor U3780 (N_3780,N_331,N_812);
nand U3781 (N_3781,N_1375,N_1389);
and U3782 (N_3782,N_576,N_1052);
or U3783 (N_3783,N_726,N_42);
nor U3784 (N_3784,N_994,N_1446);
nor U3785 (N_3785,N_429,N_156);
or U3786 (N_3786,N_603,N_1495);
nor U3787 (N_3787,N_536,N_1017);
and U3788 (N_3788,N_869,N_1129);
nand U3789 (N_3789,N_1695,N_359);
or U3790 (N_3790,N_210,N_1136);
nand U3791 (N_3791,N_335,N_1011);
nand U3792 (N_3792,N_61,N_374);
or U3793 (N_3793,N_253,N_296);
nor U3794 (N_3794,N_584,N_418);
nor U3795 (N_3795,N_1031,N_1438);
and U3796 (N_3796,N_1133,N_527);
and U3797 (N_3797,N_400,N_1452);
nor U3798 (N_3798,N_1183,N_1240);
nor U3799 (N_3799,N_460,N_1146);
nor U3800 (N_3800,N_1180,N_1691);
nand U3801 (N_3801,N_347,N_1744);
or U3802 (N_3802,N_300,N_1457);
nand U3803 (N_3803,N_903,N_272);
or U3804 (N_3804,N_994,N_1445);
or U3805 (N_3805,N_13,N_1262);
nor U3806 (N_3806,N_49,N_95);
or U3807 (N_3807,N_198,N_432);
nand U3808 (N_3808,N_1444,N_77);
and U3809 (N_3809,N_1276,N_1063);
and U3810 (N_3810,N_669,N_1844);
and U3811 (N_3811,N_1631,N_246);
xor U3812 (N_3812,N_331,N_1169);
nor U3813 (N_3813,N_688,N_727);
nand U3814 (N_3814,N_1630,N_588);
nor U3815 (N_3815,N_1330,N_569);
or U3816 (N_3816,N_904,N_1294);
and U3817 (N_3817,N_1197,N_1483);
nand U3818 (N_3818,N_845,N_58);
or U3819 (N_3819,N_1580,N_823);
nand U3820 (N_3820,N_1978,N_931);
nand U3821 (N_3821,N_1192,N_940);
nand U3822 (N_3822,N_988,N_1995);
nor U3823 (N_3823,N_224,N_848);
nor U3824 (N_3824,N_453,N_871);
and U3825 (N_3825,N_6,N_1595);
or U3826 (N_3826,N_423,N_970);
nand U3827 (N_3827,N_199,N_1924);
and U3828 (N_3828,N_1030,N_1698);
nor U3829 (N_3829,N_1772,N_1457);
and U3830 (N_3830,N_1743,N_732);
nand U3831 (N_3831,N_1433,N_1828);
nor U3832 (N_3832,N_1432,N_429);
and U3833 (N_3833,N_1366,N_1999);
nand U3834 (N_3834,N_114,N_1982);
nor U3835 (N_3835,N_1991,N_93);
and U3836 (N_3836,N_548,N_1475);
nand U3837 (N_3837,N_409,N_184);
or U3838 (N_3838,N_522,N_1615);
and U3839 (N_3839,N_1028,N_1468);
and U3840 (N_3840,N_1050,N_1515);
or U3841 (N_3841,N_498,N_1928);
and U3842 (N_3842,N_571,N_811);
nand U3843 (N_3843,N_1116,N_1799);
and U3844 (N_3844,N_1951,N_711);
nor U3845 (N_3845,N_1058,N_996);
and U3846 (N_3846,N_1855,N_801);
and U3847 (N_3847,N_37,N_1299);
and U3848 (N_3848,N_448,N_1476);
and U3849 (N_3849,N_1410,N_466);
nand U3850 (N_3850,N_880,N_1989);
nor U3851 (N_3851,N_1873,N_486);
or U3852 (N_3852,N_149,N_1845);
or U3853 (N_3853,N_1768,N_579);
nand U3854 (N_3854,N_520,N_93);
and U3855 (N_3855,N_877,N_1906);
nor U3856 (N_3856,N_844,N_1888);
or U3857 (N_3857,N_332,N_1325);
nand U3858 (N_3858,N_979,N_996);
nand U3859 (N_3859,N_109,N_16);
and U3860 (N_3860,N_600,N_1300);
nand U3861 (N_3861,N_565,N_1130);
nand U3862 (N_3862,N_1057,N_489);
nor U3863 (N_3863,N_267,N_1179);
nand U3864 (N_3864,N_964,N_389);
and U3865 (N_3865,N_316,N_839);
or U3866 (N_3866,N_995,N_482);
nand U3867 (N_3867,N_1539,N_827);
nor U3868 (N_3868,N_1486,N_1503);
and U3869 (N_3869,N_732,N_670);
nor U3870 (N_3870,N_288,N_370);
nor U3871 (N_3871,N_1844,N_713);
or U3872 (N_3872,N_263,N_1903);
nor U3873 (N_3873,N_1604,N_422);
nand U3874 (N_3874,N_1154,N_1809);
nor U3875 (N_3875,N_141,N_646);
or U3876 (N_3876,N_715,N_677);
and U3877 (N_3877,N_499,N_1018);
nand U3878 (N_3878,N_128,N_1141);
nand U3879 (N_3879,N_1477,N_524);
and U3880 (N_3880,N_198,N_735);
xnor U3881 (N_3881,N_1882,N_426);
and U3882 (N_3882,N_1346,N_301);
nand U3883 (N_3883,N_182,N_129);
or U3884 (N_3884,N_1972,N_1954);
nand U3885 (N_3885,N_1750,N_371);
and U3886 (N_3886,N_226,N_955);
nor U3887 (N_3887,N_1966,N_664);
nor U3888 (N_3888,N_983,N_876);
nand U3889 (N_3889,N_334,N_32);
nor U3890 (N_3890,N_275,N_777);
or U3891 (N_3891,N_1213,N_771);
nor U3892 (N_3892,N_307,N_228);
and U3893 (N_3893,N_1443,N_1273);
nor U3894 (N_3894,N_1248,N_1875);
or U3895 (N_3895,N_1834,N_1035);
nand U3896 (N_3896,N_1459,N_1833);
nand U3897 (N_3897,N_1508,N_201);
nand U3898 (N_3898,N_1587,N_1489);
or U3899 (N_3899,N_1359,N_1023);
nand U3900 (N_3900,N_915,N_1532);
and U3901 (N_3901,N_508,N_1924);
and U3902 (N_3902,N_1532,N_770);
or U3903 (N_3903,N_376,N_617);
and U3904 (N_3904,N_294,N_1847);
and U3905 (N_3905,N_930,N_1356);
nor U3906 (N_3906,N_747,N_288);
nor U3907 (N_3907,N_918,N_1605);
nor U3908 (N_3908,N_1516,N_660);
or U3909 (N_3909,N_1173,N_370);
nor U3910 (N_3910,N_937,N_1765);
nor U3911 (N_3911,N_902,N_1905);
nor U3912 (N_3912,N_939,N_1417);
or U3913 (N_3913,N_836,N_283);
nand U3914 (N_3914,N_811,N_472);
nand U3915 (N_3915,N_1739,N_137);
and U3916 (N_3916,N_1354,N_1936);
or U3917 (N_3917,N_1865,N_58);
nand U3918 (N_3918,N_1674,N_553);
or U3919 (N_3919,N_82,N_1988);
nand U3920 (N_3920,N_1203,N_181);
nor U3921 (N_3921,N_1167,N_882);
nor U3922 (N_3922,N_152,N_1265);
and U3923 (N_3923,N_1160,N_388);
nand U3924 (N_3924,N_454,N_291);
xor U3925 (N_3925,N_1886,N_467);
nor U3926 (N_3926,N_1928,N_1463);
or U3927 (N_3927,N_1180,N_37);
and U3928 (N_3928,N_1090,N_1396);
nor U3929 (N_3929,N_1550,N_768);
xnor U3930 (N_3930,N_1637,N_356);
and U3931 (N_3931,N_680,N_892);
nor U3932 (N_3932,N_1044,N_1733);
or U3933 (N_3933,N_377,N_1025);
nand U3934 (N_3934,N_1302,N_1845);
or U3935 (N_3935,N_620,N_1902);
and U3936 (N_3936,N_58,N_1393);
nand U3937 (N_3937,N_1724,N_1701);
and U3938 (N_3938,N_441,N_1126);
nand U3939 (N_3939,N_534,N_1739);
or U3940 (N_3940,N_1947,N_1466);
and U3941 (N_3941,N_379,N_228);
nor U3942 (N_3942,N_1080,N_999);
nor U3943 (N_3943,N_199,N_992);
nor U3944 (N_3944,N_242,N_1961);
or U3945 (N_3945,N_542,N_1664);
nand U3946 (N_3946,N_23,N_1299);
or U3947 (N_3947,N_1526,N_1959);
and U3948 (N_3948,N_1774,N_1295);
and U3949 (N_3949,N_822,N_1193);
nor U3950 (N_3950,N_183,N_1054);
nor U3951 (N_3951,N_378,N_317);
nand U3952 (N_3952,N_393,N_1751);
and U3953 (N_3953,N_1975,N_1870);
or U3954 (N_3954,N_455,N_981);
and U3955 (N_3955,N_1426,N_1360);
and U3956 (N_3956,N_1860,N_1276);
nor U3957 (N_3957,N_1333,N_1183);
or U3958 (N_3958,N_363,N_1156);
or U3959 (N_3959,N_1593,N_1588);
and U3960 (N_3960,N_1735,N_428);
and U3961 (N_3961,N_1689,N_810);
nor U3962 (N_3962,N_1325,N_1101);
nor U3963 (N_3963,N_1997,N_1233);
and U3964 (N_3964,N_1355,N_1591);
xor U3965 (N_3965,N_1985,N_1962);
nor U3966 (N_3966,N_1864,N_259);
nor U3967 (N_3967,N_1424,N_284);
nand U3968 (N_3968,N_410,N_1450);
xor U3969 (N_3969,N_876,N_1549);
nand U3970 (N_3970,N_1435,N_533);
nand U3971 (N_3971,N_1665,N_1598);
or U3972 (N_3972,N_1802,N_1373);
or U3973 (N_3973,N_1576,N_1211);
or U3974 (N_3974,N_1854,N_1902);
nor U3975 (N_3975,N_1078,N_442);
and U3976 (N_3976,N_549,N_12);
nand U3977 (N_3977,N_766,N_404);
or U3978 (N_3978,N_1449,N_1478);
nand U3979 (N_3979,N_1523,N_1693);
nand U3980 (N_3980,N_1371,N_1511);
nor U3981 (N_3981,N_1396,N_979);
nand U3982 (N_3982,N_1992,N_344);
nand U3983 (N_3983,N_526,N_1472);
and U3984 (N_3984,N_1233,N_434);
nor U3985 (N_3985,N_1634,N_1359);
nor U3986 (N_3986,N_1177,N_715);
nand U3987 (N_3987,N_1365,N_1949);
nand U3988 (N_3988,N_375,N_3);
nor U3989 (N_3989,N_1702,N_1567);
or U3990 (N_3990,N_472,N_1042);
nor U3991 (N_3991,N_370,N_600);
nand U3992 (N_3992,N_558,N_1609);
nor U3993 (N_3993,N_645,N_315);
and U3994 (N_3994,N_746,N_719);
and U3995 (N_3995,N_619,N_1821);
or U3996 (N_3996,N_1299,N_1466);
and U3997 (N_3997,N_1167,N_1665);
or U3998 (N_3998,N_732,N_1171);
nand U3999 (N_3999,N_764,N_1794);
and U4000 (N_4000,N_2419,N_2945);
or U4001 (N_4001,N_2999,N_3473);
and U4002 (N_4002,N_2857,N_3248);
and U4003 (N_4003,N_2613,N_3531);
and U4004 (N_4004,N_3826,N_3467);
nand U4005 (N_4005,N_3852,N_2767);
nand U4006 (N_4006,N_3650,N_2818);
nor U4007 (N_4007,N_3639,N_2038);
or U4008 (N_4008,N_3934,N_2731);
or U4009 (N_4009,N_2189,N_2651);
nand U4010 (N_4010,N_2155,N_3770);
nor U4011 (N_4011,N_3270,N_3478);
or U4012 (N_4012,N_2582,N_2796);
or U4013 (N_4013,N_2789,N_2183);
nand U4014 (N_4014,N_2678,N_2751);
nor U4015 (N_4015,N_2441,N_3711);
nand U4016 (N_4016,N_3456,N_2050);
or U4017 (N_4017,N_2361,N_3106);
nand U4018 (N_4018,N_3325,N_2943);
or U4019 (N_4019,N_2550,N_3028);
nand U4020 (N_4020,N_3805,N_3312);
and U4021 (N_4021,N_3888,N_3517);
nand U4022 (N_4022,N_2477,N_2688);
and U4023 (N_4023,N_3387,N_3245);
nor U4024 (N_4024,N_3524,N_3273);
nand U4025 (N_4025,N_3902,N_2983);
nor U4026 (N_4026,N_3876,N_3862);
nor U4027 (N_4027,N_2640,N_2641);
and U4028 (N_4028,N_3768,N_2209);
nor U4029 (N_4029,N_3115,N_2741);
nand U4030 (N_4030,N_2971,N_2330);
nor U4031 (N_4031,N_3544,N_2736);
or U4032 (N_4032,N_2236,N_3059);
and U4033 (N_4033,N_3729,N_2667);
nor U4034 (N_4034,N_2828,N_2383);
or U4035 (N_4035,N_2699,N_3803);
nor U4036 (N_4036,N_2542,N_3165);
and U4037 (N_4037,N_3297,N_2339);
and U4038 (N_4038,N_2884,N_3151);
or U4039 (N_4039,N_2822,N_3860);
and U4040 (N_4040,N_2481,N_3533);
and U4041 (N_4041,N_3501,N_3956);
and U4042 (N_4042,N_2043,N_2494);
nor U4043 (N_4043,N_2358,N_3882);
nand U4044 (N_4044,N_3961,N_3199);
or U4045 (N_4045,N_2355,N_3430);
nor U4046 (N_4046,N_3782,N_2394);
and U4047 (N_4047,N_2514,N_3017);
nand U4048 (N_4048,N_3205,N_3884);
nor U4049 (N_4049,N_2961,N_3013);
or U4050 (N_4050,N_2469,N_2933);
nor U4051 (N_4051,N_3575,N_2516);
and U4052 (N_4052,N_2829,N_2920);
and U4053 (N_4053,N_2401,N_2825);
or U4054 (N_4054,N_3943,N_3764);
nand U4055 (N_4055,N_3692,N_3640);
and U4056 (N_4056,N_3084,N_3583);
nor U4057 (N_4057,N_2471,N_3033);
or U4058 (N_4058,N_3474,N_2010);
and U4059 (N_4059,N_2041,N_3459);
and U4060 (N_4060,N_2763,N_2118);
xnor U4061 (N_4061,N_2785,N_2913);
and U4062 (N_4062,N_3322,N_2738);
nor U4063 (N_4063,N_3872,N_3847);
nand U4064 (N_4064,N_2562,N_2128);
or U4065 (N_4065,N_3584,N_2004);
and U4066 (N_4066,N_3655,N_3225);
and U4067 (N_4067,N_3874,N_3586);
and U4068 (N_4068,N_3182,N_3565);
or U4069 (N_4069,N_3713,N_2690);
nor U4070 (N_4070,N_3632,N_3579);
and U4071 (N_4071,N_2359,N_3893);
nor U4072 (N_4072,N_3966,N_3851);
and U4073 (N_4073,N_2325,N_2534);
and U4074 (N_4074,N_3564,N_3004);
nor U4075 (N_4075,N_3492,N_2179);
nand U4076 (N_4076,N_2243,N_2342);
and U4077 (N_4077,N_3078,N_2385);
and U4078 (N_4078,N_3491,N_3259);
or U4079 (N_4079,N_3070,N_3587);
nand U4080 (N_4080,N_2080,N_3923);
and U4081 (N_4081,N_3117,N_3614);
or U4082 (N_4082,N_3175,N_3236);
nand U4083 (N_4083,N_3742,N_3975);
nand U4084 (N_4084,N_2484,N_2865);
and U4085 (N_4085,N_2107,N_3056);
nor U4086 (N_4086,N_3897,N_2980);
or U4087 (N_4087,N_3170,N_2122);
or U4088 (N_4088,N_2743,N_3889);
nor U4089 (N_4089,N_2096,N_2705);
or U4090 (N_4090,N_2332,N_2695);
or U4091 (N_4091,N_3947,N_3853);
nor U4092 (N_4092,N_2021,N_3686);
or U4093 (N_4093,N_3690,N_3986);
nand U4094 (N_4094,N_3087,N_2490);
nand U4095 (N_4095,N_2259,N_2430);
nor U4096 (N_4096,N_3712,N_2996);
and U4097 (N_4097,N_3415,N_3815);
nor U4098 (N_4098,N_2252,N_3667);
and U4099 (N_4099,N_2614,N_2827);
nand U4100 (N_4100,N_3073,N_2292);
and U4101 (N_4101,N_3453,N_3879);
nand U4102 (N_4102,N_2347,N_2926);
nand U4103 (N_4103,N_2574,N_3468);
nand U4104 (N_4104,N_3145,N_2526);
nor U4105 (N_4105,N_3880,N_2852);
or U4106 (N_4106,N_2815,N_2120);
or U4107 (N_4107,N_2257,N_3323);
nand U4108 (N_4108,N_2165,N_3562);
and U4109 (N_4109,N_3052,N_3445);
or U4110 (N_4110,N_2079,N_3103);
or U4111 (N_4111,N_3654,N_3792);
nand U4112 (N_4112,N_3948,N_3649);
nand U4113 (N_4113,N_3168,N_2282);
or U4114 (N_4114,N_3385,N_3334);
nor U4115 (N_4115,N_2657,N_2584);
or U4116 (N_4116,N_3623,N_3597);
or U4117 (N_4117,N_2217,N_2171);
or U4118 (N_4118,N_2501,N_2173);
and U4119 (N_4119,N_2020,N_3974);
or U4120 (N_4120,N_3911,N_3596);
and U4121 (N_4121,N_3790,N_2253);
and U4122 (N_4122,N_3025,N_2664);
nand U4123 (N_4123,N_3133,N_3946);
and U4124 (N_4124,N_2957,N_2451);
and U4125 (N_4125,N_2934,N_2150);
and U4126 (N_4126,N_2024,N_3003);
nor U4127 (N_4127,N_3723,N_3341);
nand U4128 (N_4128,N_3027,N_3613);
nor U4129 (N_4129,N_2305,N_2098);
or U4130 (N_4130,N_2679,N_2851);
and U4131 (N_4131,N_3337,N_2406);
nor U4132 (N_4132,N_2517,N_2721);
nor U4133 (N_4133,N_2775,N_3828);
and U4134 (N_4134,N_2476,N_2571);
nor U4135 (N_4135,N_2119,N_3443);
nor U4136 (N_4136,N_2124,N_2007);
nand U4137 (N_4137,N_2046,N_2917);
or U4138 (N_4138,N_2753,N_3725);
or U4139 (N_4139,N_3209,N_2662);
or U4140 (N_4140,N_2057,N_3189);
nor U4141 (N_4141,N_3231,N_2085);
nor U4142 (N_4142,N_3605,N_2212);
nand U4143 (N_4143,N_3539,N_3120);
or U4144 (N_4144,N_2612,N_2223);
nor U4145 (N_4145,N_2340,N_3012);
or U4146 (N_4146,N_3938,N_3959);
nand U4147 (N_4147,N_2137,N_3124);
nand U4148 (N_4148,N_3881,N_2138);
nand U4149 (N_4149,N_2877,N_2569);
nand U4150 (N_4150,N_3286,N_2161);
nand U4151 (N_4151,N_3043,N_3775);
or U4152 (N_4152,N_3202,N_2938);
nand U4153 (N_4153,N_2345,N_2166);
nor U4154 (N_4154,N_2962,N_2949);
and U4155 (N_4155,N_2802,N_3557);
nor U4156 (N_4156,N_3651,N_3169);
nand U4157 (N_4157,N_3740,N_2411);
nor U4158 (N_4158,N_2047,N_2814);
and U4159 (N_4159,N_3353,N_3919);
or U4160 (N_4160,N_3525,N_3053);
or U4161 (N_4161,N_3212,N_3736);
nand U4162 (N_4162,N_3714,N_3419);
xnor U4163 (N_4163,N_2812,N_2849);
nand U4164 (N_4164,N_3294,N_3185);
nand U4165 (N_4165,N_2027,N_2054);
or U4166 (N_4166,N_2101,N_2693);
and U4167 (N_4167,N_3598,N_3984);
nor U4168 (N_4168,N_3247,N_3755);
nor U4169 (N_4169,N_3767,N_2283);
nor U4170 (N_4170,N_2296,N_2072);
nand U4171 (N_4171,N_3235,N_2400);
nand U4172 (N_4172,N_3561,N_2391);
nor U4173 (N_4173,N_3018,N_2931);
nor U4174 (N_4174,N_3771,N_2579);
or U4175 (N_4175,N_2228,N_2914);
or U4176 (N_4176,N_3239,N_2220);
nand U4177 (N_4177,N_3549,N_3754);
and U4178 (N_4178,N_2899,N_2384);
and U4179 (N_4179,N_2982,N_3995);
nor U4180 (N_4180,N_3519,N_3455);
nand U4181 (N_4181,N_3305,N_3858);
or U4182 (N_4182,N_2109,N_3252);
or U4183 (N_4183,N_3748,N_3645);
nand U4184 (N_4184,N_2858,N_2280);
and U4185 (N_4185,N_3854,N_3421);
nor U4186 (N_4186,N_2370,N_2218);
or U4187 (N_4187,N_3931,N_3431);
or U4188 (N_4188,N_2639,N_3843);
nor U4189 (N_4189,N_3657,N_3300);
nor U4190 (N_4190,N_3410,N_3681);
nand U4191 (N_4191,N_3724,N_3555);
and U4192 (N_4192,N_3972,N_2442);
or U4193 (N_4193,N_3777,N_2556);
nand U4194 (N_4194,N_3976,N_3733);
or U4195 (N_4195,N_3011,N_3745);
and U4196 (N_4196,N_3497,N_3634);
nor U4197 (N_4197,N_3253,N_2337);
nand U4198 (N_4198,N_3275,N_2434);
or U4199 (N_4199,N_2671,N_3905);
or U4200 (N_4200,N_3469,N_2134);
or U4201 (N_4201,N_2308,N_2285);
and U4202 (N_4202,N_2397,N_3261);
and U4203 (N_4203,N_2486,N_2258);
or U4204 (N_4204,N_2774,N_2300);
and U4205 (N_4205,N_2364,N_3585);
nor U4206 (N_4206,N_3857,N_3730);
nand U4207 (N_4207,N_3656,N_3024);
xnor U4208 (N_4208,N_2276,N_2927);
nand U4209 (N_4209,N_3167,N_2642);
and U4210 (N_4210,N_3232,N_3908);
nor U4211 (N_4211,N_2061,N_3265);
nand U4212 (N_4212,N_3765,N_2859);
nor U4213 (N_4213,N_2843,N_3753);
or U4214 (N_4214,N_2089,N_2866);
and U4215 (N_4215,N_3841,N_2868);
or U4216 (N_4216,N_3763,N_3154);
nand U4217 (N_4217,N_3950,N_2127);
nand U4218 (N_4218,N_2942,N_3664);
and U4219 (N_4219,N_3532,N_2413);
or U4220 (N_4220,N_2352,N_2807);
or U4221 (N_4221,N_3296,N_2928);
and U4222 (N_4222,N_3999,N_2316);
nor U4223 (N_4223,N_2696,N_3118);
nand U4224 (N_4224,N_3307,N_3174);
nor U4225 (N_4225,N_3920,N_3652);
and U4226 (N_4226,N_2402,N_3008);
and U4227 (N_4227,N_3551,N_3941);
nor U4228 (N_4228,N_3869,N_3490);
or U4229 (N_4229,N_2555,N_3509);
or U4230 (N_4230,N_3479,N_2718);
nor U4231 (N_4231,N_3391,N_2620);
xnor U4232 (N_4232,N_2299,N_2398);
nand U4233 (N_4233,N_2950,N_3394);
nand U4234 (N_4234,N_3816,N_3176);
nor U4235 (N_4235,N_3140,N_3503);
nor U4236 (N_4236,N_2488,N_3371);
nand U4237 (N_4237,N_3684,N_3206);
or U4238 (N_4238,N_2460,N_2691);
and U4239 (N_4239,N_2269,N_2029);
nor U4240 (N_4240,N_2604,N_3338);
and U4241 (N_4241,N_3475,N_3592);
nand U4242 (N_4242,N_3488,N_3835);
nor U4243 (N_4243,N_2543,N_2200);
and U4244 (N_4244,N_2395,N_3599);
nor U4245 (N_4245,N_2680,N_2005);
or U4246 (N_4246,N_2947,N_2674);
and U4247 (N_4247,N_2649,N_3345);
or U4248 (N_4248,N_3116,N_3347);
nand U4249 (N_4249,N_2341,N_3727);
and U4250 (N_4250,N_3703,N_3216);
nor U4251 (N_4251,N_2525,N_3061);
nand U4252 (N_4252,N_2372,N_2745);
or U4253 (N_4253,N_3360,N_3303);
nand U4254 (N_4254,N_3412,N_3126);
or U4255 (N_4255,N_3991,N_2362);
nor U4256 (N_4256,N_2954,N_3958);
and U4257 (N_4257,N_3643,N_3207);
or U4258 (N_4258,N_2765,N_2675);
or U4259 (N_4259,N_2133,N_2512);
and U4260 (N_4260,N_3507,N_2870);
nand U4261 (N_4261,N_3721,N_3311);
xor U4262 (N_4262,N_3791,N_3179);
nor U4263 (N_4263,N_2764,N_2194);
and U4264 (N_4264,N_2353,N_3595);
nand U4265 (N_4265,N_3160,N_2433);
or U4266 (N_4266,N_3363,N_2723);
nand U4267 (N_4267,N_3466,N_2226);
or U4268 (N_4268,N_3554,N_2506);
or U4269 (N_4269,N_2030,N_3899);
and U4270 (N_4270,N_2686,N_3158);
nand U4271 (N_4271,N_2909,N_2169);
nand U4272 (N_4272,N_2539,N_2523);
and U4273 (N_4273,N_3228,N_2412);
xnor U4274 (N_4274,N_2702,N_3617);
nor U4275 (N_4275,N_3821,N_2777);
and U4276 (N_4276,N_2130,N_3498);
nand U4277 (N_4277,N_3437,N_3255);
nand U4278 (N_4278,N_3540,N_3611);
nand U4279 (N_4279,N_2066,N_3336);
and U4280 (N_4280,N_3688,N_2214);
nand U4281 (N_4281,N_3258,N_2875);
or U4282 (N_4282,N_3400,N_3372);
nand U4283 (N_4283,N_3653,N_2132);
nand U4284 (N_4284,N_3054,N_2633);
and U4285 (N_4285,N_3386,N_2676);
nor U4286 (N_4286,N_2483,N_2952);
xor U4287 (N_4287,N_2912,N_2034);
and U4288 (N_4288,N_3057,N_3393);
or U4289 (N_4289,N_3982,N_2895);
or U4290 (N_4290,N_2896,N_3600);
nor U4291 (N_4291,N_3355,N_2991);
xnor U4292 (N_4292,N_2554,N_3382);
nand U4293 (N_4293,N_2951,N_2988);
or U4294 (N_4294,N_2421,N_2575);
and U4295 (N_4295,N_2164,N_2627);
nand U4296 (N_4296,N_3229,N_3785);
nor U4297 (N_4297,N_2320,N_3834);
or U4298 (N_4298,N_2146,N_2975);
or U4299 (N_4299,N_3081,N_3499);
and U4300 (N_4300,N_3060,N_3354);
nand U4301 (N_4301,N_3788,N_3728);
and U4302 (N_4302,N_3058,N_3493);
nor U4303 (N_4303,N_3864,N_2423);
nand U4304 (N_4304,N_2873,N_2845);
nand U4305 (N_4305,N_3241,N_2968);
nor U4306 (N_4306,N_2624,N_3074);
or U4307 (N_4307,N_3448,N_2443);
nand U4308 (N_4308,N_3100,N_2199);
nand U4309 (N_4309,N_3369,N_3090);
nand U4310 (N_4310,N_2022,N_3648);
nand U4311 (N_4311,N_2496,N_2193);
nand U4312 (N_4312,N_3641,N_2136);
and U4313 (N_4313,N_3996,N_3750);
and U4314 (N_4314,N_3020,N_2668);
xor U4315 (N_4315,N_3002,N_3271);
nand U4316 (N_4316,N_3240,N_2198);
and U4317 (N_4317,N_3547,N_3662);
nand U4318 (N_4318,N_3997,N_2778);
nand U4319 (N_4319,N_3045,N_3146);
and U4320 (N_4320,N_3756,N_3527);
or U4321 (N_4321,N_2800,N_2681);
nor U4322 (N_4322,N_2515,N_2069);
nand U4323 (N_4323,N_3510,N_2908);
or U4324 (N_4324,N_2206,N_2302);
nor U4325 (N_4325,N_2608,N_2768);
and U4326 (N_4326,N_3395,N_2771);
or U4327 (N_4327,N_2256,N_2861);
nor U4328 (N_4328,N_3365,N_3514);
nand U4329 (N_4329,N_2151,N_3898);
or U4330 (N_4330,N_2502,N_3687);
and U4331 (N_4331,N_3178,N_2769);
or U4332 (N_4332,N_3238,N_2810);
or U4333 (N_4333,N_3779,N_2918);
and U4334 (N_4334,N_2560,N_3041);
or U4335 (N_4335,N_2026,N_2883);
or U4336 (N_4336,N_2694,N_3942);
or U4337 (N_4337,N_2240,N_2637);
or U4338 (N_4338,N_3715,N_3401);
nand U4339 (N_4339,N_3695,N_2708);
nor U4340 (N_4340,N_3113,N_3769);
or U4341 (N_4341,N_3197,N_2363);
or U4342 (N_4342,N_3726,N_2598);
nor U4343 (N_4343,N_3486,N_3739);
nor U4344 (N_4344,N_2487,N_3685);
and U4345 (N_4345,N_2375,N_3374);
nand U4346 (N_4346,N_3761,N_3553);
and U4347 (N_4347,N_2946,N_3870);
nor U4348 (N_4348,N_3424,N_3744);
and U4349 (N_4349,N_3282,N_2500);
and U4350 (N_4350,N_3161,N_2255);
and U4351 (N_4351,N_2507,N_3604);
or U4352 (N_4352,N_2333,N_3556);
and U4353 (N_4353,N_2905,N_3977);
nand U4354 (N_4354,N_2530,N_2653);
or U4355 (N_4355,N_2035,N_2463);
and U4356 (N_4356,N_2188,N_2561);
or U4357 (N_4357,N_3180,N_3254);
nand U4358 (N_4358,N_2660,N_3505);
nand U4359 (N_4359,N_2087,N_2491);
nor U4360 (N_4360,N_2354,N_3917);
or U4361 (N_4361,N_3625,N_2297);
nor U4362 (N_4362,N_3675,N_2730);
nor U4363 (N_4363,N_2794,N_2279);
and U4364 (N_4364,N_3464,N_2060);
or U4365 (N_4365,N_3506,N_3978);
nor U4366 (N_4366,N_3181,N_2251);
nand U4367 (N_4367,N_3831,N_2075);
nor U4368 (N_4368,N_3629,N_2091);
and U4369 (N_4369,N_2838,N_3211);
or U4370 (N_4370,N_2545,N_3198);
or U4371 (N_4371,N_2840,N_3998);
and U4372 (N_4372,N_2470,N_3062);
or U4373 (N_4373,N_3227,N_2365);
or U4374 (N_4374,N_3993,N_2230);
nor U4375 (N_4375,N_2626,N_3030);
and U4376 (N_4376,N_3313,N_3083);
nand U4377 (N_4377,N_3447,N_3287);
nor U4378 (N_4378,N_2016,N_2823);
nor U4379 (N_4379,N_2860,N_2650);
nor U4380 (N_4380,N_2468,N_2659);
nor U4381 (N_4381,N_3940,N_2714);
or U4382 (N_4382,N_3331,N_2710);
and U4383 (N_4383,N_3795,N_3992);
nand U4384 (N_4384,N_2622,N_2735);
nand U4385 (N_4385,N_3064,N_3191);
and U4386 (N_4386,N_2467,N_3251);
and U4387 (N_4387,N_3086,N_2634);
or U4388 (N_4388,N_2281,N_2303);
nor U4389 (N_4389,N_2605,N_3536);
and U4390 (N_4390,N_3077,N_3717);
nor U4391 (N_4391,N_2254,N_3523);
and U4392 (N_4392,N_3789,N_2816);
or U4393 (N_4393,N_3289,N_3148);
nand U4394 (N_4394,N_2290,N_2770);
nor U4395 (N_4395,N_2479,N_3042);
nand U4396 (N_4396,N_2009,N_3516);
nand U4397 (N_4397,N_3809,N_2454);
nand U4398 (N_4398,N_3183,N_3280);
or U4399 (N_4399,N_2655,N_3637);
and U4400 (N_4400,N_2930,N_2819);
nand U4401 (N_4401,N_3633,N_2242);
and U4402 (N_4402,N_3927,N_3856);
or U4403 (N_4403,N_3576,N_2772);
nand U4404 (N_4404,N_2963,N_3438);
nor U4405 (N_4405,N_2033,N_3379);
nor U4406 (N_4406,N_2513,N_3051);
or U4407 (N_4407,N_2453,N_3746);
nand U4408 (N_4408,N_3827,N_2040);
nor U4409 (N_4409,N_2168,N_3694);
nand U4410 (N_4410,N_2184,N_2204);
and U4411 (N_4411,N_3339,N_2638);
nor U4412 (N_4412,N_2915,N_2094);
or U4413 (N_4413,N_3719,N_2288);
nand U4414 (N_4414,N_3925,N_2139);
or U4415 (N_4415,N_3463,N_2628);
nand U4416 (N_4416,N_3912,N_3578);
or U4417 (N_4417,N_2203,N_3906);
nor U4418 (N_4418,N_2489,N_2874);
nand U4419 (N_4419,N_3811,N_3731);
nor U4420 (N_4420,N_3244,N_2420);
nand U4421 (N_4421,N_2186,N_2504);
and U4422 (N_4422,N_3990,N_3234);
xor U4423 (N_4423,N_2399,N_2601);
nand U4424 (N_4424,N_2011,N_2611);
xnor U4425 (N_4425,N_3166,N_3718);
nand U4426 (N_4426,N_2238,N_3502);
or U4427 (N_4427,N_3967,N_3328);
nand U4428 (N_4428,N_2386,N_3836);
or U4429 (N_4429,N_3356,N_3094);
xnor U4430 (N_4430,N_2939,N_2196);
nor U4431 (N_4431,N_2371,N_3132);
nand U4432 (N_4432,N_2824,N_2881);
and U4433 (N_4433,N_2959,N_3817);
nand U4434 (N_4434,N_3377,N_2820);
and U4435 (N_4435,N_2058,N_2799);
nand U4436 (N_4436,N_2095,N_2744);
nor U4437 (N_4437,N_3200,N_2585);
nand U4438 (N_4438,N_2418,N_2264);
nor U4439 (N_4439,N_3440,N_3306);
nand U4440 (N_4440,N_2916,N_2644);
or U4441 (N_4441,N_2114,N_2855);
and U4442 (N_4442,N_2842,N_2336);
and U4443 (N_4443,N_2701,N_3450);
xor U4444 (N_4444,N_3432,N_2955);
and U4445 (N_4445,N_2672,N_3699);
or U4446 (N_4446,N_3658,N_2956);
nor U4447 (N_4447,N_3034,N_3281);
nand U4448 (N_4448,N_3630,N_3333);
and U4449 (N_4449,N_2856,N_3659);
or U4450 (N_4450,N_2459,N_3163);
or U4451 (N_4451,N_3968,N_3392);
nor U4452 (N_4452,N_3952,N_2278);
nor U4453 (N_4453,N_2833,N_3171);
and U4454 (N_4454,N_3276,N_2306);
and U4455 (N_4455,N_3204,N_3546);
and U4456 (N_4456,N_3482,N_2110);
or U4457 (N_4457,N_2967,N_2703);
nand U4458 (N_4458,N_3226,N_2910);
nand U4459 (N_4459,N_2301,N_3308);
nand U4460 (N_4460,N_2783,N_3773);
or U4461 (N_4461,N_3707,N_2792);
nand U4462 (N_4462,N_3568,N_2053);
nand U4463 (N_4463,N_2289,N_2937);
and U4464 (N_4464,N_3314,N_2329);
nand U4465 (N_4465,N_2602,N_2607);
and U4466 (N_4466,N_2103,N_3644);
nand U4467 (N_4467,N_2586,N_2093);
or U4468 (N_4468,N_3760,N_2304);
and U4469 (N_4469,N_2392,N_3384);
nand U4470 (N_4470,N_3112,N_2935);
xor U4471 (N_4471,N_3367,N_2902);
nor U4472 (N_4472,N_3177,N_3679);
nor U4473 (N_4473,N_2176,N_3786);
xor U4474 (N_4474,N_2588,N_2958);
or U4475 (N_4475,N_3065,N_3677);
nor U4476 (N_4476,N_2563,N_3939);
nor U4477 (N_4477,N_3678,N_3570);
or U4478 (N_4478,N_2998,N_2064);
and U4479 (N_4479,N_3890,N_2781);
and U4480 (N_4480,N_2415,N_2482);
and U4481 (N_4481,N_3357,N_2984);
and U4482 (N_4482,N_3573,N_3368);
nor U4483 (N_4483,N_2153,N_2779);
nand U4484 (N_4484,N_2813,N_3137);
nor U4485 (N_4485,N_2493,N_3264);
nand U4486 (N_4486,N_2112,N_2941);
or U4487 (N_4487,N_3928,N_2629);
or U4488 (N_4488,N_3190,N_3285);
nor U4489 (N_4489,N_3196,N_3672);
and U4490 (N_4490,N_2263,N_3612);
or U4491 (N_4491,N_3622,N_2177);
nor U4492 (N_4492,N_2158,N_2717);
nand U4493 (N_4493,N_3388,N_3309);
or U4494 (N_4494,N_2396,N_2245);
or U4495 (N_4495,N_2044,N_2900);
nand U4496 (N_4496,N_3518,N_2893);
and U4497 (N_4497,N_2427,N_3411);
and U4498 (N_4498,N_2791,N_3621);
nand U4499 (N_4499,N_2190,N_3500);
nor U4500 (N_4500,N_2167,N_3219);
or U4501 (N_4501,N_2437,N_2898);
or U4502 (N_4502,N_3830,N_3208);
nor U4503 (N_4503,N_3218,N_2536);
nor U4504 (N_4504,N_3751,N_3955);
or U4505 (N_4505,N_3416,N_3543);
or U4506 (N_4506,N_2734,N_3125);
nand U4507 (N_4507,N_2076,N_2826);
and U4508 (N_4508,N_2172,N_3315);
and U4509 (N_4509,N_2558,N_2994);
nand U4510 (N_4510,N_2760,N_3960);
and U4511 (N_4511,N_2405,N_2393);
xor U4512 (N_4512,N_2338,N_2887);
nand U4513 (N_4513,N_2234,N_3566);
nand U4514 (N_4514,N_3104,N_3980);
nand U4515 (N_4515,N_2367,N_2636);
and U4516 (N_4516,N_2716,N_3038);
xnor U4517 (N_4517,N_3068,N_2284);
nand U4518 (N_4518,N_3048,N_3710);
or U4519 (N_4519,N_3855,N_2548);
or U4520 (N_4520,N_3953,N_3217);
or U4521 (N_4521,N_3326,N_3800);
and U4522 (N_4522,N_2082,N_2499);
or U4523 (N_4523,N_3274,N_3138);
and U4524 (N_4524,N_3577,N_2727);
and U4525 (N_4525,N_2195,N_2596);
and U4526 (N_4526,N_2403,N_2923);
nand U4527 (N_4527,N_3290,N_2692);
nand U4528 (N_4528,N_2871,N_2964);
and U4529 (N_4529,N_3962,N_2108);
or U4530 (N_4530,N_2268,N_2140);
and U4531 (N_4531,N_3230,N_3963);
nand U4532 (N_4532,N_3627,N_2707);
nor U4533 (N_4533,N_2665,N_2201);
and U4534 (N_4534,N_3134,N_2077);
nor U4535 (N_4535,N_3607,N_3029);
or U4536 (N_4536,N_3291,N_3000);
nor U4537 (N_4537,N_2619,N_2830);
nor U4538 (N_4538,N_3263,N_2520);
nand U4539 (N_4539,N_3272,N_2677);
and U4540 (N_4540,N_3031,N_2131);
or U4541 (N_4541,N_2457,N_2888);
nand U4542 (N_4542,N_3246,N_3616);
nor U4543 (N_4543,N_2211,N_3709);
or U4544 (N_4544,N_2531,N_3863);
or U4545 (N_4545,N_2728,N_2175);
or U4546 (N_4546,N_3776,N_3620);
and U4547 (N_4547,N_3581,N_2532);
nor U4548 (N_4548,N_3608,N_3590);
nand U4549 (N_4549,N_3487,N_3414);
and U4550 (N_4550,N_3119,N_3172);
or U4551 (N_4551,N_3129,N_2348);
or U4552 (N_4552,N_3787,N_2697);
or U4553 (N_4553,N_3838,N_2786);
or U4554 (N_4554,N_3082,N_2906);
and U4555 (N_4555,N_2932,N_3873);
or U4556 (N_4556,N_2187,N_2466);
nand U4557 (N_4557,N_2689,N_3602);
or U4558 (N_4558,N_3757,N_2250);
or U4559 (N_4559,N_3351,N_2055);
xor U4560 (N_4560,N_2422,N_3403);
nand U4561 (N_4561,N_2510,N_3930);
nor U4562 (N_4562,N_2152,N_3647);
or U4563 (N_4563,N_2700,N_3066);
nor U4564 (N_4564,N_3582,N_3215);
nor U4565 (N_4565,N_3846,N_2287);
nor U4566 (N_4566,N_3628,N_2729);
or U4567 (N_4567,N_3895,N_2552);
and U4568 (N_4568,N_2989,N_2115);
and U4569 (N_4569,N_2524,N_2417);
nor U4570 (N_4570,N_2431,N_3075);
or U4571 (N_4571,N_3494,N_2557);
or U4572 (N_4572,N_3361,N_2919);
or U4573 (N_4573,N_3833,N_2215);
nor U4574 (N_4574,N_2310,N_2724);
nand U4575 (N_4575,N_2378,N_2326);
or U4576 (N_4576,N_3798,N_3909);
or U4577 (N_4577,N_2428,N_3804);
nand U4578 (N_4578,N_2948,N_3784);
nand U4579 (N_4579,N_2709,N_3472);
nor U4580 (N_4580,N_2309,N_2733);
nor U4581 (N_4581,N_2540,N_3954);
nand U4582 (N_4582,N_3673,N_3530);
nor U4583 (N_4583,N_2537,N_3601);
nand U4584 (N_4584,N_3702,N_3691);
nor U4585 (N_4585,N_3965,N_3091);
nor U4586 (N_4586,N_3439,N_3390);
and U4587 (N_4587,N_2811,N_3096);
nand U4588 (N_4588,N_2062,N_3563);
nor U4589 (N_4589,N_2973,N_3558);
nor U4590 (N_4590,N_2388,N_3548);
nor U4591 (N_4591,N_3348,N_3859);
and U4592 (N_4592,N_3781,N_3588);
and U4593 (N_4593,N_3164,N_3875);
nor U4594 (N_4594,N_3295,N_3734);
or U4595 (N_4595,N_3515,N_2074);
nor U4596 (N_4596,N_2713,N_2631);
nor U4597 (N_4597,N_3680,N_3362);
nor U4598 (N_4598,N_2635,N_3465);
and U4599 (N_4599,N_2970,N_3039);
or U4600 (N_4600,N_2685,N_2752);
and U4601 (N_4601,N_2522,N_2835);
or U4602 (N_4602,N_2117,N_2566);
or U4603 (N_4603,N_3141,N_2670);
or U4604 (N_4604,N_3454,N_3572);
and U4605 (N_4605,N_2408,N_3969);
nor U4606 (N_4606,N_3047,N_3458);
xor U4607 (N_4607,N_2995,N_3320);
nor U4608 (N_4608,N_3079,N_2897);
nor U4609 (N_4609,N_3910,N_3542);
and U4610 (N_4610,N_2615,N_3088);
or U4611 (N_4611,N_3135,N_3700);
and U4612 (N_4612,N_3267,N_3389);
nor U4613 (N_4613,N_3157,N_3526);
or U4614 (N_4614,N_3661,N_2573);
or U4615 (N_4615,N_3793,N_2616);
nor U4616 (N_4616,N_2273,N_3292);
nand U4617 (N_4617,N_3014,N_2298);
nand U4618 (N_4618,N_3642,N_3072);
nand U4619 (N_4619,N_3022,N_3105);
or U4620 (N_4620,N_2286,N_3201);
nor U4621 (N_4621,N_2045,N_2780);
and U4622 (N_4622,N_3344,N_3646);
nand U4623 (N_4623,N_3460,N_3844);
and U4624 (N_4624,N_3044,N_2452);
nand U4625 (N_4625,N_3335,N_2725);
or U4626 (N_4626,N_2368,N_3122);
nor U4627 (N_4627,N_3050,N_2202);
nand U4628 (N_4628,N_3298,N_3720);
or U4629 (N_4629,N_3871,N_3810);
and U4630 (N_4630,N_3749,N_2180);
or U4631 (N_4631,N_3921,N_3127);
nand U4632 (N_4632,N_3223,N_2597);
xor U4633 (N_4633,N_2737,N_3128);
nor U4634 (N_4634,N_2528,N_2719);
nand U4635 (N_4635,N_2003,N_2972);
and U4636 (N_4636,N_2809,N_2317);
nor U4637 (N_4637,N_2879,N_2229);
and U4638 (N_4638,N_3762,N_3373);
nand U4639 (N_4639,N_3131,N_2847);
nor U4640 (N_4640,N_3284,N_2224);
nor U4641 (N_4641,N_3937,N_2157);
nand U4642 (N_4642,N_2798,N_3089);
nor U4643 (N_4643,N_2006,N_2059);
nand U4644 (N_4644,N_2241,N_2756);
nand U4645 (N_4645,N_2652,N_2373);
nand U4646 (N_4646,N_2260,N_3915);
nand U4647 (N_4647,N_3535,N_2577);
or U4648 (N_4648,N_2880,N_3187);
or U4649 (N_4649,N_2116,N_3508);
and U4650 (N_4650,N_3704,N_3758);
nand U4651 (N_4651,N_3878,N_2836);
nand U4652 (N_4652,N_3866,N_2889);
xnor U4653 (N_4653,N_3005,N_2439);
nand U4654 (N_4654,N_2740,N_3359);
nand U4655 (N_4655,N_2429,N_3683);
and U4656 (N_4656,N_2519,N_3820);
and U4657 (N_4657,N_2037,N_2986);
and U4658 (N_4658,N_3317,N_2092);
nand U4659 (N_4659,N_2261,N_3936);
and U4660 (N_4660,N_2886,N_2225);
and U4661 (N_4661,N_3766,N_2426);
and U4662 (N_4662,N_2480,N_3111);
or U4663 (N_4663,N_3266,N_3802);
or U4664 (N_4664,N_2023,N_3147);
and U4665 (N_4665,N_2511,N_2323);
nor U4666 (N_4666,N_3901,N_3538);
nor U4667 (N_4667,N_2990,N_2684);
nor U4668 (N_4668,N_2143,N_2854);
or U4669 (N_4669,N_3885,N_2521);
nor U4670 (N_4670,N_2940,N_3689);
and U4671 (N_4671,N_3242,N_3398);
or U4672 (N_4672,N_3428,N_2232);
nor U4673 (N_4673,N_2049,N_3214);
nor U4674 (N_4674,N_2002,N_3737);
and U4675 (N_4675,N_2821,N_2063);
nor U4676 (N_4676,N_2078,N_3150);
nand U4677 (N_4677,N_2808,N_3007);
or U4678 (N_4678,N_3671,N_3698);
or U4679 (N_4679,N_3631,N_2052);
and U4680 (N_4680,N_2748,N_2028);
nand U4681 (N_4681,N_2105,N_3638);
and U4682 (N_4682,N_2156,N_3098);
and U4683 (N_4683,N_3192,N_3983);
nand U4684 (N_4684,N_2197,N_2746);
or U4685 (N_4685,N_3405,N_2381);
nor U4686 (N_4686,N_2666,N_3988);
and U4687 (N_4687,N_3867,N_3929);
nor U4688 (N_4688,N_3069,N_2307);
nor U4689 (N_4689,N_3243,N_2148);
nor U4690 (N_4690,N_3040,N_2149);
and U4691 (N_4691,N_2192,N_3708);
and U4692 (N_4692,N_3752,N_3108);
nand U4693 (N_4693,N_2581,N_2863);
or U4694 (N_4694,N_2425,N_2832);
and U4695 (N_4695,N_2135,N_2755);
and U4696 (N_4696,N_3922,N_3824);
or U4697 (N_4697,N_2546,N_2706);
or U4698 (N_4698,N_3868,N_2102);
and U4699 (N_4699,N_3848,N_2609);
nand U4700 (N_4700,N_2621,N_2014);
or U4701 (N_4701,N_3520,N_2966);
nand U4702 (N_4702,N_3896,N_2019);
nand U4703 (N_4703,N_2106,N_2788);
nor U4704 (N_4704,N_2754,N_2704);
nor U4705 (N_4705,N_3705,N_2407);
nand U4706 (N_4706,N_2065,N_2432);
or U4707 (N_4707,N_2455,N_3023);
or U4708 (N_4708,N_2018,N_2801);
nand U4709 (N_4709,N_2141,N_3021);
nand U4710 (N_4710,N_2100,N_3593);
or U4711 (N_4711,N_3496,N_2595);
and U4712 (N_4712,N_3829,N_2170);
xnor U4713 (N_4713,N_3808,N_2837);
and U4714 (N_4714,N_2377,N_2924);
nor U4715 (N_4715,N_2450,N_3340);
nand U4716 (N_4716,N_3528,N_2036);
nand U4717 (N_4717,N_3055,N_2929);
nor U4718 (N_4718,N_2445,N_2846);
nor U4719 (N_4719,N_3483,N_2698);
nand U4720 (N_4720,N_2976,N_3434);
or U4721 (N_4721,N_2017,N_3489);
nand U4722 (N_4722,N_3914,N_2599);
nor U4723 (N_4723,N_2311,N_2790);
nor U4724 (N_4724,N_3537,N_3110);
or U4725 (N_4725,N_3329,N_2762);
nand U4726 (N_4726,N_2270,N_3609);
or U4727 (N_4727,N_2125,N_2969);
or U4728 (N_4728,N_3142,N_2742);
nand U4729 (N_4729,N_3545,N_3814);
or U4730 (N_4730,N_2159,N_2549);
or U4731 (N_4731,N_2682,N_3913);
nand U4732 (N_4732,N_2349,N_3945);
nor U4733 (N_4733,N_3887,N_2366);
nand U4734 (N_4734,N_3224,N_3636);
or U4735 (N_4735,N_3376,N_3559);
nor U4736 (N_4736,N_2235,N_3550);
nand U4737 (N_4737,N_3260,N_2654);
nand U4738 (N_4738,N_3195,N_2205);
nand U4739 (N_4739,N_3932,N_2328);
nor U4740 (N_4740,N_3697,N_2646);
and U4741 (N_4741,N_3249,N_3971);
and U4742 (N_4742,N_2147,N_3095);
and U4743 (N_4743,N_2277,N_2448);
nor U4744 (N_4744,N_3409,N_3383);
or U4745 (N_4745,N_2630,N_2000);
nand U4746 (N_4746,N_2293,N_2645);
nand U4747 (N_4747,N_3102,N_3327);
nor U4748 (N_4748,N_2492,N_2025);
or U4749 (N_4749,N_2042,N_2776);
and U4750 (N_4750,N_2239,N_2099);
nand U4751 (N_4751,N_3840,N_3426);
nand U4752 (N_4752,N_2834,N_3924);
and U4753 (N_4753,N_3032,N_2804);
or U4754 (N_4754,N_3842,N_3109);
or U4755 (N_4755,N_2182,N_3288);
or U4756 (N_4756,N_3806,N_3380);
or U4757 (N_4757,N_2658,N_2795);
and U4758 (N_4758,N_3747,N_2344);
nand U4759 (N_4759,N_2568,N_3318);
nand U4760 (N_4760,N_2632,N_2334);
or U4761 (N_4761,N_2051,N_2673);
or U4762 (N_4762,N_2227,N_3822);
nand U4763 (N_4763,N_2505,N_2921);
or U4764 (N_4764,N_2862,N_3101);
nand U4765 (N_4765,N_2759,N_2623);
or U4766 (N_4766,N_3144,N_3001);
and U4767 (N_4767,N_2720,N_3063);
nand U4768 (N_4768,N_2233,N_2086);
xor U4769 (N_4769,N_2618,N_3783);
xnor U4770 (N_4770,N_3442,N_3891);
nand U4771 (N_4771,N_3153,N_2977);
nor U4772 (N_4772,N_2001,N_2346);
or U4773 (N_4773,N_2274,N_3278);
xor U4774 (N_4774,N_3046,N_3903);
nor U4775 (N_4775,N_2324,N_2529);
or U4776 (N_4776,N_3399,N_3397);
nand U4777 (N_4777,N_3660,N_2440);
nor U4778 (N_4778,N_3594,N_3188);
xnor U4779 (N_4779,N_2084,N_2872);
or U4780 (N_4780,N_3818,N_2661);
nand U4781 (N_4781,N_2464,N_2191);
or U4782 (N_4782,N_3279,N_2462);
nand U4783 (N_4783,N_3571,N_3735);
nor U4784 (N_4784,N_3574,N_3037);
xnor U4785 (N_4785,N_2656,N_2979);
and U4786 (N_4786,N_2249,N_2015);
and U4787 (N_4787,N_3987,N_2478);
and U4788 (N_4788,N_3668,N_2992);
or U4789 (N_4789,N_2891,N_3706);
and U4790 (N_4790,N_2576,N_3152);
and U4791 (N_4791,N_3504,N_3097);
nor U4792 (N_4792,N_2687,N_2113);
nand U4793 (N_4793,N_2787,N_2031);
or U4794 (N_4794,N_2465,N_3237);
nor U4795 (N_4795,N_3521,N_3396);
and U4796 (N_4796,N_3364,N_2357);
nand U4797 (N_4797,N_2551,N_2841);
and U4798 (N_4798,N_2922,N_3861);
nand U4799 (N_4799,N_2538,N_2446);
nand U4800 (N_4800,N_2248,N_2275);
nand U4801 (N_4801,N_3457,N_2162);
and U4802 (N_4802,N_3964,N_2219);
and U4803 (N_4803,N_2237,N_2294);
xor U4804 (N_4804,N_3159,N_3375);
nor U4805 (N_4805,N_3420,N_3665);
nor U4806 (N_4806,N_3471,N_3759);
and U4807 (N_4807,N_2503,N_2593);
nor U4808 (N_4808,N_2591,N_3985);
nor U4809 (N_4809,N_2965,N_3350);
nor U4810 (N_4810,N_3184,N_2570);
nand U4811 (N_4811,N_2475,N_3807);
xnor U4812 (N_4812,N_3299,N_2797);
or U4813 (N_4813,N_2784,N_2213);
nor U4814 (N_4814,N_2587,N_2295);
and U4815 (N_4815,N_3799,N_2867);
nor U4816 (N_4816,N_3310,N_2541);
nor U4817 (N_4817,N_2647,N_3370);
and U4818 (N_4818,N_2032,N_3407);
nor U4819 (N_4819,N_3476,N_2850);
or U4820 (N_4820,N_2438,N_3933);
and U4821 (N_4821,N_2314,N_3541);
nor U4822 (N_4822,N_2978,N_2711);
nor U4823 (N_4823,N_2145,N_2864);
and U4824 (N_4824,N_3552,N_3304);
and U4825 (N_4825,N_2271,N_3512);
nor U4826 (N_4826,N_3693,N_3635);
nor U4827 (N_4827,N_2313,N_2456);
or U4828 (N_4828,N_3136,N_3332);
nor U4829 (N_4829,N_3422,N_2244);
and U4830 (N_4830,N_3194,N_2567);
xor U4831 (N_4831,N_2178,N_2497);
or U4832 (N_4832,N_3427,N_3418);
nor U4833 (N_4833,N_3262,N_3220);
nand U4834 (N_4834,N_2985,N_3484);
and U4835 (N_4835,N_3378,N_3222);
xnor U4836 (N_4836,N_2123,N_3580);
nand U4837 (N_4837,N_3425,N_2960);
or U4838 (N_4838,N_3257,N_2126);
nor U4839 (N_4839,N_3301,N_3099);
xor U4840 (N_4840,N_3186,N_3293);
nor U4841 (N_4841,N_3676,N_2535);
nor U4842 (N_4842,N_2590,N_3850);
or U4843 (N_4843,N_2369,N_2533);
or U4844 (N_4844,N_3935,N_2583);
or U4845 (N_4845,N_2806,N_2758);
nor U4846 (N_4846,N_2291,N_2473);
nand U4847 (N_4847,N_2987,N_3796);
xor U4848 (N_4848,N_2210,N_3346);
nand U4849 (N_4849,N_3343,N_2174);
nor U4850 (N_4850,N_3250,N_3408);
and U4851 (N_4851,N_3534,N_3256);
nor U4852 (N_4852,N_3233,N_3477);
and U4853 (N_4853,N_3114,N_2231);
nor U4854 (N_4854,N_3435,N_3121);
nor U4855 (N_4855,N_3926,N_2208);
or U4856 (N_4856,N_3149,N_2894);
nand U4857 (N_4857,N_3210,N_2669);
or U4858 (N_4858,N_2090,N_3529);
nand U4859 (N_4859,N_2485,N_3049);
nor U4860 (N_4860,N_2410,N_2144);
nor U4861 (N_4861,N_2817,N_3522);
nor U4862 (N_4862,N_3610,N_2594);
nand U4863 (N_4863,N_2997,N_2088);
nand U4864 (N_4864,N_2683,N_2953);
nand U4865 (N_4865,N_3918,N_3404);
nand U4866 (N_4866,N_2648,N_2012);
and U4867 (N_4867,N_3813,N_3772);
or U4868 (N_4868,N_2600,N_2154);
and U4869 (N_4869,N_3618,N_3173);
or U4870 (N_4870,N_2447,N_3513);
nand U4871 (N_4871,N_3067,N_3886);
and U4872 (N_4872,N_2343,N_2163);
and U4873 (N_4873,N_2803,N_2097);
nor U4874 (N_4874,N_3774,N_3026);
nand U4875 (N_4875,N_2424,N_2911);
nand U4876 (N_4876,N_2083,N_2907);
nand U4877 (N_4877,N_3429,N_2121);
or U4878 (N_4878,N_2056,N_2322);
and U4879 (N_4879,N_2944,N_2073);
or U4880 (N_4880,N_2382,N_2509);
nor U4881 (N_4881,N_3162,N_2262);
or U4882 (N_4882,N_2974,N_3302);
and U4883 (N_4883,N_3107,N_2379);
nor U4884 (N_4884,N_3560,N_3221);
nand U4885 (N_4885,N_2142,N_3319);
and U4886 (N_4886,N_3123,N_2474);
and U4887 (N_4887,N_2458,N_2773);
nor U4888 (N_4888,N_3567,N_3778);
xor U4889 (N_4889,N_3076,N_2068);
nor U4890 (N_4890,N_3606,N_2726);
nand U4891 (N_4891,N_3780,N_3156);
or U4892 (N_4892,N_3006,N_3626);
nor U4893 (N_4893,N_2222,N_3349);
nor U4894 (N_4894,N_2266,N_3619);
or U4895 (N_4895,N_3839,N_2461);
nand U4896 (N_4896,N_3894,N_2185);
or U4897 (N_4897,N_2610,N_2221);
and U4898 (N_4898,N_2715,N_2013);
nor U4899 (N_4899,N_3823,N_2885);
and U4900 (N_4900,N_3406,N_3019);
and U4901 (N_4901,N_2414,N_2739);
nand U4902 (N_4902,N_3402,N_3904);
nor U4903 (N_4903,N_3342,N_3916);
and U4904 (N_4904,N_2878,N_3603);
nor U4905 (N_4905,N_3203,N_3812);
or U4906 (N_4906,N_3722,N_2712);
or U4907 (N_4907,N_2805,N_3837);
nand U4908 (N_4908,N_3666,N_3423);
and U4909 (N_4909,N_3316,N_3615);
or U4910 (N_4910,N_3794,N_3892);
and U4911 (N_4911,N_3269,N_2578);
and U4912 (N_4912,N_3010,N_2936);
nor U4913 (N_4913,N_3433,N_3093);
nand U4914 (N_4914,N_3036,N_2625);
nor U4915 (N_4915,N_3849,N_3449);
xor U4916 (N_4916,N_2793,N_2749);
nor U4917 (N_4917,N_2901,N_3495);
or U4918 (N_4918,N_2663,N_3085);
nand U4919 (N_4919,N_3480,N_2207);
nor U4920 (N_4920,N_3092,N_3446);
nand U4921 (N_4921,N_3462,N_2643);
nand U4922 (N_4922,N_3682,N_2247);
or U4923 (N_4923,N_2553,N_3865);
nor U4924 (N_4924,N_3674,N_2925);
nand U4925 (N_4925,N_3366,N_2436);
nand U4926 (N_4926,N_2904,N_2374);
nor U4927 (N_4927,N_3511,N_2335);
or U4928 (N_4928,N_3589,N_3981);
or U4929 (N_4929,N_3213,N_2747);
nand U4930 (N_4930,N_3900,N_2380);
or U4931 (N_4931,N_3016,N_2449);
nor U4932 (N_4932,N_3413,N_2831);
nor U4933 (N_4933,N_3321,N_2603);
and U4934 (N_4934,N_3716,N_2848);
and U4935 (N_4935,N_3324,N_2444);
and U4936 (N_4936,N_3569,N_2111);
nor U4937 (N_4937,N_3417,N_2409);
or U4938 (N_4938,N_2008,N_2312);
and U4939 (N_4939,N_3957,N_3883);
and U4940 (N_4940,N_2508,N_2048);
and U4941 (N_4941,N_3973,N_3277);
nor U4942 (N_4942,N_2882,N_2360);
and U4943 (N_4943,N_2067,N_2039);
nor U4944 (N_4944,N_3944,N_3481);
or U4945 (N_4945,N_3080,N_3358);
or U4946 (N_4946,N_2993,N_3624);
and U4947 (N_4947,N_3832,N_3970);
nand U4948 (N_4948,N_2181,N_2839);
nor U4949 (N_4949,N_2876,N_2580);
and U4950 (N_4950,N_2081,N_2782);
and U4951 (N_4951,N_3591,N_3436);
and U4952 (N_4952,N_2518,N_2404);
or U4953 (N_4953,N_3009,N_2498);
or U4954 (N_4954,N_2265,N_2071);
nand U4955 (N_4955,N_2327,N_3994);
nand U4956 (N_4956,N_3441,N_2544);
and U4957 (N_4957,N_2416,N_3452);
nand U4958 (N_4958,N_2890,N_2564);
or U4959 (N_4959,N_2351,N_2559);
and U4960 (N_4960,N_3035,N_2246);
or U4961 (N_4961,N_2267,N_2160);
and U4962 (N_4962,N_3670,N_3663);
xnor U4963 (N_4963,N_2318,N_3143);
nor U4964 (N_4964,N_3193,N_2387);
or U4965 (N_4965,N_2844,N_2757);
or U4966 (N_4966,N_2435,N_2331);
and U4967 (N_4967,N_3071,N_2350);
nor U4968 (N_4968,N_3819,N_2070);
nand U4969 (N_4969,N_3877,N_2732);
xnor U4970 (N_4970,N_3283,N_3139);
or U4971 (N_4971,N_3669,N_2766);
and U4972 (N_4972,N_3949,N_3979);
nand U4973 (N_4973,N_2892,N_3738);
nor U4974 (N_4974,N_2321,N_3461);
or U4975 (N_4975,N_3701,N_3485);
and U4976 (N_4976,N_3951,N_2216);
nand U4977 (N_4977,N_3470,N_3155);
and U4978 (N_4978,N_2722,N_3352);
nor U4979 (N_4979,N_3268,N_3801);
nor U4980 (N_4980,N_2750,N_2104);
xor U4981 (N_4981,N_3451,N_2527);
nand U4982 (N_4982,N_2981,N_3696);
or U4983 (N_4983,N_3381,N_3130);
nor U4984 (N_4984,N_2853,N_3743);
or U4985 (N_4985,N_2565,N_2547);
or U4986 (N_4986,N_2356,N_2319);
and U4987 (N_4987,N_2129,N_2272);
nor U4988 (N_4988,N_2589,N_2495);
and U4989 (N_4989,N_3732,N_3907);
nand U4990 (N_4990,N_2761,N_3330);
nand U4991 (N_4991,N_3845,N_2376);
or U4992 (N_4992,N_3015,N_2390);
nand U4993 (N_4993,N_2315,N_3797);
nand U4994 (N_4994,N_2592,N_3444);
or U4995 (N_4995,N_3989,N_2606);
xnor U4996 (N_4996,N_3741,N_3825);
and U4997 (N_4997,N_2869,N_2472);
nor U4998 (N_4998,N_2389,N_2572);
or U4999 (N_4999,N_2903,N_2617);
nor U5000 (N_5000,N_2876,N_2368);
nand U5001 (N_5001,N_3843,N_3090);
or U5002 (N_5002,N_3193,N_3432);
nor U5003 (N_5003,N_2985,N_3733);
nor U5004 (N_5004,N_2430,N_3409);
or U5005 (N_5005,N_2129,N_2070);
nand U5006 (N_5006,N_2869,N_3922);
nand U5007 (N_5007,N_2813,N_3730);
and U5008 (N_5008,N_2577,N_2290);
nor U5009 (N_5009,N_3524,N_2063);
nand U5010 (N_5010,N_2309,N_3229);
nand U5011 (N_5011,N_3687,N_2325);
nand U5012 (N_5012,N_2153,N_3115);
nor U5013 (N_5013,N_2628,N_2990);
and U5014 (N_5014,N_2901,N_2931);
or U5015 (N_5015,N_3015,N_3538);
xnor U5016 (N_5016,N_3623,N_2403);
and U5017 (N_5017,N_3948,N_2704);
or U5018 (N_5018,N_2747,N_3715);
or U5019 (N_5019,N_3109,N_3673);
or U5020 (N_5020,N_2385,N_3079);
nand U5021 (N_5021,N_3746,N_3767);
nor U5022 (N_5022,N_2175,N_3036);
nor U5023 (N_5023,N_3326,N_3043);
and U5024 (N_5024,N_3420,N_3436);
nor U5025 (N_5025,N_2340,N_3793);
and U5026 (N_5026,N_3645,N_2757);
nor U5027 (N_5027,N_3494,N_3450);
nor U5028 (N_5028,N_2452,N_3304);
nand U5029 (N_5029,N_2713,N_3804);
and U5030 (N_5030,N_2142,N_3101);
and U5031 (N_5031,N_2947,N_2358);
nor U5032 (N_5032,N_3488,N_2540);
or U5033 (N_5033,N_2483,N_3936);
and U5034 (N_5034,N_3237,N_3042);
and U5035 (N_5035,N_3834,N_2766);
or U5036 (N_5036,N_2497,N_3918);
and U5037 (N_5037,N_2295,N_2876);
xnor U5038 (N_5038,N_2599,N_3436);
nand U5039 (N_5039,N_2073,N_2736);
or U5040 (N_5040,N_2046,N_2397);
nand U5041 (N_5041,N_2778,N_3011);
or U5042 (N_5042,N_3510,N_3877);
nor U5043 (N_5043,N_2959,N_3853);
or U5044 (N_5044,N_2445,N_3647);
nor U5045 (N_5045,N_2319,N_2022);
nand U5046 (N_5046,N_3014,N_3641);
nor U5047 (N_5047,N_3978,N_2915);
nor U5048 (N_5048,N_3078,N_3927);
or U5049 (N_5049,N_2719,N_2989);
nand U5050 (N_5050,N_2770,N_2416);
and U5051 (N_5051,N_3962,N_3065);
nor U5052 (N_5052,N_2298,N_2235);
or U5053 (N_5053,N_2763,N_2370);
nand U5054 (N_5054,N_3149,N_3532);
or U5055 (N_5055,N_2296,N_2902);
or U5056 (N_5056,N_3345,N_2239);
or U5057 (N_5057,N_2940,N_2294);
and U5058 (N_5058,N_3220,N_3087);
nor U5059 (N_5059,N_2036,N_3718);
or U5060 (N_5060,N_2087,N_2272);
and U5061 (N_5061,N_3669,N_2130);
and U5062 (N_5062,N_2645,N_2898);
or U5063 (N_5063,N_3404,N_3558);
and U5064 (N_5064,N_2584,N_3315);
xor U5065 (N_5065,N_3189,N_3322);
and U5066 (N_5066,N_2342,N_3887);
and U5067 (N_5067,N_3643,N_3797);
or U5068 (N_5068,N_2790,N_3071);
xnor U5069 (N_5069,N_2157,N_3472);
and U5070 (N_5070,N_3683,N_2455);
nor U5071 (N_5071,N_3950,N_2022);
nor U5072 (N_5072,N_2294,N_2066);
nor U5073 (N_5073,N_2251,N_3065);
nand U5074 (N_5074,N_3914,N_3896);
nand U5075 (N_5075,N_2739,N_3868);
xor U5076 (N_5076,N_2228,N_3195);
nor U5077 (N_5077,N_2974,N_2971);
nand U5078 (N_5078,N_3260,N_2430);
xnor U5079 (N_5079,N_2024,N_3962);
nand U5080 (N_5080,N_3370,N_3950);
nand U5081 (N_5081,N_3249,N_2357);
nand U5082 (N_5082,N_3268,N_3568);
nor U5083 (N_5083,N_3829,N_2620);
nand U5084 (N_5084,N_3443,N_3363);
or U5085 (N_5085,N_2274,N_3095);
nand U5086 (N_5086,N_3896,N_2161);
nand U5087 (N_5087,N_2044,N_2351);
and U5088 (N_5088,N_3012,N_3700);
and U5089 (N_5089,N_2318,N_2562);
nand U5090 (N_5090,N_3377,N_2635);
nor U5091 (N_5091,N_2869,N_3313);
nor U5092 (N_5092,N_2919,N_2062);
nand U5093 (N_5093,N_3282,N_3878);
nand U5094 (N_5094,N_3636,N_3607);
nor U5095 (N_5095,N_3362,N_2552);
and U5096 (N_5096,N_2029,N_2126);
and U5097 (N_5097,N_2368,N_2925);
or U5098 (N_5098,N_3070,N_3972);
nand U5099 (N_5099,N_3048,N_2166);
and U5100 (N_5100,N_2849,N_3259);
nor U5101 (N_5101,N_2066,N_2158);
and U5102 (N_5102,N_2172,N_3317);
nor U5103 (N_5103,N_2563,N_3273);
nand U5104 (N_5104,N_2515,N_3828);
xnor U5105 (N_5105,N_3116,N_2514);
nand U5106 (N_5106,N_2591,N_2871);
and U5107 (N_5107,N_2286,N_2619);
nand U5108 (N_5108,N_2568,N_3678);
nor U5109 (N_5109,N_3730,N_3069);
nand U5110 (N_5110,N_2430,N_3194);
nand U5111 (N_5111,N_2303,N_3648);
nand U5112 (N_5112,N_2264,N_2860);
nand U5113 (N_5113,N_3809,N_2195);
nand U5114 (N_5114,N_3548,N_3983);
nor U5115 (N_5115,N_2525,N_3381);
and U5116 (N_5116,N_2605,N_3910);
nand U5117 (N_5117,N_3324,N_3613);
or U5118 (N_5118,N_3082,N_2081);
or U5119 (N_5119,N_3564,N_2437);
and U5120 (N_5120,N_2438,N_2650);
nor U5121 (N_5121,N_2046,N_3678);
and U5122 (N_5122,N_3197,N_2550);
nand U5123 (N_5123,N_3177,N_2422);
or U5124 (N_5124,N_3943,N_2064);
and U5125 (N_5125,N_3783,N_2619);
nor U5126 (N_5126,N_3323,N_3149);
nor U5127 (N_5127,N_3581,N_2423);
or U5128 (N_5128,N_2525,N_3701);
nor U5129 (N_5129,N_3196,N_2129);
nand U5130 (N_5130,N_3875,N_3530);
and U5131 (N_5131,N_3381,N_3800);
or U5132 (N_5132,N_3702,N_3113);
or U5133 (N_5133,N_2591,N_2481);
nand U5134 (N_5134,N_3127,N_2965);
and U5135 (N_5135,N_2637,N_2894);
nor U5136 (N_5136,N_2568,N_2848);
nand U5137 (N_5137,N_2281,N_3438);
and U5138 (N_5138,N_2106,N_2063);
and U5139 (N_5139,N_3825,N_3479);
nor U5140 (N_5140,N_3862,N_3355);
nand U5141 (N_5141,N_2310,N_2547);
nor U5142 (N_5142,N_3424,N_3319);
nor U5143 (N_5143,N_3933,N_3623);
nand U5144 (N_5144,N_2873,N_2841);
or U5145 (N_5145,N_3897,N_2728);
nor U5146 (N_5146,N_2968,N_2432);
or U5147 (N_5147,N_3624,N_3317);
nand U5148 (N_5148,N_2196,N_3832);
and U5149 (N_5149,N_2500,N_3798);
nand U5150 (N_5150,N_3185,N_3167);
or U5151 (N_5151,N_3779,N_3078);
or U5152 (N_5152,N_2791,N_2179);
xor U5153 (N_5153,N_2299,N_3083);
xnor U5154 (N_5154,N_2294,N_2566);
and U5155 (N_5155,N_2641,N_2622);
or U5156 (N_5156,N_3081,N_2249);
or U5157 (N_5157,N_3092,N_2142);
or U5158 (N_5158,N_3406,N_3246);
nor U5159 (N_5159,N_2161,N_3637);
and U5160 (N_5160,N_3055,N_2229);
nor U5161 (N_5161,N_2591,N_2712);
and U5162 (N_5162,N_2000,N_2279);
nand U5163 (N_5163,N_3162,N_2906);
or U5164 (N_5164,N_2684,N_2121);
nand U5165 (N_5165,N_3769,N_3086);
and U5166 (N_5166,N_2073,N_3491);
nand U5167 (N_5167,N_2868,N_2934);
or U5168 (N_5168,N_3209,N_3867);
or U5169 (N_5169,N_2742,N_3856);
and U5170 (N_5170,N_2837,N_2494);
nand U5171 (N_5171,N_3334,N_3008);
or U5172 (N_5172,N_2326,N_2597);
nor U5173 (N_5173,N_3250,N_3877);
and U5174 (N_5174,N_3777,N_2815);
or U5175 (N_5175,N_3800,N_2814);
and U5176 (N_5176,N_3888,N_2167);
or U5177 (N_5177,N_3001,N_3471);
nand U5178 (N_5178,N_3249,N_3843);
or U5179 (N_5179,N_3322,N_2940);
or U5180 (N_5180,N_3943,N_3541);
nor U5181 (N_5181,N_3596,N_3493);
nand U5182 (N_5182,N_2912,N_3758);
or U5183 (N_5183,N_2075,N_2988);
and U5184 (N_5184,N_3839,N_3550);
or U5185 (N_5185,N_3851,N_2719);
nand U5186 (N_5186,N_3395,N_2683);
nand U5187 (N_5187,N_2066,N_3731);
nand U5188 (N_5188,N_2850,N_2467);
nor U5189 (N_5189,N_2371,N_3012);
nand U5190 (N_5190,N_2714,N_2205);
and U5191 (N_5191,N_2135,N_3093);
or U5192 (N_5192,N_3223,N_3062);
or U5193 (N_5193,N_2175,N_3732);
nand U5194 (N_5194,N_3807,N_2180);
xnor U5195 (N_5195,N_3263,N_2098);
and U5196 (N_5196,N_2183,N_2646);
and U5197 (N_5197,N_3331,N_3204);
nand U5198 (N_5198,N_2024,N_2523);
and U5199 (N_5199,N_3503,N_3413);
or U5200 (N_5200,N_3229,N_2126);
or U5201 (N_5201,N_3328,N_3542);
or U5202 (N_5202,N_2882,N_3942);
nor U5203 (N_5203,N_2617,N_2108);
and U5204 (N_5204,N_2628,N_2787);
or U5205 (N_5205,N_2546,N_3699);
and U5206 (N_5206,N_2941,N_2902);
and U5207 (N_5207,N_2731,N_2951);
nor U5208 (N_5208,N_2599,N_3600);
and U5209 (N_5209,N_2587,N_3530);
and U5210 (N_5210,N_2156,N_2163);
nand U5211 (N_5211,N_2167,N_2081);
and U5212 (N_5212,N_2218,N_2770);
nand U5213 (N_5213,N_3776,N_3078);
nor U5214 (N_5214,N_3421,N_2955);
nor U5215 (N_5215,N_2689,N_2841);
and U5216 (N_5216,N_3751,N_3306);
or U5217 (N_5217,N_2382,N_3683);
xor U5218 (N_5218,N_2379,N_2805);
or U5219 (N_5219,N_2535,N_2895);
nand U5220 (N_5220,N_3151,N_3377);
xnor U5221 (N_5221,N_2698,N_3913);
nand U5222 (N_5222,N_2754,N_3844);
nand U5223 (N_5223,N_2713,N_3680);
or U5224 (N_5224,N_2118,N_3503);
or U5225 (N_5225,N_3281,N_3882);
and U5226 (N_5226,N_2487,N_3860);
nor U5227 (N_5227,N_2335,N_2654);
nand U5228 (N_5228,N_2822,N_3419);
and U5229 (N_5229,N_3988,N_2665);
and U5230 (N_5230,N_2564,N_2123);
nor U5231 (N_5231,N_2435,N_2042);
or U5232 (N_5232,N_2865,N_2399);
and U5233 (N_5233,N_3316,N_3903);
and U5234 (N_5234,N_2532,N_2715);
nand U5235 (N_5235,N_2702,N_3875);
nor U5236 (N_5236,N_3797,N_2877);
nand U5237 (N_5237,N_2987,N_3391);
and U5238 (N_5238,N_3429,N_3774);
and U5239 (N_5239,N_3288,N_3964);
and U5240 (N_5240,N_2190,N_3834);
and U5241 (N_5241,N_3658,N_2791);
nand U5242 (N_5242,N_3945,N_2352);
nor U5243 (N_5243,N_2303,N_2519);
nor U5244 (N_5244,N_3612,N_2252);
nand U5245 (N_5245,N_2843,N_2024);
nor U5246 (N_5246,N_3639,N_2361);
nor U5247 (N_5247,N_3166,N_3664);
or U5248 (N_5248,N_3435,N_3041);
nand U5249 (N_5249,N_3871,N_2726);
and U5250 (N_5250,N_2549,N_2163);
xnor U5251 (N_5251,N_3878,N_2291);
or U5252 (N_5252,N_2099,N_2828);
and U5253 (N_5253,N_2269,N_3530);
and U5254 (N_5254,N_2301,N_3498);
and U5255 (N_5255,N_3314,N_2625);
nor U5256 (N_5256,N_2999,N_2406);
nor U5257 (N_5257,N_2309,N_3687);
nand U5258 (N_5258,N_3181,N_3102);
nand U5259 (N_5259,N_2671,N_3383);
and U5260 (N_5260,N_2378,N_2481);
nor U5261 (N_5261,N_3245,N_2596);
or U5262 (N_5262,N_2198,N_3762);
nand U5263 (N_5263,N_3996,N_2912);
or U5264 (N_5264,N_2656,N_2454);
nor U5265 (N_5265,N_3124,N_3846);
xor U5266 (N_5266,N_3196,N_3012);
and U5267 (N_5267,N_2066,N_3078);
or U5268 (N_5268,N_3597,N_3567);
nor U5269 (N_5269,N_3000,N_3363);
nand U5270 (N_5270,N_2261,N_3625);
nor U5271 (N_5271,N_2451,N_3602);
and U5272 (N_5272,N_3323,N_2588);
and U5273 (N_5273,N_3809,N_3253);
xnor U5274 (N_5274,N_3280,N_2710);
or U5275 (N_5275,N_2433,N_3535);
or U5276 (N_5276,N_3109,N_3854);
or U5277 (N_5277,N_3948,N_3355);
or U5278 (N_5278,N_3081,N_3685);
or U5279 (N_5279,N_3460,N_2098);
and U5280 (N_5280,N_3142,N_3981);
and U5281 (N_5281,N_3787,N_3134);
xor U5282 (N_5282,N_2623,N_3236);
nand U5283 (N_5283,N_2875,N_2528);
or U5284 (N_5284,N_3078,N_3089);
nor U5285 (N_5285,N_2910,N_3223);
nor U5286 (N_5286,N_3883,N_3119);
or U5287 (N_5287,N_3169,N_3582);
nor U5288 (N_5288,N_2134,N_2028);
or U5289 (N_5289,N_2644,N_2886);
nand U5290 (N_5290,N_2878,N_3124);
or U5291 (N_5291,N_2133,N_2815);
nand U5292 (N_5292,N_2046,N_2375);
nor U5293 (N_5293,N_3210,N_2350);
or U5294 (N_5294,N_2555,N_3563);
nor U5295 (N_5295,N_3529,N_2184);
and U5296 (N_5296,N_3913,N_3017);
nand U5297 (N_5297,N_2990,N_3119);
and U5298 (N_5298,N_2339,N_3513);
nor U5299 (N_5299,N_2331,N_2049);
nand U5300 (N_5300,N_2805,N_2608);
and U5301 (N_5301,N_2377,N_3378);
or U5302 (N_5302,N_2235,N_2788);
nand U5303 (N_5303,N_3913,N_3470);
nand U5304 (N_5304,N_3203,N_3341);
and U5305 (N_5305,N_2782,N_3903);
or U5306 (N_5306,N_2977,N_2898);
nand U5307 (N_5307,N_3234,N_2723);
nand U5308 (N_5308,N_2122,N_2879);
or U5309 (N_5309,N_3743,N_2867);
nor U5310 (N_5310,N_3225,N_2580);
or U5311 (N_5311,N_2303,N_2623);
nor U5312 (N_5312,N_3986,N_3356);
nor U5313 (N_5313,N_3359,N_3014);
nor U5314 (N_5314,N_3277,N_2871);
nand U5315 (N_5315,N_2462,N_2050);
or U5316 (N_5316,N_2991,N_3651);
nand U5317 (N_5317,N_3976,N_2295);
or U5318 (N_5318,N_3833,N_2976);
or U5319 (N_5319,N_2990,N_2752);
nor U5320 (N_5320,N_3677,N_2788);
and U5321 (N_5321,N_2259,N_2602);
nand U5322 (N_5322,N_3371,N_3833);
or U5323 (N_5323,N_2497,N_2966);
nand U5324 (N_5324,N_2838,N_2484);
or U5325 (N_5325,N_2346,N_3015);
and U5326 (N_5326,N_2148,N_2633);
or U5327 (N_5327,N_3737,N_2448);
nor U5328 (N_5328,N_3418,N_3581);
or U5329 (N_5329,N_3991,N_2368);
and U5330 (N_5330,N_3493,N_2697);
nand U5331 (N_5331,N_2060,N_3879);
and U5332 (N_5332,N_3922,N_2282);
nand U5333 (N_5333,N_3542,N_3882);
nand U5334 (N_5334,N_3304,N_2520);
nor U5335 (N_5335,N_3470,N_2160);
or U5336 (N_5336,N_3820,N_3816);
or U5337 (N_5337,N_2500,N_2008);
nand U5338 (N_5338,N_2651,N_3077);
nor U5339 (N_5339,N_2971,N_3233);
nand U5340 (N_5340,N_2326,N_2357);
and U5341 (N_5341,N_2655,N_2020);
and U5342 (N_5342,N_2096,N_3314);
or U5343 (N_5343,N_2756,N_3928);
nor U5344 (N_5344,N_2900,N_2279);
nand U5345 (N_5345,N_3651,N_3414);
nand U5346 (N_5346,N_2792,N_3842);
or U5347 (N_5347,N_3477,N_2899);
nand U5348 (N_5348,N_3790,N_2925);
nand U5349 (N_5349,N_3964,N_2851);
or U5350 (N_5350,N_3802,N_3994);
and U5351 (N_5351,N_3357,N_2316);
nand U5352 (N_5352,N_2072,N_3005);
or U5353 (N_5353,N_3196,N_3830);
and U5354 (N_5354,N_2882,N_2843);
and U5355 (N_5355,N_3435,N_3710);
or U5356 (N_5356,N_3965,N_2286);
nand U5357 (N_5357,N_2787,N_2674);
and U5358 (N_5358,N_3289,N_2131);
or U5359 (N_5359,N_2795,N_2623);
or U5360 (N_5360,N_3888,N_2501);
and U5361 (N_5361,N_3250,N_2938);
and U5362 (N_5362,N_2244,N_3782);
or U5363 (N_5363,N_2994,N_2157);
nand U5364 (N_5364,N_3584,N_3565);
and U5365 (N_5365,N_2374,N_2460);
or U5366 (N_5366,N_3825,N_2407);
and U5367 (N_5367,N_3495,N_3913);
or U5368 (N_5368,N_3001,N_2715);
nand U5369 (N_5369,N_3138,N_2613);
nor U5370 (N_5370,N_2909,N_2213);
or U5371 (N_5371,N_2748,N_3354);
or U5372 (N_5372,N_3965,N_3409);
nand U5373 (N_5373,N_3771,N_3549);
or U5374 (N_5374,N_3100,N_2991);
nand U5375 (N_5375,N_3109,N_3564);
nand U5376 (N_5376,N_3527,N_3751);
and U5377 (N_5377,N_3690,N_3271);
or U5378 (N_5378,N_3477,N_3061);
nor U5379 (N_5379,N_3496,N_3321);
nor U5380 (N_5380,N_3097,N_2638);
nand U5381 (N_5381,N_2103,N_2356);
or U5382 (N_5382,N_3606,N_2009);
nor U5383 (N_5383,N_2235,N_2621);
or U5384 (N_5384,N_2759,N_3053);
nand U5385 (N_5385,N_3475,N_2547);
nand U5386 (N_5386,N_3011,N_3541);
or U5387 (N_5387,N_2737,N_2880);
and U5388 (N_5388,N_2290,N_3854);
and U5389 (N_5389,N_3192,N_2387);
nand U5390 (N_5390,N_3932,N_2933);
and U5391 (N_5391,N_3532,N_2314);
nand U5392 (N_5392,N_3823,N_2828);
nand U5393 (N_5393,N_2348,N_2437);
and U5394 (N_5394,N_3318,N_3695);
and U5395 (N_5395,N_3115,N_2149);
nand U5396 (N_5396,N_2319,N_3971);
and U5397 (N_5397,N_2978,N_2446);
nand U5398 (N_5398,N_3557,N_2517);
or U5399 (N_5399,N_2737,N_3765);
and U5400 (N_5400,N_2581,N_3115);
and U5401 (N_5401,N_2263,N_3177);
xnor U5402 (N_5402,N_2708,N_3516);
and U5403 (N_5403,N_3091,N_3025);
or U5404 (N_5404,N_3728,N_2092);
and U5405 (N_5405,N_2144,N_2291);
nand U5406 (N_5406,N_2206,N_2927);
nand U5407 (N_5407,N_2169,N_2109);
nand U5408 (N_5408,N_2546,N_3593);
and U5409 (N_5409,N_2762,N_2513);
and U5410 (N_5410,N_2236,N_2976);
and U5411 (N_5411,N_2688,N_2799);
or U5412 (N_5412,N_2772,N_3646);
nand U5413 (N_5413,N_3018,N_2836);
or U5414 (N_5414,N_2104,N_2113);
or U5415 (N_5415,N_3924,N_2951);
and U5416 (N_5416,N_2948,N_3427);
nand U5417 (N_5417,N_2502,N_2224);
or U5418 (N_5418,N_3261,N_3946);
nand U5419 (N_5419,N_3415,N_3117);
or U5420 (N_5420,N_2914,N_2050);
and U5421 (N_5421,N_2402,N_2112);
nor U5422 (N_5422,N_2722,N_2767);
nand U5423 (N_5423,N_3445,N_2826);
nand U5424 (N_5424,N_3290,N_3532);
and U5425 (N_5425,N_2374,N_2558);
or U5426 (N_5426,N_2610,N_2415);
nand U5427 (N_5427,N_2852,N_3825);
nor U5428 (N_5428,N_2949,N_2161);
or U5429 (N_5429,N_2286,N_3202);
nor U5430 (N_5430,N_3004,N_3470);
or U5431 (N_5431,N_3267,N_2318);
or U5432 (N_5432,N_3379,N_2422);
and U5433 (N_5433,N_3647,N_3073);
or U5434 (N_5434,N_3108,N_3288);
and U5435 (N_5435,N_3393,N_3532);
and U5436 (N_5436,N_2568,N_2706);
and U5437 (N_5437,N_2411,N_2169);
nand U5438 (N_5438,N_2223,N_3768);
nand U5439 (N_5439,N_3061,N_3998);
and U5440 (N_5440,N_2078,N_3610);
or U5441 (N_5441,N_3997,N_2030);
and U5442 (N_5442,N_2480,N_2479);
or U5443 (N_5443,N_2850,N_2701);
and U5444 (N_5444,N_2162,N_2445);
and U5445 (N_5445,N_3262,N_2758);
or U5446 (N_5446,N_2363,N_2984);
and U5447 (N_5447,N_2164,N_3988);
and U5448 (N_5448,N_2323,N_2715);
nand U5449 (N_5449,N_3088,N_3857);
or U5450 (N_5450,N_2857,N_3354);
nand U5451 (N_5451,N_3456,N_3484);
and U5452 (N_5452,N_3924,N_2363);
and U5453 (N_5453,N_2998,N_2107);
and U5454 (N_5454,N_2909,N_3859);
nor U5455 (N_5455,N_3274,N_2030);
or U5456 (N_5456,N_3441,N_2601);
or U5457 (N_5457,N_2296,N_3129);
nor U5458 (N_5458,N_3543,N_2249);
xor U5459 (N_5459,N_2193,N_2443);
or U5460 (N_5460,N_2957,N_2195);
or U5461 (N_5461,N_2131,N_2384);
nor U5462 (N_5462,N_2763,N_3090);
nor U5463 (N_5463,N_3333,N_3077);
or U5464 (N_5464,N_3192,N_3636);
and U5465 (N_5465,N_2691,N_3098);
or U5466 (N_5466,N_2395,N_2101);
or U5467 (N_5467,N_3030,N_2167);
or U5468 (N_5468,N_2984,N_2791);
and U5469 (N_5469,N_2582,N_2253);
nand U5470 (N_5470,N_2915,N_3621);
nand U5471 (N_5471,N_2802,N_3638);
nand U5472 (N_5472,N_2951,N_3999);
nand U5473 (N_5473,N_2824,N_2980);
or U5474 (N_5474,N_3338,N_2489);
xnor U5475 (N_5475,N_2553,N_3476);
nand U5476 (N_5476,N_3079,N_2636);
nor U5477 (N_5477,N_2736,N_2354);
nand U5478 (N_5478,N_2929,N_3753);
or U5479 (N_5479,N_3175,N_3640);
or U5480 (N_5480,N_2069,N_2564);
and U5481 (N_5481,N_3997,N_2786);
nand U5482 (N_5482,N_2176,N_3902);
and U5483 (N_5483,N_3339,N_3068);
nor U5484 (N_5484,N_2427,N_3478);
xor U5485 (N_5485,N_2708,N_2196);
and U5486 (N_5486,N_2226,N_2368);
nand U5487 (N_5487,N_2564,N_2313);
nor U5488 (N_5488,N_2030,N_3057);
or U5489 (N_5489,N_2079,N_3594);
nand U5490 (N_5490,N_2482,N_2486);
nand U5491 (N_5491,N_3235,N_2294);
and U5492 (N_5492,N_3854,N_3480);
or U5493 (N_5493,N_2392,N_3236);
nor U5494 (N_5494,N_2966,N_3254);
nor U5495 (N_5495,N_2363,N_2949);
or U5496 (N_5496,N_2608,N_3037);
nand U5497 (N_5497,N_2692,N_3975);
and U5498 (N_5498,N_2809,N_2942);
nand U5499 (N_5499,N_3800,N_3622);
and U5500 (N_5500,N_2781,N_2291);
or U5501 (N_5501,N_2415,N_2351);
and U5502 (N_5502,N_3617,N_3869);
nand U5503 (N_5503,N_3734,N_3675);
and U5504 (N_5504,N_3256,N_3429);
nor U5505 (N_5505,N_3524,N_3600);
and U5506 (N_5506,N_2254,N_3340);
and U5507 (N_5507,N_3260,N_2462);
nand U5508 (N_5508,N_2530,N_3696);
or U5509 (N_5509,N_3801,N_2660);
nor U5510 (N_5510,N_2620,N_2494);
nand U5511 (N_5511,N_3905,N_3977);
nand U5512 (N_5512,N_3898,N_2809);
or U5513 (N_5513,N_3565,N_2683);
or U5514 (N_5514,N_3044,N_3021);
or U5515 (N_5515,N_3792,N_3389);
or U5516 (N_5516,N_2526,N_3697);
nand U5517 (N_5517,N_3176,N_3608);
nor U5518 (N_5518,N_3041,N_2445);
nand U5519 (N_5519,N_2912,N_3254);
nor U5520 (N_5520,N_2883,N_2081);
and U5521 (N_5521,N_2238,N_3727);
or U5522 (N_5522,N_3924,N_2085);
nand U5523 (N_5523,N_3356,N_2358);
nand U5524 (N_5524,N_2363,N_2643);
nand U5525 (N_5525,N_2274,N_3727);
nor U5526 (N_5526,N_2451,N_3321);
nor U5527 (N_5527,N_3555,N_3176);
xnor U5528 (N_5528,N_2706,N_2856);
xor U5529 (N_5529,N_2425,N_3069);
and U5530 (N_5530,N_3704,N_2080);
nand U5531 (N_5531,N_3926,N_3142);
and U5532 (N_5532,N_2390,N_3184);
or U5533 (N_5533,N_2468,N_2600);
or U5534 (N_5534,N_3211,N_2244);
nand U5535 (N_5535,N_2498,N_3819);
and U5536 (N_5536,N_2834,N_3871);
and U5537 (N_5537,N_3772,N_2522);
nor U5538 (N_5538,N_3729,N_2352);
nand U5539 (N_5539,N_2702,N_3689);
nor U5540 (N_5540,N_3679,N_2321);
nand U5541 (N_5541,N_2324,N_2299);
nor U5542 (N_5542,N_3344,N_3273);
or U5543 (N_5543,N_3653,N_2456);
nand U5544 (N_5544,N_2178,N_2171);
nor U5545 (N_5545,N_2892,N_2719);
or U5546 (N_5546,N_3338,N_3854);
or U5547 (N_5547,N_3296,N_3832);
nor U5548 (N_5548,N_3206,N_2082);
nor U5549 (N_5549,N_2015,N_2089);
or U5550 (N_5550,N_2917,N_2103);
or U5551 (N_5551,N_3429,N_3620);
nand U5552 (N_5552,N_2022,N_3702);
or U5553 (N_5553,N_3296,N_2876);
and U5554 (N_5554,N_2720,N_3105);
nor U5555 (N_5555,N_3298,N_3170);
nand U5556 (N_5556,N_3334,N_3939);
xor U5557 (N_5557,N_2486,N_2119);
and U5558 (N_5558,N_3906,N_3612);
nor U5559 (N_5559,N_2565,N_3873);
nor U5560 (N_5560,N_2245,N_2526);
nor U5561 (N_5561,N_2174,N_3250);
nor U5562 (N_5562,N_3833,N_3400);
and U5563 (N_5563,N_3748,N_3564);
or U5564 (N_5564,N_3900,N_3951);
xnor U5565 (N_5565,N_3448,N_3774);
nand U5566 (N_5566,N_2152,N_3757);
and U5567 (N_5567,N_3905,N_2923);
nor U5568 (N_5568,N_3779,N_2920);
and U5569 (N_5569,N_2699,N_3788);
nor U5570 (N_5570,N_3491,N_3660);
nand U5571 (N_5571,N_3270,N_2391);
nor U5572 (N_5572,N_2877,N_3239);
nor U5573 (N_5573,N_3654,N_3544);
nand U5574 (N_5574,N_2279,N_3764);
or U5575 (N_5575,N_2679,N_3400);
or U5576 (N_5576,N_2594,N_3399);
nand U5577 (N_5577,N_2052,N_3887);
xor U5578 (N_5578,N_3022,N_3397);
nor U5579 (N_5579,N_2369,N_3095);
and U5580 (N_5580,N_3985,N_2629);
nor U5581 (N_5581,N_2133,N_2438);
or U5582 (N_5582,N_3545,N_3829);
nand U5583 (N_5583,N_2493,N_3103);
nand U5584 (N_5584,N_3670,N_2253);
nand U5585 (N_5585,N_3252,N_3301);
nand U5586 (N_5586,N_2188,N_3580);
and U5587 (N_5587,N_3372,N_3072);
and U5588 (N_5588,N_3088,N_3507);
nand U5589 (N_5589,N_3807,N_3254);
and U5590 (N_5590,N_2232,N_3877);
nor U5591 (N_5591,N_2827,N_3827);
nor U5592 (N_5592,N_2922,N_3878);
nor U5593 (N_5593,N_3104,N_2332);
nor U5594 (N_5594,N_2243,N_3490);
nor U5595 (N_5595,N_3126,N_3591);
or U5596 (N_5596,N_2166,N_3556);
or U5597 (N_5597,N_2747,N_2047);
or U5598 (N_5598,N_3030,N_2688);
and U5599 (N_5599,N_2868,N_2020);
nand U5600 (N_5600,N_2207,N_3701);
nor U5601 (N_5601,N_2490,N_3410);
and U5602 (N_5602,N_2369,N_2717);
nor U5603 (N_5603,N_2019,N_2458);
nor U5604 (N_5604,N_2069,N_2336);
and U5605 (N_5605,N_3566,N_3799);
nor U5606 (N_5606,N_2545,N_3337);
nor U5607 (N_5607,N_3902,N_2346);
xor U5608 (N_5608,N_2265,N_3310);
nand U5609 (N_5609,N_3168,N_2107);
and U5610 (N_5610,N_2127,N_2524);
or U5611 (N_5611,N_2687,N_3443);
or U5612 (N_5612,N_3397,N_3506);
and U5613 (N_5613,N_2947,N_2140);
nor U5614 (N_5614,N_3676,N_2169);
or U5615 (N_5615,N_3822,N_3249);
or U5616 (N_5616,N_3956,N_2750);
or U5617 (N_5617,N_2431,N_2300);
nor U5618 (N_5618,N_3894,N_3090);
and U5619 (N_5619,N_2231,N_3843);
nand U5620 (N_5620,N_3693,N_2336);
or U5621 (N_5621,N_2901,N_3036);
or U5622 (N_5622,N_2086,N_3218);
nand U5623 (N_5623,N_2929,N_3221);
and U5624 (N_5624,N_2251,N_2180);
nand U5625 (N_5625,N_2621,N_3366);
nor U5626 (N_5626,N_2686,N_2569);
nand U5627 (N_5627,N_2985,N_2769);
and U5628 (N_5628,N_2179,N_3757);
and U5629 (N_5629,N_3698,N_2110);
nor U5630 (N_5630,N_2962,N_2306);
nand U5631 (N_5631,N_2882,N_3508);
and U5632 (N_5632,N_2935,N_2054);
and U5633 (N_5633,N_3088,N_3524);
and U5634 (N_5634,N_3526,N_2061);
nor U5635 (N_5635,N_2247,N_2121);
nand U5636 (N_5636,N_2045,N_3912);
or U5637 (N_5637,N_2075,N_2168);
xnor U5638 (N_5638,N_3481,N_3824);
and U5639 (N_5639,N_3614,N_2991);
and U5640 (N_5640,N_2628,N_2165);
and U5641 (N_5641,N_3748,N_2043);
nor U5642 (N_5642,N_2132,N_3231);
nor U5643 (N_5643,N_2147,N_2214);
nor U5644 (N_5644,N_2284,N_3708);
and U5645 (N_5645,N_3568,N_3169);
nor U5646 (N_5646,N_3932,N_3211);
and U5647 (N_5647,N_2395,N_2765);
nor U5648 (N_5648,N_2394,N_3985);
nand U5649 (N_5649,N_2436,N_2599);
and U5650 (N_5650,N_3800,N_3888);
or U5651 (N_5651,N_2071,N_2543);
or U5652 (N_5652,N_3595,N_2006);
nor U5653 (N_5653,N_3990,N_3001);
nand U5654 (N_5654,N_2451,N_3675);
nor U5655 (N_5655,N_2339,N_2183);
and U5656 (N_5656,N_3162,N_2797);
nor U5657 (N_5657,N_3359,N_3959);
and U5658 (N_5658,N_3237,N_2941);
nand U5659 (N_5659,N_3643,N_2425);
nor U5660 (N_5660,N_2099,N_2640);
nor U5661 (N_5661,N_2073,N_3054);
or U5662 (N_5662,N_3286,N_3367);
or U5663 (N_5663,N_2469,N_2132);
nor U5664 (N_5664,N_3969,N_2791);
and U5665 (N_5665,N_3761,N_3781);
or U5666 (N_5666,N_2319,N_2809);
or U5667 (N_5667,N_2546,N_3267);
nor U5668 (N_5668,N_3442,N_3693);
nand U5669 (N_5669,N_2935,N_2607);
or U5670 (N_5670,N_2713,N_3677);
nor U5671 (N_5671,N_3924,N_2038);
or U5672 (N_5672,N_3121,N_2642);
nor U5673 (N_5673,N_2859,N_2927);
nor U5674 (N_5674,N_2864,N_2266);
and U5675 (N_5675,N_2299,N_3630);
and U5676 (N_5676,N_3524,N_3872);
nor U5677 (N_5677,N_3762,N_2159);
nor U5678 (N_5678,N_3093,N_3606);
and U5679 (N_5679,N_2365,N_2816);
nand U5680 (N_5680,N_3261,N_2899);
nor U5681 (N_5681,N_2608,N_2007);
or U5682 (N_5682,N_3130,N_3918);
nand U5683 (N_5683,N_3748,N_2022);
or U5684 (N_5684,N_3352,N_2827);
or U5685 (N_5685,N_2414,N_2463);
and U5686 (N_5686,N_3393,N_2861);
nand U5687 (N_5687,N_3494,N_2324);
or U5688 (N_5688,N_2680,N_2297);
or U5689 (N_5689,N_2252,N_3469);
nor U5690 (N_5690,N_3227,N_2890);
nand U5691 (N_5691,N_2209,N_2194);
or U5692 (N_5692,N_2082,N_3481);
or U5693 (N_5693,N_2970,N_2978);
nor U5694 (N_5694,N_2136,N_3899);
nor U5695 (N_5695,N_3085,N_2914);
or U5696 (N_5696,N_3041,N_3045);
nor U5697 (N_5697,N_2023,N_2957);
nand U5698 (N_5698,N_2062,N_3845);
or U5699 (N_5699,N_2385,N_3344);
nand U5700 (N_5700,N_3767,N_2413);
nand U5701 (N_5701,N_3348,N_2611);
nand U5702 (N_5702,N_3710,N_2538);
or U5703 (N_5703,N_3770,N_3074);
nand U5704 (N_5704,N_3449,N_3523);
or U5705 (N_5705,N_3532,N_2410);
nand U5706 (N_5706,N_3020,N_3714);
nand U5707 (N_5707,N_2206,N_2478);
or U5708 (N_5708,N_3082,N_3390);
nand U5709 (N_5709,N_2453,N_2680);
and U5710 (N_5710,N_3786,N_3535);
nand U5711 (N_5711,N_2524,N_2999);
and U5712 (N_5712,N_3450,N_3949);
and U5713 (N_5713,N_3718,N_3772);
and U5714 (N_5714,N_2535,N_2669);
nor U5715 (N_5715,N_3770,N_2859);
nor U5716 (N_5716,N_3934,N_3930);
nand U5717 (N_5717,N_3706,N_2847);
nand U5718 (N_5718,N_2028,N_2774);
or U5719 (N_5719,N_2919,N_2703);
nand U5720 (N_5720,N_3581,N_3404);
nor U5721 (N_5721,N_3560,N_3960);
nor U5722 (N_5722,N_3791,N_3161);
nand U5723 (N_5723,N_3198,N_3674);
nor U5724 (N_5724,N_2919,N_3650);
nand U5725 (N_5725,N_3629,N_3454);
or U5726 (N_5726,N_3034,N_3342);
and U5727 (N_5727,N_2915,N_3127);
nand U5728 (N_5728,N_2631,N_3406);
and U5729 (N_5729,N_3485,N_3373);
nand U5730 (N_5730,N_2544,N_2721);
and U5731 (N_5731,N_2025,N_2272);
and U5732 (N_5732,N_3189,N_2788);
nand U5733 (N_5733,N_3547,N_2787);
or U5734 (N_5734,N_3491,N_2579);
nand U5735 (N_5735,N_2620,N_3583);
and U5736 (N_5736,N_2707,N_3737);
and U5737 (N_5737,N_3912,N_2983);
nand U5738 (N_5738,N_2555,N_2387);
nand U5739 (N_5739,N_3737,N_3012);
nor U5740 (N_5740,N_2399,N_2606);
and U5741 (N_5741,N_2584,N_3230);
and U5742 (N_5742,N_3983,N_2429);
nor U5743 (N_5743,N_3238,N_3599);
nor U5744 (N_5744,N_2331,N_3677);
nand U5745 (N_5745,N_3154,N_2873);
nand U5746 (N_5746,N_2819,N_2995);
nor U5747 (N_5747,N_2517,N_3484);
and U5748 (N_5748,N_3323,N_2231);
and U5749 (N_5749,N_2502,N_3854);
or U5750 (N_5750,N_3068,N_2450);
nand U5751 (N_5751,N_2897,N_3274);
or U5752 (N_5752,N_3037,N_2164);
nand U5753 (N_5753,N_2948,N_3123);
nand U5754 (N_5754,N_3155,N_2677);
or U5755 (N_5755,N_2650,N_3302);
nand U5756 (N_5756,N_2987,N_3206);
or U5757 (N_5757,N_3243,N_3559);
and U5758 (N_5758,N_2309,N_3250);
and U5759 (N_5759,N_3381,N_2318);
nand U5760 (N_5760,N_2627,N_3571);
and U5761 (N_5761,N_3553,N_3896);
or U5762 (N_5762,N_3479,N_3455);
and U5763 (N_5763,N_2849,N_3707);
xnor U5764 (N_5764,N_3173,N_3113);
nor U5765 (N_5765,N_2623,N_3199);
nor U5766 (N_5766,N_3422,N_3072);
nor U5767 (N_5767,N_2194,N_2885);
xor U5768 (N_5768,N_2641,N_2610);
nor U5769 (N_5769,N_3214,N_3056);
and U5770 (N_5770,N_2721,N_2011);
xor U5771 (N_5771,N_2751,N_3767);
nor U5772 (N_5772,N_2585,N_2092);
xnor U5773 (N_5773,N_3186,N_3501);
or U5774 (N_5774,N_2552,N_3567);
and U5775 (N_5775,N_2080,N_2516);
and U5776 (N_5776,N_3802,N_2375);
xnor U5777 (N_5777,N_2584,N_3488);
nand U5778 (N_5778,N_3703,N_2214);
nor U5779 (N_5779,N_3025,N_3193);
nor U5780 (N_5780,N_2746,N_2788);
or U5781 (N_5781,N_3566,N_2115);
nor U5782 (N_5782,N_3501,N_2284);
or U5783 (N_5783,N_3085,N_3561);
and U5784 (N_5784,N_2674,N_3149);
nor U5785 (N_5785,N_3118,N_2658);
or U5786 (N_5786,N_2596,N_2647);
nor U5787 (N_5787,N_3698,N_3949);
nand U5788 (N_5788,N_3845,N_3974);
nand U5789 (N_5789,N_3341,N_3247);
or U5790 (N_5790,N_3343,N_3679);
and U5791 (N_5791,N_2912,N_2241);
and U5792 (N_5792,N_3124,N_3742);
and U5793 (N_5793,N_2972,N_3175);
nand U5794 (N_5794,N_3362,N_2594);
nand U5795 (N_5795,N_3403,N_3864);
nand U5796 (N_5796,N_3586,N_3173);
and U5797 (N_5797,N_3340,N_3581);
nor U5798 (N_5798,N_2645,N_3576);
nand U5799 (N_5799,N_3959,N_3918);
or U5800 (N_5800,N_2297,N_3720);
and U5801 (N_5801,N_2649,N_2768);
and U5802 (N_5802,N_3605,N_2141);
or U5803 (N_5803,N_2128,N_3592);
nand U5804 (N_5804,N_3007,N_3965);
or U5805 (N_5805,N_3463,N_2508);
nand U5806 (N_5806,N_2457,N_3535);
nor U5807 (N_5807,N_3352,N_2415);
nor U5808 (N_5808,N_2816,N_3802);
and U5809 (N_5809,N_3148,N_3831);
and U5810 (N_5810,N_3856,N_2959);
and U5811 (N_5811,N_2121,N_2351);
nor U5812 (N_5812,N_3884,N_3692);
and U5813 (N_5813,N_2117,N_2493);
and U5814 (N_5814,N_2487,N_3674);
and U5815 (N_5815,N_3535,N_2571);
or U5816 (N_5816,N_3519,N_3008);
or U5817 (N_5817,N_3855,N_2124);
nor U5818 (N_5818,N_2261,N_3288);
and U5819 (N_5819,N_3129,N_3930);
nand U5820 (N_5820,N_3161,N_2580);
nor U5821 (N_5821,N_3418,N_3768);
nor U5822 (N_5822,N_3824,N_2792);
nand U5823 (N_5823,N_3069,N_2657);
nor U5824 (N_5824,N_3552,N_2790);
nand U5825 (N_5825,N_3109,N_2904);
nor U5826 (N_5826,N_3322,N_2167);
or U5827 (N_5827,N_2782,N_3130);
or U5828 (N_5828,N_3084,N_3592);
and U5829 (N_5829,N_2338,N_3962);
nor U5830 (N_5830,N_2876,N_2970);
nand U5831 (N_5831,N_2466,N_3079);
and U5832 (N_5832,N_3151,N_2783);
nor U5833 (N_5833,N_3039,N_3722);
nor U5834 (N_5834,N_3790,N_2592);
nand U5835 (N_5835,N_2147,N_3250);
and U5836 (N_5836,N_3204,N_3361);
and U5837 (N_5837,N_2030,N_2941);
and U5838 (N_5838,N_3490,N_3850);
or U5839 (N_5839,N_2139,N_2586);
nor U5840 (N_5840,N_2709,N_3571);
and U5841 (N_5841,N_3637,N_2654);
and U5842 (N_5842,N_2147,N_2450);
or U5843 (N_5843,N_2249,N_2472);
and U5844 (N_5844,N_3657,N_2229);
nand U5845 (N_5845,N_3666,N_2773);
and U5846 (N_5846,N_3738,N_3371);
nand U5847 (N_5847,N_3956,N_2155);
and U5848 (N_5848,N_3966,N_2337);
nand U5849 (N_5849,N_3371,N_2219);
nor U5850 (N_5850,N_2127,N_3156);
nor U5851 (N_5851,N_2137,N_3328);
or U5852 (N_5852,N_2080,N_2204);
or U5853 (N_5853,N_2837,N_2270);
or U5854 (N_5854,N_2588,N_2256);
or U5855 (N_5855,N_2860,N_3901);
nor U5856 (N_5856,N_3136,N_2687);
or U5857 (N_5857,N_2565,N_2788);
nor U5858 (N_5858,N_3429,N_2249);
nor U5859 (N_5859,N_2746,N_2879);
nand U5860 (N_5860,N_2358,N_2545);
or U5861 (N_5861,N_3236,N_2883);
or U5862 (N_5862,N_3033,N_3915);
nand U5863 (N_5863,N_3551,N_2305);
nor U5864 (N_5864,N_2168,N_2974);
nor U5865 (N_5865,N_3736,N_2898);
or U5866 (N_5866,N_3157,N_3324);
or U5867 (N_5867,N_2378,N_3518);
or U5868 (N_5868,N_3830,N_3664);
nor U5869 (N_5869,N_3347,N_3922);
or U5870 (N_5870,N_2996,N_2950);
or U5871 (N_5871,N_3483,N_3867);
nor U5872 (N_5872,N_2225,N_3039);
xor U5873 (N_5873,N_2028,N_3093);
or U5874 (N_5874,N_2168,N_2148);
nand U5875 (N_5875,N_2004,N_2561);
nor U5876 (N_5876,N_3010,N_2858);
and U5877 (N_5877,N_3108,N_3443);
and U5878 (N_5878,N_3452,N_3299);
and U5879 (N_5879,N_3253,N_2797);
nor U5880 (N_5880,N_3343,N_2348);
nand U5881 (N_5881,N_2587,N_2639);
nor U5882 (N_5882,N_2507,N_3715);
or U5883 (N_5883,N_2424,N_3388);
nand U5884 (N_5884,N_3960,N_3533);
nand U5885 (N_5885,N_2723,N_2182);
or U5886 (N_5886,N_3038,N_3461);
and U5887 (N_5887,N_2538,N_3846);
or U5888 (N_5888,N_3448,N_3898);
nand U5889 (N_5889,N_3847,N_3341);
nor U5890 (N_5890,N_3314,N_3477);
or U5891 (N_5891,N_2716,N_3480);
and U5892 (N_5892,N_2283,N_3574);
and U5893 (N_5893,N_2296,N_2398);
nor U5894 (N_5894,N_2777,N_3652);
or U5895 (N_5895,N_3062,N_2822);
nor U5896 (N_5896,N_2899,N_2143);
or U5897 (N_5897,N_2508,N_2970);
nand U5898 (N_5898,N_3633,N_2177);
or U5899 (N_5899,N_2314,N_3909);
nand U5900 (N_5900,N_2447,N_2936);
or U5901 (N_5901,N_2439,N_3134);
nand U5902 (N_5902,N_2160,N_3446);
nor U5903 (N_5903,N_3437,N_3448);
nor U5904 (N_5904,N_3201,N_2321);
and U5905 (N_5905,N_3708,N_2649);
nand U5906 (N_5906,N_3934,N_2558);
and U5907 (N_5907,N_2710,N_2985);
nor U5908 (N_5908,N_3090,N_3841);
and U5909 (N_5909,N_2426,N_3272);
nand U5910 (N_5910,N_3573,N_2082);
or U5911 (N_5911,N_2002,N_3152);
nand U5912 (N_5912,N_2887,N_2555);
or U5913 (N_5913,N_3491,N_2489);
or U5914 (N_5914,N_2058,N_3945);
nand U5915 (N_5915,N_2234,N_2595);
or U5916 (N_5916,N_3635,N_3730);
or U5917 (N_5917,N_3764,N_3312);
or U5918 (N_5918,N_3516,N_3599);
nor U5919 (N_5919,N_3240,N_2921);
nor U5920 (N_5920,N_2059,N_3628);
nand U5921 (N_5921,N_2976,N_2437);
nand U5922 (N_5922,N_2092,N_3147);
nor U5923 (N_5923,N_2865,N_2277);
or U5924 (N_5924,N_2006,N_2120);
nand U5925 (N_5925,N_3767,N_2262);
nor U5926 (N_5926,N_2967,N_2586);
nor U5927 (N_5927,N_3776,N_3702);
and U5928 (N_5928,N_2731,N_3250);
nand U5929 (N_5929,N_3828,N_2711);
or U5930 (N_5930,N_2874,N_2105);
nor U5931 (N_5931,N_3102,N_3042);
nor U5932 (N_5932,N_3872,N_3967);
or U5933 (N_5933,N_3925,N_3588);
and U5934 (N_5934,N_3907,N_3882);
nor U5935 (N_5935,N_2950,N_3658);
nor U5936 (N_5936,N_2506,N_3193);
and U5937 (N_5937,N_3000,N_2130);
and U5938 (N_5938,N_2888,N_2865);
nand U5939 (N_5939,N_2531,N_2142);
or U5940 (N_5940,N_3287,N_2572);
nor U5941 (N_5941,N_2587,N_2984);
or U5942 (N_5942,N_2571,N_2238);
nand U5943 (N_5943,N_2298,N_2413);
nor U5944 (N_5944,N_2235,N_3592);
and U5945 (N_5945,N_2502,N_3260);
or U5946 (N_5946,N_3872,N_2687);
and U5947 (N_5947,N_2580,N_2273);
nor U5948 (N_5948,N_2514,N_3549);
nand U5949 (N_5949,N_3017,N_2716);
nor U5950 (N_5950,N_3876,N_3544);
nand U5951 (N_5951,N_2151,N_3554);
and U5952 (N_5952,N_2373,N_2414);
nand U5953 (N_5953,N_3260,N_2389);
nand U5954 (N_5954,N_2532,N_3448);
nor U5955 (N_5955,N_2818,N_2711);
nor U5956 (N_5956,N_3763,N_2936);
nand U5957 (N_5957,N_3625,N_3721);
and U5958 (N_5958,N_2976,N_2904);
or U5959 (N_5959,N_3976,N_3136);
or U5960 (N_5960,N_3791,N_2788);
nor U5961 (N_5961,N_3812,N_2884);
nor U5962 (N_5962,N_3793,N_2360);
nand U5963 (N_5963,N_2902,N_2880);
or U5964 (N_5964,N_2655,N_2342);
or U5965 (N_5965,N_2656,N_3397);
and U5966 (N_5966,N_3177,N_2934);
and U5967 (N_5967,N_3305,N_2638);
nor U5968 (N_5968,N_3346,N_2350);
nor U5969 (N_5969,N_3540,N_2714);
nand U5970 (N_5970,N_3578,N_2483);
nor U5971 (N_5971,N_2737,N_2725);
and U5972 (N_5972,N_3969,N_3142);
nand U5973 (N_5973,N_2719,N_3880);
and U5974 (N_5974,N_3481,N_3845);
and U5975 (N_5975,N_2572,N_3619);
and U5976 (N_5976,N_2976,N_2684);
nand U5977 (N_5977,N_2286,N_3326);
xnor U5978 (N_5978,N_2255,N_3751);
nor U5979 (N_5979,N_2395,N_2227);
or U5980 (N_5980,N_3388,N_3881);
nor U5981 (N_5981,N_2672,N_2068);
or U5982 (N_5982,N_2549,N_2271);
or U5983 (N_5983,N_2906,N_2997);
nand U5984 (N_5984,N_3600,N_3358);
nor U5985 (N_5985,N_2013,N_2744);
nor U5986 (N_5986,N_3612,N_3463);
or U5987 (N_5987,N_2319,N_2898);
nand U5988 (N_5988,N_2656,N_2837);
xor U5989 (N_5989,N_2415,N_3120);
and U5990 (N_5990,N_2853,N_3377);
nand U5991 (N_5991,N_3649,N_3845);
and U5992 (N_5992,N_3561,N_2320);
nand U5993 (N_5993,N_2046,N_2985);
and U5994 (N_5994,N_2046,N_3557);
nand U5995 (N_5995,N_3350,N_2246);
nand U5996 (N_5996,N_2026,N_2677);
and U5997 (N_5997,N_2447,N_2400);
and U5998 (N_5998,N_3903,N_2727);
and U5999 (N_5999,N_3706,N_3716);
nor U6000 (N_6000,N_4689,N_5352);
nor U6001 (N_6001,N_5479,N_4261);
xor U6002 (N_6002,N_5587,N_5768);
nand U6003 (N_6003,N_5298,N_5906);
or U6004 (N_6004,N_4072,N_4155);
or U6005 (N_6005,N_5880,N_4282);
nand U6006 (N_6006,N_4765,N_4991);
nor U6007 (N_6007,N_5738,N_5164);
or U6008 (N_6008,N_5868,N_5978);
nand U6009 (N_6009,N_5746,N_5771);
and U6010 (N_6010,N_4114,N_5297);
xnor U6011 (N_6011,N_5050,N_4253);
nand U6012 (N_6012,N_4853,N_5068);
xor U6013 (N_6013,N_4817,N_5147);
and U6014 (N_6014,N_5066,N_5913);
nor U6015 (N_6015,N_5843,N_5062);
or U6016 (N_6016,N_5891,N_4137);
nand U6017 (N_6017,N_4368,N_4482);
and U6018 (N_6018,N_4026,N_5079);
nand U6019 (N_6019,N_5275,N_5274);
nor U6020 (N_6020,N_4276,N_4949);
nand U6021 (N_6021,N_5284,N_4422);
nand U6022 (N_6022,N_4340,N_4663);
and U6023 (N_6023,N_5895,N_5128);
nor U6024 (N_6024,N_4372,N_5075);
nand U6025 (N_6025,N_4460,N_4289);
and U6026 (N_6026,N_4809,N_5134);
nor U6027 (N_6027,N_4147,N_5469);
or U6028 (N_6028,N_5825,N_4941);
xnor U6029 (N_6029,N_4583,N_4610);
nor U6030 (N_6030,N_5995,N_5010);
nor U6031 (N_6031,N_4619,N_4668);
or U6032 (N_6032,N_4326,N_5980);
nand U6033 (N_6033,N_5624,N_4281);
nor U6034 (N_6034,N_4077,N_4028);
nor U6035 (N_6035,N_4153,N_4358);
nor U6036 (N_6036,N_5862,N_4006);
nand U6037 (N_6037,N_4665,N_5860);
nand U6038 (N_6038,N_4628,N_4223);
nor U6039 (N_6039,N_5499,N_4366);
or U6040 (N_6040,N_5564,N_5721);
or U6041 (N_6041,N_5566,N_4964);
nand U6042 (N_6042,N_5626,N_4721);
nor U6043 (N_6043,N_5199,N_5729);
nor U6044 (N_6044,N_4037,N_4783);
nor U6045 (N_6045,N_4049,N_4922);
or U6046 (N_6046,N_4122,N_5679);
nor U6047 (N_6047,N_5249,N_5744);
nor U6048 (N_6048,N_4730,N_5311);
nor U6049 (N_6049,N_4321,N_4118);
nor U6050 (N_6050,N_4643,N_5046);
nor U6051 (N_6051,N_5665,N_5047);
nand U6052 (N_6052,N_5893,N_5750);
and U6053 (N_6053,N_4902,N_5481);
or U6054 (N_6054,N_5006,N_5956);
and U6055 (N_6055,N_4916,N_5095);
and U6056 (N_6056,N_4076,N_5151);
and U6057 (N_6057,N_4492,N_5556);
nor U6058 (N_6058,N_5139,N_4742);
nor U6059 (N_6059,N_4278,N_4279);
or U6060 (N_6060,N_5427,N_4310);
and U6061 (N_6061,N_4322,N_5533);
and U6062 (N_6062,N_4053,N_5247);
or U6063 (N_6063,N_5142,N_5178);
nand U6064 (N_6064,N_4557,N_5551);
nand U6065 (N_6065,N_5618,N_4824);
or U6066 (N_6066,N_5830,N_4320);
nor U6067 (N_6067,N_4085,N_5424);
nand U6068 (N_6068,N_5613,N_4869);
and U6069 (N_6069,N_5254,N_4953);
nor U6070 (N_6070,N_4345,N_5101);
or U6071 (N_6071,N_4263,N_5334);
or U6072 (N_6072,N_5214,N_4517);
nor U6073 (N_6073,N_4001,N_5033);
or U6074 (N_6074,N_4002,N_5100);
nor U6075 (N_6075,N_4044,N_4735);
or U6076 (N_6076,N_4558,N_4070);
nand U6077 (N_6077,N_4715,N_4398);
or U6078 (N_6078,N_4240,N_5790);
nor U6079 (N_6079,N_4304,N_5281);
or U6080 (N_6080,N_4490,N_5846);
nor U6081 (N_6081,N_4083,N_5554);
nor U6082 (N_6082,N_5748,N_4633);
nor U6083 (N_6083,N_4519,N_5408);
nand U6084 (N_6084,N_5337,N_5097);
and U6085 (N_6085,N_5674,N_4502);
and U6086 (N_6086,N_4720,N_4277);
and U6087 (N_6087,N_5719,N_4898);
and U6088 (N_6088,N_4795,N_4974);
xor U6089 (N_6089,N_4461,N_4634);
and U6090 (N_6090,N_5837,N_4328);
or U6091 (N_6091,N_4976,N_5728);
and U6092 (N_6092,N_4872,N_5295);
and U6093 (N_6093,N_4283,N_4676);
or U6094 (N_6094,N_5967,N_4248);
or U6095 (N_6095,N_4254,N_4882);
nor U6096 (N_6096,N_4702,N_5011);
and U6097 (N_6097,N_5042,N_4651);
nand U6098 (N_6098,N_5316,N_4164);
nand U6099 (N_6099,N_4787,N_5030);
xnor U6100 (N_6100,N_5203,N_5970);
or U6101 (N_6101,N_5892,N_4190);
nand U6102 (N_6102,N_4704,N_4833);
or U6103 (N_6103,N_5712,N_5440);
and U6104 (N_6104,N_5794,N_5362);
nor U6105 (N_6105,N_4325,N_5890);
xor U6106 (N_6106,N_5781,N_5402);
nor U6107 (N_6107,N_4291,N_4488);
and U6108 (N_6108,N_4394,N_4412);
nand U6109 (N_6109,N_5930,N_4200);
nand U6110 (N_6110,N_4951,N_5081);
and U6111 (N_6111,N_5475,N_5185);
nand U6112 (N_6112,N_5458,N_4745);
nor U6113 (N_6113,N_4140,N_4221);
xnor U6114 (N_6114,N_5834,N_4313);
and U6115 (N_6115,N_4611,N_4561);
nor U6116 (N_6116,N_5384,N_5253);
and U6117 (N_6117,N_5375,N_5169);
and U6118 (N_6118,N_5951,N_4181);
or U6119 (N_6119,N_5317,N_5314);
and U6120 (N_6120,N_4736,N_4764);
nor U6121 (N_6121,N_5355,N_5289);
nand U6122 (N_6122,N_4088,N_4798);
and U6123 (N_6123,N_5398,N_5617);
nor U6124 (N_6124,N_4970,N_5597);
and U6125 (N_6125,N_5426,N_5823);
nand U6126 (N_6126,N_4523,N_5112);
or U6127 (N_6127,N_4808,N_4344);
or U6128 (N_6128,N_5174,N_5545);
or U6129 (N_6129,N_4184,N_5129);
and U6130 (N_6130,N_5360,N_4560);
xor U6131 (N_6131,N_5237,N_4891);
nor U6132 (N_6132,N_4593,N_5325);
nor U6133 (N_6133,N_4862,N_4713);
or U6134 (N_6134,N_5236,N_4161);
or U6135 (N_6135,N_4312,N_5826);
or U6136 (N_6136,N_5664,N_5783);
nand U6137 (N_6137,N_5461,N_5922);
nand U6138 (N_6138,N_5711,N_4052);
or U6139 (N_6139,N_4838,N_5245);
nor U6140 (N_6140,N_4511,N_5114);
or U6141 (N_6141,N_5537,N_4971);
nand U6142 (N_6142,N_5944,N_5938);
or U6143 (N_6143,N_5848,N_5818);
or U6144 (N_6144,N_5889,N_4477);
nand U6145 (N_6145,N_4933,N_5421);
nor U6146 (N_6146,N_5641,N_4618);
or U6147 (N_6147,N_5077,N_4471);
or U6148 (N_6148,N_5012,N_4078);
and U6149 (N_6149,N_4532,N_4251);
nor U6150 (N_6150,N_5961,N_4057);
nor U6151 (N_6151,N_5584,N_5255);
or U6152 (N_6152,N_4586,N_4255);
nor U6153 (N_6153,N_4566,N_4400);
nor U6154 (N_6154,N_4995,N_5542);
nor U6155 (N_6155,N_4396,N_5588);
or U6156 (N_6156,N_5294,N_5125);
nor U6157 (N_6157,N_4660,N_4166);
nor U6158 (N_6158,N_5779,N_5263);
and U6159 (N_6159,N_4359,N_5106);
nand U6160 (N_6160,N_5299,N_4635);
nand U6161 (N_6161,N_5108,N_4793);
nand U6162 (N_6162,N_5739,N_5753);
and U6163 (N_6163,N_4827,N_5092);
nand U6164 (N_6164,N_5899,N_5170);
nor U6165 (N_6165,N_5792,N_4367);
and U6166 (N_6166,N_4480,N_4260);
nor U6167 (N_6167,N_5700,N_4639);
nor U6168 (N_6168,N_5844,N_5265);
and U6169 (N_6169,N_5069,N_4187);
nor U6170 (N_6170,N_5900,N_5976);
nand U6171 (N_6171,N_4284,N_5954);
nor U6172 (N_6172,N_5221,N_5871);
nand U6173 (N_6173,N_5639,N_4733);
nand U6174 (N_6174,N_5549,N_5935);
xor U6175 (N_6175,N_5575,N_4644);
nand U6176 (N_6176,N_5642,N_4840);
or U6177 (N_6177,N_5619,N_5698);
and U6178 (N_6178,N_5160,N_4476);
and U6179 (N_6179,N_5583,N_5115);
nor U6180 (N_6180,N_4516,N_5686);
nor U6181 (N_6181,N_4638,N_5672);
nor U6182 (N_6182,N_5945,N_4024);
or U6183 (N_6183,N_4867,N_4352);
and U6184 (N_6184,N_5990,N_5749);
nand U6185 (N_6185,N_4604,N_4701);
and U6186 (N_6186,N_4636,N_5804);
nor U6187 (N_6187,N_4992,N_5801);
and U6188 (N_6188,N_4485,N_5787);
or U6189 (N_6189,N_4655,N_5416);
or U6190 (N_6190,N_5725,N_4996);
nand U6191 (N_6191,N_4861,N_5778);
nor U6192 (N_6192,N_5212,N_5262);
nand U6193 (N_6193,N_4152,N_5677);
or U6194 (N_6194,N_4499,N_5697);
or U6195 (N_6195,N_4430,N_5020);
and U6196 (N_6196,N_4960,N_4339);
nor U6197 (N_6197,N_4959,N_4129);
or U6198 (N_6198,N_5336,N_4469);
xor U6199 (N_6199,N_5490,N_4497);
nor U6200 (N_6200,N_4401,N_5330);
and U6201 (N_6201,N_4271,N_4703);
nor U6202 (N_6202,N_4439,N_4998);
nand U6203 (N_6203,N_4710,N_5383);
nand U6204 (N_6204,N_4132,N_4524);
or U6205 (N_6205,N_5466,N_5213);
and U6206 (N_6206,N_4780,N_4238);
and U6207 (N_6207,N_5835,N_5879);
nand U6208 (N_6208,N_4921,N_5229);
or U6209 (N_6209,N_4536,N_5634);
nor U6210 (N_6210,N_5401,N_5026);
nor U6211 (N_6211,N_5869,N_4097);
nand U6212 (N_6212,N_4946,N_4102);
or U6213 (N_6213,N_5996,N_4025);
nor U6214 (N_6214,N_5407,N_5159);
nand U6215 (N_6215,N_5232,N_4364);
nor U6216 (N_6216,N_4059,N_4937);
and U6217 (N_6217,N_4802,N_5085);
nand U6218 (N_6218,N_5633,N_4311);
or U6219 (N_6219,N_4338,N_5054);
or U6220 (N_6220,N_4257,N_5016);
nor U6221 (N_6221,N_4903,N_5751);
or U6222 (N_6222,N_5378,N_5430);
nand U6223 (N_6223,N_5509,N_4819);
nor U6224 (N_6224,N_4332,N_5349);
nand U6225 (N_6225,N_5167,N_4148);
or U6226 (N_6226,N_5207,N_4815);
or U6227 (N_6227,N_4465,N_5568);
nand U6228 (N_6228,N_4901,N_5810);
xnor U6229 (N_6229,N_4160,N_5189);
or U6230 (N_6230,N_4656,N_4087);
nor U6231 (N_6231,N_4231,N_4151);
nand U6232 (N_6232,N_4983,N_4390);
nand U6233 (N_6233,N_5567,N_5272);
nand U6234 (N_6234,N_4080,N_5260);
and U6235 (N_6235,N_4066,N_5496);
and U6236 (N_6236,N_4444,N_4419);
nor U6237 (N_6237,N_5582,N_4011);
or U6238 (N_6238,N_4407,N_4455);
nor U6239 (N_6239,N_4095,N_4408);
nand U6240 (N_6240,N_4353,N_4875);
and U6241 (N_6241,N_5380,N_5560);
and U6242 (N_6242,N_5504,N_4449);
and U6243 (N_6243,N_5194,N_5492);
and U6244 (N_6244,N_5870,N_5840);
nand U6245 (N_6245,N_5215,N_4567);
nand U6246 (N_6246,N_4319,N_4177);
nand U6247 (N_6247,N_5415,N_5453);
or U6248 (N_6248,N_5720,N_4810);
or U6249 (N_6249,N_5628,N_5821);
and U6250 (N_6250,N_5409,N_5960);
and U6251 (N_6251,N_5552,N_4448);
or U6252 (N_6252,N_4870,N_4569);
or U6253 (N_6253,N_4487,N_5503);
and U6254 (N_6254,N_4171,N_4324);
nor U6255 (N_6255,N_4725,N_4625);
and U6256 (N_6256,N_4513,N_5484);
or U6257 (N_6257,N_5113,N_4700);
nor U6258 (N_6258,N_4664,N_4299);
nor U6259 (N_6259,N_5493,N_5894);
and U6260 (N_6260,N_5173,N_4414);
or U6261 (N_6261,N_4669,N_4609);
and U6262 (N_6262,N_4969,N_5709);
nor U6263 (N_6263,N_5457,N_5593);
nand U6264 (N_6264,N_4416,N_4197);
and U6265 (N_6265,N_5168,N_4373);
and U6266 (N_6266,N_5553,N_5116);
nor U6267 (N_6267,N_4159,N_4622);
and U6268 (N_6268,N_4799,N_4268);
and U6269 (N_6269,N_4172,N_5904);
nor U6270 (N_6270,N_4705,N_5800);
nor U6271 (N_6271,N_4017,N_5391);
or U6272 (N_6272,N_5514,N_5535);
and U6273 (N_6273,N_4968,N_4357);
nand U6274 (N_6274,N_5799,N_5694);
nor U6275 (N_6275,N_5266,N_4686);
nand U6276 (N_6276,N_4650,N_4866);
nor U6277 (N_6277,N_4158,N_5572);
or U6278 (N_6278,N_5126,N_4760);
nor U6279 (N_6279,N_5943,N_4904);
nand U6280 (N_6280,N_5495,N_4242);
and U6281 (N_6281,N_5940,N_4722);
xor U6282 (N_6282,N_4606,N_4966);
and U6283 (N_6283,N_5162,N_5140);
or U6284 (N_6284,N_4014,N_4089);
or U6285 (N_6285,N_4099,N_4112);
or U6286 (N_6286,N_4298,N_4588);
and U6287 (N_6287,N_4379,N_5186);
nor U6288 (N_6288,N_5205,N_4047);
nand U6289 (N_6289,N_4443,N_4712);
and U6290 (N_6290,N_4040,N_4830);
nor U6291 (N_6291,N_4426,N_4348);
nor U6292 (N_6292,N_4616,N_4589);
nor U6293 (N_6293,N_4544,N_5538);
nand U6294 (N_6294,N_5444,N_5797);
nor U6295 (N_6295,N_4503,N_4518);
and U6296 (N_6296,N_5141,N_4962);
or U6297 (N_6297,N_4865,N_4687);
xor U6298 (N_6298,N_5513,N_4377);
and U6299 (N_6299,N_4647,N_4111);
and U6300 (N_6300,N_4822,N_4335);
and U6301 (N_6301,N_5936,N_4192);
and U6302 (N_6302,N_4308,N_5635);
and U6303 (N_6303,N_5524,N_4521);
nor U6304 (N_6304,N_4498,N_4881);
or U6305 (N_6305,N_4842,N_4342);
and U6306 (N_6306,N_5812,N_4065);
or U6307 (N_6307,N_5534,N_5888);
nor U6308 (N_6308,N_5293,N_5002);
nand U6309 (N_6309,N_5576,N_5630);
nand U6310 (N_6310,N_4627,N_5571);
xor U6311 (N_6311,N_4209,N_5903);
or U6312 (N_6312,N_5515,N_4489);
xor U6313 (N_6313,N_5404,N_4229);
nand U6314 (N_6314,N_5829,N_5283);
nand U6315 (N_6315,N_4243,N_5569);
nor U6316 (N_6316,N_4900,N_4117);
and U6317 (N_6317,N_4621,N_5600);
and U6318 (N_6318,N_5578,N_5122);
or U6319 (N_6319,N_5278,N_5765);
nand U6320 (N_6320,N_5905,N_5096);
xnor U6321 (N_6321,N_5580,N_4370);
and U6322 (N_6322,N_5696,N_5347);
nor U6323 (N_6323,N_4110,N_5898);
nand U6324 (N_6324,N_5007,N_5972);
nand U6325 (N_6325,N_4403,N_5761);
and U6326 (N_6326,N_4559,N_5745);
and U6327 (N_6327,N_5034,N_4846);
and U6328 (N_6328,N_4692,N_5226);
or U6329 (N_6329,N_5695,N_5726);
or U6330 (N_6330,N_4607,N_5357);
and U6331 (N_6331,N_5171,N_4546);
nor U6332 (N_6332,N_5684,N_4574);
xor U6333 (N_6333,N_5094,N_5754);
or U6334 (N_6334,N_4661,N_4673);
or U6335 (N_6335,N_5279,N_5109);
or U6336 (N_6336,N_4758,N_4036);
nand U6337 (N_6337,N_5915,N_5267);
or U6338 (N_6338,N_4956,N_4107);
and U6339 (N_6339,N_4415,N_4170);
nand U6340 (N_6340,N_5521,N_5445);
nand U6341 (N_6341,N_5923,N_5747);
nand U6342 (N_6342,N_4150,N_5187);
nor U6343 (N_6343,N_5759,N_5965);
or U6344 (N_6344,N_5682,N_4167);
or U6345 (N_6345,N_4273,N_4314);
or U6346 (N_6346,N_5723,N_5688);
or U6347 (N_6347,N_4051,N_5574);
or U6348 (N_6348,N_5654,N_5313);
nand U6349 (N_6349,N_4943,N_5252);
or U6350 (N_6350,N_4806,N_5992);
nand U6351 (N_6351,N_4580,N_5015);
nor U6352 (N_6352,N_4775,N_5873);
nor U6353 (N_6353,N_5350,N_4759);
and U6354 (N_6354,N_5839,N_5381);
or U6355 (N_6355,N_4475,N_5372);
nand U6356 (N_6356,N_5942,N_4022);
nor U6357 (N_6357,N_5482,N_5780);
nor U6358 (N_6358,N_4041,N_5502);
and U6359 (N_6359,N_4029,N_5671);
nand U6360 (N_6360,N_4878,N_5271);
nand U6361 (N_6361,N_4895,N_4463);
nand U6362 (N_6362,N_4256,N_4965);
nand U6363 (N_6363,N_5373,N_5211);
and U6364 (N_6364,N_5086,N_5256);
nor U6365 (N_6365,N_5603,N_5285);
and U6366 (N_6366,N_5103,N_5713);
nor U6367 (N_6367,N_4706,N_4681);
xnor U6368 (N_6368,N_5452,N_5808);
nand U6369 (N_6369,N_5339,N_4108);
or U6370 (N_6370,N_5543,N_5158);
or U6371 (N_6371,N_5208,N_4437);
or U6372 (N_6372,N_4854,N_5831);
nor U6373 (N_6373,N_5699,N_5602);
or U6374 (N_6374,N_4615,N_4063);
and U6375 (N_6375,N_4990,N_5459);
nor U6376 (N_6376,N_4441,N_4896);
and U6377 (N_6377,N_4270,N_4678);
or U6378 (N_6378,N_5581,N_4241);
or U6379 (N_6379,N_4138,N_4402);
and U6380 (N_6380,N_4309,N_5433);
nor U6381 (N_6381,N_5150,N_5966);
or U6382 (N_6382,N_5019,N_4329);
xnor U6383 (N_6383,N_5436,N_4507);
nor U6384 (N_6384,N_4740,N_5450);
or U6385 (N_6385,N_4863,N_4699);
nand U6386 (N_6386,N_4929,N_5438);
and U6387 (N_6387,N_4794,N_5412);
nand U6388 (N_6388,N_5622,N_5851);
nand U6389 (N_6389,N_4333,N_4462);
and U6390 (N_6390,N_5286,N_5083);
nand U6391 (N_6391,N_4130,N_4384);
nor U6392 (N_6392,N_4202,N_5760);
nor U6393 (N_6393,N_4982,N_5315);
nor U6394 (N_6394,N_4018,N_5276);
nand U6395 (N_6395,N_4905,N_4930);
nor U6396 (N_6396,N_5621,N_5001);
and U6397 (N_6397,N_4911,N_5854);
and U6398 (N_6398,N_5592,N_4330);
nand U6399 (N_6399,N_4143,N_4553);
or U6400 (N_6400,N_5737,N_5057);
or U6401 (N_6401,N_4142,N_4542);
and U6402 (N_6402,N_4010,N_4979);
or U6403 (N_6403,N_5058,N_5658);
nor U6404 (N_6404,N_5070,N_4456);
nor U6405 (N_6405,N_4316,N_4747);
nand U6406 (N_6406,N_4383,N_4071);
xnor U6407 (N_6407,N_4552,N_4781);
and U6408 (N_6408,N_5987,N_5045);
or U6409 (N_6409,N_5397,N_5740);
nand U6410 (N_6410,N_4512,N_5483);
or U6411 (N_6411,N_5153,N_4382);
nand U6412 (N_6412,N_4007,N_4572);
or U6413 (N_6413,N_5312,N_5183);
and U6414 (N_6414,N_5420,N_5933);
or U6415 (N_6415,N_4351,N_5418);
nand U6416 (N_6416,N_5912,N_4932);
nand U6417 (N_6417,N_5523,N_4756);
nor U6418 (N_6418,N_5735,N_5991);
or U6419 (N_6419,N_5156,N_5919);
and U6420 (N_6420,N_5501,N_5644);
nor U6421 (N_6421,N_5071,N_5157);
nor U6422 (N_6422,N_4514,N_4790);
and U6423 (N_6423,N_4494,N_5379);
nor U6424 (N_6424,N_5029,N_4942);
nand U6425 (N_6425,N_5117,N_4918);
and U6426 (N_6426,N_4405,N_4264);
or U6427 (N_6427,N_4191,N_5488);
nand U6428 (N_6428,N_5431,N_5329);
nor U6429 (N_6429,N_4834,N_5953);
nand U6430 (N_6430,N_4723,N_5202);
or U6431 (N_6431,N_5809,N_4886);
nand U6432 (N_6432,N_5702,N_4987);
and U6433 (N_6433,N_4816,N_5040);
or U6434 (N_6434,N_4442,N_5388);
or U6435 (N_6435,N_4534,N_4180);
nor U6436 (N_6436,N_5191,N_4409);
and U6437 (N_6437,N_4548,N_4975);
and U6438 (N_6438,N_4890,N_5827);
or U6439 (N_6439,N_4061,N_4563);
and U6440 (N_6440,N_5947,N_4562);
and U6441 (N_6441,N_4208,N_4594);
and U6442 (N_6442,N_4144,N_4436);
nor U6443 (N_6443,N_4565,N_4910);
nor U6444 (N_6444,N_4131,N_5031);
nand U6445 (N_6445,N_5724,N_4349);
nand U6446 (N_6446,N_4994,N_5758);
nor U6447 (N_6447,N_5764,N_5775);
and U6448 (N_6448,N_4856,N_4391);
nor U6449 (N_6449,N_5939,N_5985);
and U6450 (N_6450,N_4098,N_4365);
and U6451 (N_6451,N_5356,N_5914);
nand U6452 (N_6452,N_5610,N_4075);
or U6453 (N_6453,N_4295,N_4757);
or U6454 (N_6454,N_5774,N_4406);
nand U6455 (N_6455,N_5302,N_5973);
and U6456 (N_6456,N_4843,N_4526);
or U6457 (N_6457,N_4529,N_4288);
and U6458 (N_6458,N_5118,N_4323);
nor U6459 (N_6459,N_4149,N_5353);
nor U6460 (N_6460,N_5763,N_5235);
nor U6461 (N_6461,N_4694,N_4698);
or U6462 (N_6462,N_4535,N_4789);
or U6463 (N_6463,N_5354,N_5365);
nand U6464 (N_6464,N_5544,N_5419);
or U6465 (N_6465,N_4290,N_4667);
nand U6466 (N_6466,N_5161,N_4473);
or U6467 (N_6467,N_5948,N_4505);
or U6468 (N_6468,N_4459,N_5119);
and U6469 (N_6469,N_5795,N_4543);
or U6470 (N_6470,N_5258,N_5123);
xor U6471 (N_6471,N_5974,N_5901);
or U6472 (N_6472,N_5474,N_5741);
and U6473 (N_6473,N_5422,N_4198);
nand U6474 (N_6474,N_4128,N_5084);
nand U6475 (N_6475,N_4575,N_5144);
or U6476 (N_6476,N_4844,N_4234);
or U6477 (N_6477,N_5363,N_5705);
or U6478 (N_6478,N_4104,N_4350);
or U6479 (N_6479,N_5620,N_4027);
nor U6480 (N_6480,N_4893,N_5874);
or U6481 (N_6481,N_5511,N_4336);
or U6482 (N_6482,N_4274,N_5146);
or U6483 (N_6483,N_5089,N_4828);
nand U6484 (N_6484,N_4458,N_4550);
nand U6485 (N_6485,N_5099,N_5073);
nor U6486 (N_6486,N_4948,N_5977);
nor U6487 (N_6487,N_4989,N_4614);
and U6488 (N_6488,N_5661,N_4748);
nand U6489 (N_6489,N_5776,N_5926);
or U6490 (N_6490,N_4297,N_5210);
and U6491 (N_6491,N_5498,N_5701);
nand U6492 (N_6492,N_4666,N_5025);
nor U6493 (N_6493,N_5107,N_4785);
nor U6494 (N_6494,N_4680,N_5604);
and U6495 (N_6495,N_4988,N_4812);
nor U6496 (N_6496,N_4214,N_4906);
and U6497 (N_6497,N_4272,N_5847);
nor U6498 (N_6498,N_5324,N_5653);
nand U6499 (N_6499,N_5277,N_5656);
nand U6500 (N_6500,N_4168,N_4582);
nand U6501 (N_6501,N_4453,N_5074);
nand U6502 (N_6502,N_5303,N_5432);
nor U6503 (N_6503,N_5786,N_4094);
or U6504 (N_6504,N_5242,N_4042);
nand U6505 (N_6505,N_5652,N_4579);
nor U6506 (N_6506,N_4768,N_5730);
and U6507 (N_6507,N_4538,N_4204);
xnor U6508 (N_6508,N_5586,N_5590);
nand U6509 (N_6509,N_5282,N_5762);
or U6510 (N_6510,N_4058,N_5611);
or U6511 (N_6511,N_5038,N_4410);
nor U6512 (N_6512,N_5439,N_4750);
and U6513 (N_6513,N_5866,N_5093);
nand U6514 (N_6514,N_4504,N_5876);
and U6515 (N_6515,N_5451,N_5090);
or U6516 (N_6516,N_4245,N_4145);
or U6517 (N_6517,N_4262,N_4734);
and U6518 (N_6518,N_4048,N_5154);
and U6519 (N_6519,N_4924,N_4043);
and U6520 (N_6520,N_5908,N_4163);
nor U6521 (N_6521,N_5063,N_4731);
or U6522 (N_6522,N_4719,N_4774);
or U6523 (N_6523,N_5605,N_5929);
nor U6524 (N_6524,N_4860,N_5819);
nor U6525 (N_6525,N_4124,N_5342);
and U6526 (N_6526,N_4912,N_5660);
nand U6527 (N_6527,N_5878,N_4825);
or U6528 (N_6528,N_5640,N_4973);
nand U6529 (N_6529,N_4244,N_5013);
nand U6530 (N_6530,N_4954,N_4568);
and U6531 (N_6531,N_4707,N_4908);
nor U6532 (N_6532,N_5527,N_5941);
and U6533 (N_6533,N_5060,N_5039);
nor U6534 (N_6534,N_5952,N_5454);
or U6535 (N_6535,N_5305,N_4788);
nor U6536 (N_6536,N_5177,N_5756);
nor U6537 (N_6537,N_4624,N_5824);
nor U6538 (N_6538,N_4592,N_4226);
xor U6539 (N_6539,N_5842,N_4600);
and U6540 (N_6540,N_5984,N_5927);
nor U6541 (N_6541,N_4729,N_5670);
nor U6542 (N_6542,N_4837,N_5023);
nand U6543 (N_6543,N_5668,N_5536);
or U6544 (N_6544,N_5009,N_5770);
nor U6545 (N_6545,N_5924,N_4623);
and U6546 (N_6546,N_5198,N_4091);
nand U6547 (N_6547,N_4800,N_4845);
or U6548 (N_6548,N_5814,N_4716);
nand U6549 (N_6549,N_5707,N_5393);
nor U6550 (N_6550,N_5200,N_4892);
and U6551 (N_6551,N_5143,N_4986);
and U6552 (N_6552,N_4897,N_5884);
or U6553 (N_6553,N_4728,N_5184);
nor U6554 (N_6554,N_5338,N_5309);
nand U6555 (N_6555,N_4346,N_5322);
nand U6556 (N_6556,N_4763,N_5632);
or U6557 (N_6557,N_4228,N_4612);
or U6558 (N_6558,N_5838,N_4506);
nand U6559 (N_6559,N_5182,N_5000);
nor U6560 (N_6560,N_4779,N_5216);
or U6561 (N_6561,N_4564,N_5410);
and U6562 (N_6562,N_5949,N_5358);
nand U6563 (N_6563,N_5703,N_4105);
and U6564 (N_6564,N_4337,N_4033);
or U6565 (N_6565,N_5902,N_5963);
nand U6566 (N_6566,N_4595,N_4232);
nand U6567 (N_6567,N_4743,N_5999);
or U6568 (N_6568,N_4654,N_4907);
nand U6569 (N_6569,N_5772,N_5385);
or U6570 (N_6570,N_4302,N_4101);
nor U6571 (N_6571,N_4020,N_4019);
nor U6572 (N_6572,N_5348,N_5172);
xor U6573 (N_6573,N_4876,N_4139);
nand U6574 (N_6574,N_4090,N_5852);
nor U6575 (N_6575,N_4936,N_4885);
or U6576 (N_6576,N_5530,N_4826);
or U6577 (N_6577,N_4084,N_4103);
and U6578 (N_6578,N_4626,N_5449);
xor U6579 (N_6579,N_5218,N_4642);
nand U6580 (N_6580,N_4005,N_4212);
or U6581 (N_6581,N_4113,N_5371);
and U6582 (N_6582,N_4418,N_4420);
xor U6583 (N_6583,N_4913,N_4852);
nand U6584 (N_6584,N_4183,N_5364);
xor U6585 (N_6585,N_4481,N_4165);
and U6586 (N_6586,N_5120,N_5557);
nor U6587 (N_6587,N_4649,N_5691);
xnor U6588 (N_6588,N_4360,N_5918);
or U6589 (N_6589,N_4522,N_5246);
nand U6590 (N_6590,N_4193,N_5248);
and U6591 (N_6591,N_4958,N_4068);
nor U6592 (N_6592,N_4064,N_5230);
and U6593 (N_6593,N_5014,N_5647);
nand U6594 (N_6594,N_4280,N_4549);
and U6595 (N_6595,N_4591,N_4801);
xnor U6596 (N_6596,N_4726,N_4935);
or U6597 (N_6597,N_5021,N_5306);
and U6598 (N_6598,N_4275,N_4176);
nand U6599 (N_6599,N_5429,N_5163);
or U6600 (N_6600,N_4012,N_5845);
nor U6601 (N_6601,N_4467,N_5310);
or U6602 (N_6602,N_5024,N_4008);
nand U6603 (N_6603,N_5505,N_5041);
nor U6604 (N_6604,N_4361,N_4685);
and U6605 (N_6605,N_5414,N_4858);
and U6606 (N_6606,N_5676,N_5718);
nor U6607 (N_6607,N_5693,N_4186);
nand U6608 (N_6608,N_5896,N_4292);
nor U6609 (N_6609,N_5962,N_5480);
and U6610 (N_6610,N_5064,N_5320);
nand U6611 (N_6611,N_4570,N_4727);
nand U6612 (N_6612,N_5596,N_5130);
nor U6613 (N_6613,N_4447,N_4015);
and U6614 (N_6614,N_4474,N_4981);
nor U6615 (N_6615,N_5997,N_4013);
nand U6616 (N_6616,N_4035,N_4841);
and U6617 (N_6617,N_4438,N_5478);
and U6618 (N_6618,N_4672,N_5268);
nor U6619 (N_6619,N_4690,N_4541);
and U6620 (N_6620,N_5403,N_4045);
and U6621 (N_6621,N_4156,N_4752);
or U6622 (N_6622,N_5528,N_4670);
nand U6623 (N_6623,N_5290,N_5645);
nor U6624 (N_6624,N_5098,N_4450);
xor U6625 (N_6625,N_4205,N_5206);
nand U6626 (N_6626,N_4452,N_4934);
nor U6627 (N_6627,N_4301,N_4784);
or U6628 (N_6628,N_4446,N_5231);
nor U6629 (N_6629,N_4985,N_5225);
or U6630 (N_6630,N_4100,N_5601);
and U6631 (N_6631,N_5833,N_4708);
or U6632 (N_6632,N_5998,N_5287);
nor U6633 (N_6633,N_5369,N_5755);
nor U6634 (N_6634,N_4931,N_4738);
nor U6635 (N_6635,N_4034,N_5072);
nand U6636 (N_6636,N_4873,N_4468);
or U6637 (N_6637,N_5018,N_5598);
and U6638 (N_6638,N_5508,N_4116);
or U6639 (N_6639,N_5149,N_4836);
xor U6640 (N_6640,N_5065,N_4317);
and U6641 (N_6641,N_5055,N_5570);
and U6642 (N_6642,N_4617,N_4864);
or U6643 (N_6643,N_4486,N_4947);
and U6644 (N_6644,N_5957,N_5223);
nand U6645 (N_6645,N_5562,N_5732);
or U6646 (N_6646,N_4950,N_4877);
and U6647 (N_6647,N_4381,N_5875);
or U6648 (N_6648,N_4578,N_5958);
and U6649 (N_6649,N_5005,N_5417);
nand U6650 (N_6650,N_5222,N_4851);
or U6651 (N_6651,N_5993,N_5983);
nand U6652 (N_6652,N_5710,N_5468);
or U6653 (N_6653,N_4773,N_4531);
or U6654 (N_6654,N_5657,N_5863);
and U6655 (N_6655,N_4374,N_4376);
or U6656 (N_6656,N_5111,N_5637);
nor U6657 (N_6657,N_4424,N_5638);
or U6658 (N_6658,N_4849,N_5043);
or U6659 (N_6659,N_5959,N_4818);
nand U6660 (N_6660,N_4369,N_5340);
and U6661 (N_6661,N_4684,N_5080);
or U6662 (N_6662,N_4509,N_5692);
and U6663 (N_6663,N_4296,N_4879);
xnor U6664 (N_6664,N_4032,N_5616);
and U6665 (N_6665,N_5341,N_5540);
nand U6666 (N_6666,N_5500,N_5916);
or U6667 (N_6667,N_5526,N_5301);
and U6668 (N_6668,N_5425,N_5179);
and U6669 (N_6669,N_5708,N_4859);
nor U6670 (N_6670,N_4755,N_4055);
or U6671 (N_6671,N_4031,N_4909);
nor U6672 (N_6672,N_4030,N_4547);
or U6673 (N_6673,N_5121,N_4792);
nor U6674 (N_6674,N_4196,N_5625);
or U6675 (N_6675,N_4079,N_5667);
or U6676 (N_6676,N_5928,N_4293);
or U6677 (N_6677,N_4265,N_5486);
or U6678 (N_6678,N_5558,N_4926);
nor U6679 (N_6679,N_5531,N_5811);
nand U6680 (N_6680,N_4433,N_5321);
nand U6681 (N_6681,N_4215,N_4829);
and U6682 (N_6682,N_5532,N_4749);
and U6683 (N_6683,N_5591,N_5399);
or U6684 (N_6684,N_5806,N_5437);
nand U6685 (N_6685,N_5607,N_4435);
and U6686 (N_6686,N_5510,N_4237);
nor U6687 (N_6687,N_4510,N_5877);
nand U6688 (N_6688,N_5752,N_5176);
nor U6689 (N_6689,N_5376,N_4637);
and U6690 (N_6690,N_5886,N_4327);
and U6691 (N_6691,N_4889,N_5651);
and U6692 (N_6692,N_5465,N_4127);
nand U6693 (N_6693,N_4484,N_4919);
or U6694 (N_6694,N_4201,N_4630);
and U6695 (N_6695,N_5022,N_5784);
nor U6696 (N_6696,N_4977,N_5685);
nor U6697 (N_6697,N_5742,N_5273);
nand U6698 (N_6698,N_4303,N_5017);
or U6699 (N_6699,N_4092,N_4318);
nand U6700 (N_6700,N_4537,N_5224);
nor U6701 (N_6701,N_5390,N_5476);
or U6702 (N_6702,N_5932,N_5446);
nand U6703 (N_6703,N_5455,N_5217);
nor U6704 (N_6704,N_4219,N_5102);
or U6705 (N_6705,N_4984,N_4754);
and U6706 (N_6706,N_5518,N_4778);
nor U6707 (N_6707,N_4252,N_4884);
or U6708 (N_6708,N_5233,N_5802);
nand U6709 (N_6709,N_4658,N_5318);
nor U6710 (N_6710,N_5333,N_4696);
or U6711 (N_6711,N_4454,N_5327);
and U6712 (N_6712,N_5377,N_4203);
or U6713 (N_6713,N_4224,N_5241);
or U6714 (N_6714,N_5411,N_4807);
nor U6715 (N_6715,N_5907,N_4923);
or U6716 (N_6716,N_4955,N_4813);
nand U6717 (N_6717,N_5855,N_4967);
or U6718 (N_6718,N_4608,N_4411);
xnor U6719 (N_6719,N_4945,N_5982);
or U6720 (N_6720,N_4805,N_4831);
nor U6721 (N_6721,N_4753,N_5793);
or U6722 (N_6722,N_4199,N_5673);
and U6723 (N_6723,N_4239,N_4046);
nor U6724 (N_6724,N_4004,N_5548);
or U6725 (N_6725,N_4782,N_5374);
and U6726 (N_6726,N_4938,N_5175);
and U6727 (N_6727,N_4598,N_4393);
and U6728 (N_6728,N_5165,N_5257);
and U6729 (N_6729,N_5579,N_5608);
nand U6730 (N_6730,N_5386,N_5423);
nand U6731 (N_6731,N_5447,N_4133);
and U6732 (N_6732,N_5201,N_5332);
nand U6733 (N_6733,N_4993,N_4233);
nor U6734 (N_6734,N_5881,N_5589);
or U6735 (N_6735,N_4371,N_5828);
and U6736 (N_6736,N_5269,N_4395);
nand U6737 (N_6737,N_4175,N_5507);
nand U6738 (N_6738,N_4082,N_4652);
and U6739 (N_6739,N_5239,N_5872);
and U6740 (N_6740,N_4417,N_4573);
nor U6741 (N_6741,N_5406,N_5220);
or U6742 (N_6742,N_5714,N_5925);
or U6743 (N_6743,N_4645,N_5462);
nor U6744 (N_6744,N_4683,N_5850);
or U6745 (N_6745,N_5132,N_4429);
xnor U6746 (N_6746,N_4096,N_5003);
nor U6747 (N_6747,N_5238,N_4646);
nand U6748 (N_6748,N_4590,N_5849);
xnor U6749 (N_6749,N_5816,N_5678);
nand U6750 (N_6750,N_4470,N_5680);
nor U6751 (N_6751,N_4732,N_4141);
nor U6752 (N_6752,N_4533,N_4691);
and U6753 (N_6753,N_5773,N_5529);
or U6754 (N_6754,N_5088,N_4258);
and U6755 (N_6755,N_4629,N_4392);
or U6756 (N_6756,N_5456,N_4767);
xor U6757 (N_6757,N_4054,N_4266);
and U6758 (N_6758,N_5472,N_5815);
and U6759 (N_6759,N_5988,N_4525);
or U6760 (N_6760,N_5032,N_5234);
nor U6761 (N_6761,N_5803,N_4093);
nor U6762 (N_6762,N_4556,N_4648);
nor U6763 (N_6763,N_4675,N_5920);
nand U6764 (N_6764,N_5887,N_4899);
nor U6765 (N_6765,N_5777,N_4584);
nor U6766 (N_6766,N_5937,N_5131);
and U6767 (N_6767,N_5209,N_5623);
or U6768 (N_6768,N_5785,N_4939);
nand U6769 (N_6769,N_4375,N_4387);
nor U6770 (N_6770,N_4355,N_5757);
nor U6771 (N_6771,N_5650,N_5689);
nor U6772 (N_6772,N_4603,N_4928);
or U6773 (N_6773,N_5841,N_5615);
nand U6774 (N_6774,N_5629,N_4285);
and U6775 (N_6775,N_4814,N_4331);
or U6776 (N_6776,N_4220,N_5614);
nand U6777 (N_6777,N_5865,N_4464);
and U6778 (N_6778,N_5690,N_5736);
nand U6779 (N_6779,N_5636,N_5048);
nand U6780 (N_6780,N_5190,N_5251);
nand U6781 (N_6781,N_5733,N_4761);
and U6782 (N_6782,N_5727,N_5789);
nor U6783 (N_6783,N_4527,N_5460);
nand U6784 (N_6784,N_5969,N_5219);
or U6785 (N_6785,N_5706,N_4925);
nor U6786 (N_6786,N_4999,N_4599);
or U6787 (N_6787,N_5734,N_5413);
or U6788 (N_6788,N_4213,N_5968);
or U6789 (N_6789,N_4300,N_5517);
nand U6790 (N_6790,N_4404,N_5135);
and U6791 (N_6791,N_5489,N_5137);
nand U6792 (N_6792,N_4472,N_5441);
nor U6793 (N_6793,N_5512,N_5300);
and U6794 (N_6794,N_4178,N_4188);
nor U6795 (N_6795,N_5981,N_4770);
or U6796 (N_6796,N_4334,N_4021);
nor U6797 (N_6797,N_5052,N_4530);
nand U6798 (N_6798,N_5485,N_4920);
or U6799 (N_6799,N_4307,N_5817);
nand U6800 (N_6800,N_4210,N_4551);
nand U6801 (N_6801,N_4601,N_4528);
or U6802 (N_6802,N_4978,N_4653);
nor U6803 (N_6803,N_5934,N_5195);
or U6804 (N_6804,N_4855,N_4380);
and U6805 (N_6805,N_4056,N_4997);
or U6806 (N_6806,N_4545,N_5261);
nand U6807 (N_6807,N_4363,N_5565);
nor U6808 (N_6808,N_5813,N_5563);
nor U6809 (N_6809,N_4820,N_5766);
nand U6810 (N_6810,N_4106,N_5516);
nand U6811 (N_6811,N_4587,N_4847);
and U6812 (N_6812,N_5487,N_5304);
and U6813 (N_6813,N_4086,N_5442);
nor U6814 (N_6814,N_5405,N_5782);
nand U6815 (N_6815,N_4602,N_5836);
and U6816 (N_6816,N_5008,N_4211);
or U6817 (N_6817,N_4388,N_4362);
xnor U6818 (N_6818,N_5148,N_5288);
nor U6819 (N_6819,N_5497,N_4539);
nand U6820 (N_6820,N_4674,N_4000);
nand U6821 (N_6821,N_4440,N_5463);
and U6822 (N_6822,N_5240,N_4741);
and U6823 (N_6823,N_5344,N_5599);
or U6824 (N_6824,N_4389,N_4832);
or U6825 (N_6825,N_4249,N_4341);
nor U6826 (N_6826,N_5704,N_5471);
nand U6827 (N_6827,N_4154,N_4620);
and U6828 (N_6828,N_5767,N_4554);
nor U6829 (N_6829,N_5181,N_4697);
or U6830 (N_6830,N_4835,N_5559);
nor U6831 (N_6831,N_4421,N_5539);
or U6832 (N_6832,N_5382,N_4169);
nand U6833 (N_6833,N_5400,N_4009);
or U6834 (N_6834,N_4023,N_4385);
nand U6835 (N_6835,N_5359,N_4179);
and U6836 (N_6836,N_4746,N_4431);
and U6837 (N_6837,N_4927,N_4121);
or U6838 (N_6838,N_5264,N_4250);
nor U6839 (N_6839,N_5180,N_4776);
nor U6840 (N_6840,N_4136,N_5028);
nand U6841 (N_6841,N_4038,N_5585);
nand U6842 (N_6842,N_4123,N_4597);
nand U6843 (N_6843,N_4717,N_5396);
nand U6844 (N_6844,N_4577,N_4399);
nand U6845 (N_6845,N_5856,N_4073);
nand U6846 (N_6846,N_4267,N_5110);
nand U6847 (N_6847,N_4804,N_4478);
and U6848 (N_6848,N_5494,N_4632);
and U6849 (N_6849,N_4688,N_5683);
nand U6850 (N_6850,N_4796,N_5188);
or U6851 (N_6851,N_5051,N_4247);
or U6852 (N_6852,N_5428,N_4839);
nand U6853 (N_6853,N_4520,N_4466);
nor U6854 (N_6854,N_5986,N_5520);
nand U6855 (N_6855,N_4495,N_5078);
nor U6856 (N_6856,N_4236,N_4016);
or U6857 (N_6857,N_4883,N_4718);
nor U6858 (N_6858,N_5506,N_4555);
nor U6859 (N_6859,N_5392,N_5715);
nand U6860 (N_6860,N_4803,N_5292);
nor U6861 (N_6861,N_5822,N_5145);
or U6862 (N_6862,N_5788,N_4677);
or U6863 (N_6863,N_5104,N_5859);
nand U6864 (N_6864,N_5395,N_5227);
nand U6865 (N_6865,N_4120,N_4115);
and U6866 (N_6866,N_5435,N_4182);
nor U6867 (N_6867,N_4605,N_4207);
or U6868 (N_6868,N_4003,N_5917);
or U6869 (N_6869,N_4766,N_4952);
and U6870 (N_6870,N_5270,N_5681);
or U6871 (N_6871,N_5594,N_4917);
and U6872 (N_6872,N_4894,N_5166);
and U6873 (N_6873,N_5627,N_5864);
or U6874 (N_6874,N_4772,N_4693);
nor U6875 (N_6875,N_4657,N_5722);
nor U6876 (N_6876,N_4496,N_5946);
nand U6877 (N_6877,N_4771,N_4146);
nand U6878 (N_6878,N_4501,N_4356);
or U6879 (N_6879,N_5326,N_4425);
and U6880 (N_6880,N_5197,N_4915);
or U6881 (N_6881,N_5193,N_5649);
and U6882 (N_6882,N_5858,N_5643);
nor U6883 (N_6883,N_4871,N_5883);
nand U6884 (N_6884,N_5675,N_5291);
nand U6885 (N_6885,N_4039,N_5550);
and U6886 (N_6886,N_5882,N_4714);
nand U6887 (N_6887,N_4315,N_4386);
or U6888 (N_6888,N_5082,N_4631);
and U6889 (N_6889,N_4682,N_5127);
and U6890 (N_6890,N_4347,N_5044);
or U6891 (N_6891,N_4194,N_4119);
or U6892 (N_6892,N_5955,N_5910);
and U6893 (N_6893,N_4135,N_4797);
and U6894 (N_6894,N_5911,N_4413);
and U6895 (N_6895,N_4493,N_4662);
nor U6896 (N_6896,N_5368,N_5731);
nor U6897 (N_6897,N_4961,N_5921);
and U6898 (N_6898,N_5631,N_5663);
or U6899 (N_6899,N_5087,N_5434);
and U6900 (N_6900,N_5448,N_4821);
nand U6901 (N_6901,N_5467,N_4515);
nor U6902 (N_6902,N_4857,N_5798);
nor U6903 (N_6903,N_4944,N_4483);
nor U6904 (N_6904,N_5004,N_5323);
nand U6905 (N_6905,N_4081,N_5971);
and U6906 (N_6906,N_5662,N_4343);
and U6907 (N_6907,N_4222,N_5561);
nor U6908 (N_6908,N_4887,N_4581);
nor U6909 (N_6909,N_5387,N_4491);
or U6910 (N_6910,N_5152,N_5138);
nor U6911 (N_6911,N_5820,N_5155);
nand U6912 (N_6912,N_4225,N_5717);
nand U6913 (N_6913,N_4259,N_4500);
or U6914 (N_6914,N_4508,N_4074);
or U6915 (N_6915,N_5769,N_5931);
or U6916 (N_6916,N_4134,N_4173);
and U6917 (N_6917,N_4848,N_5443);
and U6918 (N_6918,N_4427,N_5308);
or U6919 (N_6919,N_4235,N_4540);
and U6920 (N_6920,N_4874,N_5909);
and U6921 (N_6921,N_4868,N_4880);
and U6922 (N_6922,N_5204,N_4060);
nand U6923 (N_6923,N_5525,N_4786);
or U6924 (N_6924,N_4576,N_5335);
or U6925 (N_6925,N_5648,N_4963);
or U6926 (N_6926,N_4695,N_4162);
and U6927 (N_6927,N_4218,N_5331);
and U6928 (N_6928,N_5035,N_5716);
and U6929 (N_6929,N_5243,N_5345);
or U6930 (N_6930,N_5470,N_5105);
and U6931 (N_6931,N_4671,N_5464);
nor U6932 (N_6932,N_4457,N_4972);
nor U6933 (N_6933,N_4378,N_5867);
nand U6934 (N_6934,N_5027,N_4428);
and U6935 (N_6935,N_4434,N_5547);
nand U6936 (N_6936,N_4125,N_4062);
nor U6937 (N_6937,N_4067,N_4744);
and U6938 (N_6938,N_4246,N_5666);
and U6939 (N_6939,N_5367,N_5228);
nor U6940 (N_6940,N_4109,N_4286);
nor U6941 (N_6941,N_5196,N_4888);
or U6942 (N_6942,N_4640,N_4940);
nor U6943 (N_6943,N_5975,N_5646);
nor U6944 (N_6944,N_4737,N_5053);
nor U6945 (N_6945,N_4811,N_5857);
nor U6946 (N_6946,N_4157,N_4957);
nor U6947 (N_6947,N_5546,N_5067);
and U6948 (N_6948,N_5994,N_5612);
or U6949 (N_6949,N_4980,N_4585);
nor U6950 (N_6950,N_4174,N_5136);
nor U6951 (N_6951,N_5061,N_4571);
or U6952 (N_6952,N_5389,N_5832);
nor U6953 (N_6953,N_5853,N_5473);
and U6954 (N_6954,N_5522,N_5743);
or U6955 (N_6955,N_4195,N_5669);
nor U6956 (N_6956,N_5346,N_5361);
nor U6957 (N_6957,N_5250,N_4659);
or U6958 (N_6958,N_4050,N_4269);
and U6959 (N_6959,N_5366,N_4777);
or U6960 (N_6960,N_4769,N_5049);
and U6961 (N_6961,N_4679,N_5655);
nand U6962 (N_6962,N_5687,N_5964);
or U6963 (N_6963,N_5609,N_5477);
or U6964 (N_6964,N_5791,N_4445);
nand U6965 (N_6965,N_4739,N_5192);
nor U6966 (N_6966,N_5328,N_5541);
and U6967 (N_6967,N_4185,N_5259);
or U6968 (N_6968,N_4217,N_5885);
and U6969 (N_6969,N_4479,N_4423);
or U6970 (N_6970,N_5519,N_4189);
nand U6971 (N_6971,N_4709,N_4432);
nand U6972 (N_6972,N_4914,N_4069);
nor U6973 (N_6973,N_5807,N_4216);
nand U6974 (N_6974,N_5124,N_5979);
or U6975 (N_6975,N_4791,N_4711);
nand U6976 (N_6976,N_4751,N_5491);
nand U6977 (N_6977,N_5343,N_5577);
and U6978 (N_6978,N_5861,N_4823);
or U6979 (N_6979,N_5573,N_5133);
and U6980 (N_6980,N_5805,N_5659);
nand U6981 (N_6981,N_5319,N_4762);
and U6982 (N_6982,N_5059,N_4641);
nor U6983 (N_6983,N_4294,N_4230);
nor U6984 (N_6984,N_4126,N_4305);
and U6985 (N_6985,N_5950,N_5370);
nand U6986 (N_6986,N_4354,N_4227);
nor U6987 (N_6987,N_5394,N_4613);
nand U6988 (N_6988,N_5595,N_4397);
or U6989 (N_6989,N_5076,N_4287);
nor U6990 (N_6990,N_4850,N_5989);
and U6991 (N_6991,N_5056,N_5897);
or U6992 (N_6992,N_5796,N_5296);
nand U6993 (N_6993,N_4306,N_4206);
or U6994 (N_6994,N_5280,N_5036);
and U6995 (N_6995,N_4596,N_4724);
and U6996 (N_6996,N_5091,N_5307);
or U6997 (N_6997,N_5606,N_5555);
or U6998 (N_6998,N_5244,N_5037);
nand U6999 (N_6999,N_5351,N_4451);
and U7000 (N_7000,N_5183,N_4051);
or U7001 (N_7001,N_4857,N_4543);
and U7002 (N_7002,N_5862,N_4907);
or U7003 (N_7003,N_4239,N_4150);
nand U7004 (N_7004,N_5783,N_5430);
and U7005 (N_7005,N_4898,N_5752);
nor U7006 (N_7006,N_4966,N_5755);
and U7007 (N_7007,N_5360,N_4689);
or U7008 (N_7008,N_5361,N_5815);
nand U7009 (N_7009,N_5916,N_5014);
and U7010 (N_7010,N_5095,N_5439);
and U7011 (N_7011,N_5514,N_4170);
or U7012 (N_7012,N_4614,N_4687);
and U7013 (N_7013,N_5605,N_4535);
and U7014 (N_7014,N_4359,N_5628);
nand U7015 (N_7015,N_5706,N_4830);
nor U7016 (N_7016,N_4596,N_4801);
nor U7017 (N_7017,N_4870,N_5240);
and U7018 (N_7018,N_5611,N_4240);
or U7019 (N_7019,N_5993,N_4742);
nor U7020 (N_7020,N_4203,N_5772);
nor U7021 (N_7021,N_4068,N_5024);
nor U7022 (N_7022,N_5355,N_5263);
xor U7023 (N_7023,N_4937,N_5219);
nor U7024 (N_7024,N_5704,N_5067);
and U7025 (N_7025,N_5268,N_5701);
nand U7026 (N_7026,N_5060,N_4550);
nor U7027 (N_7027,N_4562,N_4771);
nor U7028 (N_7028,N_4002,N_4906);
nand U7029 (N_7029,N_5852,N_4775);
nor U7030 (N_7030,N_5058,N_5615);
nand U7031 (N_7031,N_4967,N_5935);
or U7032 (N_7032,N_4418,N_4891);
xnor U7033 (N_7033,N_5715,N_5774);
nand U7034 (N_7034,N_4197,N_5505);
nand U7035 (N_7035,N_4063,N_5248);
and U7036 (N_7036,N_4002,N_5886);
nor U7037 (N_7037,N_5043,N_4790);
and U7038 (N_7038,N_5142,N_5892);
nor U7039 (N_7039,N_5330,N_4348);
and U7040 (N_7040,N_5315,N_4170);
nor U7041 (N_7041,N_4435,N_4050);
and U7042 (N_7042,N_5396,N_5823);
and U7043 (N_7043,N_4811,N_5855);
or U7044 (N_7044,N_5163,N_4602);
and U7045 (N_7045,N_5860,N_5927);
or U7046 (N_7046,N_4948,N_5865);
or U7047 (N_7047,N_5848,N_5574);
or U7048 (N_7048,N_5838,N_5474);
or U7049 (N_7049,N_4101,N_5200);
nand U7050 (N_7050,N_4835,N_4414);
and U7051 (N_7051,N_4016,N_5037);
or U7052 (N_7052,N_5164,N_4774);
nor U7053 (N_7053,N_4780,N_4400);
or U7054 (N_7054,N_4101,N_4512);
nor U7055 (N_7055,N_4721,N_5971);
or U7056 (N_7056,N_5136,N_4855);
and U7057 (N_7057,N_5836,N_4808);
nand U7058 (N_7058,N_5189,N_5034);
nor U7059 (N_7059,N_5902,N_5741);
nor U7060 (N_7060,N_5885,N_4753);
nor U7061 (N_7061,N_4363,N_5366);
nand U7062 (N_7062,N_5385,N_4424);
nand U7063 (N_7063,N_5447,N_4447);
and U7064 (N_7064,N_4293,N_5738);
or U7065 (N_7065,N_5999,N_4966);
nor U7066 (N_7066,N_5060,N_4699);
nand U7067 (N_7067,N_5449,N_5433);
and U7068 (N_7068,N_5414,N_4917);
nand U7069 (N_7069,N_4058,N_4038);
or U7070 (N_7070,N_4673,N_5046);
and U7071 (N_7071,N_5722,N_5921);
nand U7072 (N_7072,N_4023,N_5753);
and U7073 (N_7073,N_5885,N_5978);
nand U7074 (N_7074,N_4502,N_4302);
nor U7075 (N_7075,N_5564,N_5711);
and U7076 (N_7076,N_4260,N_5323);
or U7077 (N_7077,N_5193,N_4253);
nand U7078 (N_7078,N_4166,N_4074);
nand U7079 (N_7079,N_4122,N_4510);
and U7080 (N_7080,N_4138,N_4830);
nor U7081 (N_7081,N_4109,N_4637);
nor U7082 (N_7082,N_4738,N_5080);
nor U7083 (N_7083,N_4784,N_5192);
nand U7084 (N_7084,N_4144,N_5750);
and U7085 (N_7085,N_5743,N_4551);
and U7086 (N_7086,N_4329,N_5938);
nor U7087 (N_7087,N_5503,N_4556);
or U7088 (N_7088,N_4885,N_5179);
nand U7089 (N_7089,N_5740,N_4960);
nand U7090 (N_7090,N_4029,N_4743);
and U7091 (N_7091,N_4462,N_4886);
nand U7092 (N_7092,N_5255,N_4253);
nand U7093 (N_7093,N_4376,N_4385);
nor U7094 (N_7094,N_5668,N_4760);
nor U7095 (N_7095,N_4622,N_5984);
xor U7096 (N_7096,N_5296,N_4066);
nand U7097 (N_7097,N_5441,N_5890);
nand U7098 (N_7098,N_5473,N_4641);
nor U7099 (N_7099,N_5547,N_5624);
nor U7100 (N_7100,N_4794,N_4472);
nor U7101 (N_7101,N_4345,N_4198);
nand U7102 (N_7102,N_5687,N_4089);
and U7103 (N_7103,N_4237,N_4961);
nand U7104 (N_7104,N_4976,N_4625);
xnor U7105 (N_7105,N_4115,N_5545);
or U7106 (N_7106,N_4546,N_5091);
and U7107 (N_7107,N_4815,N_4308);
or U7108 (N_7108,N_4526,N_5651);
nand U7109 (N_7109,N_5097,N_5632);
and U7110 (N_7110,N_4763,N_5857);
nor U7111 (N_7111,N_4794,N_4220);
or U7112 (N_7112,N_4057,N_4476);
or U7113 (N_7113,N_5962,N_5403);
and U7114 (N_7114,N_4854,N_5568);
or U7115 (N_7115,N_4484,N_4504);
and U7116 (N_7116,N_5797,N_4906);
or U7117 (N_7117,N_4844,N_4525);
and U7118 (N_7118,N_5776,N_5731);
and U7119 (N_7119,N_5060,N_4921);
and U7120 (N_7120,N_4620,N_4521);
and U7121 (N_7121,N_4218,N_5186);
xor U7122 (N_7122,N_4929,N_4127);
nand U7123 (N_7123,N_5226,N_4463);
nor U7124 (N_7124,N_5637,N_5287);
nand U7125 (N_7125,N_5772,N_5253);
or U7126 (N_7126,N_5255,N_4079);
nor U7127 (N_7127,N_4417,N_5274);
nor U7128 (N_7128,N_5313,N_4858);
or U7129 (N_7129,N_5742,N_4334);
or U7130 (N_7130,N_5830,N_4553);
nand U7131 (N_7131,N_4498,N_5425);
or U7132 (N_7132,N_4678,N_5646);
or U7133 (N_7133,N_4576,N_5639);
nand U7134 (N_7134,N_5791,N_4737);
or U7135 (N_7135,N_5615,N_4215);
nand U7136 (N_7136,N_4745,N_5081);
nor U7137 (N_7137,N_5639,N_5983);
nand U7138 (N_7138,N_5004,N_5336);
and U7139 (N_7139,N_5198,N_4825);
xor U7140 (N_7140,N_4263,N_5220);
nor U7141 (N_7141,N_4910,N_4626);
and U7142 (N_7142,N_5231,N_4797);
nand U7143 (N_7143,N_5800,N_4286);
nor U7144 (N_7144,N_5044,N_5228);
nor U7145 (N_7145,N_5595,N_5323);
or U7146 (N_7146,N_5777,N_5413);
nand U7147 (N_7147,N_4571,N_5709);
and U7148 (N_7148,N_5936,N_4405);
and U7149 (N_7149,N_4190,N_4446);
or U7150 (N_7150,N_5121,N_4721);
nor U7151 (N_7151,N_4113,N_4667);
nor U7152 (N_7152,N_5013,N_4008);
or U7153 (N_7153,N_5539,N_4797);
nor U7154 (N_7154,N_5576,N_5197);
or U7155 (N_7155,N_4113,N_4005);
and U7156 (N_7156,N_4343,N_5178);
nand U7157 (N_7157,N_5165,N_4694);
nor U7158 (N_7158,N_4752,N_5057);
and U7159 (N_7159,N_4995,N_4172);
and U7160 (N_7160,N_4986,N_5054);
or U7161 (N_7161,N_4768,N_5705);
nand U7162 (N_7162,N_5995,N_4769);
nand U7163 (N_7163,N_4594,N_5620);
nand U7164 (N_7164,N_4104,N_4484);
nand U7165 (N_7165,N_5795,N_5811);
nand U7166 (N_7166,N_5961,N_4275);
xor U7167 (N_7167,N_4974,N_4128);
nand U7168 (N_7168,N_4777,N_4750);
and U7169 (N_7169,N_5684,N_5680);
nor U7170 (N_7170,N_4909,N_5885);
or U7171 (N_7171,N_5637,N_4423);
nor U7172 (N_7172,N_5159,N_5797);
and U7173 (N_7173,N_5732,N_5508);
nand U7174 (N_7174,N_4305,N_4293);
or U7175 (N_7175,N_4842,N_4359);
or U7176 (N_7176,N_4145,N_5767);
nand U7177 (N_7177,N_5494,N_5833);
and U7178 (N_7178,N_4362,N_5373);
nor U7179 (N_7179,N_4508,N_5345);
nor U7180 (N_7180,N_5055,N_5422);
and U7181 (N_7181,N_5678,N_4646);
or U7182 (N_7182,N_5682,N_5414);
nor U7183 (N_7183,N_5492,N_4969);
nor U7184 (N_7184,N_4851,N_4833);
or U7185 (N_7185,N_5977,N_5775);
nor U7186 (N_7186,N_4528,N_4079);
or U7187 (N_7187,N_4498,N_5548);
nand U7188 (N_7188,N_5453,N_4759);
or U7189 (N_7189,N_5283,N_4640);
nand U7190 (N_7190,N_4033,N_4711);
or U7191 (N_7191,N_5275,N_4757);
nor U7192 (N_7192,N_5575,N_5951);
or U7193 (N_7193,N_4953,N_5004);
and U7194 (N_7194,N_5978,N_5417);
nor U7195 (N_7195,N_4727,N_5488);
nand U7196 (N_7196,N_4859,N_4596);
and U7197 (N_7197,N_4519,N_5646);
or U7198 (N_7198,N_4280,N_4180);
nand U7199 (N_7199,N_5529,N_5798);
and U7200 (N_7200,N_4334,N_5112);
and U7201 (N_7201,N_4871,N_4737);
nand U7202 (N_7202,N_5157,N_5376);
and U7203 (N_7203,N_4832,N_4742);
nand U7204 (N_7204,N_4606,N_4998);
or U7205 (N_7205,N_4973,N_4523);
nand U7206 (N_7206,N_5811,N_4212);
and U7207 (N_7207,N_5086,N_5573);
nand U7208 (N_7208,N_4538,N_4931);
nor U7209 (N_7209,N_5967,N_4639);
nand U7210 (N_7210,N_4761,N_5433);
or U7211 (N_7211,N_4372,N_4131);
nand U7212 (N_7212,N_5890,N_5651);
and U7213 (N_7213,N_4080,N_4765);
nor U7214 (N_7214,N_4652,N_5510);
nor U7215 (N_7215,N_5550,N_5650);
or U7216 (N_7216,N_4276,N_5025);
or U7217 (N_7217,N_4834,N_4537);
nor U7218 (N_7218,N_5662,N_4361);
and U7219 (N_7219,N_4595,N_5870);
or U7220 (N_7220,N_4392,N_5761);
or U7221 (N_7221,N_5891,N_5081);
xnor U7222 (N_7222,N_5294,N_4076);
and U7223 (N_7223,N_5342,N_5805);
nand U7224 (N_7224,N_5046,N_5985);
nand U7225 (N_7225,N_5405,N_4209);
nor U7226 (N_7226,N_4569,N_5990);
and U7227 (N_7227,N_5616,N_4251);
or U7228 (N_7228,N_4340,N_4801);
or U7229 (N_7229,N_4037,N_5245);
nor U7230 (N_7230,N_4553,N_5100);
or U7231 (N_7231,N_4020,N_5885);
nor U7232 (N_7232,N_4129,N_5606);
nand U7233 (N_7233,N_5078,N_4979);
or U7234 (N_7234,N_4932,N_4033);
and U7235 (N_7235,N_5517,N_4962);
or U7236 (N_7236,N_5057,N_5483);
xnor U7237 (N_7237,N_4295,N_5038);
nand U7238 (N_7238,N_4392,N_4139);
and U7239 (N_7239,N_4838,N_5267);
nand U7240 (N_7240,N_4040,N_5053);
and U7241 (N_7241,N_4713,N_5667);
and U7242 (N_7242,N_4368,N_4353);
or U7243 (N_7243,N_5452,N_4883);
and U7244 (N_7244,N_5853,N_5774);
and U7245 (N_7245,N_4229,N_5402);
or U7246 (N_7246,N_4835,N_5472);
or U7247 (N_7247,N_4046,N_5709);
or U7248 (N_7248,N_5137,N_5971);
nand U7249 (N_7249,N_4212,N_4396);
nor U7250 (N_7250,N_5894,N_4825);
nand U7251 (N_7251,N_5525,N_4051);
nor U7252 (N_7252,N_5103,N_4016);
or U7253 (N_7253,N_5257,N_5028);
and U7254 (N_7254,N_5491,N_5011);
and U7255 (N_7255,N_5396,N_4176);
or U7256 (N_7256,N_4906,N_5014);
nand U7257 (N_7257,N_4422,N_5975);
or U7258 (N_7258,N_5301,N_5118);
nand U7259 (N_7259,N_5872,N_5833);
nor U7260 (N_7260,N_4022,N_4745);
nor U7261 (N_7261,N_4038,N_4587);
nor U7262 (N_7262,N_5307,N_5718);
and U7263 (N_7263,N_5906,N_5855);
or U7264 (N_7264,N_5322,N_4292);
or U7265 (N_7265,N_4473,N_4363);
and U7266 (N_7266,N_5786,N_5772);
nor U7267 (N_7267,N_4923,N_5721);
nor U7268 (N_7268,N_5223,N_4341);
and U7269 (N_7269,N_4131,N_5194);
nand U7270 (N_7270,N_5591,N_5251);
nor U7271 (N_7271,N_5104,N_5436);
or U7272 (N_7272,N_5541,N_5013);
nand U7273 (N_7273,N_5824,N_4797);
nor U7274 (N_7274,N_5419,N_5256);
or U7275 (N_7275,N_5329,N_5160);
or U7276 (N_7276,N_4459,N_5138);
nand U7277 (N_7277,N_4009,N_4171);
nor U7278 (N_7278,N_4472,N_4160);
or U7279 (N_7279,N_4195,N_4864);
nand U7280 (N_7280,N_4822,N_4804);
xor U7281 (N_7281,N_5998,N_5473);
or U7282 (N_7282,N_5149,N_5977);
nor U7283 (N_7283,N_5610,N_4240);
and U7284 (N_7284,N_5221,N_4773);
nor U7285 (N_7285,N_4090,N_4594);
and U7286 (N_7286,N_4840,N_4057);
nor U7287 (N_7287,N_4009,N_4913);
and U7288 (N_7288,N_5239,N_5704);
or U7289 (N_7289,N_5507,N_4510);
or U7290 (N_7290,N_4995,N_5004);
nand U7291 (N_7291,N_4991,N_5849);
nor U7292 (N_7292,N_4610,N_4395);
and U7293 (N_7293,N_5731,N_4451);
or U7294 (N_7294,N_5616,N_5418);
nand U7295 (N_7295,N_4155,N_5838);
nand U7296 (N_7296,N_5069,N_5425);
nand U7297 (N_7297,N_4115,N_4020);
and U7298 (N_7298,N_4234,N_4837);
nor U7299 (N_7299,N_5644,N_4614);
or U7300 (N_7300,N_4560,N_5462);
nand U7301 (N_7301,N_4298,N_4719);
or U7302 (N_7302,N_5855,N_5268);
and U7303 (N_7303,N_4495,N_5711);
nand U7304 (N_7304,N_5841,N_5212);
xor U7305 (N_7305,N_4622,N_4008);
and U7306 (N_7306,N_4227,N_4690);
nor U7307 (N_7307,N_4008,N_5600);
nor U7308 (N_7308,N_4409,N_4287);
nor U7309 (N_7309,N_5578,N_4247);
nand U7310 (N_7310,N_4886,N_5345);
and U7311 (N_7311,N_5475,N_4940);
or U7312 (N_7312,N_5485,N_4488);
nor U7313 (N_7313,N_5852,N_5627);
and U7314 (N_7314,N_5131,N_4180);
nor U7315 (N_7315,N_4196,N_5698);
or U7316 (N_7316,N_4363,N_4686);
nand U7317 (N_7317,N_5429,N_5049);
nor U7318 (N_7318,N_5865,N_5816);
and U7319 (N_7319,N_5599,N_4722);
and U7320 (N_7320,N_4519,N_4029);
nand U7321 (N_7321,N_4510,N_5626);
nand U7322 (N_7322,N_5911,N_4025);
nand U7323 (N_7323,N_4060,N_4839);
nor U7324 (N_7324,N_4233,N_4258);
or U7325 (N_7325,N_5894,N_5673);
or U7326 (N_7326,N_5598,N_4209);
xor U7327 (N_7327,N_4051,N_4973);
or U7328 (N_7328,N_4889,N_4079);
or U7329 (N_7329,N_4637,N_5956);
nor U7330 (N_7330,N_4734,N_4719);
nor U7331 (N_7331,N_4592,N_4493);
nand U7332 (N_7332,N_4955,N_4789);
and U7333 (N_7333,N_5817,N_5640);
nor U7334 (N_7334,N_5206,N_4343);
xor U7335 (N_7335,N_4853,N_4088);
or U7336 (N_7336,N_5991,N_4092);
nor U7337 (N_7337,N_4986,N_4070);
xor U7338 (N_7338,N_5663,N_4853);
nor U7339 (N_7339,N_5015,N_5876);
nand U7340 (N_7340,N_4670,N_4629);
nand U7341 (N_7341,N_5650,N_5999);
or U7342 (N_7342,N_5369,N_4568);
or U7343 (N_7343,N_5156,N_5680);
xnor U7344 (N_7344,N_4278,N_4722);
and U7345 (N_7345,N_5523,N_4249);
nor U7346 (N_7346,N_5787,N_4306);
and U7347 (N_7347,N_4886,N_5714);
nand U7348 (N_7348,N_4244,N_5589);
and U7349 (N_7349,N_5401,N_5040);
nor U7350 (N_7350,N_4825,N_5834);
and U7351 (N_7351,N_4686,N_5490);
and U7352 (N_7352,N_4224,N_5118);
or U7353 (N_7353,N_5442,N_4884);
nor U7354 (N_7354,N_4310,N_5607);
nand U7355 (N_7355,N_4024,N_4406);
nor U7356 (N_7356,N_4972,N_4492);
and U7357 (N_7357,N_4815,N_4312);
and U7358 (N_7358,N_4798,N_4279);
nor U7359 (N_7359,N_4556,N_5143);
and U7360 (N_7360,N_4760,N_5889);
and U7361 (N_7361,N_4646,N_5911);
nand U7362 (N_7362,N_4923,N_4963);
and U7363 (N_7363,N_5080,N_5075);
xor U7364 (N_7364,N_4131,N_4260);
nand U7365 (N_7365,N_4042,N_4933);
and U7366 (N_7366,N_4359,N_5645);
nor U7367 (N_7367,N_4888,N_4560);
and U7368 (N_7368,N_4593,N_5686);
nand U7369 (N_7369,N_4332,N_4859);
or U7370 (N_7370,N_5970,N_5388);
nand U7371 (N_7371,N_4848,N_5681);
nor U7372 (N_7372,N_4458,N_4715);
and U7373 (N_7373,N_4524,N_4644);
nand U7374 (N_7374,N_5891,N_4006);
nand U7375 (N_7375,N_5024,N_4174);
nor U7376 (N_7376,N_5865,N_4353);
nand U7377 (N_7377,N_5950,N_4894);
nand U7378 (N_7378,N_4354,N_4154);
or U7379 (N_7379,N_4150,N_4299);
or U7380 (N_7380,N_4401,N_5898);
nand U7381 (N_7381,N_4772,N_5859);
or U7382 (N_7382,N_4420,N_5918);
nor U7383 (N_7383,N_4985,N_4535);
nand U7384 (N_7384,N_4152,N_4073);
and U7385 (N_7385,N_4628,N_4489);
nor U7386 (N_7386,N_4242,N_5267);
and U7387 (N_7387,N_5326,N_5255);
and U7388 (N_7388,N_5641,N_4659);
nand U7389 (N_7389,N_5235,N_5889);
or U7390 (N_7390,N_5607,N_4995);
nand U7391 (N_7391,N_5453,N_4207);
or U7392 (N_7392,N_5135,N_4667);
or U7393 (N_7393,N_5584,N_4414);
or U7394 (N_7394,N_4915,N_4527);
nand U7395 (N_7395,N_5354,N_5230);
nor U7396 (N_7396,N_4447,N_4516);
nand U7397 (N_7397,N_5706,N_5754);
and U7398 (N_7398,N_5278,N_4742);
or U7399 (N_7399,N_5872,N_5163);
and U7400 (N_7400,N_4807,N_4768);
and U7401 (N_7401,N_4076,N_4789);
nand U7402 (N_7402,N_4473,N_4305);
and U7403 (N_7403,N_5411,N_4823);
nor U7404 (N_7404,N_5423,N_4799);
or U7405 (N_7405,N_5741,N_5926);
and U7406 (N_7406,N_4556,N_5856);
nand U7407 (N_7407,N_5243,N_4565);
nand U7408 (N_7408,N_4692,N_5046);
and U7409 (N_7409,N_5672,N_5624);
or U7410 (N_7410,N_5011,N_5847);
and U7411 (N_7411,N_5808,N_4726);
or U7412 (N_7412,N_5679,N_5524);
or U7413 (N_7413,N_5776,N_5627);
or U7414 (N_7414,N_5426,N_5491);
or U7415 (N_7415,N_5976,N_4648);
and U7416 (N_7416,N_4509,N_4400);
or U7417 (N_7417,N_5674,N_4738);
nand U7418 (N_7418,N_5024,N_5946);
or U7419 (N_7419,N_5102,N_4990);
and U7420 (N_7420,N_5396,N_4578);
or U7421 (N_7421,N_5915,N_4179);
and U7422 (N_7422,N_5084,N_4058);
or U7423 (N_7423,N_5745,N_5525);
nor U7424 (N_7424,N_4999,N_5956);
nand U7425 (N_7425,N_4437,N_4442);
and U7426 (N_7426,N_4660,N_5605);
or U7427 (N_7427,N_4052,N_4678);
and U7428 (N_7428,N_4886,N_5837);
nand U7429 (N_7429,N_4609,N_4699);
or U7430 (N_7430,N_4392,N_5073);
and U7431 (N_7431,N_5974,N_5339);
nor U7432 (N_7432,N_5680,N_4769);
nor U7433 (N_7433,N_5469,N_4537);
nand U7434 (N_7434,N_5576,N_4234);
or U7435 (N_7435,N_4399,N_5014);
or U7436 (N_7436,N_4733,N_4206);
and U7437 (N_7437,N_4552,N_4262);
or U7438 (N_7438,N_5332,N_5070);
nor U7439 (N_7439,N_4563,N_5749);
or U7440 (N_7440,N_4682,N_5158);
and U7441 (N_7441,N_4256,N_5796);
nor U7442 (N_7442,N_4480,N_5158);
nand U7443 (N_7443,N_5509,N_5093);
nor U7444 (N_7444,N_4793,N_5786);
or U7445 (N_7445,N_4149,N_5532);
nor U7446 (N_7446,N_5986,N_4915);
or U7447 (N_7447,N_4649,N_4066);
and U7448 (N_7448,N_5238,N_5111);
or U7449 (N_7449,N_5123,N_5081);
and U7450 (N_7450,N_5323,N_5766);
nand U7451 (N_7451,N_5695,N_4661);
and U7452 (N_7452,N_4163,N_5640);
or U7453 (N_7453,N_5033,N_5114);
nand U7454 (N_7454,N_5108,N_5539);
nand U7455 (N_7455,N_5694,N_4006);
or U7456 (N_7456,N_4058,N_4099);
or U7457 (N_7457,N_5777,N_5835);
and U7458 (N_7458,N_5087,N_5938);
and U7459 (N_7459,N_5878,N_4035);
or U7460 (N_7460,N_5347,N_5388);
and U7461 (N_7461,N_4699,N_5120);
nand U7462 (N_7462,N_4650,N_5715);
and U7463 (N_7463,N_5655,N_5993);
nor U7464 (N_7464,N_4683,N_5868);
or U7465 (N_7465,N_4397,N_5971);
or U7466 (N_7466,N_4606,N_4065);
and U7467 (N_7467,N_4142,N_4498);
or U7468 (N_7468,N_4168,N_5015);
nand U7469 (N_7469,N_4783,N_5460);
nor U7470 (N_7470,N_4530,N_4082);
and U7471 (N_7471,N_4381,N_5027);
nand U7472 (N_7472,N_5880,N_4489);
nand U7473 (N_7473,N_5247,N_4616);
nor U7474 (N_7474,N_4436,N_4833);
nor U7475 (N_7475,N_5849,N_4946);
nor U7476 (N_7476,N_5557,N_4021);
nand U7477 (N_7477,N_4223,N_4801);
xnor U7478 (N_7478,N_5831,N_4702);
nor U7479 (N_7479,N_4622,N_5653);
nand U7480 (N_7480,N_4484,N_5106);
nor U7481 (N_7481,N_4161,N_5760);
nor U7482 (N_7482,N_5378,N_4677);
or U7483 (N_7483,N_4168,N_4056);
and U7484 (N_7484,N_4085,N_5864);
and U7485 (N_7485,N_5359,N_4331);
and U7486 (N_7486,N_5368,N_5531);
nand U7487 (N_7487,N_5073,N_4356);
or U7488 (N_7488,N_4249,N_5174);
nand U7489 (N_7489,N_5625,N_4922);
or U7490 (N_7490,N_4790,N_4740);
or U7491 (N_7491,N_4597,N_4590);
or U7492 (N_7492,N_4908,N_5188);
nand U7493 (N_7493,N_5140,N_4191);
xor U7494 (N_7494,N_4458,N_4511);
and U7495 (N_7495,N_4073,N_5601);
and U7496 (N_7496,N_5500,N_5901);
and U7497 (N_7497,N_4469,N_5924);
nor U7498 (N_7498,N_4885,N_5342);
and U7499 (N_7499,N_5493,N_4877);
and U7500 (N_7500,N_4303,N_5039);
or U7501 (N_7501,N_5069,N_4503);
and U7502 (N_7502,N_4842,N_5134);
nor U7503 (N_7503,N_5374,N_5842);
nand U7504 (N_7504,N_5186,N_5566);
and U7505 (N_7505,N_4148,N_5478);
nand U7506 (N_7506,N_5004,N_5490);
and U7507 (N_7507,N_5504,N_4707);
or U7508 (N_7508,N_4757,N_5334);
nor U7509 (N_7509,N_4618,N_5928);
nor U7510 (N_7510,N_5242,N_4661);
and U7511 (N_7511,N_5064,N_5946);
nor U7512 (N_7512,N_5852,N_4203);
or U7513 (N_7513,N_4253,N_5582);
nor U7514 (N_7514,N_4202,N_5936);
nor U7515 (N_7515,N_4367,N_4595);
or U7516 (N_7516,N_4567,N_5918);
or U7517 (N_7517,N_4232,N_5628);
nand U7518 (N_7518,N_5903,N_4421);
and U7519 (N_7519,N_5019,N_4566);
and U7520 (N_7520,N_4368,N_5289);
and U7521 (N_7521,N_5648,N_4506);
and U7522 (N_7522,N_5474,N_4306);
or U7523 (N_7523,N_5705,N_4939);
or U7524 (N_7524,N_4565,N_4079);
or U7525 (N_7525,N_5334,N_4432);
nor U7526 (N_7526,N_5873,N_4063);
xor U7527 (N_7527,N_5419,N_4904);
and U7528 (N_7528,N_4217,N_5307);
and U7529 (N_7529,N_4700,N_4246);
nand U7530 (N_7530,N_5865,N_4864);
nand U7531 (N_7531,N_5006,N_5110);
nand U7532 (N_7532,N_4427,N_5065);
and U7533 (N_7533,N_4318,N_5259);
and U7534 (N_7534,N_4614,N_4980);
nor U7535 (N_7535,N_5898,N_4953);
nand U7536 (N_7536,N_4733,N_4869);
nand U7537 (N_7537,N_4736,N_5195);
nand U7538 (N_7538,N_5859,N_5349);
and U7539 (N_7539,N_5480,N_5001);
nand U7540 (N_7540,N_5568,N_5004);
nor U7541 (N_7541,N_4730,N_4064);
and U7542 (N_7542,N_5796,N_4357);
and U7543 (N_7543,N_5328,N_4282);
or U7544 (N_7544,N_4768,N_4504);
or U7545 (N_7545,N_4051,N_5882);
nand U7546 (N_7546,N_5305,N_4031);
nor U7547 (N_7547,N_4357,N_4554);
or U7548 (N_7548,N_4259,N_5480);
or U7549 (N_7549,N_4724,N_5464);
nand U7550 (N_7550,N_5954,N_4365);
and U7551 (N_7551,N_4849,N_5615);
nand U7552 (N_7552,N_5598,N_4853);
or U7553 (N_7553,N_4510,N_5441);
nor U7554 (N_7554,N_5392,N_4005);
nor U7555 (N_7555,N_4769,N_4608);
nor U7556 (N_7556,N_5990,N_5013);
nand U7557 (N_7557,N_4279,N_4732);
and U7558 (N_7558,N_4007,N_4311);
and U7559 (N_7559,N_4813,N_5355);
nand U7560 (N_7560,N_4715,N_4098);
nand U7561 (N_7561,N_5378,N_5653);
and U7562 (N_7562,N_5932,N_5445);
and U7563 (N_7563,N_4879,N_4420);
and U7564 (N_7564,N_5287,N_4506);
nand U7565 (N_7565,N_4448,N_5714);
and U7566 (N_7566,N_5923,N_5361);
or U7567 (N_7567,N_5479,N_4626);
and U7568 (N_7568,N_5107,N_4433);
and U7569 (N_7569,N_5747,N_4842);
nor U7570 (N_7570,N_5994,N_4670);
nor U7571 (N_7571,N_4607,N_5085);
and U7572 (N_7572,N_4313,N_5678);
and U7573 (N_7573,N_4508,N_4390);
nor U7574 (N_7574,N_5307,N_4770);
and U7575 (N_7575,N_5374,N_4848);
or U7576 (N_7576,N_4467,N_4660);
xor U7577 (N_7577,N_4028,N_5984);
nand U7578 (N_7578,N_5816,N_4556);
or U7579 (N_7579,N_5241,N_5102);
nand U7580 (N_7580,N_5400,N_4592);
nor U7581 (N_7581,N_4519,N_5727);
nand U7582 (N_7582,N_4359,N_4634);
or U7583 (N_7583,N_4540,N_4383);
and U7584 (N_7584,N_5696,N_5094);
nand U7585 (N_7585,N_4457,N_5229);
nand U7586 (N_7586,N_5035,N_5862);
nand U7587 (N_7587,N_4836,N_4985);
nand U7588 (N_7588,N_5862,N_4211);
and U7589 (N_7589,N_4659,N_4766);
nand U7590 (N_7590,N_4733,N_5719);
or U7591 (N_7591,N_4861,N_5096);
or U7592 (N_7592,N_5156,N_4222);
or U7593 (N_7593,N_4057,N_4451);
nor U7594 (N_7594,N_4003,N_4327);
and U7595 (N_7595,N_4490,N_5121);
nor U7596 (N_7596,N_5500,N_5145);
and U7597 (N_7597,N_4678,N_4343);
and U7598 (N_7598,N_5334,N_5635);
nor U7599 (N_7599,N_4273,N_4449);
nor U7600 (N_7600,N_4675,N_4823);
nor U7601 (N_7601,N_5823,N_5212);
nor U7602 (N_7602,N_5564,N_4743);
nor U7603 (N_7603,N_5522,N_5104);
and U7604 (N_7604,N_5140,N_5900);
nor U7605 (N_7605,N_5957,N_5684);
nand U7606 (N_7606,N_5337,N_5981);
nand U7607 (N_7607,N_4668,N_5349);
nor U7608 (N_7608,N_4469,N_4126);
nand U7609 (N_7609,N_4649,N_4056);
or U7610 (N_7610,N_4803,N_4331);
or U7611 (N_7611,N_5370,N_4872);
nand U7612 (N_7612,N_4691,N_4082);
nand U7613 (N_7613,N_5551,N_5664);
nor U7614 (N_7614,N_5168,N_5256);
and U7615 (N_7615,N_5715,N_4603);
nand U7616 (N_7616,N_4244,N_4739);
and U7617 (N_7617,N_5737,N_5259);
nor U7618 (N_7618,N_5197,N_5394);
or U7619 (N_7619,N_5631,N_4809);
or U7620 (N_7620,N_5231,N_4193);
nor U7621 (N_7621,N_5909,N_5572);
nor U7622 (N_7622,N_5712,N_4923);
nand U7623 (N_7623,N_4394,N_5094);
and U7624 (N_7624,N_4801,N_5231);
or U7625 (N_7625,N_5719,N_4889);
nor U7626 (N_7626,N_4955,N_5731);
nand U7627 (N_7627,N_4596,N_4236);
or U7628 (N_7628,N_5423,N_4343);
and U7629 (N_7629,N_4389,N_5479);
nand U7630 (N_7630,N_4885,N_5726);
or U7631 (N_7631,N_5106,N_4281);
nor U7632 (N_7632,N_5108,N_4632);
nor U7633 (N_7633,N_5578,N_5643);
and U7634 (N_7634,N_4657,N_5474);
or U7635 (N_7635,N_5465,N_4500);
or U7636 (N_7636,N_4027,N_5057);
or U7637 (N_7637,N_4199,N_5568);
and U7638 (N_7638,N_4061,N_5404);
and U7639 (N_7639,N_4844,N_5240);
nand U7640 (N_7640,N_4357,N_4211);
and U7641 (N_7641,N_5824,N_5866);
and U7642 (N_7642,N_5259,N_4446);
or U7643 (N_7643,N_4875,N_4040);
or U7644 (N_7644,N_5318,N_4364);
nor U7645 (N_7645,N_5428,N_4036);
nor U7646 (N_7646,N_4626,N_4133);
nor U7647 (N_7647,N_4509,N_5957);
nor U7648 (N_7648,N_4594,N_4533);
nor U7649 (N_7649,N_4784,N_5278);
nand U7650 (N_7650,N_4393,N_5328);
nor U7651 (N_7651,N_5971,N_5445);
or U7652 (N_7652,N_5684,N_5289);
nand U7653 (N_7653,N_4005,N_5739);
nor U7654 (N_7654,N_4834,N_4570);
nor U7655 (N_7655,N_5997,N_5707);
xnor U7656 (N_7656,N_5880,N_4978);
and U7657 (N_7657,N_4213,N_5118);
nor U7658 (N_7658,N_5702,N_4246);
nand U7659 (N_7659,N_4169,N_4958);
or U7660 (N_7660,N_5256,N_5046);
nand U7661 (N_7661,N_4609,N_5163);
or U7662 (N_7662,N_5975,N_4114);
nor U7663 (N_7663,N_5030,N_4845);
and U7664 (N_7664,N_4263,N_4491);
nand U7665 (N_7665,N_5178,N_4426);
nor U7666 (N_7666,N_5950,N_5013);
nor U7667 (N_7667,N_5542,N_5483);
or U7668 (N_7668,N_4923,N_5482);
or U7669 (N_7669,N_5174,N_4061);
and U7670 (N_7670,N_5972,N_5683);
nand U7671 (N_7671,N_4913,N_4008);
xnor U7672 (N_7672,N_5793,N_4600);
xor U7673 (N_7673,N_4230,N_5734);
or U7674 (N_7674,N_4014,N_4605);
and U7675 (N_7675,N_4511,N_5550);
and U7676 (N_7676,N_4451,N_5647);
and U7677 (N_7677,N_5971,N_5233);
or U7678 (N_7678,N_5166,N_4119);
and U7679 (N_7679,N_5984,N_5089);
or U7680 (N_7680,N_4968,N_5440);
xnor U7681 (N_7681,N_4390,N_5683);
nand U7682 (N_7682,N_5223,N_5543);
nand U7683 (N_7683,N_4078,N_4192);
nand U7684 (N_7684,N_5894,N_5562);
nor U7685 (N_7685,N_4382,N_4581);
and U7686 (N_7686,N_5764,N_5097);
or U7687 (N_7687,N_4083,N_4917);
and U7688 (N_7688,N_4642,N_5230);
nor U7689 (N_7689,N_5294,N_5078);
nand U7690 (N_7690,N_4993,N_5527);
nand U7691 (N_7691,N_5428,N_5822);
nand U7692 (N_7692,N_4232,N_4110);
nand U7693 (N_7693,N_4170,N_5012);
nor U7694 (N_7694,N_5075,N_4998);
nor U7695 (N_7695,N_4519,N_5370);
nand U7696 (N_7696,N_4300,N_5709);
and U7697 (N_7697,N_5606,N_4388);
and U7698 (N_7698,N_4813,N_5722);
nand U7699 (N_7699,N_4601,N_4201);
or U7700 (N_7700,N_5042,N_4261);
nand U7701 (N_7701,N_4680,N_4245);
or U7702 (N_7702,N_5310,N_4718);
nand U7703 (N_7703,N_4478,N_5985);
xor U7704 (N_7704,N_4149,N_4002);
nor U7705 (N_7705,N_5709,N_5001);
or U7706 (N_7706,N_4388,N_5195);
or U7707 (N_7707,N_5754,N_4476);
and U7708 (N_7708,N_4604,N_4933);
and U7709 (N_7709,N_4994,N_5154);
and U7710 (N_7710,N_4878,N_4796);
or U7711 (N_7711,N_4649,N_5567);
or U7712 (N_7712,N_4265,N_5812);
nand U7713 (N_7713,N_5011,N_4714);
or U7714 (N_7714,N_4733,N_5838);
or U7715 (N_7715,N_4677,N_5501);
or U7716 (N_7716,N_4374,N_5721);
or U7717 (N_7717,N_5149,N_5048);
and U7718 (N_7718,N_4269,N_4934);
and U7719 (N_7719,N_4974,N_4197);
or U7720 (N_7720,N_5538,N_4830);
or U7721 (N_7721,N_4452,N_4731);
nor U7722 (N_7722,N_5108,N_4502);
or U7723 (N_7723,N_4316,N_4515);
nor U7724 (N_7724,N_5192,N_4011);
or U7725 (N_7725,N_5446,N_5476);
or U7726 (N_7726,N_5620,N_5632);
and U7727 (N_7727,N_5874,N_5995);
nand U7728 (N_7728,N_4327,N_4739);
nor U7729 (N_7729,N_5522,N_5685);
nor U7730 (N_7730,N_4394,N_5250);
nor U7731 (N_7731,N_4378,N_5432);
nor U7732 (N_7732,N_5013,N_4231);
or U7733 (N_7733,N_4027,N_4327);
nand U7734 (N_7734,N_5522,N_4432);
nand U7735 (N_7735,N_4090,N_4474);
and U7736 (N_7736,N_4236,N_4109);
nor U7737 (N_7737,N_4377,N_5239);
or U7738 (N_7738,N_5845,N_5100);
nand U7739 (N_7739,N_4001,N_5079);
and U7740 (N_7740,N_4476,N_4080);
nand U7741 (N_7741,N_5342,N_4300);
and U7742 (N_7742,N_5007,N_4569);
and U7743 (N_7743,N_5531,N_5044);
or U7744 (N_7744,N_5371,N_4422);
nand U7745 (N_7745,N_5854,N_4684);
nor U7746 (N_7746,N_4949,N_5748);
nand U7747 (N_7747,N_5488,N_4901);
or U7748 (N_7748,N_5075,N_4651);
nand U7749 (N_7749,N_4715,N_5654);
and U7750 (N_7750,N_4716,N_4527);
nand U7751 (N_7751,N_4491,N_4801);
nor U7752 (N_7752,N_4768,N_5392);
and U7753 (N_7753,N_5276,N_5925);
and U7754 (N_7754,N_5750,N_4697);
or U7755 (N_7755,N_4089,N_5368);
nor U7756 (N_7756,N_4469,N_5530);
and U7757 (N_7757,N_5492,N_5924);
or U7758 (N_7758,N_5209,N_5832);
or U7759 (N_7759,N_5001,N_4751);
nand U7760 (N_7760,N_4260,N_4119);
xor U7761 (N_7761,N_5868,N_5288);
nand U7762 (N_7762,N_4101,N_5152);
and U7763 (N_7763,N_5436,N_4972);
or U7764 (N_7764,N_5158,N_4213);
nor U7765 (N_7765,N_4252,N_4602);
and U7766 (N_7766,N_5922,N_5776);
nor U7767 (N_7767,N_4146,N_4139);
and U7768 (N_7768,N_4753,N_5939);
nand U7769 (N_7769,N_5906,N_5963);
nand U7770 (N_7770,N_4303,N_5830);
and U7771 (N_7771,N_5683,N_5699);
or U7772 (N_7772,N_5085,N_5150);
nand U7773 (N_7773,N_4913,N_5208);
nor U7774 (N_7774,N_4247,N_5296);
and U7775 (N_7775,N_4053,N_5696);
and U7776 (N_7776,N_4167,N_5965);
nor U7777 (N_7777,N_5423,N_5186);
or U7778 (N_7778,N_5282,N_5201);
or U7779 (N_7779,N_4466,N_5698);
nand U7780 (N_7780,N_4296,N_5778);
nor U7781 (N_7781,N_5487,N_5016);
nand U7782 (N_7782,N_4923,N_5890);
or U7783 (N_7783,N_5807,N_4796);
nand U7784 (N_7784,N_5882,N_4084);
nor U7785 (N_7785,N_4504,N_5078);
nand U7786 (N_7786,N_5955,N_5726);
and U7787 (N_7787,N_4301,N_5990);
or U7788 (N_7788,N_4878,N_4341);
or U7789 (N_7789,N_4365,N_5025);
nand U7790 (N_7790,N_5183,N_5176);
nor U7791 (N_7791,N_4986,N_4932);
nand U7792 (N_7792,N_5901,N_4302);
nor U7793 (N_7793,N_4813,N_5132);
nor U7794 (N_7794,N_5323,N_4663);
nand U7795 (N_7795,N_4632,N_5334);
nor U7796 (N_7796,N_5764,N_5953);
and U7797 (N_7797,N_4998,N_5039);
nor U7798 (N_7798,N_4762,N_4354);
nand U7799 (N_7799,N_4592,N_5662);
xnor U7800 (N_7800,N_5557,N_5505);
nor U7801 (N_7801,N_5582,N_4840);
or U7802 (N_7802,N_4930,N_5372);
nor U7803 (N_7803,N_5464,N_5640);
and U7804 (N_7804,N_5092,N_4375);
nor U7805 (N_7805,N_5526,N_5814);
nand U7806 (N_7806,N_5403,N_4457);
and U7807 (N_7807,N_4608,N_5940);
nand U7808 (N_7808,N_4237,N_4492);
nand U7809 (N_7809,N_5460,N_5063);
nand U7810 (N_7810,N_5674,N_4005);
or U7811 (N_7811,N_4027,N_4476);
or U7812 (N_7812,N_5980,N_4218);
and U7813 (N_7813,N_5740,N_5660);
and U7814 (N_7814,N_4976,N_4761);
and U7815 (N_7815,N_4675,N_5371);
nor U7816 (N_7816,N_5748,N_4918);
and U7817 (N_7817,N_4262,N_4593);
or U7818 (N_7818,N_4789,N_5618);
nand U7819 (N_7819,N_4536,N_5860);
and U7820 (N_7820,N_5030,N_4467);
or U7821 (N_7821,N_4496,N_4779);
or U7822 (N_7822,N_5097,N_5074);
nand U7823 (N_7823,N_4028,N_5278);
nor U7824 (N_7824,N_5291,N_4465);
or U7825 (N_7825,N_5901,N_4136);
nand U7826 (N_7826,N_4396,N_4451);
nor U7827 (N_7827,N_4277,N_4632);
nand U7828 (N_7828,N_5479,N_4790);
nor U7829 (N_7829,N_5033,N_5031);
nor U7830 (N_7830,N_5749,N_5418);
nor U7831 (N_7831,N_4575,N_5156);
or U7832 (N_7832,N_4625,N_4823);
or U7833 (N_7833,N_5552,N_5005);
nor U7834 (N_7834,N_4562,N_5231);
nor U7835 (N_7835,N_5977,N_4874);
nand U7836 (N_7836,N_4625,N_5727);
nand U7837 (N_7837,N_5386,N_5721);
nor U7838 (N_7838,N_5253,N_5231);
nand U7839 (N_7839,N_5340,N_5628);
nor U7840 (N_7840,N_4343,N_5642);
xnor U7841 (N_7841,N_5020,N_4769);
and U7842 (N_7842,N_5954,N_5281);
nand U7843 (N_7843,N_5925,N_4492);
nor U7844 (N_7844,N_5703,N_4017);
nand U7845 (N_7845,N_5302,N_5373);
nor U7846 (N_7846,N_4785,N_4206);
nor U7847 (N_7847,N_4148,N_5132);
nand U7848 (N_7848,N_5973,N_5234);
and U7849 (N_7849,N_5216,N_4160);
or U7850 (N_7850,N_4017,N_5139);
or U7851 (N_7851,N_4551,N_5140);
nand U7852 (N_7852,N_5014,N_5284);
nand U7853 (N_7853,N_5379,N_5309);
or U7854 (N_7854,N_4567,N_5846);
nor U7855 (N_7855,N_4011,N_5396);
nand U7856 (N_7856,N_5670,N_5391);
and U7857 (N_7857,N_5101,N_4751);
nand U7858 (N_7858,N_5556,N_5515);
or U7859 (N_7859,N_5529,N_4150);
or U7860 (N_7860,N_4820,N_5410);
nand U7861 (N_7861,N_4134,N_4841);
or U7862 (N_7862,N_4955,N_5334);
and U7863 (N_7863,N_4107,N_4587);
and U7864 (N_7864,N_4580,N_5677);
nor U7865 (N_7865,N_4578,N_4868);
and U7866 (N_7866,N_4638,N_5343);
nor U7867 (N_7867,N_5657,N_5027);
xor U7868 (N_7868,N_4340,N_5985);
or U7869 (N_7869,N_5619,N_5900);
and U7870 (N_7870,N_5060,N_5952);
or U7871 (N_7871,N_4831,N_5929);
or U7872 (N_7872,N_5113,N_5359);
nand U7873 (N_7873,N_5657,N_4205);
and U7874 (N_7874,N_4013,N_4745);
nand U7875 (N_7875,N_5857,N_4277);
or U7876 (N_7876,N_4202,N_5438);
and U7877 (N_7877,N_4580,N_5137);
nor U7878 (N_7878,N_4333,N_4493);
nand U7879 (N_7879,N_5468,N_5913);
or U7880 (N_7880,N_4475,N_5895);
or U7881 (N_7881,N_4498,N_5769);
nand U7882 (N_7882,N_5560,N_4317);
and U7883 (N_7883,N_5176,N_4971);
nor U7884 (N_7884,N_4708,N_5685);
and U7885 (N_7885,N_4595,N_5837);
or U7886 (N_7886,N_5646,N_4143);
and U7887 (N_7887,N_4179,N_5268);
and U7888 (N_7888,N_4419,N_4168);
or U7889 (N_7889,N_4449,N_5679);
or U7890 (N_7890,N_5340,N_5249);
nor U7891 (N_7891,N_5144,N_4895);
xor U7892 (N_7892,N_5897,N_5197);
nand U7893 (N_7893,N_4661,N_4976);
xnor U7894 (N_7894,N_5413,N_4052);
or U7895 (N_7895,N_5754,N_4235);
nor U7896 (N_7896,N_5533,N_5537);
or U7897 (N_7897,N_4979,N_4288);
nand U7898 (N_7898,N_5057,N_4180);
and U7899 (N_7899,N_5855,N_4395);
nor U7900 (N_7900,N_4334,N_5858);
nor U7901 (N_7901,N_5185,N_5094);
and U7902 (N_7902,N_5979,N_5301);
nor U7903 (N_7903,N_4091,N_4305);
or U7904 (N_7904,N_4689,N_5734);
nor U7905 (N_7905,N_5805,N_4714);
and U7906 (N_7906,N_5596,N_4569);
xnor U7907 (N_7907,N_5206,N_5230);
nor U7908 (N_7908,N_5302,N_4471);
nor U7909 (N_7909,N_5431,N_5107);
and U7910 (N_7910,N_5244,N_5605);
nor U7911 (N_7911,N_5752,N_5709);
nand U7912 (N_7912,N_4035,N_5692);
and U7913 (N_7913,N_5644,N_5535);
nand U7914 (N_7914,N_5377,N_5903);
nor U7915 (N_7915,N_4400,N_5981);
nor U7916 (N_7916,N_4272,N_5272);
nor U7917 (N_7917,N_4278,N_5387);
and U7918 (N_7918,N_5611,N_5827);
and U7919 (N_7919,N_5987,N_4615);
nand U7920 (N_7920,N_5350,N_4569);
and U7921 (N_7921,N_4896,N_5539);
nand U7922 (N_7922,N_5133,N_4756);
nand U7923 (N_7923,N_4341,N_5038);
or U7924 (N_7924,N_5739,N_5654);
nor U7925 (N_7925,N_4325,N_4552);
nor U7926 (N_7926,N_4079,N_4076);
nand U7927 (N_7927,N_5748,N_5407);
nor U7928 (N_7928,N_5693,N_4938);
nand U7929 (N_7929,N_4531,N_4195);
nand U7930 (N_7930,N_4780,N_4924);
nor U7931 (N_7931,N_5242,N_5600);
and U7932 (N_7932,N_4041,N_5767);
xor U7933 (N_7933,N_5534,N_5299);
or U7934 (N_7934,N_4985,N_4609);
and U7935 (N_7935,N_4311,N_5132);
nand U7936 (N_7936,N_5732,N_4777);
and U7937 (N_7937,N_4712,N_5523);
or U7938 (N_7938,N_5642,N_4473);
or U7939 (N_7939,N_5383,N_4719);
nand U7940 (N_7940,N_5656,N_4794);
nand U7941 (N_7941,N_5044,N_4363);
nand U7942 (N_7942,N_4027,N_5604);
nand U7943 (N_7943,N_4897,N_5919);
or U7944 (N_7944,N_4423,N_4349);
and U7945 (N_7945,N_5458,N_4442);
nand U7946 (N_7946,N_4223,N_4180);
and U7947 (N_7947,N_4215,N_5969);
or U7948 (N_7948,N_5506,N_4602);
nand U7949 (N_7949,N_5324,N_4916);
and U7950 (N_7950,N_5689,N_4238);
xnor U7951 (N_7951,N_4365,N_5132);
nor U7952 (N_7952,N_4696,N_4446);
and U7953 (N_7953,N_5143,N_5040);
nor U7954 (N_7954,N_4373,N_5503);
or U7955 (N_7955,N_5521,N_5014);
or U7956 (N_7956,N_5584,N_5289);
nor U7957 (N_7957,N_4733,N_4011);
or U7958 (N_7958,N_5947,N_5346);
or U7959 (N_7959,N_4910,N_4419);
and U7960 (N_7960,N_5397,N_4930);
and U7961 (N_7961,N_4097,N_5119);
nor U7962 (N_7962,N_5964,N_4333);
nor U7963 (N_7963,N_4681,N_5578);
xor U7964 (N_7964,N_4563,N_5300);
nor U7965 (N_7965,N_4187,N_5422);
nor U7966 (N_7966,N_4358,N_4767);
and U7967 (N_7967,N_4401,N_4553);
or U7968 (N_7968,N_5578,N_4150);
nor U7969 (N_7969,N_5549,N_4835);
and U7970 (N_7970,N_5891,N_4897);
nand U7971 (N_7971,N_4672,N_5723);
or U7972 (N_7972,N_4783,N_4845);
nand U7973 (N_7973,N_4323,N_5462);
nor U7974 (N_7974,N_5138,N_5912);
or U7975 (N_7975,N_5422,N_5876);
or U7976 (N_7976,N_5188,N_5337);
and U7977 (N_7977,N_5191,N_5397);
and U7978 (N_7978,N_5430,N_4097);
or U7979 (N_7979,N_4978,N_4019);
nand U7980 (N_7980,N_4506,N_5653);
nand U7981 (N_7981,N_4222,N_4563);
xnor U7982 (N_7982,N_4259,N_5424);
nor U7983 (N_7983,N_4569,N_4947);
and U7984 (N_7984,N_5333,N_5409);
nand U7985 (N_7985,N_5820,N_4573);
nor U7986 (N_7986,N_5164,N_5636);
and U7987 (N_7987,N_5629,N_4897);
nand U7988 (N_7988,N_5874,N_4820);
or U7989 (N_7989,N_5647,N_5226);
nand U7990 (N_7990,N_4317,N_5456);
and U7991 (N_7991,N_4555,N_5593);
nand U7992 (N_7992,N_4507,N_5121);
or U7993 (N_7993,N_4575,N_5953);
and U7994 (N_7994,N_5416,N_5926);
nor U7995 (N_7995,N_4949,N_4167);
or U7996 (N_7996,N_4945,N_4995);
nor U7997 (N_7997,N_5023,N_5402);
and U7998 (N_7998,N_4050,N_5265);
and U7999 (N_7999,N_5880,N_4772);
nand U8000 (N_8000,N_6780,N_7326);
nor U8001 (N_8001,N_7204,N_6089);
nand U8002 (N_8002,N_7580,N_6087);
xnor U8003 (N_8003,N_6139,N_7633);
and U8004 (N_8004,N_6913,N_7291);
nand U8005 (N_8005,N_7346,N_7160);
or U8006 (N_8006,N_7371,N_6372);
and U8007 (N_8007,N_7313,N_7329);
or U8008 (N_8008,N_6324,N_7208);
nor U8009 (N_8009,N_7861,N_7819);
or U8010 (N_8010,N_7450,N_6597);
nand U8011 (N_8011,N_7288,N_6776);
or U8012 (N_8012,N_7853,N_6393);
or U8013 (N_8013,N_7140,N_6265);
or U8014 (N_8014,N_6009,N_6959);
and U8015 (N_8015,N_6330,N_7395);
nand U8016 (N_8016,N_7424,N_6226);
nand U8017 (N_8017,N_7079,N_7656);
and U8018 (N_8018,N_6269,N_7597);
nand U8019 (N_8019,N_6351,N_6361);
and U8020 (N_8020,N_7068,N_6564);
or U8021 (N_8021,N_7579,N_6063);
xor U8022 (N_8022,N_6537,N_6478);
nor U8023 (N_8023,N_6266,N_7728);
nand U8024 (N_8024,N_7862,N_6876);
nor U8025 (N_8025,N_6108,N_6604);
nor U8026 (N_8026,N_7349,N_6781);
nand U8027 (N_8027,N_7891,N_6456);
nand U8028 (N_8028,N_6504,N_7441);
nand U8029 (N_8029,N_7363,N_6156);
and U8030 (N_8030,N_7578,N_7784);
nor U8031 (N_8031,N_6484,N_6255);
nor U8032 (N_8032,N_6539,N_7671);
nor U8033 (N_8033,N_6020,N_7024);
or U8034 (N_8034,N_7178,N_6169);
or U8035 (N_8035,N_6841,N_7296);
or U8036 (N_8036,N_7158,N_7331);
nor U8037 (N_8037,N_7487,N_7546);
nand U8038 (N_8038,N_7491,N_6948);
nor U8039 (N_8039,N_7351,N_6662);
or U8040 (N_8040,N_7110,N_7096);
nor U8041 (N_8041,N_7589,N_7634);
and U8042 (N_8042,N_6785,N_7867);
nor U8043 (N_8043,N_7593,N_7167);
and U8044 (N_8044,N_6856,N_7482);
nand U8045 (N_8045,N_6234,N_7956);
or U8046 (N_8046,N_7653,N_7754);
nor U8047 (N_8047,N_7590,N_6793);
nor U8048 (N_8048,N_6246,N_7301);
nand U8049 (N_8049,N_7536,N_6096);
nor U8050 (N_8050,N_6782,N_7198);
and U8051 (N_8051,N_6652,N_7774);
or U8052 (N_8052,N_6617,N_7155);
and U8053 (N_8053,N_6395,N_7129);
xor U8054 (N_8054,N_6445,N_7782);
nand U8055 (N_8055,N_7674,N_6195);
nand U8056 (N_8056,N_6198,N_7779);
nand U8057 (N_8057,N_7503,N_7021);
nor U8058 (N_8058,N_6526,N_6424);
nor U8059 (N_8059,N_7695,N_7071);
nand U8060 (N_8060,N_7391,N_6495);
or U8061 (N_8061,N_7324,N_7289);
nor U8062 (N_8062,N_6595,N_6531);
xnor U8063 (N_8063,N_7666,N_6426);
or U8064 (N_8064,N_6520,N_7554);
nor U8065 (N_8065,N_7984,N_7412);
nor U8066 (N_8066,N_7568,N_7176);
nand U8067 (N_8067,N_7628,N_7881);
nor U8068 (N_8068,N_6575,N_6306);
nor U8069 (N_8069,N_7105,N_6006);
nor U8070 (N_8070,N_6568,N_7910);
nor U8071 (N_8071,N_7453,N_7623);
nor U8072 (N_8072,N_6873,N_7494);
nor U8073 (N_8073,N_6134,N_6955);
or U8074 (N_8074,N_6309,N_6586);
and U8075 (N_8075,N_7271,N_6251);
nand U8076 (N_8076,N_6362,N_7355);
nor U8077 (N_8077,N_7828,N_7461);
or U8078 (N_8078,N_7547,N_6899);
or U8079 (N_8079,N_6143,N_6055);
nand U8080 (N_8080,N_7283,N_6429);
or U8081 (N_8081,N_7570,N_6416);
or U8082 (N_8082,N_6190,N_7928);
nand U8083 (N_8083,N_6705,N_6562);
and U8084 (N_8084,N_7997,N_7419);
or U8085 (N_8085,N_7660,N_7452);
nand U8086 (N_8086,N_6485,N_7814);
or U8087 (N_8087,N_7768,N_7272);
nor U8088 (N_8088,N_7255,N_7353);
or U8089 (N_8089,N_6852,N_6256);
or U8090 (N_8090,N_7733,N_6970);
and U8091 (N_8091,N_6216,N_6584);
nor U8092 (N_8092,N_6350,N_7918);
or U8093 (N_8093,N_6165,N_6448);
and U8094 (N_8094,N_7221,N_7852);
nor U8095 (N_8095,N_7912,N_6197);
nand U8096 (N_8096,N_6206,N_7875);
or U8097 (N_8097,N_6925,N_7199);
and U8098 (N_8098,N_6798,N_6936);
nor U8099 (N_8099,N_7892,N_7937);
or U8100 (N_8100,N_6942,N_7783);
xnor U8101 (N_8101,N_6675,N_7599);
or U8102 (N_8102,N_6104,N_6867);
and U8103 (N_8103,N_7745,N_6649);
or U8104 (N_8104,N_7507,N_6613);
nand U8105 (N_8105,N_6267,N_6308);
xnor U8106 (N_8106,N_6981,N_6039);
and U8107 (N_8107,N_7835,N_7818);
and U8108 (N_8108,N_7934,N_6137);
nand U8109 (N_8109,N_6072,N_6455);
nor U8110 (N_8110,N_6561,N_7392);
or U8111 (N_8111,N_6240,N_6446);
and U8112 (N_8112,N_6615,N_6797);
nand U8113 (N_8113,N_7330,N_6807);
nand U8114 (N_8114,N_7126,N_6703);
nand U8115 (N_8115,N_7793,N_7706);
nand U8116 (N_8116,N_6067,N_7484);
or U8117 (N_8117,N_7517,N_6033);
and U8118 (N_8118,N_6605,N_6287);
or U8119 (N_8119,N_7583,N_6441);
nor U8120 (N_8120,N_7926,N_7707);
nor U8121 (N_8121,N_7145,N_6706);
nor U8122 (N_8122,N_6657,N_6228);
nand U8123 (N_8123,N_6976,N_7498);
nand U8124 (N_8124,N_6522,N_6032);
or U8125 (N_8125,N_6721,N_7383);
or U8126 (N_8126,N_6378,N_6784);
or U8127 (N_8127,N_7552,N_6634);
nor U8128 (N_8128,N_6930,N_7943);
nand U8129 (N_8129,N_7239,N_6203);
or U8130 (N_8130,N_6028,N_6326);
nor U8131 (N_8131,N_6843,N_6607);
or U8132 (N_8132,N_6903,N_6535);
nor U8133 (N_8133,N_7615,N_6822);
nand U8134 (N_8134,N_6693,N_7059);
and U8135 (N_8135,N_7955,N_6835);
nor U8136 (N_8136,N_7254,N_6133);
nor U8137 (N_8137,N_6831,N_6029);
and U8138 (N_8138,N_6659,N_7033);
or U8139 (N_8139,N_7090,N_7977);
nor U8140 (N_8140,N_6406,N_6789);
nor U8141 (N_8141,N_7462,N_6052);
and U8142 (N_8142,N_6842,N_7716);
nand U8143 (N_8143,N_6518,N_6479);
or U8144 (N_8144,N_6099,N_6453);
or U8145 (N_8145,N_6892,N_6689);
nor U8146 (N_8146,N_7212,N_7222);
or U8147 (N_8147,N_6650,N_6130);
and U8148 (N_8148,N_7763,N_7545);
and U8149 (N_8149,N_7605,N_7323);
nor U8150 (N_8150,N_7258,N_6210);
nand U8151 (N_8151,N_6157,N_7164);
and U8152 (N_8152,N_7177,N_7640);
and U8153 (N_8153,N_7531,N_7407);
or U8154 (N_8154,N_6428,N_7135);
and U8155 (N_8155,N_6297,N_6548);
or U8156 (N_8156,N_7297,N_6149);
or U8157 (N_8157,N_7719,N_7738);
and U8158 (N_8158,N_6180,N_6179);
or U8159 (N_8159,N_7979,N_7084);
or U8160 (N_8160,N_7118,N_7659);
or U8161 (N_8161,N_6219,N_7172);
nand U8162 (N_8162,N_6400,N_7099);
or U8163 (N_8163,N_7304,N_6624);
nand U8164 (N_8164,N_7077,N_7809);
and U8165 (N_8165,N_7932,N_6944);
nor U8166 (N_8166,N_6836,N_7005);
and U8167 (N_8167,N_6223,N_6606);
or U8168 (N_8168,N_6191,N_7729);
nor U8169 (N_8169,N_6128,N_7527);
nor U8170 (N_8170,N_7770,N_6722);
nand U8171 (N_8171,N_7534,N_6321);
nand U8172 (N_8172,N_7134,N_7566);
and U8173 (N_8173,N_6150,N_7974);
or U8174 (N_8174,N_7053,N_6685);
and U8175 (N_8175,N_6305,N_6972);
nand U8176 (N_8176,N_7944,N_7133);
or U8177 (N_8177,N_6135,N_6608);
nor U8178 (N_8178,N_6720,N_7231);
or U8179 (N_8179,N_7332,N_6768);
nor U8180 (N_8180,N_6473,N_7121);
nand U8181 (N_8181,N_6550,N_6603);
nand U8182 (N_8182,N_7730,N_7540);
nand U8183 (N_8183,N_7844,N_7714);
nor U8184 (N_8184,N_6227,N_6519);
or U8185 (N_8185,N_6475,N_6728);
and U8186 (N_8186,N_6771,N_6735);
nand U8187 (N_8187,N_7769,N_7207);
or U8188 (N_8188,N_6923,N_6048);
nand U8189 (N_8189,N_7696,N_7182);
nor U8190 (N_8190,N_6639,N_7665);
nor U8191 (N_8191,N_7873,N_7505);
or U8192 (N_8192,N_7613,N_7797);
and U8193 (N_8193,N_7264,N_7420);
nand U8194 (N_8194,N_7841,N_7490);
or U8195 (N_8195,N_6060,N_7905);
and U8196 (N_8196,N_6314,N_6431);
nor U8197 (N_8197,N_6742,N_7334);
nor U8198 (N_8198,N_6885,N_7286);
or U8199 (N_8199,N_7107,N_6779);
nor U8200 (N_8200,N_7617,N_6958);
and U8201 (N_8201,N_6224,N_7029);
and U8202 (N_8202,N_7727,N_6168);
nor U8203 (N_8203,N_7193,N_6131);
and U8204 (N_8204,N_6820,N_7376);
nor U8205 (N_8205,N_6816,N_7495);
or U8206 (N_8206,N_7691,N_7180);
and U8207 (N_8207,N_6295,N_7646);
nand U8208 (N_8208,N_7661,N_7043);
or U8209 (N_8209,N_6275,N_7612);
or U8210 (N_8210,N_6369,N_7981);
nand U8211 (N_8211,N_6310,N_6941);
and U8212 (N_8212,N_6552,N_7935);
and U8213 (N_8213,N_7279,N_7447);
nor U8214 (N_8214,N_7806,N_7522);
and U8215 (N_8215,N_7576,N_6381);
or U8216 (N_8216,N_6532,N_7973);
or U8217 (N_8217,N_7645,N_6946);
nand U8218 (N_8218,N_6846,N_6124);
nor U8219 (N_8219,N_6962,N_6402);
and U8220 (N_8220,N_7183,N_6623);
or U8221 (N_8221,N_7972,N_7907);
nor U8222 (N_8222,N_6702,N_6949);
nand U8223 (N_8223,N_6733,N_6025);
nand U8224 (N_8224,N_6364,N_7202);
or U8225 (N_8225,N_7585,N_6138);
and U8226 (N_8226,N_7734,N_7845);
nor U8227 (N_8227,N_7992,N_7149);
and U8228 (N_8228,N_6422,N_7667);
nand U8229 (N_8229,N_6368,N_7139);
or U8230 (N_8230,N_6963,N_6126);
nand U8231 (N_8231,N_7606,N_6337);
nor U8232 (N_8232,N_6682,N_7896);
or U8233 (N_8233,N_6098,N_6817);
nor U8234 (N_8234,N_6286,N_7889);
nand U8235 (N_8235,N_7868,N_7871);
nor U8236 (N_8236,N_7810,N_6500);
nor U8237 (N_8237,N_7650,N_6420);
and U8238 (N_8238,N_7378,N_7312);
nand U8239 (N_8239,N_6917,N_6580);
xor U8240 (N_8240,N_6747,N_7635);
or U8241 (N_8241,N_7314,N_7037);
and U8242 (N_8242,N_7532,N_6984);
nor U8243 (N_8243,N_7595,N_7725);
or U8244 (N_8244,N_7169,N_6759);
nand U8245 (N_8245,N_7776,N_6411);
and U8246 (N_8246,N_6902,N_6289);
or U8247 (N_8247,N_6523,N_7842);
and U8248 (N_8248,N_7712,N_6524);
and U8249 (N_8249,N_7676,N_6094);
nand U8250 (N_8250,N_6392,N_7808);
or U8251 (N_8251,N_7571,N_7075);
nor U8252 (N_8252,N_6794,N_7632);
nor U8253 (N_8253,N_7726,N_7048);
nand U8254 (N_8254,N_7700,N_6463);
nor U8255 (N_8255,N_7924,N_7902);
nand U8256 (N_8256,N_7173,N_6663);
and U8257 (N_8257,N_7270,N_6494);
nor U8258 (N_8258,N_7216,N_6013);
nand U8259 (N_8259,N_7409,N_6574);
and U8260 (N_8260,N_7227,N_6185);
or U8261 (N_8261,N_6172,N_6756);
nand U8262 (N_8262,N_7174,N_7601);
nor U8263 (N_8263,N_7752,N_6989);
and U8264 (N_8264,N_6937,N_6648);
and U8265 (N_8265,N_6935,N_7639);
and U8266 (N_8266,N_7524,N_6920);
nand U8267 (N_8267,N_6427,N_6162);
nor U8268 (N_8268,N_7120,N_6491);
and U8269 (N_8269,N_6074,N_7614);
xnor U8270 (N_8270,N_7865,N_6430);
and U8271 (N_8271,N_7829,N_6881);
and U8272 (N_8272,N_6090,N_6610);
and U8273 (N_8273,N_6398,N_6601);
and U8274 (N_8274,N_6215,N_6417);
xnor U8275 (N_8275,N_6960,N_6696);
nand U8276 (N_8276,N_6612,N_7751);
nand U8277 (N_8277,N_6844,N_7826);
or U8278 (N_8278,N_7884,N_7663);
nand U8279 (N_8279,N_7074,N_7057);
or U8280 (N_8280,N_7234,N_6977);
xnor U8281 (N_8281,N_6818,N_7125);
and U8282 (N_8282,N_7338,N_7022);
or U8283 (N_8283,N_7906,N_7306);
nand U8284 (N_8284,N_7781,N_6540);
or U8285 (N_8285,N_6184,N_7577);
and U8286 (N_8286,N_7011,N_7750);
xor U8287 (N_8287,N_7106,N_6196);
or U8288 (N_8288,N_6085,N_7224);
nor U8289 (N_8289,N_6263,N_7115);
and U8290 (N_8290,N_6670,N_6783);
and U8291 (N_8291,N_6283,N_6775);
and U8292 (N_8292,N_6405,N_6750);
nand U8293 (N_8293,N_7230,N_7559);
nand U8294 (N_8294,N_6071,N_6837);
nor U8295 (N_8295,N_7898,N_7122);
and U8296 (N_8296,N_7220,N_6510);
nor U8297 (N_8297,N_7654,N_7235);
and U8298 (N_8298,N_6027,N_6258);
nand U8299 (N_8299,N_7062,N_6152);
nand U8300 (N_8300,N_6515,N_6008);
or U8301 (N_8301,N_6987,N_6023);
or U8302 (N_8302,N_6298,N_7916);
or U8303 (N_8303,N_6585,N_7909);
and U8304 (N_8304,N_7007,N_7496);
nor U8305 (N_8305,N_7697,N_6672);
xnor U8306 (N_8306,N_7539,N_7843);
nand U8307 (N_8307,N_6905,N_7015);
and U8308 (N_8308,N_7066,N_7367);
and U8309 (N_8309,N_6752,N_7146);
nor U8310 (N_8310,N_6095,N_7170);
nand U8311 (N_8311,N_6651,N_7247);
and U8312 (N_8312,N_6912,N_6854);
or U8313 (N_8313,N_6450,N_7433);
nand U8314 (N_8314,N_6017,N_7526);
nor U8315 (N_8315,N_6285,N_7919);
or U8316 (N_8316,N_7374,N_7214);
and U8317 (N_8317,N_6953,N_7192);
nand U8318 (N_8318,N_7786,N_7294);
and U8319 (N_8319,N_6501,N_6080);
or U8320 (N_8320,N_6932,N_7815);
and U8321 (N_8321,N_6155,N_7631);
nand U8322 (N_8322,N_7347,N_6331);
and U8323 (N_8323,N_6916,N_6254);
or U8324 (N_8324,N_7563,N_7194);
or U8325 (N_8325,N_6301,N_6145);
nor U8326 (N_8326,N_7701,N_7856);
xor U8327 (N_8327,N_6810,N_6377);
and U8328 (N_8328,N_7269,N_6909);
and U8329 (N_8329,N_7248,N_6734);
nand U8330 (N_8330,N_6581,N_6767);
and U8331 (N_8331,N_7885,N_7893);
and U8332 (N_8332,N_7791,N_6993);
nor U8333 (N_8333,N_6587,N_6105);
xor U8334 (N_8334,N_6965,N_7747);
and U8335 (N_8335,N_6231,N_6778);
nor U8336 (N_8336,N_7780,N_7483);
and U8337 (N_8337,N_6622,N_7930);
nand U8338 (N_8338,N_6154,N_7673);
nand U8339 (N_8339,N_7850,N_7915);
and U8340 (N_8340,N_6863,N_6824);
or U8341 (N_8341,N_6700,N_6387);
or U8342 (N_8342,N_7245,N_6140);
or U8343 (N_8343,N_6961,N_6665);
nand U8344 (N_8344,N_6966,N_6037);
nand U8345 (N_8345,N_7732,N_7390);
and U8346 (N_8346,N_6897,N_6273);
nand U8347 (N_8347,N_6808,N_6760);
and U8348 (N_8348,N_7113,N_7558);
nor U8349 (N_8349,N_7644,N_6712);
or U8350 (N_8350,N_7764,N_7280);
nor U8351 (N_8351,N_7000,N_7510);
and U8352 (N_8352,N_6503,N_6765);
and U8353 (N_8353,N_6732,N_7200);
or U8354 (N_8354,N_7693,N_7410);
nand U8355 (N_8355,N_7888,N_6744);
or U8356 (N_8356,N_6952,N_6136);
and U8357 (N_8357,N_6001,N_7813);
nand U8358 (N_8358,N_7816,N_6870);
or U8359 (N_8359,N_7963,N_6697);
xnor U8360 (N_8360,N_7088,N_7460);
nand U8361 (N_8361,N_6329,N_7857);
and U8362 (N_8362,N_7765,N_6718);
or U8363 (N_8363,N_6829,N_6667);
and U8364 (N_8364,N_7012,N_6076);
or U8365 (N_8365,N_6466,N_7243);
and U8366 (N_8366,N_6158,N_7851);
nor U8367 (N_8367,N_6117,N_7310);
and U8368 (N_8368,N_6147,N_6741);
nand U8369 (N_8369,N_7249,N_6316);
nor U8370 (N_8370,N_7056,N_6928);
nand U8371 (N_8371,N_7569,N_7073);
nand U8372 (N_8372,N_7166,N_6051);
and U8373 (N_8373,N_6279,N_7587);
and U8374 (N_8374,N_6262,N_6882);
nand U8375 (N_8375,N_7013,N_7352);
and U8376 (N_8376,N_7027,N_6694);
nand U8377 (N_8377,N_7790,N_6618);
and U8378 (N_8378,N_6739,N_6790);
and U8379 (N_8379,N_7834,N_7445);
and U8380 (N_8380,N_6969,N_7394);
nor U8381 (N_8381,N_7672,N_7238);
nand U8382 (N_8382,N_7290,N_7058);
nand U8383 (N_8383,N_6823,N_6338);
or U8384 (N_8384,N_7381,N_7171);
nand U8385 (N_8385,N_6806,N_7070);
nand U8386 (N_8386,N_6100,N_6115);
or U8387 (N_8387,N_6452,N_6677);
and U8388 (N_8388,N_6483,N_6040);
nand U8389 (N_8389,N_6214,N_6508);
nand U8390 (N_8390,N_7377,N_7308);
and U8391 (N_8391,N_6260,N_6218);
or U8392 (N_8392,N_6986,N_6335);
nor U8393 (N_8393,N_7025,N_7685);
or U8394 (N_8394,N_7699,N_7690);
and U8395 (N_8395,N_7602,N_6724);
nand U8396 (N_8396,N_6443,N_7803);
nor U8397 (N_8397,N_6035,N_7575);
nand U8398 (N_8398,N_7050,N_7993);
or U8399 (N_8399,N_6924,N_7114);
and U8400 (N_8400,N_7508,N_6645);
nor U8401 (N_8401,N_6904,N_6014);
and U8402 (N_8402,N_7925,N_7513);
nor U8403 (N_8403,N_7209,N_7807);
or U8404 (N_8404,N_7282,N_7939);
nand U8405 (N_8405,N_7603,N_7237);
and U8406 (N_8406,N_6571,N_6795);
xor U8407 (N_8407,N_6288,N_7836);
or U8408 (N_8408,N_6695,N_6110);
nor U8409 (N_8409,N_6166,N_6509);
nand U8410 (N_8410,N_7703,N_7225);
nand U8411 (N_8411,N_6281,N_6636);
and U8412 (N_8412,N_7913,N_7922);
nand U8413 (N_8413,N_6069,N_7232);
nor U8414 (N_8414,N_6159,N_7041);
or U8415 (N_8415,N_6643,N_6872);
and U8416 (N_8416,N_7970,N_6878);
nor U8417 (N_8417,N_7983,N_6049);
and U8418 (N_8418,N_7165,N_6865);
nor U8419 (N_8419,N_7968,N_7863);
or U8420 (N_8420,N_7159,N_6628);
and U8421 (N_8421,N_7018,N_6235);
and U8422 (N_8422,N_7380,N_7434);
nor U8423 (N_8423,N_7092,N_6527);
or U8424 (N_8424,N_7327,N_6352);
xnor U8425 (N_8425,N_6171,N_6058);
nor U8426 (N_8426,N_7138,N_6077);
or U8427 (N_8427,N_7211,N_7206);
nand U8428 (N_8428,N_7362,N_6187);
nand U8429 (N_8429,N_7933,N_7448);
nand U8430 (N_8430,N_7649,N_6259);
nand U8431 (N_8431,N_7111,N_6056);
nand U8432 (N_8432,N_7564,N_6304);
or U8433 (N_8433,N_7257,N_7026);
or U8434 (N_8434,N_6188,N_6481);
nand U8435 (N_8435,N_6850,N_6918);
nand U8436 (N_8436,N_7273,N_7422);
nor U8437 (N_8437,N_6082,N_6701);
nor U8438 (N_8438,N_6474,N_7032);
or U8439 (N_8439,N_6546,N_7455);
or U8440 (N_8440,N_6717,N_6616);
or U8441 (N_8441,N_7415,N_7426);
nor U8442 (N_8442,N_6079,N_7343);
nor U8443 (N_8443,N_6896,N_6141);
or U8444 (N_8444,N_6861,N_6553);
nor U8445 (N_8445,N_6536,N_7303);
or U8446 (N_8446,N_6974,N_7824);
and U8447 (N_8447,N_6176,N_6011);
nand U8448 (N_8448,N_6342,N_7610);
nand U8449 (N_8449,N_7181,N_6911);
xor U8450 (N_8450,N_6307,N_7618);
or U8451 (N_8451,N_6237,N_6556);
nand U8452 (N_8452,N_6669,N_6341);
or U8453 (N_8453,N_6549,N_6164);
nor U8454 (N_8454,N_7655,N_7356);
and U8455 (N_8455,N_6964,N_7616);
xnor U8456 (N_8456,N_7196,N_7630);
or U8457 (N_8457,N_7778,N_6044);
nor U8458 (N_8458,N_6207,N_7827);
nand U8459 (N_8459,N_7624,N_6743);
or U8460 (N_8460,N_6512,N_7525);
and U8461 (N_8461,N_7830,N_6467);
nor U8462 (N_8462,N_7389,N_6253);
nand U8463 (N_8463,N_7792,N_6005);
and U8464 (N_8464,N_7203,N_6769);
and U8465 (N_8465,N_7832,N_7556);
or U8466 (N_8466,N_7384,N_7004);
nor U8467 (N_8467,N_7592,N_6995);
nand U8468 (N_8468,N_6192,N_6723);
or U8469 (N_8469,N_6233,N_6890);
nor U8470 (N_8470,N_7082,N_7694);
nor U8471 (N_8471,N_6163,N_7444);
or U8472 (N_8472,N_7123,N_6653);
and U8473 (N_8473,N_6632,N_7477);
or U8474 (N_8474,N_6367,N_7064);
nor U8475 (N_8475,N_6022,N_7757);
xnor U8476 (N_8476,N_6579,N_7911);
or U8477 (N_8477,N_6749,N_7931);
and U8478 (N_8478,N_7945,N_7975);
or U8479 (N_8479,N_6748,N_6458);
nand U8480 (N_8480,N_6353,N_6629);
or U8481 (N_8481,N_7512,N_6070);
nand U8482 (N_8482,N_7677,N_6004);
and U8483 (N_8483,N_6018,N_7318);
nor U8484 (N_8484,N_7954,N_6895);
and U8485 (N_8485,N_7076,N_7591);
nor U8486 (N_8486,N_7350,N_6112);
nor U8487 (N_8487,N_7112,N_7801);
and U8488 (N_8488,N_6371,N_7360);
or U8489 (N_8489,N_7094,N_6840);
nor U8490 (N_8490,N_7989,N_6088);
nand U8491 (N_8491,N_7572,N_7600);
nor U8492 (N_8492,N_6302,N_7320);
nor U8493 (N_8493,N_6588,N_6684);
nor U8494 (N_8494,N_7473,N_7357);
nand U8495 (N_8495,N_7967,N_7416);
nand U8496 (N_8496,N_7551,N_7152);
nor U8497 (N_8497,N_6413,N_6699);
or U8498 (N_8498,N_6738,N_7263);
or U8499 (N_8499,N_6438,N_7811);
nand U8500 (N_8500,N_7128,N_6193);
or U8501 (N_8501,N_7488,N_7960);
nor U8502 (N_8502,N_7354,N_6346);
or U8503 (N_8503,N_6340,N_7500);
nand U8504 (N_8504,N_6967,N_7398);
nor U8505 (N_8505,N_7880,N_6399);
nand U8506 (N_8506,N_6252,N_6386);
and U8507 (N_8507,N_7557,N_7476);
nor U8508 (N_8508,N_6591,N_7019);
nand U8509 (N_8509,N_6016,N_7951);
or U8510 (N_8510,N_7217,N_7731);
nand U8511 (N_8511,N_7718,N_7197);
and U8512 (N_8512,N_7305,N_7017);
nand U8513 (N_8513,N_7034,N_6708);
nand U8514 (N_8514,N_7874,N_6528);
nor U8515 (N_8515,N_6208,N_7962);
and U8516 (N_8516,N_7516,N_7798);
or U8517 (N_8517,N_6146,N_6887);
and U8518 (N_8518,N_7756,N_6686);
or U8519 (N_8519,N_6469,N_6291);
and U8520 (N_8520,N_7087,N_7493);
nand U8521 (N_8521,N_7311,N_7103);
or U8522 (N_8522,N_7521,N_6664);
or U8523 (N_8523,N_6833,N_7582);
or U8524 (N_8524,N_6621,N_7949);
and U8525 (N_8525,N_7847,N_6534);
and U8526 (N_8526,N_6333,N_6366);
nand U8527 (N_8527,N_7777,N_7098);
nor U8528 (N_8528,N_7344,N_6800);
or U8529 (N_8529,N_7386,N_6811);
and U8530 (N_8530,N_6038,N_7788);
nand U8531 (N_8531,N_6225,N_6715);
nor U8532 (N_8532,N_7292,N_7795);
or U8533 (N_8533,N_6065,N_7904);
nand U8534 (N_8534,N_7368,N_7504);
nand U8535 (N_8535,N_7086,N_6919);
or U8536 (N_8536,N_7952,N_6397);
and U8537 (N_8537,N_6186,N_6951);
nand U8538 (N_8538,N_6002,N_7567);
nor U8539 (N_8539,N_7063,N_7501);
nor U8540 (N_8540,N_6596,N_6476);
and U8541 (N_8541,N_7300,N_6194);
and U8542 (N_8542,N_7102,N_7787);
and U8543 (N_8543,N_6646,N_7767);
nor U8544 (N_8544,N_6906,N_6619);
nand U8545 (N_8545,N_7439,N_6127);
or U8546 (N_8546,N_6637,N_6660);
nor U8547 (N_8547,N_6915,N_7657);
and U8548 (N_8548,N_6736,N_7722);
nand U8549 (N_8549,N_6323,N_6204);
xor U8550 (N_8550,N_6726,N_7449);
nand U8551 (N_8551,N_7016,N_6938);
or U8552 (N_8552,N_6183,N_6360);
nor U8553 (N_8553,N_6773,N_6030);
nand U8554 (N_8554,N_6280,N_7643);
nor U8555 (N_8555,N_6418,N_7533);
nor U8556 (N_8556,N_7317,N_6167);
nand U8557 (N_8557,N_7233,N_6365);
nor U8558 (N_8558,N_7621,N_6415);
or U8559 (N_8559,N_6404,N_7328);
or U8560 (N_8560,N_6328,N_6753);
nand U8561 (N_8561,N_7994,N_7213);
nor U8562 (N_8562,N_6983,N_6294);
xnor U8563 (N_8563,N_7201,N_6161);
nor U8564 (N_8564,N_7443,N_6589);
or U8565 (N_8565,N_6551,N_7872);
nor U8566 (N_8566,N_6940,N_7802);
and U8567 (N_8567,N_7668,N_7831);
nor U8568 (N_8568,N_7812,N_7085);
or U8569 (N_8569,N_6673,N_6103);
nand U8570 (N_8570,N_6274,N_7261);
and U8571 (N_8571,N_7511,N_6713);
or U8572 (N_8572,N_6620,N_6370);
or U8573 (N_8573,N_6182,N_6497);
or U8574 (N_8574,N_6812,N_7978);
nor U8575 (N_8575,N_7325,N_7988);
and U8576 (N_8576,N_6412,N_6973);
xor U8577 (N_8577,N_7372,N_6683);
and U8578 (N_8578,N_7980,N_7620);
or U8579 (N_8579,N_6336,N_7837);
or U8580 (N_8580,N_6626,N_6727);
and U8581 (N_8581,N_6988,N_7596);
nor U8582 (N_8582,N_6858,N_6356);
or U8583 (N_8583,N_6676,N_6354);
or U8584 (N_8584,N_6862,N_7143);
and U8585 (N_8585,N_7638,N_7142);
or U8586 (N_8586,N_7562,N_6921);
nor U8587 (N_8587,N_7268,N_6982);
and U8588 (N_8588,N_7965,N_6499);
or U8589 (N_8589,N_7437,N_7375);
nand U8590 (N_8590,N_6496,N_7748);
nand U8591 (N_8591,N_6177,N_6151);
or U8592 (N_8592,N_6121,N_7849);
or U8593 (N_8593,N_6414,N_7822);
nand U8594 (N_8594,N_6910,N_6786);
nand U8595 (N_8595,N_6423,N_7870);
and U8596 (N_8596,N_6658,N_6655);
nor U8597 (N_8597,N_6382,N_7883);
and U8598 (N_8598,N_7038,N_6543);
or U8599 (N_8599,N_6477,N_6250);
nand U8600 (N_8600,N_7299,N_7957);
and U8601 (N_8601,N_7771,N_7370);
or U8602 (N_8602,N_7523,N_6189);
nor U8603 (N_8603,N_6838,N_6692);
nor U8604 (N_8604,N_7061,N_6238);
or U8605 (N_8605,N_7014,N_6012);
or U8606 (N_8606,N_6710,N_6066);
or U8607 (N_8607,N_6142,N_6498);
xor U8608 (N_8608,N_6565,N_6893);
and U8609 (N_8609,N_6502,N_7509);
and U8610 (N_8610,N_6631,N_6679);
and U8611 (N_8611,N_7711,N_6407);
and U8612 (N_8612,N_7855,N_6451);
xnor U8613 (N_8613,N_7028,N_7162);
or U8614 (N_8614,N_6687,N_7987);
xor U8615 (N_8615,N_7109,N_6106);
nor U8616 (N_8616,N_6389,N_6839);
and U8617 (N_8617,N_7717,N_6081);
and U8618 (N_8618,N_7151,N_6891);
or U8619 (N_8619,N_6109,N_7340);
nor U8620 (N_8620,N_7117,N_7608);
or U8621 (N_8621,N_7446,N_6201);
and U8622 (N_8622,N_6078,N_6933);
nor U8623 (N_8623,N_7474,N_6827);
or U8624 (N_8624,N_6444,N_7080);
and U8625 (N_8625,N_6563,N_6554);
or U8626 (N_8626,N_7281,N_6971);
nor U8627 (N_8627,N_6007,N_7069);
xor U8628 (N_8628,N_7277,N_6880);
nand U8629 (N_8629,N_7267,N_7772);
nor U8630 (N_8630,N_7894,N_7541);
and U8631 (N_8631,N_6757,N_7799);
nand U8632 (N_8632,N_6764,N_7382);
and U8633 (N_8633,N_7427,N_7914);
and U8634 (N_8634,N_6107,N_6492);
nor U8635 (N_8635,N_6711,N_6900);
nor U8636 (N_8636,N_7373,N_6123);
nand U8637 (N_8637,N_7744,N_6674);
and U8638 (N_8638,N_7917,N_7698);
and U8639 (N_8639,N_7396,N_7259);
and U8640 (N_8640,N_6440,N_7953);
nor U8641 (N_8641,N_6249,N_6318);
nor U8642 (N_8642,N_7250,N_7680);
or U8643 (N_8643,N_7083,N_6690);
and U8644 (N_8644,N_6488,N_6057);
and U8645 (N_8645,N_7402,N_6375);
and U8646 (N_8646,N_6654,N_6122);
or U8647 (N_8647,N_7342,N_6435);
nand U8648 (N_8648,N_6383,N_6101);
or U8649 (N_8649,N_7423,N_7215);
nor U8650 (N_8650,N_7430,N_6229);
or U8651 (N_8651,N_7740,N_7148);
nor U8652 (N_8652,N_6410,N_6200);
or U8653 (N_8653,N_6871,N_7895);
and U8654 (N_8654,N_7679,N_6999);
nand U8655 (N_8655,N_7081,N_7403);
nand U8656 (N_8656,N_6388,N_6222);
nor U8657 (N_8657,N_7187,N_7464);
or U8658 (N_8658,N_6821,N_6573);
or U8659 (N_8659,N_7555,N_7549);
and U8660 (N_8660,N_6355,N_7899);
nand U8661 (N_8661,N_6506,N_6344);
xnor U8662 (N_8662,N_7805,N_7042);
and U8663 (N_8663,N_6471,N_7959);
nand U8664 (N_8664,N_6529,N_7168);
nor U8665 (N_8665,N_6868,N_6614);
nand U8666 (N_8666,N_6086,N_6758);
nor U8667 (N_8667,N_6533,N_6879);
nor U8668 (N_8668,N_6541,N_7266);
nor U8669 (N_8669,N_6855,N_7358);
nand U8670 (N_8670,N_6181,N_6801);
and U8671 (N_8671,N_7049,N_6530);
and U8672 (N_8672,N_6437,N_6243);
nor U8673 (N_8673,N_7116,N_7361);
nor U8674 (N_8674,N_6602,N_7417);
nand U8675 (N_8675,N_6054,N_7467);
or U8676 (N_8676,N_6947,N_6763);
nand U8677 (N_8677,N_7859,N_6447);
nand U8678 (N_8678,N_6385,N_7542);
or U8679 (N_8679,N_6513,N_6391);
or U8680 (N_8680,N_7295,N_7990);
nor U8681 (N_8681,N_6472,N_6635);
and U8682 (N_8682,N_7619,N_6311);
and U8683 (N_8683,N_7506,N_7020);
or U8684 (N_8684,N_7669,N_6943);
or U8685 (N_8685,N_7759,N_6442);
or U8686 (N_8686,N_7132,N_6053);
or U8687 (N_8687,N_6019,N_6047);
or U8688 (N_8688,N_7119,N_6347);
or U8689 (N_8689,N_7497,N_7724);
and U8690 (N_8690,N_6026,N_7766);
nor U8691 (N_8691,N_7065,N_6849);
or U8692 (N_8692,N_6825,N_7218);
or U8693 (N_8693,N_6834,N_6317);
and U8694 (N_8694,N_6791,N_6041);
or U8695 (N_8695,N_7921,N_7886);
nor U8696 (N_8696,N_6465,N_7466);
nand U8697 (N_8697,N_7359,N_6860);
xnor U8698 (N_8698,N_7762,N_7093);
or U8699 (N_8699,N_6592,N_7369);
nor U8700 (N_8700,N_6097,N_7520);
nor U8701 (N_8701,N_6857,N_6576);
nor U8702 (N_8702,N_6125,N_6931);
or U8703 (N_8703,N_7996,N_6809);
nand U8704 (N_8704,N_7629,N_6647);
and U8705 (N_8705,N_7008,N_7435);
or U8706 (N_8706,N_7502,N_6874);
nand U8707 (N_8707,N_7223,N_6754);
and U8708 (N_8708,N_7130,N_7794);
nor U8709 (N_8709,N_7401,N_7047);
and U8710 (N_8710,N_7274,N_7561);
nand U8711 (N_8711,N_7739,N_6593);
nor U8712 (N_8712,N_6292,N_6577);
and U8713 (N_8713,N_6379,N_6598);
and U8714 (N_8714,N_6996,N_6170);
or U8715 (N_8715,N_7594,N_6482);
nor U8716 (N_8716,N_7961,N_7789);
xnor U8717 (N_8717,N_7648,N_6464);
nor U8718 (N_8718,N_7055,N_7854);
and U8719 (N_8719,N_6990,N_6792);
nor U8720 (N_8720,N_6102,N_6828);
and U8721 (N_8721,N_7941,N_6869);
and U8722 (N_8722,N_6908,N_6050);
and U8723 (N_8723,N_7936,N_6992);
and U8724 (N_8724,N_7705,N_6678);
and U8725 (N_8725,N_7458,N_7923);
or U8726 (N_8726,N_6042,N_7753);
or U8727 (N_8727,N_7537,N_6489);
nor U8728 (N_8728,N_7746,N_7157);
nand U8729 (N_8729,N_7581,N_7682);
nor U8730 (N_8730,N_7339,N_7030);
nand U8731 (N_8731,N_7364,N_6034);
nand U8732 (N_8732,N_6630,N_7136);
nor U8733 (N_8733,N_7438,N_7345);
and U8734 (N_8734,N_6572,N_6538);
nand U8735 (N_8735,N_7365,N_6363);
and U8736 (N_8736,N_6221,N_7878);
and U8737 (N_8737,N_7366,N_7947);
nor U8738 (N_8738,N_6583,N_6359);
nand U8739 (N_8739,N_7336,N_7565);
or U8740 (N_8740,N_6119,N_7036);
nor U8741 (N_8741,N_6242,N_7385);
and U8742 (N_8742,N_7869,N_6901);
or U8743 (N_8743,N_6178,N_6507);
and U8744 (N_8744,N_7067,N_6627);
or U8745 (N_8745,N_6954,N_6745);
or U8746 (N_8746,N_7651,N_6848);
nand U8747 (N_8747,N_7393,N_6325);
or U8748 (N_8748,N_6772,N_7278);
nand U8749 (N_8749,N_6641,N_7518);
or U8750 (N_8750,N_6303,N_7627);
or U8751 (N_8751,N_7642,N_7607);
and U8752 (N_8752,N_7256,N_7413);
or U8753 (N_8753,N_7710,N_6640);
or U8754 (N_8754,N_7486,N_6907);
nand U8755 (N_8755,N_7003,N_7713);
nand U8756 (N_8756,N_7877,N_7195);
nor U8757 (N_8757,N_6609,N_7252);
nand U8758 (N_8758,N_7229,N_7039);
nor U8759 (N_8759,N_7472,N_6212);
nand U8760 (N_8760,N_7054,N_7626);
nor U8761 (N_8761,N_6211,N_6244);
nand U8762 (N_8762,N_7184,N_6557);
nor U8763 (N_8763,N_7141,N_7432);
or U8764 (N_8764,N_7302,N_6408);
nor U8765 (N_8765,N_7436,N_7584);
or U8766 (N_8766,N_7966,N_7839);
and U8767 (N_8767,N_7678,N_7760);
nor U8768 (N_8768,N_6116,N_7457);
nand U8769 (N_8769,N_6740,N_6468);
nand U8770 (N_8770,N_7469,N_6462);
nor U8771 (N_8771,N_7275,N_7226);
nand U8772 (N_8772,N_7901,N_7387);
nor U8773 (N_8773,N_6994,N_6642);
nand U8774 (N_8774,N_6374,N_6401);
or U8775 (N_8775,N_6220,N_7108);
nand U8776 (N_8776,N_6725,N_6064);
or U8777 (N_8777,N_7662,N_7101);
and U8778 (N_8778,N_7800,N_7408);
and U8779 (N_8779,N_6661,N_7950);
and U8780 (N_8780,N_6770,N_7514);
and U8781 (N_8781,N_7920,N_7709);
and U8782 (N_8782,N_6315,N_6707);
nand U8783 (N_8783,N_6144,N_6633);
or U8784 (N_8784,N_6460,N_6799);
or U8785 (N_8785,N_6118,N_6068);
nand U8786 (N_8786,N_6805,N_6819);
nand U8787 (N_8787,N_7775,N_7276);
nand U8788 (N_8788,N_6120,N_6245);
nand U8789 (N_8789,N_7051,N_7031);
nor U8790 (N_8790,N_6569,N_7091);
nor U8791 (N_8791,N_7188,N_6024);
nand U8792 (N_8792,N_6457,N_7485);
and U8793 (N_8793,N_6886,N_6845);
xnor U8794 (N_8794,N_6599,N_7456);
nand U8795 (N_8795,N_6815,N_6236);
nand U8796 (N_8796,N_7287,N_7796);
nand U8797 (N_8797,N_6175,N_7210);
or U8798 (N_8798,N_6046,N_6148);
nand U8799 (N_8799,N_6433,N_7337);
or U8800 (N_8800,N_6173,N_7175);
nor U8801 (N_8801,N_7316,N_6888);
nand U8802 (N_8802,N_7150,N_6091);
and U8803 (N_8803,N_6525,N_7573);
nor U8804 (N_8804,N_6376,N_6875);
and U8805 (N_8805,N_7470,N_7823);
and U8806 (N_8806,N_6209,N_7046);
or U8807 (N_8807,N_6567,N_6380);
or U8808 (N_8808,N_6671,N_6582);
and U8809 (N_8809,N_7240,N_6322);
and U8810 (N_8810,N_6349,N_7471);
nor U8811 (N_8811,N_6991,N_6681);
nand U8812 (N_8812,N_7887,N_7897);
nand U8813 (N_8813,N_7652,N_7958);
and U8814 (N_8814,N_6113,N_6691);
nand U8815 (N_8815,N_6968,N_7708);
nor U8816 (N_8816,N_7675,N_7251);
nand U8817 (N_8817,N_7131,N_7285);
nor U8818 (N_8818,N_7499,N_6559);
and U8819 (N_8819,N_6950,N_7189);
and U8820 (N_8820,N_6021,N_6409);
nand U8821 (N_8821,N_6788,N_7147);
nand U8822 (N_8822,N_7773,N_7689);
and U8823 (N_8823,N_6594,N_6980);
or U8824 (N_8824,N_7658,N_7241);
or U8825 (N_8825,N_7072,N_7846);
nor U8826 (N_8826,N_6339,N_7010);
nor U8827 (N_8827,N_7636,N_6787);
nand U8828 (N_8828,N_6160,N_7242);
nor U8829 (N_8829,N_6555,N_7478);
nand U8830 (N_8830,N_6814,N_6480);
nand U8831 (N_8831,N_7692,N_6114);
nor U8832 (N_8832,N_7244,N_6059);
or U8833 (N_8833,N_6003,N_7089);
nand U8834 (N_8834,N_6985,N_6929);
or U8835 (N_8835,N_6092,N_6277);
or U8836 (N_8836,N_7161,N_6320);
or U8837 (N_8837,N_7664,N_7454);
and U8838 (N_8838,N_7519,N_6545);
nor U8839 (N_8839,N_6517,N_7262);
or U8840 (N_8840,N_7406,N_7840);
or U8841 (N_8841,N_7104,N_7687);
nor U8842 (N_8842,N_6714,N_7817);
and U8843 (N_8843,N_6230,N_7929);
nor U8844 (N_8844,N_6600,N_7670);
and U8845 (N_8845,N_7544,N_7598);
nand U8846 (N_8846,N_6547,N_7948);
or U8847 (N_8847,N_7876,N_7451);
nand U8848 (N_8848,N_6241,N_7588);
and U8849 (N_8849,N_6866,N_6439);
or U8850 (N_8850,N_6486,N_7858);
nand U8851 (N_8851,N_6319,N_7538);
nand U8852 (N_8852,N_7761,N_7431);
or U8853 (N_8853,N_6830,N_6851);
nand U8854 (N_8854,N_7535,N_6544);
or U8855 (N_8855,N_6638,N_6449);
nand U8856 (N_8856,N_7489,N_7321);
and U8857 (N_8857,N_6847,N_7927);
xor U8858 (N_8858,N_6232,N_7397);
or U8859 (N_8859,N_7341,N_7002);
nand U8860 (N_8860,N_6384,N_7400);
and U8861 (N_8861,N_6296,N_7179);
or U8862 (N_8862,N_7681,N_7418);
and U8863 (N_8863,N_6036,N_6083);
or U8864 (N_8864,N_6487,N_6373);
nand U8865 (N_8865,N_7543,N_6282);
nor U8866 (N_8866,N_6278,N_7480);
or U8867 (N_8867,N_7848,N_6217);
nand U8868 (N_8868,N_7964,N_7625);
nand U8869 (N_8869,N_7530,N_7723);
nor U8870 (N_8870,N_7553,N_6884);
and U8871 (N_8871,N_7405,N_7804);
nor U8872 (N_8872,N_7720,N_7641);
and U8873 (N_8873,N_6202,N_7688);
or U8874 (N_8874,N_6709,N_6514);
and U8875 (N_8875,N_6421,N_6000);
or U8876 (N_8876,N_6390,N_7293);
and U8877 (N_8877,N_6313,N_6975);
nand U8878 (N_8878,N_6766,N_6290);
nor U8879 (N_8879,N_6813,N_7866);
nor U8880 (N_8880,N_7999,N_6459);
and U8881 (N_8881,N_7421,N_6111);
nand U8882 (N_8882,N_7284,N_7322);
nor U8883 (N_8883,N_7686,N_7785);
nor U8884 (N_8884,N_6894,N_7154);
xnor U8885 (N_8885,N_6578,N_7414);
nand U8886 (N_8886,N_6666,N_7399);
nand U8887 (N_8887,N_6731,N_7219);
nand U8888 (N_8888,N_7985,N_7404);
or U8889 (N_8889,N_7006,N_7045);
nand U8890 (N_8890,N_6045,N_6300);
nor U8891 (N_8891,N_6343,N_7529);
nand U8892 (N_8892,N_7127,N_7044);
or U8893 (N_8893,N_6394,N_7468);
nand U8894 (N_8894,N_6644,N_6796);
nand U8895 (N_8895,N_6516,N_6432);
and U8896 (N_8896,N_7560,N_6490);
nand U8897 (N_8897,N_7463,N_6061);
nand U8898 (N_8898,N_6927,N_6570);
nor U8899 (N_8899,N_6883,N_6668);
nand U8900 (N_8900,N_7946,N_7298);
and U8901 (N_8901,N_7982,N_7736);
or U8902 (N_8902,N_6248,N_7683);
and U8903 (N_8903,N_6755,N_7991);
nor U8904 (N_8904,N_7492,N_7260);
nor U8905 (N_8905,N_7715,N_7124);
or U8906 (N_8906,N_7060,N_7702);
nor U8907 (N_8907,N_6505,N_7144);
nor U8908 (N_8908,N_7735,N_6357);
or U8909 (N_8909,N_7908,N_6730);
and U8910 (N_8910,N_6877,N_7335);
and U8911 (N_8911,N_7153,N_6271);
and U8912 (N_8912,N_7190,N_7319);
or U8913 (N_8913,N_6205,N_6542);
nand U8914 (N_8914,N_7986,N_6257);
nand U8915 (N_8915,N_7040,N_7900);
xnor U8916 (N_8916,N_6898,N_6276);
nor U8917 (N_8917,N_6716,N_6719);
and U8918 (N_8918,N_7741,N_7940);
nor U8919 (N_8919,N_6084,N_6093);
nand U8920 (N_8920,N_6043,N_6031);
or U8921 (N_8921,N_7586,N_7191);
and U8922 (N_8922,N_6656,N_7246);
and U8923 (N_8923,N_6680,N_6015);
or U8924 (N_8924,N_6327,N_7755);
nand U8925 (N_8925,N_7743,N_6403);
and U8926 (N_8926,N_6826,N_6312);
nand U8927 (N_8927,N_6270,N_7622);
or U8928 (N_8928,N_7095,N_6560);
nor U8929 (N_8929,N_6247,N_7879);
nor U8930 (N_8930,N_7442,N_7609);
and U8931 (N_8931,N_7035,N_7704);
or U8932 (N_8932,N_6332,N_6461);
or U8933 (N_8933,N_6945,N_7388);
and U8934 (N_8934,N_6777,N_6956);
nand U8935 (N_8935,N_6521,N_6174);
nor U8936 (N_8936,N_7611,N_7475);
nand U8937 (N_8937,N_6611,N_6345);
or U8938 (N_8938,N_6832,N_6396);
nand U8939 (N_8939,N_6239,N_7890);
or U8940 (N_8940,N_6348,N_7156);
and U8941 (N_8941,N_6859,N_6213);
or U8942 (N_8942,N_6751,N_7838);
nand U8943 (N_8943,N_6957,N_7825);
or U8944 (N_8944,N_6284,N_7903);
and U8945 (N_8945,N_6704,N_6199);
and U8946 (N_8946,N_6922,N_6293);
nor U8947 (N_8947,N_6272,N_7023);
nor U8948 (N_8948,N_6761,N_7821);
and U8949 (N_8949,N_7009,N_6299);
nand U8950 (N_8950,N_6804,N_7758);
nand U8951 (N_8951,N_7971,N_6998);
nand U8952 (N_8952,N_6688,N_6934);
or U8953 (N_8953,N_7515,N_6132);
or U8954 (N_8954,N_6075,N_7185);
and U8955 (N_8955,N_7528,N_6978);
nor U8956 (N_8956,N_7550,N_6889);
nor U8957 (N_8957,N_6737,N_6425);
nor U8958 (N_8958,N_7938,N_6511);
nand U8959 (N_8959,N_6073,N_6746);
or U8960 (N_8960,N_6264,N_7205);
or U8961 (N_8961,N_7481,N_6470);
nor U8962 (N_8962,N_7440,N_7749);
nor U8963 (N_8963,N_7737,N_7860);
nor U8964 (N_8964,N_6590,N_7998);
nand U8965 (N_8965,N_7637,N_6914);
nand U8966 (N_8966,N_7969,N_6803);
nand U8967 (N_8967,N_6434,N_6153);
nand U8968 (N_8968,N_7604,N_7942);
or U8969 (N_8969,N_7820,N_7078);
and U8970 (N_8970,N_6762,N_7100);
nand U8971 (N_8971,N_6566,N_6729);
nand U8972 (N_8972,N_6926,N_7882);
and U8973 (N_8973,N_7265,N_6625);
nor U8974 (N_8974,N_6558,N_6493);
nand U8975 (N_8975,N_7684,N_6261);
nor U8976 (N_8976,N_6268,N_6853);
nor U8977 (N_8977,N_7548,N_6698);
nor U8978 (N_8978,N_6419,N_7186);
and U8979 (N_8979,N_6774,N_7309);
nand U8980 (N_8980,N_7307,N_7465);
nor U8981 (N_8981,N_6334,N_7425);
or U8982 (N_8982,N_7236,N_6129);
nor U8983 (N_8983,N_7163,N_7864);
nand U8984 (N_8984,N_7742,N_6802);
and U8985 (N_8985,N_7052,N_7137);
or U8986 (N_8986,N_7429,N_7647);
nor U8987 (N_8987,N_7459,N_7097);
or U8988 (N_8988,N_7228,N_7995);
or U8989 (N_8989,N_7315,N_6939);
nand U8990 (N_8990,N_7333,N_6997);
nor U8991 (N_8991,N_7721,N_7348);
nor U8992 (N_8992,N_7411,N_7976);
or U8993 (N_8993,N_7379,N_6436);
nor U8994 (N_8994,N_7833,N_7574);
or U8995 (N_8995,N_6010,N_7001);
nand U8996 (N_8996,N_7253,N_6062);
nor U8997 (N_8997,N_7479,N_6454);
xor U8998 (N_8998,N_6864,N_7428);
or U8999 (N_8999,N_6358,N_6979);
nor U9000 (N_9000,N_6596,N_6214);
nand U9001 (N_9001,N_7796,N_7079);
nor U9002 (N_9002,N_7396,N_6547);
and U9003 (N_9003,N_7795,N_7787);
and U9004 (N_9004,N_7802,N_6497);
and U9005 (N_9005,N_6023,N_6446);
and U9006 (N_9006,N_7865,N_6283);
nor U9007 (N_9007,N_7628,N_6820);
nand U9008 (N_9008,N_6692,N_6693);
nand U9009 (N_9009,N_7625,N_6797);
and U9010 (N_9010,N_7228,N_7796);
nand U9011 (N_9011,N_7765,N_7616);
nor U9012 (N_9012,N_7155,N_7420);
or U9013 (N_9013,N_6980,N_7991);
nor U9014 (N_9014,N_7505,N_6106);
nand U9015 (N_9015,N_7473,N_6518);
and U9016 (N_9016,N_6862,N_7736);
and U9017 (N_9017,N_7878,N_6413);
or U9018 (N_9018,N_7099,N_7767);
nand U9019 (N_9019,N_7496,N_6401);
and U9020 (N_9020,N_7253,N_6432);
nor U9021 (N_9021,N_6217,N_6753);
or U9022 (N_9022,N_6634,N_6415);
nor U9023 (N_9023,N_7613,N_7377);
nand U9024 (N_9024,N_7735,N_7579);
nor U9025 (N_9025,N_7060,N_7735);
or U9026 (N_9026,N_7881,N_6186);
nor U9027 (N_9027,N_7162,N_6039);
or U9028 (N_9028,N_6724,N_6081);
nor U9029 (N_9029,N_6033,N_7515);
nor U9030 (N_9030,N_7772,N_6614);
or U9031 (N_9031,N_6247,N_7455);
and U9032 (N_9032,N_7070,N_6514);
nor U9033 (N_9033,N_6780,N_6968);
xnor U9034 (N_9034,N_6639,N_6169);
nand U9035 (N_9035,N_6680,N_6787);
nor U9036 (N_9036,N_7462,N_6070);
or U9037 (N_9037,N_7145,N_7702);
xor U9038 (N_9038,N_6600,N_7233);
and U9039 (N_9039,N_6243,N_6838);
nor U9040 (N_9040,N_7658,N_7636);
nor U9041 (N_9041,N_7295,N_6836);
nor U9042 (N_9042,N_6286,N_7024);
or U9043 (N_9043,N_6161,N_6961);
nand U9044 (N_9044,N_7659,N_6748);
nor U9045 (N_9045,N_7361,N_7962);
or U9046 (N_9046,N_7504,N_6138);
nand U9047 (N_9047,N_7479,N_6472);
or U9048 (N_9048,N_6841,N_7806);
and U9049 (N_9049,N_6168,N_7545);
nor U9050 (N_9050,N_6174,N_7410);
or U9051 (N_9051,N_6921,N_6798);
and U9052 (N_9052,N_7029,N_6611);
and U9053 (N_9053,N_6400,N_7309);
and U9054 (N_9054,N_7485,N_7197);
and U9055 (N_9055,N_6594,N_7548);
nor U9056 (N_9056,N_7651,N_6418);
nor U9057 (N_9057,N_6339,N_6755);
nor U9058 (N_9058,N_7064,N_6373);
nand U9059 (N_9059,N_6369,N_7196);
and U9060 (N_9060,N_7692,N_7795);
nand U9061 (N_9061,N_6748,N_6380);
and U9062 (N_9062,N_7126,N_7321);
or U9063 (N_9063,N_7121,N_6996);
and U9064 (N_9064,N_6385,N_6320);
and U9065 (N_9065,N_6846,N_6137);
or U9066 (N_9066,N_6263,N_6443);
and U9067 (N_9067,N_7743,N_6389);
nand U9068 (N_9068,N_7307,N_7667);
and U9069 (N_9069,N_6272,N_7681);
or U9070 (N_9070,N_6417,N_7179);
or U9071 (N_9071,N_7051,N_7482);
and U9072 (N_9072,N_7686,N_6143);
nand U9073 (N_9073,N_7520,N_6246);
and U9074 (N_9074,N_6689,N_7775);
or U9075 (N_9075,N_6013,N_6475);
or U9076 (N_9076,N_6115,N_6450);
or U9077 (N_9077,N_6232,N_6676);
nor U9078 (N_9078,N_6650,N_7999);
nor U9079 (N_9079,N_7585,N_7922);
and U9080 (N_9080,N_6910,N_7828);
or U9081 (N_9081,N_6763,N_6800);
and U9082 (N_9082,N_6080,N_6962);
and U9083 (N_9083,N_6470,N_7426);
nand U9084 (N_9084,N_6630,N_7000);
or U9085 (N_9085,N_6224,N_6837);
nor U9086 (N_9086,N_6240,N_7968);
and U9087 (N_9087,N_7941,N_7402);
nor U9088 (N_9088,N_7565,N_6420);
nor U9089 (N_9089,N_6744,N_6428);
or U9090 (N_9090,N_6234,N_6456);
or U9091 (N_9091,N_7036,N_7117);
nor U9092 (N_9092,N_6367,N_6103);
nand U9093 (N_9093,N_7025,N_7513);
nor U9094 (N_9094,N_6572,N_6635);
and U9095 (N_9095,N_6466,N_7038);
and U9096 (N_9096,N_6494,N_7347);
and U9097 (N_9097,N_6562,N_7800);
and U9098 (N_9098,N_7248,N_6672);
or U9099 (N_9099,N_6719,N_6440);
and U9100 (N_9100,N_7059,N_7389);
nor U9101 (N_9101,N_6096,N_7278);
or U9102 (N_9102,N_7573,N_6067);
and U9103 (N_9103,N_7530,N_6908);
nor U9104 (N_9104,N_6305,N_6180);
and U9105 (N_9105,N_7326,N_6909);
or U9106 (N_9106,N_6464,N_6720);
or U9107 (N_9107,N_6687,N_7011);
nand U9108 (N_9108,N_7789,N_7486);
nand U9109 (N_9109,N_7026,N_6710);
nor U9110 (N_9110,N_6641,N_6450);
nor U9111 (N_9111,N_6194,N_7685);
nand U9112 (N_9112,N_7425,N_7787);
and U9113 (N_9113,N_7518,N_7693);
or U9114 (N_9114,N_7079,N_6338);
nand U9115 (N_9115,N_6917,N_7028);
nor U9116 (N_9116,N_6020,N_7277);
and U9117 (N_9117,N_7022,N_7803);
nand U9118 (N_9118,N_6981,N_6439);
and U9119 (N_9119,N_7922,N_7550);
nor U9120 (N_9120,N_6289,N_6302);
nor U9121 (N_9121,N_6910,N_6179);
nor U9122 (N_9122,N_7183,N_7201);
and U9123 (N_9123,N_6859,N_6383);
and U9124 (N_9124,N_6648,N_7032);
nor U9125 (N_9125,N_7764,N_7691);
nor U9126 (N_9126,N_7239,N_6548);
and U9127 (N_9127,N_7733,N_7689);
nor U9128 (N_9128,N_6119,N_7762);
nor U9129 (N_9129,N_6907,N_7390);
nand U9130 (N_9130,N_6710,N_6758);
nand U9131 (N_9131,N_7134,N_7986);
nand U9132 (N_9132,N_6913,N_7746);
nand U9133 (N_9133,N_6957,N_6642);
nand U9134 (N_9134,N_6923,N_6878);
nand U9135 (N_9135,N_6497,N_6610);
and U9136 (N_9136,N_6788,N_6534);
nand U9137 (N_9137,N_7973,N_7154);
or U9138 (N_9138,N_6688,N_7845);
nor U9139 (N_9139,N_6954,N_7828);
or U9140 (N_9140,N_7176,N_7834);
and U9141 (N_9141,N_7650,N_7132);
nand U9142 (N_9142,N_7559,N_6293);
nand U9143 (N_9143,N_6649,N_6499);
nor U9144 (N_9144,N_7572,N_7471);
or U9145 (N_9145,N_7866,N_7601);
and U9146 (N_9146,N_6849,N_6307);
or U9147 (N_9147,N_7414,N_7396);
nand U9148 (N_9148,N_6447,N_6962);
and U9149 (N_9149,N_6487,N_7707);
nand U9150 (N_9150,N_6157,N_7151);
nand U9151 (N_9151,N_7952,N_7521);
and U9152 (N_9152,N_6947,N_6630);
nand U9153 (N_9153,N_7271,N_7938);
or U9154 (N_9154,N_6154,N_7688);
nor U9155 (N_9155,N_7274,N_7091);
nor U9156 (N_9156,N_6451,N_6426);
nor U9157 (N_9157,N_6742,N_6290);
nor U9158 (N_9158,N_7396,N_7606);
and U9159 (N_9159,N_7234,N_7570);
or U9160 (N_9160,N_7042,N_6044);
or U9161 (N_9161,N_6294,N_7223);
nand U9162 (N_9162,N_6780,N_6849);
and U9163 (N_9163,N_6895,N_7020);
or U9164 (N_9164,N_6132,N_7234);
or U9165 (N_9165,N_7821,N_6470);
or U9166 (N_9166,N_6790,N_6593);
nor U9167 (N_9167,N_7196,N_6374);
or U9168 (N_9168,N_7339,N_6230);
nor U9169 (N_9169,N_6622,N_6642);
or U9170 (N_9170,N_6484,N_6518);
and U9171 (N_9171,N_7049,N_6304);
xor U9172 (N_9172,N_6930,N_7753);
nor U9173 (N_9173,N_7115,N_6973);
or U9174 (N_9174,N_7217,N_6721);
nor U9175 (N_9175,N_6786,N_6355);
xnor U9176 (N_9176,N_7051,N_6770);
nor U9177 (N_9177,N_7950,N_7058);
nor U9178 (N_9178,N_6621,N_6804);
nor U9179 (N_9179,N_6330,N_7654);
and U9180 (N_9180,N_7447,N_6309);
nor U9181 (N_9181,N_6534,N_7282);
or U9182 (N_9182,N_7417,N_6256);
nor U9183 (N_9183,N_7161,N_6831);
nand U9184 (N_9184,N_6445,N_6954);
and U9185 (N_9185,N_7675,N_7556);
and U9186 (N_9186,N_6940,N_6872);
or U9187 (N_9187,N_6405,N_7778);
nor U9188 (N_9188,N_6470,N_6018);
or U9189 (N_9189,N_6392,N_7022);
and U9190 (N_9190,N_7591,N_7451);
nor U9191 (N_9191,N_7741,N_6098);
nor U9192 (N_9192,N_7844,N_6116);
and U9193 (N_9193,N_6432,N_6500);
nand U9194 (N_9194,N_7884,N_7529);
or U9195 (N_9195,N_6360,N_7517);
and U9196 (N_9196,N_7693,N_7412);
or U9197 (N_9197,N_6424,N_7488);
or U9198 (N_9198,N_6426,N_7508);
or U9199 (N_9199,N_6242,N_6938);
and U9200 (N_9200,N_7002,N_6419);
nand U9201 (N_9201,N_6270,N_6473);
nand U9202 (N_9202,N_6925,N_6864);
nand U9203 (N_9203,N_7955,N_6903);
nand U9204 (N_9204,N_7090,N_6976);
or U9205 (N_9205,N_7026,N_7237);
or U9206 (N_9206,N_6168,N_7355);
nand U9207 (N_9207,N_7381,N_6763);
and U9208 (N_9208,N_7706,N_6419);
and U9209 (N_9209,N_6488,N_7569);
and U9210 (N_9210,N_6972,N_7727);
nand U9211 (N_9211,N_7404,N_6234);
or U9212 (N_9212,N_6700,N_6228);
nand U9213 (N_9213,N_7950,N_7236);
nor U9214 (N_9214,N_7644,N_6774);
or U9215 (N_9215,N_6162,N_6277);
and U9216 (N_9216,N_6725,N_7814);
and U9217 (N_9217,N_6902,N_6045);
and U9218 (N_9218,N_6327,N_6919);
and U9219 (N_9219,N_7987,N_7379);
or U9220 (N_9220,N_7630,N_6040);
and U9221 (N_9221,N_6158,N_6436);
nor U9222 (N_9222,N_6896,N_7109);
and U9223 (N_9223,N_6530,N_7058);
nand U9224 (N_9224,N_6716,N_7038);
nand U9225 (N_9225,N_6946,N_7762);
nor U9226 (N_9226,N_6444,N_7467);
nand U9227 (N_9227,N_7064,N_6311);
and U9228 (N_9228,N_7574,N_6040);
or U9229 (N_9229,N_6961,N_7747);
nand U9230 (N_9230,N_7220,N_7476);
and U9231 (N_9231,N_7768,N_7913);
nand U9232 (N_9232,N_6118,N_6885);
and U9233 (N_9233,N_6729,N_7800);
and U9234 (N_9234,N_7132,N_6798);
nand U9235 (N_9235,N_7405,N_6930);
nand U9236 (N_9236,N_7790,N_7077);
and U9237 (N_9237,N_6069,N_7868);
nor U9238 (N_9238,N_6224,N_7888);
nand U9239 (N_9239,N_6005,N_6672);
or U9240 (N_9240,N_7279,N_6238);
or U9241 (N_9241,N_7917,N_7031);
nand U9242 (N_9242,N_6022,N_6039);
or U9243 (N_9243,N_7443,N_7037);
or U9244 (N_9244,N_6224,N_7516);
nand U9245 (N_9245,N_6127,N_7564);
or U9246 (N_9246,N_7338,N_6260);
or U9247 (N_9247,N_7521,N_7714);
xor U9248 (N_9248,N_7684,N_7767);
or U9249 (N_9249,N_7655,N_7180);
nor U9250 (N_9250,N_6249,N_6567);
or U9251 (N_9251,N_6656,N_6657);
or U9252 (N_9252,N_6591,N_6864);
or U9253 (N_9253,N_6445,N_6505);
nand U9254 (N_9254,N_7096,N_6038);
nor U9255 (N_9255,N_6669,N_7841);
nor U9256 (N_9256,N_7264,N_6463);
or U9257 (N_9257,N_6223,N_7647);
or U9258 (N_9258,N_6181,N_6039);
and U9259 (N_9259,N_6511,N_6151);
nand U9260 (N_9260,N_6131,N_7327);
or U9261 (N_9261,N_6758,N_6202);
and U9262 (N_9262,N_6675,N_7266);
and U9263 (N_9263,N_7409,N_6657);
and U9264 (N_9264,N_6136,N_6406);
or U9265 (N_9265,N_6707,N_6847);
nor U9266 (N_9266,N_6958,N_6535);
nor U9267 (N_9267,N_6065,N_6997);
nor U9268 (N_9268,N_6644,N_7279);
nor U9269 (N_9269,N_6145,N_7642);
nor U9270 (N_9270,N_6866,N_6593);
nand U9271 (N_9271,N_6337,N_6701);
nand U9272 (N_9272,N_7369,N_7855);
nand U9273 (N_9273,N_7866,N_6749);
and U9274 (N_9274,N_6594,N_7559);
nor U9275 (N_9275,N_7405,N_6126);
or U9276 (N_9276,N_7398,N_6872);
nor U9277 (N_9277,N_7878,N_6353);
and U9278 (N_9278,N_6924,N_7319);
or U9279 (N_9279,N_6022,N_7080);
and U9280 (N_9280,N_6178,N_6453);
nand U9281 (N_9281,N_6429,N_6896);
or U9282 (N_9282,N_7843,N_6121);
nor U9283 (N_9283,N_7304,N_7699);
nand U9284 (N_9284,N_6979,N_6476);
nand U9285 (N_9285,N_6283,N_6399);
nor U9286 (N_9286,N_6072,N_6148);
or U9287 (N_9287,N_7274,N_6698);
or U9288 (N_9288,N_7449,N_6761);
or U9289 (N_9289,N_6901,N_6031);
nand U9290 (N_9290,N_6730,N_6148);
nor U9291 (N_9291,N_7842,N_7315);
or U9292 (N_9292,N_6608,N_7584);
and U9293 (N_9293,N_7060,N_6435);
or U9294 (N_9294,N_7107,N_7757);
or U9295 (N_9295,N_7384,N_7292);
or U9296 (N_9296,N_7203,N_6173);
nand U9297 (N_9297,N_7695,N_7476);
or U9298 (N_9298,N_7348,N_7600);
nand U9299 (N_9299,N_6406,N_7050);
or U9300 (N_9300,N_7869,N_6384);
and U9301 (N_9301,N_7386,N_7698);
and U9302 (N_9302,N_6658,N_6321);
nor U9303 (N_9303,N_7911,N_6979);
or U9304 (N_9304,N_7055,N_7185);
nand U9305 (N_9305,N_7551,N_6717);
nand U9306 (N_9306,N_7486,N_6481);
nor U9307 (N_9307,N_6808,N_7081);
and U9308 (N_9308,N_7727,N_7873);
or U9309 (N_9309,N_7748,N_7941);
or U9310 (N_9310,N_6758,N_6729);
or U9311 (N_9311,N_7229,N_7063);
nand U9312 (N_9312,N_7310,N_6062);
and U9313 (N_9313,N_7156,N_7746);
nor U9314 (N_9314,N_7122,N_7550);
nand U9315 (N_9315,N_6228,N_6483);
nand U9316 (N_9316,N_6235,N_7693);
and U9317 (N_9317,N_7271,N_6163);
and U9318 (N_9318,N_7251,N_7154);
and U9319 (N_9319,N_7405,N_7943);
nand U9320 (N_9320,N_7298,N_7380);
nand U9321 (N_9321,N_6326,N_6004);
or U9322 (N_9322,N_6464,N_7029);
or U9323 (N_9323,N_6613,N_7309);
nand U9324 (N_9324,N_6737,N_7169);
nand U9325 (N_9325,N_7147,N_6043);
nand U9326 (N_9326,N_6172,N_6637);
and U9327 (N_9327,N_6446,N_7307);
or U9328 (N_9328,N_6106,N_6366);
and U9329 (N_9329,N_6649,N_7476);
nand U9330 (N_9330,N_6357,N_6922);
or U9331 (N_9331,N_7593,N_7278);
nand U9332 (N_9332,N_7829,N_6943);
nor U9333 (N_9333,N_6025,N_7825);
nor U9334 (N_9334,N_6669,N_7282);
xnor U9335 (N_9335,N_6330,N_6883);
nor U9336 (N_9336,N_6398,N_7561);
nand U9337 (N_9337,N_7502,N_7725);
nand U9338 (N_9338,N_7711,N_6472);
and U9339 (N_9339,N_7910,N_6388);
nor U9340 (N_9340,N_6595,N_7897);
nand U9341 (N_9341,N_7242,N_7089);
or U9342 (N_9342,N_7911,N_7947);
nand U9343 (N_9343,N_6160,N_6991);
nor U9344 (N_9344,N_6599,N_7976);
or U9345 (N_9345,N_7420,N_7491);
nor U9346 (N_9346,N_6442,N_7127);
nor U9347 (N_9347,N_7772,N_7583);
nand U9348 (N_9348,N_6371,N_6631);
nor U9349 (N_9349,N_6451,N_7911);
or U9350 (N_9350,N_6295,N_6396);
and U9351 (N_9351,N_6730,N_7980);
or U9352 (N_9352,N_7528,N_7300);
nand U9353 (N_9353,N_7739,N_6398);
nand U9354 (N_9354,N_7566,N_7199);
xor U9355 (N_9355,N_7394,N_7090);
or U9356 (N_9356,N_6043,N_7578);
and U9357 (N_9357,N_7595,N_7427);
nand U9358 (N_9358,N_7803,N_7366);
and U9359 (N_9359,N_7125,N_6692);
and U9360 (N_9360,N_7681,N_6250);
or U9361 (N_9361,N_6899,N_6601);
nand U9362 (N_9362,N_7063,N_7489);
or U9363 (N_9363,N_7314,N_6520);
nor U9364 (N_9364,N_6668,N_6230);
nor U9365 (N_9365,N_7647,N_6092);
and U9366 (N_9366,N_7408,N_7250);
xnor U9367 (N_9367,N_7867,N_7749);
or U9368 (N_9368,N_7892,N_6402);
and U9369 (N_9369,N_7759,N_6189);
nand U9370 (N_9370,N_7966,N_6349);
and U9371 (N_9371,N_7768,N_7473);
and U9372 (N_9372,N_7299,N_7098);
xor U9373 (N_9373,N_7103,N_7616);
nand U9374 (N_9374,N_7795,N_7760);
nand U9375 (N_9375,N_7981,N_7246);
nand U9376 (N_9376,N_7228,N_7255);
and U9377 (N_9377,N_6506,N_7273);
nand U9378 (N_9378,N_7021,N_6392);
nand U9379 (N_9379,N_6820,N_6999);
or U9380 (N_9380,N_6840,N_6275);
nor U9381 (N_9381,N_6803,N_7158);
or U9382 (N_9382,N_6799,N_6715);
or U9383 (N_9383,N_7352,N_6477);
nand U9384 (N_9384,N_6364,N_6138);
or U9385 (N_9385,N_6021,N_7137);
nor U9386 (N_9386,N_6667,N_6792);
xor U9387 (N_9387,N_7903,N_7468);
nand U9388 (N_9388,N_7238,N_6880);
and U9389 (N_9389,N_6266,N_6220);
and U9390 (N_9390,N_6127,N_7449);
nor U9391 (N_9391,N_7763,N_7699);
or U9392 (N_9392,N_6311,N_6928);
nor U9393 (N_9393,N_7701,N_7963);
and U9394 (N_9394,N_7192,N_7380);
and U9395 (N_9395,N_6623,N_6705);
nor U9396 (N_9396,N_6794,N_6565);
nand U9397 (N_9397,N_6496,N_7175);
nor U9398 (N_9398,N_6192,N_6627);
or U9399 (N_9399,N_6819,N_6843);
nand U9400 (N_9400,N_7302,N_7129);
or U9401 (N_9401,N_7376,N_7148);
or U9402 (N_9402,N_6733,N_6081);
or U9403 (N_9403,N_7029,N_6046);
xor U9404 (N_9404,N_7403,N_6060);
nand U9405 (N_9405,N_6792,N_7910);
nand U9406 (N_9406,N_7078,N_7698);
and U9407 (N_9407,N_7384,N_7492);
and U9408 (N_9408,N_6802,N_6040);
or U9409 (N_9409,N_7710,N_6817);
and U9410 (N_9410,N_7138,N_6244);
nand U9411 (N_9411,N_6358,N_6246);
xor U9412 (N_9412,N_7340,N_7866);
and U9413 (N_9413,N_6349,N_7378);
or U9414 (N_9414,N_6884,N_7805);
nand U9415 (N_9415,N_6541,N_7129);
nor U9416 (N_9416,N_6175,N_7821);
nand U9417 (N_9417,N_6958,N_6384);
and U9418 (N_9418,N_6903,N_6495);
nand U9419 (N_9419,N_6087,N_7899);
or U9420 (N_9420,N_7556,N_6603);
or U9421 (N_9421,N_7969,N_6392);
nand U9422 (N_9422,N_6861,N_7868);
nor U9423 (N_9423,N_6768,N_6264);
nand U9424 (N_9424,N_6419,N_7029);
and U9425 (N_9425,N_6674,N_7754);
nand U9426 (N_9426,N_7292,N_7074);
or U9427 (N_9427,N_6038,N_7780);
and U9428 (N_9428,N_7106,N_6399);
nand U9429 (N_9429,N_6954,N_7549);
nand U9430 (N_9430,N_6238,N_7947);
nor U9431 (N_9431,N_6719,N_7635);
nand U9432 (N_9432,N_6597,N_6522);
nand U9433 (N_9433,N_7353,N_7404);
and U9434 (N_9434,N_6344,N_6474);
and U9435 (N_9435,N_6355,N_6126);
nand U9436 (N_9436,N_7778,N_7162);
or U9437 (N_9437,N_7236,N_7069);
nor U9438 (N_9438,N_6367,N_6638);
or U9439 (N_9439,N_7075,N_7009);
nand U9440 (N_9440,N_6248,N_7823);
and U9441 (N_9441,N_6742,N_6496);
nor U9442 (N_9442,N_6858,N_6575);
and U9443 (N_9443,N_6365,N_6439);
or U9444 (N_9444,N_7481,N_7131);
or U9445 (N_9445,N_6817,N_7103);
or U9446 (N_9446,N_7443,N_7848);
nor U9447 (N_9447,N_7135,N_6074);
nand U9448 (N_9448,N_6154,N_7743);
or U9449 (N_9449,N_7587,N_7515);
nand U9450 (N_9450,N_6047,N_7945);
nand U9451 (N_9451,N_6170,N_7593);
or U9452 (N_9452,N_7546,N_7916);
or U9453 (N_9453,N_7178,N_7577);
nor U9454 (N_9454,N_6326,N_6197);
or U9455 (N_9455,N_7544,N_6685);
nand U9456 (N_9456,N_7658,N_6846);
nand U9457 (N_9457,N_6961,N_7562);
nand U9458 (N_9458,N_7659,N_7492);
nand U9459 (N_9459,N_7389,N_7428);
nor U9460 (N_9460,N_7877,N_6167);
and U9461 (N_9461,N_6038,N_6063);
nor U9462 (N_9462,N_7755,N_6085);
nor U9463 (N_9463,N_7442,N_7497);
and U9464 (N_9464,N_6878,N_7923);
and U9465 (N_9465,N_7849,N_6788);
nand U9466 (N_9466,N_7223,N_6044);
or U9467 (N_9467,N_6290,N_6657);
nor U9468 (N_9468,N_6770,N_6765);
or U9469 (N_9469,N_6926,N_6265);
and U9470 (N_9470,N_7361,N_7778);
nor U9471 (N_9471,N_7883,N_7633);
nand U9472 (N_9472,N_6697,N_7823);
and U9473 (N_9473,N_6724,N_7309);
nand U9474 (N_9474,N_6262,N_6595);
xor U9475 (N_9475,N_6304,N_6592);
nor U9476 (N_9476,N_7485,N_7840);
and U9477 (N_9477,N_7042,N_6158);
and U9478 (N_9478,N_6890,N_7747);
and U9479 (N_9479,N_7066,N_7745);
or U9480 (N_9480,N_7165,N_6013);
or U9481 (N_9481,N_7188,N_7603);
and U9482 (N_9482,N_6508,N_6727);
or U9483 (N_9483,N_7868,N_6650);
and U9484 (N_9484,N_7837,N_6598);
nor U9485 (N_9485,N_7955,N_7670);
and U9486 (N_9486,N_7154,N_6935);
and U9487 (N_9487,N_6202,N_7945);
and U9488 (N_9488,N_7660,N_6287);
nor U9489 (N_9489,N_6635,N_6262);
xor U9490 (N_9490,N_7172,N_7245);
and U9491 (N_9491,N_6311,N_6654);
nand U9492 (N_9492,N_6240,N_6650);
nor U9493 (N_9493,N_7310,N_7462);
xnor U9494 (N_9494,N_7653,N_6577);
and U9495 (N_9495,N_7060,N_6601);
and U9496 (N_9496,N_7646,N_6152);
or U9497 (N_9497,N_7715,N_7661);
and U9498 (N_9498,N_7106,N_6312);
and U9499 (N_9499,N_7438,N_6437);
or U9500 (N_9500,N_7955,N_7739);
nor U9501 (N_9501,N_6669,N_7223);
or U9502 (N_9502,N_7858,N_7045);
nor U9503 (N_9503,N_6726,N_6125);
and U9504 (N_9504,N_6946,N_6505);
nor U9505 (N_9505,N_7857,N_7173);
or U9506 (N_9506,N_7990,N_6172);
nand U9507 (N_9507,N_6662,N_7134);
and U9508 (N_9508,N_7734,N_7372);
and U9509 (N_9509,N_7044,N_6995);
or U9510 (N_9510,N_7912,N_7427);
nand U9511 (N_9511,N_7333,N_6964);
and U9512 (N_9512,N_6483,N_6138);
and U9513 (N_9513,N_7085,N_7340);
or U9514 (N_9514,N_6320,N_7579);
nor U9515 (N_9515,N_7686,N_7767);
and U9516 (N_9516,N_6006,N_6674);
or U9517 (N_9517,N_6514,N_6692);
and U9518 (N_9518,N_6860,N_6904);
nor U9519 (N_9519,N_6729,N_6258);
nor U9520 (N_9520,N_7560,N_7153);
nor U9521 (N_9521,N_6560,N_6525);
nand U9522 (N_9522,N_6563,N_6820);
nand U9523 (N_9523,N_7226,N_6028);
and U9524 (N_9524,N_6888,N_6907);
xor U9525 (N_9525,N_7392,N_7968);
or U9526 (N_9526,N_7175,N_7613);
and U9527 (N_9527,N_6744,N_7071);
or U9528 (N_9528,N_7632,N_6481);
nand U9529 (N_9529,N_7443,N_7921);
nand U9530 (N_9530,N_7109,N_6835);
nor U9531 (N_9531,N_7887,N_7743);
or U9532 (N_9532,N_6364,N_7654);
and U9533 (N_9533,N_6629,N_6426);
nand U9534 (N_9534,N_6923,N_7173);
nor U9535 (N_9535,N_7177,N_7830);
or U9536 (N_9536,N_6931,N_6522);
nor U9537 (N_9537,N_7787,N_6371);
or U9538 (N_9538,N_6629,N_7971);
nor U9539 (N_9539,N_7130,N_7443);
or U9540 (N_9540,N_7947,N_6843);
nand U9541 (N_9541,N_6461,N_7285);
nand U9542 (N_9542,N_6738,N_7639);
nand U9543 (N_9543,N_7916,N_7268);
and U9544 (N_9544,N_7773,N_7951);
nor U9545 (N_9545,N_7303,N_7792);
nand U9546 (N_9546,N_7665,N_6180);
and U9547 (N_9547,N_7358,N_7408);
or U9548 (N_9548,N_7178,N_7347);
or U9549 (N_9549,N_6351,N_7211);
nand U9550 (N_9550,N_6208,N_6514);
xor U9551 (N_9551,N_7530,N_6126);
nor U9552 (N_9552,N_6443,N_6984);
nor U9553 (N_9553,N_6622,N_6053);
and U9554 (N_9554,N_6186,N_7092);
and U9555 (N_9555,N_7274,N_6680);
nand U9556 (N_9556,N_7984,N_7500);
nor U9557 (N_9557,N_6223,N_7731);
nor U9558 (N_9558,N_7583,N_6432);
nand U9559 (N_9559,N_7279,N_6236);
or U9560 (N_9560,N_6710,N_6839);
nor U9561 (N_9561,N_7871,N_7299);
and U9562 (N_9562,N_7710,N_7078);
or U9563 (N_9563,N_7013,N_6422);
nor U9564 (N_9564,N_6370,N_6952);
or U9565 (N_9565,N_6337,N_7666);
and U9566 (N_9566,N_7423,N_7580);
and U9567 (N_9567,N_6073,N_7220);
nor U9568 (N_9568,N_6918,N_6960);
or U9569 (N_9569,N_7777,N_6196);
xor U9570 (N_9570,N_7229,N_7287);
xnor U9571 (N_9571,N_7311,N_7685);
nand U9572 (N_9572,N_6249,N_6145);
nand U9573 (N_9573,N_6119,N_6366);
nor U9574 (N_9574,N_6655,N_6334);
or U9575 (N_9575,N_7088,N_6163);
nand U9576 (N_9576,N_6469,N_6164);
or U9577 (N_9577,N_7828,N_6847);
nor U9578 (N_9578,N_7746,N_7421);
and U9579 (N_9579,N_6969,N_7826);
or U9580 (N_9580,N_7187,N_6850);
nand U9581 (N_9581,N_6648,N_6244);
nor U9582 (N_9582,N_6303,N_6108);
nand U9583 (N_9583,N_7660,N_7672);
and U9584 (N_9584,N_6527,N_6632);
or U9585 (N_9585,N_6857,N_7015);
nand U9586 (N_9586,N_7627,N_7351);
nor U9587 (N_9587,N_6414,N_6299);
nand U9588 (N_9588,N_6353,N_6941);
nand U9589 (N_9589,N_6292,N_7638);
and U9590 (N_9590,N_7175,N_6135);
nor U9591 (N_9591,N_7002,N_7078);
and U9592 (N_9592,N_7815,N_7775);
nor U9593 (N_9593,N_7580,N_6230);
nor U9594 (N_9594,N_7059,N_7211);
and U9595 (N_9595,N_6336,N_7511);
nor U9596 (N_9596,N_6982,N_7424);
and U9597 (N_9597,N_7138,N_6358);
and U9598 (N_9598,N_6462,N_7656);
and U9599 (N_9599,N_7003,N_7891);
and U9600 (N_9600,N_6047,N_7853);
nor U9601 (N_9601,N_6723,N_6576);
nand U9602 (N_9602,N_7946,N_7598);
nor U9603 (N_9603,N_6480,N_7142);
or U9604 (N_9604,N_7728,N_6856);
or U9605 (N_9605,N_7780,N_6984);
nand U9606 (N_9606,N_6469,N_7024);
or U9607 (N_9607,N_6021,N_6631);
or U9608 (N_9608,N_7837,N_7555);
nor U9609 (N_9609,N_6840,N_7879);
nand U9610 (N_9610,N_6175,N_7504);
and U9611 (N_9611,N_6359,N_7995);
or U9612 (N_9612,N_6255,N_6198);
nor U9613 (N_9613,N_7368,N_7330);
and U9614 (N_9614,N_6642,N_6618);
nor U9615 (N_9615,N_7985,N_7145);
and U9616 (N_9616,N_6036,N_7305);
nor U9617 (N_9617,N_7693,N_6995);
nand U9618 (N_9618,N_7888,N_7425);
and U9619 (N_9619,N_7951,N_7836);
nand U9620 (N_9620,N_7142,N_6314);
or U9621 (N_9621,N_7235,N_7172);
and U9622 (N_9622,N_6704,N_7032);
nand U9623 (N_9623,N_6071,N_7100);
or U9624 (N_9624,N_6895,N_6114);
nor U9625 (N_9625,N_7704,N_6994);
nor U9626 (N_9626,N_6733,N_6985);
nor U9627 (N_9627,N_6980,N_7808);
nand U9628 (N_9628,N_6322,N_7174);
and U9629 (N_9629,N_6398,N_6981);
and U9630 (N_9630,N_7647,N_6192);
and U9631 (N_9631,N_7012,N_7607);
and U9632 (N_9632,N_6981,N_6995);
and U9633 (N_9633,N_6251,N_6221);
nor U9634 (N_9634,N_7704,N_7049);
nor U9635 (N_9635,N_7062,N_7234);
and U9636 (N_9636,N_6588,N_6178);
and U9637 (N_9637,N_6618,N_7842);
nor U9638 (N_9638,N_6425,N_7494);
or U9639 (N_9639,N_6957,N_6277);
and U9640 (N_9640,N_6936,N_6315);
or U9641 (N_9641,N_7143,N_6020);
and U9642 (N_9642,N_7987,N_7721);
or U9643 (N_9643,N_6215,N_6963);
or U9644 (N_9644,N_6198,N_7805);
and U9645 (N_9645,N_7477,N_7302);
nor U9646 (N_9646,N_7732,N_7501);
and U9647 (N_9647,N_6655,N_6353);
or U9648 (N_9648,N_7176,N_7883);
nand U9649 (N_9649,N_7386,N_7854);
or U9650 (N_9650,N_6439,N_7910);
and U9651 (N_9651,N_6170,N_6041);
or U9652 (N_9652,N_7982,N_6267);
and U9653 (N_9653,N_6829,N_7056);
and U9654 (N_9654,N_6405,N_7831);
or U9655 (N_9655,N_6589,N_6095);
xor U9656 (N_9656,N_6889,N_6633);
and U9657 (N_9657,N_7645,N_6507);
nor U9658 (N_9658,N_7634,N_6273);
or U9659 (N_9659,N_7007,N_6802);
and U9660 (N_9660,N_7625,N_7971);
nor U9661 (N_9661,N_6540,N_7216);
nand U9662 (N_9662,N_7671,N_6543);
nor U9663 (N_9663,N_6062,N_6493);
nor U9664 (N_9664,N_7757,N_6803);
nor U9665 (N_9665,N_6662,N_7600);
nor U9666 (N_9666,N_6791,N_6777);
nand U9667 (N_9667,N_7238,N_6295);
or U9668 (N_9668,N_6258,N_6450);
nor U9669 (N_9669,N_6412,N_6016);
nor U9670 (N_9670,N_6390,N_6394);
or U9671 (N_9671,N_6036,N_6695);
nand U9672 (N_9672,N_7250,N_6293);
nand U9673 (N_9673,N_6652,N_7327);
or U9674 (N_9674,N_7318,N_7831);
xnor U9675 (N_9675,N_6374,N_7750);
nand U9676 (N_9676,N_6927,N_7827);
and U9677 (N_9677,N_6256,N_7358);
or U9678 (N_9678,N_6919,N_7312);
nor U9679 (N_9679,N_7278,N_6577);
and U9680 (N_9680,N_7740,N_7661);
and U9681 (N_9681,N_6364,N_7485);
nand U9682 (N_9682,N_7743,N_7610);
nor U9683 (N_9683,N_7824,N_7762);
nor U9684 (N_9684,N_7805,N_7815);
and U9685 (N_9685,N_7271,N_7250);
nor U9686 (N_9686,N_6909,N_6500);
and U9687 (N_9687,N_6525,N_6673);
nor U9688 (N_9688,N_6991,N_7936);
nor U9689 (N_9689,N_6405,N_7169);
nand U9690 (N_9690,N_7209,N_6079);
and U9691 (N_9691,N_6059,N_7017);
and U9692 (N_9692,N_6717,N_6461);
or U9693 (N_9693,N_6817,N_6651);
nor U9694 (N_9694,N_7843,N_7877);
or U9695 (N_9695,N_6413,N_6918);
nor U9696 (N_9696,N_6200,N_7396);
nor U9697 (N_9697,N_7122,N_6418);
nand U9698 (N_9698,N_6414,N_6175);
or U9699 (N_9699,N_6374,N_6522);
nand U9700 (N_9700,N_7348,N_6485);
and U9701 (N_9701,N_6624,N_6528);
nand U9702 (N_9702,N_6822,N_7794);
and U9703 (N_9703,N_6998,N_6050);
nor U9704 (N_9704,N_6619,N_6357);
and U9705 (N_9705,N_7399,N_6869);
or U9706 (N_9706,N_6479,N_7408);
or U9707 (N_9707,N_7939,N_7138);
or U9708 (N_9708,N_7281,N_7676);
nor U9709 (N_9709,N_7771,N_7261);
or U9710 (N_9710,N_6113,N_7384);
nor U9711 (N_9711,N_6657,N_6437);
nand U9712 (N_9712,N_6781,N_7626);
and U9713 (N_9713,N_7800,N_7738);
nand U9714 (N_9714,N_6733,N_7471);
nand U9715 (N_9715,N_7032,N_7324);
xnor U9716 (N_9716,N_6468,N_6259);
or U9717 (N_9717,N_7046,N_6637);
nor U9718 (N_9718,N_7408,N_7898);
nor U9719 (N_9719,N_6912,N_7545);
nor U9720 (N_9720,N_6039,N_7978);
and U9721 (N_9721,N_6666,N_6580);
and U9722 (N_9722,N_6543,N_7788);
and U9723 (N_9723,N_6677,N_7462);
nand U9724 (N_9724,N_6831,N_7053);
nand U9725 (N_9725,N_7548,N_7208);
nor U9726 (N_9726,N_6842,N_7791);
nand U9727 (N_9727,N_6997,N_6599);
and U9728 (N_9728,N_7506,N_6095);
and U9729 (N_9729,N_6351,N_7581);
and U9730 (N_9730,N_6414,N_6811);
nor U9731 (N_9731,N_6037,N_7781);
or U9732 (N_9732,N_6000,N_7397);
or U9733 (N_9733,N_7349,N_6012);
or U9734 (N_9734,N_6344,N_6312);
nor U9735 (N_9735,N_6737,N_6975);
xnor U9736 (N_9736,N_6430,N_6911);
nor U9737 (N_9737,N_7243,N_7985);
nor U9738 (N_9738,N_6841,N_6679);
and U9739 (N_9739,N_7853,N_6092);
or U9740 (N_9740,N_7760,N_7311);
nor U9741 (N_9741,N_6052,N_7622);
and U9742 (N_9742,N_7410,N_7652);
nor U9743 (N_9743,N_6090,N_6716);
and U9744 (N_9744,N_7773,N_6717);
nand U9745 (N_9745,N_7421,N_6054);
and U9746 (N_9746,N_6273,N_7238);
nand U9747 (N_9747,N_6743,N_6715);
and U9748 (N_9748,N_6216,N_6393);
and U9749 (N_9749,N_6991,N_7459);
nor U9750 (N_9750,N_7744,N_6141);
xor U9751 (N_9751,N_7690,N_7451);
or U9752 (N_9752,N_6781,N_7498);
and U9753 (N_9753,N_6494,N_7036);
and U9754 (N_9754,N_6119,N_6698);
nor U9755 (N_9755,N_6371,N_7927);
or U9756 (N_9756,N_7081,N_6182);
nand U9757 (N_9757,N_7651,N_6858);
and U9758 (N_9758,N_6133,N_6441);
and U9759 (N_9759,N_7871,N_7071);
and U9760 (N_9760,N_7247,N_6775);
nor U9761 (N_9761,N_7102,N_6145);
or U9762 (N_9762,N_6085,N_6570);
or U9763 (N_9763,N_7086,N_7051);
nand U9764 (N_9764,N_6103,N_6968);
and U9765 (N_9765,N_7468,N_7850);
nand U9766 (N_9766,N_7397,N_7858);
and U9767 (N_9767,N_7226,N_7398);
nor U9768 (N_9768,N_6942,N_6499);
nand U9769 (N_9769,N_7792,N_6431);
and U9770 (N_9770,N_7183,N_6549);
or U9771 (N_9771,N_7185,N_6555);
nand U9772 (N_9772,N_7860,N_7359);
nor U9773 (N_9773,N_6800,N_6114);
nand U9774 (N_9774,N_6192,N_7879);
nor U9775 (N_9775,N_7332,N_6754);
xor U9776 (N_9776,N_6339,N_6484);
nor U9777 (N_9777,N_7213,N_6347);
or U9778 (N_9778,N_7208,N_7141);
nor U9779 (N_9779,N_6819,N_6457);
and U9780 (N_9780,N_7589,N_7891);
nor U9781 (N_9781,N_7620,N_6630);
xnor U9782 (N_9782,N_6987,N_6998);
nand U9783 (N_9783,N_7254,N_6384);
or U9784 (N_9784,N_6574,N_7278);
nor U9785 (N_9785,N_6955,N_6737);
nor U9786 (N_9786,N_6533,N_7574);
or U9787 (N_9787,N_6990,N_7148);
and U9788 (N_9788,N_6058,N_6688);
and U9789 (N_9789,N_6455,N_7111);
nor U9790 (N_9790,N_7609,N_6576);
and U9791 (N_9791,N_6169,N_6195);
or U9792 (N_9792,N_6932,N_7211);
and U9793 (N_9793,N_6163,N_7160);
nor U9794 (N_9794,N_7911,N_6557);
nor U9795 (N_9795,N_6212,N_7732);
nor U9796 (N_9796,N_7056,N_6139);
or U9797 (N_9797,N_6284,N_6399);
nand U9798 (N_9798,N_6178,N_6340);
nand U9799 (N_9799,N_7396,N_6137);
and U9800 (N_9800,N_6290,N_7960);
nand U9801 (N_9801,N_7495,N_7319);
nor U9802 (N_9802,N_7891,N_6643);
or U9803 (N_9803,N_6865,N_6610);
and U9804 (N_9804,N_7775,N_6979);
nor U9805 (N_9805,N_6962,N_6289);
nor U9806 (N_9806,N_7291,N_6192);
and U9807 (N_9807,N_6514,N_7258);
nor U9808 (N_9808,N_7187,N_6739);
or U9809 (N_9809,N_6790,N_7095);
nand U9810 (N_9810,N_7476,N_6897);
xnor U9811 (N_9811,N_6548,N_7482);
and U9812 (N_9812,N_6091,N_6098);
nor U9813 (N_9813,N_7132,N_7617);
and U9814 (N_9814,N_6301,N_6105);
or U9815 (N_9815,N_6099,N_6410);
nand U9816 (N_9816,N_6410,N_6836);
nor U9817 (N_9817,N_7056,N_7352);
and U9818 (N_9818,N_7862,N_6597);
or U9819 (N_9819,N_7581,N_7672);
or U9820 (N_9820,N_7438,N_7049);
and U9821 (N_9821,N_7818,N_6705);
nor U9822 (N_9822,N_6878,N_7607);
and U9823 (N_9823,N_7809,N_7354);
nand U9824 (N_9824,N_7755,N_7664);
or U9825 (N_9825,N_7344,N_7919);
and U9826 (N_9826,N_7765,N_6195);
nand U9827 (N_9827,N_7194,N_6631);
nor U9828 (N_9828,N_7339,N_7718);
and U9829 (N_9829,N_6649,N_7335);
nand U9830 (N_9830,N_6725,N_7080);
nor U9831 (N_9831,N_6825,N_6910);
and U9832 (N_9832,N_7462,N_7613);
nor U9833 (N_9833,N_6780,N_6309);
or U9834 (N_9834,N_7236,N_6672);
nand U9835 (N_9835,N_6669,N_6848);
nor U9836 (N_9836,N_7397,N_6521);
and U9837 (N_9837,N_6147,N_7314);
nand U9838 (N_9838,N_7735,N_6605);
nor U9839 (N_9839,N_7800,N_7099);
nand U9840 (N_9840,N_6606,N_7618);
nor U9841 (N_9841,N_6506,N_7309);
nor U9842 (N_9842,N_6498,N_6343);
and U9843 (N_9843,N_6655,N_7583);
or U9844 (N_9844,N_6969,N_6497);
or U9845 (N_9845,N_7257,N_7520);
nand U9846 (N_9846,N_7129,N_7592);
nand U9847 (N_9847,N_7763,N_6043);
nor U9848 (N_9848,N_7785,N_7113);
and U9849 (N_9849,N_6505,N_7881);
nor U9850 (N_9850,N_6683,N_7125);
nand U9851 (N_9851,N_6637,N_7578);
or U9852 (N_9852,N_7346,N_6939);
and U9853 (N_9853,N_6312,N_6995);
nand U9854 (N_9854,N_6109,N_6439);
nor U9855 (N_9855,N_7496,N_6538);
xor U9856 (N_9856,N_7518,N_7164);
xnor U9857 (N_9857,N_6415,N_7630);
nand U9858 (N_9858,N_7392,N_6392);
or U9859 (N_9859,N_6209,N_6920);
or U9860 (N_9860,N_6620,N_7825);
nand U9861 (N_9861,N_6490,N_6618);
and U9862 (N_9862,N_7268,N_7628);
nand U9863 (N_9863,N_7083,N_7084);
nor U9864 (N_9864,N_7609,N_7748);
and U9865 (N_9865,N_7887,N_7111);
and U9866 (N_9866,N_6138,N_7485);
nand U9867 (N_9867,N_6044,N_6654);
nand U9868 (N_9868,N_6453,N_7381);
or U9869 (N_9869,N_7371,N_7356);
nand U9870 (N_9870,N_6356,N_7747);
nand U9871 (N_9871,N_6067,N_7417);
xor U9872 (N_9872,N_6262,N_6400);
nand U9873 (N_9873,N_6589,N_6537);
and U9874 (N_9874,N_6450,N_6932);
nor U9875 (N_9875,N_6501,N_6181);
and U9876 (N_9876,N_6313,N_6565);
and U9877 (N_9877,N_6960,N_6101);
nand U9878 (N_9878,N_6905,N_6697);
nor U9879 (N_9879,N_6198,N_6135);
or U9880 (N_9880,N_6834,N_7940);
and U9881 (N_9881,N_6581,N_6584);
nor U9882 (N_9882,N_7339,N_6561);
or U9883 (N_9883,N_6263,N_6570);
or U9884 (N_9884,N_7850,N_7066);
nor U9885 (N_9885,N_7246,N_7602);
nand U9886 (N_9886,N_7091,N_7786);
and U9887 (N_9887,N_6784,N_6952);
or U9888 (N_9888,N_6453,N_6843);
and U9889 (N_9889,N_7855,N_7045);
nand U9890 (N_9890,N_6147,N_7984);
or U9891 (N_9891,N_6033,N_7422);
or U9892 (N_9892,N_6188,N_7664);
nand U9893 (N_9893,N_6136,N_6122);
nand U9894 (N_9894,N_6668,N_6236);
and U9895 (N_9895,N_7121,N_7574);
or U9896 (N_9896,N_6204,N_6386);
and U9897 (N_9897,N_6571,N_6792);
and U9898 (N_9898,N_7412,N_7138);
and U9899 (N_9899,N_7601,N_7502);
or U9900 (N_9900,N_7437,N_6896);
nand U9901 (N_9901,N_7593,N_7306);
nor U9902 (N_9902,N_7067,N_7584);
or U9903 (N_9903,N_7298,N_7457);
nand U9904 (N_9904,N_6725,N_7323);
or U9905 (N_9905,N_7187,N_6704);
xor U9906 (N_9906,N_6119,N_7313);
nand U9907 (N_9907,N_7806,N_7260);
nor U9908 (N_9908,N_7621,N_6023);
and U9909 (N_9909,N_6062,N_7048);
or U9910 (N_9910,N_6454,N_7436);
or U9911 (N_9911,N_7242,N_7596);
and U9912 (N_9912,N_7496,N_6864);
and U9913 (N_9913,N_6507,N_6032);
nand U9914 (N_9914,N_7632,N_6702);
nand U9915 (N_9915,N_6036,N_7075);
or U9916 (N_9916,N_7646,N_6263);
and U9917 (N_9917,N_6045,N_6793);
nand U9918 (N_9918,N_7618,N_6005);
nand U9919 (N_9919,N_6942,N_6209);
or U9920 (N_9920,N_6944,N_7538);
or U9921 (N_9921,N_7733,N_7344);
nand U9922 (N_9922,N_6209,N_7162);
or U9923 (N_9923,N_6899,N_7047);
nand U9924 (N_9924,N_7626,N_7176);
and U9925 (N_9925,N_6945,N_6156);
or U9926 (N_9926,N_6637,N_6295);
and U9927 (N_9927,N_7365,N_7799);
nor U9928 (N_9928,N_7276,N_7260);
or U9929 (N_9929,N_7577,N_7492);
or U9930 (N_9930,N_6109,N_6885);
or U9931 (N_9931,N_7169,N_7166);
and U9932 (N_9932,N_7878,N_7353);
nand U9933 (N_9933,N_6726,N_6728);
nand U9934 (N_9934,N_7945,N_6266);
and U9935 (N_9935,N_6941,N_7784);
or U9936 (N_9936,N_7903,N_6215);
nor U9937 (N_9937,N_7084,N_7422);
or U9938 (N_9938,N_6527,N_7880);
nor U9939 (N_9939,N_6575,N_6832);
and U9940 (N_9940,N_6989,N_6017);
nand U9941 (N_9941,N_7467,N_7206);
nand U9942 (N_9942,N_6463,N_7780);
or U9943 (N_9943,N_6186,N_6572);
or U9944 (N_9944,N_7512,N_7209);
xnor U9945 (N_9945,N_7369,N_7195);
xor U9946 (N_9946,N_6013,N_7936);
and U9947 (N_9947,N_7389,N_6961);
or U9948 (N_9948,N_7886,N_7699);
nor U9949 (N_9949,N_7780,N_7751);
and U9950 (N_9950,N_6451,N_6824);
or U9951 (N_9951,N_7933,N_7626);
or U9952 (N_9952,N_7446,N_6004);
nor U9953 (N_9953,N_6377,N_7341);
nand U9954 (N_9954,N_7123,N_6623);
nor U9955 (N_9955,N_7671,N_7361);
nand U9956 (N_9956,N_6677,N_7417);
or U9957 (N_9957,N_6083,N_6530);
and U9958 (N_9958,N_7341,N_7247);
nor U9959 (N_9959,N_6552,N_7677);
or U9960 (N_9960,N_7275,N_7627);
and U9961 (N_9961,N_6038,N_6817);
nand U9962 (N_9962,N_7438,N_6417);
or U9963 (N_9963,N_7785,N_6058);
nand U9964 (N_9964,N_6172,N_7178);
nand U9965 (N_9965,N_6093,N_6728);
nor U9966 (N_9966,N_6886,N_6252);
nor U9967 (N_9967,N_7192,N_7385);
nor U9968 (N_9968,N_6214,N_6436);
nand U9969 (N_9969,N_6857,N_7600);
and U9970 (N_9970,N_6399,N_7221);
xor U9971 (N_9971,N_7020,N_6863);
nor U9972 (N_9972,N_7505,N_6617);
xnor U9973 (N_9973,N_6042,N_7847);
and U9974 (N_9974,N_6754,N_7197);
nor U9975 (N_9975,N_6526,N_6854);
or U9976 (N_9976,N_6948,N_6170);
nand U9977 (N_9977,N_6087,N_7597);
nor U9978 (N_9978,N_7591,N_6986);
and U9979 (N_9979,N_6918,N_6420);
or U9980 (N_9980,N_6193,N_6155);
nand U9981 (N_9981,N_7799,N_7618);
nor U9982 (N_9982,N_7295,N_6654);
or U9983 (N_9983,N_7136,N_6672);
and U9984 (N_9984,N_7831,N_6745);
or U9985 (N_9985,N_6378,N_7561);
nor U9986 (N_9986,N_6314,N_6673);
nand U9987 (N_9987,N_6027,N_6517);
and U9988 (N_9988,N_7441,N_6594);
nand U9989 (N_9989,N_6064,N_6072);
nor U9990 (N_9990,N_7022,N_6940);
nand U9991 (N_9991,N_6030,N_6890);
nand U9992 (N_9992,N_6965,N_6815);
or U9993 (N_9993,N_6738,N_6158);
nor U9994 (N_9994,N_6277,N_7409);
nor U9995 (N_9995,N_7251,N_7356);
nand U9996 (N_9996,N_6259,N_6334);
nor U9997 (N_9997,N_7373,N_6381);
and U9998 (N_9998,N_6720,N_7456);
and U9999 (N_9999,N_7467,N_7349);
nand UO_0 (O_0,N_9519,N_8295);
nor UO_1 (O_1,N_9407,N_9740);
or UO_2 (O_2,N_9548,N_8912);
nor UO_3 (O_3,N_8302,N_8571);
and UO_4 (O_4,N_9493,N_9172);
xnor UO_5 (O_5,N_9244,N_9657);
or UO_6 (O_6,N_9863,N_9791);
or UO_7 (O_7,N_9742,N_8144);
nor UO_8 (O_8,N_9369,N_8921);
and UO_9 (O_9,N_9653,N_9646);
nor UO_10 (O_10,N_8748,N_8862);
nand UO_11 (O_11,N_8187,N_8966);
xor UO_12 (O_12,N_9212,N_9660);
nor UO_13 (O_13,N_8611,N_9809);
or UO_14 (O_14,N_8873,N_9403);
or UO_15 (O_15,N_9040,N_9089);
or UO_16 (O_16,N_8035,N_9192);
or UO_17 (O_17,N_8657,N_8037);
xor UO_18 (O_18,N_9782,N_8649);
nor UO_19 (O_19,N_8304,N_9434);
or UO_20 (O_20,N_8797,N_8338);
and UO_21 (O_21,N_9523,N_8936);
and UO_22 (O_22,N_8301,N_9537);
and UO_23 (O_23,N_9639,N_9303);
or UO_24 (O_24,N_9920,N_8993);
or UO_25 (O_25,N_8164,N_9743);
nand UO_26 (O_26,N_8746,N_8360);
or UO_27 (O_27,N_9812,N_9534);
nor UO_28 (O_28,N_9643,N_9163);
or UO_29 (O_29,N_9905,N_9277);
nor UO_30 (O_30,N_9227,N_9363);
and UO_31 (O_31,N_9293,N_9087);
nand UO_32 (O_32,N_9855,N_9757);
nand UO_33 (O_33,N_8800,N_8781);
nor UO_34 (O_34,N_8169,N_9746);
and UO_35 (O_35,N_8305,N_9845);
or UO_36 (O_36,N_8745,N_9268);
nor UO_37 (O_37,N_9883,N_8581);
nand UO_38 (O_38,N_8809,N_8947);
nand UO_39 (O_39,N_8499,N_8109);
or UO_40 (O_40,N_9627,N_9889);
nand UO_41 (O_41,N_9980,N_9781);
nor UO_42 (O_42,N_9335,N_9432);
and UO_43 (O_43,N_9825,N_8510);
or UO_44 (O_44,N_8971,N_8630);
and UO_45 (O_45,N_9551,N_8703);
nor UO_46 (O_46,N_9157,N_9998);
and UO_47 (O_47,N_9071,N_8551);
nor UO_48 (O_48,N_9839,N_8944);
nand UO_49 (O_49,N_8776,N_9304);
nor UO_50 (O_50,N_8612,N_9535);
xnor UO_51 (O_51,N_9923,N_9602);
and UO_52 (O_52,N_9215,N_9490);
nand UO_53 (O_53,N_8167,N_9704);
nor UO_54 (O_54,N_9968,N_8048);
and UO_55 (O_55,N_8973,N_8440);
or UO_56 (O_56,N_9271,N_9794);
or UO_57 (O_57,N_8885,N_9961);
and UO_58 (O_58,N_8521,N_8516);
nor UO_59 (O_59,N_8327,N_9665);
and UO_60 (O_60,N_9651,N_8369);
nand UO_61 (O_61,N_8057,N_9895);
nor UO_62 (O_62,N_9934,N_8892);
or UO_63 (O_63,N_8165,N_8861);
or UO_64 (O_64,N_8455,N_8962);
nand UO_65 (O_65,N_9382,N_9378);
nor UO_66 (O_66,N_9406,N_9722);
or UO_67 (O_67,N_8215,N_8420);
and UO_68 (O_68,N_8867,N_8595);
xor UO_69 (O_69,N_9272,N_9582);
or UO_70 (O_70,N_8284,N_9566);
and UO_71 (O_71,N_8162,N_8210);
nor UO_72 (O_72,N_9255,N_9978);
nor UO_73 (O_73,N_8832,N_9579);
nor UO_74 (O_74,N_9321,N_8489);
or UO_75 (O_75,N_9325,N_9001);
or UO_76 (O_76,N_9530,N_8391);
nor UO_77 (O_77,N_8761,N_8193);
xnor UO_78 (O_78,N_9195,N_9360);
nor UO_79 (O_79,N_9836,N_9636);
xor UO_80 (O_80,N_9066,N_9715);
or UO_81 (O_81,N_9750,N_8474);
or UO_82 (O_82,N_8254,N_8032);
or UO_83 (O_83,N_8352,N_9739);
or UO_84 (O_84,N_8730,N_9465);
nor UO_85 (O_85,N_9332,N_8677);
nand UO_86 (O_86,N_9572,N_8212);
and UO_87 (O_87,N_9090,N_8805);
and UO_88 (O_88,N_9785,N_8206);
or UO_89 (O_89,N_9076,N_8505);
nor UO_90 (O_90,N_8839,N_8774);
and UO_91 (O_91,N_8603,N_8874);
nor UO_92 (O_92,N_8398,N_9614);
or UO_93 (O_93,N_8722,N_8726);
or UO_94 (O_94,N_8752,N_9446);
and UO_95 (O_95,N_9494,N_9786);
nor UO_96 (O_96,N_8158,N_8219);
nand UO_97 (O_97,N_9435,N_8729);
nor UO_98 (O_98,N_9638,N_9858);
and UO_99 (O_99,N_9240,N_8299);
nand UO_100 (O_100,N_8423,N_8765);
or UO_101 (O_101,N_8685,N_9184);
and UO_102 (O_102,N_9034,N_9995);
nor UO_103 (O_103,N_8842,N_9075);
nand UO_104 (O_104,N_8552,N_9754);
or UO_105 (O_105,N_9984,N_8363);
xor UO_106 (O_106,N_9028,N_8593);
and UO_107 (O_107,N_8564,N_9874);
nand UO_108 (O_108,N_9868,N_9104);
and UO_109 (O_109,N_8740,N_8655);
or UO_110 (O_110,N_8239,N_9383);
nand UO_111 (O_111,N_8633,N_8563);
nor UO_112 (O_112,N_8848,N_8309);
nand UO_113 (O_113,N_8123,N_9591);
or UO_114 (O_114,N_8869,N_8487);
xor UO_115 (O_115,N_9402,N_8427);
nor UO_116 (O_116,N_8207,N_8555);
nand UO_117 (O_117,N_9395,N_9064);
and UO_118 (O_118,N_9205,N_9211);
nor UO_119 (O_119,N_8733,N_9928);
nand UO_120 (O_120,N_8412,N_9840);
nand UO_121 (O_121,N_9916,N_8393);
and UO_122 (O_122,N_9124,N_8188);
and UO_123 (O_123,N_8897,N_9849);
nor UO_124 (O_124,N_9732,N_8335);
or UO_125 (O_125,N_8246,N_9831);
or UO_126 (O_126,N_8775,N_9977);
nor UO_127 (O_127,N_8168,N_8434);
nor UO_128 (O_128,N_8233,N_8678);
nor UO_129 (O_129,N_9964,N_9941);
nor UO_130 (O_130,N_8846,N_9527);
or UO_131 (O_131,N_9570,N_9381);
nor UO_132 (O_132,N_9476,N_9733);
nand UO_133 (O_133,N_8705,N_8736);
nor UO_134 (O_134,N_8528,N_8609);
nand UO_135 (O_135,N_8969,N_8511);
nor UO_136 (O_136,N_9896,N_9899);
and UO_137 (O_137,N_8602,N_9397);
or UO_138 (O_138,N_8791,N_9426);
nor UO_139 (O_139,N_9654,N_8985);
nand UO_140 (O_140,N_9692,N_8712);
nor UO_141 (O_141,N_8665,N_8371);
and UO_142 (O_142,N_8941,N_8990);
and UO_143 (O_143,N_9241,N_8131);
nand UO_144 (O_144,N_9190,N_8699);
nor UO_145 (O_145,N_8222,N_9596);
nor UO_146 (O_146,N_8554,N_8461);
or UO_147 (O_147,N_8700,N_9738);
and UO_148 (O_148,N_8820,N_9698);
and UO_149 (O_149,N_9857,N_9433);
nand UO_150 (O_150,N_8436,N_8813);
or UO_151 (O_151,N_8640,N_9324);
and UO_152 (O_152,N_9982,N_9186);
nand UO_153 (O_153,N_9790,N_8586);
or UO_154 (O_154,N_8606,N_9776);
nand UO_155 (O_155,N_8545,N_9078);
and UO_156 (O_156,N_9800,N_8515);
or UO_157 (O_157,N_8961,N_8069);
nand UO_158 (O_158,N_8986,N_9218);
nor UO_159 (O_159,N_9538,N_8597);
or UO_160 (O_160,N_8448,N_9228);
nand UO_161 (O_161,N_8672,N_8179);
nor UO_162 (O_162,N_8946,N_8843);
or UO_163 (O_163,N_9118,N_8468);
nor UO_164 (O_164,N_9972,N_9237);
or UO_165 (O_165,N_8670,N_8428);
or UO_166 (O_166,N_8875,N_8263);
or UO_167 (O_167,N_9238,N_9827);
nor UO_168 (O_168,N_8014,N_8098);
and UO_169 (O_169,N_9346,N_9290);
nand UO_170 (O_170,N_8177,N_9055);
nand UO_171 (O_171,N_9209,N_9930);
nor UO_172 (O_172,N_9488,N_8668);
nor UO_173 (O_173,N_8697,N_9142);
and UO_174 (O_174,N_8830,N_9243);
and UO_175 (O_175,N_9297,N_8856);
nand UO_176 (O_176,N_8495,N_9497);
or UO_177 (O_177,N_9664,N_8326);
and UO_178 (O_178,N_9291,N_8824);
nor UO_179 (O_179,N_9338,N_9510);
nand UO_180 (O_180,N_9234,N_9187);
or UO_181 (O_181,N_9761,N_8536);
nor UO_182 (O_182,N_8804,N_8099);
or UO_183 (O_183,N_9797,N_9684);
nand UO_184 (O_184,N_9992,N_8477);
and UO_185 (O_185,N_9901,N_8562);
nand UO_186 (O_186,N_9856,N_8561);
nor UO_187 (O_187,N_8084,N_8227);
and UO_188 (O_188,N_9261,N_9128);
nor UO_189 (O_189,N_9460,N_8818);
nand UO_190 (O_190,N_9219,N_8339);
and UO_191 (O_191,N_9808,N_9966);
nor UO_192 (O_192,N_9342,N_9796);
xnor UO_193 (O_193,N_8955,N_9137);
nand UO_194 (O_194,N_9189,N_9015);
or UO_195 (O_195,N_9178,N_9216);
nand UO_196 (O_196,N_8321,N_9278);
and UO_197 (O_197,N_8808,N_9037);
nor UO_198 (O_198,N_9613,N_9960);
nand UO_199 (O_199,N_8506,N_8568);
and UO_200 (O_200,N_9140,N_9070);
and UO_201 (O_201,N_9852,N_8421);
and UO_202 (O_202,N_8977,N_8180);
nor UO_203 (O_203,N_9046,N_8322);
and UO_204 (O_204,N_9221,N_8980);
nand UO_205 (O_205,N_8275,N_9604);
nor UO_206 (O_206,N_8900,N_8402);
and UO_207 (O_207,N_9181,N_9688);
or UO_208 (O_208,N_9152,N_8934);
nand UO_209 (O_209,N_9640,N_8930);
nand UO_210 (O_210,N_9377,N_9105);
and UO_211 (O_211,N_9439,N_8807);
nor UO_212 (O_212,N_8950,N_9632);
and UO_213 (O_213,N_8509,N_9807);
xor UO_214 (O_214,N_8323,N_9597);
nand UO_215 (O_215,N_8992,N_8949);
xor UO_216 (O_216,N_9100,N_9479);
or UO_217 (O_217,N_8520,N_8894);
and UO_218 (O_218,N_9888,N_9296);
and UO_219 (O_219,N_9929,N_9714);
nor UO_220 (O_220,N_8294,N_9410);
and UO_221 (O_221,N_9544,N_9884);
nor UO_222 (O_222,N_8674,N_8376);
or UO_223 (O_223,N_8134,N_8952);
xor UO_224 (O_224,N_9974,N_9116);
nor UO_225 (O_225,N_8447,N_9663);
and UO_226 (O_226,N_9667,N_8956);
nor UO_227 (O_227,N_8981,N_9676);
nor UO_228 (O_228,N_9220,N_8261);
and UO_229 (O_229,N_9292,N_9173);
or UO_230 (O_230,N_8285,N_8580);
nor UO_231 (O_231,N_9991,N_8147);
nor UO_232 (O_232,N_8146,N_8715);
nor UO_233 (O_233,N_8105,N_9576);
xnor UO_234 (O_234,N_8837,N_9083);
nand UO_235 (O_235,N_9322,N_8163);
nor UO_236 (O_236,N_9354,N_8145);
or UO_237 (O_237,N_8415,N_8344);
and UO_238 (O_238,N_8409,N_9803);
and UO_239 (O_239,N_8160,N_8850);
nand UO_240 (O_240,N_8313,N_8074);
and UO_241 (O_241,N_8693,N_9489);
xor UO_242 (O_242,N_9758,N_8358);
xnor UO_243 (O_243,N_8410,N_8132);
and UO_244 (O_244,N_9623,N_8799);
nor UO_245 (O_245,N_9760,N_9133);
and UO_246 (O_246,N_8435,N_9280);
and UO_247 (O_247,N_8021,N_9230);
and UO_248 (O_248,N_9343,N_8334);
nor UO_249 (O_249,N_8978,N_8919);
and UO_250 (O_250,N_8368,N_9699);
or UO_251 (O_251,N_8664,N_9029);
and UO_252 (O_252,N_9557,N_8652);
and UO_253 (O_253,N_8011,N_9609);
and UO_254 (O_254,N_9107,N_9771);
or UO_255 (O_255,N_9482,N_8333);
and UO_256 (O_256,N_9666,N_9817);
and UO_257 (O_257,N_8001,N_9717);
and UO_258 (O_258,N_8248,N_9906);
and UO_259 (O_259,N_9198,N_9298);
nor UO_260 (O_260,N_9952,N_9486);
nor UO_261 (O_261,N_9353,N_9917);
nand UO_262 (O_262,N_8152,N_9824);
nor UO_263 (O_263,N_9775,N_9429);
and UO_264 (O_264,N_8538,N_9097);
nor UO_265 (O_265,N_9415,N_8596);
and UO_266 (O_266,N_8346,N_8111);
nor UO_267 (O_267,N_9314,N_8493);
or UO_268 (O_268,N_8221,N_8871);
or UO_269 (O_269,N_8046,N_9861);
nand UO_270 (O_270,N_8567,N_9787);
or UO_271 (O_271,N_8548,N_8078);
or UO_272 (O_272,N_8779,N_9832);
or UO_273 (O_273,N_8938,N_9970);
nor UO_274 (O_274,N_8267,N_8063);
or UO_275 (O_275,N_8728,N_8470);
or UO_276 (O_276,N_9512,N_8385);
nand UO_277 (O_277,N_8269,N_9119);
nor UO_278 (O_278,N_9235,N_9351);
nand UO_279 (O_279,N_9263,N_9110);
nor UO_280 (O_280,N_9645,N_8795);
nor UO_281 (O_281,N_9958,N_8137);
nand UO_282 (O_282,N_9449,N_8406);
or UO_283 (O_283,N_8810,N_8546);
nor UO_284 (O_284,N_9870,N_9724);
nand UO_285 (O_285,N_9532,N_9223);
and UO_286 (O_286,N_8324,N_8059);
and UO_287 (O_287,N_8345,N_8072);
or UO_288 (O_288,N_9180,N_8095);
nor UO_289 (O_289,N_8384,N_9368);
nor UO_290 (O_290,N_9169,N_8920);
nand UO_291 (O_291,N_9553,N_8517);
and UO_292 (O_292,N_9391,N_8082);
or UO_293 (O_293,N_9253,N_9678);
or UO_294 (O_294,N_9096,N_9748);
and UO_295 (O_295,N_9601,N_8300);
or UO_296 (O_296,N_9965,N_9860);
nand UO_297 (O_297,N_9333,N_8401);
nand UO_298 (O_298,N_8598,N_8311);
or UO_299 (O_299,N_9248,N_8646);
and UO_300 (O_300,N_8620,N_9751);
and UO_301 (O_301,N_9686,N_8821);
nor UO_302 (O_302,N_8120,N_9979);
nor UO_303 (O_303,N_8058,N_9561);
nor UO_304 (O_304,N_9252,N_9203);
nand UO_305 (O_305,N_9649,N_9127);
xor UO_306 (O_306,N_9508,N_9162);
and UO_307 (O_307,N_9681,N_8594);
or UO_308 (O_308,N_8692,N_9361);
or UO_309 (O_309,N_8783,N_9072);
nand UO_310 (O_310,N_8130,N_9425);
and UO_311 (O_311,N_8236,N_9607);
or UO_312 (O_312,N_9295,N_9113);
nand UO_313 (O_313,N_8656,N_8784);
or UO_314 (O_314,N_8591,N_8836);
nor UO_315 (O_315,N_8866,N_8342);
nand UO_316 (O_316,N_9661,N_9320);
or UO_317 (O_317,N_8577,N_9515);
nand UO_318 (O_318,N_8708,N_8631);
or UO_319 (O_319,N_9364,N_9370);
nand UO_320 (O_320,N_8354,N_9080);
nand UO_321 (O_321,N_8004,N_8676);
nor UO_322 (O_322,N_9329,N_9495);
nand UO_323 (O_323,N_9996,N_8068);
nand UO_324 (O_324,N_8768,N_8079);
nor UO_325 (O_325,N_9625,N_8191);
and UO_326 (O_326,N_8259,N_8876);
nand UO_327 (O_327,N_9583,N_9554);
nor UO_328 (O_328,N_8007,N_8583);
nor UO_329 (O_329,N_9466,N_8793);
nand UO_330 (O_330,N_8653,N_8484);
nand UO_331 (O_331,N_9158,N_9062);
or UO_332 (O_332,N_9716,N_8588);
nor UO_333 (O_333,N_9741,N_9662);
or UO_334 (O_334,N_8426,N_8033);
nor UO_335 (O_335,N_8174,N_9975);
or UO_336 (O_336,N_9229,N_8296);
nor UO_337 (O_337,N_8743,N_9111);
nor UO_338 (O_338,N_9086,N_9441);
nor UO_339 (O_339,N_9835,N_8518);
xnor UO_340 (O_340,N_9409,N_8457);
or UO_341 (O_341,N_8318,N_8245);
nor UO_342 (O_342,N_8887,N_8560);
or UO_343 (O_343,N_9848,N_9683);
or UO_344 (O_344,N_9559,N_8929);
and UO_345 (O_345,N_8332,N_8018);
nor UO_346 (O_346,N_9438,N_8811);
or UO_347 (O_347,N_9079,N_8757);
and UO_348 (O_348,N_9050,N_9287);
nor UO_349 (O_349,N_8417,N_9430);
nand UO_350 (O_350,N_9918,N_8009);
nand UO_351 (O_351,N_9872,N_8140);
and UO_352 (O_352,N_8899,N_8159);
and UO_353 (O_353,N_8075,N_9174);
and UO_354 (O_354,N_8405,N_8803);
nor UO_355 (O_355,N_8438,N_8937);
nor UO_356 (O_356,N_8917,N_8717);
and UO_357 (O_357,N_8277,N_9769);
nor UO_358 (O_358,N_9307,N_9658);
and UO_359 (O_359,N_8467,N_8156);
and UO_360 (O_360,N_8533,N_8539);
nand UO_361 (O_361,N_8094,N_9125);
and UO_362 (O_362,N_9997,N_9258);
nor UO_363 (O_363,N_9467,N_9131);
nor UO_364 (O_364,N_8349,N_8103);
nand UO_365 (O_365,N_8397,N_9682);
and UO_366 (O_366,N_8582,N_9386);
nor UO_367 (O_367,N_9331,N_8619);
xor UO_368 (O_368,N_9772,N_9310);
and UO_369 (O_369,N_9084,N_8320);
nor UO_370 (O_370,N_9674,N_9841);
or UO_371 (O_371,N_8241,N_8835);
nand UO_372 (O_372,N_9052,N_9630);
and UO_373 (O_373,N_8661,N_9077);
or UO_374 (O_374,N_9756,N_9257);
nor UO_375 (O_375,N_9008,N_9359);
nand UO_376 (O_376,N_8050,N_9233);
nor UO_377 (O_377,N_8698,N_8407);
and UO_378 (O_378,N_8953,N_9024);
or UO_379 (O_379,N_8465,N_8189);
nor UO_380 (O_380,N_8689,N_8466);
and UO_381 (O_381,N_8176,N_9514);
nand UO_382 (O_382,N_9091,N_8823);
and UO_383 (O_383,N_8356,N_9045);
xnor UO_384 (O_384,N_9898,N_9428);
or UO_385 (O_385,N_9069,N_9815);
nand UO_386 (O_386,N_8043,N_9014);
nor UO_387 (O_387,N_9371,N_9471);
and UO_388 (O_388,N_9491,N_9197);
nor UO_389 (O_389,N_9365,N_8359);
and UO_390 (O_390,N_9529,N_9610);
nor UO_391 (O_391,N_9621,N_9988);
or UO_392 (O_392,N_8997,N_8303);
or UO_393 (O_393,N_8149,N_9633);
and UO_394 (O_394,N_8201,N_9939);
and UO_395 (O_395,N_9585,N_8010);
and UO_396 (O_396,N_8576,N_8610);
and UO_397 (O_397,N_8599,N_9562);
or UO_398 (O_398,N_8411,N_8016);
nor UO_399 (O_399,N_8879,N_9616);
and UO_400 (O_400,N_8558,N_8904);
or UO_401 (O_401,N_8119,N_9723);
nor UO_402 (O_402,N_9286,N_8788);
nor UO_403 (O_403,N_8044,N_9893);
or UO_404 (O_404,N_8822,N_9702);
and UO_405 (O_405,N_9915,N_8274);
and UO_406 (O_406,N_9249,N_9690);
nand UO_407 (O_407,N_8880,N_8796);
and UO_408 (O_408,N_8787,N_9517);
nand UO_409 (O_409,N_8651,N_8306);
nand UO_410 (O_410,N_8557,N_8151);
nand UO_411 (O_411,N_9679,N_8272);
nor UO_412 (O_412,N_8225,N_8666);
and UO_413 (O_413,N_8827,N_9094);
and UO_414 (O_414,N_9013,N_9210);
nand UO_415 (O_415,N_8170,N_9573);
nor UO_416 (O_416,N_9634,N_8999);
or UO_417 (O_417,N_8175,N_9440);
nor UO_418 (O_418,N_9867,N_8654);
nor UO_419 (O_419,N_8199,N_8660);
nand UO_420 (O_420,N_9165,N_8996);
nand UO_421 (O_421,N_9328,N_8624);
nand UO_422 (O_422,N_8110,N_9183);
and UO_423 (O_423,N_8290,N_9766);
nand UO_424 (O_424,N_9725,N_9109);
or UO_425 (O_425,N_9151,N_9017);
nand UO_426 (O_426,N_9085,N_8903);
nand UO_427 (O_427,N_9171,N_9422);
or UO_428 (O_428,N_9762,N_9200);
and UO_429 (O_429,N_9925,N_8896);
and UO_430 (O_430,N_9671,N_9236);
nand UO_431 (O_431,N_8198,N_9470);
and UO_432 (O_432,N_9545,N_9049);
nor UO_433 (O_433,N_9894,N_8378);
and UO_434 (O_434,N_8325,N_8542);
or UO_435 (O_435,N_8255,N_9865);
nor UO_436 (O_436,N_8350,N_9294);
and UO_437 (O_437,N_8645,N_8556);
nor UO_438 (O_438,N_8723,N_9020);
and UO_439 (O_439,N_8954,N_8200);
xnor UO_440 (O_440,N_8719,N_9047);
nand UO_441 (O_441,N_9012,N_8143);
nor UO_442 (O_442,N_9226,N_9955);
nor UO_443 (O_443,N_9763,N_8315);
nand UO_444 (O_444,N_8860,N_8750);
or UO_445 (O_445,N_9413,N_9647);
nor UO_446 (O_446,N_9710,N_9039);
and UO_447 (O_447,N_9708,N_9744);
and UO_448 (O_448,N_9199,N_9374);
and UO_449 (O_449,N_9357,N_9876);
nand UO_450 (O_450,N_8459,N_9480);
nor UO_451 (O_451,N_9408,N_8456);
nand UO_452 (O_452,N_8065,N_9902);
and UO_453 (O_453,N_8605,N_9507);
xor UO_454 (O_454,N_9935,N_8307);
xnor UO_455 (O_455,N_8863,N_8943);
xor UO_456 (O_456,N_8403,N_9141);
and UO_457 (O_457,N_9689,N_8702);
nand UO_458 (O_458,N_9801,N_8989);
and UO_459 (O_459,N_8641,N_9469);
nand UO_460 (O_460,N_9416,N_9315);
nand UO_461 (O_461,N_8983,N_9204);
and UO_462 (O_462,N_8782,N_8347);
nand UO_463 (O_463,N_8927,N_8844);
and UO_464 (O_464,N_9834,N_8491);
nor UO_465 (O_465,N_8229,N_8348);
nand UO_466 (O_466,N_8613,N_8994);
and UO_467 (O_467,N_8450,N_8424);
and UO_468 (O_468,N_9642,N_9299);
and UO_469 (O_469,N_8639,N_8008);
nor UO_470 (O_470,N_8283,N_8250);
and UO_471 (O_471,N_9010,N_9810);
and UO_472 (O_472,N_9811,N_8578);
or UO_473 (O_473,N_8638,N_9818);
nand UO_474 (O_474,N_8673,N_8445);
nand UO_475 (O_475,N_9574,N_9528);
nand UO_476 (O_476,N_8279,N_9945);
xor UO_477 (O_477,N_8507,N_9475);
nand UO_478 (O_478,N_8392,N_9267);
or UO_479 (O_479,N_9700,N_8483);
and UO_480 (O_480,N_8724,N_9018);
or UO_481 (O_481,N_9112,N_8907);
or UO_482 (O_482,N_9164,N_9672);
nor UO_483 (O_483,N_8847,N_9345);
nor UO_484 (O_484,N_8462,N_8727);
and UO_485 (O_485,N_8683,N_9033);
nand UO_486 (O_486,N_9129,N_9316);
nand UO_487 (O_487,N_8939,N_8735);
and UO_488 (O_488,N_9730,N_9814);
and UO_489 (O_489,N_8133,N_8530);
nor UO_490 (O_490,N_9673,N_9457);
and UO_491 (O_491,N_8553,N_9146);
nor UO_492 (O_492,N_8963,N_8413);
nand UO_493 (O_493,N_8504,N_8831);
nor UO_494 (O_494,N_8497,N_9436);
nor UO_495 (O_495,N_8379,N_8370);
or UO_496 (O_496,N_9259,N_9547);
nand UO_497 (O_497,N_9838,N_9875);
nor UO_498 (O_498,N_8453,N_8107);
or UO_499 (O_499,N_9948,N_8042);
nor UO_500 (O_500,N_8845,N_9058);
xor UO_501 (O_501,N_9731,N_9092);
nor UO_502 (O_502,N_8756,N_8377);
or UO_503 (O_503,N_8680,N_8090);
nand UO_504 (O_504,N_9726,N_8083);
and UO_505 (O_505,N_9897,N_9994);
or UO_506 (O_506,N_8209,N_9619);
nand UO_507 (O_507,N_9755,N_8389);
or UO_508 (O_508,N_9492,N_9273);
and UO_509 (O_509,N_9399,N_8020);
or UO_510 (O_510,N_8731,N_9102);
nor UO_511 (O_511,N_8073,N_9260);
or UO_512 (O_512,N_9445,N_9516);
or UO_513 (O_513,N_9269,N_8265);
or UO_514 (O_514,N_9712,N_8298);
and UO_515 (O_515,N_8884,N_9334);
nand UO_516 (O_516,N_8889,N_9264);
or UO_517 (O_517,N_8029,N_9504);
or UO_518 (O_518,N_9536,N_9276);
nor UO_519 (O_519,N_8760,N_9976);
nand UO_520 (O_520,N_9463,N_9877);
and UO_521 (O_521,N_9414,N_8235);
nand UO_522 (O_522,N_8153,N_8908);
nor UO_523 (O_523,N_8237,N_9944);
nand UO_524 (O_524,N_9886,N_8262);
and UO_525 (O_525,N_9558,N_8604);
and UO_526 (O_526,N_9038,N_9586);
and UO_527 (O_527,N_9830,N_8849);
and UO_528 (O_528,N_9780,N_9611);
and UO_529 (O_529,N_8650,N_9362);
or UO_530 (O_530,N_9011,N_8960);
and UO_531 (O_531,N_9160,N_8819);
and UO_532 (O_532,N_9485,N_9932);
nand UO_533 (O_533,N_8291,N_8282);
xnor UO_534 (O_534,N_8725,N_8481);
and UO_535 (O_535,N_8374,N_8418);
or UO_536 (O_536,N_8469,N_9950);
nor UO_537 (O_537,N_8473,N_8482);
and UO_538 (O_538,N_9908,N_9301);
nor UO_539 (O_539,N_8527,N_8534);
or UO_540 (O_540,N_9522,N_9176);
or UO_541 (O_541,N_8476,N_8251);
and UO_542 (O_542,N_8270,N_9032);
nor UO_543 (O_543,N_8328,N_9615);
nand UO_544 (O_544,N_8138,N_9478);
nand UO_545 (O_545,N_9161,N_8223);
nand UO_546 (O_546,N_9130,N_9159);
or UO_547 (O_547,N_9477,N_9390);
and UO_548 (O_548,N_9454,N_9891);
or UO_549 (O_549,N_9612,N_9282);
or UO_550 (O_550,N_9349,N_9793);
nor UO_551 (O_551,N_8289,N_8437);
and UO_552 (O_552,N_8957,N_8851);
nand UO_553 (O_553,N_9135,N_8959);
nand UO_554 (O_554,N_9859,N_8127);
and UO_555 (O_555,N_9594,N_9580);
or UO_556 (O_556,N_8310,N_9608);
or UO_557 (O_557,N_9387,N_8769);
nand UO_558 (O_558,N_8012,N_8738);
nor UO_559 (O_559,N_9853,N_8431);
or UO_560 (O_560,N_8154,N_8060);
or UO_561 (O_561,N_9957,N_8353);
nand UO_562 (O_562,N_9588,N_8025);
nor UO_563 (O_563,N_8062,N_8688);
nor UO_564 (O_564,N_9424,N_8070);
nand UO_565 (O_565,N_9396,N_9498);
and UO_566 (O_566,N_8502,N_9022);
or UO_567 (O_567,N_9552,N_9392);
nor UO_568 (O_568,N_9341,N_9617);
and UO_569 (O_569,N_8135,N_8118);
nor UO_570 (O_570,N_8341,N_8355);
and UO_571 (O_571,N_9016,N_9412);
nand UO_572 (O_572,N_8987,N_8991);
nand UO_573 (O_573,N_9777,N_8742);
nand UO_574 (O_574,N_9231,N_9088);
or UO_575 (O_575,N_9644,N_8935);
nor UO_576 (O_576,N_8911,N_9912);
and UO_577 (O_577,N_8224,N_8883);
nor UO_578 (O_578,N_8316,N_9549);
nor UO_579 (O_579,N_8388,N_8789);
or UO_580 (O_580,N_9251,N_8815);
and UO_581 (O_581,N_8732,N_8579);
or UO_582 (O_582,N_9265,N_9520);
or UO_583 (O_583,N_9985,N_8617);
nand UO_584 (O_584,N_9366,N_8524);
nor UO_585 (O_585,N_9207,N_9053);
and UO_586 (O_586,N_8093,N_9217);
nand UO_587 (O_587,N_9384,N_8240);
nand UO_588 (O_588,N_8053,N_9000);
or UO_589 (O_589,N_8113,N_9624);
nand UO_590 (O_590,N_9822,N_9373);
nand UO_591 (O_591,N_9347,N_8096);
and UO_592 (O_592,N_8027,N_9182);
or UO_593 (O_593,N_8701,N_9458);
and UO_594 (O_594,N_8629,N_8669);
nor UO_595 (O_595,N_9194,N_9031);
or UO_596 (O_596,N_8829,N_9641);
or UO_597 (O_597,N_9222,N_8675);
and UO_598 (O_598,N_8622,N_9605);
nor UO_599 (O_599,N_8951,N_8125);
nor UO_600 (O_600,N_8399,N_9006);
or UO_601 (O_601,N_8475,N_8535);
and UO_602 (O_602,N_9735,N_9879);
and UO_603 (O_603,N_9348,N_8964);
nand UO_604 (O_604,N_9940,N_8928);
nand UO_605 (O_605,N_8139,N_8914);
nand UO_606 (O_606,N_9472,N_8190);
nor UO_607 (O_607,N_8566,N_9765);
nor UO_608 (O_608,N_9474,N_9914);
and UO_609 (O_609,N_9266,N_9541);
or UO_610 (O_610,N_8519,N_9311);
nor UO_611 (O_611,N_8643,N_8858);
nand UO_612 (O_612,N_8792,N_8031);
nand UO_613 (O_613,N_8051,N_9202);
and UO_614 (O_614,N_9170,N_8565);
and UO_615 (O_615,N_8872,N_8901);
nand UO_616 (O_616,N_9821,N_9456);
nor UO_617 (O_617,N_8460,N_9509);
and UO_618 (O_618,N_8034,N_8704);
nand UO_619 (O_619,N_8681,N_9419);
nor UO_620 (O_620,N_8514,N_8888);
nand UO_621 (O_621,N_8117,N_8047);
and UO_622 (O_622,N_8982,N_9595);
and UO_623 (O_623,N_8129,N_9042);
and UO_624 (O_624,N_9637,N_9355);
and UO_625 (O_625,N_9820,N_8375);
nand UO_626 (O_626,N_9444,N_8394);
nor UO_627 (O_627,N_8893,N_9330);
nor UO_628 (O_628,N_8408,N_9943);
nand UO_629 (O_629,N_9697,N_8264);
nand UO_630 (O_630,N_8891,N_8976);
or UO_631 (O_631,N_8054,N_9878);
nor UO_632 (O_632,N_9224,N_9035);
and UO_633 (O_633,N_9284,N_8764);
nor UO_634 (O_634,N_9082,N_8513);
or UO_635 (O_635,N_8780,N_8572);
and UO_636 (O_636,N_8454,N_8287);
or UO_637 (O_637,N_9956,N_8532);
nand UO_638 (O_638,N_8003,N_9191);
and UO_639 (O_639,N_9309,N_8439);
nor UO_640 (O_640,N_8902,N_9919);
or UO_641 (O_641,N_8293,N_8228);
xor UO_642 (O_642,N_9168,N_8045);
or UO_643 (O_643,N_8080,N_8806);
nand UO_644 (O_644,N_9123,N_9563);
nor UO_645 (O_645,N_8711,N_8608);
or UO_646 (O_646,N_8569,N_8432);
and UO_647 (O_647,N_8798,N_9973);
xor UO_648 (O_648,N_9262,N_8737);
nor UO_649 (O_649,N_8485,N_9675);
and UO_650 (O_650,N_9752,N_9656);
nor UO_651 (O_651,N_9375,N_9687);
nor UO_652 (O_652,N_8772,N_8762);
nor UO_653 (O_653,N_8970,N_8441);
nor UO_654 (O_654,N_8451,N_8744);
or UO_655 (O_655,N_9188,N_9881);
nor UO_656 (O_656,N_9242,N_9890);
nand UO_657 (O_657,N_9021,N_8244);
or UO_658 (O_658,N_8471,N_8136);
nor UO_659 (O_659,N_8525,N_9136);
nand UO_660 (O_660,N_8647,N_8816);
or UO_661 (O_661,N_8178,N_9779);
xnor UO_662 (O_662,N_8721,N_8659);
or UO_663 (O_663,N_8121,N_8855);
and UO_664 (O_664,N_8755,N_9778);
or UO_665 (O_665,N_9336,N_8496);
nand UO_666 (O_666,N_8286,N_9462);
nand UO_667 (O_667,N_8231,N_8771);
nand UO_668 (O_668,N_9376,N_9073);
nor UO_669 (O_669,N_8501,N_8214);
nand UO_670 (O_670,N_9317,N_9312);
nor UO_671 (O_671,N_8770,N_8751);
nand UO_672 (O_672,N_8238,N_9628);
or UO_673 (O_673,N_9533,N_8794);
nand UO_674 (O_674,N_8208,N_9706);
or UO_675 (O_675,N_8621,N_8707);
nor UO_676 (O_676,N_8965,N_8585);
nor UO_677 (O_677,N_9959,N_8023);
or UO_678 (O_678,N_8243,N_9805);
nor UO_679 (O_679,N_9705,N_8226);
or UO_680 (O_680,N_9056,N_8157);
and UO_681 (O_681,N_9461,N_9759);
nor UO_682 (O_682,N_9340,N_8242);
nand UO_683 (O_683,N_8890,N_8918);
and UO_684 (O_684,N_9792,N_8092);
and UO_685 (O_685,N_8442,N_9156);
nand UO_686 (O_686,N_8644,N_8091);
nor UO_687 (O_687,N_8574,N_8101);
nor UO_688 (O_688,N_9565,N_9420);
nand UO_689 (O_689,N_9149,N_9421);
nand UO_690 (O_690,N_9115,N_9442);
or UO_691 (O_691,N_9289,N_8252);
nand UO_692 (O_692,N_9826,N_8104);
and UO_693 (O_693,N_8974,N_9864);
or UO_694 (O_694,N_9962,N_8882);
nand UO_695 (O_695,N_8182,N_9885);
nand UO_696 (O_696,N_8706,N_9843);
xor UO_697 (O_697,N_9828,N_9450);
or UO_698 (O_698,N_9768,N_8933);
or UO_699 (O_699,N_8383,N_8691);
or UO_700 (O_700,N_9967,N_8192);
nor UO_701 (O_701,N_8030,N_8217);
nand UO_702 (O_702,N_8380,N_8940);
and UO_703 (O_703,N_9926,N_8365);
nor UO_704 (O_704,N_9987,N_8028);
or UO_705 (O_705,N_8747,N_8230);
or UO_706 (O_706,N_9933,N_9484);
nor UO_707 (O_707,N_8988,N_9947);
and UO_708 (O_708,N_9813,N_8479);
nand UO_709 (O_709,N_8694,N_9589);
nand UO_710 (O_710,N_8817,N_9448);
and UO_711 (O_711,N_9339,N_8512);
or UO_712 (O_712,N_9804,N_8449);
or UO_713 (O_713,N_9677,N_8425);
nand UO_714 (O_714,N_9862,N_8150);
and UO_715 (O_715,N_9693,N_9145);
or UO_716 (O_716,N_9728,N_8767);
or UO_717 (O_717,N_9963,N_9098);
nor UO_718 (O_718,N_8202,N_8979);
or UO_719 (O_719,N_9575,N_8537);
nand UO_720 (O_720,N_8592,N_8913);
nor UO_721 (O_721,N_8634,N_8623);
nand UO_722 (O_722,N_8181,N_9372);
and UO_723 (O_723,N_9060,N_8958);
or UO_724 (O_724,N_8801,N_8864);
or UO_725 (O_725,N_9106,N_9213);
nor UO_726 (O_726,N_8329,N_9153);
and UO_727 (O_727,N_8718,N_8232);
or UO_728 (O_728,N_8749,N_9719);
nand UO_729 (O_729,N_9620,N_9007);
nand UO_730 (O_730,N_8587,N_8531);
nand UO_731 (O_731,N_8559,N_9513);
and UO_732 (O_732,N_8590,N_9306);
and UO_733 (O_733,N_8336,N_9540);
or UO_734 (O_734,N_9208,N_9727);
and UO_735 (O_735,N_9578,N_9747);
and UO_736 (O_736,N_9126,N_9851);
and UO_737 (O_737,N_9065,N_9670);
or UO_738 (O_738,N_8463,N_9592);
nand UO_739 (O_739,N_9405,N_8684);
and UO_740 (O_740,N_9270,N_9019);
and UO_741 (O_741,N_9953,N_9138);
nor UO_742 (O_742,N_9009,N_9577);
and UO_743 (O_743,N_8877,N_8387);
or UO_744 (O_744,N_9385,N_9318);
nor UO_745 (O_745,N_8886,N_9367);
and UO_746 (O_746,N_9525,N_8066);
or UO_747 (O_747,N_9938,N_9542);
nor UO_748 (O_748,N_8696,N_8024);
or UO_749 (O_749,N_9483,N_9166);
or UO_750 (O_750,N_8662,N_9846);
or UO_751 (O_751,N_9358,N_9668);
and UO_752 (O_752,N_8253,N_8503);
or UO_753 (O_753,N_9201,N_9256);
or UO_754 (O_754,N_8273,N_9989);
or UO_755 (O_755,N_8687,N_8122);
nand UO_756 (O_756,N_8626,N_9036);
nand UO_757 (O_757,N_9027,N_9239);
nand UO_758 (O_758,N_8161,N_9121);
nand UO_759 (O_759,N_9927,N_8052);
and UO_760 (O_760,N_8635,N_9063);
nor UO_761 (O_761,N_8922,N_9556);
and UO_762 (O_762,N_9954,N_8256);
nor UO_763 (O_763,N_8834,N_9054);
or UO_764 (O_764,N_9880,N_9584);
nor UO_765 (O_765,N_8422,N_9518);
nor UO_766 (O_766,N_9788,N_8071);
nand UO_767 (O_767,N_9949,N_8716);
and UO_768 (O_768,N_9539,N_8984);
or UO_769 (O_769,N_8600,N_8280);
nand UO_770 (O_770,N_8865,N_9911);
and UO_771 (O_771,N_8364,N_9829);
xor UO_772 (O_772,N_8695,N_9869);
nor UO_773 (O_773,N_9511,N_9274);
or UO_774 (O_774,N_9749,N_9784);
nand UO_775 (O_775,N_9951,N_8573);
nor UO_776 (O_776,N_9319,N_9503);
and UO_777 (O_777,N_8276,N_9764);
nand UO_778 (O_778,N_8627,N_8100);
nand UO_779 (O_779,N_9150,N_8446);
nand UO_780 (O_780,N_8404,N_8373);
and UO_781 (O_781,N_9305,N_8494);
or UO_782 (O_782,N_9887,N_8452);
or UO_783 (O_783,N_8734,N_9942);
nand UO_784 (O_784,N_8679,N_9225);
or UO_785 (O_785,N_9026,N_8840);
or UO_786 (O_786,N_8340,N_9337);
nand UO_787 (O_787,N_8763,N_9600);
and UO_788 (O_788,N_9737,N_9631);
and UO_789 (O_789,N_9394,N_9499);
or UO_790 (O_790,N_8085,N_8636);
or UO_791 (O_791,N_9025,N_8615);
nor UO_792 (O_792,N_9931,N_8658);
and UO_793 (O_793,N_9175,N_8036);
and UO_794 (O_794,N_8281,N_8637);
nor UO_795 (O_795,N_9833,N_8337);
or UO_796 (O_796,N_8297,N_8895);
and UO_797 (O_797,N_9389,N_9114);
and UO_798 (O_798,N_8642,N_9143);
and UO_799 (O_799,N_8308,N_9568);
and UO_800 (O_800,N_9521,N_8926);
xnor UO_801 (O_801,N_9379,N_9981);
nor UO_802 (O_802,N_9543,N_8381);
nor UO_803 (O_803,N_9819,N_9459);
and UO_804 (O_804,N_8197,N_9718);
nand UO_805 (O_805,N_9404,N_8108);
or UO_806 (O_806,N_9067,N_8838);
or UO_807 (O_807,N_8923,N_8759);
and UO_808 (O_808,N_8942,N_9774);
or UO_809 (O_809,N_8216,N_9250);
nor UO_810 (O_810,N_8141,N_8601);
or UO_811 (O_811,N_8975,N_9999);
and UO_812 (O_812,N_8881,N_9167);
and UO_813 (O_813,N_9041,N_8686);
or UO_814 (O_814,N_8218,N_8766);
and UO_815 (O_815,N_9144,N_8859);
nor UO_816 (O_816,N_9411,N_8268);
nor UO_817 (O_817,N_9795,N_8773);
or UO_818 (O_818,N_9924,N_8112);
nor UO_819 (O_819,N_8115,N_8614);
and UO_820 (O_820,N_9567,N_9352);
nand UO_821 (O_821,N_8852,N_9753);
and UO_822 (O_822,N_9904,N_8575);
nor UO_823 (O_823,N_8825,N_9496);
nand UO_824 (O_824,N_8271,N_8833);
nor UO_825 (O_825,N_8019,N_9427);
and UO_826 (O_826,N_9873,N_8814);
nor UO_827 (O_827,N_8331,N_8247);
nor UO_828 (O_828,N_9986,N_8211);
and UO_829 (O_829,N_9900,N_8488);
nor UO_830 (O_830,N_8972,N_9468);
nor UO_831 (O_831,N_8203,N_8086);
and UO_832 (O_832,N_8522,N_8968);
nor UO_833 (O_833,N_8529,N_8915);
and UO_834 (O_834,N_9179,N_8292);
nand UO_835 (O_835,N_9767,N_8317);
nor UO_836 (O_836,N_8540,N_9401);
and UO_837 (O_837,N_8102,N_8171);
nor UO_838 (O_838,N_9806,N_8857);
and UO_839 (O_839,N_8330,N_9288);
nand UO_840 (O_840,N_8064,N_9302);
nor UO_841 (O_841,N_9275,N_9850);
and UO_842 (O_842,N_8087,N_9720);
nor UO_843 (O_843,N_8351,N_8458);
and UO_844 (O_844,N_9400,N_9481);
and UO_845 (O_845,N_8549,N_9907);
nor UO_846 (O_846,N_8386,N_9866);
or UO_847 (O_847,N_8173,N_8416);
nor UO_848 (O_848,N_9685,N_9326);
and UO_849 (O_849,N_9648,N_9206);
or UO_850 (O_850,N_8114,N_9526);
nand UO_851 (O_851,N_9308,N_8155);
or UO_852 (O_852,N_8395,N_9734);
nand UO_853 (O_853,N_8878,N_8400);
nor UO_854 (O_854,N_9074,N_9844);
nand UO_855 (O_855,N_8372,N_8945);
nand UO_856 (O_856,N_9344,N_8257);
xor UO_857 (O_857,N_9117,N_9745);
nand UO_858 (O_858,N_8089,N_9655);
nor UO_859 (O_859,N_8015,N_9023);
nand UO_860 (O_860,N_8049,N_8005);
or UO_861 (O_861,N_9629,N_8002);
nand UO_862 (O_862,N_9283,N_9936);
and UO_863 (O_863,N_9423,N_9707);
nor UO_864 (O_864,N_9892,N_9502);
nor UO_865 (O_865,N_8910,N_8667);
nand UO_866 (O_866,N_9214,N_8430);
nand UO_867 (O_867,N_9464,N_8056);
or UO_868 (O_868,N_9971,N_8464);
nor UO_869 (O_869,N_8786,N_9603);
or UO_870 (O_870,N_8472,N_9132);
nor UO_871 (O_871,N_9789,N_9560);
nand UO_872 (O_872,N_8061,N_8258);
and UO_873 (O_873,N_9356,N_8898);
nand UO_874 (O_874,N_9593,N_8266);
or UO_875 (O_875,N_8948,N_9903);
or UO_876 (O_876,N_9969,N_8357);
nor UO_877 (O_877,N_9043,N_9099);
nand UO_878 (O_878,N_9232,N_8000);
or UO_879 (O_879,N_8648,N_8812);
and UO_880 (O_880,N_9455,N_9691);
nor UO_881 (O_881,N_8905,N_8390);
or UO_882 (O_882,N_9871,N_9196);
or UO_883 (O_883,N_9418,N_9120);
nor UO_884 (O_884,N_9081,N_8543);
or UO_885 (O_885,N_9555,N_9618);
and UO_886 (O_886,N_8607,N_8205);
nand UO_887 (O_887,N_9599,N_9193);
or UO_888 (O_888,N_8826,N_8088);
or UO_889 (O_889,N_9185,N_8142);
or UO_890 (O_890,N_8278,N_9550);
nor UO_891 (O_891,N_8486,N_8739);
or UO_892 (O_892,N_8343,N_8013);
or UO_893 (O_893,N_9652,N_8870);
nor UO_894 (O_894,N_8067,N_8444);
and UO_895 (O_895,N_8116,N_9937);
nand UO_896 (O_896,N_8366,N_9281);
or UO_897 (O_897,N_8628,N_8998);
and UO_898 (O_898,N_9452,N_9134);
and UO_899 (O_899,N_9254,N_8741);
xor UO_900 (O_900,N_8508,N_9093);
nor UO_901 (O_901,N_8126,N_8183);
nand UO_902 (O_902,N_8777,N_9388);
and UO_903 (O_903,N_9798,N_9546);
or UO_904 (O_904,N_8550,N_8186);
or UO_905 (O_905,N_8498,N_8790);
or UO_906 (O_906,N_8414,N_8632);
and UO_907 (O_907,N_8841,N_9736);
xnor UO_908 (O_908,N_9773,N_9473);
nand UO_909 (O_909,N_9061,N_9245);
nor UO_910 (O_910,N_9500,N_9350);
or UO_911 (O_911,N_9659,N_8213);
nor UO_912 (O_912,N_8932,N_9279);
nand UO_913 (O_913,N_9922,N_9506);
and UO_914 (O_914,N_9095,N_8260);
and UO_915 (O_915,N_9327,N_8026);
and UO_916 (O_916,N_8361,N_8204);
nor UO_917 (O_917,N_8220,N_9837);
nand UO_918 (O_918,N_8128,N_9453);
or UO_919 (O_919,N_9398,N_8040);
nand UO_920 (O_920,N_9155,N_8319);
nor UO_921 (O_921,N_9285,N_9606);
or UO_922 (O_922,N_8185,N_9057);
nand UO_923 (O_923,N_9823,N_9447);
nand UO_924 (O_924,N_9680,N_9177);
nand UO_925 (O_925,N_8081,N_9068);
and UO_926 (O_926,N_9581,N_9417);
nand UO_927 (O_927,N_8663,N_9695);
nand UO_928 (O_928,N_8166,N_9854);
and UO_929 (O_929,N_8547,N_9993);
and UO_930 (O_930,N_8249,N_8396);
and UO_931 (O_931,N_9380,N_8584);
xor UO_932 (O_932,N_8828,N_9694);
or UO_933 (O_933,N_8526,N_8753);
and UO_934 (O_934,N_8802,N_8312);
nand UO_935 (O_935,N_9990,N_8570);
and UO_936 (O_936,N_9783,N_9770);
nor UO_937 (O_937,N_9313,N_8854);
nor UO_938 (O_938,N_8006,N_9635);
nor UO_939 (O_939,N_9909,N_9799);
nor UO_940 (O_940,N_9703,N_8909);
and UO_941 (O_941,N_9051,N_8924);
or UO_942 (O_942,N_9622,N_9437);
nand UO_943 (O_943,N_9044,N_8234);
or UO_944 (O_944,N_8616,N_8916);
nand UO_945 (O_945,N_8690,N_8124);
or UO_946 (O_946,N_8367,N_8097);
nor UO_947 (O_947,N_9059,N_9005);
or UO_948 (O_948,N_8492,N_9431);
and UO_949 (O_949,N_8288,N_9847);
and UO_950 (O_950,N_8778,N_9571);
and UO_951 (O_951,N_9139,N_8995);
or UO_952 (O_952,N_8017,N_9300);
nand UO_953 (O_953,N_8106,N_8758);
nand UO_954 (O_954,N_9122,N_9983);
nor UO_955 (O_955,N_8625,N_9590);
and UO_956 (O_956,N_8076,N_8041);
or UO_957 (O_957,N_8443,N_8906);
and UO_958 (O_958,N_9696,N_9048);
or UO_959 (O_959,N_9729,N_9147);
or UO_960 (O_960,N_9393,N_8196);
nand UO_961 (O_961,N_9910,N_9030);
nor UO_962 (O_962,N_9802,N_8589);
or UO_963 (O_963,N_9247,N_9531);
nand UO_964 (O_964,N_8714,N_9003);
or UO_965 (O_965,N_8785,N_8720);
nor UO_966 (O_966,N_9709,N_9108);
or UO_967 (O_967,N_9598,N_9913);
or UO_968 (O_968,N_8500,N_9564);
or UO_969 (O_969,N_8853,N_8967);
nor UO_970 (O_970,N_8868,N_8713);
or UO_971 (O_971,N_8184,N_9626);
and UO_972 (O_972,N_8490,N_9816);
or UO_973 (O_973,N_8931,N_8671);
or UO_974 (O_974,N_9002,N_8682);
or UO_975 (O_975,N_9103,N_8382);
or UO_976 (O_976,N_8038,N_8478);
nand UO_977 (O_977,N_8314,N_9501);
xnor UO_978 (O_978,N_9443,N_9246);
nand UO_979 (O_979,N_9713,N_8172);
nor UO_980 (O_980,N_9669,N_8055);
and UO_981 (O_981,N_8077,N_8480);
or UO_982 (O_982,N_9451,N_8541);
or UO_983 (O_983,N_9701,N_9004);
and UO_984 (O_984,N_8925,N_8022);
nand UO_985 (O_985,N_8709,N_9721);
nor UO_986 (O_986,N_9505,N_8523);
nor UO_987 (O_987,N_9148,N_9569);
and UO_988 (O_988,N_8429,N_9842);
nor UO_989 (O_989,N_9487,N_8039);
or UO_990 (O_990,N_8194,N_9101);
and UO_991 (O_991,N_8544,N_8195);
nand UO_992 (O_992,N_9882,N_8754);
nand UO_993 (O_993,N_8419,N_9524);
nor UO_994 (O_994,N_8618,N_8362);
or UO_995 (O_995,N_9711,N_8148);
nand UO_996 (O_996,N_8710,N_9154);
nand UO_997 (O_997,N_8433,N_9323);
and UO_998 (O_998,N_9650,N_9946);
or UO_999 (O_999,N_9587,N_9921);
nand UO_1000 (O_1000,N_9711,N_8608);
and UO_1001 (O_1001,N_9345,N_9189);
or UO_1002 (O_1002,N_8166,N_9203);
nand UO_1003 (O_1003,N_9916,N_9454);
and UO_1004 (O_1004,N_8250,N_8886);
nand UO_1005 (O_1005,N_8197,N_8403);
nand UO_1006 (O_1006,N_9643,N_9025);
nand UO_1007 (O_1007,N_9659,N_9545);
and UO_1008 (O_1008,N_8050,N_9294);
nand UO_1009 (O_1009,N_9762,N_8469);
and UO_1010 (O_1010,N_9429,N_8917);
nand UO_1011 (O_1011,N_8044,N_8913);
or UO_1012 (O_1012,N_8571,N_8777);
or UO_1013 (O_1013,N_9638,N_9158);
or UO_1014 (O_1014,N_8168,N_8259);
nor UO_1015 (O_1015,N_8504,N_8926);
nand UO_1016 (O_1016,N_8536,N_8293);
nor UO_1017 (O_1017,N_9549,N_9947);
nor UO_1018 (O_1018,N_9740,N_8036);
xor UO_1019 (O_1019,N_8937,N_9016);
and UO_1020 (O_1020,N_9015,N_8133);
or UO_1021 (O_1021,N_8629,N_8073);
or UO_1022 (O_1022,N_8911,N_8811);
or UO_1023 (O_1023,N_9355,N_9106);
nand UO_1024 (O_1024,N_9997,N_9486);
nand UO_1025 (O_1025,N_8819,N_8872);
and UO_1026 (O_1026,N_8382,N_9016);
and UO_1027 (O_1027,N_8659,N_9522);
and UO_1028 (O_1028,N_8412,N_8532);
or UO_1029 (O_1029,N_8132,N_9297);
nor UO_1030 (O_1030,N_9402,N_8683);
nor UO_1031 (O_1031,N_8199,N_9929);
nand UO_1032 (O_1032,N_9618,N_9643);
nor UO_1033 (O_1033,N_8567,N_8872);
nor UO_1034 (O_1034,N_9288,N_8531);
nand UO_1035 (O_1035,N_8872,N_9434);
nor UO_1036 (O_1036,N_9344,N_9603);
and UO_1037 (O_1037,N_9535,N_9547);
nor UO_1038 (O_1038,N_8072,N_8417);
or UO_1039 (O_1039,N_8760,N_8826);
nor UO_1040 (O_1040,N_9847,N_8654);
nor UO_1041 (O_1041,N_8981,N_8955);
and UO_1042 (O_1042,N_8826,N_8774);
xnor UO_1043 (O_1043,N_8936,N_9906);
or UO_1044 (O_1044,N_9934,N_9285);
nor UO_1045 (O_1045,N_9717,N_9380);
or UO_1046 (O_1046,N_9081,N_9288);
nand UO_1047 (O_1047,N_8889,N_9841);
nor UO_1048 (O_1048,N_9302,N_9044);
xnor UO_1049 (O_1049,N_8883,N_9751);
or UO_1050 (O_1050,N_9352,N_8413);
nor UO_1051 (O_1051,N_8026,N_8912);
or UO_1052 (O_1052,N_8622,N_9971);
nor UO_1053 (O_1053,N_9582,N_9949);
xor UO_1054 (O_1054,N_8790,N_9849);
nand UO_1055 (O_1055,N_9032,N_9091);
nor UO_1056 (O_1056,N_9195,N_9372);
or UO_1057 (O_1057,N_9652,N_9455);
or UO_1058 (O_1058,N_8249,N_8007);
nor UO_1059 (O_1059,N_8009,N_9284);
nand UO_1060 (O_1060,N_8375,N_9895);
nand UO_1061 (O_1061,N_8613,N_8974);
or UO_1062 (O_1062,N_8511,N_8627);
nand UO_1063 (O_1063,N_8651,N_8386);
nor UO_1064 (O_1064,N_8949,N_9541);
or UO_1065 (O_1065,N_9227,N_9601);
xnor UO_1066 (O_1066,N_9489,N_9515);
nand UO_1067 (O_1067,N_8664,N_8146);
and UO_1068 (O_1068,N_9930,N_8590);
nand UO_1069 (O_1069,N_8652,N_8693);
nand UO_1070 (O_1070,N_8964,N_9259);
and UO_1071 (O_1071,N_9786,N_8010);
or UO_1072 (O_1072,N_8701,N_8171);
nand UO_1073 (O_1073,N_9539,N_8452);
nand UO_1074 (O_1074,N_9418,N_9619);
nor UO_1075 (O_1075,N_9277,N_8425);
or UO_1076 (O_1076,N_9880,N_8582);
and UO_1077 (O_1077,N_8605,N_8766);
nand UO_1078 (O_1078,N_8095,N_9255);
or UO_1079 (O_1079,N_9354,N_8591);
or UO_1080 (O_1080,N_9687,N_9207);
or UO_1081 (O_1081,N_9135,N_8463);
and UO_1082 (O_1082,N_9762,N_9229);
nor UO_1083 (O_1083,N_8290,N_9768);
nand UO_1084 (O_1084,N_8125,N_9660);
nor UO_1085 (O_1085,N_9692,N_8806);
nand UO_1086 (O_1086,N_9153,N_8378);
or UO_1087 (O_1087,N_9287,N_8426);
and UO_1088 (O_1088,N_9742,N_8928);
or UO_1089 (O_1089,N_8832,N_8653);
nor UO_1090 (O_1090,N_8180,N_9463);
and UO_1091 (O_1091,N_9412,N_9336);
and UO_1092 (O_1092,N_8120,N_8730);
nand UO_1093 (O_1093,N_8711,N_8920);
nand UO_1094 (O_1094,N_8562,N_8221);
and UO_1095 (O_1095,N_9616,N_8904);
nand UO_1096 (O_1096,N_8795,N_9302);
and UO_1097 (O_1097,N_9997,N_8620);
nor UO_1098 (O_1098,N_8908,N_8150);
nor UO_1099 (O_1099,N_9460,N_9277);
nand UO_1100 (O_1100,N_8621,N_9557);
nor UO_1101 (O_1101,N_8157,N_9666);
or UO_1102 (O_1102,N_8332,N_8726);
nand UO_1103 (O_1103,N_9245,N_8040);
xnor UO_1104 (O_1104,N_9324,N_9665);
nor UO_1105 (O_1105,N_9099,N_9213);
nor UO_1106 (O_1106,N_9082,N_9064);
or UO_1107 (O_1107,N_9757,N_9238);
or UO_1108 (O_1108,N_9724,N_9756);
nor UO_1109 (O_1109,N_8118,N_8101);
or UO_1110 (O_1110,N_8431,N_8650);
or UO_1111 (O_1111,N_9300,N_9534);
nor UO_1112 (O_1112,N_8206,N_8269);
or UO_1113 (O_1113,N_9048,N_9368);
nor UO_1114 (O_1114,N_8642,N_9911);
or UO_1115 (O_1115,N_8120,N_9039);
nor UO_1116 (O_1116,N_9079,N_8763);
nand UO_1117 (O_1117,N_8069,N_8852);
nand UO_1118 (O_1118,N_8878,N_9381);
nor UO_1119 (O_1119,N_8455,N_8609);
nand UO_1120 (O_1120,N_9583,N_9172);
nor UO_1121 (O_1121,N_8110,N_8759);
nand UO_1122 (O_1122,N_9274,N_9921);
nand UO_1123 (O_1123,N_9424,N_9661);
nand UO_1124 (O_1124,N_8537,N_9058);
and UO_1125 (O_1125,N_8400,N_8243);
xnor UO_1126 (O_1126,N_8043,N_9652);
or UO_1127 (O_1127,N_9753,N_8962);
nand UO_1128 (O_1128,N_9709,N_9258);
nand UO_1129 (O_1129,N_8250,N_8285);
and UO_1130 (O_1130,N_8651,N_8968);
nor UO_1131 (O_1131,N_8279,N_8074);
or UO_1132 (O_1132,N_8083,N_8097);
nor UO_1133 (O_1133,N_9035,N_9667);
and UO_1134 (O_1134,N_8428,N_9342);
or UO_1135 (O_1135,N_8862,N_8106);
nor UO_1136 (O_1136,N_8512,N_8233);
or UO_1137 (O_1137,N_8630,N_9889);
and UO_1138 (O_1138,N_8900,N_9125);
nor UO_1139 (O_1139,N_8687,N_8918);
nand UO_1140 (O_1140,N_9183,N_9560);
and UO_1141 (O_1141,N_9310,N_9546);
nor UO_1142 (O_1142,N_9635,N_8226);
or UO_1143 (O_1143,N_9183,N_9672);
nor UO_1144 (O_1144,N_9877,N_9745);
and UO_1145 (O_1145,N_9123,N_8723);
nor UO_1146 (O_1146,N_8461,N_8179);
or UO_1147 (O_1147,N_8241,N_8283);
or UO_1148 (O_1148,N_9576,N_9979);
nand UO_1149 (O_1149,N_8006,N_8407);
or UO_1150 (O_1150,N_8005,N_9847);
and UO_1151 (O_1151,N_8565,N_8722);
nor UO_1152 (O_1152,N_9914,N_8481);
or UO_1153 (O_1153,N_9732,N_9583);
nor UO_1154 (O_1154,N_9236,N_9557);
nor UO_1155 (O_1155,N_8996,N_9392);
and UO_1156 (O_1156,N_8614,N_9034);
nor UO_1157 (O_1157,N_9272,N_8041);
nand UO_1158 (O_1158,N_9487,N_8936);
or UO_1159 (O_1159,N_8297,N_8899);
nand UO_1160 (O_1160,N_8423,N_9700);
nand UO_1161 (O_1161,N_9897,N_9162);
or UO_1162 (O_1162,N_8381,N_8741);
nand UO_1163 (O_1163,N_8548,N_8614);
xnor UO_1164 (O_1164,N_8647,N_9468);
and UO_1165 (O_1165,N_9165,N_8660);
nand UO_1166 (O_1166,N_9875,N_8394);
nor UO_1167 (O_1167,N_8631,N_9264);
nand UO_1168 (O_1168,N_8558,N_8204);
or UO_1169 (O_1169,N_9859,N_8601);
nor UO_1170 (O_1170,N_9389,N_9124);
nor UO_1171 (O_1171,N_9968,N_8772);
or UO_1172 (O_1172,N_9983,N_8399);
nand UO_1173 (O_1173,N_8139,N_9001);
or UO_1174 (O_1174,N_8401,N_9473);
nor UO_1175 (O_1175,N_9236,N_9874);
nand UO_1176 (O_1176,N_8572,N_9679);
or UO_1177 (O_1177,N_9650,N_9274);
nor UO_1178 (O_1178,N_8014,N_9149);
nand UO_1179 (O_1179,N_8984,N_9834);
nand UO_1180 (O_1180,N_8157,N_8749);
and UO_1181 (O_1181,N_9094,N_9087);
xnor UO_1182 (O_1182,N_8600,N_9954);
nor UO_1183 (O_1183,N_8609,N_8138);
nand UO_1184 (O_1184,N_9201,N_8447);
nor UO_1185 (O_1185,N_9569,N_8516);
nor UO_1186 (O_1186,N_9700,N_8269);
nand UO_1187 (O_1187,N_8397,N_9398);
xor UO_1188 (O_1188,N_8650,N_9811);
and UO_1189 (O_1189,N_9583,N_8149);
or UO_1190 (O_1190,N_8819,N_9672);
nor UO_1191 (O_1191,N_8114,N_9792);
and UO_1192 (O_1192,N_8450,N_9336);
nand UO_1193 (O_1193,N_9931,N_8555);
or UO_1194 (O_1194,N_8292,N_8636);
nand UO_1195 (O_1195,N_8202,N_9560);
nor UO_1196 (O_1196,N_8002,N_9836);
nor UO_1197 (O_1197,N_8424,N_8584);
nor UO_1198 (O_1198,N_8045,N_8914);
or UO_1199 (O_1199,N_8910,N_8102);
and UO_1200 (O_1200,N_9738,N_9952);
and UO_1201 (O_1201,N_8491,N_9262);
or UO_1202 (O_1202,N_9426,N_8362);
or UO_1203 (O_1203,N_8266,N_9517);
nand UO_1204 (O_1204,N_9604,N_8001);
or UO_1205 (O_1205,N_8534,N_9613);
nor UO_1206 (O_1206,N_8244,N_8663);
nand UO_1207 (O_1207,N_9868,N_8289);
or UO_1208 (O_1208,N_8711,N_9873);
nand UO_1209 (O_1209,N_9390,N_8489);
nor UO_1210 (O_1210,N_8807,N_8716);
nor UO_1211 (O_1211,N_8596,N_8458);
or UO_1212 (O_1212,N_9954,N_8194);
and UO_1213 (O_1213,N_8041,N_9706);
and UO_1214 (O_1214,N_8088,N_8791);
nor UO_1215 (O_1215,N_8392,N_8433);
nand UO_1216 (O_1216,N_9007,N_9539);
or UO_1217 (O_1217,N_8487,N_8358);
nor UO_1218 (O_1218,N_9921,N_8836);
and UO_1219 (O_1219,N_9825,N_9064);
nand UO_1220 (O_1220,N_8505,N_8723);
and UO_1221 (O_1221,N_8053,N_9130);
and UO_1222 (O_1222,N_8485,N_8674);
nor UO_1223 (O_1223,N_8905,N_9809);
and UO_1224 (O_1224,N_9740,N_8958);
nand UO_1225 (O_1225,N_9376,N_8955);
or UO_1226 (O_1226,N_8360,N_8872);
or UO_1227 (O_1227,N_8497,N_8542);
xnor UO_1228 (O_1228,N_8417,N_9937);
nand UO_1229 (O_1229,N_9617,N_9356);
nor UO_1230 (O_1230,N_9107,N_8672);
and UO_1231 (O_1231,N_9508,N_8100);
or UO_1232 (O_1232,N_9726,N_9111);
or UO_1233 (O_1233,N_9011,N_8202);
or UO_1234 (O_1234,N_8397,N_8834);
or UO_1235 (O_1235,N_9088,N_8473);
or UO_1236 (O_1236,N_8930,N_8226);
or UO_1237 (O_1237,N_9616,N_9724);
nor UO_1238 (O_1238,N_8312,N_9548);
and UO_1239 (O_1239,N_8673,N_8117);
or UO_1240 (O_1240,N_9869,N_9457);
nor UO_1241 (O_1241,N_9886,N_8528);
or UO_1242 (O_1242,N_8350,N_8301);
nor UO_1243 (O_1243,N_9974,N_8638);
and UO_1244 (O_1244,N_9910,N_9456);
or UO_1245 (O_1245,N_9017,N_9899);
and UO_1246 (O_1246,N_9024,N_9023);
or UO_1247 (O_1247,N_8226,N_9986);
or UO_1248 (O_1248,N_8050,N_9303);
nor UO_1249 (O_1249,N_8594,N_9986);
or UO_1250 (O_1250,N_9131,N_9779);
and UO_1251 (O_1251,N_8403,N_8990);
nand UO_1252 (O_1252,N_8293,N_8742);
nor UO_1253 (O_1253,N_9007,N_9466);
nor UO_1254 (O_1254,N_9853,N_8159);
and UO_1255 (O_1255,N_8935,N_8738);
nand UO_1256 (O_1256,N_9489,N_8531);
nand UO_1257 (O_1257,N_9967,N_9366);
or UO_1258 (O_1258,N_8683,N_8654);
nand UO_1259 (O_1259,N_8882,N_9696);
nor UO_1260 (O_1260,N_9058,N_9662);
and UO_1261 (O_1261,N_9939,N_8631);
and UO_1262 (O_1262,N_8940,N_9131);
nand UO_1263 (O_1263,N_8573,N_9455);
and UO_1264 (O_1264,N_9109,N_9240);
or UO_1265 (O_1265,N_9042,N_8463);
nand UO_1266 (O_1266,N_8938,N_9508);
or UO_1267 (O_1267,N_8615,N_8357);
nand UO_1268 (O_1268,N_8279,N_9717);
or UO_1269 (O_1269,N_8969,N_9926);
nand UO_1270 (O_1270,N_8656,N_8445);
and UO_1271 (O_1271,N_8203,N_8637);
and UO_1272 (O_1272,N_9874,N_8919);
and UO_1273 (O_1273,N_9428,N_9100);
or UO_1274 (O_1274,N_8903,N_8500);
nand UO_1275 (O_1275,N_8983,N_9600);
nor UO_1276 (O_1276,N_9930,N_9871);
and UO_1277 (O_1277,N_8661,N_8871);
nand UO_1278 (O_1278,N_9576,N_9567);
nor UO_1279 (O_1279,N_8810,N_8852);
nand UO_1280 (O_1280,N_8367,N_9930);
nor UO_1281 (O_1281,N_8237,N_9988);
nor UO_1282 (O_1282,N_9386,N_9103);
or UO_1283 (O_1283,N_8374,N_9772);
and UO_1284 (O_1284,N_8270,N_8306);
nand UO_1285 (O_1285,N_9653,N_8764);
nand UO_1286 (O_1286,N_9308,N_9167);
and UO_1287 (O_1287,N_8036,N_8194);
and UO_1288 (O_1288,N_9169,N_8228);
and UO_1289 (O_1289,N_9473,N_8510);
nand UO_1290 (O_1290,N_8168,N_9070);
xor UO_1291 (O_1291,N_9866,N_9848);
nor UO_1292 (O_1292,N_9297,N_9556);
and UO_1293 (O_1293,N_9883,N_8618);
or UO_1294 (O_1294,N_9118,N_9067);
and UO_1295 (O_1295,N_9640,N_8150);
xnor UO_1296 (O_1296,N_9660,N_9772);
or UO_1297 (O_1297,N_8355,N_9209);
nand UO_1298 (O_1298,N_9881,N_9000);
nand UO_1299 (O_1299,N_9563,N_8300);
nor UO_1300 (O_1300,N_9339,N_9035);
nor UO_1301 (O_1301,N_8418,N_9472);
nor UO_1302 (O_1302,N_8510,N_8585);
or UO_1303 (O_1303,N_9115,N_9253);
nor UO_1304 (O_1304,N_9967,N_8830);
or UO_1305 (O_1305,N_9706,N_9278);
or UO_1306 (O_1306,N_9093,N_9149);
and UO_1307 (O_1307,N_9923,N_9391);
nor UO_1308 (O_1308,N_8410,N_8049);
and UO_1309 (O_1309,N_8395,N_9068);
nor UO_1310 (O_1310,N_9215,N_9717);
nand UO_1311 (O_1311,N_9725,N_9016);
nor UO_1312 (O_1312,N_9711,N_9168);
or UO_1313 (O_1313,N_9843,N_9861);
or UO_1314 (O_1314,N_9362,N_9198);
or UO_1315 (O_1315,N_8331,N_8745);
nand UO_1316 (O_1316,N_8340,N_8319);
nor UO_1317 (O_1317,N_8915,N_8299);
nor UO_1318 (O_1318,N_8922,N_8971);
and UO_1319 (O_1319,N_8809,N_8512);
or UO_1320 (O_1320,N_9753,N_8396);
nor UO_1321 (O_1321,N_9019,N_9268);
nand UO_1322 (O_1322,N_8851,N_8358);
and UO_1323 (O_1323,N_8570,N_8052);
or UO_1324 (O_1324,N_9532,N_9159);
nor UO_1325 (O_1325,N_9102,N_9772);
nand UO_1326 (O_1326,N_9536,N_8194);
nor UO_1327 (O_1327,N_8900,N_9463);
and UO_1328 (O_1328,N_9637,N_9318);
xnor UO_1329 (O_1329,N_9000,N_9284);
or UO_1330 (O_1330,N_8287,N_9232);
or UO_1331 (O_1331,N_9361,N_9730);
nand UO_1332 (O_1332,N_9946,N_8633);
and UO_1333 (O_1333,N_9911,N_9953);
or UO_1334 (O_1334,N_9585,N_8832);
and UO_1335 (O_1335,N_9792,N_8013);
or UO_1336 (O_1336,N_9251,N_8631);
and UO_1337 (O_1337,N_9767,N_9802);
nor UO_1338 (O_1338,N_8499,N_8559);
and UO_1339 (O_1339,N_9135,N_9066);
nand UO_1340 (O_1340,N_8969,N_8401);
xor UO_1341 (O_1341,N_8637,N_8399);
or UO_1342 (O_1342,N_8058,N_8324);
nor UO_1343 (O_1343,N_9063,N_9032);
and UO_1344 (O_1344,N_8689,N_8923);
and UO_1345 (O_1345,N_8741,N_9040);
or UO_1346 (O_1346,N_9491,N_9229);
or UO_1347 (O_1347,N_9619,N_8168);
and UO_1348 (O_1348,N_8901,N_8489);
nand UO_1349 (O_1349,N_9693,N_9953);
nor UO_1350 (O_1350,N_9497,N_9245);
nor UO_1351 (O_1351,N_9160,N_8570);
nand UO_1352 (O_1352,N_8373,N_9565);
nor UO_1353 (O_1353,N_8044,N_9344);
nor UO_1354 (O_1354,N_9436,N_8766);
or UO_1355 (O_1355,N_9124,N_8959);
or UO_1356 (O_1356,N_9361,N_8327);
and UO_1357 (O_1357,N_8182,N_8283);
nand UO_1358 (O_1358,N_8633,N_8130);
nand UO_1359 (O_1359,N_9978,N_8200);
and UO_1360 (O_1360,N_9148,N_9606);
and UO_1361 (O_1361,N_8929,N_9699);
nand UO_1362 (O_1362,N_9354,N_8102);
and UO_1363 (O_1363,N_9463,N_8583);
or UO_1364 (O_1364,N_8238,N_8007);
and UO_1365 (O_1365,N_8228,N_9741);
nor UO_1366 (O_1366,N_8474,N_8632);
or UO_1367 (O_1367,N_9863,N_8041);
and UO_1368 (O_1368,N_8343,N_8317);
xor UO_1369 (O_1369,N_9902,N_8554);
and UO_1370 (O_1370,N_9613,N_9926);
or UO_1371 (O_1371,N_8074,N_8112);
and UO_1372 (O_1372,N_9068,N_8355);
and UO_1373 (O_1373,N_8554,N_8409);
nor UO_1374 (O_1374,N_8493,N_8222);
nor UO_1375 (O_1375,N_9570,N_8066);
and UO_1376 (O_1376,N_8804,N_8851);
and UO_1377 (O_1377,N_9967,N_8360);
or UO_1378 (O_1378,N_9867,N_9740);
nand UO_1379 (O_1379,N_8838,N_8880);
nor UO_1380 (O_1380,N_8825,N_9609);
xnor UO_1381 (O_1381,N_8320,N_9351);
nor UO_1382 (O_1382,N_9631,N_9769);
or UO_1383 (O_1383,N_9868,N_9837);
or UO_1384 (O_1384,N_9006,N_8744);
nand UO_1385 (O_1385,N_8518,N_8384);
and UO_1386 (O_1386,N_8684,N_9730);
nor UO_1387 (O_1387,N_8908,N_8592);
or UO_1388 (O_1388,N_8339,N_9088);
xnor UO_1389 (O_1389,N_8118,N_8300);
and UO_1390 (O_1390,N_8715,N_8778);
or UO_1391 (O_1391,N_8214,N_9446);
nand UO_1392 (O_1392,N_9605,N_8023);
nor UO_1393 (O_1393,N_8908,N_9481);
or UO_1394 (O_1394,N_9385,N_8037);
nand UO_1395 (O_1395,N_9573,N_9493);
nand UO_1396 (O_1396,N_9548,N_8634);
and UO_1397 (O_1397,N_9638,N_8078);
nor UO_1398 (O_1398,N_8396,N_9538);
nand UO_1399 (O_1399,N_9722,N_9183);
nand UO_1400 (O_1400,N_8663,N_8838);
or UO_1401 (O_1401,N_9851,N_8076);
and UO_1402 (O_1402,N_9694,N_9987);
or UO_1403 (O_1403,N_8441,N_9935);
or UO_1404 (O_1404,N_9095,N_9448);
nand UO_1405 (O_1405,N_8034,N_9751);
and UO_1406 (O_1406,N_9091,N_8740);
nor UO_1407 (O_1407,N_8113,N_9389);
nand UO_1408 (O_1408,N_8316,N_9561);
nor UO_1409 (O_1409,N_8829,N_8324);
and UO_1410 (O_1410,N_8847,N_9787);
nand UO_1411 (O_1411,N_9259,N_9356);
nand UO_1412 (O_1412,N_8180,N_9218);
nand UO_1413 (O_1413,N_9152,N_8378);
nand UO_1414 (O_1414,N_8474,N_9675);
and UO_1415 (O_1415,N_8519,N_9966);
and UO_1416 (O_1416,N_9093,N_9770);
and UO_1417 (O_1417,N_8647,N_9476);
nor UO_1418 (O_1418,N_8905,N_8600);
nor UO_1419 (O_1419,N_8603,N_9654);
or UO_1420 (O_1420,N_9971,N_9489);
or UO_1421 (O_1421,N_9653,N_8162);
nand UO_1422 (O_1422,N_9285,N_9973);
or UO_1423 (O_1423,N_8046,N_9820);
nor UO_1424 (O_1424,N_8814,N_8290);
nand UO_1425 (O_1425,N_8899,N_8541);
nor UO_1426 (O_1426,N_8921,N_9780);
nor UO_1427 (O_1427,N_8654,N_8164);
nand UO_1428 (O_1428,N_8104,N_9393);
and UO_1429 (O_1429,N_9102,N_8633);
or UO_1430 (O_1430,N_8260,N_9292);
and UO_1431 (O_1431,N_8253,N_8968);
nor UO_1432 (O_1432,N_9183,N_9505);
or UO_1433 (O_1433,N_8632,N_9720);
or UO_1434 (O_1434,N_8605,N_9436);
and UO_1435 (O_1435,N_8335,N_9034);
or UO_1436 (O_1436,N_8068,N_9862);
xor UO_1437 (O_1437,N_9222,N_9935);
or UO_1438 (O_1438,N_8125,N_9256);
and UO_1439 (O_1439,N_8136,N_8806);
and UO_1440 (O_1440,N_9147,N_9684);
nor UO_1441 (O_1441,N_9660,N_9825);
or UO_1442 (O_1442,N_9646,N_9426);
nor UO_1443 (O_1443,N_9252,N_9021);
nor UO_1444 (O_1444,N_8117,N_9246);
nand UO_1445 (O_1445,N_9394,N_8099);
nand UO_1446 (O_1446,N_9352,N_8234);
or UO_1447 (O_1447,N_8801,N_9844);
or UO_1448 (O_1448,N_8771,N_8934);
nor UO_1449 (O_1449,N_9146,N_8607);
and UO_1450 (O_1450,N_9629,N_8951);
nor UO_1451 (O_1451,N_8461,N_8253);
and UO_1452 (O_1452,N_9197,N_8585);
and UO_1453 (O_1453,N_9106,N_9021);
or UO_1454 (O_1454,N_8385,N_8807);
or UO_1455 (O_1455,N_9689,N_9435);
nand UO_1456 (O_1456,N_8551,N_8288);
and UO_1457 (O_1457,N_8732,N_9634);
nand UO_1458 (O_1458,N_8418,N_9459);
nand UO_1459 (O_1459,N_9196,N_8663);
and UO_1460 (O_1460,N_9498,N_8987);
or UO_1461 (O_1461,N_9514,N_8589);
nand UO_1462 (O_1462,N_8715,N_8038);
nand UO_1463 (O_1463,N_9979,N_9431);
or UO_1464 (O_1464,N_9060,N_8968);
and UO_1465 (O_1465,N_8773,N_9424);
or UO_1466 (O_1466,N_9680,N_9141);
nand UO_1467 (O_1467,N_9622,N_9579);
and UO_1468 (O_1468,N_8074,N_9032);
or UO_1469 (O_1469,N_8309,N_8529);
and UO_1470 (O_1470,N_9361,N_9311);
or UO_1471 (O_1471,N_9318,N_8437);
nand UO_1472 (O_1472,N_8584,N_8219);
and UO_1473 (O_1473,N_9860,N_9171);
nor UO_1474 (O_1474,N_8931,N_9644);
xor UO_1475 (O_1475,N_8040,N_9450);
and UO_1476 (O_1476,N_8253,N_8025);
or UO_1477 (O_1477,N_9771,N_8230);
nor UO_1478 (O_1478,N_8447,N_8983);
and UO_1479 (O_1479,N_8324,N_9892);
or UO_1480 (O_1480,N_8881,N_9283);
or UO_1481 (O_1481,N_8654,N_8160);
nand UO_1482 (O_1482,N_9049,N_8623);
nand UO_1483 (O_1483,N_9492,N_8024);
xor UO_1484 (O_1484,N_8582,N_8358);
or UO_1485 (O_1485,N_9465,N_8572);
or UO_1486 (O_1486,N_9234,N_8715);
nand UO_1487 (O_1487,N_8483,N_9015);
nor UO_1488 (O_1488,N_9474,N_9602);
and UO_1489 (O_1489,N_9512,N_9198);
or UO_1490 (O_1490,N_9115,N_9459);
or UO_1491 (O_1491,N_9908,N_9362);
and UO_1492 (O_1492,N_8131,N_8063);
and UO_1493 (O_1493,N_8990,N_8338);
nand UO_1494 (O_1494,N_8254,N_9307);
and UO_1495 (O_1495,N_9732,N_8007);
and UO_1496 (O_1496,N_9434,N_8237);
and UO_1497 (O_1497,N_9162,N_8096);
xnor UO_1498 (O_1498,N_8785,N_9856);
nand UO_1499 (O_1499,N_9933,N_9818);
endmodule