module basic_500_3000_500_15_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_281,In_462);
or U1 (N_1,In_231,In_271);
nand U2 (N_2,In_471,In_356);
or U3 (N_3,In_273,In_106);
xor U4 (N_4,In_151,In_67);
nor U5 (N_5,In_393,In_154);
and U6 (N_6,In_195,In_191);
or U7 (N_7,In_40,In_410);
xnor U8 (N_8,In_58,In_98);
nand U9 (N_9,In_325,In_310);
or U10 (N_10,In_433,In_158);
or U11 (N_11,In_201,In_181);
or U12 (N_12,In_254,In_62);
and U13 (N_13,In_155,In_172);
or U14 (N_14,In_402,In_129);
and U15 (N_15,In_403,In_488);
nand U16 (N_16,In_329,In_25);
nand U17 (N_17,In_17,In_441);
and U18 (N_18,In_100,In_318);
or U19 (N_19,In_194,In_282);
nor U20 (N_20,In_364,In_35);
and U21 (N_21,In_414,In_82);
and U22 (N_22,In_304,In_164);
and U23 (N_23,In_37,In_114);
and U24 (N_24,In_493,In_406);
xnor U25 (N_25,In_293,In_352);
nand U26 (N_26,In_361,In_419);
and U27 (N_27,In_336,In_322);
nand U28 (N_28,In_59,In_122);
or U29 (N_29,In_171,In_245);
or U30 (N_30,In_187,In_456);
nor U31 (N_31,In_355,In_207);
xor U32 (N_32,In_341,In_237);
and U33 (N_33,In_220,In_50);
nand U34 (N_34,In_418,In_306);
and U35 (N_35,In_308,In_54);
or U36 (N_36,In_320,In_430);
nor U37 (N_37,In_286,In_330);
nand U38 (N_38,In_264,In_449);
nor U39 (N_39,In_261,In_463);
nor U40 (N_40,In_338,In_112);
nor U41 (N_41,In_2,In_119);
and U42 (N_42,In_460,In_485);
nor U43 (N_43,In_285,In_380);
nand U44 (N_44,In_262,In_77);
or U45 (N_45,In_452,In_97);
nand U46 (N_46,In_468,In_91);
and U47 (N_47,In_335,In_227);
and U48 (N_48,In_190,In_210);
nor U49 (N_49,In_305,In_126);
or U50 (N_50,In_121,In_69);
and U51 (N_51,In_168,In_76);
nand U52 (N_52,In_75,In_226);
or U53 (N_53,In_357,In_133);
nor U54 (N_54,In_369,In_302);
nand U55 (N_55,In_202,In_477);
nand U56 (N_56,In_358,In_412);
or U57 (N_57,In_115,In_211);
nor U58 (N_58,In_379,In_385);
and U59 (N_59,In_61,In_426);
nand U60 (N_60,In_491,In_32);
or U61 (N_61,In_346,In_185);
nor U62 (N_62,In_22,In_255);
or U63 (N_63,In_478,In_177);
and U64 (N_64,In_221,In_86);
xnor U65 (N_65,In_57,In_103);
nand U66 (N_66,In_323,In_213);
nor U67 (N_67,In_267,In_182);
nand U68 (N_68,In_333,In_311);
nand U69 (N_69,In_301,In_38);
nor U70 (N_70,In_464,In_107);
nand U71 (N_71,In_21,In_8);
and U72 (N_72,In_28,In_81);
or U73 (N_73,In_139,In_291);
or U74 (N_74,In_295,In_328);
nor U75 (N_75,In_499,In_170);
and U76 (N_76,In_140,In_319);
nand U77 (N_77,In_162,In_425);
and U78 (N_78,In_391,In_399);
nand U79 (N_79,In_206,In_496);
nor U80 (N_80,In_455,In_334);
and U81 (N_81,In_242,In_395);
nor U82 (N_82,In_365,In_321);
nand U83 (N_83,In_152,In_367);
nor U84 (N_84,In_36,In_376);
and U85 (N_85,In_439,In_431);
nand U86 (N_86,In_197,In_117);
and U87 (N_87,In_483,In_189);
or U88 (N_88,In_396,In_290);
nand U89 (N_89,In_183,In_422);
nor U90 (N_90,In_363,In_146);
and U91 (N_91,In_85,In_224);
xor U92 (N_92,In_7,In_157);
or U93 (N_93,In_176,In_249);
nand U94 (N_94,In_490,In_84);
and U95 (N_95,In_470,In_1);
nor U96 (N_96,In_52,In_444);
nor U97 (N_97,In_179,In_10);
nand U98 (N_98,In_467,In_386);
nand U99 (N_99,In_186,In_437);
or U100 (N_100,In_108,In_448);
nor U101 (N_101,In_174,In_150);
and U102 (N_102,In_299,In_457);
and U103 (N_103,In_400,In_70);
and U104 (N_104,In_474,In_287);
nor U105 (N_105,In_482,In_34);
nand U106 (N_106,In_26,In_284);
nand U107 (N_107,In_347,In_266);
nor U108 (N_108,In_178,In_229);
nand U109 (N_109,In_368,In_411);
and U110 (N_110,In_390,In_349);
nor U111 (N_111,In_15,In_199);
and U112 (N_112,In_447,In_198);
nand U113 (N_113,In_331,In_353);
nand U114 (N_114,In_23,In_292);
nand U115 (N_115,In_99,In_248);
or U116 (N_116,In_53,In_337);
or U117 (N_117,In_72,In_359);
nand U118 (N_118,In_317,In_120);
and U119 (N_119,In_332,In_200);
or U120 (N_120,In_461,In_388);
nor U121 (N_121,In_424,In_298);
nor U122 (N_122,In_88,In_90);
nor U123 (N_123,In_49,In_5);
nor U124 (N_124,In_175,In_89);
nand U125 (N_125,In_279,In_445);
or U126 (N_126,In_79,In_41);
xor U127 (N_127,In_165,In_137);
and U128 (N_128,In_124,In_263);
nand U129 (N_129,In_345,In_453);
and U130 (N_130,In_394,In_135);
and U131 (N_131,In_381,In_173);
nand U132 (N_132,In_494,In_458);
nand U133 (N_133,In_472,In_180);
nor U134 (N_134,In_459,In_87);
nor U135 (N_135,In_233,In_428);
or U136 (N_136,In_475,In_436);
nor U137 (N_137,In_236,In_71);
nand U138 (N_138,In_143,In_476);
and U139 (N_139,In_343,In_16);
nor U140 (N_140,In_232,In_392);
nand U141 (N_141,In_313,In_9);
nand U142 (N_142,In_169,In_94);
nor U143 (N_143,In_148,In_111);
xor U144 (N_144,In_272,In_141);
and U145 (N_145,In_276,In_372);
nor U146 (N_146,In_66,In_6);
or U147 (N_147,In_442,In_203);
nor U148 (N_148,In_193,In_127);
and U149 (N_149,In_132,In_309);
or U150 (N_150,In_404,In_218);
nand U151 (N_151,In_300,In_465);
or U152 (N_152,In_450,In_217);
and U153 (N_153,In_209,In_373);
nor U154 (N_154,In_405,In_487);
nor U155 (N_155,In_13,In_134);
nand U156 (N_156,In_486,In_149);
or U157 (N_157,In_131,In_366);
or U158 (N_158,In_223,In_253);
and U159 (N_159,In_116,In_407);
and U160 (N_160,In_113,In_382);
or U161 (N_161,In_110,In_219);
and U162 (N_162,In_244,In_238);
nor U163 (N_163,In_344,In_225);
nand U164 (N_164,In_257,In_20);
nand U165 (N_165,In_326,In_409);
nand U166 (N_166,In_294,In_147);
and U167 (N_167,In_283,In_440);
nor U168 (N_168,In_351,In_446);
nor U169 (N_169,In_275,In_316);
and U170 (N_170,In_327,In_39);
and U171 (N_171,In_130,In_56);
or U172 (N_172,In_350,In_280);
or U173 (N_173,In_212,In_105);
xor U174 (N_174,In_469,In_63);
or U175 (N_175,In_4,In_128);
or U176 (N_176,In_214,In_297);
or U177 (N_177,In_51,In_0);
nor U178 (N_178,In_246,In_205);
nor U179 (N_179,In_64,In_289);
and U180 (N_180,In_401,In_136);
nor U181 (N_181,In_378,In_166);
nand U182 (N_182,In_55,In_167);
and U183 (N_183,In_83,In_427);
nand U184 (N_184,In_270,In_435);
xnor U185 (N_185,In_312,In_420);
nor U186 (N_186,In_259,In_315);
nor U187 (N_187,In_278,In_204);
xor U188 (N_188,In_479,In_239);
or U189 (N_189,In_473,In_118);
and U190 (N_190,In_222,In_415);
nand U191 (N_191,In_397,In_288);
nor U192 (N_192,In_234,In_159);
and U193 (N_193,In_432,In_241);
nand U194 (N_194,In_413,In_48);
or U195 (N_195,In_296,In_434);
and U196 (N_196,In_268,In_389);
and U197 (N_197,In_78,In_14);
xnor U198 (N_198,In_342,In_11);
nand U199 (N_199,In_163,In_123);
nand U200 (N_200,N_83,N_131);
and U201 (N_201,N_102,N_30);
or U202 (N_202,In_421,N_133);
or U203 (N_203,N_14,N_110);
nor U204 (N_204,N_18,N_104);
and U205 (N_205,N_29,N_101);
xnor U206 (N_206,N_90,In_95);
nand U207 (N_207,N_4,In_258);
nor U208 (N_208,N_116,In_495);
nand U209 (N_209,N_132,N_144);
or U210 (N_210,N_49,N_135);
and U211 (N_211,In_42,N_92);
nand U212 (N_212,N_6,N_169);
nand U213 (N_213,N_158,N_123);
nand U214 (N_214,N_122,N_148);
nand U215 (N_215,N_74,N_59);
nand U216 (N_216,In_274,N_86);
nand U217 (N_217,N_114,N_126);
or U218 (N_218,N_195,In_144);
nor U219 (N_219,N_143,N_38);
nand U220 (N_220,In_354,N_198);
or U221 (N_221,N_188,In_438);
nor U222 (N_222,N_16,N_137);
or U223 (N_223,N_165,N_176);
nor U224 (N_224,In_489,N_52);
nor U225 (N_225,N_28,N_31);
and U226 (N_226,In_247,N_163);
nor U227 (N_227,In_43,In_33);
and U228 (N_228,N_51,N_111);
nand U229 (N_229,N_178,N_24);
nor U230 (N_230,N_109,In_348);
nand U231 (N_231,N_68,N_182);
nor U232 (N_232,In_497,N_50);
nor U233 (N_233,In_160,N_61);
nand U234 (N_234,N_11,N_120);
or U235 (N_235,In_145,N_22);
nor U236 (N_236,N_112,N_185);
or U237 (N_237,In_153,In_31);
nand U238 (N_238,In_138,N_177);
nand U239 (N_239,In_92,In_73);
and U240 (N_240,In_429,N_119);
nor U241 (N_241,N_89,N_161);
or U242 (N_242,N_121,N_162);
or U243 (N_243,In_3,In_18);
or U244 (N_244,N_125,N_67);
nand U245 (N_245,In_377,In_68);
nor U246 (N_246,N_80,In_340);
or U247 (N_247,N_150,N_147);
and U248 (N_248,N_19,In_47);
nand U249 (N_249,N_48,N_3);
and U250 (N_250,N_7,N_85);
nor U251 (N_251,N_26,N_155);
or U252 (N_252,In_481,In_375);
and U253 (N_253,N_186,N_136);
nand U254 (N_254,In_96,In_216);
and U255 (N_255,In_45,N_97);
nor U256 (N_256,N_175,N_1);
and U257 (N_257,N_94,In_104);
nor U258 (N_258,In_314,In_101);
or U259 (N_259,N_187,In_228);
nand U260 (N_260,N_70,N_12);
and U261 (N_261,N_69,N_39);
and U262 (N_262,In_252,In_188);
and U263 (N_263,In_240,N_42);
nor U264 (N_264,N_34,In_30);
xor U265 (N_265,N_8,In_492);
nor U266 (N_266,N_32,N_15);
or U267 (N_267,N_160,N_103);
or U268 (N_268,In_260,N_99);
xnor U269 (N_269,In_208,N_105);
and U270 (N_270,In_484,N_25);
and U271 (N_271,In_12,N_145);
nor U272 (N_272,N_33,N_134);
and U273 (N_273,In_109,N_192);
nand U274 (N_274,N_5,N_157);
nand U275 (N_275,N_193,N_9);
or U276 (N_276,N_139,In_417);
nor U277 (N_277,In_80,N_167);
and U278 (N_278,In_362,In_370);
nand U279 (N_279,N_91,N_181);
and U280 (N_280,N_66,N_172);
nand U281 (N_281,N_130,N_17);
nand U282 (N_282,N_196,In_243);
or U283 (N_283,In_192,In_498);
nand U284 (N_284,In_265,In_451);
and U285 (N_285,N_168,N_153);
nor U286 (N_286,In_374,In_184);
or U287 (N_287,N_164,In_125);
and U288 (N_288,N_191,N_53);
nor U289 (N_289,In_387,N_190);
and U290 (N_290,N_45,N_95);
or U291 (N_291,N_63,N_118);
xor U292 (N_292,N_71,N_107);
and U293 (N_293,N_152,N_76);
nor U294 (N_294,In_324,N_170);
nand U295 (N_295,N_142,N_141);
nand U296 (N_296,N_149,N_2);
nand U297 (N_297,N_82,N_146);
nor U298 (N_298,N_75,N_40);
nand U299 (N_299,N_128,In_74);
nand U300 (N_300,In_65,N_78);
nor U301 (N_301,N_20,In_230);
or U302 (N_302,N_81,N_73);
nand U303 (N_303,N_84,In_303);
nor U304 (N_304,N_36,In_102);
nand U305 (N_305,N_21,N_179);
nor U306 (N_306,N_98,In_398);
or U307 (N_307,In_250,N_106);
nand U308 (N_308,N_46,In_277);
or U309 (N_309,In_60,N_184);
or U310 (N_310,N_199,N_88);
nand U311 (N_311,N_13,N_37);
or U312 (N_312,N_180,N_55);
or U313 (N_313,N_113,In_44);
or U314 (N_314,N_58,In_215);
and U315 (N_315,In_443,In_307);
nand U316 (N_316,In_235,N_43);
nor U317 (N_317,In_384,N_0);
nor U318 (N_318,In_156,N_60);
nor U319 (N_319,In_383,In_93);
or U320 (N_320,In_423,N_72);
or U321 (N_321,In_19,In_29);
or U322 (N_322,In_196,N_174);
nor U323 (N_323,In_27,N_62);
or U324 (N_324,N_87,N_173);
nor U325 (N_325,In_256,In_466);
and U326 (N_326,N_117,N_154);
and U327 (N_327,N_64,N_129);
and U328 (N_328,N_138,N_77);
nor U329 (N_329,N_10,N_27);
or U330 (N_330,In_480,N_115);
and U331 (N_331,N_41,N_140);
or U332 (N_332,N_96,N_197);
or U333 (N_333,N_54,N_183);
nand U334 (N_334,N_108,In_142);
nand U335 (N_335,N_159,In_408);
nor U336 (N_336,N_100,N_57);
or U337 (N_337,N_47,N_35);
or U338 (N_338,In_46,N_189);
or U339 (N_339,N_124,In_269);
nor U340 (N_340,In_416,N_56);
nand U341 (N_341,In_24,In_360);
nor U342 (N_342,In_454,In_371);
nor U343 (N_343,N_93,N_151);
and U344 (N_344,In_339,In_251);
nor U345 (N_345,N_156,N_194);
or U346 (N_346,In_161,N_127);
nor U347 (N_347,N_44,N_65);
and U348 (N_348,N_23,N_171);
nand U349 (N_349,N_79,N_166);
nor U350 (N_350,In_416,N_99);
nor U351 (N_351,N_18,In_417);
nor U352 (N_352,N_49,N_192);
or U353 (N_353,In_481,N_40);
and U354 (N_354,N_187,In_125);
nand U355 (N_355,In_145,In_269);
nand U356 (N_356,N_158,N_184);
xor U357 (N_357,N_132,N_15);
nor U358 (N_358,N_181,N_6);
and U359 (N_359,In_161,N_57);
or U360 (N_360,N_51,N_77);
and U361 (N_361,N_20,N_153);
nor U362 (N_362,N_74,N_14);
nand U363 (N_363,N_161,In_497);
nor U364 (N_364,N_39,In_92);
or U365 (N_365,N_24,In_408);
and U366 (N_366,N_192,N_51);
nor U367 (N_367,In_184,N_62);
and U368 (N_368,N_45,In_354);
nand U369 (N_369,N_106,N_82);
and U370 (N_370,N_10,In_31);
nor U371 (N_371,In_80,N_53);
xnor U372 (N_372,In_384,In_451);
nand U373 (N_373,N_61,In_33);
or U374 (N_374,N_75,In_398);
nor U375 (N_375,N_55,N_76);
nor U376 (N_376,In_3,N_158);
nor U377 (N_377,N_190,In_43);
nand U378 (N_378,In_12,In_92);
nor U379 (N_379,In_362,In_454);
nor U380 (N_380,In_429,N_41);
or U381 (N_381,N_109,N_57);
nand U382 (N_382,N_157,In_12);
nand U383 (N_383,In_480,In_19);
nand U384 (N_384,N_64,N_24);
nand U385 (N_385,In_362,N_196);
and U386 (N_386,N_87,In_377);
and U387 (N_387,In_247,In_256);
nor U388 (N_388,N_38,N_40);
nor U389 (N_389,In_256,N_187);
nor U390 (N_390,In_80,N_5);
and U391 (N_391,N_54,N_163);
and U392 (N_392,N_122,N_133);
or U393 (N_393,N_172,N_160);
or U394 (N_394,N_18,N_125);
nand U395 (N_395,In_398,In_230);
or U396 (N_396,N_68,N_79);
or U397 (N_397,In_443,In_498);
nand U398 (N_398,In_383,In_92);
nor U399 (N_399,N_89,N_30);
or U400 (N_400,N_243,N_282);
nor U401 (N_401,N_383,N_257);
nand U402 (N_402,N_202,N_399);
and U403 (N_403,N_318,N_274);
and U404 (N_404,N_323,N_371);
nand U405 (N_405,N_375,N_290);
nand U406 (N_406,N_298,N_292);
nor U407 (N_407,N_222,N_204);
nand U408 (N_408,N_254,N_273);
nand U409 (N_409,N_310,N_379);
and U410 (N_410,N_262,N_213);
or U411 (N_411,N_387,N_330);
nor U412 (N_412,N_229,N_244);
or U413 (N_413,N_289,N_281);
or U414 (N_414,N_346,N_258);
nand U415 (N_415,N_362,N_252);
nand U416 (N_416,N_238,N_391);
nor U417 (N_417,N_361,N_333);
and U418 (N_418,N_317,N_366);
or U419 (N_419,N_363,N_340);
and U420 (N_420,N_368,N_339);
nor U421 (N_421,N_219,N_311);
nor U422 (N_422,N_315,N_269);
nand U423 (N_423,N_365,N_265);
nor U424 (N_424,N_327,N_230);
nor U425 (N_425,N_291,N_306);
nand U426 (N_426,N_266,N_297);
nand U427 (N_427,N_216,N_344);
or U428 (N_428,N_353,N_351);
or U429 (N_429,N_296,N_329);
nor U430 (N_430,N_369,N_355);
and U431 (N_431,N_287,N_388);
nor U432 (N_432,N_264,N_343);
xor U433 (N_433,N_386,N_352);
or U434 (N_434,N_232,N_381);
and U435 (N_435,N_288,N_247);
nand U436 (N_436,N_338,N_201);
and U437 (N_437,N_218,N_356);
and U438 (N_438,N_337,N_332);
xnor U439 (N_439,N_320,N_223);
and U440 (N_440,N_276,N_234);
and U441 (N_441,N_205,N_284);
or U442 (N_442,N_253,N_240);
or U443 (N_443,N_305,N_394);
or U444 (N_444,N_294,N_303);
nand U445 (N_445,N_396,N_220);
or U446 (N_446,N_380,N_341);
nor U447 (N_447,N_331,N_214);
nand U448 (N_448,N_259,N_349);
and U449 (N_449,N_228,N_283);
and U450 (N_450,N_279,N_233);
nand U451 (N_451,N_250,N_312);
or U452 (N_452,N_326,N_207);
nor U453 (N_453,N_321,N_256);
nor U454 (N_454,N_384,N_248);
nor U455 (N_455,N_300,N_322);
and U456 (N_456,N_370,N_374);
nand U457 (N_457,N_357,N_308);
nand U458 (N_458,N_324,N_200);
nand U459 (N_459,N_307,N_313);
nand U460 (N_460,N_389,N_293);
or U461 (N_461,N_237,N_221);
nand U462 (N_462,N_302,N_268);
nand U463 (N_463,N_226,N_208);
nand U464 (N_464,N_398,N_249);
nor U465 (N_465,N_217,N_325);
or U466 (N_466,N_342,N_359);
nor U467 (N_467,N_206,N_285);
or U468 (N_468,N_319,N_328);
nand U469 (N_469,N_203,N_275);
and U470 (N_470,N_367,N_316);
and U471 (N_471,N_295,N_397);
nand U472 (N_472,N_260,N_372);
nand U473 (N_473,N_224,N_314);
nand U474 (N_474,N_278,N_382);
nand U475 (N_475,N_212,N_280);
nor U476 (N_476,N_345,N_211);
nor U477 (N_477,N_286,N_245);
nor U478 (N_478,N_227,N_377);
and U479 (N_479,N_239,N_309);
nand U480 (N_480,N_373,N_231);
nand U481 (N_481,N_263,N_225);
and U482 (N_482,N_364,N_336);
and U483 (N_483,N_390,N_236);
nor U484 (N_484,N_235,N_304);
and U485 (N_485,N_360,N_251);
nor U486 (N_486,N_277,N_299);
nor U487 (N_487,N_385,N_215);
or U488 (N_488,N_271,N_334);
or U489 (N_489,N_358,N_209);
nand U490 (N_490,N_392,N_241);
nor U491 (N_491,N_246,N_270);
or U492 (N_492,N_267,N_301);
or U493 (N_493,N_350,N_395);
nor U494 (N_494,N_378,N_210);
or U495 (N_495,N_393,N_261);
and U496 (N_496,N_348,N_354);
xnor U497 (N_497,N_272,N_242);
and U498 (N_498,N_255,N_347);
or U499 (N_499,N_335,N_376);
nor U500 (N_500,N_338,N_394);
and U501 (N_501,N_304,N_319);
and U502 (N_502,N_236,N_345);
nand U503 (N_503,N_273,N_308);
nor U504 (N_504,N_392,N_370);
nand U505 (N_505,N_245,N_241);
and U506 (N_506,N_365,N_245);
and U507 (N_507,N_234,N_264);
nand U508 (N_508,N_377,N_334);
or U509 (N_509,N_215,N_354);
xor U510 (N_510,N_326,N_302);
or U511 (N_511,N_348,N_356);
or U512 (N_512,N_223,N_259);
and U513 (N_513,N_382,N_395);
nand U514 (N_514,N_371,N_281);
or U515 (N_515,N_363,N_236);
xnor U516 (N_516,N_308,N_260);
or U517 (N_517,N_229,N_252);
nor U518 (N_518,N_208,N_377);
and U519 (N_519,N_241,N_293);
nand U520 (N_520,N_294,N_220);
or U521 (N_521,N_328,N_345);
nand U522 (N_522,N_242,N_204);
or U523 (N_523,N_273,N_303);
or U524 (N_524,N_337,N_384);
nor U525 (N_525,N_234,N_261);
or U526 (N_526,N_272,N_330);
nand U527 (N_527,N_228,N_216);
nor U528 (N_528,N_397,N_364);
and U529 (N_529,N_218,N_387);
or U530 (N_530,N_386,N_335);
nor U531 (N_531,N_358,N_248);
nand U532 (N_532,N_248,N_341);
nand U533 (N_533,N_385,N_316);
and U534 (N_534,N_356,N_333);
and U535 (N_535,N_270,N_215);
or U536 (N_536,N_209,N_325);
nand U537 (N_537,N_329,N_222);
nand U538 (N_538,N_254,N_344);
or U539 (N_539,N_201,N_237);
nor U540 (N_540,N_387,N_357);
nor U541 (N_541,N_330,N_214);
or U542 (N_542,N_398,N_327);
nor U543 (N_543,N_312,N_217);
xnor U544 (N_544,N_224,N_293);
nor U545 (N_545,N_352,N_373);
nor U546 (N_546,N_388,N_223);
nor U547 (N_547,N_362,N_215);
nand U548 (N_548,N_291,N_275);
nand U549 (N_549,N_239,N_367);
or U550 (N_550,N_248,N_349);
nor U551 (N_551,N_273,N_312);
nand U552 (N_552,N_367,N_327);
or U553 (N_553,N_258,N_389);
and U554 (N_554,N_371,N_248);
nand U555 (N_555,N_392,N_331);
or U556 (N_556,N_387,N_222);
and U557 (N_557,N_241,N_398);
and U558 (N_558,N_282,N_233);
or U559 (N_559,N_248,N_246);
nand U560 (N_560,N_282,N_238);
or U561 (N_561,N_330,N_327);
nor U562 (N_562,N_229,N_386);
xor U563 (N_563,N_389,N_298);
nor U564 (N_564,N_363,N_395);
nand U565 (N_565,N_338,N_301);
or U566 (N_566,N_374,N_261);
nor U567 (N_567,N_313,N_231);
and U568 (N_568,N_217,N_276);
nor U569 (N_569,N_388,N_345);
nand U570 (N_570,N_351,N_211);
or U571 (N_571,N_284,N_301);
nand U572 (N_572,N_270,N_340);
and U573 (N_573,N_239,N_388);
nor U574 (N_574,N_241,N_257);
or U575 (N_575,N_312,N_330);
and U576 (N_576,N_332,N_394);
nor U577 (N_577,N_393,N_214);
nor U578 (N_578,N_370,N_288);
or U579 (N_579,N_312,N_387);
nor U580 (N_580,N_249,N_363);
nand U581 (N_581,N_256,N_364);
nor U582 (N_582,N_275,N_279);
and U583 (N_583,N_311,N_384);
and U584 (N_584,N_388,N_291);
nand U585 (N_585,N_291,N_295);
xor U586 (N_586,N_223,N_218);
nor U587 (N_587,N_390,N_276);
nor U588 (N_588,N_235,N_201);
and U589 (N_589,N_315,N_376);
nor U590 (N_590,N_321,N_380);
nand U591 (N_591,N_272,N_209);
or U592 (N_592,N_200,N_237);
nor U593 (N_593,N_302,N_233);
nor U594 (N_594,N_397,N_251);
nor U595 (N_595,N_205,N_251);
or U596 (N_596,N_245,N_201);
and U597 (N_597,N_223,N_214);
nand U598 (N_598,N_292,N_325);
or U599 (N_599,N_293,N_327);
nor U600 (N_600,N_426,N_534);
nor U601 (N_601,N_500,N_563);
nand U602 (N_602,N_495,N_553);
or U603 (N_603,N_415,N_531);
or U604 (N_604,N_570,N_412);
xnor U605 (N_605,N_581,N_505);
or U606 (N_606,N_428,N_576);
nand U607 (N_607,N_431,N_424);
nand U608 (N_608,N_434,N_451);
or U609 (N_609,N_556,N_487);
or U610 (N_610,N_488,N_536);
nand U611 (N_611,N_577,N_420);
and U612 (N_612,N_520,N_594);
nand U613 (N_613,N_566,N_506);
or U614 (N_614,N_462,N_441);
or U615 (N_615,N_513,N_467);
nor U616 (N_616,N_571,N_548);
nand U617 (N_617,N_464,N_564);
or U618 (N_618,N_579,N_552);
xor U619 (N_619,N_595,N_419);
and U620 (N_620,N_546,N_459);
nand U621 (N_621,N_458,N_519);
nand U622 (N_622,N_423,N_489);
or U623 (N_623,N_475,N_549);
nor U624 (N_624,N_522,N_509);
nor U625 (N_625,N_598,N_568);
xnor U626 (N_626,N_528,N_562);
nand U627 (N_627,N_599,N_471);
and U628 (N_628,N_468,N_514);
nand U629 (N_629,N_532,N_446);
nand U630 (N_630,N_518,N_438);
nand U631 (N_631,N_567,N_422);
nor U632 (N_632,N_547,N_413);
and U633 (N_633,N_511,N_502);
or U634 (N_634,N_590,N_477);
nor U635 (N_635,N_524,N_486);
nor U636 (N_636,N_478,N_507);
nor U637 (N_637,N_543,N_515);
nor U638 (N_638,N_410,N_510);
and U639 (N_639,N_448,N_504);
nor U640 (N_640,N_530,N_542);
xnor U641 (N_641,N_596,N_593);
and U642 (N_642,N_527,N_537);
and U643 (N_643,N_481,N_587);
nor U644 (N_644,N_592,N_417);
or U645 (N_645,N_597,N_421);
nand U646 (N_646,N_484,N_470);
nor U647 (N_647,N_432,N_578);
nand U648 (N_648,N_582,N_437);
nand U649 (N_649,N_472,N_491);
nor U650 (N_650,N_474,N_463);
and U651 (N_651,N_516,N_435);
xor U652 (N_652,N_411,N_540);
or U653 (N_653,N_580,N_402);
nor U654 (N_654,N_447,N_541);
nand U655 (N_655,N_405,N_538);
nand U656 (N_656,N_400,N_430);
or U657 (N_657,N_450,N_454);
or U658 (N_658,N_457,N_558);
or U659 (N_659,N_429,N_469);
or U660 (N_660,N_533,N_535);
nand U661 (N_661,N_501,N_512);
nor U662 (N_662,N_574,N_452);
and U663 (N_663,N_529,N_557);
or U664 (N_664,N_465,N_496);
nor U665 (N_665,N_569,N_499);
nor U666 (N_666,N_401,N_550);
nor U667 (N_667,N_554,N_443);
nand U668 (N_668,N_503,N_460);
nand U669 (N_669,N_455,N_480);
or U670 (N_670,N_497,N_456);
xor U671 (N_671,N_584,N_427);
or U672 (N_672,N_561,N_485);
nand U673 (N_673,N_404,N_523);
nand U674 (N_674,N_589,N_433);
nor U675 (N_675,N_555,N_418);
or U676 (N_676,N_479,N_440);
and U677 (N_677,N_407,N_439);
nand U678 (N_678,N_409,N_575);
or U679 (N_679,N_508,N_573);
nor U680 (N_680,N_559,N_588);
nand U681 (N_681,N_493,N_545);
xor U682 (N_682,N_408,N_526);
nor U683 (N_683,N_414,N_585);
or U684 (N_684,N_416,N_544);
and U685 (N_685,N_591,N_539);
or U686 (N_686,N_473,N_572);
or U687 (N_687,N_442,N_517);
nor U688 (N_688,N_551,N_453);
nor U689 (N_689,N_436,N_461);
nand U690 (N_690,N_466,N_494);
nand U691 (N_691,N_406,N_483);
nor U692 (N_692,N_521,N_490);
nor U693 (N_693,N_560,N_444);
nor U694 (N_694,N_403,N_449);
and U695 (N_695,N_586,N_498);
and U696 (N_696,N_425,N_482);
nand U697 (N_697,N_476,N_492);
or U698 (N_698,N_565,N_445);
nor U699 (N_699,N_525,N_583);
nor U700 (N_700,N_585,N_571);
or U701 (N_701,N_458,N_450);
and U702 (N_702,N_537,N_440);
nor U703 (N_703,N_431,N_548);
or U704 (N_704,N_573,N_577);
nand U705 (N_705,N_542,N_514);
or U706 (N_706,N_533,N_519);
xor U707 (N_707,N_561,N_580);
or U708 (N_708,N_570,N_460);
nor U709 (N_709,N_583,N_565);
nand U710 (N_710,N_521,N_552);
and U711 (N_711,N_580,N_418);
nor U712 (N_712,N_542,N_522);
or U713 (N_713,N_549,N_509);
and U714 (N_714,N_542,N_470);
or U715 (N_715,N_483,N_513);
or U716 (N_716,N_431,N_513);
nand U717 (N_717,N_477,N_533);
or U718 (N_718,N_506,N_418);
xnor U719 (N_719,N_596,N_500);
nor U720 (N_720,N_592,N_556);
and U721 (N_721,N_453,N_558);
or U722 (N_722,N_463,N_473);
nand U723 (N_723,N_446,N_454);
nor U724 (N_724,N_408,N_484);
and U725 (N_725,N_562,N_584);
and U726 (N_726,N_540,N_449);
nor U727 (N_727,N_520,N_438);
and U728 (N_728,N_405,N_403);
nor U729 (N_729,N_492,N_529);
nand U730 (N_730,N_475,N_594);
and U731 (N_731,N_431,N_430);
nand U732 (N_732,N_405,N_524);
or U733 (N_733,N_470,N_582);
nor U734 (N_734,N_586,N_512);
nand U735 (N_735,N_561,N_568);
and U736 (N_736,N_524,N_550);
or U737 (N_737,N_536,N_585);
and U738 (N_738,N_503,N_565);
xor U739 (N_739,N_429,N_550);
and U740 (N_740,N_432,N_417);
or U741 (N_741,N_556,N_421);
nor U742 (N_742,N_432,N_437);
nor U743 (N_743,N_493,N_470);
nand U744 (N_744,N_567,N_466);
nor U745 (N_745,N_525,N_543);
and U746 (N_746,N_543,N_429);
nor U747 (N_747,N_461,N_417);
or U748 (N_748,N_510,N_489);
nand U749 (N_749,N_464,N_413);
and U750 (N_750,N_521,N_482);
and U751 (N_751,N_510,N_566);
nor U752 (N_752,N_454,N_442);
and U753 (N_753,N_570,N_592);
or U754 (N_754,N_460,N_599);
nor U755 (N_755,N_484,N_495);
or U756 (N_756,N_553,N_451);
nor U757 (N_757,N_459,N_453);
nand U758 (N_758,N_455,N_486);
nand U759 (N_759,N_408,N_465);
or U760 (N_760,N_477,N_525);
nand U761 (N_761,N_501,N_588);
or U762 (N_762,N_518,N_567);
xnor U763 (N_763,N_504,N_587);
nor U764 (N_764,N_506,N_417);
nand U765 (N_765,N_407,N_529);
and U766 (N_766,N_515,N_472);
or U767 (N_767,N_547,N_414);
nor U768 (N_768,N_451,N_513);
or U769 (N_769,N_432,N_568);
nand U770 (N_770,N_459,N_439);
nand U771 (N_771,N_533,N_507);
and U772 (N_772,N_496,N_502);
or U773 (N_773,N_462,N_431);
nor U774 (N_774,N_565,N_422);
nor U775 (N_775,N_562,N_482);
and U776 (N_776,N_428,N_481);
nand U777 (N_777,N_482,N_591);
nand U778 (N_778,N_431,N_472);
nor U779 (N_779,N_599,N_435);
and U780 (N_780,N_448,N_586);
or U781 (N_781,N_463,N_431);
or U782 (N_782,N_567,N_570);
nand U783 (N_783,N_421,N_452);
nand U784 (N_784,N_587,N_459);
and U785 (N_785,N_537,N_417);
or U786 (N_786,N_532,N_502);
or U787 (N_787,N_497,N_579);
and U788 (N_788,N_446,N_569);
and U789 (N_789,N_478,N_418);
nor U790 (N_790,N_424,N_546);
xnor U791 (N_791,N_454,N_465);
nor U792 (N_792,N_432,N_466);
nor U793 (N_793,N_442,N_597);
nand U794 (N_794,N_573,N_402);
or U795 (N_795,N_592,N_454);
or U796 (N_796,N_597,N_439);
or U797 (N_797,N_538,N_586);
and U798 (N_798,N_576,N_546);
or U799 (N_799,N_402,N_420);
and U800 (N_800,N_606,N_657);
nor U801 (N_801,N_719,N_616);
nand U802 (N_802,N_627,N_776);
nor U803 (N_803,N_758,N_687);
nor U804 (N_804,N_675,N_750);
and U805 (N_805,N_619,N_706);
or U806 (N_806,N_645,N_771);
nor U807 (N_807,N_726,N_666);
and U808 (N_808,N_612,N_664);
and U809 (N_809,N_621,N_790);
nor U810 (N_810,N_695,N_755);
and U811 (N_811,N_744,N_669);
nand U812 (N_812,N_791,N_780);
and U813 (N_813,N_743,N_681);
nand U814 (N_814,N_752,N_734);
nand U815 (N_815,N_697,N_635);
nand U816 (N_816,N_717,N_650);
and U817 (N_817,N_633,N_673);
nand U818 (N_818,N_689,N_703);
or U819 (N_819,N_761,N_602);
or U820 (N_820,N_660,N_764);
nand U821 (N_821,N_668,N_763);
or U822 (N_822,N_756,N_715);
xnor U823 (N_823,N_747,N_672);
nor U824 (N_824,N_654,N_759);
nor U825 (N_825,N_735,N_708);
nor U826 (N_826,N_642,N_722);
or U827 (N_827,N_655,N_624);
or U828 (N_828,N_623,N_682);
and U829 (N_829,N_614,N_658);
nand U830 (N_830,N_607,N_725);
nand U831 (N_831,N_718,N_659);
nand U832 (N_832,N_617,N_630);
and U833 (N_833,N_638,N_685);
or U834 (N_834,N_772,N_696);
nand U835 (N_835,N_698,N_622);
nand U836 (N_836,N_766,N_647);
or U837 (N_837,N_733,N_707);
and U838 (N_838,N_637,N_694);
nor U839 (N_839,N_667,N_782);
and U840 (N_840,N_693,N_649);
and U841 (N_841,N_680,N_628);
and U842 (N_842,N_720,N_605);
nor U843 (N_843,N_787,N_721);
and U844 (N_844,N_651,N_674);
or U845 (N_845,N_727,N_652);
and U846 (N_846,N_710,N_795);
and U847 (N_847,N_610,N_777);
nor U848 (N_848,N_736,N_737);
nand U849 (N_849,N_792,N_789);
nor U850 (N_850,N_705,N_670);
nor U851 (N_851,N_634,N_648);
nand U852 (N_852,N_701,N_671);
nor U853 (N_853,N_778,N_676);
nor U854 (N_854,N_631,N_641);
nor U855 (N_855,N_793,N_765);
nand U856 (N_856,N_760,N_656);
nand U857 (N_857,N_691,N_798);
and U858 (N_858,N_751,N_769);
or U859 (N_859,N_746,N_677);
or U860 (N_860,N_644,N_709);
nor U861 (N_861,N_723,N_797);
nand U862 (N_862,N_714,N_609);
nand U863 (N_863,N_662,N_704);
or U864 (N_864,N_712,N_732);
nand U865 (N_865,N_601,N_740);
and U866 (N_866,N_640,N_724);
nand U867 (N_867,N_779,N_702);
nor U868 (N_868,N_742,N_690);
and U869 (N_869,N_653,N_773);
nand U870 (N_870,N_794,N_679);
and U871 (N_871,N_786,N_783);
nand U872 (N_872,N_731,N_613);
nor U873 (N_873,N_762,N_788);
nand U874 (N_874,N_741,N_781);
or U875 (N_875,N_745,N_775);
and U876 (N_876,N_618,N_713);
nand U877 (N_877,N_770,N_684);
and U878 (N_878,N_604,N_620);
nor U879 (N_879,N_785,N_636);
and U880 (N_880,N_753,N_799);
nor U881 (N_881,N_629,N_646);
or U882 (N_882,N_615,N_688);
nor U883 (N_883,N_716,N_728);
and U884 (N_884,N_711,N_639);
nand U885 (N_885,N_796,N_663);
nor U886 (N_886,N_757,N_748);
and U887 (N_887,N_774,N_767);
nor U888 (N_888,N_739,N_643);
or U889 (N_889,N_608,N_611);
nor U890 (N_890,N_700,N_626);
or U891 (N_891,N_665,N_600);
nor U892 (N_892,N_632,N_754);
or U893 (N_893,N_784,N_730);
nand U894 (N_894,N_625,N_749);
nor U895 (N_895,N_738,N_603);
and U896 (N_896,N_692,N_699);
nand U897 (N_897,N_678,N_683);
and U898 (N_898,N_661,N_686);
nand U899 (N_899,N_768,N_729);
nor U900 (N_900,N_751,N_749);
and U901 (N_901,N_642,N_719);
nand U902 (N_902,N_735,N_641);
nor U903 (N_903,N_745,N_735);
nand U904 (N_904,N_600,N_735);
nand U905 (N_905,N_724,N_647);
and U906 (N_906,N_799,N_783);
or U907 (N_907,N_648,N_611);
nand U908 (N_908,N_602,N_772);
or U909 (N_909,N_690,N_775);
and U910 (N_910,N_747,N_625);
or U911 (N_911,N_770,N_734);
nand U912 (N_912,N_735,N_698);
nand U913 (N_913,N_747,N_648);
nand U914 (N_914,N_794,N_733);
nand U915 (N_915,N_642,N_621);
and U916 (N_916,N_740,N_635);
or U917 (N_917,N_619,N_742);
and U918 (N_918,N_668,N_726);
nor U919 (N_919,N_659,N_622);
and U920 (N_920,N_786,N_737);
or U921 (N_921,N_696,N_726);
nand U922 (N_922,N_675,N_784);
and U923 (N_923,N_671,N_738);
nand U924 (N_924,N_605,N_692);
or U925 (N_925,N_622,N_689);
xnor U926 (N_926,N_756,N_685);
or U927 (N_927,N_778,N_644);
and U928 (N_928,N_645,N_740);
or U929 (N_929,N_632,N_706);
nor U930 (N_930,N_650,N_606);
or U931 (N_931,N_691,N_634);
nor U932 (N_932,N_698,N_633);
and U933 (N_933,N_690,N_696);
xor U934 (N_934,N_701,N_722);
nand U935 (N_935,N_608,N_793);
or U936 (N_936,N_700,N_728);
nor U937 (N_937,N_786,N_729);
nor U938 (N_938,N_774,N_703);
nand U939 (N_939,N_682,N_626);
nor U940 (N_940,N_662,N_781);
nand U941 (N_941,N_757,N_737);
or U942 (N_942,N_651,N_617);
nand U943 (N_943,N_747,N_652);
nor U944 (N_944,N_646,N_623);
nand U945 (N_945,N_642,N_626);
nor U946 (N_946,N_614,N_696);
or U947 (N_947,N_689,N_739);
nand U948 (N_948,N_791,N_771);
nand U949 (N_949,N_688,N_726);
or U950 (N_950,N_757,N_702);
or U951 (N_951,N_777,N_727);
nor U952 (N_952,N_677,N_699);
nor U953 (N_953,N_746,N_792);
and U954 (N_954,N_773,N_637);
and U955 (N_955,N_667,N_703);
xnor U956 (N_956,N_638,N_646);
nand U957 (N_957,N_670,N_751);
or U958 (N_958,N_779,N_610);
and U959 (N_959,N_622,N_747);
nor U960 (N_960,N_604,N_607);
nand U961 (N_961,N_613,N_622);
nand U962 (N_962,N_701,N_662);
nand U963 (N_963,N_695,N_771);
or U964 (N_964,N_670,N_606);
nand U965 (N_965,N_787,N_720);
nand U966 (N_966,N_634,N_723);
nor U967 (N_967,N_750,N_690);
nand U968 (N_968,N_609,N_784);
xnor U969 (N_969,N_606,N_701);
nand U970 (N_970,N_764,N_662);
and U971 (N_971,N_712,N_722);
nor U972 (N_972,N_736,N_684);
and U973 (N_973,N_638,N_718);
nand U974 (N_974,N_679,N_647);
nor U975 (N_975,N_764,N_692);
xnor U976 (N_976,N_781,N_713);
nand U977 (N_977,N_670,N_774);
or U978 (N_978,N_668,N_609);
nand U979 (N_979,N_727,N_683);
nor U980 (N_980,N_621,N_794);
nand U981 (N_981,N_702,N_769);
nand U982 (N_982,N_734,N_608);
nand U983 (N_983,N_624,N_662);
and U984 (N_984,N_719,N_737);
nand U985 (N_985,N_768,N_700);
and U986 (N_986,N_683,N_677);
nand U987 (N_987,N_708,N_751);
nand U988 (N_988,N_684,N_712);
or U989 (N_989,N_634,N_628);
nand U990 (N_990,N_776,N_684);
and U991 (N_991,N_703,N_709);
and U992 (N_992,N_631,N_785);
or U993 (N_993,N_623,N_729);
nor U994 (N_994,N_727,N_714);
nor U995 (N_995,N_771,N_661);
nand U996 (N_996,N_794,N_680);
nor U997 (N_997,N_719,N_721);
nand U998 (N_998,N_631,N_671);
and U999 (N_999,N_601,N_789);
or U1000 (N_1000,N_869,N_828);
and U1001 (N_1001,N_810,N_979);
or U1002 (N_1002,N_934,N_957);
or U1003 (N_1003,N_862,N_885);
nor U1004 (N_1004,N_803,N_981);
nor U1005 (N_1005,N_903,N_879);
nand U1006 (N_1006,N_834,N_887);
or U1007 (N_1007,N_889,N_893);
and U1008 (N_1008,N_839,N_856);
nor U1009 (N_1009,N_909,N_827);
nand U1010 (N_1010,N_987,N_994);
or U1011 (N_1011,N_884,N_843);
nand U1012 (N_1012,N_938,N_992);
nor U1013 (N_1013,N_896,N_949);
nor U1014 (N_1014,N_875,N_921);
or U1015 (N_1015,N_932,N_814);
and U1016 (N_1016,N_940,N_806);
nand U1017 (N_1017,N_818,N_958);
or U1018 (N_1018,N_945,N_824);
or U1019 (N_1019,N_937,N_815);
or U1020 (N_1020,N_941,N_916);
nand U1021 (N_1021,N_933,N_939);
nand U1022 (N_1022,N_892,N_836);
or U1023 (N_1023,N_956,N_978);
or U1024 (N_1024,N_913,N_915);
nor U1025 (N_1025,N_983,N_831);
or U1026 (N_1026,N_975,N_817);
or U1027 (N_1027,N_841,N_870);
nand U1028 (N_1028,N_891,N_936);
or U1029 (N_1029,N_962,N_928);
nor U1030 (N_1030,N_861,N_942);
and U1031 (N_1031,N_919,N_801);
nor U1032 (N_1032,N_972,N_966);
nand U1033 (N_1033,N_811,N_982);
nand U1034 (N_1034,N_859,N_820);
nor U1035 (N_1035,N_840,N_904);
or U1036 (N_1036,N_851,N_922);
or U1037 (N_1037,N_822,N_873);
and U1038 (N_1038,N_930,N_947);
nand U1039 (N_1039,N_901,N_865);
or U1040 (N_1040,N_849,N_914);
and U1041 (N_1041,N_995,N_826);
or U1042 (N_1042,N_882,N_895);
nand U1043 (N_1043,N_969,N_805);
and U1044 (N_1044,N_918,N_813);
and U1045 (N_1045,N_809,N_844);
and U1046 (N_1046,N_980,N_905);
nand U1047 (N_1047,N_943,N_830);
nand U1048 (N_1048,N_973,N_876);
nand U1049 (N_1049,N_886,N_991);
and U1050 (N_1050,N_935,N_967);
nor U1051 (N_1051,N_931,N_816);
nand U1052 (N_1052,N_977,N_868);
or U1053 (N_1053,N_976,N_911);
or U1054 (N_1054,N_898,N_883);
or U1055 (N_1055,N_946,N_954);
nor U1056 (N_1056,N_961,N_974);
or U1057 (N_1057,N_990,N_866);
or U1058 (N_1058,N_854,N_833);
nand U1059 (N_1059,N_800,N_852);
or U1060 (N_1060,N_965,N_952);
xnor U1061 (N_1061,N_984,N_855);
and U1062 (N_1062,N_920,N_821);
nand U1063 (N_1063,N_874,N_845);
nand U1064 (N_1064,N_917,N_912);
or U1065 (N_1065,N_910,N_835);
nand U1066 (N_1066,N_996,N_857);
nand U1067 (N_1067,N_838,N_871);
nor U1068 (N_1068,N_900,N_897);
nand U1069 (N_1069,N_877,N_899);
or U1070 (N_1070,N_823,N_890);
or U1071 (N_1071,N_825,N_960);
or U1072 (N_1072,N_986,N_955);
and U1073 (N_1073,N_858,N_927);
or U1074 (N_1074,N_950,N_880);
nor U1075 (N_1075,N_997,N_988);
nor U1076 (N_1076,N_964,N_999);
nand U1077 (N_1077,N_860,N_944);
nand U1078 (N_1078,N_863,N_894);
or U1079 (N_1079,N_832,N_878);
xnor U1080 (N_1080,N_872,N_985);
nor U1081 (N_1081,N_808,N_867);
or U1082 (N_1082,N_881,N_968);
nor U1083 (N_1083,N_802,N_829);
and U1084 (N_1084,N_929,N_902);
and U1085 (N_1085,N_847,N_959);
or U1086 (N_1086,N_837,N_953);
nand U1087 (N_1087,N_924,N_807);
or U1088 (N_1088,N_812,N_864);
or U1089 (N_1089,N_850,N_925);
nand U1090 (N_1090,N_998,N_906);
nand U1091 (N_1091,N_907,N_951);
nand U1092 (N_1092,N_989,N_908);
nand U1093 (N_1093,N_963,N_971);
or U1094 (N_1094,N_993,N_970);
nor U1095 (N_1095,N_926,N_948);
nor U1096 (N_1096,N_853,N_848);
and U1097 (N_1097,N_819,N_804);
and U1098 (N_1098,N_888,N_923);
nor U1099 (N_1099,N_846,N_842);
and U1100 (N_1100,N_808,N_901);
nor U1101 (N_1101,N_957,N_847);
or U1102 (N_1102,N_868,N_847);
xnor U1103 (N_1103,N_944,N_929);
and U1104 (N_1104,N_966,N_953);
and U1105 (N_1105,N_813,N_867);
nor U1106 (N_1106,N_837,N_878);
nand U1107 (N_1107,N_895,N_897);
or U1108 (N_1108,N_884,N_895);
nand U1109 (N_1109,N_820,N_890);
nor U1110 (N_1110,N_923,N_804);
or U1111 (N_1111,N_899,N_912);
nand U1112 (N_1112,N_840,N_902);
nand U1113 (N_1113,N_953,N_969);
and U1114 (N_1114,N_965,N_803);
nor U1115 (N_1115,N_978,N_895);
nand U1116 (N_1116,N_900,N_876);
or U1117 (N_1117,N_819,N_946);
or U1118 (N_1118,N_841,N_937);
nand U1119 (N_1119,N_988,N_882);
and U1120 (N_1120,N_932,N_809);
nand U1121 (N_1121,N_998,N_885);
or U1122 (N_1122,N_880,N_870);
nand U1123 (N_1123,N_813,N_932);
nor U1124 (N_1124,N_904,N_848);
nand U1125 (N_1125,N_875,N_903);
nand U1126 (N_1126,N_979,N_912);
and U1127 (N_1127,N_903,N_987);
nand U1128 (N_1128,N_810,N_827);
nand U1129 (N_1129,N_994,N_967);
and U1130 (N_1130,N_926,N_873);
or U1131 (N_1131,N_961,N_892);
nor U1132 (N_1132,N_880,N_884);
and U1133 (N_1133,N_942,N_860);
or U1134 (N_1134,N_826,N_886);
nand U1135 (N_1135,N_879,N_906);
or U1136 (N_1136,N_955,N_931);
nand U1137 (N_1137,N_992,N_869);
or U1138 (N_1138,N_834,N_908);
and U1139 (N_1139,N_965,N_848);
nand U1140 (N_1140,N_975,N_978);
or U1141 (N_1141,N_900,N_820);
nand U1142 (N_1142,N_852,N_941);
nand U1143 (N_1143,N_946,N_839);
or U1144 (N_1144,N_940,N_824);
or U1145 (N_1145,N_955,N_935);
nor U1146 (N_1146,N_823,N_820);
or U1147 (N_1147,N_912,N_937);
nor U1148 (N_1148,N_907,N_832);
and U1149 (N_1149,N_953,N_877);
or U1150 (N_1150,N_855,N_904);
nor U1151 (N_1151,N_983,N_824);
nor U1152 (N_1152,N_888,N_905);
and U1153 (N_1153,N_875,N_900);
nor U1154 (N_1154,N_806,N_814);
nor U1155 (N_1155,N_839,N_919);
and U1156 (N_1156,N_850,N_863);
or U1157 (N_1157,N_938,N_939);
nor U1158 (N_1158,N_945,N_907);
nor U1159 (N_1159,N_810,N_847);
and U1160 (N_1160,N_837,N_963);
or U1161 (N_1161,N_918,N_816);
and U1162 (N_1162,N_861,N_980);
and U1163 (N_1163,N_837,N_865);
and U1164 (N_1164,N_865,N_949);
nand U1165 (N_1165,N_878,N_880);
nand U1166 (N_1166,N_821,N_858);
and U1167 (N_1167,N_855,N_874);
or U1168 (N_1168,N_943,N_949);
and U1169 (N_1169,N_914,N_918);
nor U1170 (N_1170,N_940,N_992);
nand U1171 (N_1171,N_851,N_939);
nor U1172 (N_1172,N_895,N_833);
and U1173 (N_1173,N_960,N_862);
or U1174 (N_1174,N_968,N_916);
or U1175 (N_1175,N_880,N_862);
xnor U1176 (N_1176,N_897,N_858);
or U1177 (N_1177,N_890,N_951);
nand U1178 (N_1178,N_805,N_990);
nand U1179 (N_1179,N_961,N_808);
nor U1180 (N_1180,N_914,N_942);
nand U1181 (N_1181,N_838,N_832);
and U1182 (N_1182,N_939,N_815);
nand U1183 (N_1183,N_971,N_804);
nand U1184 (N_1184,N_965,N_822);
nand U1185 (N_1185,N_844,N_879);
nand U1186 (N_1186,N_807,N_911);
nand U1187 (N_1187,N_907,N_895);
nor U1188 (N_1188,N_988,N_992);
nor U1189 (N_1189,N_803,N_916);
nor U1190 (N_1190,N_890,N_937);
nand U1191 (N_1191,N_888,N_845);
and U1192 (N_1192,N_997,N_846);
xor U1193 (N_1193,N_857,N_901);
and U1194 (N_1194,N_909,N_854);
or U1195 (N_1195,N_945,N_957);
nor U1196 (N_1196,N_838,N_958);
nor U1197 (N_1197,N_876,N_865);
and U1198 (N_1198,N_846,N_966);
nand U1199 (N_1199,N_845,N_948);
or U1200 (N_1200,N_1153,N_1029);
or U1201 (N_1201,N_1083,N_1058);
or U1202 (N_1202,N_1109,N_1021);
nand U1203 (N_1203,N_1145,N_1057);
and U1204 (N_1204,N_1101,N_1114);
and U1205 (N_1205,N_1132,N_1089);
and U1206 (N_1206,N_1044,N_1187);
nor U1207 (N_1207,N_1139,N_1081);
nand U1208 (N_1208,N_1004,N_1036);
nand U1209 (N_1209,N_1067,N_1045);
and U1210 (N_1210,N_1129,N_1048);
nor U1211 (N_1211,N_1194,N_1174);
nand U1212 (N_1212,N_1092,N_1116);
and U1213 (N_1213,N_1049,N_1070);
nand U1214 (N_1214,N_1124,N_1150);
nor U1215 (N_1215,N_1078,N_1197);
and U1216 (N_1216,N_1010,N_1167);
nor U1217 (N_1217,N_1131,N_1025);
nor U1218 (N_1218,N_1159,N_1137);
or U1219 (N_1219,N_1123,N_1099);
or U1220 (N_1220,N_1063,N_1033);
nand U1221 (N_1221,N_1064,N_1154);
nor U1222 (N_1222,N_1051,N_1012);
nor U1223 (N_1223,N_1098,N_1176);
nand U1224 (N_1224,N_1052,N_1113);
nor U1225 (N_1225,N_1172,N_1162);
or U1226 (N_1226,N_1115,N_1108);
nor U1227 (N_1227,N_1066,N_1138);
and U1228 (N_1228,N_1195,N_1148);
nor U1229 (N_1229,N_1087,N_1095);
nand U1230 (N_1230,N_1163,N_1165);
nand U1231 (N_1231,N_1135,N_1190);
nand U1232 (N_1232,N_1017,N_1149);
nand U1233 (N_1233,N_1136,N_1074);
or U1234 (N_1234,N_1026,N_1014);
nand U1235 (N_1235,N_1024,N_1168);
or U1236 (N_1236,N_1022,N_1065);
and U1237 (N_1237,N_1133,N_1068);
nor U1238 (N_1238,N_1151,N_1047);
or U1239 (N_1239,N_1160,N_1015);
or U1240 (N_1240,N_1006,N_1055);
nand U1241 (N_1241,N_1179,N_1180);
or U1242 (N_1242,N_1102,N_1181);
nand U1243 (N_1243,N_1020,N_1001);
and U1244 (N_1244,N_1140,N_1002);
nor U1245 (N_1245,N_1091,N_1003);
or U1246 (N_1246,N_1126,N_1073);
nor U1247 (N_1247,N_1142,N_1097);
and U1248 (N_1248,N_1013,N_1103);
and U1249 (N_1249,N_1094,N_1143);
and U1250 (N_1250,N_1009,N_1127);
nor U1251 (N_1251,N_1042,N_1035);
nor U1252 (N_1252,N_1146,N_1090);
nand U1253 (N_1253,N_1037,N_1100);
nand U1254 (N_1254,N_1125,N_1188);
nor U1255 (N_1255,N_1183,N_1191);
and U1256 (N_1256,N_1059,N_1193);
or U1257 (N_1257,N_1107,N_1121);
and U1258 (N_1258,N_1186,N_1071);
or U1259 (N_1259,N_1199,N_1117);
nand U1260 (N_1260,N_1178,N_1106);
nor U1261 (N_1261,N_1040,N_1161);
or U1262 (N_1262,N_1079,N_1075);
and U1263 (N_1263,N_1104,N_1032);
or U1264 (N_1264,N_1060,N_1105);
or U1265 (N_1265,N_1118,N_1000);
or U1266 (N_1266,N_1096,N_1034);
or U1267 (N_1267,N_1011,N_1062);
nand U1268 (N_1268,N_1069,N_1158);
and U1269 (N_1269,N_1112,N_1182);
nor U1270 (N_1270,N_1085,N_1152);
nand U1271 (N_1271,N_1039,N_1076);
nand U1272 (N_1272,N_1166,N_1056);
nor U1273 (N_1273,N_1007,N_1041);
nand U1274 (N_1274,N_1005,N_1050);
xnor U1275 (N_1275,N_1027,N_1147);
nand U1276 (N_1276,N_1164,N_1061);
nor U1277 (N_1277,N_1170,N_1082);
xnor U1278 (N_1278,N_1054,N_1157);
nand U1279 (N_1279,N_1016,N_1023);
or U1280 (N_1280,N_1155,N_1008);
nand U1281 (N_1281,N_1171,N_1119);
nor U1282 (N_1282,N_1173,N_1088);
or U1283 (N_1283,N_1031,N_1189);
nor U1284 (N_1284,N_1093,N_1128);
nor U1285 (N_1285,N_1198,N_1072);
and U1286 (N_1286,N_1030,N_1084);
or U1287 (N_1287,N_1053,N_1028);
nor U1288 (N_1288,N_1086,N_1177);
and U1289 (N_1289,N_1156,N_1196);
nand U1290 (N_1290,N_1080,N_1184);
nor U1291 (N_1291,N_1185,N_1019);
nand U1292 (N_1292,N_1018,N_1043);
nor U1293 (N_1293,N_1192,N_1144);
and U1294 (N_1294,N_1038,N_1110);
nand U1295 (N_1295,N_1134,N_1120);
and U1296 (N_1296,N_1077,N_1169);
and U1297 (N_1297,N_1046,N_1175);
or U1298 (N_1298,N_1111,N_1141);
and U1299 (N_1299,N_1130,N_1122);
nor U1300 (N_1300,N_1062,N_1162);
or U1301 (N_1301,N_1147,N_1070);
xnor U1302 (N_1302,N_1042,N_1110);
nor U1303 (N_1303,N_1165,N_1080);
nor U1304 (N_1304,N_1104,N_1121);
and U1305 (N_1305,N_1060,N_1101);
nand U1306 (N_1306,N_1078,N_1083);
nor U1307 (N_1307,N_1046,N_1039);
nand U1308 (N_1308,N_1053,N_1081);
nand U1309 (N_1309,N_1143,N_1135);
nand U1310 (N_1310,N_1111,N_1068);
and U1311 (N_1311,N_1126,N_1090);
nor U1312 (N_1312,N_1176,N_1134);
or U1313 (N_1313,N_1020,N_1023);
or U1314 (N_1314,N_1028,N_1153);
or U1315 (N_1315,N_1014,N_1016);
or U1316 (N_1316,N_1135,N_1049);
and U1317 (N_1317,N_1176,N_1199);
nor U1318 (N_1318,N_1031,N_1082);
and U1319 (N_1319,N_1054,N_1159);
nor U1320 (N_1320,N_1170,N_1161);
or U1321 (N_1321,N_1138,N_1162);
or U1322 (N_1322,N_1134,N_1097);
and U1323 (N_1323,N_1072,N_1021);
and U1324 (N_1324,N_1134,N_1114);
nand U1325 (N_1325,N_1104,N_1167);
or U1326 (N_1326,N_1190,N_1016);
nor U1327 (N_1327,N_1078,N_1150);
or U1328 (N_1328,N_1169,N_1198);
nand U1329 (N_1329,N_1152,N_1097);
or U1330 (N_1330,N_1054,N_1032);
or U1331 (N_1331,N_1010,N_1155);
or U1332 (N_1332,N_1107,N_1197);
nand U1333 (N_1333,N_1027,N_1030);
nand U1334 (N_1334,N_1049,N_1088);
or U1335 (N_1335,N_1080,N_1034);
and U1336 (N_1336,N_1127,N_1051);
and U1337 (N_1337,N_1048,N_1047);
or U1338 (N_1338,N_1053,N_1120);
nor U1339 (N_1339,N_1191,N_1149);
nand U1340 (N_1340,N_1045,N_1070);
nor U1341 (N_1341,N_1114,N_1037);
nor U1342 (N_1342,N_1010,N_1126);
nor U1343 (N_1343,N_1093,N_1037);
and U1344 (N_1344,N_1162,N_1029);
and U1345 (N_1345,N_1075,N_1142);
and U1346 (N_1346,N_1088,N_1187);
nor U1347 (N_1347,N_1085,N_1096);
and U1348 (N_1348,N_1139,N_1157);
and U1349 (N_1349,N_1039,N_1118);
and U1350 (N_1350,N_1041,N_1073);
nand U1351 (N_1351,N_1091,N_1033);
or U1352 (N_1352,N_1102,N_1008);
nand U1353 (N_1353,N_1192,N_1032);
nand U1354 (N_1354,N_1110,N_1107);
nand U1355 (N_1355,N_1108,N_1005);
and U1356 (N_1356,N_1053,N_1109);
nand U1357 (N_1357,N_1165,N_1139);
nand U1358 (N_1358,N_1135,N_1141);
and U1359 (N_1359,N_1074,N_1034);
nor U1360 (N_1360,N_1065,N_1132);
and U1361 (N_1361,N_1130,N_1106);
nand U1362 (N_1362,N_1138,N_1128);
and U1363 (N_1363,N_1119,N_1186);
and U1364 (N_1364,N_1154,N_1033);
and U1365 (N_1365,N_1124,N_1122);
and U1366 (N_1366,N_1053,N_1186);
and U1367 (N_1367,N_1111,N_1161);
nand U1368 (N_1368,N_1002,N_1020);
or U1369 (N_1369,N_1036,N_1170);
xnor U1370 (N_1370,N_1157,N_1074);
nor U1371 (N_1371,N_1120,N_1143);
and U1372 (N_1372,N_1154,N_1080);
or U1373 (N_1373,N_1181,N_1113);
nor U1374 (N_1374,N_1184,N_1169);
nor U1375 (N_1375,N_1067,N_1019);
and U1376 (N_1376,N_1057,N_1032);
nand U1377 (N_1377,N_1136,N_1071);
nand U1378 (N_1378,N_1153,N_1001);
nor U1379 (N_1379,N_1118,N_1010);
nand U1380 (N_1380,N_1057,N_1078);
or U1381 (N_1381,N_1121,N_1024);
or U1382 (N_1382,N_1171,N_1016);
nor U1383 (N_1383,N_1073,N_1102);
nor U1384 (N_1384,N_1140,N_1138);
and U1385 (N_1385,N_1147,N_1086);
nand U1386 (N_1386,N_1103,N_1006);
nand U1387 (N_1387,N_1178,N_1037);
or U1388 (N_1388,N_1185,N_1175);
nor U1389 (N_1389,N_1034,N_1017);
nand U1390 (N_1390,N_1135,N_1170);
or U1391 (N_1391,N_1136,N_1070);
nor U1392 (N_1392,N_1165,N_1054);
nand U1393 (N_1393,N_1009,N_1044);
or U1394 (N_1394,N_1164,N_1092);
nand U1395 (N_1395,N_1021,N_1023);
or U1396 (N_1396,N_1197,N_1160);
xor U1397 (N_1397,N_1124,N_1079);
or U1398 (N_1398,N_1021,N_1174);
nand U1399 (N_1399,N_1053,N_1066);
and U1400 (N_1400,N_1388,N_1318);
nor U1401 (N_1401,N_1320,N_1272);
nor U1402 (N_1402,N_1246,N_1243);
or U1403 (N_1403,N_1264,N_1329);
and U1404 (N_1404,N_1295,N_1333);
nor U1405 (N_1405,N_1376,N_1286);
or U1406 (N_1406,N_1389,N_1213);
or U1407 (N_1407,N_1273,N_1350);
nand U1408 (N_1408,N_1316,N_1306);
nand U1409 (N_1409,N_1241,N_1381);
nand U1410 (N_1410,N_1282,N_1314);
nand U1411 (N_1411,N_1211,N_1308);
or U1412 (N_1412,N_1347,N_1330);
or U1413 (N_1413,N_1232,N_1359);
and U1414 (N_1414,N_1344,N_1210);
and U1415 (N_1415,N_1365,N_1342);
nor U1416 (N_1416,N_1363,N_1399);
nor U1417 (N_1417,N_1247,N_1361);
nor U1418 (N_1418,N_1251,N_1338);
nor U1419 (N_1419,N_1234,N_1343);
nor U1420 (N_1420,N_1367,N_1223);
nor U1421 (N_1421,N_1275,N_1335);
nand U1422 (N_1422,N_1301,N_1267);
nand U1423 (N_1423,N_1281,N_1229);
nor U1424 (N_1424,N_1356,N_1240);
nand U1425 (N_1425,N_1284,N_1204);
nor U1426 (N_1426,N_1292,N_1385);
or U1427 (N_1427,N_1212,N_1249);
or U1428 (N_1428,N_1315,N_1353);
nor U1429 (N_1429,N_1271,N_1391);
nand U1430 (N_1430,N_1220,N_1207);
and U1431 (N_1431,N_1341,N_1259);
nand U1432 (N_1432,N_1258,N_1305);
or U1433 (N_1433,N_1370,N_1339);
nor U1434 (N_1434,N_1224,N_1332);
nand U1435 (N_1435,N_1384,N_1307);
nand U1436 (N_1436,N_1269,N_1313);
nand U1437 (N_1437,N_1321,N_1225);
and U1438 (N_1438,N_1290,N_1252);
or U1439 (N_1439,N_1226,N_1334);
or U1440 (N_1440,N_1239,N_1379);
nand U1441 (N_1441,N_1377,N_1280);
and U1442 (N_1442,N_1257,N_1328);
and U1443 (N_1443,N_1380,N_1236);
nor U1444 (N_1444,N_1325,N_1289);
nand U1445 (N_1445,N_1358,N_1395);
or U1446 (N_1446,N_1299,N_1288);
nor U1447 (N_1447,N_1218,N_1340);
nor U1448 (N_1448,N_1302,N_1309);
nor U1449 (N_1449,N_1215,N_1250);
or U1450 (N_1450,N_1293,N_1312);
nand U1451 (N_1451,N_1245,N_1276);
xor U1452 (N_1452,N_1300,N_1235);
nor U1453 (N_1453,N_1255,N_1279);
nand U1454 (N_1454,N_1378,N_1383);
or U1455 (N_1455,N_1244,N_1230);
nand U1456 (N_1456,N_1387,N_1263);
nor U1457 (N_1457,N_1346,N_1202);
nor U1458 (N_1458,N_1216,N_1372);
or U1459 (N_1459,N_1262,N_1283);
or U1460 (N_1460,N_1374,N_1221);
nor U1461 (N_1461,N_1398,N_1364);
or U1462 (N_1462,N_1268,N_1352);
nand U1463 (N_1463,N_1233,N_1298);
nand U1464 (N_1464,N_1256,N_1254);
nor U1465 (N_1465,N_1237,N_1278);
and U1466 (N_1466,N_1354,N_1373);
nor U1467 (N_1467,N_1386,N_1362);
xnor U1468 (N_1468,N_1270,N_1253);
and U1469 (N_1469,N_1348,N_1206);
nor U1470 (N_1470,N_1324,N_1291);
and U1471 (N_1471,N_1277,N_1382);
or U1472 (N_1472,N_1397,N_1266);
nor U1473 (N_1473,N_1303,N_1227);
and U1474 (N_1474,N_1317,N_1238);
nand U1475 (N_1475,N_1296,N_1322);
nand U1476 (N_1476,N_1337,N_1208);
nand U1477 (N_1477,N_1274,N_1394);
nand U1478 (N_1478,N_1331,N_1345);
and U1479 (N_1479,N_1297,N_1393);
or U1480 (N_1480,N_1327,N_1336);
nor U1481 (N_1481,N_1323,N_1228);
and U1482 (N_1482,N_1390,N_1396);
nand U1483 (N_1483,N_1242,N_1349);
nor U1484 (N_1484,N_1214,N_1217);
and U1485 (N_1485,N_1294,N_1285);
nand U1486 (N_1486,N_1248,N_1222);
nand U1487 (N_1487,N_1368,N_1311);
and U1488 (N_1488,N_1231,N_1357);
nor U1489 (N_1489,N_1371,N_1310);
or U1490 (N_1490,N_1360,N_1205);
nor U1491 (N_1491,N_1375,N_1319);
or U1492 (N_1492,N_1261,N_1203);
nor U1493 (N_1493,N_1265,N_1355);
nand U1494 (N_1494,N_1260,N_1366);
and U1495 (N_1495,N_1219,N_1326);
or U1496 (N_1496,N_1369,N_1392);
and U1497 (N_1497,N_1287,N_1304);
nand U1498 (N_1498,N_1209,N_1201);
and U1499 (N_1499,N_1200,N_1351);
nand U1500 (N_1500,N_1280,N_1342);
nor U1501 (N_1501,N_1344,N_1367);
nand U1502 (N_1502,N_1384,N_1216);
nor U1503 (N_1503,N_1242,N_1384);
nand U1504 (N_1504,N_1225,N_1303);
nor U1505 (N_1505,N_1247,N_1383);
and U1506 (N_1506,N_1382,N_1218);
nor U1507 (N_1507,N_1365,N_1292);
nor U1508 (N_1508,N_1204,N_1237);
nand U1509 (N_1509,N_1225,N_1204);
and U1510 (N_1510,N_1368,N_1361);
and U1511 (N_1511,N_1338,N_1376);
and U1512 (N_1512,N_1284,N_1398);
or U1513 (N_1513,N_1318,N_1366);
and U1514 (N_1514,N_1368,N_1360);
or U1515 (N_1515,N_1297,N_1334);
nand U1516 (N_1516,N_1374,N_1238);
nor U1517 (N_1517,N_1397,N_1206);
and U1518 (N_1518,N_1299,N_1263);
or U1519 (N_1519,N_1285,N_1216);
nand U1520 (N_1520,N_1304,N_1385);
and U1521 (N_1521,N_1283,N_1393);
and U1522 (N_1522,N_1310,N_1395);
nand U1523 (N_1523,N_1396,N_1323);
nor U1524 (N_1524,N_1387,N_1314);
and U1525 (N_1525,N_1364,N_1336);
nor U1526 (N_1526,N_1334,N_1205);
and U1527 (N_1527,N_1284,N_1286);
nand U1528 (N_1528,N_1373,N_1340);
and U1529 (N_1529,N_1236,N_1204);
and U1530 (N_1530,N_1221,N_1338);
nand U1531 (N_1531,N_1211,N_1266);
nor U1532 (N_1532,N_1271,N_1308);
nand U1533 (N_1533,N_1253,N_1268);
nand U1534 (N_1534,N_1371,N_1288);
nand U1535 (N_1535,N_1202,N_1225);
or U1536 (N_1536,N_1243,N_1356);
nor U1537 (N_1537,N_1357,N_1230);
nand U1538 (N_1538,N_1224,N_1215);
nand U1539 (N_1539,N_1291,N_1252);
nand U1540 (N_1540,N_1399,N_1216);
and U1541 (N_1541,N_1249,N_1312);
and U1542 (N_1542,N_1298,N_1306);
nand U1543 (N_1543,N_1377,N_1327);
nand U1544 (N_1544,N_1384,N_1243);
nand U1545 (N_1545,N_1366,N_1212);
or U1546 (N_1546,N_1345,N_1285);
or U1547 (N_1547,N_1320,N_1235);
nand U1548 (N_1548,N_1339,N_1329);
or U1549 (N_1549,N_1256,N_1315);
nor U1550 (N_1550,N_1273,N_1388);
nor U1551 (N_1551,N_1207,N_1362);
or U1552 (N_1552,N_1204,N_1203);
nand U1553 (N_1553,N_1373,N_1206);
or U1554 (N_1554,N_1333,N_1353);
or U1555 (N_1555,N_1339,N_1380);
and U1556 (N_1556,N_1253,N_1243);
and U1557 (N_1557,N_1299,N_1306);
nand U1558 (N_1558,N_1304,N_1266);
nand U1559 (N_1559,N_1309,N_1246);
nand U1560 (N_1560,N_1369,N_1327);
xor U1561 (N_1561,N_1327,N_1332);
nand U1562 (N_1562,N_1322,N_1234);
or U1563 (N_1563,N_1215,N_1339);
and U1564 (N_1564,N_1217,N_1374);
nand U1565 (N_1565,N_1315,N_1302);
and U1566 (N_1566,N_1232,N_1374);
and U1567 (N_1567,N_1211,N_1203);
nand U1568 (N_1568,N_1220,N_1367);
or U1569 (N_1569,N_1210,N_1260);
or U1570 (N_1570,N_1268,N_1350);
xor U1571 (N_1571,N_1274,N_1377);
nand U1572 (N_1572,N_1229,N_1309);
nand U1573 (N_1573,N_1369,N_1207);
nand U1574 (N_1574,N_1219,N_1286);
or U1575 (N_1575,N_1259,N_1333);
nor U1576 (N_1576,N_1264,N_1231);
and U1577 (N_1577,N_1316,N_1272);
and U1578 (N_1578,N_1349,N_1246);
nor U1579 (N_1579,N_1247,N_1271);
and U1580 (N_1580,N_1344,N_1349);
or U1581 (N_1581,N_1359,N_1223);
or U1582 (N_1582,N_1385,N_1357);
and U1583 (N_1583,N_1362,N_1275);
and U1584 (N_1584,N_1273,N_1200);
xnor U1585 (N_1585,N_1264,N_1244);
or U1586 (N_1586,N_1266,N_1216);
nand U1587 (N_1587,N_1201,N_1317);
nand U1588 (N_1588,N_1377,N_1259);
and U1589 (N_1589,N_1280,N_1350);
nor U1590 (N_1590,N_1337,N_1281);
nor U1591 (N_1591,N_1324,N_1200);
nor U1592 (N_1592,N_1397,N_1383);
nor U1593 (N_1593,N_1283,N_1350);
and U1594 (N_1594,N_1386,N_1274);
nand U1595 (N_1595,N_1320,N_1269);
nand U1596 (N_1596,N_1312,N_1300);
nand U1597 (N_1597,N_1322,N_1282);
nand U1598 (N_1598,N_1296,N_1307);
or U1599 (N_1599,N_1307,N_1393);
and U1600 (N_1600,N_1418,N_1542);
or U1601 (N_1601,N_1583,N_1580);
and U1602 (N_1602,N_1473,N_1476);
nand U1603 (N_1603,N_1401,N_1484);
or U1604 (N_1604,N_1405,N_1422);
or U1605 (N_1605,N_1554,N_1563);
xor U1606 (N_1606,N_1426,N_1470);
nor U1607 (N_1607,N_1414,N_1407);
nand U1608 (N_1608,N_1423,N_1544);
and U1609 (N_1609,N_1424,N_1506);
nand U1610 (N_1610,N_1545,N_1460);
nand U1611 (N_1611,N_1540,N_1537);
and U1612 (N_1612,N_1565,N_1437);
or U1613 (N_1613,N_1570,N_1575);
nor U1614 (N_1614,N_1406,N_1450);
nor U1615 (N_1615,N_1562,N_1445);
xnor U1616 (N_1616,N_1592,N_1541);
nor U1617 (N_1617,N_1566,N_1453);
xor U1618 (N_1618,N_1515,N_1523);
nor U1619 (N_1619,N_1480,N_1493);
xor U1620 (N_1620,N_1502,N_1561);
and U1621 (N_1621,N_1411,N_1410);
nor U1622 (N_1622,N_1576,N_1485);
nand U1623 (N_1623,N_1428,N_1536);
xor U1624 (N_1624,N_1471,N_1546);
nor U1625 (N_1625,N_1577,N_1519);
nand U1626 (N_1626,N_1531,N_1511);
nand U1627 (N_1627,N_1400,N_1513);
and U1628 (N_1628,N_1558,N_1472);
or U1629 (N_1629,N_1538,N_1465);
xor U1630 (N_1630,N_1582,N_1527);
and U1631 (N_1631,N_1479,N_1594);
and U1632 (N_1632,N_1512,N_1522);
and U1633 (N_1633,N_1543,N_1595);
nand U1634 (N_1634,N_1573,N_1461);
or U1635 (N_1635,N_1477,N_1455);
nor U1636 (N_1636,N_1481,N_1514);
xnor U1637 (N_1637,N_1408,N_1579);
nand U1638 (N_1638,N_1596,N_1469);
and U1639 (N_1639,N_1413,N_1483);
xnor U1640 (N_1640,N_1448,N_1475);
or U1641 (N_1641,N_1505,N_1507);
nand U1642 (N_1642,N_1551,N_1462);
nor U1643 (N_1643,N_1417,N_1436);
nor U1644 (N_1644,N_1482,N_1593);
nand U1645 (N_1645,N_1499,N_1464);
nand U1646 (N_1646,N_1572,N_1509);
nand U1647 (N_1647,N_1520,N_1454);
nand U1648 (N_1648,N_1466,N_1404);
xor U1649 (N_1649,N_1571,N_1487);
or U1650 (N_1650,N_1447,N_1433);
or U1651 (N_1651,N_1589,N_1549);
or U1652 (N_1652,N_1456,N_1495);
or U1653 (N_1653,N_1432,N_1489);
nand U1654 (N_1654,N_1528,N_1496);
or U1655 (N_1655,N_1442,N_1510);
nor U1656 (N_1656,N_1567,N_1556);
and U1657 (N_1657,N_1458,N_1501);
nor U1658 (N_1658,N_1599,N_1584);
nand U1659 (N_1659,N_1498,N_1524);
xnor U1660 (N_1660,N_1439,N_1588);
nand U1661 (N_1661,N_1500,N_1597);
or U1662 (N_1662,N_1492,N_1463);
xor U1663 (N_1663,N_1503,N_1585);
nand U1664 (N_1664,N_1440,N_1434);
or U1665 (N_1665,N_1560,N_1488);
nand U1666 (N_1666,N_1449,N_1427);
and U1667 (N_1667,N_1415,N_1555);
and U1668 (N_1668,N_1581,N_1486);
nand U1669 (N_1669,N_1539,N_1429);
nand U1670 (N_1670,N_1552,N_1517);
nor U1671 (N_1671,N_1403,N_1430);
nor U1672 (N_1672,N_1553,N_1420);
or U1673 (N_1673,N_1508,N_1548);
xor U1674 (N_1674,N_1416,N_1452);
and U1675 (N_1675,N_1468,N_1533);
nand U1676 (N_1676,N_1518,N_1419);
nor U1677 (N_1677,N_1550,N_1474);
nor U1678 (N_1678,N_1591,N_1459);
or U1679 (N_1679,N_1421,N_1491);
xnor U1680 (N_1680,N_1504,N_1535);
nor U1681 (N_1681,N_1443,N_1587);
or U1682 (N_1682,N_1534,N_1559);
nor U1683 (N_1683,N_1497,N_1516);
nor U1684 (N_1684,N_1478,N_1402);
nor U1685 (N_1685,N_1425,N_1409);
or U1686 (N_1686,N_1564,N_1490);
and U1687 (N_1687,N_1438,N_1435);
and U1688 (N_1688,N_1525,N_1547);
nor U1689 (N_1689,N_1444,N_1451);
or U1690 (N_1690,N_1529,N_1569);
and U1691 (N_1691,N_1446,N_1598);
and U1692 (N_1692,N_1526,N_1441);
or U1693 (N_1693,N_1494,N_1578);
and U1694 (N_1694,N_1590,N_1532);
nand U1695 (N_1695,N_1557,N_1568);
nor U1696 (N_1696,N_1457,N_1521);
nor U1697 (N_1697,N_1530,N_1431);
nor U1698 (N_1698,N_1412,N_1467);
nand U1699 (N_1699,N_1574,N_1586);
nand U1700 (N_1700,N_1544,N_1551);
nand U1701 (N_1701,N_1579,N_1570);
nand U1702 (N_1702,N_1481,N_1549);
or U1703 (N_1703,N_1414,N_1456);
nor U1704 (N_1704,N_1581,N_1445);
and U1705 (N_1705,N_1568,N_1493);
nor U1706 (N_1706,N_1538,N_1487);
and U1707 (N_1707,N_1515,N_1447);
nand U1708 (N_1708,N_1498,N_1415);
nand U1709 (N_1709,N_1417,N_1484);
or U1710 (N_1710,N_1455,N_1447);
or U1711 (N_1711,N_1497,N_1425);
nor U1712 (N_1712,N_1559,N_1406);
nand U1713 (N_1713,N_1530,N_1439);
and U1714 (N_1714,N_1570,N_1513);
nand U1715 (N_1715,N_1418,N_1413);
nand U1716 (N_1716,N_1417,N_1576);
or U1717 (N_1717,N_1462,N_1464);
nor U1718 (N_1718,N_1435,N_1442);
nand U1719 (N_1719,N_1540,N_1409);
and U1720 (N_1720,N_1494,N_1591);
nor U1721 (N_1721,N_1546,N_1516);
nand U1722 (N_1722,N_1517,N_1589);
nor U1723 (N_1723,N_1454,N_1455);
nand U1724 (N_1724,N_1569,N_1554);
nand U1725 (N_1725,N_1516,N_1513);
or U1726 (N_1726,N_1507,N_1493);
or U1727 (N_1727,N_1432,N_1545);
or U1728 (N_1728,N_1423,N_1456);
and U1729 (N_1729,N_1496,N_1418);
and U1730 (N_1730,N_1449,N_1560);
and U1731 (N_1731,N_1465,N_1567);
nor U1732 (N_1732,N_1402,N_1403);
and U1733 (N_1733,N_1535,N_1486);
nand U1734 (N_1734,N_1471,N_1578);
nor U1735 (N_1735,N_1443,N_1467);
and U1736 (N_1736,N_1467,N_1414);
and U1737 (N_1737,N_1498,N_1581);
nand U1738 (N_1738,N_1466,N_1435);
nor U1739 (N_1739,N_1450,N_1588);
or U1740 (N_1740,N_1438,N_1507);
or U1741 (N_1741,N_1424,N_1522);
nor U1742 (N_1742,N_1426,N_1401);
or U1743 (N_1743,N_1567,N_1435);
nor U1744 (N_1744,N_1565,N_1564);
nor U1745 (N_1745,N_1444,N_1480);
nor U1746 (N_1746,N_1477,N_1561);
nand U1747 (N_1747,N_1499,N_1515);
or U1748 (N_1748,N_1495,N_1514);
xnor U1749 (N_1749,N_1447,N_1452);
nor U1750 (N_1750,N_1508,N_1463);
and U1751 (N_1751,N_1514,N_1419);
or U1752 (N_1752,N_1499,N_1420);
nor U1753 (N_1753,N_1588,N_1591);
and U1754 (N_1754,N_1595,N_1462);
nor U1755 (N_1755,N_1554,N_1573);
or U1756 (N_1756,N_1571,N_1527);
or U1757 (N_1757,N_1502,N_1509);
or U1758 (N_1758,N_1542,N_1487);
or U1759 (N_1759,N_1526,N_1452);
or U1760 (N_1760,N_1515,N_1507);
or U1761 (N_1761,N_1590,N_1569);
nand U1762 (N_1762,N_1457,N_1570);
nor U1763 (N_1763,N_1412,N_1432);
or U1764 (N_1764,N_1590,N_1478);
and U1765 (N_1765,N_1438,N_1570);
nor U1766 (N_1766,N_1476,N_1433);
or U1767 (N_1767,N_1435,N_1547);
xnor U1768 (N_1768,N_1441,N_1549);
xor U1769 (N_1769,N_1481,N_1413);
or U1770 (N_1770,N_1406,N_1426);
nand U1771 (N_1771,N_1500,N_1585);
or U1772 (N_1772,N_1563,N_1429);
nor U1773 (N_1773,N_1485,N_1422);
or U1774 (N_1774,N_1475,N_1584);
or U1775 (N_1775,N_1437,N_1406);
and U1776 (N_1776,N_1410,N_1552);
nand U1777 (N_1777,N_1578,N_1493);
and U1778 (N_1778,N_1450,N_1486);
nand U1779 (N_1779,N_1503,N_1476);
or U1780 (N_1780,N_1515,N_1417);
or U1781 (N_1781,N_1463,N_1409);
or U1782 (N_1782,N_1412,N_1443);
nor U1783 (N_1783,N_1495,N_1574);
or U1784 (N_1784,N_1448,N_1574);
nand U1785 (N_1785,N_1414,N_1501);
nor U1786 (N_1786,N_1449,N_1547);
and U1787 (N_1787,N_1471,N_1588);
or U1788 (N_1788,N_1466,N_1431);
or U1789 (N_1789,N_1405,N_1431);
and U1790 (N_1790,N_1501,N_1516);
or U1791 (N_1791,N_1524,N_1515);
nor U1792 (N_1792,N_1408,N_1450);
and U1793 (N_1793,N_1582,N_1409);
and U1794 (N_1794,N_1555,N_1529);
nor U1795 (N_1795,N_1408,N_1445);
nor U1796 (N_1796,N_1578,N_1536);
nand U1797 (N_1797,N_1409,N_1574);
and U1798 (N_1798,N_1597,N_1536);
nand U1799 (N_1799,N_1461,N_1578);
and U1800 (N_1800,N_1623,N_1621);
nand U1801 (N_1801,N_1778,N_1605);
and U1802 (N_1802,N_1782,N_1775);
nor U1803 (N_1803,N_1776,N_1793);
or U1804 (N_1804,N_1626,N_1644);
or U1805 (N_1805,N_1680,N_1692);
and U1806 (N_1806,N_1651,N_1766);
xor U1807 (N_1807,N_1697,N_1629);
or U1808 (N_1808,N_1601,N_1660);
or U1809 (N_1809,N_1722,N_1640);
nor U1810 (N_1810,N_1693,N_1764);
or U1811 (N_1811,N_1733,N_1795);
nand U1812 (N_1812,N_1649,N_1701);
and U1813 (N_1813,N_1689,N_1750);
or U1814 (N_1814,N_1740,N_1672);
nand U1815 (N_1815,N_1675,N_1661);
nand U1816 (N_1816,N_1785,N_1742);
or U1817 (N_1817,N_1737,N_1671);
or U1818 (N_1818,N_1657,N_1665);
nor U1819 (N_1819,N_1708,N_1602);
nor U1820 (N_1820,N_1687,N_1760);
or U1821 (N_1821,N_1631,N_1790);
or U1822 (N_1822,N_1768,N_1719);
or U1823 (N_1823,N_1705,N_1718);
or U1824 (N_1824,N_1736,N_1632);
nor U1825 (N_1825,N_1707,N_1646);
nand U1826 (N_1826,N_1659,N_1624);
and U1827 (N_1827,N_1636,N_1704);
or U1828 (N_1828,N_1769,N_1744);
and U1829 (N_1829,N_1630,N_1772);
or U1830 (N_1830,N_1754,N_1645);
and U1831 (N_1831,N_1668,N_1798);
and U1832 (N_1832,N_1603,N_1789);
nand U1833 (N_1833,N_1723,N_1677);
or U1834 (N_1834,N_1783,N_1741);
nor U1835 (N_1835,N_1779,N_1622);
or U1836 (N_1836,N_1690,N_1606);
or U1837 (N_1837,N_1788,N_1797);
or U1838 (N_1838,N_1669,N_1745);
or U1839 (N_1839,N_1676,N_1610);
nand U1840 (N_1840,N_1667,N_1673);
nand U1841 (N_1841,N_1647,N_1663);
nand U1842 (N_1842,N_1633,N_1721);
or U1843 (N_1843,N_1634,N_1729);
nor U1844 (N_1844,N_1739,N_1749);
nand U1845 (N_1845,N_1607,N_1696);
nand U1846 (N_1846,N_1714,N_1748);
or U1847 (N_1847,N_1648,N_1787);
nor U1848 (N_1848,N_1747,N_1699);
xnor U1849 (N_1849,N_1735,N_1796);
nor U1850 (N_1850,N_1717,N_1618);
xor U1851 (N_1851,N_1780,N_1670);
or U1852 (N_1852,N_1688,N_1734);
nand U1853 (N_1853,N_1738,N_1679);
nand U1854 (N_1854,N_1686,N_1619);
or U1855 (N_1855,N_1753,N_1724);
nand U1856 (N_1856,N_1639,N_1781);
or U1857 (N_1857,N_1643,N_1628);
nor U1858 (N_1858,N_1641,N_1691);
nor U1859 (N_1859,N_1774,N_1720);
nand U1860 (N_1860,N_1650,N_1759);
and U1861 (N_1861,N_1751,N_1617);
nor U1862 (N_1862,N_1730,N_1611);
nor U1863 (N_1863,N_1726,N_1608);
and U1864 (N_1864,N_1683,N_1609);
nor U1865 (N_1865,N_1711,N_1713);
nand U1866 (N_1866,N_1702,N_1755);
nor U1867 (N_1867,N_1706,N_1761);
nand U1868 (N_1868,N_1620,N_1627);
nand U1869 (N_1869,N_1625,N_1655);
or U1870 (N_1870,N_1616,N_1799);
nor U1871 (N_1871,N_1604,N_1715);
nor U1872 (N_1872,N_1638,N_1600);
nand U1873 (N_1873,N_1681,N_1700);
nor U1874 (N_1874,N_1770,N_1666);
and U1875 (N_1875,N_1727,N_1767);
nor U1876 (N_1876,N_1678,N_1695);
or U1877 (N_1877,N_1709,N_1682);
nand U1878 (N_1878,N_1757,N_1756);
or U1879 (N_1879,N_1712,N_1725);
or U1880 (N_1880,N_1664,N_1731);
and U1881 (N_1881,N_1612,N_1685);
xnor U1882 (N_1882,N_1656,N_1752);
xor U1883 (N_1883,N_1784,N_1732);
and U1884 (N_1884,N_1746,N_1716);
and U1885 (N_1885,N_1694,N_1614);
nand U1886 (N_1886,N_1652,N_1674);
nor U1887 (N_1887,N_1763,N_1777);
and U1888 (N_1888,N_1794,N_1743);
nand U1889 (N_1889,N_1773,N_1762);
nor U1890 (N_1890,N_1662,N_1653);
and U1891 (N_1891,N_1635,N_1703);
nor U1892 (N_1892,N_1684,N_1786);
nand U1893 (N_1893,N_1710,N_1771);
nand U1894 (N_1894,N_1765,N_1728);
nor U1895 (N_1895,N_1698,N_1758);
nand U1896 (N_1896,N_1613,N_1791);
nand U1897 (N_1897,N_1642,N_1658);
nor U1898 (N_1898,N_1615,N_1654);
and U1899 (N_1899,N_1637,N_1792);
xor U1900 (N_1900,N_1676,N_1658);
nor U1901 (N_1901,N_1638,N_1668);
and U1902 (N_1902,N_1630,N_1667);
or U1903 (N_1903,N_1605,N_1675);
nor U1904 (N_1904,N_1686,N_1707);
or U1905 (N_1905,N_1623,N_1673);
nand U1906 (N_1906,N_1745,N_1643);
and U1907 (N_1907,N_1799,N_1774);
nor U1908 (N_1908,N_1776,N_1791);
nand U1909 (N_1909,N_1751,N_1636);
xnor U1910 (N_1910,N_1798,N_1671);
nor U1911 (N_1911,N_1713,N_1765);
and U1912 (N_1912,N_1711,N_1686);
nor U1913 (N_1913,N_1734,N_1723);
nor U1914 (N_1914,N_1633,N_1671);
nor U1915 (N_1915,N_1660,N_1608);
or U1916 (N_1916,N_1749,N_1725);
nor U1917 (N_1917,N_1793,N_1720);
nor U1918 (N_1918,N_1747,N_1701);
and U1919 (N_1919,N_1667,N_1602);
nand U1920 (N_1920,N_1662,N_1611);
or U1921 (N_1921,N_1726,N_1796);
nor U1922 (N_1922,N_1727,N_1625);
and U1923 (N_1923,N_1603,N_1725);
or U1924 (N_1924,N_1741,N_1716);
or U1925 (N_1925,N_1698,N_1606);
nand U1926 (N_1926,N_1613,N_1699);
nand U1927 (N_1927,N_1753,N_1751);
or U1928 (N_1928,N_1636,N_1743);
or U1929 (N_1929,N_1746,N_1713);
or U1930 (N_1930,N_1772,N_1737);
and U1931 (N_1931,N_1672,N_1690);
xnor U1932 (N_1932,N_1673,N_1759);
or U1933 (N_1933,N_1720,N_1627);
nor U1934 (N_1934,N_1698,N_1795);
nand U1935 (N_1935,N_1750,N_1757);
nor U1936 (N_1936,N_1682,N_1773);
and U1937 (N_1937,N_1603,N_1694);
and U1938 (N_1938,N_1726,N_1724);
nand U1939 (N_1939,N_1754,N_1760);
and U1940 (N_1940,N_1729,N_1797);
nand U1941 (N_1941,N_1779,N_1743);
nor U1942 (N_1942,N_1675,N_1651);
nor U1943 (N_1943,N_1627,N_1634);
nor U1944 (N_1944,N_1687,N_1650);
or U1945 (N_1945,N_1627,N_1754);
or U1946 (N_1946,N_1620,N_1668);
and U1947 (N_1947,N_1693,N_1688);
and U1948 (N_1948,N_1603,N_1760);
nor U1949 (N_1949,N_1677,N_1661);
or U1950 (N_1950,N_1689,N_1657);
and U1951 (N_1951,N_1709,N_1630);
and U1952 (N_1952,N_1640,N_1600);
or U1953 (N_1953,N_1648,N_1765);
nor U1954 (N_1954,N_1694,N_1602);
nor U1955 (N_1955,N_1694,N_1648);
nor U1956 (N_1956,N_1638,N_1608);
and U1957 (N_1957,N_1731,N_1694);
nor U1958 (N_1958,N_1731,N_1750);
and U1959 (N_1959,N_1728,N_1734);
and U1960 (N_1960,N_1650,N_1696);
and U1961 (N_1961,N_1739,N_1742);
nand U1962 (N_1962,N_1627,N_1692);
or U1963 (N_1963,N_1601,N_1637);
nor U1964 (N_1964,N_1691,N_1639);
or U1965 (N_1965,N_1738,N_1697);
and U1966 (N_1966,N_1625,N_1677);
nor U1967 (N_1967,N_1707,N_1785);
or U1968 (N_1968,N_1771,N_1614);
and U1969 (N_1969,N_1681,N_1632);
and U1970 (N_1970,N_1689,N_1625);
or U1971 (N_1971,N_1616,N_1746);
nand U1972 (N_1972,N_1635,N_1763);
or U1973 (N_1973,N_1698,N_1694);
and U1974 (N_1974,N_1769,N_1658);
nor U1975 (N_1975,N_1692,N_1735);
nor U1976 (N_1976,N_1688,N_1673);
nand U1977 (N_1977,N_1725,N_1655);
nand U1978 (N_1978,N_1741,N_1738);
nor U1979 (N_1979,N_1681,N_1747);
nor U1980 (N_1980,N_1669,N_1767);
or U1981 (N_1981,N_1774,N_1662);
and U1982 (N_1982,N_1606,N_1611);
or U1983 (N_1983,N_1664,N_1665);
or U1984 (N_1984,N_1712,N_1763);
nor U1985 (N_1985,N_1795,N_1796);
nand U1986 (N_1986,N_1654,N_1758);
nor U1987 (N_1987,N_1722,N_1751);
or U1988 (N_1988,N_1733,N_1601);
nand U1989 (N_1989,N_1778,N_1701);
or U1990 (N_1990,N_1697,N_1657);
or U1991 (N_1991,N_1711,N_1793);
or U1992 (N_1992,N_1691,N_1631);
nand U1993 (N_1993,N_1765,N_1684);
nor U1994 (N_1994,N_1675,N_1780);
nor U1995 (N_1995,N_1603,N_1771);
and U1996 (N_1996,N_1623,N_1750);
nor U1997 (N_1997,N_1779,N_1655);
and U1998 (N_1998,N_1614,N_1721);
or U1999 (N_1999,N_1615,N_1695);
nand U2000 (N_2000,N_1905,N_1928);
or U2001 (N_2001,N_1961,N_1889);
nand U2002 (N_2002,N_1955,N_1996);
nor U2003 (N_2003,N_1865,N_1985);
nor U2004 (N_2004,N_1898,N_1845);
and U2005 (N_2005,N_1976,N_1967);
and U2006 (N_2006,N_1969,N_1988);
nand U2007 (N_2007,N_1904,N_1948);
or U2008 (N_2008,N_1916,N_1930);
nand U2009 (N_2009,N_1949,N_1841);
nor U2010 (N_2010,N_1920,N_1887);
nor U2011 (N_2011,N_1844,N_1881);
and U2012 (N_2012,N_1848,N_1859);
nor U2013 (N_2013,N_1831,N_1863);
nor U2014 (N_2014,N_1899,N_1915);
or U2015 (N_2015,N_1924,N_1903);
or U2016 (N_2016,N_1897,N_1980);
or U2017 (N_2017,N_1836,N_1989);
and U2018 (N_2018,N_1882,N_1921);
xor U2019 (N_2019,N_1927,N_1929);
or U2020 (N_2020,N_1872,N_1869);
or U2021 (N_2021,N_1926,N_1805);
and U2022 (N_2022,N_1829,N_1974);
and U2023 (N_2023,N_1938,N_1819);
nor U2024 (N_2024,N_1942,N_1971);
or U2025 (N_2025,N_1876,N_1995);
nand U2026 (N_2026,N_1802,N_1817);
and U2027 (N_2027,N_1963,N_1934);
or U2028 (N_2028,N_1851,N_1807);
nor U2029 (N_2029,N_1827,N_1983);
or U2030 (N_2030,N_1909,N_1809);
or U2031 (N_2031,N_1861,N_1939);
xnor U2032 (N_2032,N_1896,N_1830);
or U2033 (N_2033,N_1981,N_1825);
and U2034 (N_2034,N_1853,N_1879);
or U2035 (N_2035,N_1864,N_1925);
and U2036 (N_2036,N_1834,N_1990);
and U2037 (N_2037,N_1975,N_1919);
xor U2038 (N_2038,N_1945,N_1936);
nand U2039 (N_2039,N_1801,N_1873);
nor U2040 (N_2040,N_1843,N_1890);
nand U2041 (N_2041,N_1842,N_1857);
nand U2042 (N_2042,N_1866,N_1913);
or U2043 (N_2043,N_1892,N_1947);
or U2044 (N_2044,N_1855,N_1914);
or U2045 (N_2045,N_1858,N_1912);
or U2046 (N_2046,N_1822,N_1895);
and U2047 (N_2047,N_1838,N_1960);
nand U2048 (N_2048,N_1806,N_1986);
nor U2049 (N_2049,N_1810,N_1815);
nand U2050 (N_2050,N_1957,N_1972);
or U2051 (N_2051,N_1835,N_1824);
nand U2052 (N_2052,N_1893,N_1943);
nand U2053 (N_2053,N_1908,N_1870);
nor U2054 (N_2054,N_1868,N_1901);
or U2055 (N_2055,N_1918,N_1952);
and U2056 (N_2056,N_1966,N_1977);
or U2057 (N_2057,N_1852,N_1854);
or U2058 (N_2058,N_1837,N_1997);
or U2059 (N_2059,N_1820,N_1877);
or U2060 (N_2060,N_1956,N_1811);
and U2061 (N_2061,N_1946,N_1911);
nand U2062 (N_2062,N_1880,N_1856);
xnor U2063 (N_2063,N_1833,N_1964);
and U2064 (N_2064,N_1816,N_1821);
or U2065 (N_2065,N_1917,N_1944);
nand U2066 (N_2066,N_1803,N_1999);
nor U2067 (N_2067,N_1954,N_1888);
and U2068 (N_2068,N_1878,N_1839);
or U2069 (N_2069,N_1940,N_1849);
nor U2070 (N_2070,N_1818,N_1958);
and U2071 (N_2071,N_1937,N_1832);
nor U2072 (N_2072,N_1907,N_1970);
nor U2073 (N_2073,N_1850,N_1840);
xor U2074 (N_2074,N_1987,N_1900);
nand U2075 (N_2075,N_1935,N_1933);
nand U2076 (N_2076,N_1826,N_1808);
nor U2077 (N_2077,N_1968,N_1922);
or U2078 (N_2078,N_1886,N_1979);
nand U2079 (N_2079,N_1847,N_1804);
nor U2080 (N_2080,N_1800,N_1871);
and U2081 (N_2081,N_1931,N_1894);
and U2082 (N_2082,N_1973,N_1951);
nand U2083 (N_2083,N_1813,N_1884);
and U2084 (N_2084,N_1910,N_1953);
or U2085 (N_2085,N_1965,N_1994);
or U2086 (N_2086,N_1814,N_1862);
nor U2087 (N_2087,N_1950,N_1984);
or U2088 (N_2088,N_1923,N_1823);
nor U2089 (N_2089,N_1906,N_1860);
nor U2090 (N_2090,N_1941,N_1812);
or U2091 (N_2091,N_1883,N_1932);
or U2092 (N_2092,N_1885,N_1959);
nor U2093 (N_2093,N_1998,N_1874);
or U2094 (N_2094,N_1891,N_1828);
nand U2095 (N_2095,N_1993,N_1902);
or U2096 (N_2096,N_1982,N_1962);
and U2097 (N_2097,N_1846,N_1875);
nor U2098 (N_2098,N_1867,N_1992);
or U2099 (N_2099,N_1978,N_1991);
nor U2100 (N_2100,N_1906,N_1896);
nor U2101 (N_2101,N_1986,N_1982);
nand U2102 (N_2102,N_1820,N_1821);
and U2103 (N_2103,N_1992,N_1925);
nand U2104 (N_2104,N_1894,N_1972);
nor U2105 (N_2105,N_1989,N_1819);
nor U2106 (N_2106,N_1954,N_1971);
or U2107 (N_2107,N_1892,N_1979);
nor U2108 (N_2108,N_1888,N_1834);
nand U2109 (N_2109,N_1980,N_1931);
nand U2110 (N_2110,N_1808,N_1903);
and U2111 (N_2111,N_1907,N_1813);
nor U2112 (N_2112,N_1860,N_1821);
nand U2113 (N_2113,N_1889,N_1845);
and U2114 (N_2114,N_1964,N_1984);
nand U2115 (N_2115,N_1978,N_1990);
and U2116 (N_2116,N_1853,N_1922);
or U2117 (N_2117,N_1881,N_1974);
nor U2118 (N_2118,N_1913,N_1912);
nand U2119 (N_2119,N_1895,N_1877);
and U2120 (N_2120,N_1893,N_1835);
nand U2121 (N_2121,N_1904,N_1833);
or U2122 (N_2122,N_1856,N_1822);
nor U2123 (N_2123,N_1831,N_1950);
or U2124 (N_2124,N_1957,N_1941);
or U2125 (N_2125,N_1830,N_1952);
and U2126 (N_2126,N_1923,N_1969);
and U2127 (N_2127,N_1969,N_1889);
and U2128 (N_2128,N_1884,N_1989);
nor U2129 (N_2129,N_1897,N_1852);
nor U2130 (N_2130,N_1929,N_1841);
and U2131 (N_2131,N_1995,N_1971);
and U2132 (N_2132,N_1881,N_1804);
nor U2133 (N_2133,N_1993,N_1962);
and U2134 (N_2134,N_1912,N_1840);
or U2135 (N_2135,N_1859,N_1971);
or U2136 (N_2136,N_1930,N_1821);
nand U2137 (N_2137,N_1992,N_1940);
or U2138 (N_2138,N_1850,N_1887);
nand U2139 (N_2139,N_1938,N_1914);
nor U2140 (N_2140,N_1976,N_1853);
nor U2141 (N_2141,N_1806,N_1834);
or U2142 (N_2142,N_1901,N_1986);
or U2143 (N_2143,N_1842,N_1986);
or U2144 (N_2144,N_1932,N_1880);
and U2145 (N_2145,N_1986,N_1925);
or U2146 (N_2146,N_1848,N_1997);
nor U2147 (N_2147,N_1801,N_1811);
nor U2148 (N_2148,N_1989,N_1953);
nor U2149 (N_2149,N_1867,N_1903);
nand U2150 (N_2150,N_1911,N_1921);
or U2151 (N_2151,N_1877,N_1835);
xnor U2152 (N_2152,N_1889,N_1852);
xnor U2153 (N_2153,N_1899,N_1895);
or U2154 (N_2154,N_1827,N_1931);
nand U2155 (N_2155,N_1948,N_1954);
nor U2156 (N_2156,N_1914,N_1869);
or U2157 (N_2157,N_1924,N_1809);
or U2158 (N_2158,N_1995,N_1889);
or U2159 (N_2159,N_1973,N_1920);
or U2160 (N_2160,N_1945,N_1847);
and U2161 (N_2161,N_1820,N_1991);
nand U2162 (N_2162,N_1899,N_1844);
or U2163 (N_2163,N_1870,N_1854);
or U2164 (N_2164,N_1855,N_1959);
and U2165 (N_2165,N_1919,N_1992);
and U2166 (N_2166,N_1877,N_1920);
nor U2167 (N_2167,N_1985,N_1921);
nor U2168 (N_2168,N_1944,N_1860);
nor U2169 (N_2169,N_1896,N_1840);
or U2170 (N_2170,N_1802,N_1928);
or U2171 (N_2171,N_1873,N_1851);
and U2172 (N_2172,N_1908,N_1868);
or U2173 (N_2173,N_1917,N_1847);
nand U2174 (N_2174,N_1966,N_1888);
and U2175 (N_2175,N_1865,N_1861);
or U2176 (N_2176,N_1940,N_1853);
and U2177 (N_2177,N_1958,N_1832);
and U2178 (N_2178,N_1958,N_1836);
and U2179 (N_2179,N_1846,N_1889);
nor U2180 (N_2180,N_1975,N_1903);
and U2181 (N_2181,N_1871,N_1980);
nand U2182 (N_2182,N_1866,N_1853);
xor U2183 (N_2183,N_1821,N_1810);
and U2184 (N_2184,N_1890,N_1939);
nor U2185 (N_2185,N_1956,N_1862);
nand U2186 (N_2186,N_1952,N_1915);
nor U2187 (N_2187,N_1952,N_1910);
nor U2188 (N_2188,N_1970,N_1877);
or U2189 (N_2189,N_1986,N_1941);
nand U2190 (N_2190,N_1942,N_1841);
nand U2191 (N_2191,N_1802,N_1996);
or U2192 (N_2192,N_1922,N_1948);
xor U2193 (N_2193,N_1844,N_1938);
or U2194 (N_2194,N_1999,N_1996);
or U2195 (N_2195,N_1910,N_1827);
and U2196 (N_2196,N_1965,N_1916);
or U2197 (N_2197,N_1895,N_1982);
or U2198 (N_2198,N_1884,N_1950);
nor U2199 (N_2199,N_1806,N_1815);
nor U2200 (N_2200,N_2095,N_2008);
nor U2201 (N_2201,N_2066,N_2121);
xor U2202 (N_2202,N_2043,N_2104);
nor U2203 (N_2203,N_2153,N_2054);
xor U2204 (N_2204,N_2186,N_2004);
nor U2205 (N_2205,N_2035,N_2116);
or U2206 (N_2206,N_2126,N_2156);
nor U2207 (N_2207,N_2003,N_2030);
nand U2208 (N_2208,N_2047,N_2110);
xor U2209 (N_2209,N_2005,N_2185);
or U2210 (N_2210,N_2197,N_2036);
or U2211 (N_2211,N_2042,N_2015);
and U2212 (N_2212,N_2044,N_2103);
nand U2213 (N_2213,N_2049,N_2175);
nor U2214 (N_2214,N_2006,N_2134);
nand U2215 (N_2215,N_2083,N_2196);
and U2216 (N_2216,N_2070,N_2100);
or U2217 (N_2217,N_2016,N_2065);
nor U2218 (N_2218,N_2188,N_2084);
and U2219 (N_2219,N_2141,N_2086);
or U2220 (N_2220,N_2020,N_2027);
and U2221 (N_2221,N_2055,N_2187);
nor U2222 (N_2222,N_2058,N_2085);
or U2223 (N_2223,N_2099,N_2052);
or U2224 (N_2224,N_2023,N_2146);
nor U2225 (N_2225,N_2076,N_2077);
nor U2226 (N_2226,N_2041,N_2031);
and U2227 (N_2227,N_2078,N_2170);
nor U2228 (N_2228,N_2046,N_2051);
nand U2229 (N_2229,N_2140,N_2122);
or U2230 (N_2230,N_2081,N_2133);
nor U2231 (N_2231,N_2087,N_2168);
and U2232 (N_2232,N_2163,N_2117);
nand U2233 (N_2233,N_2011,N_2136);
xnor U2234 (N_2234,N_2181,N_2067);
or U2235 (N_2235,N_2106,N_2165);
nor U2236 (N_2236,N_2190,N_2022);
or U2237 (N_2237,N_2164,N_2032);
xnor U2238 (N_2238,N_2040,N_2069);
nor U2239 (N_2239,N_2137,N_2152);
nor U2240 (N_2240,N_2151,N_2159);
nand U2241 (N_2241,N_2193,N_2033);
nor U2242 (N_2242,N_2108,N_2111);
nor U2243 (N_2243,N_2002,N_2098);
nor U2244 (N_2244,N_2123,N_2142);
nor U2245 (N_2245,N_2192,N_2092);
nor U2246 (N_2246,N_2180,N_2045);
nand U2247 (N_2247,N_2102,N_2009);
and U2248 (N_2248,N_2174,N_2028);
or U2249 (N_2249,N_2183,N_2158);
xor U2250 (N_2250,N_2177,N_2178);
nand U2251 (N_2251,N_2073,N_2029);
or U2252 (N_2252,N_2112,N_2176);
nor U2253 (N_2253,N_2072,N_2160);
and U2254 (N_2254,N_2089,N_2129);
nor U2255 (N_2255,N_2101,N_2144);
nor U2256 (N_2256,N_2161,N_2063);
nand U2257 (N_2257,N_2056,N_2132);
and U2258 (N_2258,N_2019,N_2050);
and U2259 (N_2259,N_2057,N_2012);
or U2260 (N_2260,N_2039,N_2115);
nand U2261 (N_2261,N_2082,N_2167);
nor U2262 (N_2262,N_2071,N_2088);
nor U2263 (N_2263,N_2091,N_2169);
nor U2264 (N_2264,N_2097,N_2128);
or U2265 (N_2265,N_2109,N_2155);
or U2266 (N_2266,N_2162,N_2172);
nor U2267 (N_2267,N_2173,N_2107);
nor U2268 (N_2268,N_2191,N_2124);
nor U2269 (N_2269,N_2120,N_2079);
or U2270 (N_2270,N_2113,N_2138);
and U2271 (N_2271,N_2189,N_2148);
or U2272 (N_2272,N_2135,N_2038);
or U2273 (N_2273,N_2171,N_2096);
nand U2274 (N_2274,N_2025,N_2194);
and U2275 (N_2275,N_2064,N_2127);
nand U2276 (N_2276,N_2053,N_2198);
and U2277 (N_2277,N_2018,N_2010);
nand U2278 (N_2278,N_2149,N_2150);
nor U2279 (N_2279,N_2000,N_2017);
and U2280 (N_2280,N_2059,N_2094);
nor U2281 (N_2281,N_2130,N_2139);
nor U2282 (N_2282,N_2037,N_2074);
nor U2283 (N_2283,N_2034,N_2199);
nand U2284 (N_2284,N_2060,N_2001);
xor U2285 (N_2285,N_2125,N_2090);
or U2286 (N_2286,N_2182,N_2119);
nor U2287 (N_2287,N_2154,N_2179);
nor U2288 (N_2288,N_2007,N_2195);
and U2289 (N_2289,N_2157,N_2131);
nor U2290 (N_2290,N_2024,N_2143);
nand U2291 (N_2291,N_2145,N_2068);
xor U2292 (N_2292,N_2061,N_2062);
nor U2293 (N_2293,N_2105,N_2013);
and U2294 (N_2294,N_2093,N_2114);
and U2295 (N_2295,N_2075,N_2048);
nand U2296 (N_2296,N_2147,N_2026);
nor U2297 (N_2297,N_2014,N_2166);
nor U2298 (N_2298,N_2184,N_2021);
nor U2299 (N_2299,N_2118,N_2080);
nor U2300 (N_2300,N_2055,N_2135);
and U2301 (N_2301,N_2036,N_2177);
and U2302 (N_2302,N_2162,N_2027);
or U2303 (N_2303,N_2055,N_2107);
nand U2304 (N_2304,N_2027,N_2131);
nor U2305 (N_2305,N_2141,N_2067);
nor U2306 (N_2306,N_2167,N_2033);
and U2307 (N_2307,N_2036,N_2077);
nand U2308 (N_2308,N_2010,N_2089);
and U2309 (N_2309,N_2041,N_2157);
or U2310 (N_2310,N_2115,N_2107);
or U2311 (N_2311,N_2165,N_2095);
and U2312 (N_2312,N_2191,N_2163);
or U2313 (N_2313,N_2027,N_2090);
nor U2314 (N_2314,N_2156,N_2115);
or U2315 (N_2315,N_2147,N_2152);
nand U2316 (N_2316,N_2116,N_2065);
nand U2317 (N_2317,N_2115,N_2040);
and U2318 (N_2318,N_2077,N_2084);
and U2319 (N_2319,N_2179,N_2086);
or U2320 (N_2320,N_2171,N_2095);
and U2321 (N_2321,N_2149,N_2058);
nand U2322 (N_2322,N_2146,N_2009);
or U2323 (N_2323,N_2115,N_2103);
and U2324 (N_2324,N_2132,N_2118);
nor U2325 (N_2325,N_2008,N_2188);
or U2326 (N_2326,N_2179,N_2003);
or U2327 (N_2327,N_2064,N_2034);
nand U2328 (N_2328,N_2074,N_2129);
or U2329 (N_2329,N_2105,N_2003);
or U2330 (N_2330,N_2081,N_2183);
and U2331 (N_2331,N_2017,N_2026);
nor U2332 (N_2332,N_2007,N_2043);
nor U2333 (N_2333,N_2055,N_2060);
nand U2334 (N_2334,N_2115,N_2155);
or U2335 (N_2335,N_2116,N_2043);
and U2336 (N_2336,N_2023,N_2162);
and U2337 (N_2337,N_2112,N_2196);
or U2338 (N_2338,N_2171,N_2164);
and U2339 (N_2339,N_2025,N_2034);
or U2340 (N_2340,N_2137,N_2180);
nor U2341 (N_2341,N_2064,N_2097);
and U2342 (N_2342,N_2001,N_2151);
nand U2343 (N_2343,N_2064,N_2071);
nand U2344 (N_2344,N_2112,N_2197);
and U2345 (N_2345,N_2077,N_2061);
nor U2346 (N_2346,N_2173,N_2191);
and U2347 (N_2347,N_2043,N_2108);
or U2348 (N_2348,N_2176,N_2113);
and U2349 (N_2349,N_2037,N_2068);
nor U2350 (N_2350,N_2172,N_2179);
and U2351 (N_2351,N_2012,N_2076);
nand U2352 (N_2352,N_2122,N_2074);
nand U2353 (N_2353,N_2163,N_2044);
nand U2354 (N_2354,N_2078,N_2126);
nor U2355 (N_2355,N_2058,N_2146);
and U2356 (N_2356,N_2141,N_2156);
and U2357 (N_2357,N_2199,N_2187);
and U2358 (N_2358,N_2036,N_2168);
nor U2359 (N_2359,N_2107,N_2010);
or U2360 (N_2360,N_2162,N_2160);
or U2361 (N_2361,N_2107,N_2194);
nor U2362 (N_2362,N_2116,N_2192);
or U2363 (N_2363,N_2188,N_2187);
nand U2364 (N_2364,N_2006,N_2107);
and U2365 (N_2365,N_2193,N_2148);
or U2366 (N_2366,N_2142,N_2126);
or U2367 (N_2367,N_2029,N_2099);
nor U2368 (N_2368,N_2121,N_2159);
and U2369 (N_2369,N_2190,N_2132);
or U2370 (N_2370,N_2118,N_2116);
or U2371 (N_2371,N_2028,N_2088);
xor U2372 (N_2372,N_2154,N_2138);
nand U2373 (N_2373,N_2015,N_2154);
nor U2374 (N_2374,N_2031,N_2037);
nor U2375 (N_2375,N_2058,N_2176);
nor U2376 (N_2376,N_2050,N_2070);
nor U2377 (N_2377,N_2017,N_2130);
and U2378 (N_2378,N_2133,N_2073);
and U2379 (N_2379,N_2152,N_2176);
nand U2380 (N_2380,N_2109,N_2191);
nand U2381 (N_2381,N_2007,N_2129);
nor U2382 (N_2382,N_2171,N_2034);
and U2383 (N_2383,N_2163,N_2134);
or U2384 (N_2384,N_2067,N_2017);
and U2385 (N_2385,N_2046,N_2091);
and U2386 (N_2386,N_2060,N_2183);
and U2387 (N_2387,N_2011,N_2147);
nor U2388 (N_2388,N_2074,N_2048);
nor U2389 (N_2389,N_2180,N_2143);
and U2390 (N_2390,N_2038,N_2021);
and U2391 (N_2391,N_2061,N_2167);
and U2392 (N_2392,N_2001,N_2156);
and U2393 (N_2393,N_2071,N_2023);
or U2394 (N_2394,N_2106,N_2075);
or U2395 (N_2395,N_2015,N_2103);
or U2396 (N_2396,N_2119,N_2076);
nand U2397 (N_2397,N_2051,N_2013);
and U2398 (N_2398,N_2008,N_2158);
and U2399 (N_2399,N_2037,N_2139);
nor U2400 (N_2400,N_2342,N_2394);
nand U2401 (N_2401,N_2332,N_2236);
or U2402 (N_2402,N_2320,N_2358);
and U2403 (N_2403,N_2334,N_2223);
nand U2404 (N_2404,N_2323,N_2273);
or U2405 (N_2405,N_2248,N_2216);
nor U2406 (N_2406,N_2286,N_2207);
or U2407 (N_2407,N_2372,N_2232);
or U2408 (N_2408,N_2234,N_2349);
and U2409 (N_2409,N_2222,N_2264);
and U2410 (N_2410,N_2270,N_2231);
and U2411 (N_2411,N_2239,N_2240);
or U2412 (N_2412,N_2296,N_2322);
xor U2413 (N_2413,N_2289,N_2250);
or U2414 (N_2414,N_2368,N_2283);
nor U2415 (N_2415,N_2374,N_2268);
nand U2416 (N_2416,N_2346,N_2399);
or U2417 (N_2417,N_2365,N_2330);
and U2418 (N_2418,N_2241,N_2350);
and U2419 (N_2419,N_2314,N_2307);
nand U2420 (N_2420,N_2274,N_2335);
nand U2421 (N_2421,N_2254,N_2381);
or U2422 (N_2422,N_2285,N_2306);
or U2423 (N_2423,N_2391,N_2353);
nand U2424 (N_2424,N_2218,N_2300);
nor U2425 (N_2425,N_2352,N_2347);
nand U2426 (N_2426,N_2356,N_2235);
nand U2427 (N_2427,N_2221,N_2313);
nor U2428 (N_2428,N_2384,N_2291);
nor U2429 (N_2429,N_2263,N_2355);
nor U2430 (N_2430,N_2382,N_2380);
nor U2431 (N_2431,N_2233,N_2398);
nand U2432 (N_2432,N_2348,N_2371);
nor U2433 (N_2433,N_2298,N_2258);
nor U2434 (N_2434,N_2267,N_2249);
nand U2435 (N_2435,N_2311,N_2279);
nand U2436 (N_2436,N_2272,N_2308);
nand U2437 (N_2437,N_2376,N_2345);
nand U2438 (N_2438,N_2359,N_2315);
xnor U2439 (N_2439,N_2328,N_2238);
and U2440 (N_2440,N_2393,N_2357);
nor U2441 (N_2441,N_2369,N_2303);
or U2442 (N_2442,N_2282,N_2287);
nor U2443 (N_2443,N_2225,N_2210);
nor U2444 (N_2444,N_2310,N_2378);
and U2445 (N_2445,N_2229,N_2230);
nand U2446 (N_2446,N_2251,N_2265);
or U2447 (N_2447,N_2226,N_2275);
or U2448 (N_2448,N_2209,N_2375);
nor U2449 (N_2449,N_2325,N_2312);
or U2450 (N_2450,N_2329,N_2338);
nor U2451 (N_2451,N_2200,N_2284);
or U2452 (N_2452,N_2259,N_2295);
nand U2453 (N_2453,N_2260,N_2321);
nand U2454 (N_2454,N_2363,N_2302);
nor U2455 (N_2455,N_2361,N_2253);
or U2456 (N_2456,N_2214,N_2219);
or U2457 (N_2457,N_2336,N_2280);
and U2458 (N_2458,N_2388,N_2318);
nor U2459 (N_2459,N_2213,N_2206);
nand U2460 (N_2460,N_2304,N_2212);
nand U2461 (N_2461,N_2331,N_2324);
nor U2462 (N_2462,N_2337,N_2217);
nor U2463 (N_2463,N_2370,N_2367);
nor U2464 (N_2464,N_2228,N_2255);
and U2465 (N_2465,N_2262,N_2392);
nor U2466 (N_2466,N_2341,N_2354);
or U2467 (N_2467,N_2243,N_2379);
nor U2468 (N_2468,N_2340,N_2339);
xor U2469 (N_2469,N_2397,N_2386);
and U2470 (N_2470,N_2377,N_2290);
nor U2471 (N_2471,N_2294,N_2364);
nand U2472 (N_2472,N_2333,N_2395);
nor U2473 (N_2473,N_2373,N_2389);
nor U2474 (N_2474,N_2256,N_2396);
nor U2475 (N_2475,N_2385,N_2208);
nand U2476 (N_2476,N_2344,N_2204);
nor U2477 (N_2477,N_2343,N_2242);
and U2478 (N_2478,N_2319,N_2317);
and U2479 (N_2479,N_2245,N_2390);
and U2480 (N_2480,N_2305,N_2244);
and U2481 (N_2481,N_2293,N_2309);
or U2482 (N_2482,N_2327,N_2215);
nor U2483 (N_2483,N_2301,N_2281);
nor U2484 (N_2484,N_2269,N_2237);
nor U2485 (N_2485,N_2220,N_2366);
nand U2486 (N_2486,N_2383,N_2266);
and U2487 (N_2487,N_2362,N_2205);
and U2488 (N_2488,N_2326,N_2224);
nand U2489 (N_2489,N_2297,N_2360);
or U2490 (N_2490,N_2257,N_2227);
nand U2491 (N_2491,N_2203,N_2276);
nand U2492 (N_2492,N_2202,N_2246);
and U2493 (N_2493,N_2252,N_2271);
or U2494 (N_2494,N_2261,N_2387);
nand U2495 (N_2495,N_2247,N_2277);
and U2496 (N_2496,N_2299,N_2292);
nor U2497 (N_2497,N_2278,N_2316);
nand U2498 (N_2498,N_2211,N_2201);
nor U2499 (N_2499,N_2288,N_2351);
or U2500 (N_2500,N_2275,N_2387);
or U2501 (N_2501,N_2201,N_2392);
nor U2502 (N_2502,N_2238,N_2297);
nand U2503 (N_2503,N_2331,N_2352);
nor U2504 (N_2504,N_2379,N_2258);
or U2505 (N_2505,N_2303,N_2356);
nand U2506 (N_2506,N_2306,N_2227);
and U2507 (N_2507,N_2268,N_2256);
and U2508 (N_2508,N_2378,N_2206);
or U2509 (N_2509,N_2323,N_2205);
and U2510 (N_2510,N_2254,N_2275);
nor U2511 (N_2511,N_2226,N_2283);
and U2512 (N_2512,N_2352,N_2385);
nor U2513 (N_2513,N_2313,N_2241);
nand U2514 (N_2514,N_2261,N_2356);
or U2515 (N_2515,N_2201,N_2337);
and U2516 (N_2516,N_2264,N_2286);
and U2517 (N_2517,N_2296,N_2217);
nor U2518 (N_2518,N_2252,N_2263);
and U2519 (N_2519,N_2314,N_2342);
nor U2520 (N_2520,N_2261,N_2301);
and U2521 (N_2521,N_2246,N_2313);
and U2522 (N_2522,N_2282,N_2295);
nand U2523 (N_2523,N_2229,N_2214);
or U2524 (N_2524,N_2313,N_2344);
nor U2525 (N_2525,N_2293,N_2292);
nand U2526 (N_2526,N_2305,N_2335);
or U2527 (N_2527,N_2249,N_2225);
nor U2528 (N_2528,N_2323,N_2331);
and U2529 (N_2529,N_2348,N_2287);
and U2530 (N_2530,N_2397,N_2232);
nand U2531 (N_2531,N_2200,N_2227);
and U2532 (N_2532,N_2265,N_2398);
or U2533 (N_2533,N_2222,N_2275);
and U2534 (N_2534,N_2291,N_2264);
or U2535 (N_2535,N_2248,N_2254);
and U2536 (N_2536,N_2229,N_2222);
or U2537 (N_2537,N_2237,N_2289);
nand U2538 (N_2538,N_2211,N_2281);
nand U2539 (N_2539,N_2375,N_2377);
or U2540 (N_2540,N_2356,N_2333);
nand U2541 (N_2541,N_2395,N_2224);
nor U2542 (N_2542,N_2249,N_2274);
xnor U2543 (N_2543,N_2228,N_2297);
or U2544 (N_2544,N_2203,N_2226);
nor U2545 (N_2545,N_2393,N_2258);
and U2546 (N_2546,N_2306,N_2295);
nand U2547 (N_2547,N_2356,N_2324);
or U2548 (N_2548,N_2301,N_2222);
or U2549 (N_2549,N_2316,N_2262);
nand U2550 (N_2550,N_2396,N_2247);
and U2551 (N_2551,N_2284,N_2213);
nand U2552 (N_2552,N_2233,N_2241);
nor U2553 (N_2553,N_2366,N_2393);
nand U2554 (N_2554,N_2387,N_2222);
and U2555 (N_2555,N_2375,N_2220);
or U2556 (N_2556,N_2311,N_2323);
xnor U2557 (N_2557,N_2354,N_2274);
or U2558 (N_2558,N_2218,N_2277);
nor U2559 (N_2559,N_2379,N_2264);
and U2560 (N_2560,N_2290,N_2355);
nand U2561 (N_2561,N_2279,N_2227);
nor U2562 (N_2562,N_2367,N_2242);
and U2563 (N_2563,N_2360,N_2260);
or U2564 (N_2564,N_2394,N_2395);
nor U2565 (N_2565,N_2349,N_2298);
and U2566 (N_2566,N_2213,N_2326);
nand U2567 (N_2567,N_2240,N_2273);
or U2568 (N_2568,N_2284,N_2272);
nor U2569 (N_2569,N_2371,N_2333);
nand U2570 (N_2570,N_2276,N_2359);
nor U2571 (N_2571,N_2398,N_2300);
and U2572 (N_2572,N_2229,N_2321);
nor U2573 (N_2573,N_2202,N_2218);
and U2574 (N_2574,N_2341,N_2257);
nor U2575 (N_2575,N_2255,N_2374);
or U2576 (N_2576,N_2315,N_2281);
or U2577 (N_2577,N_2276,N_2242);
or U2578 (N_2578,N_2389,N_2262);
and U2579 (N_2579,N_2268,N_2291);
nand U2580 (N_2580,N_2251,N_2377);
and U2581 (N_2581,N_2200,N_2357);
nor U2582 (N_2582,N_2334,N_2369);
nand U2583 (N_2583,N_2318,N_2313);
or U2584 (N_2584,N_2375,N_2248);
or U2585 (N_2585,N_2236,N_2336);
nor U2586 (N_2586,N_2296,N_2396);
or U2587 (N_2587,N_2203,N_2339);
nand U2588 (N_2588,N_2274,N_2373);
nor U2589 (N_2589,N_2339,N_2346);
nor U2590 (N_2590,N_2388,N_2369);
nand U2591 (N_2591,N_2262,N_2396);
and U2592 (N_2592,N_2203,N_2202);
or U2593 (N_2593,N_2342,N_2362);
nand U2594 (N_2594,N_2379,N_2372);
and U2595 (N_2595,N_2261,N_2341);
or U2596 (N_2596,N_2248,N_2261);
and U2597 (N_2597,N_2210,N_2367);
and U2598 (N_2598,N_2227,N_2335);
nand U2599 (N_2599,N_2307,N_2358);
and U2600 (N_2600,N_2552,N_2407);
and U2601 (N_2601,N_2563,N_2573);
and U2602 (N_2602,N_2421,N_2450);
nor U2603 (N_2603,N_2591,N_2577);
and U2604 (N_2604,N_2442,N_2504);
xnor U2605 (N_2605,N_2477,N_2571);
or U2606 (N_2606,N_2439,N_2433);
and U2607 (N_2607,N_2443,N_2444);
and U2608 (N_2608,N_2466,N_2454);
nor U2609 (N_2609,N_2546,N_2515);
and U2610 (N_2610,N_2523,N_2536);
or U2611 (N_2611,N_2413,N_2501);
nor U2612 (N_2612,N_2514,N_2550);
and U2613 (N_2613,N_2570,N_2446);
and U2614 (N_2614,N_2489,N_2415);
nand U2615 (N_2615,N_2425,N_2568);
nand U2616 (N_2616,N_2426,N_2435);
or U2617 (N_2617,N_2558,N_2512);
and U2618 (N_2618,N_2499,N_2471);
nand U2619 (N_2619,N_2434,N_2592);
nand U2620 (N_2620,N_2566,N_2447);
or U2621 (N_2621,N_2596,N_2493);
nor U2622 (N_2622,N_2500,N_2430);
and U2623 (N_2623,N_2508,N_2498);
or U2624 (N_2624,N_2428,N_2467);
nand U2625 (N_2625,N_2470,N_2409);
and U2626 (N_2626,N_2416,N_2559);
nor U2627 (N_2627,N_2551,N_2495);
and U2628 (N_2628,N_2438,N_2507);
and U2629 (N_2629,N_2457,N_2494);
xor U2630 (N_2630,N_2548,N_2528);
or U2631 (N_2631,N_2530,N_2429);
nor U2632 (N_2632,N_2448,N_2517);
xnor U2633 (N_2633,N_2565,N_2532);
nand U2634 (N_2634,N_2583,N_2572);
nand U2635 (N_2635,N_2486,N_2585);
and U2636 (N_2636,N_2518,N_2455);
or U2637 (N_2637,N_2414,N_2516);
or U2638 (N_2638,N_2574,N_2549);
nor U2639 (N_2639,N_2474,N_2488);
or U2640 (N_2640,N_2529,N_2436);
nand U2641 (N_2641,N_2403,N_2458);
nor U2642 (N_2642,N_2555,N_2598);
nand U2643 (N_2643,N_2543,N_2535);
and U2644 (N_2644,N_2479,N_2408);
nor U2645 (N_2645,N_2424,N_2472);
nor U2646 (N_2646,N_2581,N_2513);
xor U2647 (N_2647,N_2589,N_2502);
or U2648 (N_2648,N_2449,N_2402);
and U2649 (N_2649,N_2561,N_2483);
or U2650 (N_2650,N_2463,N_2460);
nand U2651 (N_2651,N_2554,N_2491);
or U2652 (N_2652,N_2468,N_2484);
nand U2653 (N_2653,N_2580,N_2509);
nand U2654 (N_2654,N_2497,N_2410);
and U2655 (N_2655,N_2478,N_2419);
and U2656 (N_2656,N_2441,N_2593);
or U2657 (N_2657,N_2553,N_2576);
nor U2658 (N_2658,N_2562,N_2462);
nor U2659 (N_2659,N_2496,N_2584);
or U2660 (N_2660,N_2503,N_2524);
nor U2661 (N_2661,N_2437,N_2542);
nand U2662 (N_2662,N_2545,N_2431);
or U2663 (N_2663,N_2459,N_2588);
and U2664 (N_2664,N_2420,N_2445);
nand U2665 (N_2665,N_2567,N_2505);
nand U2666 (N_2666,N_2586,N_2534);
nor U2667 (N_2667,N_2531,N_2487);
or U2668 (N_2668,N_2527,N_2511);
nand U2669 (N_2669,N_2520,N_2476);
and U2670 (N_2670,N_2564,N_2556);
or U2671 (N_2671,N_2599,N_2453);
nor U2672 (N_2672,N_2506,N_2539);
nand U2673 (N_2673,N_2537,N_2473);
and U2674 (N_2674,N_2575,N_2490);
nor U2675 (N_2675,N_2522,N_2461);
nand U2676 (N_2676,N_2417,N_2579);
and U2677 (N_2677,N_2406,N_2540);
and U2678 (N_2678,N_2469,N_2481);
nand U2679 (N_2679,N_2526,N_2485);
nor U2680 (N_2680,N_2475,N_2451);
and U2681 (N_2681,N_2412,N_2594);
and U2682 (N_2682,N_2557,N_2465);
nor U2683 (N_2683,N_2423,N_2578);
nor U2684 (N_2684,N_2405,N_2541);
nand U2685 (N_2685,N_2533,N_2560);
and U2686 (N_2686,N_2525,N_2482);
or U2687 (N_2687,N_2440,N_2492);
and U2688 (N_2688,N_2401,N_2427);
nand U2689 (N_2689,N_2510,N_2521);
nor U2690 (N_2690,N_2480,N_2569);
nor U2691 (N_2691,N_2582,N_2597);
or U2692 (N_2692,N_2590,N_2452);
and U2693 (N_2693,N_2418,N_2538);
or U2694 (N_2694,N_2404,N_2456);
nor U2695 (N_2695,N_2547,N_2544);
nand U2696 (N_2696,N_2422,N_2464);
and U2697 (N_2697,N_2432,N_2595);
or U2698 (N_2698,N_2400,N_2411);
nand U2699 (N_2699,N_2519,N_2587);
nand U2700 (N_2700,N_2534,N_2594);
nand U2701 (N_2701,N_2476,N_2508);
nand U2702 (N_2702,N_2595,N_2532);
nand U2703 (N_2703,N_2489,N_2485);
nand U2704 (N_2704,N_2589,N_2421);
nand U2705 (N_2705,N_2568,N_2582);
nor U2706 (N_2706,N_2442,N_2464);
nand U2707 (N_2707,N_2487,N_2436);
nand U2708 (N_2708,N_2532,N_2437);
and U2709 (N_2709,N_2506,N_2557);
or U2710 (N_2710,N_2562,N_2479);
or U2711 (N_2711,N_2469,N_2420);
or U2712 (N_2712,N_2466,N_2451);
and U2713 (N_2713,N_2450,N_2595);
nand U2714 (N_2714,N_2473,N_2485);
and U2715 (N_2715,N_2445,N_2579);
nor U2716 (N_2716,N_2556,N_2586);
and U2717 (N_2717,N_2473,N_2557);
nor U2718 (N_2718,N_2502,N_2483);
nor U2719 (N_2719,N_2589,N_2596);
nand U2720 (N_2720,N_2554,N_2447);
or U2721 (N_2721,N_2597,N_2448);
or U2722 (N_2722,N_2556,N_2515);
or U2723 (N_2723,N_2468,N_2506);
or U2724 (N_2724,N_2494,N_2496);
nor U2725 (N_2725,N_2460,N_2550);
or U2726 (N_2726,N_2581,N_2500);
or U2727 (N_2727,N_2580,N_2412);
nand U2728 (N_2728,N_2504,N_2405);
or U2729 (N_2729,N_2516,N_2444);
nor U2730 (N_2730,N_2554,N_2577);
nand U2731 (N_2731,N_2502,N_2592);
nand U2732 (N_2732,N_2418,N_2502);
nor U2733 (N_2733,N_2537,N_2453);
and U2734 (N_2734,N_2598,N_2465);
nand U2735 (N_2735,N_2501,N_2401);
or U2736 (N_2736,N_2540,N_2563);
or U2737 (N_2737,N_2454,N_2506);
or U2738 (N_2738,N_2407,N_2423);
and U2739 (N_2739,N_2416,N_2582);
nor U2740 (N_2740,N_2543,N_2441);
and U2741 (N_2741,N_2437,N_2534);
nor U2742 (N_2742,N_2459,N_2426);
or U2743 (N_2743,N_2513,N_2431);
xnor U2744 (N_2744,N_2558,N_2509);
nand U2745 (N_2745,N_2482,N_2530);
or U2746 (N_2746,N_2402,N_2465);
and U2747 (N_2747,N_2583,N_2490);
nand U2748 (N_2748,N_2498,N_2496);
nand U2749 (N_2749,N_2582,N_2487);
and U2750 (N_2750,N_2534,N_2585);
nor U2751 (N_2751,N_2419,N_2490);
nand U2752 (N_2752,N_2559,N_2469);
nor U2753 (N_2753,N_2525,N_2560);
nand U2754 (N_2754,N_2458,N_2553);
and U2755 (N_2755,N_2520,N_2596);
and U2756 (N_2756,N_2528,N_2550);
nand U2757 (N_2757,N_2454,N_2445);
nand U2758 (N_2758,N_2471,N_2520);
nand U2759 (N_2759,N_2545,N_2581);
and U2760 (N_2760,N_2557,N_2433);
nor U2761 (N_2761,N_2409,N_2588);
or U2762 (N_2762,N_2471,N_2549);
nand U2763 (N_2763,N_2479,N_2533);
nand U2764 (N_2764,N_2407,N_2581);
or U2765 (N_2765,N_2566,N_2497);
and U2766 (N_2766,N_2553,N_2511);
nor U2767 (N_2767,N_2478,N_2501);
nand U2768 (N_2768,N_2575,N_2468);
nor U2769 (N_2769,N_2447,N_2574);
nor U2770 (N_2770,N_2501,N_2531);
and U2771 (N_2771,N_2442,N_2581);
nor U2772 (N_2772,N_2543,N_2516);
nand U2773 (N_2773,N_2554,N_2597);
nor U2774 (N_2774,N_2418,N_2575);
nand U2775 (N_2775,N_2438,N_2500);
or U2776 (N_2776,N_2529,N_2571);
or U2777 (N_2777,N_2587,N_2449);
or U2778 (N_2778,N_2495,N_2499);
nand U2779 (N_2779,N_2509,N_2575);
or U2780 (N_2780,N_2417,N_2599);
and U2781 (N_2781,N_2536,N_2572);
nor U2782 (N_2782,N_2425,N_2472);
nor U2783 (N_2783,N_2519,N_2460);
or U2784 (N_2784,N_2592,N_2463);
nor U2785 (N_2785,N_2411,N_2405);
or U2786 (N_2786,N_2549,N_2414);
or U2787 (N_2787,N_2595,N_2540);
nand U2788 (N_2788,N_2517,N_2546);
nor U2789 (N_2789,N_2453,N_2433);
nand U2790 (N_2790,N_2424,N_2455);
or U2791 (N_2791,N_2425,N_2449);
or U2792 (N_2792,N_2508,N_2583);
nand U2793 (N_2793,N_2561,N_2530);
nor U2794 (N_2794,N_2467,N_2466);
nand U2795 (N_2795,N_2567,N_2579);
or U2796 (N_2796,N_2448,N_2443);
nor U2797 (N_2797,N_2408,N_2599);
and U2798 (N_2798,N_2489,N_2488);
and U2799 (N_2799,N_2472,N_2459);
xnor U2800 (N_2800,N_2686,N_2692);
nand U2801 (N_2801,N_2709,N_2630);
nand U2802 (N_2802,N_2677,N_2687);
nor U2803 (N_2803,N_2729,N_2769);
nor U2804 (N_2804,N_2675,N_2740);
or U2805 (N_2805,N_2705,N_2738);
and U2806 (N_2806,N_2690,N_2639);
nand U2807 (N_2807,N_2606,N_2614);
nor U2808 (N_2808,N_2652,N_2715);
and U2809 (N_2809,N_2615,N_2607);
and U2810 (N_2810,N_2665,N_2622);
nand U2811 (N_2811,N_2646,N_2793);
and U2812 (N_2812,N_2758,N_2695);
or U2813 (N_2813,N_2696,N_2643);
and U2814 (N_2814,N_2693,N_2795);
nand U2815 (N_2815,N_2689,N_2697);
or U2816 (N_2816,N_2703,N_2633);
or U2817 (N_2817,N_2678,N_2766);
and U2818 (N_2818,N_2787,N_2747);
or U2819 (N_2819,N_2628,N_2604);
or U2820 (N_2820,N_2711,N_2702);
nand U2821 (N_2821,N_2650,N_2620);
nand U2822 (N_2822,N_2717,N_2799);
or U2823 (N_2823,N_2656,N_2765);
or U2824 (N_2824,N_2760,N_2618);
and U2825 (N_2825,N_2624,N_2636);
or U2826 (N_2826,N_2726,N_2660);
or U2827 (N_2827,N_2716,N_2623);
xor U2828 (N_2828,N_2775,N_2776);
nor U2829 (N_2829,N_2786,N_2701);
or U2830 (N_2830,N_2757,N_2661);
nand U2831 (N_2831,N_2704,N_2626);
or U2832 (N_2832,N_2640,N_2791);
xnor U2833 (N_2833,N_2772,N_2730);
or U2834 (N_2834,N_2753,N_2649);
nor U2835 (N_2835,N_2669,N_2631);
or U2836 (N_2836,N_2610,N_2632);
and U2837 (N_2837,N_2612,N_2780);
or U2838 (N_2838,N_2684,N_2714);
xnor U2839 (N_2839,N_2733,N_2790);
or U2840 (N_2840,N_2625,N_2641);
or U2841 (N_2841,N_2655,N_2731);
nor U2842 (N_2842,N_2601,N_2779);
nor U2843 (N_2843,N_2768,N_2734);
nor U2844 (N_2844,N_2764,N_2739);
or U2845 (N_2845,N_2647,N_2736);
nor U2846 (N_2846,N_2763,N_2755);
nor U2847 (N_2847,N_2611,N_2627);
or U2848 (N_2848,N_2629,N_2666);
or U2849 (N_2849,N_2659,N_2635);
and U2850 (N_2850,N_2648,N_2712);
and U2851 (N_2851,N_2746,N_2663);
or U2852 (N_2852,N_2638,N_2671);
nand U2853 (N_2853,N_2685,N_2699);
nand U2854 (N_2854,N_2676,N_2613);
nand U2855 (N_2855,N_2688,N_2708);
and U2856 (N_2856,N_2745,N_2681);
and U2857 (N_2857,N_2720,N_2670);
nor U2858 (N_2858,N_2721,N_2773);
and U2859 (N_2859,N_2789,N_2744);
nor U2860 (N_2860,N_2771,N_2637);
or U2861 (N_2861,N_2683,N_2707);
nor U2862 (N_2862,N_2735,N_2634);
and U2863 (N_2863,N_2698,N_2674);
or U2864 (N_2864,N_2722,N_2718);
or U2865 (N_2865,N_2759,N_2784);
xor U2866 (N_2866,N_2651,N_2602);
nor U2867 (N_2867,N_2658,N_2619);
or U2868 (N_2868,N_2668,N_2706);
and U2869 (N_2869,N_2737,N_2644);
and U2870 (N_2870,N_2751,N_2798);
nand U2871 (N_2871,N_2761,N_2617);
nor U2872 (N_2872,N_2605,N_2667);
nor U2873 (N_2873,N_2792,N_2672);
nand U2874 (N_2874,N_2742,N_2725);
and U2875 (N_2875,N_2788,N_2682);
nand U2876 (N_2876,N_2794,N_2741);
nand U2877 (N_2877,N_2694,N_2750);
and U2878 (N_2878,N_2783,N_2608);
nor U2879 (N_2879,N_2654,N_2645);
xnor U2880 (N_2880,N_2728,N_2785);
nor U2881 (N_2881,N_2621,N_2782);
nor U2882 (N_2882,N_2748,N_2662);
and U2883 (N_2883,N_2691,N_2664);
nor U2884 (N_2884,N_2754,N_2673);
xor U2885 (N_2885,N_2710,N_2723);
nand U2886 (N_2886,N_2713,N_2749);
nor U2887 (N_2887,N_2680,N_2732);
and U2888 (N_2888,N_2653,N_2767);
and U2889 (N_2889,N_2603,N_2724);
or U2890 (N_2890,N_2657,N_2700);
nand U2891 (N_2891,N_2752,N_2727);
or U2892 (N_2892,N_2781,N_2762);
and U2893 (N_2893,N_2600,N_2797);
or U2894 (N_2894,N_2770,N_2616);
nand U2895 (N_2895,N_2719,N_2774);
nand U2896 (N_2896,N_2756,N_2778);
or U2897 (N_2897,N_2743,N_2642);
nand U2898 (N_2898,N_2777,N_2609);
or U2899 (N_2899,N_2679,N_2796);
nor U2900 (N_2900,N_2753,N_2694);
nand U2901 (N_2901,N_2656,N_2784);
and U2902 (N_2902,N_2795,N_2779);
or U2903 (N_2903,N_2742,N_2702);
and U2904 (N_2904,N_2715,N_2776);
nor U2905 (N_2905,N_2668,N_2709);
and U2906 (N_2906,N_2713,N_2720);
nor U2907 (N_2907,N_2790,N_2685);
and U2908 (N_2908,N_2676,N_2748);
and U2909 (N_2909,N_2606,N_2605);
and U2910 (N_2910,N_2735,N_2654);
and U2911 (N_2911,N_2774,N_2627);
nor U2912 (N_2912,N_2781,N_2645);
or U2913 (N_2913,N_2722,N_2736);
nor U2914 (N_2914,N_2645,N_2633);
and U2915 (N_2915,N_2717,N_2780);
nor U2916 (N_2916,N_2624,N_2667);
nand U2917 (N_2917,N_2751,N_2787);
or U2918 (N_2918,N_2786,N_2737);
nand U2919 (N_2919,N_2744,N_2763);
nor U2920 (N_2920,N_2684,N_2645);
and U2921 (N_2921,N_2765,N_2763);
nand U2922 (N_2922,N_2661,N_2690);
nand U2923 (N_2923,N_2630,N_2663);
or U2924 (N_2924,N_2677,N_2662);
nor U2925 (N_2925,N_2700,N_2611);
and U2926 (N_2926,N_2619,N_2702);
or U2927 (N_2927,N_2791,N_2730);
or U2928 (N_2928,N_2743,N_2661);
or U2929 (N_2929,N_2774,N_2695);
nand U2930 (N_2930,N_2794,N_2688);
or U2931 (N_2931,N_2679,N_2617);
nor U2932 (N_2932,N_2718,N_2710);
nor U2933 (N_2933,N_2678,N_2730);
nor U2934 (N_2934,N_2701,N_2731);
or U2935 (N_2935,N_2723,N_2799);
or U2936 (N_2936,N_2651,N_2737);
and U2937 (N_2937,N_2640,N_2684);
nand U2938 (N_2938,N_2661,N_2602);
and U2939 (N_2939,N_2766,N_2777);
nor U2940 (N_2940,N_2662,N_2719);
nor U2941 (N_2941,N_2753,N_2792);
nand U2942 (N_2942,N_2710,N_2651);
or U2943 (N_2943,N_2648,N_2729);
xnor U2944 (N_2944,N_2715,N_2707);
nor U2945 (N_2945,N_2788,N_2793);
nor U2946 (N_2946,N_2661,N_2708);
nand U2947 (N_2947,N_2669,N_2625);
or U2948 (N_2948,N_2626,N_2602);
or U2949 (N_2949,N_2686,N_2610);
or U2950 (N_2950,N_2780,N_2636);
or U2951 (N_2951,N_2650,N_2762);
or U2952 (N_2952,N_2684,N_2736);
or U2953 (N_2953,N_2665,N_2701);
or U2954 (N_2954,N_2796,N_2602);
and U2955 (N_2955,N_2629,N_2785);
and U2956 (N_2956,N_2745,N_2649);
or U2957 (N_2957,N_2679,N_2766);
nor U2958 (N_2958,N_2666,N_2646);
and U2959 (N_2959,N_2626,N_2694);
or U2960 (N_2960,N_2652,N_2644);
nor U2961 (N_2961,N_2725,N_2652);
nand U2962 (N_2962,N_2624,N_2660);
xnor U2963 (N_2963,N_2612,N_2719);
and U2964 (N_2964,N_2751,N_2749);
nor U2965 (N_2965,N_2728,N_2716);
nand U2966 (N_2966,N_2747,N_2698);
nand U2967 (N_2967,N_2790,N_2724);
nor U2968 (N_2968,N_2633,N_2615);
nand U2969 (N_2969,N_2778,N_2651);
or U2970 (N_2970,N_2616,N_2645);
or U2971 (N_2971,N_2607,N_2742);
nor U2972 (N_2972,N_2792,N_2697);
nor U2973 (N_2973,N_2776,N_2644);
xor U2974 (N_2974,N_2726,N_2779);
or U2975 (N_2975,N_2612,N_2666);
nand U2976 (N_2976,N_2633,N_2647);
nand U2977 (N_2977,N_2779,N_2663);
nor U2978 (N_2978,N_2609,N_2749);
and U2979 (N_2979,N_2688,N_2752);
nor U2980 (N_2980,N_2776,N_2793);
nand U2981 (N_2981,N_2765,N_2761);
and U2982 (N_2982,N_2692,N_2788);
nor U2983 (N_2983,N_2743,N_2673);
nor U2984 (N_2984,N_2602,N_2652);
or U2985 (N_2985,N_2676,N_2671);
or U2986 (N_2986,N_2796,N_2734);
nand U2987 (N_2987,N_2786,N_2617);
or U2988 (N_2988,N_2757,N_2700);
nor U2989 (N_2989,N_2743,N_2733);
or U2990 (N_2990,N_2702,N_2699);
nor U2991 (N_2991,N_2725,N_2747);
and U2992 (N_2992,N_2700,N_2721);
nor U2993 (N_2993,N_2717,N_2612);
nand U2994 (N_2994,N_2772,N_2691);
nand U2995 (N_2995,N_2682,N_2735);
and U2996 (N_2996,N_2618,N_2608);
nand U2997 (N_2997,N_2759,N_2774);
or U2998 (N_2998,N_2752,N_2656);
nor U2999 (N_2999,N_2608,N_2620);
nand UO_0 (O_0,N_2879,N_2928);
or UO_1 (O_1,N_2853,N_2826);
and UO_2 (O_2,N_2944,N_2867);
nor UO_3 (O_3,N_2852,N_2830);
nor UO_4 (O_4,N_2838,N_2962);
and UO_5 (O_5,N_2903,N_2803);
nor UO_6 (O_6,N_2976,N_2883);
and UO_7 (O_7,N_2851,N_2896);
or UO_8 (O_8,N_2990,N_2835);
or UO_9 (O_9,N_2902,N_2824);
nand UO_10 (O_10,N_2884,N_2829);
nor UO_11 (O_11,N_2865,N_2897);
nor UO_12 (O_12,N_2961,N_2987);
nor UO_13 (O_13,N_2887,N_2832);
or UO_14 (O_14,N_2945,N_2818);
or UO_15 (O_15,N_2996,N_2871);
nor UO_16 (O_16,N_2842,N_2959);
nand UO_17 (O_17,N_2821,N_2979);
and UO_18 (O_18,N_2825,N_2918);
and UO_19 (O_19,N_2877,N_2828);
nor UO_20 (O_20,N_2983,N_2814);
and UO_21 (O_21,N_2864,N_2890);
nor UO_22 (O_22,N_2866,N_2977);
and UO_23 (O_23,N_2822,N_2857);
nand UO_24 (O_24,N_2949,N_2910);
nor UO_25 (O_25,N_2809,N_2938);
nor UO_26 (O_26,N_2966,N_2982);
nor UO_27 (O_27,N_2882,N_2974);
nor UO_28 (O_28,N_2827,N_2833);
nand UO_29 (O_29,N_2817,N_2837);
nor UO_30 (O_30,N_2813,N_2885);
nand UO_31 (O_31,N_2820,N_2940);
and UO_32 (O_32,N_2873,N_2800);
and UO_33 (O_33,N_2921,N_2901);
nand UO_34 (O_34,N_2964,N_2891);
or UO_35 (O_35,N_2823,N_2971);
nor UO_36 (O_36,N_2954,N_2908);
nor UO_37 (O_37,N_2839,N_2915);
nor UO_38 (O_38,N_2973,N_2953);
and UO_39 (O_39,N_2899,N_2920);
nor UO_40 (O_40,N_2952,N_2812);
and UO_41 (O_41,N_2846,N_2948);
and UO_42 (O_42,N_2854,N_2937);
and UO_43 (O_43,N_2926,N_2863);
nand UO_44 (O_44,N_2845,N_2930);
and UO_45 (O_45,N_2840,N_2925);
nor UO_46 (O_46,N_2975,N_2931);
and UO_47 (O_47,N_2900,N_2980);
or UO_48 (O_48,N_2893,N_2965);
nor UO_49 (O_49,N_2984,N_2881);
or UO_50 (O_50,N_2905,N_2811);
nor UO_51 (O_51,N_2993,N_2988);
nor UO_52 (O_52,N_2922,N_2889);
xnor UO_53 (O_53,N_2859,N_2956);
and UO_54 (O_54,N_2861,N_2967);
nand UO_55 (O_55,N_2841,N_2894);
xnor UO_56 (O_56,N_2935,N_2994);
or UO_57 (O_57,N_2955,N_2860);
and UO_58 (O_58,N_2815,N_2880);
nor UO_59 (O_59,N_2950,N_2816);
nand UO_60 (O_60,N_2913,N_2942);
and UO_61 (O_61,N_2912,N_2892);
or UO_62 (O_62,N_2936,N_2986);
and UO_63 (O_63,N_2998,N_2907);
xnor UO_64 (O_64,N_2849,N_2848);
nand UO_65 (O_65,N_2963,N_2970);
nor UO_66 (O_66,N_2939,N_2991);
and UO_67 (O_67,N_2904,N_2801);
nand UO_68 (O_68,N_2909,N_2929);
nor UO_69 (O_69,N_2927,N_2947);
or UO_70 (O_70,N_2810,N_2850);
and UO_71 (O_71,N_2878,N_2856);
or UO_72 (O_72,N_2847,N_2951);
nand UO_73 (O_73,N_2888,N_2981);
nand UO_74 (O_74,N_2958,N_2834);
nor UO_75 (O_75,N_2968,N_2868);
and UO_76 (O_76,N_2872,N_2992);
nand UO_77 (O_77,N_2911,N_2844);
nand UO_78 (O_78,N_2919,N_2855);
nor UO_79 (O_79,N_2933,N_2836);
nor UO_80 (O_80,N_2924,N_2819);
and UO_81 (O_81,N_2802,N_2869);
nor UO_82 (O_82,N_2999,N_2916);
nor UO_83 (O_83,N_2960,N_2862);
nor UO_84 (O_84,N_2876,N_2808);
nor UO_85 (O_85,N_2875,N_2805);
nand UO_86 (O_86,N_2946,N_2858);
nand UO_87 (O_87,N_2804,N_2870);
or UO_88 (O_88,N_2941,N_2985);
or UO_89 (O_89,N_2807,N_2917);
and UO_90 (O_90,N_2995,N_2895);
or UO_91 (O_91,N_2932,N_2914);
xnor UO_92 (O_92,N_2898,N_2957);
or UO_93 (O_93,N_2806,N_2843);
nor UO_94 (O_94,N_2923,N_2997);
nand UO_95 (O_95,N_2906,N_2874);
nand UO_96 (O_96,N_2831,N_2978);
nand UO_97 (O_97,N_2989,N_2934);
nor UO_98 (O_98,N_2972,N_2943);
and UO_99 (O_99,N_2969,N_2886);
or UO_100 (O_100,N_2935,N_2903);
nor UO_101 (O_101,N_2861,N_2868);
and UO_102 (O_102,N_2960,N_2921);
nor UO_103 (O_103,N_2850,N_2861);
nand UO_104 (O_104,N_2912,N_2957);
nor UO_105 (O_105,N_2963,N_2810);
or UO_106 (O_106,N_2815,N_2848);
xor UO_107 (O_107,N_2946,N_2979);
or UO_108 (O_108,N_2969,N_2991);
nand UO_109 (O_109,N_2811,N_2936);
or UO_110 (O_110,N_2947,N_2931);
nand UO_111 (O_111,N_2938,N_2939);
nand UO_112 (O_112,N_2936,N_2958);
xnor UO_113 (O_113,N_2912,N_2956);
nor UO_114 (O_114,N_2911,N_2940);
or UO_115 (O_115,N_2995,N_2944);
and UO_116 (O_116,N_2833,N_2869);
or UO_117 (O_117,N_2907,N_2956);
nand UO_118 (O_118,N_2900,N_2838);
nand UO_119 (O_119,N_2858,N_2893);
and UO_120 (O_120,N_2948,N_2855);
and UO_121 (O_121,N_2871,N_2907);
and UO_122 (O_122,N_2860,N_2949);
nor UO_123 (O_123,N_2833,N_2968);
nand UO_124 (O_124,N_2852,N_2813);
nor UO_125 (O_125,N_2894,N_2876);
nor UO_126 (O_126,N_2803,N_2962);
and UO_127 (O_127,N_2940,N_2904);
and UO_128 (O_128,N_2832,N_2883);
nor UO_129 (O_129,N_2898,N_2949);
nand UO_130 (O_130,N_2937,N_2941);
nor UO_131 (O_131,N_2871,N_2828);
nor UO_132 (O_132,N_2905,N_2948);
nand UO_133 (O_133,N_2908,N_2880);
nor UO_134 (O_134,N_2929,N_2915);
nand UO_135 (O_135,N_2976,N_2941);
or UO_136 (O_136,N_2816,N_2828);
nand UO_137 (O_137,N_2856,N_2961);
or UO_138 (O_138,N_2810,N_2847);
or UO_139 (O_139,N_2874,N_2960);
or UO_140 (O_140,N_2993,N_2913);
and UO_141 (O_141,N_2973,N_2841);
and UO_142 (O_142,N_2894,N_2882);
nand UO_143 (O_143,N_2876,N_2994);
nor UO_144 (O_144,N_2939,N_2956);
xnor UO_145 (O_145,N_2956,N_2806);
xor UO_146 (O_146,N_2856,N_2841);
nand UO_147 (O_147,N_2895,N_2937);
and UO_148 (O_148,N_2948,N_2871);
or UO_149 (O_149,N_2969,N_2865);
and UO_150 (O_150,N_2889,N_2878);
and UO_151 (O_151,N_2859,N_2955);
or UO_152 (O_152,N_2994,N_2885);
nand UO_153 (O_153,N_2831,N_2813);
nor UO_154 (O_154,N_2984,N_2863);
and UO_155 (O_155,N_2867,N_2923);
nor UO_156 (O_156,N_2947,N_2894);
nor UO_157 (O_157,N_2888,N_2827);
and UO_158 (O_158,N_2847,N_2836);
nor UO_159 (O_159,N_2928,N_2906);
nor UO_160 (O_160,N_2943,N_2944);
or UO_161 (O_161,N_2826,N_2827);
and UO_162 (O_162,N_2843,N_2814);
and UO_163 (O_163,N_2911,N_2864);
or UO_164 (O_164,N_2911,N_2944);
nand UO_165 (O_165,N_2918,N_2904);
nor UO_166 (O_166,N_2915,N_2986);
nand UO_167 (O_167,N_2975,N_2863);
or UO_168 (O_168,N_2871,N_2951);
and UO_169 (O_169,N_2949,N_2806);
nand UO_170 (O_170,N_2939,N_2868);
and UO_171 (O_171,N_2803,N_2958);
and UO_172 (O_172,N_2974,N_2913);
and UO_173 (O_173,N_2816,N_2837);
and UO_174 (O_174,N_2868,N_2832);
and UO_175 (O_175,N_2849,N_2929);
nand UO_176 (O_176,N_2938,N_2808);
or UO_177 (O_177,N_2811,N_2964);
or UO_178 (O_178,N_2930,N_2829);
nor UO_179 (O_179,N_2863,N_2837);
nor UO_180 (O_180,N_2838,N_2972);
nor UO_181 (O_181,N_2811,N_2924);
xor UO_182 (O_182,N_2946,N_2826);
or UO_183 (O_183,N_2912,N_2879);
nand UO_184 (O_184,N_2911,N_2834);
and UO_185 (O_185,N_2887,N_2851);
nor UO_186 (O_186,N_2860,N_2847);
and UO_187 (O_187,N_2986,N_2882);
nor UO_188 (O_188,N_2942,N_2840);
nand UO_189 (O_189,N_2839,N_2853);
nor UO_190 (O_190,N_2920,N_2854);
nor UO_191 (O_191,N_2883,N_2990);
and UO_192 (O_192,N_2896,N_2962);
or UO_193 (O_193,N_2850,N_2976);
nand UO_194 (O_194,N_2861,N_2878);
nand UO_195 (O_195,N_2872,N_2975);
nand UO_196 (O_196,N_2986,N_2920);
or UO_197 (O_197,N_2821,N_2868);
and UO_198 (O_198,N_2863,N_2935);
and UO_199 (O_199,N_2907,N_2850);
and UO_200 (O_200,N_2913,N_2995);
nand UO_201 (O_201,N_2947,N_2831);
nand UO_202 (O_202,N_2970,N_2886);
or UO_203 (O_203,N_2868,N_2844);
or UO_204 (O_204,N_2814,N_2882);
nor UO_205 (O_205,N_2848,N_2887);
and UO_206 (O_206,N_2928,N_2940);
nand UO_207 (O_207,N_2801,N_2813);
nor UO_208 (O_208,N_2825,N_2926);
or UO_209 (O_209,N_2896,N_2976);
nand UO_210 (O_210,N_2945,N_2911);
or UO_211 (O_211,N_2827,N_2975);
and UO_212 (O_212,N_2897,N_2985);
and UO_213 (O_213,N_2858,N_2904);
nor UO_214 (O_214,N_2897,N_2887);
nand UO_215 (O_215,N_2874,N_2828);
or UO_216 (O_216,N_2936,N_2869);
or UO_217 (O_217,N_2972,N_2814);
and UO_218 (O_218,N_2952,N_2978);
nand UO_219 (O_219,N_2877,N_2961);
nor UO_220 (O_220,N_2834,N_2818);
or UO_221 (O_221,N_2885,N_2904);
and UO_222 (O_222,N_2929,N_2923);
nor UO_223 (O_223,N_2974,N_2973);
and UO_224 (O_224,N_2847,N_2830);
and UO_225 (O_225,N_2843,N_2916);
nand UO_226 (O_226,N_2937,N_2812);
or UO_227 (O_227,N_2936,N_2902);
nand UO_228 (O_228,N_2939,N_2913);
nand UO_229 (O_229,N_2838,N_2955);
nand UO_230 (O_230,N_2965,N_2996);
and UO_231 (O_231,N_2845,N_2931);
nand UO_232 (O_232,N_2819,N_2949);
nor UO_233 (O_233,N_2881,N_2865);
nor UO_234 (O_234,N_2943,N_2930);
or UO_235 (O_235,N_2965,N_2803);
or UO_236 (O_236,N_2894,N_2878);
and UO_237 (O_237,N_2807,N_2830);
or UO_238 (O_238,N_2911,N_2822);
nand UO_239 (O_239,N_2950,N_2896);
and UO_240 (O_240,N_2976,N_2954);
or UO_241 (O_241,N_2889,N_2932);
nor UO_242 (O_242,N_2930,N_2865);
nand UO_243 (O_243,N_2937,N_2990);
nand UO_244 (O_244,N_2841,N_2955);
nor UO_245 (O_245,N_2974,N_2838);
and UO_246 (O_246,N_2864,N_2982);
nand UO_247 (O_247,N_2823,N_2926);
nand UO_248 (O_248,N_2824,N_2959);
nor UO_249 (O_249,N_2849,N_2869);
and UO_250 (O_250,N_2920,N_2942);
nor UO_251 (O_251,N_2808,N_2842);
or UO_252 (O_252,N_2957,N_2985);
nand UO_253 (O_253,N_2828,N_2833);
and UO_254 (O_254,N_2948,N_2879);
or UO_255 (O_255,N_2825,N_2850);
or UO_256 (O_256,N_2908,N_2887);
nand UO_257 (O_257,N_2937,N_2908);
or UO_258 (O_258,N_2840,N_2927);
and UO_259 (O_259,N_2925,N_2991);
nand UO_260 (O_260,N_2896,N_2927);
nand UO_261 (O_261,N_2878,N_2839);
nand UO_262 (O_262,N_2873,N_2979);
xnor UO_263 (O_263,N_2914,N_2858);
nand UO_264 (O_264,N_2999,N_2921);
nor UO_265 (O_265,N_2854,N_2804);
nor UO_266 (O_266,N_2824,N_2864);
nor UO_267 (O_267,N_2915,N_2987);
nand UO_268 (O_268,N_2824,N_2913);
and UO_269 (O_269,N_2896,N_2848);
or UO_270 (O_270,N_2984,N_2824);
and UO_271 (O_271,N_2938,N_2984);
or UO_272 (O_272,N_2999,N_2893);
and UO_273 (O_273,N_2823,N_2915);
nand UO_274 (O_274,N_2864,N_2934);
or UO_275 (O_275,N_2829,N_2837);
nor UO_276 (O_276,N_2900,N_2918);
nand UO_277 (O_277,N_2903,N_2996);
or UO_278 (O_278,N_2804,N_2921);
or UO_279 (O_279,N_2829,N_2989);
and UO_280 (O_280,N_2820,N_2989);
or UO_281 (O_281,N_2919,N_2984);
nand UO_282 (O_282,N_2969,N_2989);
nor UO_283 (O_283,N_2901,N_2907);
nand UO_284 (O_284,N_2970,N_2999);
and UO_285 (O_285,N_2937,N_2953);
and UO_286 (O_286,N_2913,N_2945);
xnor UO_287 (O_287,N_2845,N_2925);
nor UO_288 (O_288,N_2926,N_2810);
and UO_289 (O_289,N_2993,N_2916);
or UO_290 (O_290,N_2830,N_2939);
nor UO_291 (O_291,N_2810,N_2892);
nor UO_292 (O_292,N_2825,N_2885);
or UO_293 (O_293,N_2866,N_2834);
and UO_294 (O_294,N_2991,N_2839);
or UO_295 (O_295,N_2861,N_2820);
nand UO_296 (O_296,N_2993,N_2975);
or UO_297 (O_297,N_2900,N_2906);
nand UO_298 (O_298,N_2801,N_2875);
and UO_299 (O_299,N_2866,N_2855);
nand UO_300 (O_300,N_2932,N_2915);
or UO_301 (O_301,N_2854,N_2929);
nor UO_302 (O_302,N_2924,N_2813);
or UO_303 (O_303,N_2977,N_2921);
and UO_304 (O_304,N_2870,N_2808);
or UO_305 (O_305,N_2886,N_2974);
xnor UO_306 (O_306,N_2898,N_2829);
nor UO_307 (O_307,N_2933,N_2812);
nand UO_308 (O_308,N_2878,N_2871);
nand UO_309 (O_309,N_2884,N_2863);
nor UO_310 (O_310,N_2913,N_2873);
and UO_311 (O_311,N_2990,N_2804);
nor UO_312 (O_312,N_2926,N_2999);
or UO_313 (O_313,N_2965,N_2941);
and UO_314 (O_314,N_2815,N_2827);
or UO_315 (O_315,N_2898,N_2999);
nor UO_316 (O_316,N_2863,N_2894);
and UO_317 (O_317,N_2928,N_2916);
nor UO_318 (O_318,N_2999,N_2951);
nand UO_319 (O_319,N_2860,N_2859);
nor UO_320 (O_320,N_2957,N_2965);
xnor UO_321 (O_321,N_2979,N_2955);
nor UO_322 (O_322,N_2801,N_2966);
and UO_323 (O_323,N_2826,N_2808);
nand UO_324 (O_324,N_2953,N_2869);
nor UO_325 (O_325,N_2890,N_2885);
nand UO_326 (O_326,N_2920,N_2950);
or UO_327 (O_327,N_2916,N_2888);
nand UO_328 (O_328,N_2941,N_2882);
and UO_329 (O_329,N_2967,N_2834);
nor UO_330 (O_330,N_2867,N_2917);
and UO_331 (O_331,N_2800,N_2889);
or UO_332 (O_332,N_2904,N_2928);
and UO_333 (O_333,N_2841,N_2933);
nand UO_334 (O_334,N_2922,N_2808);
or UO_335 (O_335,N_2945,N_2831);
nand UO_336 (O_336,N_2885,N_2990);
and UO_337 (O_337,N_2866,N_2918);
or UO_338 (O_338,N_2884,N_2959);
and UO_339 (O_339,N_2878,N_2847);
nand UO_340 (O_340,N_2930,N_2899);
and UO_341 (O_341,N_2900,N_2803);
or UO_342 (O_342,N_2826,N_2995);
and UO_343 (O_343,N_2831,N_2883);
nor UO_344 (O_344,N_2969,N_2807);
nand UO_345 (O_345,N_2998,N_2975);
and UO_346 (O_346,N_2859,N_2928);
and UO_347 (O_347,N_2876,N_2996);
or UO_348 (O_348,N_2857,N_2852);
and UO_349 (O_349,N_2906,N_2963);
and UO_350 (O_350,N_2845,N_2820);
and UO_351 (O_351,N_2979,N_2895);
nor UO_352 (O_352,N_2837,N_2951);
nor UO_353 (O_353,N_2946,N_2840);
nor UO_354 (O_354,N_2892,N_2928);
nand UO_355 (O_355,N_2899,N_2951);
or UO_356 (O_356,N_2935,N_2995);
or UO_357 (O_357,N_2851,N_2897);
and UO_358 (O_358,N_2838,N_2927);
nor UO_359 (O_359,N_2945,N_2832);
and UO_360 (O_360,N_2969,N_2983);
or UO_361 (O_361,N_2829,N_2846);
and UO_362 (O_362,N_2851,N_2980);
and UO_363 (O_363,N_2891,N_2988);
and UO_364 (O_364,N_2800,N_2835);
and UO_365 (O_365,N_2857,N_2883);
and UO_366 (O_366,N_2961,N_2941);
or UO_367 (O_367,N_2837,N_2982);
nor UO_368 (O_368,N_2955,N_2840);
or UO_369 (O_369,N_2966,N_2928);
nor UO_370 (O_370,N_2945,N_2987);
nand UO_371 (O_371,N_2946,N_2838);
and UO_372 (O_372,N_2811,N_2888);
and UO_373 (O_373,N_2835,N_2923);
nand UO_374 (O_374,N_2956,N_2817);
or UO_375 (O_375,N_2932,N_2906);
nor UO_376 (O_376,N_2969,N_2809);
and UO_377 (O_377,N_2890,N_2853);
or UO_378 (O_378,N_2869,N_2946);
and UO_379 (O_379,N_2893,N_2875);
nand UO_380 (O_380,N_2958,N_2987);
nand UO_381 (O_381,N_2922,N_2822);
or UO_382 (O_382,N_2817,N_2949);
or UO_383 (O_383,N_2921,N_2964);
or UO_384 (O_384,N_2956,N_2973);
nor UO_385 (O_385,N_2984,N_2878);
and UO_386 (O_386,N_2917,N_2941);
nand UO_387 (O_387,N_2953,N_2936);
xnor UO_388 (O_388,N_2972,N_2860);
nand UO_389 (O_389,N_2951,N_2894);
nand UO_390 (O_390,N_2882,N_2904);
nor UO_391 (O_391,N_2813,N_2920);
nand UO_392 (O_392,N_2883,N_2907);
and UO_393 (O_393,N_2855,N_2956);
nand UO_394 (O_394,N_2849,N_2879);
nand UO_395 (O_395,N_2945,N_2814);
or UO_396 (O_396,N_2874,N_2800);
nand UO_397 (O_397,N_2852,N_2972);
and UO_398 (O_398,N_2897,N_2893);
nor UO_399 (O_399,N_2942,N_2906);
and UO_400 (O_400,N_2857,N_2876);
nand UO_401 (O_401,N_2939,N_2858);
nand UO_402 (O_402,N_2971,N_2829);
or UO_403 (O_403,N_2996,N_2834);
nand UO_404 (O_404,N_2929,N_2866);
or UO_405 (O_405,N_2928,N_2816);
nand UO_406 (O_406,N_2969,N_2999);
nand UO_407 (O_407,N_2908,N_2925);
or UO_408 (O_408,N_2892,N_2815);
nor UO_409 (O_409,N_2888,N_2961);
or UO_410 (O_410,N_2875,N_2903);
nand UO_411 (O_411,N_2840,N_2848);
or UO_412 (O_412,N_2854,N_2868);
and UO_413 (O_413,N_2890,N_2868);
nor UO_414 (O_414,N_2875,N_2972);
or UO_415 (O_415,N_2866,N_2853);
nand UO_416 (O_416,N_2874,N_2868);
nand UO_417 (O_417,N_2911,N_2878);
xor UO_418 (O_418,N_2827,N_2937);
or UO_419 (O_419,N_2806,N_2856);
and UO_420 (O_420,N_2824,N_2953);
nor UO_421 (O_421,N_2861,N_2996);
or UO_422 (O_422,N_2827,N_2821);
nor UO_423 (O_423,N_2838,N_2916);
or UO_424 (O_424,N_2914,N_2995);
and UO_425 (O_425,N_2923,N_2870);
nor UO_426 (O_426,N_2887,N_2870);
and UO_427 (O_427,N_2957,N_2861);
nor UO_428 (O_428,N_2831,N_2941);
and UO_429 (O_429,N_2989,N_2880);
xnor UO_430 (O_430,N_2817,N_2946);
xnor UO_431 (O_431,N_2967,N_2921);
nand UO_432 (O_432,N_2815,N_2930);
nor UO_433 (O_433,N_2933,N_2806);
or UO_434 (O_434,N_2984,N_2972);
xor UO_435 (O_435,N_2814,N_2967);
nand UO_436 (O_436,N_2813,N_2881);
and UO_437 (O_437,N_2996,N_2873);
nor UO_438 (O_438,N_2842,N_2868);
nand UO_439 (O_439,N_2979,N_2858);
or UO_440 (O_440,N_2993,N_2942);
nand UO_441 (O_441,N_2953,N_2961);
xor UO_442 (O_442,N_2887,N_2952);
and UO_443 (O_443,N_2822,N_2975);
nand UO_444 (O_444,N_2842,N_2858);
nand UO_445 (O_445,N_2959,N_2809);
or UO_446 (O_446,N_2984,N_2963);
nand UO_447 (O_447,N_2989,N_2936);
or UO_448 (O_448,N_2972,N_2854);
nor UO_449 (O_449,N_2940,N_2885);
and UO_450 (O_450,N_2826,N_2876);
and UO_451 (O_451,N_2900,N_2979);
nand UO_452 (O_452,N_2935,N_2804);
or UO_453 (O_453,N_2987,N_2828);
nor UO_454 (O_454,N_2908,N_2897);
and UO_455 (O_455,N_2927,N_2827);
or UO_456 (O_456,N_2804,N_2919);
and UO_457 (O_457,N_2891,N_2919);
nand UO_458 (O_458,N_2895,N_2830);
nand UO_459 (O_459,N_2965,N_2843);
and UO_460 (O_460,N_2991,N_2860);
nand UO_461 (O_461,N_2922,N_2838);
nor UO_462 (O_462,N_2896,N_2949);
nand UO_463 (O_463,N_2998,N_2903);
nor UO_464 (O_464,N_2824,N_2819);
nand UO_465 (O_465,N_2974,N_2832);
nor UO_466 (O_466,N_2825,N_2920);
nor UO_467 (O_467,N_2894,N_2848);
nand UO_468 (O_468,N_2995,N_2905);
and UO_469 (O_469,N_2997,N_2962);
nand UO_470 (O_470,N_2889,N_2972);
and UO_471 (O_471,N_2943,N_2875);
nor UO_472 (O_472,N_2873,N_2974);
xor UO_473 (O_473,N_2900,N_2830);
nand UO_474 (O_474,N_2975,N_2900);
nand UO_475 (O_475,N_2909,N_2978);
nand UO_476 (O_476,N_2969,N_2870);
nand UO_477 (O_477,N_2914,N_2803);
nor UO_478 (O_478,N_2938,N_2830);
nand UO_479 (O_479,N_2972,N_2827);
or UO_480 (O_480,N_2856,N_2952);
and UO_481 (O_481,N_2997,N_2844);
and UO_482 (O_482,N_2869,N_2864);
xnor UO_483 (O_483,N_2858,N_2887);
nor UO_484 (O_484,N_2993,N_2972);
nand UO_485 (O_485,N_2972,N_2987);
nand UO_486 (O_486,N_2832,N_2839);
nor UO_487 (O_487,N_2907,N_2820);
or UO_488 (O_488,N_2983,N_2873);
nor UO_489 (O_489,N_2885,N_2822);
nor UO_490 (O_490,N_2951,N_2821);
nor UO_491 (O_491,N_2875,N_2958);
or UO_492 (O_492,N_2931,N_2871);
nor UO_493 (O_493,N_2913,N_2990);
or UO_494 (O_494,N_2930,N_2848);
or UO_495 (O_495,N_2872,N_2922);
nor UO_496 (O_496,N_2940,N_2991);
or UO_497 (O_497,N_2983,N_2994);
nand UO_498 (O_498,N_2957,N_2914);
nand UO_499 (O_499,N_2821,N_2957);
endmodule