module basic_1500_15000_2000_50_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_1257,In_69);
nor U1 (N_1,In_763,In_172);
xor U2 (N_2,In_498,In_798);
or U3 (N_3,In_570,In_425);
xor U4 (N_4,In_795,In_484);
nor U5 (N_5,In_326,In_1436);
nand U6 (N_6,In_1241,In_1495);
nand U7 (N_7,In_538,In_292);
xor U8 (N_8,In_879,In_449);
nor U9 (N_9,In_847,In_1156);
xnor U10 (N_10,In_413,In_1008);
or U11 (N_11,In_1045,In_835);
nand U12 (N_12,In_1086,In_286);
nand U13 (N_13,In_1073,In_1012);
nor U14 (N_14,In_350,In_399);
or U15 (N_15,In_1147,In_689);
xnor U16 (N_16,In_625,In_1379);
nor U17 (N_17,In_1101,In_71);
xor U18 (N_18,In_802,In_1102);
and U19 (N_19,In_80,In_132);
or U20 (N_20,In_1234,In_607);
nand U21 (N_21,In_608,In_151);
nand U22 (N_22,In_181,In_1480);
xor U23 (N_23,In_412,In_1233);
xor U24 (N_24,In_336,In_693);
or U25 (N_25,In_78,In_0);
or U26 (N_26,In_444,In_446);
and U27 (N_27,In_964,In_909);
and U28 (N_28,In_300,In_1454);
and U29 (N_29,In_233,In_388);
nand U30 (N_30,In_230,In_772);
and U31 (N_31,In_908,In_1395);
and U32 (N_32,In_176,In_1343);
or U33 (N_33,In_916,In_248);
nor U34 (N_34,In_255,In_59);
or U35 (N_35,In_1449,In_457);
and U36 (N_36,In_1448,In_800);
nor U37 (N_37,In_1238,In_1444);
nor U38 (N_38,In_330,In_1085);
or U39 (N_39,In_1129,In_1410);
nand U40 (N_40,In_976,In_518);
nor U41 (N_41,In_1093,In_384);
nand U42 (N_42,In_1050,In_749);
and U43 (N_43,In_1182,In_488);
nand U44 (N_44,In_673,In_118);
xnor U45 (N_45,In_953,In_219);
and U46 (N_46,In_242,In_373);
nor U47 (N_47,In_1382,In_161);
nand U48 (N_48,In_1419,In_512);
nand U49 (N_49,In_823,In_454);
nor U50 (N_50,In_676,In_77);
nor U51 (N_51,In_23,In_1161);
xnor U52 (N_52,In_808,In_1036);
nand U53 (N_53,In_1431,In_604);
nor U54 (N_54,In_470,In_474);
nand U55 (N_55,In_1385,In_1069);
or U56 (N_56,In_1130,In_787);
nor U57 (N_57,In_790,In_1322);
xnor U58 (N_58,In_825,In_1330);
nand U59 (N_59,In_936,In_641);
xor U60 (N_60,In_244,In_386);
nand U61 (N_61,In_1415,In_1174);
and U62 (N_62,In_647,In_681);
or U63 (N_63,In_258,In_539);
or U64 (N_64,In_812,In_391);
or U65 (N_65,In_682,In_901);
nor U66 (N_66,In_955,In_443);
and U67 (N_67,In_893,In_840);
nor U68 (N_68,In_1004,In_626);
nand U69 (N_69,In_1317,In_349);
nor U70 (N_70,In_1010,In_1024);
or U71 (N_71,In_862,In_1178);
nand U72 (N_72,In_465,In_48);
and U73 (N_73,In_563,In_1397);
nor U74 (N_74,In_369,In_651);
or U75 (N_75,In_536,In_714);
nand U76 (N_76,In_387,In_1294);
nor U77 (N_77,In_528,In_1175);
nand U78 (N_78,In_270,In_1487);
xor U79 (N_79,In_523,In_1357);
xnor U80 (N_80,In_366,In_503);
nor U81 (N_81,In_13,In_169);
and U82 (N_82,In_685,In_1212);
xor U83 (N_83,In_1001,In_707);
and U84 (N_84,In_1398,In_264);
nand U85 (N_85,In_533,In_754);
nand U86 (N_86,In_588,In_302);
nand U87 (N_87,In_586,In_1467);
and U88 (N_88,In_510,In_278);
nor U89 (N_89,In_1099,In_281);
xor U90 (N_90,In_94,In_1181);
or U91 (N_91,In_390,In_1095);
and U92 (N_92,In_111,In_837);
or U93 (N_93,In_917,In_1341);
xnor U94 (N_94,In_1346,In_1263);
nand U95 (N_95,In_476,In_128);
and U96 (N_96,In_485,In_722);
nor U97 (N_97,In_1446,In_757);
xnor U98 (N_98,In_796,In_730);
xnor U99 (N_99,In_1370,In_434);
xor U100 (N_100,In_50,In_271);
xnor U101 (N_101,In_514,In_594);
and U102 (N_102,In_1116,In_260);
xnor U103 (N_103,In_114,In_715);
nand U104 (N_104,In_635,In_502);
nand U105 (N_105,In_110,In_1460);
nand U106 (N_106,In_598,In_634);
xnor U107 (N_107,In_891,In_506);
nor U108 (N_108,In_1076,In_895);
and U109 (N_109,In_938,In_582);
xnor U110 (N_110,In_229,In_605);
xnor U111 (N_111,In_419,In_1319);
or U112 (N_112,In_746,In_1450);
and U113 (N_113,In_195,In_1328);
nor U114 (N_114,In_117,In_1042);
and U115 (N_115,In_564,In_401);
xor U116 (N_116,In_265,In_686);
nor U117 (N_117,In_619,In_1259);
nor U118 (N_118,In_1165,In_257);
xor U119 (N_119,In_1087,In_814);
or U120 (N_120,In_1109,In_1310);
and U121 (N_121,In_717,In_755);
and U122 (N_122,In_876,In_1164);
and U123 (N_123,In_1123,In_791);
or U124 (N_124,In_438,In_324);
xnor U125 (N_125,In_227,In_587);
and U126 (N_126,In_1363,In_88);
xnor U127 (N_127,In_1474,In_656);
nor U128 (N_128,In_750,In_427);
nor U129 (N_129,In_453,In_898);
nand U130 (N_130,In_269,In_308);
or U131 (N_131,In_140,In_252);
nand U132 (N_132,In_241,In_226);
nor U133 (N_133,In_1275,In_989);
nor U134 (N_134,In_663,In_985);
nand U135 (N_135,In_482,In_1268);
nor U136 (N_136,In_534,In_843);
nor U137 (N_137,In_1137,In_896);
nor U138 (N_138,In_68,In_1476);
and U139 (N_139,In_313,In_312);
nor U140 (N_140,In_1336,In_551);
or U141 (N_141,In_1132,In_335);
nor U142 (N_142,In_836,In_452);
or U143 (N_143,In_396,In_273);
nor U144 (N_144,In_553,In_1283);
nand U145 (N_145,In_1272,In_708);
nor U146 (N_146,In_356,In_127);
or U147 (N_147,In_321,In_142);
and U148 (N_148,In_1245,In_1314);
nand U149 (N_149,In_725,In_713);
nand U150 (N_150,In_54,In_674);
and U151 (N_151,In_329,In_462);
and U152 (N_152,In_305,In_93);
nand U153 (N_153,In_801,In_395);
or U154 (N_154,In_952,In_285);
or U155 (N_155,In_737,In_418);
and U156 (N_156,In_747,In_1166);
or U157 (N_157,In_1288,In_1141);
and U158 (N_158,In_609,In_84);
or U159 (N_159,In_1171,In_96);
nand U160 (N_160,In_430,In_1189);
xor U161 (N_161,In_403,In_1145);
and U162 (N_162,In_379,In_1311);
xnor U163 (N_163,In_716,In_112);
nor U164 (N_164,In_1228,In_845);
or U165 (N_165,In_1381,In_466);
nor U166 (N_166,In_779,In_1368);
xor U167 (N_167,In_73,In_1224);
nor U168 (N_168,In_1117,In_1463);
xor U169 (N_169,In_977,In_995);
and U170 (N_170,In_659,In_789);
or U171 (N_171,In_753,In_507);
and U172 (N_172,In_1409,In_939);
or U173 (N_173,In_189,In_188);
nand U174 (N_174,In_495,In_14);
nand U175 (N_175,In_874,In_1389);
nor U176 (N_176,In_639,In_1329);
or U177 (N_177,In_1289,In_1106);
or U178 (N_178,In_643,In_519);
nor U179 (N_179,In_1456,In_1096);
or U180 (N_180,In_556,In_1030);
nand U181 (N_181,In_578,In_775);
xor U182 (N_182,In_199,In_81);
and U183 (N_183,In_1140,In_1038);
xnor U184 (N_184,In_704,In_614);
nand U185 (N_185,In_591,In_149);
nand U186 (N_186,In_618,In_1088);
and U187 (N_187,In_352,In_66);
xor U188 (N_188,In_150,In_1061);
or U189 (N_189,In_832,In_1492);
xnor U190 (N_190,In_1033,In_575);
nand U191 (N_191,In_1218,In_178);
xor U192 (N_192,In_125,In_1425);
nand U193 (N_193,In_692,In_1100);
and U194 (N_194,In_416,In_782);
nor U195 (N_195,In_794,In_1285);
or U196 (N_196,In_670,In_212);
and U197 (N_197,In_831,In_1120);
or U198 (N_198,In_1347,In_1316);
and U199 (N_199,In_1404,In_1458);
nor U200 (N_200,In_839,In_975);
nand U201 (N_201,In_1361,In_1376);
xor U202 (N_202,In_815,In_355);
and U203 (N_203,In_41,In_525);
and U204 (N_204,In_1139,In_475);
or U205 (N_205,In_818,In_1380);
and U206 (N_206,In_1274,In_319);
xor U207 (N_207,In_1249,In_1104);
nor U208 (N_208,In_500,In_709);
nand U209 (N_209,In_239,In_1170);
xor U210 (N_210,In_1269,In_742);
nand U211 (N_211,In_201,In_383);
nor U212 (N_212,In_522,In_1352);
and U213 (N_213,In_906,In_655);
nor U214 (N_214,In_882,In_919);
nand U215 (N_215,In_306,In_788);
and U216 (N_216,In_834,In_268);
and U217 (N_217,In_1442,In_649);
nand U218 (N_218,In_279,In_22);
nor U219 (N_219,In_365,In_1197);
and U220 (N_220,In_496,In_727);
or U221 (N_221,In_345,In_6);
nor U222 (N_222,In_1367,In_1258);
nand U223 (N_223,In_535,In_1348);
or U224 (N_224,In_1437,In_973);
xnor U225 (N_225,In_698,In_147);
or U226 (N_226,In_4,In_943);
xor U227 (N_227,In_728,In_7);
nand U228 (N_228,In_407,In_758);
nor U229 (N_229,In_1133,In_284);
or U230 (N_230,In_833,In_1154);
or U231 (N_231,In_348,In_912);
xnor U232 (N_232,In_610,In_543);
xor U233 (N_233,In_1159,In_364);
and U234 (N_234,In_826,In_1220);
nand U235 (N_235,In_211,In_1342);
nand U236 (N_236,In_1060,In_422);
or U237 (N_237,In_504,In_1411);
or U238 (N_238,In_1453,In_1452);
nor U239 (N_239,In_338,In_1253);
xor U240 (N_240,In_424,In_1119);
or U241 (N_241,In_1455,In_1215);
or U242 (N_242,In_561,In_1021);
or U243 (N_243,In_409,In_163);
xor U244 (N_244,In_1282,In_940);
xor U245 (N_245,In_8,In_283);
nor U246 (N_246,In_203,In_1468);
and U247 (N_247,In_771,In_1418);
nand U248 (N_248,In_380,In_932);
nand U249 (N_249,In_1185,In_1052);
or U250 (N_250,In_417,In_571);
nand U251 (N_251,In_810,In_861);
nor U252 (N_252,In_5,In_648);
xnor U253 (N_253,In_1127,In_1051);
nand U254 (N_254,In_961,In_696);
nand U255 (N_255,In_972,In_852);
or U256 (N_256,In_328,In_342);
nor U257 (N_257,In_90,In_694);
xnor U258 (N_258,In_947,In_56);
or U259 (N_259,In_723,In_1040);
nand U260 (N_260,In_527,In_145);
nand U261 (N_261,In_867,In_954);
and U262 (N_262,In_235,In_1375);
xnor U263 (N_263,In_565,In_1135);
xor U264 (N_264,In_1313,In_339);
nand U265 (N_265,In_645,In_1445);
xnor U266 (N_266,In_942,In_785);
and U267 (N_267,In_773,In_115);
nand U268 (N_268,In_1094,In_202);
nor U269 (N_269,In_253,In_585);
and U270 (N_270,In_472,In_180);
and U271 (N_271,In_95,In_1018);
nand U272 (N_272,In_16,In_17);
xnor U273 (N_273,In_1320,In_559);
or U274 (N_274,In_1183,In_259);
and U275 (N_275,In_478,In_318);
nand U276 (N_276,In_1110,In_983);
xor U277 (N_277,In_894,In_1190);
or U278 (N_278,In_1150,In_662);
or U279 (N_279,In_45,In_860);
xor U280 (N_280,In_516,In_293);
nor U281 (N_281,In_397,In_873);
nor U282 (N_282,In_376,In_1136);
and U283 (N_283,In_375,In_428);
nand U284 (N_284,In_589,In_654);
or U285 (N_285,In_385,In_680);
and U286 (N_286,In_137,In_524);
nand U287 (N_287,In_930,In_851);
xnor U288 (N_288,In_592,In_666);
nor U289 (N_289,In_1002,In_1200);
nand U290 (N_290,In_629,In_1429);
nand U291 (N_291,In_381,In_144);
or U292 (N_292,In_1432,In_617);
or U293 (N_293,In_344,In_710);
nor U294 (N_294,In_471,In_751);
or U295 (N_295,In_36,In_568);
xnor U296 (N_296,In_492,In_827);
or U297 (N_297,In_1196,In_351);
and U298 (N_298,In_892,In_1155);
nor U299 (N_299,In_1325,In_1488);
xnor U300 (N_300,In_1303,In_911);
or U301 (N_301,In_1058,In_1198);
and U302 (N_302,N_74,In_872);
and U303 (N_303,In_1401,In_389);
xnor U304 (N_304,In_208,In_148);
nor U305 (N_305,In_764,In_1118);
nand U306 (N_306,In_346,N_104);
nand U307 (N_307,N_155,In_703);
xor U308 (N_308,In_200,In_455);
or U309 (N_309,N_269,In_613);
or U310 (N_310,In_1273,In_623);
or U311 (N_311,N_60,N_190);
nand U312 (N_312,In_549,In_711);
and U313 (N_313,In_573,In_1406);
and U314 (N_314,In_797,N_135);
nand U315 (N_315,In_38,In_1078);
or U316 (N_316,In_1459,In_1089);
xnor U317 (N_317,N_27,N_242);
or U318 (N_318,In_1423,N_230);
or U319 (N_319,In_256,In_1235);
nand U320 (N_320,In_327,In_433);
xnor U321 (N_321,In_473,N_258);
nand U322 (N_322,In_205,In_915);
nor U323 (N_323,N_195,In_738);
or U324 (N_324,In_40,N_28);
nand U325 (N_325,In_1478,In_1337);
nand U326 (N_326,In_621,N_96);
nor U327 (N_327,N_194,In_1434);
xor U328 (N_328,In_245,In_1248);
nor U329 (N_329,In_545,In_1338);
or U330 (N_330,In_60,In_1428);
or U331 (N_331,In_1278,In_1365);
xor U332 (N_332,In_695,In_875);
and U333 (N_333,In_931,In_1121);
nand U334 (N_334,In_1063,In_899);
or U335 (N_335,In_999,In_101);
and U336 (N_336,In_544,In_1022);
and U337 (N_337,In_170,In_1219);
or U338 (N_338,N_247,N_113);
or U339 (N_339,In_334,In_741);
nand U340 (N_340,N_46,N_47);
nor U341 (N_341,In_864,In_405);
xor U342 (N_342,N_265,In_1353);
or U343 (N_343,In_432,In_431);
or U344 (N_344,In_679,In_1494);
nor U345 (N_345,In_234,In_646);
xnor U346 (N_346,N_131,In_547);
nand U347 (N_347,N_156,In_1312);
nor U348 (N_348,In_370,In_51);
nand U349 (N_349,In_542,In_190);
nand U350 (N_350,In_1202,N_215);
or U351 (N_351,In_765,In_1451);
xor U352 (N_352,In_804,In_841);
and U353 (N_353,In_450,In_1373);
nand U354 (N_354,In_177,In_274);
xnor U355 (N_355,In_672,In_290);
xor U356 (N_356,In_108,In_770);
or U357 (N_357,N_173,N_102);
nand U358 (N_358,In_706,N_226);
or U359 (N_359,In_85,In_499);
and U360 (N_360,N_14,N_151);
and U361 (N_361,N_43,In_530);
nand U362 (N_362,In_1037,In_98);
nand U363 (N_363,In_687,In_291);
xor U364 (N_364,N_207,In_984);
and U365 (N_365,N_216,In_167);
or U366 (N_366,N_177,In_1225);
xor U367 (N_367,N_280,In_1262);
nand U368 (N_368,In_567,N_277);
xnor U369 (N_369,In_844,In_1394);
xor U370 (N_370,In_1019,N_183);
xor U371 (N_371,N_134,In_1015);
or U372 (N_372,In_353,In_632);
and U373 (N_373,In_1149,N_111);
nor U374 (N_374,In_640,In_1465);
nor U375 (N_375,In_581,In_941);
nand U376 (N_376,In_237,In_1205);
nor U377 (N_377,In_1059,In_529);
or U378 (N_378,In_1240,N_70);
or U379 (N_379,In_1413,N_110);
nand U380 (N_380,In_1482,N_236);
nand U381 (N_381,In_1206,In_799);
nand U382 (N_382,N_241,In_1359);
or U383 (N_383,In_669,N_148);
or U384 (N_384,In_143,In_1195);
and U385 (N_385,In_821,In_1261);
and U386 (N_386,In_220,In_842);
and U387 (N_387,In_266,In_631);
xnor U388 (N_388,In_988,In_74);
or U389 (N_389,In_691,In_323);
nor U390 (N_390,In_562,In_951);
or U391 (N_391,In_904,In_849);
or U392 (N_392,In_209,In_521);
and U393 (N_393,In_331,In_358);
nor U394 (N_394,In_236,N_120);
xnor U395 (N_395,In_119,N_7);
nor U396 (N_396,N_15,N_72);
or U397 (N_397,In_574,N_145);
nand U398 (N_398,In_1390,In_122);
xor U399 (N_399,In_1481,In_1080);
nand U400 (N_400,N_39,N_33);
or U401 (N_401,In_310,In_949);
nand U402 (N_402,In_1326,In_620);
nor U403 (N_403,In_1281,N_117);
and U404 (N_404,In_1499,In_925);
xnor U405 (N_405,In_1469,In_1180);
or U406 (N_406,In_1247,N_142);
xor U407 (N_407,In_566,In_3);
xor U408 (N_408,N_119,In_1386);
or U409 (N_409,In_1270,N_167);
or U410 (N_410,In_155,In_67);
xor U411 (N_411,In_314,In_572);
or U412 (N_412,N_23,In_540);
xnor U413 (N_413,In_158,N_146);
xor U414 (N_414,N_246,In_905);
nor U415 (N_415,In_1286,N_138);
xor U416 (N_416,In_107,In_813);
and U417 (N_417,In_1470,In_637);
or U418 (N_418,In_79,In_1324);
nor U419 (N_419,In_287,In_1340);
nor U420 (N_420,In_1304,In_333);
and U421 (N_421,In_865,In_1188);
nor U422 (N_422,N_103,In_1177);
and U423 (N_423,N_31,In_126);
nor U424 (N_424,In_1114,In_732);
and U425 (N_425,In_1296,N_214);
nand U426 (N_426,N_271,In_1256);
or U427 (N_427,In_809,In_340);
xnor U428 (N_428,In_1242,N_80);
or U429 (N_429,In_1366,In_250);
or U430 (N_430,In_1387,In_304);
nor U431 (N_431,In_44,N_181);
nor U432 (N_432,In_885,N_57);
and U433 (N_433,In_690,In_400);
or U434 (N_434,N_91,In_596);
nor U435 (N_435,In_1143,In_548);
nor U436 (N_436,In_1062,In_214);
nor U437 (N_437,In_213,In_1392);
and U438 (N_438,In_776,In_30);
and U439 (N_439,In_661,In_817);
xor U440 (N_440,N_164,In_166);
and U441 (N_441,N_55,In_426);
and U442 (N_442,In_301,In_783);
xor U443 (N_443,In_828,In_1077);
xor U444 (N_444,N_232,N_196);
xnor U445 (N_445,In_394,In_962);
and U446 (N_446,In_152,In_981);
nand U447 (N_447,N_185,In_322);
or U448 (N_448,N_275,In_429);
xnor U449 (N_449,In_766,In_857);
xor U450 (N_450,N_82,N_253);
or U451 (N_451,In_660,N_254);
nand U452 (N_452,In_1108,In_251);
and U453 (N_453,In_1276,In_1351);
nor U454 (N_454,In_109,In_719);
or U455 (N_455,In_929,In_246);
xor U456 (N_456,N_235,In_1230);
or U457 (N_457,In_1491,In_91);
and U458 (N_458,In_1345,In_1280);
or U459 (N_459,In_1067,In_1407);
nand U460 (N_460,In_1414,In_1138);
xor U461 (N_461,N_152,In_900);
and U462 (N_462,N_9,In_1057);
xnor U463 (N_463,In_531,In_1157);
or U464 (N_464,In_1302,In_1405);
nand U465 (N_465,In_97,In_1321);
nor U466 (N_466,N_95,In_1493);
nor U467 (N_467,In_458,In_1065);
nand U468 (N_468,In_683,N_58);
nand U469 (N_469,In_1403,In_697);
nor U470 (N_470,N_282,N_288);
and U471 (N_471,In_467,N_250);
nand U472 (N_472,In_218,In_1292);
xor U473 (N_473,In_558,In_459);
nor U474 (N_474,In_910,In_731);
and U475 (N_475,In_793,In_1284);
and U476 (N_476,In_1462,N_67);
or U477 (N_477,In_990,In_1243);
xor U478 (N_478,In_511,In_299);
or U479 (N_479,In_374,In_658);
nor U480 (N_480,In_806,In_1232);
xnor U481 (N_481,N_175,In_602);
or U482 (N_482,In_935,In_440);
or U483 (N_483,In_890,In_371);
nand U484 (N_484,N_127,In_830);
xnor U485 (N_485,In_1227,In_688);
nor U486 (N_486,In_675,N_83);
xor U487 (N_487,In_33,In_2);
nor U488 (N_488,N_218,In_480);
and U489 (N_489,N_182,In_1013);
xnor U490 (N_490,In_89,In_24);
and U491 (N_491,In_684,In_1162);
nand U492 (N_492,In_295,In_1327);
nor U493 (N_493,In_856,In_1246);
xor U494 (N_494,In_1301,In_1017);
xnor U495 (N_495,N_30,In_436);
xnor U496 (N_496,In_1186,In_1029);
nand U497 (N_497,In_792,In_616);
xnor U498 (N_498,In_414,N_56);
nor U499 (N_499,N_294,N_249);
or U500 (N_500,In_924,In_720);
or U501 (N_501,In_1124,N_211);
or U502 (N_502,In_555,In_958);
and U503 (N_503,In_316,In_886);
xnor U504 (N_504,N_123,In_421);
nor U505 (N_505,In_934,In_1318);
nand U506 (N_506,In_878,In_311);
and U507 (N_507,In_37,In_1092);
and U508 (N_508,N_228,In_1041);
or U509 (N_509,N_61,N_34);
or U510 (N_510,In_28,In_223);
xor U511 (N_511,In_508,N_8);
and U512 (N_512,N_264,In_1027);
nand U513 (N_513,In_597,In_1128);
xnor U514 (N_514,In_1354,In_638);
nand U515 (N_515,N_150,N_272);
or U516 (N_516,In_146,In_1417);
nor U517 (N_517,In_1176,In_1028);
or U518 (N_518,In_1194,N_2);
nand U519 (N_519,In_667,In_721);
xor U520 (N_520,N_179,In_206);
and U521 (N_521,In_702,In_194);
nor U522 (N_522,In_991,In_970);
nor U523 (N_523,In_652,N_36);
nand U524 (N_524,In_367,In_282);
nor U525 (N_525,In_1421,N_71);
and U526 (N_526,In_52,N_42);
nand U527 (N_527,In_859,In_665);
nand U528 (N_528,In_1412,N_212);
nor U529 (N_529,N_1,In_998);
and U530 (N_530,In_1356,In_11);
nand U531 (N_531,In_185,N_126);
or U532 (N_532,In_1362,N_237);
nand U533 (N_533,In_959,In_1107);
or U534 (N_534,In_1221,N_136);
or U535 (N_535,In_1371,In_729);
and U536 (N_536,In_541,In_1231);
nand U537 (N_537,N_193,N_22);
nand U538 (N_538,In_1360,In_249);
nand U539 (N_539,In_70,In_994);
and U540 (N_540,In_1323,N_180);
nand U541 (N_541,N_251,N_125);
nand U542 (N_542,In_778,N_229);
nand U543 (N_543,In_969,In_1298);
and U544 (N_544,In_599,In_1184);
nand U545 (N_545,In_131,In_1169);
or U546 (N_546,In_1393,In_343);
and U547 (N_547,In_442,In_838);
nand U548 (N_548,In_19,N_203);
nor U549 (N_549,N_144,In_1031);
nand U550 (N_550,In_739,In_113);
or U551 (N_551,In_577,N_18);
nand U552 (N_552,In_784,In_1430);
and U553 (N_553,In_486,In_846);
or U554 (N_554,In_341,N_92);
nor U555 (N_555,N_243,N_105);
nor U556 (N_556,In_767,In_1307);
nand U557 (N_557,N_44,N_132);
xnor U558 (N_558,In_1016,In_58);
nand U559 (N_559,N_192,N_293);
and U560 (N_560,In_848,N_141);
or U561 (N_561,N_159,In_829);
nand U562 (N_562,N_163,In_32);
or U563 (N_563,In_398,In_769);
or U564 (N_564,In_337,In_923);
and U565 (N_565,In_464,In_1193);
and U566 (N_566,In_858,In_967);
nor U567 (N_567,In_65,In_1433);
and U568 (N_568,N_154,In_1032);
and U569 (N_569,N_32,In_277);
nor U570 (N_570,In_483,In_1152);
nand U571 (N_571,In_595,In_10);
nand U572 (N_572,In_76,In_1374);
or U573 (N_573,N_130,N_40);
xnor U574 (N_574,In_628,In_781);
and U575 (N_575,N_0,In_1372);
and U576 (N_576,In_1277,In_1112);
and U577 (N_577,In_406,In_1427);
and U578 (N_578,In_15,In_477);
nand U579 (N_579,In_12,N_238);
xor U580 (N_580,In_996,In_197);
nand U581 (N_581,In_854,N_133);
or U582 (N_582,In_497,In_204);
and U583 (N_583,In_1204,N_205);
nor U584 (N_584,N_107,In_1475);
xnor U585 (N_585,In_468,In_1383);
nand U586 (N_586,In_82,In_807);
or U587 (N_587,N_78,In_238);
xor U588 (N_588,In_1334,In_263);
or U589 (N_589,N_77,In_920);
nand U590 (N_590,In_26,In_1229);
nand U591 (N_591,In_1034,In_1199);
or U592 (N_592,N_279,In_46);
nor U593 (N_593,In_678,In_913);
or U594 (N_594,In_974,N_172);
or U595 (N_595,In_756,In_1264);
or U596 (N_596,In_1167,In_966);
or U597 (N_597,In_1213,In_701);
or U598 (N_598,N_101,In_1293);
nor U599 (N_599,N_62,In_183);
nor U600 (N_600,In_1447,In_1300);
xor U601 (N_601,In_39,N_479);
xor U602 (N_602,In_1146,In_887);
nand U603 (N_603,In_1011,N_198);
or U604 (N_604,N_415,In_883);
nor U605 (N_605,N_301,N_116);
xnor U606 (N_606,In_1126,In_718);
nand U607 (N_607,In_105,N_583);
nand U608 (N_608,In_410,N_485);
nor U609 (N_609,In_1006,In_1217);
or U610 (N_610,In_1291,In_1489);
xor U611 (N_611,In_1265,In_1111);
nand U612 (N_612,N_477,In_103);
xor U613 (N_613,N_295,N_309);
or U614 (N_614,N_303,N_423);
and U615 (N_615,N_115,N_576);
nand U616 (N_616,In_552,In_871);
nor U617 (N_617,In_86,In_992);
xor U618 (N_618,N_586,N_300);
and U619 (N_619,In_42,In_160);
nand U620 (N_620,N_65,N_86);
nor U621 (N_621,N_387,In_642);
nor U622 (N_622,In_853,In_490);
xnor U623 (N_623,In_135,N_526);
nand U624 (N_624,N_171,N_376);
or U625 (N_625,N_455,N_347);
and U626 (N_626,In_650,N_377);
nor U627 (N_627,N_231,In_1074);
xor U628 (N_628,In_83,N_45);
nor U629 (N_629,N_529,N_370);
nor U630 (N_630,In_130,N_561);
and U631 (N_631,N_574,N_436);
and U632 (N_632,N_286,In_1483);
and U633 (N_633,N_433,In_903);
and U634 (N_634,In_1399,In_171);
xnor U635 (N_635,In_487,N_284);
nand U636 (N_636,N_499,In_134);
and U637 (N_637,In_415,In_590);
and U638 (N_638,N_447,N_197);
and U639 (N_639,N_558,In_120);
and U640 (N_640,In_554,N_496);
nand U641 (N_641,N_474,In_1055);
xor U642 (N_642,N_397,In_382);
or U643 (N_643,In_57,N_542);
xnor U644 (N_644,In_816,In_1142);
nor U645 (N_645,N_350,In_1009);
nor U646 (N_646,In_517,In_997);
or U647 (N_647,In_580,N_311);
and U648 (N_648,N_245,N_490);
and U649 (N_649,In_1158,In_956);
nor U650 (N_650,In_1237,In_532);
or U651 (N_651,N_210,In_1426);
or U652 (N_652,N_458,In_1250);
xor U653 (N_653,N_128,In_489);
nor U654 (N_654,In_1440,N_352);
and U655 (N_655,In_786,N_502);
or U656 (N_656,N_188,N_153);
or U657 (N_657,In_863,N_590);
nand U658 (N_658,In_191,N_52);
and U659 (N_659,In_215,In_1072);
or U660 (N_660,In_420,In_1223);
nor U661 (N_661,In_1295,N_491);
and U662 (N_662,N_430,N_261);
nand U663 (N_663,N_596,N_339);
nand U664 (N_664,N_266,In_154);
xor U665 (N_665,In_1484,N_332);
and U666 (N_666,N_262,N_354);
nand U667 (N_667,N_140,N_362);
xnor U668 (N_668,In_121,In_393);
xnor U669 (N_669,In_1103,In_907);
or U670 (N_670,In_1244,In_1201);
nor U671 (N_671,In_877,N_298);
nor U672 (N_672,In_1000,N_308);
nor U673 (N_673,In_445,In_978);
nand U674 (N_674,N_554,N_404);
and U675 (N_675,In_1064,N_438);
xnor U676 (N_676,In_1306,In_1408);
and U677 (N_677,In_884,N_76);
or U678 (N_678,N_21,N_533);
xnor U679 (N_679,N_158,In_933);
xor U680 (N_680,In_627,N_324);
and U681 (N_681,N_396,In_957);
nand U682 (N_682,In_1115,N_444);
or U683 (N_683,In_1441,In_243);
or U684 (N_684,N_505,In_272);
nor U685 (N_685,In_902,In_179);
and U686 (N_686,In_937,In_636);
and U687 (N_687,In_493,In_34);
and U688 (N_688,N_544,In_743);
xor U689 (N_689,In_1279,N_165);
nor U690 (N_690,N_336,In_1416);
and U691 (N_691,N_368,In_1222);
nor U692 (N_692,N_375,N_79);
nor U693 (N_693,In_579,N_472);
nor U694 (N_694,In_1497,N_147);
nand U695 (N_695,N_456,N_522);
nor U696 (N_696,In_61,N_527);
and U697 (N_697,N_547,In_193);
and U698 (N_698,N_568,N_318);
or U699 (N_699,In_240,In_262);
xor U700 (N_700,In_1191,In_404);
xnor U701 (N_701,In_437,In_133);
xor U702 (N_702,N_537,In_1466);
nand U703 (N_703,N_276,In_21);
nand U704 (N_704,In_777,In_173);
xnor U705 (N_705,In_736,In_569);
or U706 (N_706,In_980,In_1486);
nor U707 (N_707,N_516,N_338);
or U708 (N_708,N_199,N_98);
and U709 (N_709,N_334,N_97);
and U710 (N_710,In_479,In_1496);
nor U711 (N_711,N_285,N_89);
xnor U712 (N_712,In_1349,N_509);
nand U713 (N_713,In_1267,N_10);
xor U714 (N_714,N_90,In_228);
or U715 (N_715,N_240,N_220);
nor U716 (N_716,In_1091,In_805);
or U717 (N_717,N_143,N_12);
nand U718 (N_718,In_27,In_1333);
or U719 (N_719,N_442,N_552);
and U720 (N_720,N_316,N_457);
and U721 (N_721,N_227,In_124);
xnor U722 (N_722,N_528,In_733);
nor U723 (N_723,In_1255,In_1043);
nor U724 (N_724,In_803,N_248);
or U725 (N_725,N_588,N_422);
nor U726 (N_726,In_881,In_1023);
and U727 (N_727,In_1378,N_428);
nand U728 (N_728,In_889,N_88);
or U729 (N_729,In_1020,N_593);
and U730 (N_730,N_466,N_584);
or U731 (N_731,N_26,In_1097);
or U732 (N_732,N_287,In_320);
nor U733 (N_733,N_359,In_198);
nor U734 (N_734,In_1039,In_439);
xnor U735 (N_735,N_340,In_950);
and U736 (N_736,N_538,N_297);
nor U737 (N_737,In_1350,N_383);
or U738 (N_738,N_333,N_478);
nor U739 (N_739,In_1208,N_35);
or U740 (N_740,In_63,In_501);
nand U741 (N_741,In_748,N_506);
or U742 (N_742,N_186,N_380);
nand U743 (N_743,In_1046,N_233);
nand U744 (N_744,N_160,N_384);
nand U745 (N_745,N_418,In_761);
nor U746 (N_746,In_1025,N_99);
nor U747 (N_747,In_1260,In_232);
or U748 (N_748,In_207,In_354);
and U749 (N_749,N_461,In_762);
nand U750 (N_750,In_1490,In_136);
nand U751 (N_751,N_393,In_986);
and U752 (N_752,N_551,In_1083);
and U753 (N_753,N_508,In_515);
nand U754 (N_754,In_123,In_35);
or U755 (N_755,In_408,N_577);
xnor U756 (N_756,N_365,N_412);
xnor U757 (N_757,In_1007,N_589);
nor U758 (N_758,N_459,In_469);
and U759 (N_759,In_948,N_501);
or U760 (N_760,In_1344,N_470);
nand U761 (N_761,In_402,N_304);
or U762 (N_762,N_392,In_159);
and U763 (N_763,In_1400,N_571);
nor U764 (N_764,N_201,N_11);
and U765 (N_765,In_196,N_585);
xnor U766 (N_766,In_1168,In_1236);
nand U767 (N_767,In_1214,In_1090);
nand U768 (N_768,In_156,In_25);
nor U769 (N_769,N_524,In_921);
nor U770 (N_770,N_566,In_315);
xnor U771 (N_771,N_471,N_575);
nand U772 (N_772,In_1335,In_744);
nor U773 (N_773,N_513,In_378);
or U774 (N_774,In_1438,N_222);
xnor U775 (N_775,In_1035,N_108);
or U776 (N_776,In_460,N_530);
nand U777 (N_777,In_1439,N_379);
or U778 (N_778,In_1498,N_323);
xor U779 (N_779,N_582,N_578);
xor U780 (N_780,N_356,In_922);
or U781 (N_781,In_116,N_268);
and U782 (N_782,In_1266,In_1239);
or U783 (N_783,N_217,N_515);
or U784 (N_784,N_398,In_1369);
nand U785 (N_785,In_868,In_1014);
nor U786 (N_786,N_5,N_520);
xor U787 (N_787,N_555,N_382);
nor U788 (N_788,N_451,N_389);
or U789 (N_789,In_1420,In_824);
or U790 (N_790,In_9,In_1);
or U791 (N_791,N_480,In_1210);
nand U792 (N_792,N_489,N_413);
nor U793 (N_793,N_407,N_346);
nand U794 (N_794,In_780,N_435);
nand U795 (N_795,N_353,In_92);
or U796 (N_796,In_222,In_576);
nand U797 (N_797,In_624,N_419);
or U798 (N_798,N_208,N_579);
nand U799 (N_799,N_426,In_700);
or U800 (N_800,In_537,N_511);
or U801 (N_801,N_20,N_410);
nand U802 (N_802,In_1443,N_361);
and U803 (N_803,In_1355,In_162);
xor U804 (N_804,N_441,N_341);
nand U805 (N_805,In_72,N_209);
nand U806 (N_806,N_567,In_165);
xnor U807 (N_807,N_112,In_254);
xnor U808 (N_808,In_494,N_87);
and U809 (N_809,N_325,In_280);
or U810 (N_810,In_64,N_189);
xor U811 (N_811,In_1377,N_168);
nor U812 (N_812,N_521,N_437);
and U813 (N_813,In_1464,In_368);
nor U814 (N_814,N_469,N_349);
xnor U815 (N_815,In_971,In_448);
nor U816 (N_816,N_570,In_275);
xor U817 (N_817,In_435,In_1098);
and U818 (N_818,N_409,N_114);
and U819 (N_819,N_307,In_735);
and U820 (N_820,In_1187,In_47);
nand U821 (N_821,N_344,In_360);
or U822 (N_822,N_19,In_1287);
nand U823 (N_823,N_306,In_1254);
or U824 (N_824,In_153,N_273);
and U825 (N_825,N_532,In_317);
xor U826 (N_826,In_1315,In_657);
or U827 (N_827,N_59,In_1391);
nor U828 (N_828,In_1422,N_518);
nor U829 (N_829,In_593,N_595);
nand U830 (N_830,N_274,N_594);
or U831 (N_831,N_432,In_584);
nand U832 (N_832,In_461,In_1079);
and U833 (N_833,In_1457,In_768);
and U834 (N_834,N_68,In_601);
nor U835 (N_835,N_371,In_1435);
xor U836 (N_836,N_504,N_507);
nor U837 (N_837,N_494,In_1048);
and U838 (N_838,In_357,N_374);
nand U839 (N_839,N_270,N_473);
and U840 (N_840,N_400,In_49);
nor U841 (N_841,N_260,N_395);
and U842 (N_842,N_257,N_93);
nor U843 (N_843,N_66,N_424);
and U844 (N_844,In_926,N_176);
xnor U845 (N_845,N_452,N_394);
or U846 (N_846,In_164,N_481);
xor U847 (N_847,N_427,In_611);
and U848 (N_848,In_1207,N_16);
xor U849 (N_849,In_644,N_124);
or U850 (N_850,N_321,In_1290);
nor U851 (N_851,In_1125,In_946);
xor U852 (N_852,In_129,N_543);
and U853 (N_853,In_87,In_1160);
or U854 (N_854,In_192,In_267);
xnor U855 (N_855,In_441,In_392);
or U856 (N_856,N_355,N_534);
xnor U857 (N_857,In_1251,N_557);
or U858 (N_858,N_391,In_1331);
xor U859 (N_859,N_364,In_759);
or U860 (N_860,N_373,N_525);
xnor U861 (N_861,N_302,N_580);
and U862 (N_862,In_1473,In_372);
or U863 (N_863,N_581,In_968);
xor U864 (N_864,In_622,In_752);
or U865 (N_865,N_434,N_514);
and U866 (N_866,In_1364,In_1131);
nor U867 (N_867,N_37,In_927);
or U868 (N_868,N_483,In_1332);
and U869 (N_869,N_255,In_1384);
and U870 (N_870,N_367,N_283);
nand U871 (N_871,In_18,In_1005);
and U872 (N_872,N_545,N_549);
nor U873 (N_873,In_456,N_462);
nand U874 (N_874,In_855,In_276);
xor U875 (N_875,In_224,In_822);
and U876 (N_876,In_918,In_1216);
nor U877 (N_877,N_17,In_99);
xor U878 (N_878,N_331,N_573);
nor U879 (N_879,N_546,In_210);
nand U880 (N_880,N_417,In_993);
nand U881 (N_881,In_1054,In_982);
nor U882 (N_882,N_224,In_216);
xnor U883 (N_883,N_406,In_309);
nor U884 (N_884,In_653,In_481);
nand U885 (N_885,In_1172,N_291);
nor U886 (N_886,In_1388,In_361);
xor U887 (N_887,N_157,N_4);
and U888 (N_888,In_712,N_169);
nor U889 (N_889,N_326,N_244);
and U890 (N_890,In_1084,N_358);
and U891 (N_891,In_819,N_357);
or U892 (N_892,In_1026,In_106);
or U893 (N_893,N_263,N_386);
and U894 (N_894,N_223,In_1144);
nand U895 (N_895,N_360,N_421);
or U896 (N_896,In_362,In_1081);
xor U897 (N_897,In_1082,N_497);
nor U898 (N_898,N_317,N_492);
and U899 (N_899,N_64,N_445);
or U900 (N_900,N_343,N_337);
nor U901 (N_901,In_677,In_557);
nand U902 (N_902,N_822,N_663);
nor U903 (N_903,N_314,N_899);
xnor U904 (N_904,N_764,In_75);
and U905 (N_905,N_722,N_801);
nand U906 (N_906,N_841,N_863);
xor U907 (N_907,N_603,N_684);
and U908 (N_908,In_55,In_944);
and U909 (N_909,N_829,N_772);
xnor U910 (N_910,In_1192,N_896);
nand U911 (N_911,In_724,N_850);
and U912 (N_912,N_493,N_882);
nor U913 (N_913,N_744,N_797);
xor U914 (N_914,N_655,N_765);
xor U915 (N_915,N_741,N_870);
nand U916 (N_916,N_742,N_674);
nor U917 (N_917,N_675,N_756);
nor U918 (N_918,N_75,N_363);
or U919 (N_919,N_618,N_219);
or U920 (N_920,N_548,N_840);
nor U921 (N_921,N_789,N_845);
nor U922 (N_922,In_1226,N_673);
and U923 (N_923,N_487,In_307);
and U924 (N_924,In_174,In_1305);
xnor U925 (N_925,In_62,N_783);
nand U926 (N_926,In_296,N_745);
nand U927 (N_927,N_833,N_642);
nor U928 (N_928,N_166,N_69);
nor U929 (N_929,N_625,N_616);
and U930 (N_930,N_627,N_500);
nand U931 (N_931,N_751,In_671);
or U932 (N_932,N_556,In_820);
or U933 (N_933,N_335,N_289);
xor U934 (N_934,In_1479,In_247);
nor U935 (N_935,N_329,N_685);
nor U936 (N_936,N_414,N_846);
and U937 (N_937,N_401,N_869);
xnor U938 (N_938,N_564,N_785);
nor U939 (N_939,N_611,In_1105);
or U940 (N_940,N_867,In_1309);
or U941 (N_941,N_718,N_750);
or U942 (N_942,N_702,N_443);
xor U943 (N_943,N_884,In_1068);
or U944 (N_944,N_697,N_440);
nand U945 (N_945,N_784,N_823);
nor U946 (N_946,In_1153,In_550);
nand U947 (N_947,N_777,N_752);
and U948 (N_948,N_319,In_1047);
nor U949 (N_949,N_835,N_687);
nor U950 (N_950,N_615,N_234);
xnor U951 (N_951,N_861,N_898);
or U952 (N_952,N_312,N_626);
or U953 (N_953,N_680,N_631);
nand U954 (N_954,N_369,N_877);
and U955 (N_955,N_184,N_681);
nand U956 (N_956,N_420,N_715);
or U957 (N_957,N_820,N_106);
nand U958 (N_958,N_121,N_623);
xor U959 (N_959,In_217,N_811);
xnor U960 (N_960,N_629,N_607);
nor U961 (N_961,In_411,N_503);
nor U962 (N_962,N_672,N_688);
or U963 (N_963,N_149,N_791);
nor U964 (N_964,N_239,In_104);
nand U965 (N_965,In_325,N_605);
xnor U966 (N_966,In_546,N_894);
or U967 (N_967,N_747,In_633);
xor U968 (N_968,N_644,N_664);
nand U969 (N_969,N_512,N_812);
or U970 (N_970,N_854,In_513);
nor U971 (N_971,In_1339,N_843);
nor U972 (N_972,N_740,In_447);
xnor U973 (N_973,N_837,In_1472);
nand U974 (N_974,N_880,N_206);
or U975 (N_975,In_509,In_1053);
or U976 (N_976,N_608,N_617);
nand U977 (N_977,N_572,N_178);
xnor U978 (N_978,N_599,N_453);
nand U979 (N_979,N_719,N_731);
nand U980 (N_980,N_63,N_893);
nand U981 (N_981,In_583,N_191);
and U982 (N_982,In_1044,N_597);
xnor U983 (N_983,N_723,N_844);
nand U984 (N_984,N_738,In_1271);
or U985 (N_985,N_310,N_888);
nand U986 (N_986,N_768,N_773);
or U987 (N_987,N_460,N_6);
and U988 (N_988,In_774,N_818);
nand U989 (N_989,N_29,N_842);
or U990 (N_990,In_31,N_776);
and U991 (N_991,N_536,N_531);
xnor U992 (N_992,N_775,N_299);
and U993 (N_993,In_1056,N_849);
nand U994 (N_994,N_798,N_292);
and U995 (N_995,N_25,N_620);
and U996 (N_996,N_523,In_221);
or U997 (N_997,N_799,N_665);
nand U998 (N_998,N_320,N_656);
nand U999 (N_999,N_637,N_633);
and U1000 (N_1000,N_628,N_848);
nand U1001 (N_1001,N_488,N_614);
and U1002 (N_1002,N_692,N_780);
nand U1003 (N_1003,N_475,In_914);
and U1004 (N_1004,N_710,N_847);
xnor U1005 (N_1005,N_225,N_743);
nor U1006 (N_1006,In_1151,In_29);
or U1007 (N_1007,N_660,N_385);
xor U1008 (N_1008,N_602,In_463);
or U1009 (N_1009,In_175,N_735);
nor U1010 (N_1010,N_711,In_1122);
or U1011 (N_1011,N_351,N_468);
or U1012 (N_1012,N_803,In_184);
or U1013 (N_1013,N_598,N_495);
nor U1014 (N_1014,N_94,N_290);
xor U1015 (N_1015,N_305,In_866);
nand U1016 (N_1016,In_987,In_734);
or U1017 (N_1017,N_454,N_759);
nor U1018 (N_1018,N_781,N_476);
xnor U1019 (N_1019,N_643,N_405);
or U1020 (N_1020,N_486,In_603);
and U1021 (N_1021,N_795,N_832);
or U1022 (N_1022,In_1070,N_563);
or U1023 (N_1023,N_885,In_43);
or U1024 (N_1024,In_760,N_221);
xor U1025 (N_1025,In_699,N_640);
xnor U1026 (N_1026,N_827,N_624);
or U1027 (N_1027,N_786,N_313);
and U1028 (N_1028,N_484,N_402);
nor U1029 (N_1029,N_638,In_141);
nand U1030 (N_1030,N_632,N_782);
and U1031 (N_1031,N_714,N_856);
or U1032 (N_1032,In_630,N_650);
nor U1033 (N_1033,N_569,N_698);
nor U1034 (N_1034,N_878,In_332);
xnor U1035 (N_1035,N_830,In_520);
or U1036 (N_1036,N_647,In_186);
or U1037 (N_1037,In_1173,In_1471);
nor U1038 (N_1038,N_467,N_559);
or U1039 (N_1039,N_41,N_429);
nor U1040 (N_1040,N_771,N_540);
or U1041 (N_1041,N_690,N_834);
and U1042 (N_1042,In_288,N_54);
nor U1043 (N_1043,In_168,In_1297);
nand U1044 (N_1044,N_796,N_259);
nand U1045 (N_1045,N_591,N_860);
or U1046 (N_1046,N_762,N_706);
nand U1047 (N_1047,N_814,In_1477);
nand U1048 (N_1048,In_138,N_204);
and U1049 (N_1049,In_1075,N_748);
xor U1050 (N_1050,In_423,N_661);
nor U1051 (N_1051,N_709,N_881);
and U1052 (N_1052,N_622,In_139);
or U1053 (N_1053,In_945,In_187);
xor U1054 (N_1054,In_298,In_668);
or U1055 (N_1055,N_129,N_736);
or U1056 (N_1056,In_505,N_256);
nor U1057 (N_1057,N_694,In_303);
or U1058 (N_1058,In_1003,N_679);
xor U1059 (N_1059,N_758,N_3);
nor U1060 (N_1060,N_851,N_252);
or U1061 (N_1061,In_294,N_817);
and U1062 (N_1062,N_691,N_606);
and U1063 (N_1063,N_778,In_1424);
and U1064 (N_1064,N_859,N_202);
xor U1065 (N_1065,N_821,In_965);
and U1066 (N_1066,N_872,N_874);
nand U1067 (N_1067,N_315,N_865);
xor U1068 (N_1068,N_749,N_648);
nor U1069 (N_1069,N_707,N_13);
and U1070 (N_1070,N_450,In_100);
nor U1071 (N_1071,N_81,N_800);
and U1072 (N_1072,In_289,N_712);
or U1073 (N_1073,In_1113,N_122);
xnor U1074 (N_1074,N_378,N_787);
nand U1075 (N_1075,In_347,N_724);
xnor U1076 (N_1076,N_838,N_510);
nor U1077 (N_1077,N_671,In_1148);
nor U1078 (N_1078,N_826,In_615);
and U1079 (N_1079,N_891,In_850);
nor U1080 (N_1080,In_363,N_200);
or U1081 (N_1081,In_1252,N_411);
nor U1082 (N_1082,N_733,N_635);
or U1083 (N_1083,In_664,N_621);
nor U1084 (N_1084,N_892,N_170);
or U1085 (N_1085,N_600,In_182);
and U1086 (N_1086,In_560,N_828);
or U1087 (N_1087,N_446,N_696);
and U1088 (N_1088,In_526,In_451);
or U1089 (N_1089,N_788,N_636);
nor U1090 (N_1090,In_705,N_824);
nand U1091 (N_1091,N_734,In_102);
or U1092 (N_1092,N_682,N_883);
and U1093 (N_1093,N_658,N_448);
nor U1094 (N_1094,N_322,In_880);
xnor U1095 (N_1095,N_730,N_858);
xor U1096 (N_1096,N_793,In_963);
nand U1097 (N_1097,N_852,N_431);
xor U1098 (N_1098,N_693,N_550);
nor U1099 (N_1099,N_729,In_1179);
nand U1100 (N_1100,N_416,In_740);
xnor U1101 (N_1101,N_839,N_609);
and U1102 (N_1102,N_654,N_100);
nor U1103 (N_1103,N_853,N_732);
and U1104 (N_1104,N_695,In_1049);
nor U1105 (N_1105,N_754,In_869);
nand U1106 (N_1106,In_53,N_560);
xnor U1107 (N_1107,N_345,N_553);
or U1108 (N_1108,In_225,N_716);
and U1109 (N_1109,N_587,N_864);
and U1110 (N_1110,N_855,N_562);
nand U1111 (N_1111,In_726,In_1203);
and U1112 (N_1112,N_541,N_825);
or U1113 (N_1113,N_613,N_755);
or U1114 (N_1114,N_109,N_727);
nand U1115 (N_1115,In_1358,N_213);
or U1116 (N_1116,In_960,In_745);
xor U1117 (N_1117,N_704,N_808);
or U1118 (N_1118,In_612,N_794);
and U1119 (N_1119,N_139,N_408);
nor U1120 (N_1120,N_425,N_720);
nor U1121 (N_1121,In_1209,N_769);
and U1122 (N_1122,N_831,N_763);
xnor U1123 (N_1123,N_84,N_739);
xnor U1124 (N_1124,In_811,In_888);
and U1125 (N_1125,N_757,In_870);
and U1126 (N_1126,N_701,N_705);
or U1127 (N_1127,N_639,N_498);
and U1128 (N_1128,N_670,N_871);
xor U1129 (N_1129,N_667,In_491);
nor U1130 (N_1130,N_753,N_403);
nand U1131 (N_1131,N_770,N_463);
xor U1132 (N_1132,N_700,N_24);
nand U1133 (N_1133,N_689,N_85);
or U1134 (N_1134,N_868,In_1211);
nand U1135 (N_1135,N_399,N_73);
nand U1136 (N_1136,N_699,N_653);
xnor U1137 (N_1137,In_359,In_1134);
or U1138 (N_1138,N_816,N_49);
nand U1139 (N_1139,N_612,N_565);
or U1140 (N_1140,N_807,N_390);
nand U1141 (N_1141,N_889,N_809);
xor U1142 (N_1142,N_519,N_296);
or U1143 (N_1143,N_652,N_118);
or U1144 (N_1144,N_449,N_806);
and U1145 (N_1145,N_651,N_802);
and U1146 (N_1146,N_649,N_726);
or U1147 (N_1147,N_774,N_592);
nand U1148 (N_1148,N_879,N_662);
xnor U1149 (N_1149,N_646,N_728);
xor U1150 (N_1150,N_48,N_676);
and U1151 (N_1151,N_666,N_539);
and U1152 (N_1152,N_174,N_875);
nor U1153 (N_1153,N_876,N_342);
xnor U1154 (N_1154,N_761,N_657);
nand U1155 (N_1155,N_677,N_630);
nand U1156 (N_1156,N_721,N_348);
and U1157 (N_1157,N_766,N_895);
and U1158 (N_1158,N_890,N_887);
xnor U1159 (N_1159,N_372,N_641);
and U1160 (N_1160,N_668,N_187);
nand U1161 (N_1161,N_645,N_866);
or U1162 (N_1162,N_137,N_779);
or U1163 (N_1163,N_38,In_1299);
nor U1164 (N_1164,N_813,In_231);
nand U1165 (N_1165,N_683,N_482);
nor U1166 (N_1166,N_604,N_873);
nor U1167 (N_1167,In_600,In_1402);
or U1168 (N_1168,N_713,N_51);
or U1169 (N_1169,N_792,N_717);
nor U1170 (N_1170,N_746,N_161);
or U1171 (N_1171,N_464,N_366);
nand U1172 (N_1172,N_267,N_610);
and U1173 (N_1173,In_979,In_20);
nor U1174 (N_1174,In_297,N_281);
nand U1175 (N_1175,In_928,In_1485);
xnor U1176 (N_1176,N_53,N_804);
nor U1177 (N_1177,N_535,In_1066);
xor U1178 (N_1178,N_810,N_760);
nand U1179 (N_1179,In_897,N_162);
or U1180 (N_1180,In_261,N_737);
and U1181 (N_1181,N_517,N_327);
or U1182 (N_1182,In_157,N_669);
and U1183 (N_1183,N_659,In_1163);
and U1184 (N_1184,N_897,In_1071);
and U1185 (N_1185,N_278,N_725);
xnor U1186 (N_1186,N_465,In_1308);
and U1187 (N_1187,N_678,N_328);
and U1188 (N_1188,N_819,N_790);
or U1189 (N_1189,N_708,N_857);
nand U1190 (N_1190,N_805,In_1396);
xnor U1191 (N_1191,N_634,N_330);
nor U1192 (N_1192,N_703,N_886);
or U1193 (N_1193,N_601,N_50);
xnor U1194 (N_1194,N_381,N_836);
nor U1195 (N_1195,N_862,N_619);
or U1196 (N_1196,N_686,In_606);
and U1197 (N_1197,In_1461,N_815);
nor U1198 (N_1198,N_388,In_377);
xor U1199 (N_1199,N_767,N_439);
or U1200 (N_1200,N_1105,N_1004);
and U1201 (N_1201,N_1114,N_1092);
xnor U1202 (N_1202,N_947,N_1184);
and U1203 (N_1203,N_1175,N_1159);
xnor U1204 (N_1204,N_904,N_986);
nand U1205 (N_1205,N_968,N_1029);
nand U1206 (N_1206,N_1100,N_1053);
or U1207 (N_1207,N_932,N_1199);
nor U1208 (N_1208,N_1066,N_1194);
or U1209 (N_1209,N_956,N_980);
xor U1210 (N_1210,N_1189,N_1112);
nor U1211 (N_1211,N_1026,N_1145);
xnor U1212 (N_1212,N_1065,N_931);
or U1213 (N_1213,N_1115,N_1193);
nor U1214 (N_1214,N_1085,N_989);
and U1215 (N_1215,N_1182,N_1137);
and U1216 (N_1216,N_1014,N_1169);
xor U1217 (N_1217,N_1106,N_997);
or U1218 (N_1218,N_942,N_1118);
and U1219 (N_1219,N_1140,N_940);
or U1220 (N_1220,N_936,N_1099);
and U1221 (N_1221,N_984,N_955);
nand U1222 (N_1222,N_1186,N_1183);
nand U1223 (N_1223,N_954,N_1149);
or U1224 (N_1224,N_1061,N_1016);
and U1225 (N_1225,N_1018,N_951);
nand U1226 (N_1226,N_1077,N_1088);
and U1227 (N_1227,N_1000,N_1042);
xor U1228 (N_1228,N_925,N_1009);
nand U1229 (N_1229,N_982,N_1120);
nand U1230 (N_1230,N_1075,N_916);
or U1231 (N_1231,N_1177,N_1127);
nor U1232 (N_1232,N_923,N_1156);
nor U1233 (N_1233,N_1017,N_914);
and U1234 (N_1234,N_1068,N_1096);
or U1235 (N_1235,N_1025,N_1073);
and U1236 (N_1236,N_909,N_1166);
nand U1237 (N_1237,N_976,N_1072);
and U1238 (N_1238,N_929,N_1122);
and U1239 (N_1239,N_1171,N_958);
nand U1240 (N_1240,N_977,N_907);
or U1241 (N_1241,N_933,N_1113);
xnor U1242 (N_1242,N_1128,N_1070);
nand U1243 (N_1243,N_981,N_961);
nand U1244 (N_1244,N_922,N_1083);
or U1245 (N_1245,N_1136,N_1172);
and U1246 (N_1246,N_1086,N_1008);
or U1247 (N_1247,N_1154,N_1067);
xnor U1248 (N_1248,N_1142,N_1069);
xnor U1249 (N_1249,N_948,N_1050);
xnor U1250 (N_1250,N_1147,N_1150);
and U1251 (N_1251,N_1091,N_1165);
or U1252 (N_1252,N_1045,N_1121);
nor U1253 (N_1253,N_974,N_1058);
xnor U1254 (N_1254,N_1013,N_910);
xor U1255 (N_1255,N_1176,N_1101);
and U1256 (N_1256,N_971,N_1002);
nor U1257 (N_1257,N_999,N_1080);
nor U1258 (N_1258,N_1163,N_1117);
and U1259 (N_1259,N_930,N_1129);
xnor U1260 (N_1260,N_1144,N_902);
and U1261 (N_1261,N_1049,N_1041);
xor U1262 (N_1262,N_915,N_1152);
nor U1263 (N_1263,N_1051,N_917);
nand U1264 (N_1264,N_1012,N_1059);
or U1265 (N_1265,N_1043,N_965);
nor U1266 (N_1266,N_1030,N_957);
nor U1267 (N_1267,N_1191,N_995);
xnor U1268 (N_1268,N_1040,N_1039);
and U1269 (N_1269,N_1153,N_1035);
nand U1270 (N_1270,N_905,N_900);
xnor U1271 (N_1271,N_962,N_1021);
or U1272 (N_1272,N_1055,N_1010);
nand U1273 (N_1273,N_1123,N_1052);
xnor U1274 (N_1274,N_946,N_1146);
nor U1275 (N_1275,N_1098,N_913);
nand U1276 (N_1276,N_1031,N_1195);
or U1277 (N_1277,N_1160,N_1056);
xnor U1278 (N_1278,N_988,N_1158);
or U1279 (N_1279,N_960,N_1170);
xnor U1280 (N_1280,N_1047,N_998);
or U1281 (N_1281,N_983,N_1119);
nand U1282 (N_1282,N_1108,N_1187);
and U1283 (N_1283,N_1020,N_1179);
nand U1284 (N_1284,N_969,N_1139);
xnor U1285 (N_1285,N_964,N_941);
nor U1286 (N_1286,N_943,N_973);
nor U1287 (N_1287,N_1157,N_959);
or U1288 (N_1288,N_987,N_919);
and U1289 (N_1289,N_994,N_1033);
and U1290 (N_1290,N_1103,N_967);
xor U1291 (N_1291,N_921,N_991);
nand U1292 (N_1292,N_1078,N_990);
nand U1293 (N_1293,N_1110,N_1174);
and U1294 (N_1294,N_1022,N_949);
nand U1295 (N_1295,N_1102,N_1046);
xor U1296 (N_1296,N_937,N_1093);
nand U1297 (N_1297,N_945,N_1082);
xor U1298 (N_1298,N_1130,N_993);
xnor U1299 (N_1299,N_927,N_1131);
nand U1300 (N_1300,N_1135,N_1003);
xnor U1301 (N_1301,N_1109,N_1005);
and U1302 (N_1302,N_1062,N_1060);
nand U1303 (N_1303,N_950,N_918);
xnor U1304 (N_1304,N_903,N_944);
nor U1305 (N_1305,N_1196,N_1133);
xor U1306 (N_1306,N_935,N_1006);
or U1307 (N_1307,N_1197,N_1173);
and U1308 (N_1308,N_1027,N_1074);
nor U1309 (N_1309,N_1037,N_1063);
and U1310 (N_1310,N_1132,N_924);
nand U1311 (N_1311,N_963,N_1028);
nand U1312 (N_1312,N_1071,N_1104);
and U1313 (N_1313,N_1097,N_966);
or U1314 (N_1314,N_1034,N_1095);
nand U1315 (N_1315,N_912,N_1168);
nor U1316 (N_1316,N_1185,N_992);
nor U1317 (N_1317,N_908,N_1090);
xnor U1318 (N_1318,N_1036,N_1138);
xor U1319 (N_1319,N_1081,N_1054);
xor U1320 (N_1320,N_901,N_1032);
nand U1321 (N_1321,N_1190,N_1180);
nor U1322 (N_1322,N_1161,N_972);
or U1323 (N_1323,N_1188,N_1007);
and U1324 (N_1324,N_979,N_1084);
or U1325 (N_1325,N_911,N_1198);
or U1326 (N_1326,N_1124,N_953);
nand U1327 (N_1327,N_1148,N_1126);
nor U1328 (N_1328,N_1001,N_978);
and U1329 (N_1329,N_1038,N_1164);
and U1330 (N_1330,N_1019,N_928);
nand U1331 (N_1331,N_952,N_1076);
or U1332 (N_1332,N_938,N_1167);
and U1333 (N_1333,N_1162,N_1094);
and U1334 (N_1334,N_1155,N_1064);
or U1335 (N_1335,N_1089,N_1015);
nand U1336 (N_1336,N_1134,N_1141);
xor U1337 (N_1337,N_1181,N_1023);
xor U1338 (N_1338,N_1079,N_1143);
or U1339 (N_1339,N_1048,N_1024);
or U1340 (N_1340,N_934,N_1192);
nor U1341 (N_1341,N_1057,N_1111);
and U1342 (N_1342,N_1011,N_1178);
and U1343 (N_1343,N_1107,N_1044);
or U1344 (N_1344,N_906,N_939);
nor U1345 (N_1345,N_970,N_996);
and U1346 (N_1346,N_975,N_985);
and U1347 (N_1347,N_1151,N_1116);
nor U1348 (N_1348,N_920,N_1125);
or U1349 (N_1349,N_926,N_1087);
nor U1350 (N_1350,N_1158,N_1047);
xnor U1351 (N_1351,N_985,N_1085);
nor U1352 (N_1352,N_970,N_1146);
and U1353 (N_1353,N_1010,N_1125);
nand U1354 (N_1354,N_1183,N_1086);
or U1355 (N_1355,N_1074,N_1005);
or U1356 (N_1356,N_1028,N_1121);
nor U1357 (N_1357,N_1066,N_1062);
nand U1358 (N_1358,N_1075,N_1103);
or U1359 (N_1359,N_1052,N_1097);
xor U1360 (N_1360,N_1141,N_1155);
nor U1361 (N_1361,N_1038,N_1026);
or U1362 (N_1362,N_966,N_992);
or U1363 (N_1363,N_1037,N_995);
or U1364 (N_1364,N_1096,N_939);
or U1365 (N_1365,N_1126,N_1035);
nand U1366 (N_1366,N_900,N_999);
nand U1367 (N_1367,N_1146,N_915);
or U1368 (N_1368,N_922,N_1195);
and U1369 (N_1369,N_1163,N_1154);
nor U1370 (N_1370,N_1055,N_1045);
nor U1371 (N_1371,N_1180,N_1041);
or U1372 (N_1372,N_1111,N_1147);
nand U1373 (N_1373,N_1067,N_1151);
nor U1374 (N_1374,N_1072,N_1174);
or U1375 (N_1375,N_955,N_977);
xor U1376 (N_1376,N_1019,N_946);
xnor U1377 (N_1377,N_1192,N_1037);
and U1378 (N_1378,N_1197,N_1118);
xnor U1379 (N_1379,N_1080,N_1156);
nor U1380 (N_1380,N_1116,N_927);
and U1381 (N_1381,N_931,N_1024);
and U1382 (N_1382,N_1020,N_1195);
or U1383 (N_1383,N_1132,N_1058);
nand U1384 (N_1384,N_1091,N_1036);
and U1385 (N_1385,N_1098,N_1054);
and U1386 (N_1386,N_1166,N_1049);
and U1387 (N_1387,N_927,N_981);
xor U1388 (N_1388,N_1014,N_1086);
or U1389 (N_1389,N_1189,N_1197);
and U1390 (N_1390,N_1013,N_1125);
and U1391 (N_1391,N_1114,N_907);
nand U1392 (N_1392,N_1116,N_1167);
xor U1393 (N_1393,N_1061,N_1193);
or U1394 (N_1394,N_964,N_1028);
xnor U1395 (N_1395,N_1008,N_925);
nand U1396 (N_1396,N_1153,N_950);
nand U1397 (N_1397,N_1169,N_1037);
or U1398 (N_1398,N_1036,N_1025);
nand U1399 (N_1399,N_996,N_1084);
nand U1400 (N_1400,N_1139,N_1161);
xnor U1401 (N_1401,N_1196,N_1082);
and U1402 (N_1402,N_1065,N_1008);
xor U1403 (N_1403,N_1037,N_1035);
nand U1404 (N_1404,N_1090,N_991);
or U1405 (N_1405,N_937,N_1197);
nor U1406 (N_1406,N_1147,N_940);
or U1407 (N_1407,N_1149,N_1014);
and U1408 (N_1408,N_908,N_1089);
or U1409 (N_1409,N_996,N_1177);
nor U1410 (N_1410,N_917,N_1156);
and U1411 (N_1411,N_926,N_1116);
nor U1412 (N_1412,N_1002,N_1003);
and U1413 (N_1413,N_1104,N_906);
nor U1414 (N_1414,N_914,N_1029);
xnor U1415 (N_1415,N_952,N_1003);
or U1416 (N_1416,N_932,N_985);
xnor U1417 (N_1417,N_1007,N_1191);
xnor U1418 (N_1418,N_1188,N_1099);
nor U1419 (N_1419,N_997,N_1183);
and U1420 (N_1420,N_945,N_1079);
or U1421 (N_1421,N_923,N_1198);
and U1422 (N_1422,N_1194,N_912);
xor U1423 (N_1423,N_1140,N_1000);
or U1424 (N_1424,N_1115,N_1179);
nand U1425 (N_1425,N_924,N_902);
xnor U1426 (N_1426,N_1083,N_1161);
and U1427 (N_1427,N_1080,N_902);
and U1428 (N_1428,N_926,N_1012);
xor U1429 (N_1429,N_1198,N_964);
or U1430 (N_1430,N_1144,N_943);
and U1431 (N_1431,N_909,N_1127);
nand U1432 (N_1432,N_1155,N_1050);
and U1433 (N_1433,N_1192,N_1091);
nand U1434 (N_1434,N_1035,N_1199);
xor U1435 (N_1435,N_1198,N_993);
nor U1436 (N_1436,N_917,N_960);
nand U1437 (N_1437,N_1028,N_994);
xor U1438 (N_1438,N_1157,N_1145);
xnor U1439 (N_1439,N_986,N_1179);
or U1440 (N_1440,N_1136,N_1132);
and U1441 (N_1441,N_1018,N_1153);
and U1442 (N_1442,N_1185,N_943);
and U1443 (N_1443,N_1166,N_1021);
xor U1444 (N_1444,N_1066,N_1150);
xor U1445 (N_1445,N_909,N_1153);
and U1446 (N_1446,N_1186,N_1062);
or U1447 (N_1447,N_1105,N_1021);
xnor U1448 (N_1448,N_950,N_1124);
xnor U1449 (N_1449,N_1168,N_967);
or U1450 (N_1450,N_961,N_1053);
nand U1451 (N_1451,N_1148,N_1046);
and U1452 (N_1452,N_1053,N_1022);
nand U1453 (N_1453,N_1014,N_1194);
nor U1454 (N_1454,N_935,N_1055);
nand U1455 (N_1455,N_1115,N_1110);
nor U1456 (N_1456,N_936,N_1195);
or U1457 (N_1457,N_1166,N_1162);
nor U1458 (N_1458,N_900,N_1033);
and U1459 (N_1459,N_1037,N_1013);
xor U1460 (N_1460,N_1060,N_972);
xnor U1461 (N_1461,N_1091,N_945);
or U1462 (N_1462,N_911,N_1052);
xnor U1463 (N_1463,N_938,N_1102);
or U1464 (N_1464,N_957,N_1109);
nor U1465 (N_1465,N_935,N_1191);
xor U1466 (N_1466,N_916,N_1057);
or U1467 (N_1467,N_971,N_1051);
or U1468 (N_1468,N_1143,N_943);
xor U1469 (N_1469,N_1014,N_928);
or U1470 (N_1470,N_956,N_976);
nand U1471 (N_1471,N_918,N_1152);
and U1472 (N_1472,N_1174,N_1075);
nand U1473 (N_1473,N_1000,N_1032);
nor U1474 (N_1474,N_1127,N_1065);
xnor U1475 (N_1475,N_1150,N_1114);
and U1476 (N_1476,N_1024,N_1063);
xnor U1477 (N_1477,N_954,N_1182);
and U1478 (N_1478,N_1133,N_1189);
and U1479 (N_1479,N_952,N_1177);
and U1480 (N_1480,N_1184,N_1159);
nand U1481 (N_1481,N_1169,N_1125);
xor U1482 (N_1482,N_939,N_1005);
nor U1483 (N_1483,N_1010,N_1072);
or U1484 (N_1484,N_1150,N_981);
or U1485 (N_1485,N_1123,N_1015);
xor U1486 (N_1486,N_1181,N_975);
xnor U1487 (N_1487,N_1059,N_993);
nor U1488 (N_1488,N_1140,N_901);
nor U1489 (N_1489,N_1167,N_1096);
and U1490 (N_1490,N_962,N_978);
nand U1491 (N_1491,N_953,N_992);
or U1492 (N_1492,N_929,N_944);
nand U1493 (N_1493,N_1007,N_1012);
and U1494 (N_1494,N_1117,N_1006);
xor U1495 (N_1495,N_1148,N_1123);
and U1496 (N_1496,N_976,N_1050);
nor U1497 (N_1497,N_986,N_1154);
or U1498 (N_1498,N_924,N_1000);
nand U1499 (N_1499,N_1105,N_911);
nor U1500 (N_1500,N_1239,N_1287);
or U1501 (N_1501,N_1477,N_1434);
nor U1502 (N_1502,N_1328,N_1384);
nor U1503 (N_1503,N_1448,N_1277);
or U1504 (N_1504,N_1376,N_1294);
and U1505 (N_1505,N_1467,N_1402);
xnor U1506 (N_1506,N_1285,N_1338);
xor U1507 (N_1507,N_1469,N_1413);
nor U1508 (N_1508,N_1236,N_1224);
xor U1509 (N_1509,N_1279,N_1386);
nand U1510 (N_1510,N_1385,N_1461);
nand U1511 (N_1511,N_1257,N_1201);
and U1512 (N_1512,N_1489,N_1301);
or U1513 (N_1513,N_1395,N_1255);
nor U1514 (N_1514,N_1425,N_1443);
nor U1515 (N_1515,N_1412,N_1289);
or U1516 (N_1516,N_1280,N_1311);
nand U1517 (N_1517,N_1407,N_1358);
nor U1518 (N_1518,N_1292,N_1284);
nor U1519 (N_1519,N_1453,N_1482);
xnor U1520 (N_1520,N_1221,N_1403);
nor U1521 (N_1521,N_1213,N_1392);
nand U1522 (N_1522,N_1209,N_1488);
and U1523 (N_1523,N_1423,N_1444);
xnor U1524 (N_1524,N_1445,N_1336);
nand U1525 (N_1525,N_1238,N_1200);
xnor U1526 (N_1526,N_1315,N_1272);
and U1527 (N_1527,N_1281,N_1430);
nand U1528 (N_1528,N_1473,N_1278);
nor U1529 (N_1529,N_1442,N_1410);
and U1530 (N_1530,N_1370,N_1388);
and U1531 (N_1531,N_1214,N_1494);
xor U1532 (N_1532,N_1490,N_1433);
nor U1533 (N_1533,N_1310,N_1334);
and U1534 (N_1534,N_1458,N_1431);
nor U1535 (N_1535,N_1229,N_1233);
nor U1536 (N_1536,N_1265,N_1231);
xor U1537 (N_1537,N_1228,N_1266);
nor U1538 (N_1538,N_1223,N_1344);
or U1539 (N_1539,N_1339,N_1378);
or U1540 (N_1540,N_1372,N_1220);
xnor U1541 (N_1541,N_1424,N_1299);
nor U1542 (N_1542,N_1422,N_1426);
and U1543 (N_1543,N_1393,N_1457);
and U1544 (N_1544,N_1227,N_1212);
or U1545 (N_1545,N_1359,N_1319);
and U1546 (N_1546,N_1296,N_1234);
xor U1547 (N_1547,N_1364,N_1436);
xor U1548 (N_1548,N_1248,N_1268);
xor U1549 (N_1549,N_1346,N_1377);
xnor U1550 (N_1550,N_1345,N_1274);
or U1551 (N_1551,N_1361,N_1355);
and U1552 (N_1552,N_1454,N_1455);
nand U1553 (N_1553,N_1303,N_1493);
nor U1554 (N_1554,N_1232,N_1318);
xor U1555 (N_1555,N_1379,N_1235);
nand U1556 (N_1556,N_1230,N_1207);
nand U1557 (N_1557,N_1270,N_1219);
nand U1558 (N_1558,N_1373,N_1288);
and U1559 (N_1559,N_1365,N_1332);
nand U1560 (N_1560,N_1374,N_1481);
nand U1561 (N_1561,N_1251,N_1350);
nand U1562 (N_1562,N_1308,N_1399);
xnor U1563 (N_1563,N_1419,N_1499);
xnor U1564 (N_1564,N_1406,N_1456);
xnor U1565 (N_1565,N_1449,N_1471);
nand U1566 (N_1566,N_1450,N_1324);
and U1567 (N_1567,N_1447,N_1240);
or U1568 (N_1568,N_1258,N_1254);
or U1569 (N_1569,N_1371,N_1389);
nand U1570 (N_1570,N_1452,N_1275);
or U1571 (N_1571,N_1316,N_1269);
and U1572 (N_1572,N_1380,N_1253);
nand U1573 (N_1573,N_1416,N_1210);
nand U1574 (N_1574,N_1307,N_1331);
and U1575 (N_1575,N_1304,N_1252);
or U1576 (N_1576,N_1335,N_1362);
or U1577 (N_1577,N_1400,N_1263);
nor U1578 (N_1578,N_1330,N_1463);
and U1579 (N_1579,N_1347,N_1492);
nor U1580 (N_1580,N_1256,N_1405);
or U1581 (N_1581,N_1478,N_1348);
xor U1582 (N_1582,N_1421,N_1241);
or U1583 (N_1583,N_1203,N_1474);
nand U1584 (N_1584,N_1483,N_1353);
and U1585 (N_1585,N_1313,N_1205);
and U1586 (N_1586,N_1267,N_1367);
nor U1587 (N_1587,N_1320,N_1259);
and U1588 (N_1588,N_1298,N_1306);
or U1589 (N_1589,N_1498,N_1293);
and U1590 (N_1590,N_1390,N_1208);
xnor U1591 (N_1591,N_1475,N_1211);
and U1592 (N_1592,N_1391,N_1357);
nand U1593 (N_1593,N_1242,N_1437);
nand U1594 (N_1594,N_1446,N_1246);
or U1595 (N_1595,N_1343,N_1387);
nor U1596 (N_1596,N_1312,N_1354);
xor U1597 (N_1597,N_1322,N_1472);
xor U1598 (N_1598,N_1366,N_1314);
nor U1599 (N_1599,N_1369,N_1480);
nand U1600 (N_1600,N_1438,N_1414);
xnor U1601 (N_1601,N_1411,N_1394);
xor U1602 (N_1602,N_1262,N_1497);
nand U1603 (N_1603,N_1368,N_1300);
or U1604 (N_1604,N_1432,N_1290);
or U1605 (N_1605,N_1349,N_1427);
nor U1606 (N_1606,N_1382,N_1496);
nor U1607 (N_1607,N_1226,N_1476);
nor U1608 (N_1608,N_1282,N_1317);
xnor U1609 (N_1609,N_1360,N_1409);
or U1610 (N_1610,N_1225,N_1283);
nand U1611 (N_1611,N_1323,N_1460);
nor U1612 (N_1612,N_1273,N_1462);
nor U1613 (N_1613,N_1398,N_1222);
nor U1614 (N_1614,N_1217,N_1218);
xnor U1615 (N_1615,N_1479,N_1295);
xnor U1616 (N_1616,N_1491,N_1352);
and U1617 (N_1617,N_1381,N_1250);
or U1618 (N_1618,N_1291,N_1286);
nand U1619 (N_1619,N_1341,N_1487);
nor U1620 (N_1620,N_1356,N_1249);
and U1621 (N_1621,N_1351,N_1340);
and U1622 (N_1622,N_1302,N_1428);
or U1623 (N_1623,N_1363,N_1401);
or U1624 (N_1624,N_1260,N_1321);
nor U1625 (N_1625,N_1261,N_1325);
or U1626 (N_1626,N_1439,N_1297);
nand U1627 (N_1627,N_1429,N_1216);
and U1628 (N_1628,N_1276,N_1329);
and U1629 (N_1629,N_1206,N_1202);
xor U1630 (N_1630,N_1408,N_1237);
or U1631 (N_1631,N_1466,N_1465);
nor U1632 (N_1632,N_1396,N_1495);
nand U1633 (N_1633,N_1271,N_1459);
nor U1634 (N_1634,N_1342,N_1245);
and U1635 (N_1635,N_1418,N_1337);
nor U1636 (N_1636,N_1420,N_1435);
nor U1637 (N_1637,N_1486,N_1441);
nand U1638 (N_1638,N_1247,N_1451);
nor U1639 (N_1639,N_1204,N_1468);
xor U1640 (N_1640,N_1417,N_1404);
xnor U1641 (N_1641,N_1470,N_1243);
and U1642 (N_1642,N_1215,N_1464);
and U1643 (N_1643,N_1415,N_1397);
and U1644 (N_1644,N_1485,N_1244);
and U1645 (N_1645,N_1264,N_1327);
nand U1646 (N_1646,N_1333,N_1484);
nor U1647 (N_1647,N_1305,N_1309);
xor U1648 (N_1648,N_1383,N_1375);
or U1649 (N_1649,N_1440,N_1326);
nand U1650 (N_1650,N_1283,N_1434);
nor U1651 (N_1651,N_1270,N_1403);
or U1652 (N_1652,N_1435,N_1348);
or U1653 (N_1653,N_1282,N_1289);
nand U1654 (N_1654,N_1357,N_1392);
or U1655 (N_1655,N_1323,N_1445);
nand U1656 (N_1656,N_1363,N_1327);
nand U1657 (N_1657,N_1473,N_1474);
xor U1658 (N_1658,N_1364,N_1343);
nand U1659 (N_1659,N_1211,N_1253);
and U1660 (N_1660,N_1235,N_1484);
nand U1661 (N_1661,N_1435,N_1417);
nand U1662 (N_1662,N_1444,N_1275);
or U1663 (N_1663,N_1223,N_1222);
and U1664 (N_1664,N_1433,N_1275);
xnor U1665 (N_1665,N_1474,N_1208);
xnor U1666 (N_1666,N_1421,N_1488);
and U1667 (N_1667,N_1251,N_1442);
nand U1668 (N_1668,N_1498,N_1447);
or U1669 (N_1669,N_1339,N_1428);
and U1670 (N_1670,N_1492,N_1331);
xor U1671 (N_1671,N_1250,N_1448);
xor U1672 (N_1672,N_1416,N_1375);
and U1673 (N_1673,N_1347,N_1456);
xnor U1674 (N_1674,N_1377,N_1351);
xnor U1675 (N_1675,N_1399,N_1423);
nand U1676 (N_1676,N_1350,N_1312);
or U1677 (N_1677,N_1230,N_1210);
nand U1678 (N_1678,N_1347,N_1255);
nor U1679 (N_1679,N_1281,N_1210);
and U1680 (N_1680,N_1301,N_1317);
nand U1681 (N_1681,N_1327,N_1308);
and U1682 (N_1682,N_1312,N_1453);
and U1683 (N_1683,N_1498,N_1390);
xor U1684 (N_1684,N_1205,N_1432);
xor U1685 (N_1685,N_1483,N_1485);
nor U1686 (N_1686,N_1202,N_1335);
or U1687 (N_1687,N_1253,N_1422);
nor U1688 (N_1688,N_1336,N_1332);
xor U1689 (N_1689,N_1454,N_1270);
or U1690 (N_1690,N_1234,N_1345);
or U1691 (N_1691,N_1349,N_1246);
nor U1692 (N_1692,N_1403,N_1303);
or U1693 (N_1693,N_1201,N_1401);
xor U1694 (N_1694,N_1448,N_1441);
and U1695 (N_1695,N_1465,N_1346);
and U1696 (N_1696,N_1392,N_1367);
nor U1697 (N_1697,N_1459,N_1360);
and U1698 (N_1698,N_1264,N_1257);
nor U1699 (N_1699,N_1483,N_1410);
xor U1700 (N_1700,N_1257,N_1463);
nand U1701 (N_1701,N_1391,N_1306);
nand U1702 (N_1702,N_1371,N_1257);
and U1703 (N_1703,N_1336,N_1219);
and U1704 (N_1704,N_1460,N_1499);
and U1705 (N_1705,N_1276,N_1442);
xor U1706 (N_1706,N_1499,N_1334);
nand U1707 (N_1707,N_1291,N_1393);
xnor U1708 (N_1708,N_1332,N_1316);
xnor U1709 (N_1709,N_1489,N_1274);
and U1710 (N_1710,N_1457,N_1422);
and U1711 (N_1711,N_1206,N_1295);
or U1712 (N_1712,N_1294,N_1330);
nor U1713 (N_1713,N_1226,N_1376);
xnor U1714 (N_1714,N_1480,N_1259);
xor U1715 (N_1715,N_1304,N_1413);
nor U1716 (N_1716,N_1463,N_1250);
or U1717 (N_1717,N_1393,N_1469);
or U1718 (N_1718,N_1339,N_1442);
and U1719 (N_1719,N_1393,N_1320);
or U1720 (N_1720,N_1234,N_1287);
nor U1721 (N_1721,N_1303,N_1200);
nor U1722 (N_1722,N_1434,N_1255);
xnor U1723 (N_1723,N_1224,N_1210);
and U1724 (N_1724,N_1215,N_1445);
nand U1725 (N_1725,N_1454,N_1252);
nand U1726 (N_1726,N_1348,N_1215);
or U1727 (N_1727,N_1424,N_1202);
nor U1728 (N_1728,N_1385,N_1257);
xor U1729 (N_1729,N_1465,N_1449);
xor U1730 (N_1730,N_1267,N_1376);
nor U1731 (N_1731,N_1308,N_1407);
nand U1732 (N_1732,N_1225,N_1411);
nand U1733 (N_1733,N_1277,N_1411);
xnor U1734 (N_1734,N_1277,N_1325);
and U1735 (N_1735,N_1452,N_1289);
nand U1736 (N_1736,N_1223,N_1259);
or U1737 (N_1737,N_1232,N_1498);
or U1738 (N_1738,N_1218,N_1239);
nand U1739 (N_1739,N_1377,N_1256);
and U1740 (N_1740,N_1213,N_1316);
xor U1741 (N_1741,N_1287,N_1473);
nand U1742 (N_1742,N_1469,N_1429);
nor U1743 (N_1743,N_1458,N_1280);
nor U1744 (N_1744,N_1393,N_1383);
or U1745 (N_1745,N_1336,N_1448);
nor U1746 (N_1746,N_1393,N_1390);
xor U1747 (N_1747,N_1437,N_1260);
or U1748 (N_1748,N_1323,N_1209);
and U1749 (N_1749,N_1353,N_1497);
nand U1750 (N_1750,N_1208,N_1439);
xnor U1751 (N_1751,N_1247,N_1419);
nor U1752 (N_1752,N_1492,N_1297);
or U1753 (N_1753,N_1276,N_1447);
xor U1754 (N_1754,N_1241,N_1411);
nor U1755 (N_1755,N_1204,N_1447);
nor U1756 (N_1756,N_1386,N_1472);
nor U1757 (N_1757,N_1207,N_1297);
nor U1758 (N_1758,N_1436,N_1387);
nand U1759 (N_1759,N_1462,N_1439);
nand U1760 (N_1760,N_1399,N_1236);
and U1761 (N_1761,N_1236,N_1325);
and U1762 (N_1762,N_1290,N_1465);
nand U1763 (N_1763,N_1243,N_1314);
nor U1764 (N_1764,N_1440,N_1201);
xnor U1765 (N_1765,N_1408,N_1205);
nor U1766 (N_1766,N_1375,N_1349);
xnor U1767 (N_1767,N_1271,N_1219);
or U1768 (N_1768,N_1276,N_1467);
nand U1769 (N_1769,N_1446,N_1448);
xor U1770 (N_1770,N_1257,N_1482);
nor U1771 (N_1771,N_1287,N_1483);
nor U1772 (N_1772,N_1461,N_1293);
xor U1773 (N_1773,N_1363,N_1294);
nor U1774 (N_1774,N_1398,N_1271);
and U1775 (N_1775,N_1363,N_1292);
or U1776 (N_1776,N_1376,N_1305);
nand U1777 (N_1777,N_1406,N_1209);
nor U1778 (N_1778,N_1288,N_1230);
xor U1779 (N_1779,N_1209,N_1208);
xnor U1780 (N_1780,N_1346,N_1278);
and U1781 (N_1781,N_1331,N_1282);
or U1782 (N_1782,N_1322,N_1435);
or U1783 (N_1783,N_1433,N_1345);
xnor U1784 (N_1784,N_1378,N_1413);
nor U1785 (N_1785,N_1316,N_1266);
nand U1786 (N_1786,N_1331,N_1323);
xor U1787 (N_1787,N_1420,N_1300);
nand U1788 (N_1788,N_1214,N_1222);
or U1789 (N_1789,N_1215,N_1259);
or U1790 (N_1790,N_1477,N_1312);
nor U1791 (N_1791,N_1341,N_1486);
or U1792 (N_1792,N_1288,N_1474);
or U1793 (N_1793,N_1245,N_1460);
nor U1794 (N_1794,N_1476,N_1373);
nand U1795 (N_1795,N_1233,N_1270);
xnor U1796 (N_1796,N_1276,N_1389);
xnor U1797 (N_1797,N_1412,N_1465);
and U1798 (N_1798,N_1423,N_1359);
nand U1799 (N_1799,N_1347,N_1237);
nor U1800 (N_1800,N_1768,N_1590);
nor U1801 (N_1801,N_1558,N_1535);
nor U1802 (N_1802,N_1625,N_1614);
xor U1803 (N_1803,N_1512,N_1545);
xnor U1804 (N_1804,N_1751,N_1774);
or U1805 (N_1805,N_1728,N_1583);
and U1806 (N_1806,N_1563,N_1561);
and U1807 (N_1807,N_1607,N_1679);
or U1808 (N_1808,N_1662,N_1784);
nand U1809 (N_1809,N_1640,N_1668);
or U1810 (N_1810,N_1566,N_1788);
and U1811 (N_1811,N_1783,N_1584);
or U1812 (N_1812,N_1622,N_1579);
and U1813 (N_1813,N_1691,N_1792);
or U1814 (N_1814,N_1671,N_1652);
nor U1815 (N_1815,N_1616,N_1582);
nor U1816 (N_1816,N_1639,N_1743);
and U1817 (N_1817,N_1505,N_1696);
xor U1818 (N_1818,N_1504,N_1771);
and U1819 (N_1819,N_1531,N_1528);
xnor U1820 (N_1820,N_1565,N_1739);
nor U1821 (N_1821,N_1549,N_1663);
and U1822 (N_1822,N_1723,N_1572);
nor U1823 (N_1823,N_1740,N_1519);
xor U1824 (N_1824,N_1627,N_1514);
xor U1825 (N_1825,N_1536,N_1611);
or U1826 (N_1826,N_1715,N_1653);
xnor U1827 (N_1827,N_1559,N_1560);
nand U1828 (N_1828,N_1593,N_1576);
and U1829 (N_1829,N_1626,N_1721);
or U1830 (N_1830,N_1642,N_1608);
xnor U1831 (N_1831,N_1730,N_1704);
and U1832 (N_1832,N_1580,N_1508);
nand U1833 (N_1833,N_1754,N_1797);
or U1834 (N_1834,N_1568,N_1647);
and U1835 (N_1835,N_1676,N_1592);
xor U1836 (N_1836,N_1588,N_1620);
nand U1837 (N_1837,N_1746,N_1524);
and U1838 (N_1838,N_1760,N_1513);
xnor U1839 (N_1839,N_1795,N_1769);
nand U1840 (N_1840,N_1711,N_1610);
xnor U1841 (N_1841,N_1683,N_1602);
or U1842 (N_1842,N_1507,N_1726);
xor U1843 (N_1843,N_1598,N_1701);
and U1844 (N_1844,N_1537,N_1681);
nor U1845 (N_1845,N_1776,N_1775);
nor U1846 (N_1846,N_1687,N_1707);
or U1847 (N_1847,N_1510,N_1578);
nor U1848 (N_1848,N_1621,N_1694);
xnor U1849 (N_1849,N_1667,N_1759);
xnor U1850 (N_1850,N_1778,N_1752);
or U1851 (N_1851,N_1717,N_1773);
and U1852 (N_1852,N_1757,N_1596);
or U1853 (N_1853,N_1678,N_1737);
nand U1854 (N_1854,N_1664,N_1722);
nor U1855 (N_1855,N_1539,N_1591);
or U1856 (N_1856,N_1511,N_1503);
or U1857 (N_1857,N_1782,N_1571);
nand U1858 (N_1858,N_1673,N_1601);
and U1859 (N_1859,N_1628,N_1762);
and U1860 (N_1860,N_1523,N_1763);
xor U1861 (N_1861,N_1789,N_1686);
nand U1862 (N_1862,N_1644,N_1706);
or U1863 (N_1863,N_1660,N_1731);
and U1864 (N_1864,N_1574,N_1506);
nand U1865 (N_1865,N_1680,N_1518);
or U1866 (N_1866,N_1509,N_1594);
or U1867 (N_1867,N_1700,N_1542);
and U1868 (N_1868,N_1765,N_1713);
xor U1869 (N_1869,N_1597,N_1648);
nor U1870 (N_1870,N_1793,N_1770);
nand U1871 (N_1871,N_1637,N_1570);
or U1872 (N_1872,N_1530,N_1650);
nand U1873 (N_1873,N_1780,N_1645);
and U1874 (N_1874,N_1636,N_1745);
nand U1875 (N_1875,N_1712,N_1781);
nand U1876 (N_1876,N_1716,N_1585);
or U1877 (N_1877,N_1693,N_1688);
nand U1878 (N_1878,N_1672,N_1556);
nand U1879 (N_1879,N_1538,N_1532);
or U1880 (N_1880,N_1738,N_1761);
nor U1881 (N_1881,N_1790,N_1682);
nor U1882 (N_1882,N_1695,N_1791);
nand U1883 (N_1883,N_1655,N_1777);
xnor U1884 (N_1884,N_1517,N_1697);
nand U1885 (N_1885,N_1744,N_1750);
or U1886 (N_1886,N_1675,N_1665);
and U1887 (N_1887,N_1548,N_1742);
or U1888 (N_1888,N_1562,N_1515);
xor U1889 (N_1889,N_1658,N_1699);
or U1890 (N_1890,N_1609,N_1547);
nand U1891 (N_1891,N_1719,N_1550);
and U1892 (N_1892,N_1500,N_1729);
and U1893 (N_1893,N_1689,N_1604);
and U1894 (N_1894,N_1555,N_1674);
nor U1895 (N_1895,N_1600,N_1618);
and U1896 (N_1896,N_1564,N_1657);
or U1897 (N_1897,N_1787,N_1613);
nor U1898 (N_1898,N_1772,N_1629);
and U1899 (N_1899,N_1641,N_1724);
or U1900 (N_1900,N_1573,N_1702);
and U1901 (N_1901,N_1794,N_1685);
xor U1902 (N_1902,N_1632,N_1534);
nor U1903 (N_1903,N_1525,N_1799);
or U1904 (N_1904,N_1755,N_1516);
nand U1905 (N_1905,N_1612,N_1522);
xor U1906 (N_1906,N_1698,N_1581);
or U1907 (N_1907,N_1748,N_1520);
or U1908 (N_1908,N_1714,N_1661);
nand U1909 (N_1909,N_1638,N_1786);
and U1910 (N_1910,N_1623,N_1521);
and U1911 (N_1911,N_1646,N_1654);
nand U1912 (N_1912,N_1669,N_1708);
and U1913 (N_1913,N_1684,N_1586);
nand U1914 (N_1914,N_1798,N_1753);
or U1915 (N_1915,N_1554,N_1533);
nor U1916 (N_1916,N_1734,N_1589);
and U1917 (N_1917,N_1587,N_1633);
xnor U1918 (N_1918,N_1599,N_1756);
nor U1919 (N_1919,N_1732,N_1736);
nor U1920 (N_1920,N_1552,N_1785);
and U1921 (N_1921,N_1649,N_1767);
or U1922 (N_1922,N_1619,N_1779);
or U1923 (N_1923,N_1569,N_1656);
nor U1924 (N_1924,N_1617,N_1544);
xnor U1925 (N_1925,N_1710,N_1630);
nor U1926 (N_1926,N_1615,N_1635);
nand U1927 (N_1927,N_1557,N_1709);
xnor U1928 (N_1928,N_1718,N_1546);
nor U1929 (N_1929,N_1595,N_1540);
and U1930 (N_1930,N_1670,N_1727);
nor U1931 (N_1931,N_1766,N_1733);
xnor U1932 (N_1932,N_1567,N_1501);
or U1933 (N_1933,N_1741,N_1677);
nand U1934 (N_1934,N_1551,N_1575);
or U1935 (N_1935,N_1758,N_1631);
nand U1936 (N_1936,N_1541,N_1692);
nand U1937 (N_1937,N_1543,N_1526);
xnor U1938 (N_1938,N_1703,N_1634);
nor U1939 (N_1939,N_1747,N_1603);
nand U1940 (N_1940,N_1764,N_1666);
nor U1941 (N_1941,N_1651,N_1553);
or U1942 (N_1942,N_1720,N_1527);
and U1943 (N_1943,N_1624,N_1606);
or U1944 (N_1944,N_1577,N_1529);
or U1945 (N_1945,N_1690,N_1643);
or U1946 (N_1946,N_1796,N_1605);
or U1947 (N_1947,N_1502,N_1705);
and U1948 (N_1948,N_1659,N_1749);
nor U1949 (N_1949,N_1735,N_1725);
or U1950 (N_1950,N_1706,N_1509);
nand U1951 (N_1951,N_1722,N_1587);
nand U1952 (N_1952,N_1584,N_1755);
or U1953 (N_1953,N_1573,N_1565);
xnor U1954 (N_1954,N_1560,N_1644);
nor U1955 (N_1955,N_1742,N_1505);
nand U1956 (N_1956,N_1523,N_1760);
xnor U1957 (N_1957,N_1570,N_1769);
and U1958 (N_1958,N_1536,N_1604);
nand U1959 (N_1959,N_1660,N_1629);
xnor U1960 (N_1960,N_1694,N_1709);
and U1961 (N_1961,N_1688,N_1638);
nand U1962 (N_1962,N_1783,N_1709);
xor U1963 (N_1963,N_1721,N_1504);
nand U1964 (N_1964,N_1633,N_1683);
nand U1965 (N_1965,N_1532,N_1793);
and U1966 (N_1966,N_1583,N_1589);
nand U1967 (N_1967,N_1626,N_1517);
nor U1968 (N_1968,N_1706,N_1769);
xor U1969 (N_1969,N_1544,N_1761);
or U1970 (N_1970,N_1775,N_1579);
and U1971 (N_1971,N_1645,N_1671);
or U1972 (N_1972,N_1591,N_1586);
nor U1973 (N_1973,N_1710,N_1793);
and U1974 (N_1974,N_1771,N_1681);
nand U1975 (N_1975,N_1679,N_1601);
and U1976 (N_1976,N_1690,N_1769);
nor U1977 (N_1977,N_1570,N_1614);
xnor U1978 (N_1978,N_1687,N_1771);
or U1979 (N_1979,N_1756,N_1798);
nor U1980 (N_1980,N_1631,N_1533);
or U1981 (N_1981,N_1638,N_1628);
xnor U1982 (N_1982,N_1504,N_1697);
xnor U1983 (N_1983,N_1788,N_1681);
and U1984 (N_1984,N_1726,N_1647);
and U1985 (N_1985,N_1707,N_1695);
nor U1986 (N_1986,N_1617,N_1586);
nor U1987 (N_1987,N_1730,N_1794);
nor U1988 (N_1988,N_1690,N_1758);
nand U1989 (N_1989,N_1607,N_1587);
nand U1990 (N_1990,N_1792,N_1502);
xnor U1991 (N_1991,N_1749,N_1796);
nand U1992 (N_1992,N_1556,N_1655);
or U1993 (N_1993,N_1618,N_1522);
nand U1994 (N_1994,N_1646,N_1603);
nand U1995 (N_1995,N_1709,N_1639);
xor U1996 (N_1996,N_1690,N_1749);
nand U1997 (N_1997,N_1538,N_1706);
nand U1998 (N_1998,N_1635,N_1781);
or U1999 (N_1999,N_1665,N_1500);
or U2000 (N_2000,N_1621,N_1606);
xor U2001 (N_2001,N_1762,N_1699);
nand U2002 (N_2002,N_1794,N_1533);
nand U2003 (N_2003,N_1700,N_1515);
xnor U2004 (N_2004,N_1722,N_1525);
and U2005 (N_2005,N_1794,N_1787);
nand U2006 (N_2006,N_1727,N_1712);
xnor U2007 (N_2007,N_1619,N_1615);
and U2008 (N_2008,N_1726,N_1644);
and U2009 (N_2009,N_1648,N_1609);
nand U2010 (N_2010,N_1571,N_1518);
or U2011 (N_2011,N_1649,N_1597);
or U2012 (N_2012,N_1692,N_1735);
xor U2013 (N_2013,N_1734,N_1713);
nor U2014 (N_2014,N_1681,N_1526);
and U2015 (N_2015,N_1539,N_1789);
nor U2016 (N_2016,N_1727,N_1545);
and U2017 (N_2017,N_1525,N_1765);
nor U2018 (N_2018,N_1507,N_1637);
or U2019 (N_2019,N_1737,N_1696);
and U2020 (N_2020,N_1633,N_1626);
and U2021 (N_2021,N_1555,N_1788);
and U2022 (N_2022,N_1774,N_1604);
and U2023 (N_2023,N_1790,N_1572);
nor U2024 (N_2024,N_1676,N_1784);
and U2025 (N_2025,N_1756,N_1762);
nand U2026 (N_2026,N_1519,N_1765);
xor U2027 (N_2027,N_1581,N_1593);
nand U2028 (N_2028,N_1705,N_1712);
or U2029 (N_2029,N_1746,N_1749);
nor U2030 (N_2030,N_1744,N_1608);
nor U2031 (N_2031,N_1788,N_1725);
xnor U2032 (N_2032,N_1686,N_1584);
or U2033 (N_2033,N_1696,N_1604);
nand U2034 (N_2034,N_1538,N_1679);
xnor U2035 (N_2035,N_1761,N_1655);
nand U2036 (N_2036,N_1510,N_1769);
xnor U2037 (N_2037,N_1680,N_1780);
and U2038 (N_2038,N_1608,N_1792);
xnor U2039 (N_2039,N_1532,N_1614);
xnor U2040 (N_2040,N_1733,N_1520);
xor U2041 (N_2041,N_1645,N_1578);
xor U2042 (N_2042,N_1509,N_1739);
nor U2043 (N_2043,N_1793,N_1641);
nor U2044 (N_2044,N_1642,N_1510);
or U2045 (N_2045,N_1743,N_1580);
or U2046 (N_2046,N_1638,N_1778);
or U2047 (N_2047,N_1732,N_1712);
xor U2048 (N_2048,N_1769,N_1506);
xnor U2049 (N_2049,N_1647,N_1784);
nand U2050 (N_2050,N_1545,N_1687);
nor U2051 (N_2051,N_1617,N_1721);
or U2052 (N_2052,N_1564,N_1663);
xnor U2053 (N_2053,N_1713,N_1692);
and U2054 (N_2054,N_1630,N_1755);
nand U2055 (N_2055,N_1519,N_1782);
xor U2056 (N_2056,N_1668,N_1641);
xnor U2057 (N_2057,N_1651,N_1708);
xor U2058 (N_2058,N_1654,N_1572);
and U2059 (N_2059,N_1783,N_1683);
and U2060 (N_2060,N_1624,N_1500);
and U2061 (N_2061,N_1505,N_1509);
xor U2062 (N_2062,N_1658,N_1534);
and U2063 (N_2063,N_1632,N_1790);
or U2064 (N_2064,N_1651,N_1539);
nor U2065 (N_2065,N_1540,N_1754);
nand U2066 (N_2066,N_1701,N_1690);
nand U2067 (N_2067,N_1752,N_1618);
and U2068 (N_2068,N_1659,N_1761);
and U2069 (N_2069,N_1762,N_1748);
and U2070 (N_2070,N_1609,N_1720);
nand U2071 (N_2071,N_1668,N_1655);
nand U2072 (N_2072,N_1622,N_1751);
xor U2073 (N_2073,N_1583,N_1601);
xnor U2074 (N_2074,N_1757,N_1681);
nor U2075 (N_2075,N_1676,N_1563);
nand U2076 (N_2076,N_1759,N_1601);
nand U2077 (N_2077,N_1755,N_1716);
nand U2078 (N_2078,N_1559,N_1672);
or U2079 (N_2079,N_1526,N_1636);
xnor U2080 (N_2080,N_1502,N_1682);
nand U2081 (N_2081,N_1565,N_1662);
and U2082 (N_2082,N_1663,N_1576);
or U2083 (N_2083,N_1675,N_1733);
nor U2084 (N_2084,N_1608,N_1633);
or U2085 (N_2085,N_1542,N_1590);
nor U2086 (N_2086,N_1549,N_1585);
xor U2087 (N_2087,N_1694,N_1533);
xnor U2088 (N_2088,N_1529,N_1563);
nand U2089 (N_2089,N_1506,N_1731);
and U2090 (N_2090,N_1759,N_1746);
nor U2091 (N_2091,N_1629,N_1756);
nor U2092 (N_2092,N_1634,N_1669);
and U2093 (N_2093,N_1584,N_1600);
or U2094 (N_2094,N_1538,N_1591);
or U2095 (N_2095,N_1679,N_1517);
nand U2096 (N_2096,N_1789,N_1558);
nand U2097 (N_2097,N_1639,N_1661);
and U2098 (N_2098,N_1735,N_1637);
xnor U2099 (N_2099,N_1728,N_1727);
nand U2100 (N_2100,N_2007,N_2055);
and U2101 (N_2101,N_2043,N_1928);
nor U2102 (N_2102,N_2077,N_1889);
nor U2103 (N_2103,N_1999,N_1997);
or U2104 (N_2104,N_2065,N_1850);
and U2105 (N_2105,N_1977,N_1884);
nand U2106 (N_2106,N_1992,N_1892);
nor U2107 (N_2107,N_1930,N_1949);
or U2108 (N_2108,N_2023,N_1905);
and U2109 (N_2109,N_2045,N_2068);
nor U2110 (N_2110,N_1953,N_1980);
nor U2111 (N_2111,N_2099,N_2024);
or U2112 (N_2112,N_2053,N_2057);
nor U2113 (N_2113,N_1899,N_1860);
or U2114 (N_2114,N_2091,N_1918);
xnor U2115 (N_2115,N_1983,N_2036);
xor U2116 (N_2116,N_2079,N_1841);
xnor U2117 (N_2117,N_1950,N_1811);
or U2118 (N_2118,N_1969,N_1966);
or U2119 (N_2119,N_2031,N_1991);
nor U2120 (N_2120,N_1874,N_2019);
nor U2121 (N_2121,N_1978,N_1971);
or U2122 (N_2122,N_1847,N_1832);
or U2123 (N_2123,N_1931,N_2022);
and U2124 (N_2124,N_1806,N_1948);
nand U2125 (N_2125,N_2064,N_1984);
or U2126 (N_2126,N_2012,N_2062);
nand U2127 (N_2127,N_1946,N_2011);
and U2128 (N_2128,N_1943,N_2032);
and U2129 (N_2129,N_1820,N_1848);
or U2130 (N_2130,N_1907,N_2049);
xor U2131 (N_2131,N_2074,N_1976);
xnor U2132 (N_2132,N_1834,N_1888);
and U2133 (N_2133,N_1803,N_2084);
and U2134 (N_2134,N_2014,N_1814);
and U2135 (N_2135,N_1817,N_2020);
nand U2136 (N_2136,N_1898,N_2004);
and U2137 (N_2137,N_1939,N_1895);
or U2138 (N_2138,N_1944,N_2013);
and U2139 (N_2139,N_2039,N_1998);
nand U2140 (N_2140,N_1843,N_1925);
and U2141 (N_2141,N_1807,N_1990);
and U2142 (N_2142,N_1979,N_1871);
nor U2143 (N_2143,N_2001,N_1824);
nor U2144 (N_2144,N_1861,N_2086);
xor U2145 (N_2145,N_1970,N_1858);
nand U2146 (N_2146,N_1896,N_1813);
nor U2147 (N_2147,N_1972,N_1805);
nor U2148 (N_2148,N_2090,N_2080);
or U2149 (N_2149,N_1937,N_1800);
xnor U2150 (N_2150,N_2008,N_1870);
and U2151 (N_2151,N_2052,N_2009);
or U2152 (N_2152,N_1849,N_1873);
or U2153 (N_2153,N_2069,N_1965);
and U2154 (N_2154,N_1818,N_1879);
nand U2155 (N_2155,N_2070,N_2034);
nor U2156 (N_2156,N_1826,N_2076);
nand U2157 (N_2157,N_2054,N_1844);
and U2158 (N_2158,N_1919,N_1900);
or U2159 (N_2159,N_1866,N_2056);
xor U2160 (N_2160,N_1869,N_1904);
nor U2161 (N_2161,N_1938,N_1880);
and U2162 (N_2162,N_1961,N_1862);
nor U2163 (N_2163,N_1868,N_1819);
or U2164 (N_2164,N_1917,N_2025);
nor U2165 (N_2165,N_1893,N_2037);
xnor U2166 (N_2166,N_1973,N_1887);
xor U2167 (N_2167,N_1876,N_2047);
or U2168 (N_2168,N_2096,N_1962);
nand U2169 (N_2169,N_1902,N_1875);
xor U2170 (N_2170,N_1901,N_1822);
or U2171 (N_2171,N_1897,N_2067);
xor U2172 (N_2172,N_1957,N_2038);
nand U2173 (N_2173,N_1838,N_1994);
and U2174 (N_2174,N_1837,N_2033);
nor U2175 (N_2175,N_1906,N_1996);
nor U2176 (N_2176,N_1955,N_1926);
nand U2177 (N_2177,N_1924,N_1885);
xnor U2178 (N_2178,N_1864,N_1975);
nand U2179 (N_2179,N_2015,N_1867);
or U2180 (N_2180,N_1883,N_2066);
nor U2181 (N_2181,N_1828,N_1914);
nor U2182 (N_2182,N_1865,N_1951);
and U2183 (N_2183,N_1856,N_1809);
nor U2184 (N_2184,N_1960,N_1916);
nor U2185 (N_2185,N_1827,N_1836);
xnor U2186 (N_2186,N_1815,N_1933);
nand U2187 (N_2187,N_2095,N_2073);
or U2188 (N_2188,N_2029,N_2085);
xor U2189 (N_2189,N_1855,N_2048);
or U2190 (N_2190,N_1821,N_1987);
or U2191 (N_2191,N_1968,N_1816);
nor U2192 (N_2192,N_1956,N_1891);
nand U2193 (N_2193,N_1825,N_1830);
nand U2194 (N_2194,N_1921,N_2046);
xnor U2195 (N_2195,N_2051,N_1988);
and U2196 (N_2196,N_2042,N_1839);
and U2197 (N_2197,N_1941,N_2044);
or U2198 (N_2198,N_1963,N_1908);
or U2199 (N_2199,N_1920,N_2010);
xnor U2200 (N_2200,N_2016,N_1852);
nor U2201 (N_2201,N_1964,N_1890);
and U2202 (N_2202,N_2060,N_1911);
or U2203 (N_2203,N_2002,N_1854);
nor U2204 (N_2204,N_1913,N_1877);
and U2205 (N_2205,N_2083,N_1886);
nand U2206 (N_2206,N_2093,N_2027);
and U2207 (N_2207,N_1894,N_1936);
xnor U2208 (N_2208,N_2000,N_2028);
xnor U2209 (N_2209,N_1923,N_1853);
nor U2210 (N_2210,N_2087,N_2097);
and U2211 (N_2211,N_1833,N_1910);
nand U2212 (N_2212,N_2026,N_2030);
and U2213 (N_2213,N_1823,N_1945);
or U2214 (N_2214,N_1859,N_1872);
or U2215 (N_2215,N_1857,N_2005);
or U2216 (N_2216,N_2081,N_1981);
nor U2217 (N_2217,N_1986,N_2003);
and U2218 (N_2218,N_1940,N_1929);
xnor U2219 (N_2219,N_2071,N_1954);
nor U2220 (N_2220,N_1912,N_1932);
nor U2221 (N_2221,N_1878,N_2075);
xor U2222 (N_2222,N_1927,N_2050);
or U2223 (N_2223,N_1863,N_2072);
xor U2224 (N_2224,N_1903,N_2035);
xnor U2225 (N_2225,N_2098,N_1808);
xnor U2226 (N_2226,N_2017,N_1982);
xor U2227 (N_2227,N_1802,N_1846);
nor U2228 (N_2228,N_1882,N_2059);
nor U2229 (N_2229,N_1909,N_2061);
nand U2230 (N_2230,N_2006,N_1942);
or U2231 (N_2231,N_1935,N_1842);
xnor U2232 (N_2232,N_2092,N_1810);
or U2233 (N_2233,N_1934,N_1840);
or U2234 (N_2234,N_2041,N_1967);
and U2235 (N_2235,N_2082,N_1812);
nor U2236 (N_2236,N_1989,N_1804);
nand U2237 (N_2237,N_1993,N_1835);
nand U2238 (N_2238,N_1974,N_2078);
or U2239 (N_2239,N_1922,N_2021);
nor U2240 (N_2240,N_2018,N_2089);
nor U2241 (N_2241,N_1947,N_1959);
and U2242 (N_2242,N_1801,N_1829);
nand U2243 (N_2243,N_1958,N_1995);
xor U2244 (N_2244,N_1915,N_2058);
and U2245 (N_2245,N_1952,N_2040);
nand U2246 (N_2246,N_1985,N_2094);
or U2247 (N_2247,N_2088,N_2063);
or U2248 (N_2248,N_1881,N_1851);
or U2249 (N_2249,N_1831,N_1845);
nor U2250 (N_2250,N_1846,N_2039);
and U2251 (N_2251,N_1988,N_2001);
or U2252 (N_2252,N_2004,N_2062);
and U2253 (N_2253,N_1969,N_1860);
or U2254 (N_2254,N_1958,N_1812);
nor U2255 (N_2255,N_1824,N_2007);
nand U2256 (N_2256,N_2063,N_2028);
or U2257 (N_2257,N_1875,N_2055);
nor U2258 (N_2258,N_1904,N_1811);
xnor U2259 (N_2259,N_1918,N_1914);
and U2260 (N_2260,N_1920,N_2040);
xor U2261 (N_2261,N_2053,N_2085);
nor U2262 (N_2262,N_1816,N_2008);
xor U2263 (N_2263,N_2052,N_1821);
and U2264 (N_2264,N_1899,N_2041);
or U2265 (N_2265,N_1937,N_2071);
nor U2266 (N_2266,N_1952,N_2061);
xnor U2267 (N_2267,N_1893,N_1921);
xor U2268 (N_2268,N_2003,N_1878);
or U2269 (N_2269,N_2050,N_1807);
or U2270 (N_2270,N_1808,N_2066);
xor U2271 (N_2271,N_1904,N_1900);
nor U2272 (N_2272,N_2093,N_1958);
xnor U2273 (N_2273,N_1982,N_1800);
xnor U2274 (N_2274,N_1918,N_1845);
or U2275 (N_2275,N_1874,N_2064);
nand U2276 (N_2276,N_2012,N_2035);
and U2277 (N_2277,N_1860,N_1916);
nand U2278 (N_2278,N_1899,N_2094);
nor U2279 (N_2279,N_1911,N_1859);
xnor U2280 (N_2280,N_2096,N_1826);
or U2281 (N_2281,N_1870,N_2080);
or U2282 (N_2282,N_2004,N_2011);
nor U2283 (N_2283,N_1879,N_1921);
xor U2284 (N_2284,N_2059,N_2066);
nor U2285 (N_2285,N_1938,N_2080);
nand U2286 (N_2286,N_1904,N_1918);
nand U2287 (N_2287,N_2046,N_2074);
nand U2288 (N_2288,N_1987,N_1906);
xnor U2289 (N_2289,N_2059,N_2050);
and U2290 (N_2290,N_1956,N_2079);
or U2291 (N_2291,N_1852,N_1934);
nand U2292 (N_2292,N_1914,N_2010);
xnor U2293 (N_2293,N_1863,N_1828);
or U2294 (N_2294,N_1808,N_1896);
nand U2295 (N_2295,N_1863,N_1928);
and U2296 (N_2296,N_2092,N_1953);
xnor U2297 (N_2297,N_2041,N_1895);
nand U2298 (N_2298,N_2063,N_1919);
and U2299 (N_2299,N_1841,N_2038);
or U2300 (N_2300,N_1930,N_1996);
or U2301 (N_2301,N_1880,N_2023);
xnor U2302 (N_2302,N_2014,N_1963);
and U2303 (N_2303,N_1994,N_1841);
or U2304 (N_2304,N_2086,N_1841);
and U2305 (N_2305,N_1929,N_1817);
nor U2306 (N_2306,N_1973,N_2069);
xor U2307 (N_2307,N_2061,N_2038);
xor U2308 (N_2308,N_1999,N_2027);
xnor U2309 (N_2309,N_1845,N_1886);
or U2310 (N_2310,N_2064,N_2043);
xor U2311 (N_2311,N_2058,N_1940);
nand U2312 (N_2312,N_2000,N_1826);
and U2313 (N_2313,N_2079,N_2047);
or U2314 (N_2314,N_1870,N_2030);
and U2315 (N_2315,N_1837,N_2052);
nor U2316 (N_2316,N_1960,N_1811);
and U2317 (N_2317,N_2094,N_1930);
xnor U2318 (N_2318,N_1835,N_1864);
nor U2319 (N_2319,N_2032,N_1923);
and U2320 (N_2320,N_1935,N_1986);
or U2321 (N_2321,N_1934,N_1978);
xor U2322 (N_2322,N_1902,N_1847);
xor U2323 (N_2323,N_2076,N_2048);
or U2324 (N_2324,N_1892,N_1859);
nand U2325 (N_2325,N_1933,N_1954);
nand U2326 (N_2326,N_1977,N_1957);
and U2327 (N_2327,N_1890,N_1877);
nand U2328 (N_2328,N_1834,N_1807);
xor U2329 (N_2329,N_2018,N_1854);
nand U2330 (N_2330,N_1897,N_1850);
or U2331 (N_2331,N_2020,N_1992);
nand U2332 (N_2332,N_1837,N_1850);
nand U2333 (N_2333,N_2054,N_1830);
and U2334 (N_2334,N_1803,N_1836);
or U2335 (N_2335,N_1958,N_1974);
nor U2336 (N_2336,N_1897,N_2091);
or U2337 (N_2337,N_1961,N_2090);
or U2338 (N_2338,N_2095,N_2063);
or U2339 (N_2339,N_1967,N_1984);
and U2340 (N_2340,N_1844,N_2098);
or U2341 (N_2341,N_1817,N_1849);
and U2342 (N_2342,N_2029,N_1933);
or U2343 (N_2343,N_1890,N_1830);
xnor U2344 (N_2344,N_2028,N_1893);
or U2345 (N_2345,N_2047,N_1979);
and U2346 (N_2346,N_1847,N_1813);
nor U2347 (N_2347,N_2016,N_1974);
and U2348 (N_2348,N_1926,N_2051);
nor U2349 (N_2349,N_1810,N_1891);
and U2350 (N_2350,N_1940,N_1975);
nor U2351 (N_2351,N_2010,N_2003);
xnor U2352 (N_2352,N_2032,N_1855);
nor U2353 (N_2353,N_1974,N_1962);
and U2354 (N_2354,N_1818,N_1972);
xnor U2355 (N_2355,N_1997,N_2093);
and U2356 (N_2356,N_1889,N_2081);
and U2357 (N_2357,N_1810,N_2050);
xor U2358 (N_2358,N_1928,N_2068);
nand U2359 (N_2359,N_2032,N_1881);
or U2360 (N_2360,N_2073,N_1813);
and U2361 (N_2361,N_2000,N_2089);
nand U2362 (N_2362,N_2023,N_1914);
nand U2363 (N_2363,N_1929,N_2042);
nand U2364 (N_2364,N_1994,N_1824);
nor U2365 (N_2365,N_1990,N_1919);
and U2366 (N_2366,N_1868,N_2069);
xnor U2367 (N_2367,N_2016,N_1971);
or U2368 (N_2368,N_1953,N_1835);
nor U2369 (N_2369,N_1974,N_1978);
nor U2370 (N_2370,N_1914,N_2035);
and U2371 (N_2371,N_2012,N_2092);
nor U2372 (N_2372,N_1986,N_1904);
and U2373 (N_2373,N_1971,N_1970);
and U2374 (N_2374,N_1997,N_1927);
xor U2375 (N_2375,N_1821,N_2028);
nor U2376 (N_2376,N_1991,N_1935);
nand U2377 (N_2377,N_1947,N_1896);
nand U2378 (N_2378,N_1984,N_1849);
xor U2379 (N_2379,N_1863,N_1922);
nor U2380 (N_2380,N_1943,N_1874);
xnor U2381 (N_2381,N_1967,N_1908);
nand U2382 (N_2382,N_1927,N_1888);
nand U2383 (N_2383,N_1984,N_1864);
nor U2384 (N_2384,N_1956,N_2049);
nand U2385 (N_2385,N_2065,N_2086);
and U2386 (N_2386,N_2070,N_1980);
nand U2387 (N_2387,N_1887,N_1992);
nor U2388 (N_2388,N_2022,N_1838);
and U2389 (N_2389,N_1906,N_1974);
and U2390 (N_2390,N_1941,N_2055);
nor U2391 (N_2391,N_2086,N_2079);
and U2392 (N_2392,N_1854,N_1995);
or U2393 (N_2393,N_2045,N_2087);
nor U2394 (N_2394,N_1822,N_1812);
nand U2395 (N_2395,N_2049,N_1981);
nor U2396 (N_2396,N_1999,N_1817);
nor U2397 (N_2397,N_1813,N_2039);
nand U2398 (N_2398,N_1833,N_1987);
xor U2399 (N_2399,N_2091,N_1979);
nor U2400 (N_2400,N_2193,N_2235);
nand U2401 (N_2401,N_2137,N_2290);
or U2402 (N_2402,N_2393,N_2103);
nand U2403 (N_2403,N_2231,N_2346);
or U2404 (N_2404,N_2354,N_2398);
or U2405 (N_2405,N_2143,N_2340);
nor U2406 (N_2406,N_2224,N_2311);
xnor U2407 (N_2407,N_2238,N_2180);
xnor U2408 (N_2408,N_2198,N_2306);
nor U2409 (N_2409,N_2121,N_2232);
xnor U2410 (N_2410,N_2247,N_2297);
and U2411 (N_2411,N_2135,N_2164);
xnor U2412 (N_2412,N_2183,N_2120);
nor U2413 (N_2413,N_2347,N_2361);
nor U2414 (N_2414,N_2245,N_2200);
or U2415 (N_2415,N_2329,N_2240);
nand U2416 (N_2416,N_2114,N_2187);
xor U2417 (N_2417,N_2302,N_2156);
and U2418 (N_2418,N_2327,N_2324);
or U2419 (N_2419,N_2378,N_2144);
nor U2420 (N_2420,N_2319,N_2179);
or U2421 (N_2421,N_2229,N_2264);
and U2422 (N_2422,N_2349,N_2374);
nand U2423 (N_2423,N_2281,N_2212);
nand U2424 (N_2424,N_2257,N_2266);
nor U2425 (N_2425,N_2133,N_2182);
nor U2426 (N_2426,N_2351,N_2161);
or U2427 (N_2427,N_2197,N_2333);
and U2428 (N_2428,N_2394,N_2330);
or U2429 (N_2429,N_2313,N_2376);
nor U2430 (N_2430,N_2108,N_2248);
and U2431 (N_2431,N_2256,N_2211);
nor U2432 (N_2432,N_2289,N_2316);
xnor U2433 (N_2433,N_2226,N_2242);
and U2434 (N_2434,N_2317,N_2337);
nor U2435 (N_2435,N_2189,N_2258);
nor U2436 (N_2436,N_2147,N_2388);
nand U2437 (N_2437,N_2140,N_2345);
nand U2438 (N_2438,N_2356,N_2196);
or U2439 (N_2439,N_2308,N_2268);
nand U2440 (N_2440,N_2162,N_2219);
nand U2441 (N_2441,N_2105,N_2335);
or U2442 (N_2442,N_2215,N_2271);
or U2443 (N_2443,N_2358,N_2151);
xnor U2444 (N_2444,N_2288,N_2234);
xnor U2445 (N_2445,N_2186,N_2175);
or U2446 (N_2446,N_2191,N_2125);
nand U2447 (N_2447,N_2102,N_2104);
and U2448 (N_2448,N_2174,N_2385);
xor U2449 (N_2449,N_2241,N_2277);
nor U2450 (N_2450,N_2326,N_2227);
and U2451 (N_2451,N_2254,N_2237);
nor U2452 (N_2452,N_2169,N_2177);
and U2453 (N_2453,N_2357,N_2184);
nor U2454 (N_2454,N_2249,N_2322);
or U2455 (N_2455,N_2305,N_2359);
xnor U2456 (N_2456,N_2221,N_2115);
xnor U2457 (N_2457,N_2368,N_2262);
and U2458 (N_2458,N_2118,N_2298);
nor U2459 (N_2459,N_2263,N_2282);
nor U2460 (N_2460,N_2390,N_2206);
xnor U2461 (N_2461,N_2210,N_2320);
nand U2462 (N_2462,N_2100,N_2339);
nand U2463 (N_2463,N_2158,N_2173);
nor U2464 (N_2464,N_2387,N_2218);
or U2465 (N_2465,N_2209,N_2110);
nor U2466 (N_2466,N_2252,N_2377);
nand U2467 (N_2467,N_2167,N_2286);
or U2468 (N_2468,N_2160,N_2255);
xor U2469 (N_2469,N_2373,N_2278);
xnor U2470 (N_2470,N_2284,N_2294);
and U2471 (N_2471,N_2128,N_2301);
or U2472 (N_2472,N_2343,N_2136);
xnor U2473 (N_2473,N_2287,N_2181);
or U2474 (N_2474,N_2155,N_2134);
or U2475 (N_2475,N_2366,N_2149);
nand U2476 (N_2476,N_2279,N_2190);
nor U2477 (N_2477,N_2381,N_2223);
nor U2478 (N_2478,N_2142,N_2267);
and U2479 (N_2479,N_2230,N_2342);
or U2480 (N_2480,N_2352,N_2157);
or U2481 (N_2481,N_2315,N_2362);
or U2482 (N_2482,N_2127,N_2176);
xor U2483 (N_2483,N_2382,N_2222);
or U2484 (N_2484,N_2396,N_2353);
nand U2485 (N_2485,N_2116,N_2300);
xor U2486 (N_2486,N_2341,N_2204);
nor U2487 (N_2487,N_2269,N_2153);
and U2488 (N_2488,N_2239,N_2380);
or U2489 (N_2489,N_2172,N_2216);
nor U2490 (N_2490,N_2328,N_2274);
nand U2491 (N_2491,N_2233,N_2372);
or U2492 (N_2492,N_2243,N_2228);
or U2493 (N_2493,N_2383,N_2163);
nor U2494 (N_2494,N_2208,N_2109);
or U2495 (N_2495,N_2309,N_2214);
xor U2496 (N_2496,N_2276,N_2365);
and U2497 (N_2497,N_2275,N_2360);
or U2498 (N_2498,N_2131,N_2119);
nand U2499 (N_2499,N_2272,N_2395);
and U2500 (N_2500,N_2168,N_2293);
nor U2501 (N_2501,N_2292,N_2220);
and U2502 (N_2502,N_2217,N_2391);
nor U2503 (N_2503,N_2291,N_2170);
nor U2504 (N_2504,N_2194,N_2130);
nor U2505 (N_2505,N_2379,N_2285);
nor U2506 (N_2506,N_2123,N_2107);
nand U2507 (N_2507,N_2106,N_2250);
nand U2508 (N_2508,N_2205,N_2148);
or U2509 (N_2509,N_2389,N_2203);
and U2510 (N_2510,N_2178,N_2101);
nand U2511 (N_2511,N_2371,N_2132);
xor U2512 (N_2512,N_2325,N_2364);
nor U2513 (N_2513,N_2138,N_2124);
nor U2514 (N_2514,N_2283,N_2207);
xnor U2515 (N_2515,N_2246,N_2312);
nand U2516 (N_2516,N_2338,N_2159);
nand U2517 (N_2517,N_2369,N_2273);
nor U2518 (N_2518,N_2295,N_2185);
nand U2519 (N_2519,N_2165,N_2350);
or U2520 (N_2520,N_2251,N_2129);
and U2521 (N_2521,N_2166,N_2336);
nor U2522 (N_2522,N_2265,N_2126);
nor U2523 (N_2523,N_2392,N_2318);
and U2524 (N_2524,N_2303,N_2355);
and U2525 (N_2525,N_2323,N_2171);
nor U2526 (N_2526,N_2253,N_2375);
or U2527 (N_2527,N_2225,N_2201);
xnor U2528 (N_2528,N_2202,N_2331);
and U2529 (N_2529,N_2188,N_2146);
xor U2530 (N_2530,N_2154,N_2296);
or U2531 (N_2531,N_2141,N_2113);
nor U2532 (N_2532,N_2304,N_2244);
and U2533 (N_2533,N_2270,N_2111);
nor U2534 (N_2534,N_2145,N_2363);
and U2535 (N_2535,N_2150,N_2259);
xnor U2536 (N_2536,N_2299,N_2260);
or U2537 (N_2537,N_2367,N_2384);
nand U2538 (N_2538,N_2310,N_2370);
nor U2539 (N_2539,N_2307,N_2261);
or U2540 (N_2540,N_2195,N_2139);
nor U2541 (N_2541,N_2348,N_2192);
and U2542 (N_2542,N_2152,N_2213);
nor U2543 (N_2543,N_2397,N_2122);
nor U2544 (N_2544,N_2314,N_2321);
xor U2545 (N_2545,N_2199,N_2399);
nor U2546 (N_2546,N_2236,N_2386);
nor U2547 (N_2547,N_2112,N_2332);
or U2548 (N_2548,N_2117,N_2280);
xnor U2549 (N_2549,N_2344,N_2334);
and U2550 (N_2550,N_2132,N_2365);
and U2551 (N_2551,N_2114,N_2397);
or U2552 (N_2552,N_2165,N_2122);
nand U2553 (N_2553,N_2254,N_2160);
and U2554 (N_2554,N_2385,N_2212);
nor U2555 (N_2555,N_2165,N_2130);
or U2556 (N_2556,N_2177,N_2389);
and U2557 (N_2557,N_2305,N_2342);
or U2558 (N_2558,N_2148,N_2293);
and U2559 (N_2559,N_2293,N_2253);
nand U2560 (N_2560,N_2250,N_2165);
or U2561 (N_2561,N_2321,N_2123);
nor U2562 (N_2562,N_2210,N_2311);
nor U2563 (N_2563,N_2228,N_2315);
or U2564 (N_2564,N_2199,N_2347);
xor U2565 (N_2565,N_2119,N_2301);
or U2566 (N_2566,N_2193,N_2223);
xor U2567 (N_2567,N_2341,N_2112);
nand U2568 (N_2568,N_2396,N_2300);
and U2569 (N_2569,N_2265,N_2361);
nand U2570 (N_2570,N_2265,N_2110);
xor U2571 (N_2571,N_2269,N_2300);
and U2572 (N_2572,N_2125,N_2250);
nand U2573 (N_2573,N_2254,N_2316);
nand U2574 (N_2574,N_2156,N_2399);
nor U2575 (N_2575,N_2124,N_2202);
nand U2576 (N_2576,N_2286,N_2101);
nor U2577 (N_2577,N_2118,N_2247);
or U2578 (N_2578,N_2155,N_2372);
xor U2579 (N_2579,N_2294,N_2289);
or U2580 (N_2580,N_2157,N_2107);
or U2581 (N_2581,N_2259,N_2190);
and U2582 (N_2582,N_2317,N_2350);
and U2583 (N_2583,N_2111,N_2217);
xnor U2584 (N_2584,N_2334,N_2261);
xnor U2585 (N_2585,N_2324,N_2392);
nand U2586 (N_2586,N_2356,N_2197);
or U2587 (N_2587,N_2272,N_2187);
nor U2588 (N_2588,N_2132,N_2360);
and U2589 (N_2589,N_2254,N_2155);
xnor U2590 (N_2590,N_2327,N_2319);
nand U2591 (N_2591,N_2244,N_2155);
nand U2592 (N_2592,N_2309,N_2282);
nor U2593 (N_2593,N_2297,N_2274);
and U2594 (N_2594,N_2395,N_2285);
or U2595 (N_2595,N_2280,N_2247);
nand U2596 (N_2596,N_2261,N_2218);
or U2597 (N_2597,N_2161,N_2315);
nand U2598 (N_2598,N_2172,N_2267);
nand U2599 (N_2599,N_2185,N_2388);
nor U2600 (N_2600,N_2245,N_2396);
nor U2601 (N_2601,N_2100,N_2365);
nand U2602 (N_2602,N_2218,N_2234);
xor U2603 (N_2603,N_2387,N_2196);
and U2604 (N_2604,N_2198,N_2109);
nand U2605 (N_2605,N_2387,N_2202);
and U2606 (N_2606,N_2160,N_2345);
xor U2607 (N_2607,N_2377,N_2129);
xnor U2608 (N_2608,N_2399,N_2326);
nor U2609 (N_2609,N_2130,N_2267);
or U2610 (N_2610,N_2123,N_2330);
nor U2611 (N_2611,N_2399,N_2250);
xnor U2612 (N_2612,N_2175,N_2268);
or U2613 (N_2613,N_2264,N_2212);
or U2614 (N_2614,N_2309,N_2114);
xnor U2615 (N_2615,N_2350,N_2308);
nor U2616 (N_2616,N_2325,N_2356);
nor U2617 (N_2617,N_2205,N_2343);
or U2618 (N_2618,N_2392,N_2389);
nand U2619 (N_2619,N_2304,N_2202);
and U2620 (N_2620,N_2363,N_2399);
nand U2621 (N_2621,N_2300,N_2148);
and U2622 (N_2622,N_2154,N_2120);
nor U2623 (N_2623,N_2196,N_2385);
nor U2624 (N_2624,N_2362,N_2148);
and U2625 (N_2625,N_2113,N_2148);
nand U2626 (N_2626,N_2302,N_2376);
xor U2627 (N_2627,N_2303,N_2146);
xor U2628 (N_2628,N_2167,N_2128);
nor U2629 (N_2629,N_2246,N_2172);
nand U2630 (N_2630,N_2338,N_2317);
and U2631 (N_2631,N_2101,N_2149);
nor U2632 (N_2632,N_2136,N_2219);
and U2633 (N_2633,N_2380,N_2390);
xnor U2634 (N_2634,N_2245,N_2188);
and U2635 (N_2635,N_2394,N_2196);
nand U2636 (N_2636,N_2303,N_2357);
nand U2637 (N_2637,N_2273,N_2169);
nand U2638 (N_2638,N_2195,N_2303);
or U2639 (N_2639,N_2159,N_2129);
and U2640 (N_2640,N_2225,N_2270);
or U2641 (N_2641,N_2146,N_2204);
and U2642 (N_2642,N_2130,N_2303);
xor U2643 (N_2643,N_2200,N_2159);
nor U2644 (N_2644,N_2155,N_2327);
and U2645 (N_2645,N_2290,N_2317);
xnor U2646 (N_2646,N_2120,N_2241);
or U2647 (N_2647,N_2224,N_2119);
nor U2648 (N_2648,N_2217,N_2252);
and U2649 (N_2649,N_2211,N_2347);
nand U2650 (N_2650,N_2294,N_2392);
xnor U2651 (N_2651,N_2217,N_2173);
or U2652 (N_2652,N_2215,N_2135);
xnor U2653 (N_2653,N_2160,N_2199);
nand U2654 (N_2654,N_2244,N_2279);
nor U2655 (N_2655,N_2167,N_2370);
nor U2656 (N_2656,N_2100,N_2122);
or U2657 (N_2657,N_2342,N_2163);
nand U2658 (N_2658,N_2221,N_2305);
xnor U2659 (N_2659,N_2338,N_2395);
or U2660 (N_2660,N_2219,N_2259);
or U2661 (N_2661,N_2308,N_2169);
and U2662 (N_2662,N_2273,N_2287);
nand U2663 (N_2663,N_2151,N_2388);
or U2664 (N_2664,N_2238,N_2136);
or U2665 (N_2665,N_2114,N_2347);
nor U2666 (N_2666,N_2229,N_2141);
xor U2667 (N_2667,N_2121,N_2162);
xnor U2668 (N_2668,N_2217,N_2313);
nand U2669 (N_2669,N_2335,N_2174);
xnor U2670 (N_2670,N_2318,N_2176);
or U2671 (N_2671,N_2224,N_2255);
nand U2672 (N_2672,N_2324,N_2338);
xnor U2673 (N_2673,N_2141,N_2184);
or U2674 (N_2674,N_2158,N_2365);
xor U2675 (N_2675,N_2200,N_2326);
nor U2676 (N_2676,N_2157,N_2387);
or U2677 (N_2677,N_2281,N_2331);
xor U2678 (N_2678,N_2128,N_2162);
xnor U2679 (N_2679,N_2288,N_2251);
nand U2680 (N_2680,N_2267,N_2311);
xor U2681 (N_2681,N_2180,N_2354);
nand U2682 (N_2682,N_2203,N_2107);
or U2683 (N_2683,N_2186,N_2392);
xnor U2684 (N_2684,N_2331,N_2219);
and U2685 (N_2685,N_2283,N_2279);
and U2686 (N_2686,N_2380,N_2109);
xnor U2687 (N_2687,N_2244,N_2325);
and U2688 (N_2688,N_2278,N_2143);
and U2689 (N_2689,N_2197,N_2385);
xor U2690 (N_2690,N_2186,N_2119);
nand U2691 (N_2691,N_2234,N_2107);
and U2692 (N_2692,N_2198,N_2144);
or U2693 (N_2693,N_2378,N_2354);
xor U2694 (N_2694,N_2333,N_2111);
xnor U2695 (N_2695,N_2168,N_2364);
xor U2696 (N_2696,N_2141,N_2398);
xnor U2697 (N_2697,N_2266,N_2341);
and U2698 (N_2698,N_2222,N_2304);
xnor U2699 (N_2699,N_2271,N_2209);
or U2700 (N_2700,N_2502,N_2558);
nand U2701 (N_2701,N_2404,N_2601);
xnor U2702 (N_2702,N_2631,N_2623);
nor U2703 (N_2703,N_2581,N_2605);
nand U2704 (N_2704,N_2509,N_2507);
xnor U2705 (N_2705,N_2456,N_2465);
xnor U2706 (N_2706,N_2542,N_2685);
nand U2707 (N_2707,N_2400,N_2467);
nand U2708 (N_2708,N_2622,N_2614);
or U2709 (N_2709,N_2490,N_2649);
or U2710 (N_2710,N_2556,N_2669);
nand U2711 (N_2711,N_2666,N_2479);
and U2712 (N_2712,N_2487,N_2615);
xor U2713 (N_2713,N_2547,N_2608);
or U2714 (N_2714,N_2634,N_2651);
nand U2715 (N_2715,N_2571,N_2667);
and U2716 (N_2716,N_2568,N_2443);
nand U2717 (N_2717,N_2682,N_2475);
and U2718 (N_2718,N_2514,N_2532);
nor U2719 (N_2719,N_2551,N_2597);
or U2720 (N_2720,N_2493,N_2526);
nand U2721 (N_2721,N_2454,N_2549);
or U2722 (N_2722,N_2693,N_2470);
and U2723 (N_2723,N_2662,N_2471);
and U2724 (N_2724,N_2476,N_2648);
nand U2725 (N_2725,N_2539,N_2530);
nand U2726 (N_2726,N_2420,N_2508);
xor U2727 (N_2727,N_2450,N_2403);
or U2728 (N_2728,N_2655,N_2408);
or U2729 (N_2729,N_2447,N_2519);
or U2730 (N_2730,N_2644,N_2598);
or U2731 (N_2731,N_2537,N_2457);
nor U2732 (N_2732,N_2632,N_2441);
nor U2733 (N_2733,N_2533,N_2591);
xnor U2734 (N_2734,N_2690,N_2550);
and U2735 (N_2735,N_2694,N_2676);
nor U2736 (N_2736,N_2458,N_2495);
xor U2737 (N_2737,N_2638,N_2430);
or U2738 (N_2738,N_2670,N_2578);
nand U2739 (N_2739,N_2660,N_2401);
xnor U2740 (N_2740,N_2405,N_2566);
and U2741 (N_2741,N_2580,N_2496);
xor U2742 (N_2742,N_2672,N_2462);
nand U2743 (N_2743,N_2505,N_2469);
or U2744 (N_2744,N_2427,N_2659);
or U2745 (N_2745,N_2562,N_2482);
nor U2746 (N_2746,N_2413,N_2423);
nor U2747 (N_2747,N_2517,N_2645);
or U2748 (N_2748,N_2610,N_2654);
and U2749 (N_2749,N_2503,N_2576);
nand U2750 (N_2750,N_2411,N_2563);
nand U2751 (N_2751,N_2663,N_2483);
and U2752 (N_2752,N_2545,N_2497);
xnor U2753 (N_2753,N_2438,N_2442);
nand U2754 (N_2754,N_2553,N_2692);
nand U2755 (N_2755,N_2602,N_2536);
or U2756 (N_2756,N_2565,N_2582);
xor U2757 (N_2757,N_2491,N_2414);
xor U2758 (N_2758,N_2445,N_2574);
nor U2759 (N_2759,N_2513,N_2531);
and U2760 (N_2760,N_2573,N_2646);
and U2761 (N_2761,N_2521,N_2436);
or U2762 (N_2762,N_2524,N_2455);
or U2763 (N_2763,N_2415,N_2599);
xor U2764 (N_2764,N_2564,N_2675);
or U2765 (N_2765,N_2624,N_2681);
or U2766 (N_2766,N_2554,N_2589);
xor U2767 (N_2767,N_2665,N_2656);
xor U2768 (N_2768,N_2637,N_2461);
or U2769 (N_2769,N_2439,N_2674);
nand U2770 (N_2770,N_2525,N_2612);
xnor U2771 (N_2771,N_2680,N_2412);
or U2772 (N_2772,N_2689,N_2595);
nor U2773 (N_2773,N_2544,N_2506);
and U2774 (N_2774,N_2643,N_2588);
or U2775 (N_2775,N_2688,N_2647);
xor U2776 (N_2776,N_2501,N_2569);
or U2777 (N_2777,N_2579,N_2687);
and U2778 (N_2778,N_2636,N_2590);
and U2779 (N_2779,N_2583,N_2468);
and U2780 (N_2780,N_2575,N_2419);
or U2781 (N_2781,N_2440,N_2606);
xnor U2782 (N_2782,N_2489,N_2486);
xnor U2783 (N_2783,N_2431,N_2673);
nand U2784 (N_2784,N_2668,N_2604);
nand U2785 (N_2785,N_2616,N_2686);
and U2786 (N_2786,N_2621,N_2480);
or U2787 (N_2787,N_2592,N_2548);
nand U2788 (N_2788,N_2584,N_2609);
xor U2789 (N_2789,N_2485,N_2620);
xnor U2790 (N_2790,N_2652,N_2640);
nand U2791 (N_2791,N_2698,N_2488);
nor U2792 (N_2792,N_2464,N_2658);
nand U2793 (N_2793,N_2407,N_2500);
xnor U2794 (N_2794,N_2452,N_2552);
nor U2795 (N_2795,N_2546,N_2463);
or U2796 (N_2796,N_2516,N_2515);
nand U2797 (N_2797,N_2600,N_2619);
nor U2798 (N_2798,N_2661,N_2504);
xnor U2799 (N_2799,N_2697,N_2679);
or U2800 (N_2800,N_2699,N_2429);
and U2801 (N_2801,N_2529,N_2460);
xor U2802 (N_2802,N_2523,N_2633);
and U2803 (N_2803,N_2555,N_2474);
xor U2804 (N_2804,N_2630,N_2664);
nor U2805 (N_2805,N_2473,N_2653);
and U2806 (N_2806,N_2444,N_2593);
nor U2807 (N_2807,N_2511,N_2421);
or U2808 (N_2808,N_2557,N_2696);
nand U2809 (N_2809,N_2435,N_2684);
xnor U2810 (N_2810,N_2424,N_2522);
and U2811 (N_2811,N_2434,N_2535);
nor U2812 (N_2812,N_2498,N_2409);
or U2813 (N_2813,N_2418,N_2446);
or U2814 (N_2814,N_2428,N_2540);
nand U2815 (N_2815,N_2466,N_2639);
nor U2816 (N_2816,N_2437,N_2560);
or U2817 (N_2817,N_2406,N_2432);
nand U2818 (N_2818,N_2541,N_2410);
nand U2819 (N_2819,N_2499,N_2534);
or U2820 (N_2820,N_2425,N_2478);
or U2821 (N_2821,N_2585,N_2449);
and U2822 (N_2822,N_2657,N_2618);
xor U2823 (N_2823,N_2433,N_2459);
xnor U2824 (N_2824,N_2617,N_2671);
xor U2825 (N_2825,N_2484,N_2538);
nand U2826 (N_2826,N_2625,N_2543);
nor U2827 (N_2827,N_2611,N_2561);
nand U2828 (N_2828,N_2629,N_2577);
or U2829 (N_2829,N_2627,N_2510);
or U2830 (N_2830,N_2641,N_2520);
and U2831 (N_2831,N_2613,N_2518);
and U2832 (N_2832,N_2607,N_2572);
xor U2833 (N_2833,N_2416,N_2422);
xnor U2834 (N_2834,N_2642,N_2448);
nor U2835 (N_2835,N_2512,N_2453);
or U2836 (N_2836,N_2586,N_2472);
nor U2837 (N_2837,N_2570,N_2494);
xor U2838 (N_2838,N_2628,N_2528);
nor U2839 (N_2839,N_2451,N_2626);
nor U2840 (N_2840,N_2477,N_2635);
or U2841 (N_2841,N_2678,N_2481);
xor U2842 (N_2842,N_2650,N_2596);
xnor U2843 (N_2843,N_2426,N_2559);
xor U2844 (N_2844,N_2567,N_2587);
and U2845 (N_2845,N_2527,N_2683);
or U2846 (N_2846,N_2402,N_2677);
xor U2847 (N_2847,N_2492,N_2417);
nor U2848 (N_2848,N_2695,N_2603);
xor U2849 (N_2849,N_2594,N_2691);
and U2850 (N_2850,N_2431,N_2429);
or U2851 (N_2851,N_2677,N_2585);
nor U2852 (N_2852,N_2504,N_2531);
xor U2853 (N_2853,N_2484,N_2689);
xor U2854 (N_2854,N_2569,N_2540);
or U2855 (N_2855,N_2511,N_2467);
xnor U2856 (N_2856,N_2646,N_2513);
nor U2857 (N_2857,N_2564,N_2437);
xnor U2858 (N_2858,N_2598,N_2680);
xnor U2859 (N_2859,N_2579,N_2441);
and U2860 (N_2860,N_2602,N_2638);
nand U2861 (N_2861,N_2619,N_2679);
and U2862 (N_2862,N_2476,N_2675);
nand U2863 (N_2863,N_2453,N_2525);
nor U2864 (N_2864,N_2475,N_2667);
nor U2865 (N_2865,N_2425,N_2528);
nor U2866 (N_2866,N_2504,N_2500);
xnor U2867 (N_2867,N_2500,N_2562);
or U2868 (N_2868,N_2442,N_2555);
and U2869 (N_2869,N_2535,N_2520);
xnor U2870 (N_2870,N_2602,N_2673);
or U2871 (N_2871,N_2544,N_2469);
nor U2872 (N_2872,N_2437,N_2696);
or U2873 (N_2873,N_2567,N_2564);
and U2874 (N_2874,N_2584,N_2465);
and U2875 (N_2875,N_2603,N_2457);
nand U2876 (N_2876,N_2699,N_2496);
and U2877 (N_2877,N_2419,N_2644);
or U2878 (N_2878,N_2476,N_2616);
and U2879 (N_2879,N_2541,N_2457);
and U2880 (N_2880,N_2553,N_2656);
or U2881 (N_2881,N_2406,N_2580);
nor U2882 (N_2882,N_2633,N_2577);
or U2883 (N_2883,N_2662,N_2534);
nand U2884 (N_2884,N_2697,N_2643);
nor U2885 (N_2885,N_2573,N_2430);
nand U2886 (N_2886,N_2524,N_2493);
and U2887 (N_2887,N_2413,N_2691);
and U2888 (N_2888,N_2451,N_2563);
xnor U2889 (N_2889,N_2476,N_2451);
and U2890 (N_2890,N_2493,N_2580);
and U2891 (N_2891,N_2655,N_2679);
and U2892 (N_2892,N_2570,N_2576);
or U2893 (N_2893,N_2519,N_2562);
xor U2894 (N_2894,N_2440,N_2548);
xnor U2895 (N_2895,N_2455,N_2539);
nand U2896 (N_2896,N_2504,N_2639);
and U2897 (N_2897,N_2622,N_2584);
nor U2898 (N_2898,N_2466,N_2445);
nand U2899 (N_2899,N_2693,N_2650);
nand U2900 (N_2900,N_2495,N_2471);
xor U2901 (N_2901,N_2614,N_2581);
and U2902 (N_2902,N_2584,N_2667);
or U2903 (N_2903,N_2481,N_2485);
and U2904 (N_2904,N_2507,N_2471);
nand U2905 (N_2905,N_2404,N_2449);
nor U2906 (N_2906,N_2610,N_2529);
or U2907 (N_2907,N_2626,N_2520);
nor U2908 (N_2908,N_2429,N_2469);
xnor U2909 (N_2909,N_2484,N_2442);
or U2910 (N_2910,N_2677,N_2607);
or U2911 (N_2911,N_2508,N_2464);
and U2912 (N_2912,N_2449,N_2677);
nor U2913 (N_2913,N_2639,N_2650);
nand U2914 (N_2914,N_2590,N_2694);
or U2915 (N_2915,N_2454,N_2403);
nand U2916 (N_2916,N_2482,N_2602);
nor U2917 (N_2917,N_2621,N_2489);
and U2918 (N_2918,N_2445,N_2501);
or U2919 (N_2919,N_2503,N_2690);
or U2920 (N_2920,N_2526,N_2549);
and U2921 (N_2921,N_2616,N_2519);
xnor U2922 (N_2922,N_2686,N_2517);
nor U2923 (N_2923,N_2674,N_2429);
xnor U2924 (N_2924,N_2424,N_2476);
nor U2925 (N_2925,N_2609,N_2449);
and U2926 (N_2926,N_2651,N_2421);
or U2927 (N_2927,N_2642,N_2634);
nand U2928 (N_2928,N_2424,N_2543);
nand U2929 (N_2929,N_2578,N_2520);
and U2930 (N_2930,N_2698,N_2678);
nand U2931 (N_2931,N_2599,N_2479);
nor U2932 (N_2932,N_2570,N_2686);
or U2933 (N_2933,N_2567,N_2673);
xnor U2934 (N_2934,N_2607,N_2445);
and U2935 (N_2935,N_2493,N_2624);
or U2936 (N_2936,N_2424,N_2451);
xor U2937 (N_2937,N_2670,N_2581);
and U2938 (N_2938,N_2649,N_2611);
nand U2939 (N_2939,N_2417,N_2528);
nand U2940 (N_2940,N_2582,N_2617);
nor U2941 (N_2941,N_2439,N_2668);
and U2942 (N_2942,N_2477,N_2451);
nand U2943 (N_2943,N_2628,N_2673);
xor U2944 (N_2944,N_2409,N_2428);
nand U2945 (N_2945,N_2525,N_2616);
xor U2946 (N_2946,N_2475,N_2665);
and U2947 (N_2947,N_2612,N_2578);
nor U2948 (N_2948,N_2460,N_2426);
nand U2949 (N_2949,N_2671,N_2665);
and U2950 (N_2950,N_2429,N_2525);
and U2951 (N_2951,N_2489,N_2636);
or U2952 (N_2952,N_2667,N_2646);
nand U2953 (N_2953,N_2403,N_2437);
nand U2954 (N_2954,N_2454,N_2684);
or U2955 (N_2955,N_2642,N_2691);
xnor U2956 (N_2956,N_2460,N_2546);
nor U2957 (N_2957,N_2614,N_2679);
or U2958 (N_2958,N_2534,N_2606);
xor U2959 (N_2959,N_2487,N_2458);
xor U2960 (N_2960,N_2465,N_2630);
nand U2961 (N_2961,N_2423,N_2635);
and U2962 (N_2962,N_2447,N_2616);
and U2963 (N_2963,N_2625,N_2464);
and U2964 (N_2964,N_2424,N_2488);
nor U2965 (N_2965,N_2444,N_2579);
or U2966 (N_2966,N_2555,N_2486);
or U2967 (N_2967,N_2675,N_2614);
or U2968 (N_2968,N_2465,N_2518);
nor U2969 (N_2969,N_2493,N_2560);
xor U2970 (N_2970,N_2416,N_2602);
and U2971 (N_2971,N_2611,N_2622);
xor U2972 (N_2972,N_2595,N_2611);
and U2973 (N_2973,N_2575,N_2503);
and U2974 (N_2974,N_2430,N_2489);
nand U2975 (N_2975,N_2460,N_2693);
nand U2976 (N_2976,N_2431,N_2419);
nand U2977 (N_2977,N_2457,N_2426);
nor U2978 (N_2978,N_2451,N_2677);
and U2979 (N_2979,N_2487,N_2508);
and U2980 (N_2980,N_2542,N_2412);
nor U2981 (N_2981,N_2668,N_2663);
nor U2982 (N_2982,N_2435,N_2511);
nor U2983 (N_2983,N_2634,N_2413);
and U2984 (N_2984,N_2498,N_2653);
nor U2985 (N_2985,N_2551,N_2408);
nor U2986 (N_2986,N_2458,N_2608);
nand U2987 (N_2987,N_2652,N_2515);
nand U2988 (N_2988,N_2499,N_2575);
nand U2989 (N_2989,N_2581,N_2689);
nand U2990 (N_2990,N_2609,N_2467);
nand U2991 (N_2991,N_2489,N_2635);
nor U2992 (N_2992,N_2533,N_2500);
and U2993 (N_2993,N_2656,N_2440);
xor U2994 (N_2994,N_2579,N_2562);
and U2995 (N_2995,N_2662,N_2619);
nor U2996 (N_2996,N_2547,N_2424);
nand U2997 (N_2997,N_2500,N_2517);
and U2998 (N_2998,N_2650,N_2502);
or U2999 (N_2999,N_2518,N_2485);
nor U3000 (N_3000,N_2704,N_2803);
and U3001 (N_3001,N_2915,N_2883);
nand U3002 (N_3002,N_2969,N_2921);
or U3003 (N_3003,N_2901,N_2916);
nand U3004 (N_3004,N_2760,N_2991);
nor U3005 (N_3005,N_2979,N_2796);
or U3006 (N_3006,N_2876,N_2867);
or U3007 (N_3007,N_2759,N_2936);
nor U3008 (N_3008,N_2963,N_2944);
or U3009 (N_3009,N_2861,N_2930);
nor U3010 (N_3010,N_2838,N_2855);
or U3011 (N_3011,N_2931,N_2767);
nand U3012 (N_3012,N_2721,N_2998);
nor U3013 (N_3013,N_2938,N_2731);
nor U3014 (N_3014,N_2715,N_2892);
nor U3015 (N_3015,N_2911,N_2972);
nor U3016 (N_3016,N_2987,N_2942);
nor U3017 (N_3017,N_2776,N_2723);
xnor U3018 (N_3018,N_2889,N_2707);
nor U3019 (N_3019,N_2872,N_2977);
nand U3020 (N_3020,N_2917,N_2780);
nor U3021 (N_3021,N_2877,N_2836);
and U3022 (N_3022,N_2737,N_2899);
and U3023 (N_3023,N_2860,N_2758);
xor U3024 (N_3024,N_2850,N_2747);
nor U3025 (N_3025,N_2761,N_2837);
and U3026 (N_3026,N_2878,N_2880);
or U3027 (N_3027,N_2852,N_2881);
nand U3028 (N_3028,N_2959,N_2802);
nand U3029 (N_3029,N_2742,N_2799);
xnor U3030 (N_3030,N_2893,N_2920);
nor U3031 (N_3031,N_2726,N_2912);
or U3032 (N_3032,N_2885,N_2790);
xnor U3033 (N_3033,N_2750,N_2706);
and U3034 (N_3034,N_2830,N_2862);
nor U3035 (N_3035,N_2978,N_2735);
xor U3036 (N_3036,N_2933,N_2918);
and U3037 (N_3037,N_2774,N_2746);
and U3038 (N_3038,N_2951,N_2962);
or U3039 (N_3039,N_2762,N_2809);
nor U3040 (N_3040,N_2995,N_2713);
and U3041 (N_3041,N_2795,N_2829);
nor U3042 (N_3042,N_2820,N_2833);
nor U3043 (N_3043,N_2903,N_2784);
or U3044 (N_3044,N_2769,N_2958);
or U3045 (N_3045,N_2716,N_2816);
nor U3046 (N_3046,N_2886,N_2992);
and U3047 (N_3047,N_2826,N_2825);
and U3048 (N_3048,N_2801,N_2905);
or U3049 (N_3049,N_2840,N_2924);
or U3050 (N_3050,N_2763,N_2770);
and U3051 (N_3051,N_2981,N_2922);
nor U3052 (N_3052,N_2971,N_2711);
xnor U3053 (N_3053,N_2908,N_2973);
nand U3054 (N_3054,N_2884,N_2729);
or U3055 (N_3055,N_2794,N_2964);
and U3056 (N_3056,N_2874,N_2974);
xor U3057 (N_3057,N_2875,N_2976);
xnor U3058 (N_3058,N_2736,N_2775);
and U3059 (N_3059,N_2772,N_2719);
nor U3060 (N_3060,N_2965,N_2900);
and U3061 (N_3061,N_2858,N_2952);
or U3062 (N_3062,N_2823,N_2907);
nor U3063 (N_3063,N_2859,N_2813);
or U3064 (N_3064,N_2714,N_2902);
nor U3065 (N_3065,N_2919,N_2941);
and U3066 (N_3066,N_2984,N_2946);
xnor U3067 (N_3067,N_2935,N_2817);
xnor U3068 (N_3068,N_2705,N_2989);
xor U3069 (N_3069,N_2841,N_2843);
or U3070 (N_3070,N_2948,N_2755);
xnor U3071 (N_3071,N_2819,N_2822);
nor U3072 (N_3072,N_2847,N_2785);
or U3073 (N_3073,N_2864,N_2845);
nand U3074 (N_3074,N_2894,N_2909);
nor U3075 (N_3075,N_2831,N_2710);
or U3076 (N_3076,N_2844,N_2734);
nand U3077 (N_3077,N_2709,N_2990);
nor U3078 (N_3078,N_2994,N_2955);
or U3079 (N_3079,N_2939,N_2999);
xor U3080 (N_3080,N_2882,N_2814);
xor U3081 (N_3081,N_2961,N_2754);
nand U3082 (N_3082,N_2708,N_2738);
or U3083 (N_3083,N_2842,N_2828);
nand U3084 (N_3084,N_2722,N_2777);
nand U3085 (N_3085,N_2914,N_2786);
nor U3086 (N_3086,N_2748,N_2787);
nor U3087 (N_3087,N_2986,N_2753);
nor U3088 (N_3088,N_2848,N_2895);
nand U3089 (N_3089,N_2967,N_2792);
and U3090 (N_3090,N_2839,N_2732);
or U3091 (N_3091,N_2749,N_2804);
nand U3092 (N_3092,N_2863,N_2857);
and U3093 (N_3093,N_2988,N_2851);
xor U3094 (N_3094,N_2879,N_2827);
or U3095 (N_3095,N_2788,N_2727);
nor U3096 (N_3096,N_2771,N_2997);
nand U3097 (N_3097,N_2764,N_2712);
nor U3098 (N_3098,N_2756,N_2954);
and U3099 (N_3099,N_2791,N_2983);
and U3100 (N_3100,N_2773,N_2751);
nand U3101 (N_3101,N_2993,N_2929);
xnor U3102 (N_3102,N_2868,N_2904);
nor U3103 (N_3103,N_2743,N_2937);
and U3104 (N_3104,N_2778,N_2783);
or U3105 (N_3105,N_2725,N_2968);
nand U3106 (N_3106,N_2730,N_2949);
nand U3107 (N_3107,N_2865,N_2806);
xnor U3108 (N_3108,N_2970,N_2888);
xor U3109 (N_3109,N_2849,N_2797);
or U3110 (N_3110,N_2856,N_2744);
or U3111 (N_3111,N_2781,N_2724);
nand U3112 (N_3112,N_2871,N_2869);
or U3113 (N_3113,N_2824,N_2975);
nand U3114 (N_3114,N_2940,N_2812);
nor U3115 (N_3115,N_2779,N_2789);
nor U3116 (N_3116,N_2811,N_2947);
and U3117 (N_3117,N_2782,N_2835);
or U3118 (N_3118,N_2980,N_2701);
nand U3119 (N_3119,N_2805,N_2702);
xnor U3120 (N_3120,N_2891,N_2740);
nor U3121 (N_3121,N_2739,N_2818);
and U3122 (N_3122,N_2926,N_2718);
and U3123 (N_3123,N_2728,N_2925);
nor U3124 (N_3124,N_2923,N_2898);
nor U3125 (N_3125,N_2866,N_2810);
and U3126 (N_3126,N_2793,N_2953);
nand U3127 (N_3127,N_2897,N_2800);
nor U3128 (N_3128,N_2910,N_2766);
nor U3129 (N_3129,N_2741,N_2745);
xnor U3130 (N_3130,N_2720,N_2932);
nand U3131 (N_3131,N_2957,N_2945);
or U3132 (N_3132,N_2913,N_2928);
and U3133 (N_3133,N_2815,N_2807);
xor U3134 (N_3134,N_2834,N_2985);
nand U3135 (N_3135,N_2768,N_2808);
and U3136 (N_3136,N_2927,N_2982);
nand U3137 (N_3137,N_2700,N_2890);
or U3138 (N_3138,N_2950,N_2765);
xnor U3139 (N_3139,N_2854,N_2934);
nor U3140 (N_3140,N_2757,N_2966);
xor U3141 (N_3141,N_2853,N_2887);
xnor U3142 (N_3142,N_2956,N_2906);
nand U3143 (N_3143,N_2846,N_2752);
nand U3144 (N_3144,N_2960,N_2996);
xor U3145 (N_3145,N_2873,N_2870);
nor U3146 (N_3146,N_2943,N_2703);
xnor U3147 (N_3147,N_2798,N_2832);
xnor U3148 (N_3148,N_2717,N_2896);
and U3149 (N_3149,N_2733,N_2821);
nor U3150 (N_3150,N_2903,N_2864);
nor U3151 (N_3151,N_2869,N_2803);
or U3152 (N_3152,N_2807,N_2957);
or U3153 (N_3153,N_2791,N_2836);
nand U3154 (N_3154,N_2883,N_2705);
or U3155 (N_3155,N_2941,N_2816);
or U3156 (N_3156,N_2828,N_2873);
or U3157 (N_3157,N_2748,N_2892);
and U3158 (N_3158,N_2964,N_2910);
nor U3159 (N_3159,N_2772,N_2789);
xnor U3160 (N_3160,N_2739,N_2944);
nor U3161 (N_3161,N_2827,N_2848);
and U3162 (N_3162,N_2710,N_2990);
nor U3163 (N_3163,N_2982,N_2891);
or U3164 (N_3164,N_2902,N_2995);
and U3165 (N_3165,N_2780,N_2796);
nor U3166 (N_3166,N_2860,N_2730);
or U3167 (N_3167,N_2785,N_2763);
nand U3168 (N_3168,N_2801,N_2873);
nand U3169 (N_3169,N_2982,N_2788);
and U3170 (N_3170,N_2909,N_2782);
nor U3171 (N_3171,N_2863,N_2883);
nor U3172 (N_3172,N_2956,N_2932);
xor U3173 (N_3173,N_2974,N_2960);
nand U3174 (N_3174,N_2890,N_2869);
nand U3175 (N_3175,N_2933,N_2743);
xor U3176 (N_3176,N_2718,N_2949);
or U3177 (N_3177,N_2904,N_2728);
nor U3178 (N_3178,N_2879,N_2761);
nor U3179 (N_3179,N_2915,N_2775);
nand U3180 (N_3180,N_2802,N_2993);
nand U3181 (N_3181,N_2776,N_2993);
nor U3182 (N_3182,N_2893,N_2705);
xnor U3183 (N_3183,N_2988,N_2997);
xor U3184 (N_3184,N_2818,N_2709);
and U3185 (N_3185,N_2929,N_2998);
xor U3186 (N_3186,N_2795,N_2943);
nand U3187 (N_3187,N_2893,N_2720);
nand U3188 (N_3188,N_2972,N_2714);
xnor U3189 (N_3189,N_2808,N_2867);
nor U3190 (N_3190,N_2714,N_2903);
and U3191 (N_3191,N_2715,N_2858);
nand U3192 (N_3192,N_2876,N_2888);
and U3193 (N_3193,N_2798,N_2910);
or U3194 (N_3194,N_2803,N_2955);
or U3195 (N_3195,N_2981,N_2898);
xor U3196 (N_3196,N_2762,N_2726);
and U3197 (N_3197,N_2835,N_2940);
xnor U3198 (N_3198,N_2936,N_2912);
nand U3199 (N_3199,N_2725,N_2819);
and U3200 (N_3200,N_2946,N_2951);
nor U3201 (N_3201,N_2929,N_2705);
and U3202 (N_3202,N_2988,N_2701);
or U3203 (N_3203,N_2723,N_2840);
nand U3204 (N_3204,N_2885,N_2888);
nand U3205 (N_3205,N_2710,N_2921);
nor U3206 (N_3206,N_2895,N_2703);
and U3207 (N_3207,N_2906,N_2923);
nand U3208 (N_3208,N_2956,N_2939);
and U3209 (N_3209,N_2806,N_2734);
nand U3210 (N_3210,N_2895,N_2753);
or U3211 (N_3211,N_2941,N_2743);
nor U3212 (N_3212,N_2912,N_2841);
nand U3213 (N_3213,N_2945,N_2894);
or U3214 (N_3214,N_2958,N_2919);
and U3215 (N_3215,N_2831,N_2817);
or U3216 (N_3216,N_2905,N_2767);
nor U3217 (N_3217,N_2781,N_2730);
or U3218 (N_3218,N_2851,N_2743);
xnor U3219 (N_3219,N_2954,N_2874);
nand U3220 (N_3220,N_2789,N_2737);
or U3221 (N_3221,N_2943,N_2710);
and U3222 (N_3222,N_2709,N_2907);
xor U3223 (N_3223,N_2827,N_2875);
or U3224 (N_3224,N_2720,N_2848);
nor U3225 (N_3225,N_2733,N_2946);
or U3226 (N_3226,N_2766,N_2949);
nor U3227 (N_3227,N_2706,N_2852);
or U3228 (N_3228,N_2834,N_2799);
xor U3229 (N_3229,N_2888,N_2992);
and U3230 (N_3230,N_2963,N_2789);
xnor U3231 (N_3231,N_2883,N_2851);
and U3232 (N_3232,N_2994,N_2859);
and U3233 (N_3233,N_2745,N_2744);
and U3234 (N_3234,N_2870,N_2762);
or U3235 (N_3235,N_2933,N_2992);
nand U3236 (N_3236,N_2966,N_2999);
or U3237 (N_3237,N_2965,N_2710);
or U3238 (N_3238,N_2986,N_2932);
xnor U3239 (N_3239,N_2948,N_2910);
nand U3240 (N_3240,N_2772,N_2796);
xnor U3241 (N_3241,N_2739,N_2723);
or U3242 (N_3242,N_2796,N_2814);
nor U3243 (N_3243,N_2887,N_2991);
nand U3244 (N_3244,N_2833,N_2969);
nand U3245 (N_3245,N_2837,N_2813);
xnor U3246 (N_3246,N_2825,N_2968);
nand U3247 (N_3247,N_2720,N_2815);
and U3248 (N_3248,N_2747,N_2816);
and U3249 (N_3249,N_2722,N_2930);
nand U3250 (N_3250,N_2890,N_2895);
nor U3251 (N_3251,N_2732,N_2738);
and U3252 (N_3252,N_2962,N_2786);
or U3253 (N_3253,N_2906,N_2781);
nand U3254 (N_3254,N_2906,N_2722);
and U3255 (N_3255,N_2992,N_2807);
nand U3256 (N_3256,N_2889,N_2773);
nand U3257 (N_3257,N_2909,N_2850);
and U3258 (N_3258,N_2845,N_2912);
nand U3259 (N_3259,N_2987,N_2841);
xnor U3260 (N_3260,N_2999,N_2857);
or U3261 (N_3261,N_2785,N_2714);
xnor U3262 (N_3262,N_2913,N_2897);
nand U3263 (N_3263,N_2908,N_2832);
nand U3264 (N_3264,N_2965,N_2814);
nor U3265 (N_3265,N_2718,N_2738);
or U3266 (N_3266,N_2726,N_2731);
or U3267 (N_3267,N_2889,N_2969);
and U3268 (N_3268,N_2721,N_2739);
xnor U3269 (N_3269,N_2910,N_2848);
or U3270 (N_3270,N_2977,N_2739);
nand U3271 (N_3271,N_2946,N_2704);
xor U3272 (N_3272,N_2929,N_2890);
xor U3273 (N_3273,N_2726,N_2827);
xor U3274 (N_3274,N_2731,N_2780);
and U3275 (N_3275,N_2908,N_2789);
xor U3276 (N_3276,N_2949,N_2707);
and U3277 (N_3277,N_2874,N_2766);
or U3278 (N_3278,N_2967,N_2798);
or U3279 (N_3279,N_2817,N_2829);
nand U3280 (N_3280,N_2926,N_2905);
and U3281 (N_3281,N_2768,N_2944);
nor U3282 (N_3282,N_2811,N_2827);
or U3283 (N_3283,N_2822,N_2793);
nor U3284 (N_3284,N_2777,N_2776);
nand U3285 (N_3285,N_2796,N_2921);
and U3286 (N_3286,N_2964,N_2786);
and U3287 (N_3287,N_2971,N_2904);
and U3288 (N_3288,N_2949,N_2982);
and U3289 (N_3289,N_2726,N_2980);
xnor U3290 (N_3290,N_2905,N_2772);
xnor U3291 (N_3291,N_2996,N_2857);
or U3292 (N_3292,N_2889,N_2876);
and U3293 (N_3293,N_2942,N_2868);
nand U3294 (N_3294,N_2712,N_2727);
or U3295 (N_3295,N_2929,N_2855);
or U3296 (N_3296,N_2948,N_2995);
or U3297 (N_3297,N_2954,N_2708);
xnor U3298 (N_3298,N_2915,N_2944);
nor U3299 (N_3299,N_2843,N_2814);
and U3300 (N_3300,N_3058,N_3012);
and U3301 (N_3301,N_3263,N_3022);
and U3302 (N_3302,N_3063,N_3277);
or U3303 (N_3303,N_3053,N_3249);
nand U3304 (N_3304,N_3174,N_3133);
xor U3305 (N_3305,N_3076,N_3080);
nand U3306 (N_3306,N_3056,N_3254);
or U3307 (N_3307,N_3071,N_3110);
and U3308 (N_3308,N_3121,N_3048);
nand U3309 (N_3309,N_3008,N_3234);
or U3310 (N_3310,N_3128,N_3149);
nor U3311 (N_3311,N_3052,N_3019);
xor U3312 (N_3312,N_3227,N_3079);
and U3313 (N_3313,N_3215,N_3286);
xor U3314 (N_3314,N_3132,N_3119);
nor U3315 (N_3315,N_3034,N_3273);
nor U3316 (N_3316,N_3139,N_3165);
nand U3317 (N_3317,N_3123,N_3287);
nor U3318 (N_3318,N_3045,N_3153);
nand U3319 (N_3319,N_3290,N_3252);
or U3320 (N_3320,N_3070,N_3129);
and U3321 (N_3321,N_3299,N_3037);
or U3322 (N_3322,N_3011,N_3081);
and U3323 (N_3323,N_3172,N_3142);
xnor U3324 (N_3324,N_3208,N_3031);
or U3325 (N_3325,N_3274,N_3256);
nor U3326 (N_3326,N_3216,N_3219);
nor U3327 (N_3327,N_3257,N_3127);
or U3328 (N_3328,N_3072,N_3168);
nand U3329 (N_3329,N_3138,N_3026);
xor U3330 (N_3330,N_3250,N_3155);
xnor U3331 (N_3331,N_3276,N_3248);
nand U3332 (N_3332,N_3218,N_3109);
nor U3333 (N_3333,N_3162,N_3113);
or U3334 (N_3334,N_3260,N_3203);
or U3335 (N_3335,N_3220,N_3160);
xnor U3336 (N_3336,N_3095,N_3237);
nand U3337 (N_3337,N_3244,N_3038);
xor U3338 (N_3338,N_3288,N_3261);
xor U3339 (N_3339,N_3264,N_3293);
nor U3340 (N_3340,N_3083,N_3141);
nand U3341 (N_3341,N_3151,N_3057);
xnor U3342 (N_3342,N_3201,N_3193);
and U3343 (N_3343,N_3228,N_3059);
xor U3344 (N_3344,N_3096,N_3041);
nand U3345 (N_3345,N_3164,N_3236);
nand U3346 (N_3346,N_3240,N_3066);
xnor U3347 (N_3347,N_3131,N_3242);
or U3348 (N_3348,N_3186,N_3184);
xnor U3349 (N_3349,N_3295,N_3102);
nor U3350 (N_3350,N_3170,N_3262);
xor U3351 (N_3351,N_3154,N_3029);
or U3352 (N_3352,N_3221,N_3255);
and U3353 (N_3353,N_3010,N_3136);
nand U3354 (N_3354,N_3291,N_3073);
nor U3355 (N_3355,N_3021,N_3137);
nor U3356 (N_3356,N_3181,N_3185);
nand U3357 (N_3357,N_3281,N_3084);
or U3358 (N_3358,N_3177,N_3069);
nor U3359 (N_3359,N_3157,N_3148);
xor U3360 (N_3360,N_3196,N_3206);
xor U3361 (N_3361,N_3062,N_3282);
and U3362 (N_3362,N_3229,N_3098);
and U3363 (N_3363,N_3289,N_3020);
nand U3364 (N_3364,N_3259,N_3065);
nand U3365 (N_3365,N_3000,N_3145);
nand U3366 (N_3366,N_3251,N_3099);
nand U3367 (N_3367,N_3032,N_3147);
or U3368 (N_3368,N_3088,N_3014);
xor U3369 (N_3369,N_3068,N_3006);
xnor U3370 (N_3370,N_3217,N_3214);
xnor U3371 (N_3371,N_3189,N_3187);
or U3372 (N_3372,N_3064,N_3024);
nor U3373 (N_3373,N_3258,N_3016);
nand U3374 (N_3374,N_3043,N_3051);
nor U3375 (N_3375,N_3222,N_3270);
and U3376 (N_3376,N_3265,N_3115);
nand U3377 (N_3377,N_3158,N_3223);
nand U3378 (N_3378,N_3101,N_3130);
or U3379 (N_3379,N_3209,N_3232);
xor U3380 (N_3380,N_3049,N_3194);
or U3381 (N_3381,N_3086,N_3082);
nor U3382 (N_3382,N_3192,N_3001);
nor U3383 (N_3383,N_3040,N_3042);
nand U3384 (N_3384,N_3296,N_3036);
xnor U3385 (N_3385,N_3195,N_3111);
and U3386 (N_3386,N_3004,N_3005);
xnor U3387 (N_3387,N_3007,N_3247);
xor U3388 (N_3388,N_3087,N_3278);
nand U3389 (N_3389,N_3182,N_3092);
nor U3390 (N_3390,N_3023,N_3207);
xnor U3391 (N_3391,N_3226,N_3298);
nand U3392 (N_3392,N_3002,N_3173);
nand U3393 (N_3393,N_3124,N_3167);
and U3394 (N_3394,N_3078,N_3103);
nor U3395 (N_3395,N_3180,N_3114);
and U3396 (N_3396,N_3159,N_3253);
nor U3397 (N_3397,N_3134,N_3085);
xor U3398 (N_3398,N_3191,N_3241);
or U3399 (N_3399,N_3198,N_3018);
or U3400 (N_3400,N_3175,N_3108);
xnor U3401 (N_3401,N_3003,N_3171);
or U3402 (N_3402,N_3188,N_3230);
xor U3403 (N_3403,N_3179,N_3178);
and U3404 (N_3404,N_3106,N_3211);
xnor U3405 (N_3405,N_3231,N_3015);
xnor U3406 (N_3406,N_3205,N_3035);
and U3407 (N_3407,N_3202,N_3107);
nand U3408 (N_3408,N_3033,N_3284);
and U3409 (N_3409,N_3235,N_3213);
nor U3410 (N_3410,N_3143,N_3060);
and U3411 (N_3411,N_3025,N_3163);
nand U3412 (N_3412,N_3120,N_3292);
nand U3413 (N_3413,N_3161,N_3009);
nand U3414 (N_3414,N_3156,N_3285);
xnor U3415 (N_3415,N_3116,N_3212);
xnor U3416 (N_3416,N_3112,N_3061);
or U3417 (N_3417,N_3089,N_3280);
xor U3418 (N_3418,N_3269,N_3122);
nand U3419 (N_3419,N_3017,N_3077);
or U3420 (N_3420,N_3126,N_3233);
and U3421 (N_3421,N_3271,N_3239);
or U3422 (N_3422,N_3268,N_3275);
nand U3423 (N_3423,N_3166,N_3104);
and U3424 (N_3424,N_3105,N_3144);
and U3425 (N_3425,N_3075,N_3050);
or U3426 (N_3426,N_3176,N_3097);
and U3427 (N_3427,N_3210,N_3199);
nand U3428 (N_3428,N_3027,N_3272);
nor U3429 (N_3429,N_3074,N_3146);
nand U3430 (N_3430,N_3094,N_3091);
and U3431 (N_3431,N_3266,N_3044);
xnor U3432 (N_3432,N_3013,N_3090);
nand U3433 (N_3433,N_3279,N_3297);
nor U3434 (N_3434,N_3140,N_3224);
nand U3435 (N_3435,N_3225,N_3150);
nor U3436 (N_3436,N_3093,N_3100);
nor U3437 (N_3437,N_3183,N_3030);
nor U3438 (N_3438,N_3135,N_3190);
nor U3439 (N_3439,N_3238,N_3169);
nand U3440 (N_3440,N_3118,N_3055);
nand U3441 (N_3441,N_3117,N_3243);
and U3442 (N_3442,N_3294,N_3046);
nand U3443 (N_3443,N_3054,N_3028);
and U3444 (N_3444,N_3047,N_3197);
xnor U3445 (N_3445,N_3125,N_3039);
or U3446 (N_3446,N_3246,N_3204);
and U3447 (N_3447,N_3152,N_3267);
xor U3448 (N_3448,N_3283,N_3200);
nor U3449 (N_3449,N_3245,N_3067);
and U3450 (N_3450,N_3239,N_3153);
nand U3451 (N_3451,N_3252,N_3299);
nand U3452 (N_3452,N_3165,N_3222);
or U3453 (N_3453,N_3025,N_3126);
nor U3454 (N_3454,N_3003,N_3206);
or U3455 (N_3455,N_3226,N_3261);
and U3456 (N_3456,N_3164,N_3061);
nand U3457 (N_3457,N_3249,N_3158);
nand U3458 (N_3458,N_3019,N_3054);
nor U3459 (N_3459,N_3060,N_3145);
xnor U3460 (N_3460,N_3179,N_3269);
nand U3461 (N_3461,N_3169,N_3079);
or U3462 (N_3462,N_3252,N_3298);
nand U3463 (N_3463,N_3061,N_3145);
xnor U3464 (N_3464,N_3281,N_3101);
nand U3465 (N_3465,N_3252,N_3162);
and U3466 (N_3466,N_3018,N_3040);
nor U3467 (N_3467,N_3132,N_3190);
or U3468 (N_3468,N_3041,N_3085);
nor U3469 (N_3469,N_3002,N_3079);
nand U3470 (N_3470,N_3291,N_3292);
nor U3471 (N_3471,N_3020,N_3216);
xor U3472 (N_3472,N_3143,N_3037);
and U3473 (N_3473,N_3259,N_3104);
nand U3474 (N_3474,N_3040,N_3008);
and U3475 (N_3475,N_3090,N_3163);
xor U3476 (N_3476,N_3142,N_3030);
nand U3477 (N_3477,N_3153,N_3032);
nor U3478 (N_3478,N_3012,N_3230);
xnor U3479 (N_3479,N_3269,N_3125);
nor U3480 (N_3480,N_3027,N_3016);
nand U3481 (N_3481,N_3260,N_3013);
xnor U3482 (N_3482,N_3154,N_3131);
nor U3483 (N_3483,N_3154,N_3134);
nand U3484 (N_3484,N_3194,N_3067);
nand U3485 (N_3485,N_3110,N_3195);
and U3486 (N_3486,N_3200,N_3260);
nand U3487 (N_3487,N_3037,N_3226);
xnor U3488 (N_3488,N_3148,N_3037);
nand U3489 (N_3489,N_3095,N_3259);
nand U3490 (N_3490,N_3269,N_3114);
and U3491 (N_3491,N_3280,N_3088);
nor U3492 (N_3492,N_3178,N_3093);
nand U3493 (N_3493,N_3012,N_3221);
xnor U3494 (N_3494,N_3296,N_3104);
nand U3495 (N_3495,N_3151,N_3252);
nand U3496 (N_3496,N_3213,N_3089);
nand U3497 (N_3497,N_3108,N_3052);
xor U3498 (N_3498,N_3090,N_3028);
nand U3499 (N_3499,N_3141,N_3170);
xor U3500 (N_3500,N_3009,N_3292);
nand U3501 (N_3501,N_3001,N_3097);
and U3502 (N_3502,N_3129,N_3171);
and U3503 (N_3503,N_3111,N_3155);
xor U3504 (N_3504,N_3112,N_3031);
nor U3505 (N_3505,N_3268,N_3241);
nand U3506 (N_3506,N_3089,N_3032);
xor U3507 (N_3507,N_3171,N_3057);
nor U3508 (N_3508,N_3152,N_3173);
or U3509 (N_3509,N_3235,N_3140);
nor U3510 (N_3510,N_3268,N_3085);
nand U3511 (N_3511,N_3052,N_3244);
xor U3512 (N_3512,N_3021,N_3076);
and U3513 (N_3513,N_3068,N_3083);
nand U3514 (N_3514,N_3078,N_3064);
and U3515 (N_3515,N_3251,N_3071);
or U3516 (N_3516,N_3015,N_3004);
nand U3517 (N_3517,N_3130,N_3241);
and U3518 (N_3518,N_3025,N_3205);
xnor U3519 (N_3519,N_3003,N_3106);
and U3520 (N_3520,N_3131,N_3034);
or U3521 (N_3521,N_3281,N_3167);
xor U3522 (N_3522,N_3262,N_3248);
nand U3523 (N_3523,N_3152,N_3154);
nor U3524 (N_3524,N_3271,N_3269);
nand U3525 (N_3525,N_3175,N_3296);
and U3526 (N_3526,N_3199,N_3254);
nand U3527 (N_3527,N_3050,N_3180);
or U3528 (N_3528,N_3098,N_3050);
nor U3529 (N_3529,N_3067,N_3232);
nor U3530 (N_3530,N_3285,N_3163);
nand U3531 (N_3531,N_3055,N_3296);
nor U3532 (N_3532,N_3213,N_3262);
xnor U3533 (N_3533,N_3024,N_3196);
and U3534 (N_3534,N_3207,N_3066);
xor U3535 (N_3535,N_3188,N_3045);
and U3536 (N_3536,N_3288,N_3257);
xnor U3537 (N_3537,N_3008,N_3125);
or U3538 (N_3538,N_3157,N_3263);
xor U3539 (N_3539,N_3248,N_3191);
or U3540 (N_3540,N_3226,N_3101);
and U3541 (N_3541,N_3218,N_3221);
xor U3542 (N_3542,N_3261,N_3163);
nand U3543 (N_3543,N_3122,N_3231);
nor U3544 (N_3544,N_3236,N_3055);
or U3545 (N_3545,N_3029,N_3028);
and U3546 (N_3546,N_3210,N_3252);
nor U3547 (N_3547,N_3181,N_3164);
xor U3548 (N_3548,N_3106,N_3112);
xnor U3549 (N_3549,N_3143,N_3068);
nor U3550 (N_3550,N_3207,N_3193);
or U3551 (N_3551,N_3190,N_3047);
nor U3552 (N_3552,N_3288,N_3111);
nand U3553 (N_3553,N_3096,N_3198);
nor U3554 (N_3554,N_3134,N_3044);
nor U3555 (N_3555,N_3138,N_3208);
or U3556 (N_3556,N_3026,N_3049);
nand U3557 (N_3557,N_3240,N_3238);
and U3558 (N_3558,N_3213,N_3168);
xor U3559 (N_3559,N_3075,N_3018);
xor U3560 (N_3560,N_3039,N_3290);
nand U3561 (N_3561,N_3132,N_3129);
xor U3562 (N_3562,N_3223,N_3219);
nand U3563 (N_3563,N_3073,N_3225);
nand U3564 (N_3564,N_3204,N_3068);
and U3565 (N_3565,N_3004,N_3266);
xor U3566 (N_3566,N_3230,N_3203);
or U3567 (N_3567,N_3229,N_3270);
nor U3568 (N_3568,N_3079,N_3206);
or U3569 (N_3569,N_3215,N_3138);
or U3570 (N_3570,N_3042,N_3275);
nand U3571 (N_3571,N_3156,N_3297);
xnor U3572 (N_3572,N_3088,N_3210);
or U3573 (N_3573,N_3018,N_3178);
xor U3574 (N_3574,N_3002,N_3270);
xor U3575 (N_3575,N_3278,N_3027);
or U3576 (N_3576,N_3297,N_3275);
nor U3577 (N_3577,N_3094,N_3153);
nand U3578 (N_3578,N_3183,N_3034);
and U3579 (N_3579,N_3009,N_3223);
or U3580 (N_3580,N_3219,N_3294);
nor U3581 (N_3581,N_3016,N_3052);
xnor U3582 (N_3582,N_3029,N_3092);
nand U3583 (N_3583,N_3267,N_3161);
nor U3584 (N_3584,N_3090,N_3036);
and U3585 (N_3585,N_3208,N_3203);
nor U3586 (N_3586,N_3263,N_3059);
and U3587 (N_3587,N_3036,N_3194);
nand U3588 (N_3588,N_3160,N_3138);
nand U3589 (N_3589,N_3233,N_3108);
nor U3590 (N_3590,N_3100,N_3260);
or U3591 (N_3591,N_3140,N_3227);
or U3592 (N_3592,N_3019,N_3127);
xor U3593 (N_3593,N_3072,N_3032);
xor U3594 (N_3594,N_3074,N_3022);
or U3595 (N_3595,N_3005,N_3014);
nand U3596 (N_3596,N_3041,N_3210);
or U3597 (N_3597,N_3276,N_3031);
xnor U3598 (N_3598,N_3170,N_3018);
nand U3599 (N_3599,N_3089,N_3219);
nor U3600 (N_3600,N_3489,N_3410);
nand U3601 (N_3601,N_3512,N_3497);
and U3602 (N_3602,N_3426,N_3430);
nand U3603 (N_3603,N_3386,N_3448);
nand U3604 (N_3604,N_3528,N_3445);
nand U3605 (N_3605,N_3586,N_3356);
xor U3606 (N_3606,N_3532,N_3540);
or U3607 (N_3607,N_3354,N_3382);
and U3608 (N_3608,N_3312,N_3449);
xor U3609 (N_3609,N_3504,N_3453);
and U3610 (N_3610,N_3544,N_3479);
nor U3611 (N_3611,N_3552,N_3435);
nor U3612 (N_3612,N_3587,N_3391);
nand U3613 (N_3613,N_3514,N_3402);
and U3614 (N_3614,N_3520,N_3316);
and U3615 (N_3615,N_3339,N_3451);
nor U3616 (N_3616,N_3584,N_3416);
nand U3617 (N_3617,N_3490,N_3508);
nor U3618 (N_3618,N_3358,N_3425);
xor U3619 (N_3619,N_3305,N_3379);
and U3620 (N_3620,N_3447,N_3366);
nand U3621 (N_3621,N_3424,N_3422);
and U3622 (N_3622,N_3503,N_3536);
nand U3623 (N_3623,N_3380,N_3450);
or U3624 (N_3624,N_3444,N_3590);
and U3625 (N_3625,N_3436,N_3468);
xor U3626 (N_3626,N_3392,N_3313);
xnor U3627 (N_3627,N_3480,N_3319);
and U3628 (N_3628,N_3573,N_3403);
nand U3629 (N_3629,N_3433,N_3376);
or U3630 (N_3630,N_3330,N_3335);
nand U3631 (N_3631,N_3327,N_3378);
and U3632 (N_3632,N_3355,N_3415);
nor U3633 (N_3633,N_3405,N_3343);
and U3634 (N_3634,N_3539,N_3333);
nor U3635 (N_3635,N_3462,N_3341);
nor U3636 (N_3636,N_3531,N_3345);
xor U3637 (N_3637,N_3457,N_3576);
nor U3638 (N_3638,N_3585,N_3326);
or U3639 (N_3639,N_3412,N_3318);
xor U3640 (N_3640,N_3466,N_3502);
or U3641 (N_3641,N_3400,N_3334);
xnor U3642 (N_3642,N_3452,N_3567);
or U3643 (N_3643,N_3563,N_3589);
xor U3644 (N_3644,N_3568,N_3340);
or U3645 (N_3645,N_3510,N_3509);
nand U3646 (N_3646,N_3328,N_3309);
or U3647 (N_3647,N_3495,N_3560);
xor U3648 (N_3648,N_3407,N_3353);
or U3649 (N_3649,N_3564,N_3575);
nand U3650 (N_3650,N_3454,N_3347);
nand U3651 (N_3651,N_3371,N_3519);
and U3652 (N_3652,N_3579,N_3370);
nor U3653 (N_3653,N_3525,N_3530);
nand U3654 (N_3654,N_3437,N_3308);
nor U3655 (N_3655,N_3543,N_3357);
xor U3656 (N_3656,N_3420,N_3588);
or U3657 (N_3657,N_3546,N_3307);
xor U3658 (N_3658,N_3427,N_3527);
nand U3659 (N_3659,N_3484,N_3507);
nand U3660 (N_3660,N_3396,N_3558);
xor U3661 (N_3661,N_3442,N_3320);
xor U3662 (N_3662,N_3329,N_3550);
nor U3663 (N_3663,N_3488,N_3535);
or U3664 (N_3664,N_3562,N_3361);
nor U3665 (N_3665,N_3555,N_3421);
or U3666 (N_3666,N_3346,N_3470);
or U3667 (N_3667,N_3455,N_3368);
and U3668 (N_3668,N_3311,N_3557);
or U3669 (N_3669,N_3513,N_3545);
xor U3670 (N_3670,N_3350,N_3566);
or U3671 (N_3671,N_3300,N_3526);
nor U3672 (N_3672,N_3548,N_3441);
or U3673 (N_3673,N_3314,N_3310);
or U3674 (N_3674,N_3429,N_3384);
nor U3675 (N_3675,N_3477,N_3592);
nor U3676 (N_3676,N_3516,N_3362);
or U3677 (N_3677,N_3439,N_3471);
and U3678 (N_3678,N_3317,N_3411);
xor U3679 (N_3679,N_3399,N_3352);
or U3680 (N_3680,N_3547,N_3418);
xnor U3681 (N_3681,N_3324,N_3554);
nand U3682 (N_3682,N_3332,N_3537);
nor U3683 (N_3683,N_3369,N_3593);
or U3684 (N_3684,N_3580,N_3474);
xor U3685 (N_3685,N_3482,N_3349);
or U3686 (N_3686,N_3306,N_3483);
nand U3687 (N_3687,N_3359,N_3570);
nor U3688 (N_3688,N_3553,N_3414);
nand U3689 (N_3689,N_3496,N_3473);
xor U3690 (N_3690,N_3409,N_3398);
xor U3691 (N_3691,N_3365,N_3459);
or U3692 (N_3692,N_3408,N_3385);
or U3693 (N_3693,N_3523,N_3542);
xnor U3694 (N_3694,N_3596,N_3476);
xnor U3695 (N_3695,N_3322,N_3494);
nor U3696 (N_3696,N_3446,N_3595);
or U3697 (N_3697,N_3577,N_3458);
or U3698 (N_3698,N_3381,N_3338);
and U3699 (N_3699,N_3401,N_3406);
xor U3700 (N_3700,N_3481,N_3337);
nor U3701 (N_3701,N_3561,N_3331);
nor U3702 (N_3702,N_3524,N_3517);
xor U3703 (N_3703,N_3377,N_3397);
or U3704 (N_3704,N_3487,N_3501);
xnor U3705 (N_3705,N_3388,N_3423);
nand U3706 (N_3706,N_3443,N_3475);
xnor U3707 (N_3707,N_3578,N_3598);
or U3708 (N_3708,N_3434,N_3521);
xnor U3709 (N_3709,N_3417,N_3302);
and U3710 (N_3710,N_3522,N_3478);
and U3711 (N_3711,N_3594,N_3304);
nor U3712 (N_3712,N_3342,N_3461);
nor U3713 (N_3713,N_3472,N_3493);
nand U3714 (N_3714,N_3534,N_3364);
and U3715 (N_3715,N_3556,N_3498);
xor U3716 (N_3716,N_3404,N_3387);
or U3717 (N_3717,N_3432,N_3559);
or U3718 (N_3718,N_3395,N_3372);
and U3719 (N_3719,N_3515,N_3551);
and U3720 (N_3720,N_3348,N_3393);
nor U3721 (N_3721,N_3597,N_3374);
nor U3722 (N_3722,N_3389,N_3569);
and U3723 (N_3723,N_3465,N_3344);
xor U3724 (N_3724,N_3323,N_3565);
or U3725 (N_3725,N_3583,N_3486);
xor U3726 (N_3726,N_3367,N_3336);
xnor U3727 (N_3727,N_3485,N_3591);
and U3728 (N_3728,N_3456,N_3581);
and U3729 (N_3729,N_3383,N_3571);
and U3730 (N_3730,N_3351,N_3463);
nand U3731 (N_3731,N_3491,N_3375);
nand U3732 (N_3732,N_3360,N_3469);
or U3733 (N_3733,N_3505,N_3428);
xnor U3734 (N_3734,N_3572,N_3460);
nand U3735 (N_3735,N_3549,N_3541);
or U3736 (N_3736,N_3506,N_3438);
xnor U3737 (N_3737,N_3325,N_3301);
or U3738 (N_3738,N_3529,N_3464);
and U3739 (N_3739,N_3533,N_3499);
or U3740 (N_3740,N_3413,N_3500);
or U3741 (N_3741,N_3582,N_3431);
xor U3742 (N_3742,N_3390,N_3538);
and U3743 (N_3743,N_3511,N_3440);
or U3744 (N_3744,N_3467,N_3599);
nor U3745 (N_3745,N_3303,N_3394);
and U3746 (N_3746,N_3518,N_3419);
nand U3747 (N_3747,N_3363,N_3321);
xnor U3748 (N_3748,N_3574,N_3315);
and U3749 (N_3749,N_3373,N_3492);
nand U3750 (N_3750,N_3471,N_3575);
or U3751 (N_3751,N_3544,N_3367);
nor U3752 (N_3752,N_3341,N_3514);
xnor U3753 (N_3753,N_3578,N_3400);
and U3754 (N_3754,N_3345,N_3482);
or U3755 (N_3755,N_3458,N_3473);
xnor U3756 (N_3756,N_3532,N_3397);
nor U3757 (N_3757,N_3435,N_3452);
nor U3758 (N_3758,N_3494,N_3345);
nand U3759 (N_3759,N_3362,N_3450);
nor U3760 (N_3760,N_3546,N_3574);
nor U3761 (N_3761,N_3599,N_3364);
and U3762 (N_3762,N_3339,N_3380);
nor U3763 (N_3763,N_3416,N_3373);
nand U3764 (N_3764,N_3492,N_3569);
nand U3765 (N_3765,N_3549,N_3446);
or U3766 (N_3766,N_3377,N_3518);
and U3767 (N_3767,N_3329,N_3545);
or U3768 (N_3768,N_3446,N_3368);
xor U3769 (N_3769,N_3499,N_3310);
nand U3770 (N_3770,N_3349,N_3405);
or U3771 (N_3771,N_3382,N_3375);
xnor U3772 (N_3772,N_3349,N_3436);
or U3773 (N_3773,N_3570,N_3599);
nand U3774 (N_3774,N_3456,N_3431);
nor U3775 (N_3775,N_3340,N_3320);
nand U3776 (N_3776,N_3379,N_3430);
or U3777 (N_3777,N_3531,N_3322);
or U3778 (N_3778,N_3538,N_3515);
or U3779 (N_3779,N_3434,N_3459);
xor U3780 (N_3780,N_3502,N_3507);
or U3781 (N_3781,N_3548,N_3310);
nand U3782 (N_3782,N_3567,N_3590);
nand U3783 (N_3783,N_3534,N_3573);
and U3784 (N_3784,N_3409,N_3338);
xnor U3785 (N_3785,N_3546,N_3389);
nand U3786 (N_3786,N_3589,N_3413);
or U3787 (N_3787,N_3457,N_3306);
nand U3788 (N_3788,N_3325,N_3523);
or U3789 (N_3789,N_3591,N_3598);
xnor U3790 (N_3790,N_3425,N_3581);
xor U3791 (N_3791,N_3384,N_3577);
xor U3792 (N_3792,N_3493,N_3323);
or U3793 (N_3793,N_3403,N_3368);
nor U3794 (N_3794,N_3474,N_3436);
nand U3795 (N_3795,N_3397,N_3481);
and U3796 (N_3796,N_3373,N_3409);
nor U3797 (N_3797,N_3511,N_3366);
and U3798 (N_3798,N_3327,N_3461);
xnor U3799 (N_3799,N_3301,N_3346);
nor U3800 (N_3800,N_3465,N_3423);
and U3801 (N_3801,N_3374,N_3313);
and U3802 (N_3802,N_3315,N_3525);
nor U3803 (N_3803,N_3482,N_3581);
xor U3804 (N_3804,N_3569,N_3452);
or U3805 (N_3805,N_3575,N_3328);
nand U3806 (N_3806,N_3317,N_3417);
and U3807 (N_3807,N_3591,N_3456);
nand U3808 (N_3808,N_3553,N_3516);
nor U3809 (N_3809,N_3356,N_3463);
nor U3810 (N_3810,N_3469,N_3355);
or U3811 (N_3811,N_3493,N_3585);
nor U3812 (N_3812,N_3433,N_3536);
xor U3813 (N_3813,N_3361,N_3438);
and U3814 (N_3814,N_3445,N_3541);
nor U3815 (N_3815,N_3452,N_3346);
xor U3816 (N_3816,N_3356,N_3440);
nand U3817 (N_3817,N_3363,N_3498);
or U3818 (N_3818,N_3543,N_3319);
nor U3819 (N_3819,N_3369,N_3495);
nor U3820 (N_3820,N_3392,N_3596);
xor U3821 (N_3821,N_3565,N_3309);
nor U3822 (N_3822,N_3369,N_3371);
xnor U3823 (N_3823,N_3344,N_3486);
xnor U3824 (N_3824,N_3441,N_3309);
and U3825 (N_3825,N_3521,N_3507);
nor U3826 (N_3826,N_3552,N_3534);
xor U3827 (N_3827,N_3395,N_3306);
nor U3828 (N_3828,N_3548,N_3379);
or U3829 (N_3829,N_3402,N_3544);
and U3830 (N_3830,N_3512,N_3554);
or U3831 (N_3831,N_3595,N_3487);
or U3832 (N_3832,N_3531,N_3596);
or U3833 (N_3833,N_3415,N_3335);
nand U3834 (N_3834,N_3337,N_3393);
nor U3835 (N_3835,N_3437,N_3363);
or U3836 (N_3836,N_3490,N_3465);
nor U3837 (N_3837,N_3549,N_3537);
nor U3838 (N_3838,N_3485,N_3499);
xor U3839 (N_3839,N_3322,N_3456);
or U3840 (N_3840,N_3339,N_3555);
nand U3841 (N_3841,N_3487,N_3433);
and U3842 (N_3842,N_3491,N_3328);
nand U3843 (N_3843,N_3505,N_3384);
nor U3844 (N_3844,N_3493,N_3581);
nor U3845 (N_3845,N_3303,N_3308);
xnor U3846 (N_3846,N_3389,N_3402);
and U3847 (N_3847,N_3506,N_3441);
and U3848 (N_3848,N_3470,N_3527);
xnor U3849 (N_3849,N_3429,N_3582);
and U3850 (N_3850,N_3333,N_3369);
nand U3851 (N_3851,N_3490,N_3364);
nor U3852 (N_3852,N_3478,N_3548);
or U3853 (N_3853,N_3304,N_3321);
and U3854 (N_3854,N_3400,N_3445);
nor U3855 (N_3855,N_3390,N_3417);
nand U3856 (N_3856,N_3440,N_3549);
and U3857 (N_3857,N_3353,N_3563);
xnor U3858 (N_3858,N_3415,N_3411);
xnor U3859 (N_3859,N_3599,N_3323);
or U3860 (N_3860,N_3334,N_3580);
and U3861 (N_3861,N_3372,N_3466);
nor U3862 (N_3862,N_3597,N_3506);
nor U3863 (N_3863,N_3569,N_3368);
or U3864 (N_3864,N_3337,N_3380);
nor U3865 (N_3865,N_3574,N_3485);
nor U3866 (N_3866,N_3541,N_3467);
and U3867 (N_3867,N_3532,N_3584);
nor U3868 (N_3868,N_3335,N_3580);
nor U3869 (N_3869,N_3554,N_3413);
and U3870 (N_3870,N_3350,N_3545);
nand U3871 (N_3871,N_3331,N_3537);
nand U3872 (N_3872,N_3337,N_3356);
xnor U3873 (N_3873,N_3596,N_3372);
xnor U3874 (N_3874,N_3422,N_3419);
or U3875 (N_3875,N_3475,N_3477);
nor U3876 (N_3876,N_3500,N_3544);
nor U3877 (N_3877,N_3578,N_3397);
xnor U3878 (N_3878,N_3326,N_3344);
nand U3879 (N_3879,N_3341,N_3384);
and U3880 (N_3880,N_3363,N_3540);
nand U3881 (N_3881,N_3501,N_3510);
and U3882 (N_3882,N_3556,N_3421);
or U3883 (N_3883,N_3465,N_3381);
nor U3884 (N_3884,N_3404,N_3353);
or U3885 (N_3885,N_3539,N_3331);
nor U3886 (N_3886,N_3490,N_3507);
or U3887 (N_3887,N_3491,N_3381);
or U3888 (N_3888,N_3439,N_3432);
nand U3889 (N_3889,N_3549,N_3309);
xor U3890 (N_3890,N_3581,N_3479);
xnor U3891 (N_3891,N_3531,N_3335);
nor U3892 (N_3892,N_3478,N_3346);
or U3893 (N_3893,N_3476,N_3431);
or U3894 (N_3894,N_3353,N_3509);
nand U3895 (N_3895,N_3421,N_3368);
or U3896 (N_3896,N_3472,N_3351);
xor U3897 (N_3897,N_3310,N_3492);
or U3898 (N_3898,N_3445,N_3329);
xnor U3899 (N_3899,N_3485,N_3345);
xnor U3900 (N_3900,N_3603,N_3774);
nand U3901 (N_3901,N_3627,N_3717);
nand U3902 (N_3902,N_3823,N_3758);
or U3903 (N_3903,N_3607,N_3664);
nor U3904 (N_3904,N_3643,N_3771);
and U3905 (N_3905,N_3613,N_3742);
nor U3906 (N_3906,N_3851,N_3852);
nand U3907 (N_3907,N_3676,N_3814);
nand U3908 (N_3908,N_3876,N_3672);
nand U3909 (N_3909,N_3844,N_3684);
and U3910 (N_3910,N_3864,N_3646);
nor U3911 (N_3911,N_3601,N_3700);
nand U3912 (N_3912,N_3780,N_3884);
nor U3913 (N_3913,N_3856,N_3683);
nand U3914 (N_3914,N_3785,N_3783);
nor U3915 (N_3915,N_3846,N_3795);
nand U3916 (N_3916,N_3677,N_3657);
nor U3917 (N_3917,N_3714,N_3870);
and U3918 (N_3918,N_3654,N_3631);
nand U3919 (N_3919,N_3837,N_3895);
and U3920 (N_3920,N_3635,N_3816);
xnor U3921 (N_3921,N_3609,N_3796);
and U3922 (N_3922,N_3826,N_3896);
nor U3923 (N_3923,N_3834,N_3756);
nor U3924 (N_3924,N_3655,N_3629);
nor U3925 (N_3925,N_3786,N_3812);
or U3926 (N_3926,N_3740,N_3600);
and U3927 (N_3927,N_3839,N_3855);
or U3928 (N_3928,N_3820,N_3859);
xnor U3929 (N_3929,N_3619,N_3882);
and U3930 (N_3930,N_3865,N_3668);
and U3931 (N_3931,N_3718,N_3822);
nand U3932 (N_3932,N_3848,N_3788);
or U3933 (N_3933,N_3784,N_3872);
xnor U3934 (N_3934,N_3695,N_3735);
xnor U3935 (N_3935,N_3703,N_3707);
nand U3936 (N_3936,N_3874,N_3623);
xor U3937 (N_3937,N_3806,N_3674);
or U3938 (N_3938,N_3636,N_3720);
and U3939 (N_3939,N_3817,N_3687);
and U3940 (N_3940,N_3776,N_3725);
nor U3941 (N_3941,N_3811,N_3724);
or U3942 (N_3942,N_3889,N_3626);
or U3943 (N_3943,N_3782,N_3797);
nor U3944 (N_3944,N_3857,N_3604);
nor U3945 (N_3945,N_3807,N_3800);
or U3946 (N_3946,N_3747,N_3828);
and U3947 (N_3947,N_3705,N_3688);
or U3948 (N_3948,N_3749,N_3815);
xor U3949 (N_3949,N_3781,N_3610);
or U3950 (N_3950,N_3810,N_3673);
and U3951 (N_3951,N_3743,N_3727);
nand U3952 (N_3952,N_3899,N_3692);
or U3953 (N_3953,N_3755,N_3893);
or U3954 (N_3954,N_3888,N_3632);
nor U3955 (N_3955,N_3726,N_3850);
xor U3956 (N_3956,N_3843,N_3671);
or U3957 (N_3957,N_3818,N_3711);
or U3958 (N_3958,N_3713,N_3620);
or U3959 (N_3959,N_3892,N_3836);
nor U3960 (N_3960,N_3854,N_3708);
and U3961 (N_3961,N_3805,N_3652);
and U3962 (N_3962,N_3624,N_3831);
nand U3963 (N_3963,N_3666,N_3878);
nand U3964 (N_3964,N_3883,N_3678);
nor U3965 (N_3965,N_3642,N_3875);
or U3966 (N_3966,N_3691,N_3842);
or U3967 (N_3967,N_3648,N_3869);
nor U3968 (N_3968,N_3791,N_3661);
and U3969 (N_3969,N_3794,N_3719);
and U3970 (N_3970,N_3890,N_3697);
xor U3971 (N_3971,N_3798,N_3879);
xnor U3972 (N_3972,N_3651,N_3802);
nor U3973 (N_3973,N_3829,N_3722);
nor U3974 (N_3974,N_3667,N_3845);
nor U3975 (N_3975,N_3790,N_3633);
nand U3976 (N_3976,N_3838,N_3832);
nand U3977 (N_3977,N_3803,N_3693);
or U3978 (N_3978,N_3679,N_3793);
or U3979 (N_3979,N_3721,N_3871);
nand U3980 (N_3980,N_3602,N_3751);
nor U3981 (N_3981,N_3701,N_3649);
nor U3982 (N_3982,N_3690,N_3630);
nand U3983 (N_3983,N_3741,N_3698);
xor U3984 (N_3984,N_3757,N_3885);
or U3985 (N_3985,N_3809,N_3663);
nor U3986 (N_3986,N_3863,N_3853);
nor U3987 (N_3987,N_3611,N_3825);
or U3988 (N_3988,N_3760,N_3873);
and U3989 (N_3989,N_3827,N_3670);
or U3990 (N_3990,N_3731,N_3801);
or U3991 (N_3991,N_3625,N_3841);
and U3992 (N_3992,N_3894,N_3660);
nor U3993 (N_3993,N_3681,N_3608);
or U3994 (N_3994,N_3858,N_3778);
and U3995 (N_3995,N_3868,N_3614);
xor U3996 (N_3996,N_3765,N_3659);
nand U3997 (N_3997,N_3728,N_3867);
nor U3998 (N_3998,N_3764,N_3847);
xor U3999 (N_3999,N_3641,N_3634);
and U4000 (N_4000,N_3898,N_3622);
and U4001 (N_4001,N_3824,N_3637);
xor U4002 (N_4002,N_3881,N_3887);
nand U4003 (N_4003,N_3761,N_3804);
xor U4004 (N_4004,N_3787,N_3732);
nor U4005 (N_4005,N_3833,N_3821);
xnor U4006 (N_4006,N_3897,N_3799);
nand U4007 (N_4007,N_3699,N_3754);
nand U4008 (N_4008,N_3662,N_3792);
nor U4009 (N_4009,N_3706,N_3712);
and U4010 (N_4010,N_3696,N_3777);
and U4011 (N_4011,N_3759,N_3617);
nand U4012 (N_4012,N_3762,N_3769);
or U4013 (N_4013,N_3730,N_3766);
xnor U4014 (N_4014,N_3763,N_3746);
nor U4015 (N_4015,N_3849,N_3789);
nor U4016 (N_4016,N_3737,N_3606);
xor U4017 (N_4017,N_3775,N_3639);
xnor U4018 (N_4018,N_3891,N_3709);
and U4019 (N_4019,N_3733,N_3860);
or U4020 (N_4020,N_3835,N_3689);
and U4021 (N_4021,N_3715,N_3638);
xnor U4022 (N_4022,N_3750,N_3748);
nor U4023 (N_4023,N_3615,N_3734);
nor U4024 (N_4024,N_3745,N_3644);
xor U4025 (N_4025,N_3808,N_3612);
nor U4026 (N_4026,N_3779,N_3770);
nor U4027 (N_4027,N_3621,N_3658);
and U4028 (N_4028,N_3767,N_3704);
nand U4029 (N_4029,N_3773,N_3886);
nand U4030 (N_4030,N_3669,N_3605);
nor U4031 (N_4031,N_3686,N_3616);
nor U4032 (N_4032,N_3645,N_3753);
and U4033 (N_4033,N_3682,N_3656);
nor U4034 (N_4034,N_3650,N_3819);
or U4035 (N_4035,N_3861,N_3675);
and U4036 (N_4036,N_3665,N_3877);
and U4037 (N_4037,N_3866,N_3653);
nand U4038 (N_4038,N_3710,N_3729);
nand U4039 (N_4039,N_3813,N_3772);
or U4040 (N_4040,N_3744,N_3694);
nand U4041 (N_4041,N_3840,N_3640);
and U4042 (N_4042,N_3628,N_3736);
nor U4043 (N_4043,N_3723,N_3702);
and U4044 (N_4044,N_3862,N_3685);
nor U4045 (N_4045,N_3768,N_3647);
nor U4046 (N_4046,N_3738,N_3880);
xnor U4047 (N_4047,N_3618,N_3752);
or U4048 (N_4048,N_3830,N_3680);
and U4049 (N_4049,N_3716,N_3739);
nor U4050 (N_4050,N_3746,N_3699);
xnor U4051 (N_4051,N_3753,N_3860);
and U4052 (N_4052,N_3899,N_3827);
nor U4053 (N_4053,N_3829,N_3751);
xnor U4054 (N_4054,N_3705,N_3883);
nand U4055 (N_4055,N_3658,N_3688);
nand U4056 (N_4056,N_3880,N_3792);
nor U4057 (N_4057,N_3616,N_3830);
xor U4058 (N_4058,N_3631,N_3776);
xnor U4059 (N_4059,N_3760,N_3798);
and U4060 (N_4060,N_3726,N_3875);
or U4061 (N_4061,N_3704,N_3853);
or U4062 (N_4062,N_3806,N_3664);
nor U4063 (N_4063,N_3605,N_3898);
nor U4064 (N_4064,N_3761,N_3742);
nand U4065 (N_4065,N_3755,N_3677);
xor U4066 (N_4066,N_3701,N_3622);
and U4067 (N_4067,N_3704,N_3820);
or U4068 (N_4068,N_3886,N_3672);
xor U4069 (N_4069,N_3790,N_3613);
and U4070 (N_4070,N_3825,N_3724);
xnor U4071 (N_4071,N_3662,N_3741);
xor U4072 (N_4072,N_3899,N_3704);
xor U4073 (N_4073,N_3827,N_3722);
nor U4074 (N_4074,N_3859,N_3741);
xnor U4075 (N_4075,N_3778,N_3674);
xor U4076 (N_4076,N_3764,N_3850);
and U4077 (N_4077,N_3633,N_3772);
nor U4078 (N_4078,N_3665,N_3879);
or U4079 (N_4079,N_3642,N_3848);
and U4080 (N_4080,N_3839,N_3633);
nand U4081 (N_4081,N_3845,N_3814);
or U4082 (N_4082,N_3678,N_3671);
nor U4083 (N_4083,N_3760,N_3672);
nand U4084 (N_4084,N_3824,N_3773);
or U4085 (N_4085,N_3827,N_3751);
xnor U4086 (N_4086,N_3686,N_3843);
xnor U4087 (N_4087,N_3823,N_3673);
nor U4088 (N_4088,N_3718,N_3653);
or U4089 (N_4089,N_3803,N_3721);
or U4090 (N_4090,N_3897,N_3703);
nand U4091 (N_4091,N_3787,N_3714);
nor U4092 (N_4092,N_3880,N_3704);
xnor U4093 (N_4093,N_3803,N_3643);
xor U4094 (N_4094,N_3853,N_3750);
and U4095 (N_4095,N_3819,N_3823);
and U4096 (N_4096,N_3740,N_3699);
or U4097 (N_4097,N_3726,N_3858);
nor U4098 (N_4098,N_3853,N_3673);
nor U4099 (N_4099,N_3787,N_3899);
and U4100 (N_4100,N_3792,N_3611);
or U4101 (N_4101,N_3846,N_3630);
and U4102 (N_4102,N_3891,N_3855);
nand U4103 (N_4103,N_3808,N_3695);
nand U4104 (N_4104,N_3759,N_3632);
or U4105 (N_4105,N_3820,N_3769);
and U4106 (N_4106,N_3694,N_3872);
nand U4107 (N_4107,N_3767,N_3831);
or U4108 (N_4108,N_3867,N_3767);
or U4109 (N_4109,N_3796,N_3789);
nor U4110 (N_4110,N_3710,N_3683);
nor U4111 (N_4111,N_3825,N_3717);
xor U4112 (N_4112,N_3602,N_3797);
xor U4113 (N_4113,N_3893,N_3873);
nor U4114 (N_4114,N_3879,N_3866);
or U4115 (N_4115,N_3795,N_3811);
xor U4116 (N_4116,N_3873,N_3663);
xor U4117 (N_4117,N_3605,N_3855);
nand U4118 (N_4118,N_3604,N_3763);
nor U4119 (N_4119,N_3659,N_3603);
and U4120 (N_4120,N_3738,N_3646);
xor U4121 (N_4121,N_3663,N_3847);
nand U4122 (N_4122,N_3721,N_3638);
nor U4123 (N_4123,N_3872,N_3647);
nand U4124 (N_4124,N_3663,N_3730);
xnor U4125 (N_4125,N_3834,N_3693);
xor U4126 (N_4126,N_3690,N_3706);
or U4127 (N_4127,N_3609,N_3771);
xnor U4128 (N_4128,N_3794,N_3843);
nand U4129 (N_4129,N_3737,N_3608);
xor U4130 (N_4130,N_3764,N_3738);
and U4131 (N_4131,N_3837,N_3738);
xnor U4132 (N_4132,N_3812,N_3750);
xnor U4133 (N_4133,N_3743,N_3785);
and U4134 (N_4134,N_3629,N_3823);
or U4135 (N_4135,N_3898,N_3834);
and U4136 (N_4136,N_3896,N_3627);
nor U4137 (N_4137,N_3700,N_3777);
xor U4138 (N_4138,N_3844,N_3852);
and U4139 (N_4139,N_3869,N_3831);
nand U4140 (N_4140,N_3781,N_3850);
or U4141 (N_4141,N_3726,N_3634);
xnor U4142 (N_4142,N_3860,N_3608);
nor U4143 (N_4143,N_3887,N_3625);
and U4144 (N_4144,N_3784,N_3718);
nor U4145 (N_4145,N_3830,N_3729);
and U4146 (N_4146,N_3648,N_3724);
and U4147 (N_4147,N_3600,N_3627);
or U4148 (N_4148,N_3651,N_3730);
nand U4149 (N_4149,N_3818,N_3687);
nor U4150 (N_4150,N_3830,N_3856);
or U4151 (N_4151,N_3761,N_3640);
and U4152 (N_4152,N_3640,N_3843);
xor U4153 (N_4153,N_3874,N_3601);
nand U4154 (N_4154,N_3615,N_3602);
or U4155 (N_4155,N_3852,N_3673);
xnor U4156 (N_4156,N_3633,N_3720);
xor U4157 (N_4157,N_3803,N_3685);
nand U4158 (N_4158,N_3868,N_3734);
and U4159 (N_4159,N_3670,N_3736);
nand U4160 (N_4160,N_3664,N_3663);
nand U4161 (N_4161,N_3769,N_3825);
and U4162 (N_4162,N_3619,N_3638);
nand U4163 (N_4163,N_3721,N_3815);
nand U4164 (N_4164,N_3666,N_3668);
nor U4165 (N_4165,N_3837,N_3658);
and U4166 (N_4166,N_3836,N_3806);
nor U4167 (N_4167,N_3607,N_3662);
and U4168 (N_4168,N_3646,N_3797);
nand U4169 (N_4169,N_3686,N_3878);
nor U4170 (N_4170,N_3670,N_3739);
nand U4171 (N_4171,N_3660,N_3734);
and U4172 (N_4172,N_3797,N_3747);
nor U4173 (N_4173,N_3697,N_3785);
xnor U4174 (N_4174,N_3880,N_3873);
xor U4175 (N_4175,N_3746,N_3712);
xnor U4176 (N_4176,N_3891,N_3848);
nand U4177 (N_4177,N_3811,N_3740);
and U4178 (N_4178,N_3782,N_3719);
and U4179 (N_4179,N_3737,N_3805);
xor U4180 (N_4180,N_3697,N_3876);
or U4181 (N_4181,N_3691,N_3720);
nor U4182 (N_4182,N_3663,N_3811);
and U4183 (N_4183,N_3860,N_3633);
nor U4184 (N_4184,N_3817,N_3666);
and U4185 (N_4185,N_3830,N_3621);
or U4186 (N_4186,N_3732,N_3737);
nand U4187 (N_4187,N_3821,N_3738);
xor U4188 (N_4188,N_3868,N_3798);
and U4189 (N_4189,N_3851,N_3876);
nand U4190 (N_4190,N_3799,N_3606);
nor U4191 (N_4191,N_3835,N_3809);
or U4192 (N_4192,N_3700,N_3751);
or U4193 (N_4193,N_3603,N_3805);
and U4194 (N_4194,N_3743,N_3608);
and U4195 (N_4195,N_3754,N_3711);
xor U4196 (N_4196,N_3866,N_3637);
or U4197 (N_4197,N_3798,N_3809);
nor U4198 (N_4198,N_3606,N_3816);
nor U4199 (N_4199,N_3715,N_3892);
nand U4200 (N_4200,N_4017,N_3982);
xnor U4201 (N_4201,N_3999,N_4132);
xor U4202 (N_4202,N_3932,N_3983);
nand U4203 (N_4203,N_4001,N_3970);
nor U4204 (N_4204,N_4092,N_4197);
or U4205 (N_4205,N_4008,N_3952);
xor U4206 (N_4206,N_4100,N_4124);
xnor U4207 (N_4207,N_4038,N_3926);
or U4208 (N_4208,N_4007,N_4010);
nand U4209 (N_4209,N_4168,N_4190);
nor U4210 (N_4210,N_4182,N_4166);
nand U4211 (N_4211,N_4187,N_4108);
nand U4212 (N_4212,N_4073,N_4120);
nand U4213 (N_4213,N_4026,N_4083);
xor U4214 (N_4214,N_4137,N_4150);
xnor U4215 (N_4215,N_4025,N_3940);
nand U4216 (N_4216,N_4184,N_3941);
or U4217 (N_4217,N_3908,N_4159);
and U4218 (N_4218,N_4056,N_4012);
xor U4219 (N_4219,N_4097,N_4078);
nor U4220 (N_4220,N_4054,N_4169);
xor U4221 (N_4221,N_3912,N_4185);
and U4222 (N_4222,N_4070,N_4086);
xnor U4223 (N_4223,N_4065,N_4109);
xor U4224 (N_4224,N_4134,N_3984);
nand U4225 (N_4225,N_3921,N_4121);
and U4226 (N_4226,N_3980,N_3947);
nand U4227 (N_4227,N_4045,N_4105);
xor U4228 (N_4228,N_3909,N_3988);
and U4229 (N_4229,N_4091,N_4144);
xnor U4230 (N_4230,N_3922,N_3954);
nand U4231 (N_4231,N_3938,N_4037);
xnor U4232 (N_4232,N_3950,N_3996);
xnor U4233 (N_4233,N_3987,N_4060);
xnor U4234 (N_4234,N_4021,N_3939);
nand U4235 (N_4235,N_3913,N_3963);
nand U4236 (N_4236,N_4119,N_3998);
xor U4237 (N_4237,N_4112,N_3967);
nor U4238 (N_4238,N_4002,N_4127);
or U4239 (N_4239,N_4059,N_4082);
nor U4240 (N_4240,N_4011,N_4041);
xor U4241 (N_4241,N_4103,N_3903);
xnor U4242 (N_4242,N_4055,N_4087);
or U4243 (N_4243,N_3937,N_4033);
or U4244 (N_4244,N_4135,N_3958);
nand U4245 (N_4245,N_4032,N_4035);
and U4246 (N_4246,N_4048,N_4043);
nor U4247 (N_4247,N_4183,N_4063);
nor U4248 (N_4248,N_4018,N_4198);
or U4249 (N_4249,N_4110,N_4057);
nand U4250 (N_4250,N_3977,N_4094);
or U4251 (N_4251,N_4141,N_4172);
nor U4252 (N_4252,N_3934,N_4160);
xor U4253 (N_4253,N_4020,N_3972);
or U4254 (N_4254,N_3964,N_4062);
nand U4255 (N_4255,N_4188,N_3966);
and U4256 (N_4256,N_4171,N_3927);
nor U4257 (N_4257,N_4193,N_4195);
xnor U4258 (N_4258,N_4095,N_3925);
nand U4259 (N_4259,N_4085,N_3946);
or U4260 (N_4260,N_4024,N_4016);
nor U4261 (N_4261,N_4003,N_4104);
nand U4262 (N_4262,N_3956,N_4199);
and U4263 (N_4263,N_3914,N_3917);
nor U4264 (N_4264,N_3920,N_4069);
xor U4265 (N_4265,N_3994,N_4036);
nor U4266 (N_4266,N_4167,N_4028);
xor U4267 (N_4267,N_4143,N_4170);
or U4268 (N_4268,N_4155,N_4034);
nand U4269 (N_4269,N_3981,N_4081);
nor U4270 (N_4270,N_3955,N_4089);
or U4271 (N_4271,N_3900,N_4061);
xnor U4272 (N_4272,N_3992,N_3989);
nand U4273 (N_4273,N_4080,N_4163);
nor U4274 (N_4274,N_4051,N_3904);
and U4275 (N_4275,N_4115,N_3997);
or U4276 (N_4276,N_3974,N_3957);
or U4277 (N_4277,N_4006,N_3951);
xnor U4278 (N_4278,N_4164,N_4174);
or U4279 (N_4279,N_4023,N_3915);
nor U4280 (N_4280,N_4077,N_3906);
nor U4281 (N_4281,N_3942,N_4158);
nand U4282 (N_4282,N_4153,N_3953);
and U4283 (N_4283,N_4125,N_4042);
nor U4284 (N_4284,N_4040,N_4180);
or U4285 (N_4285,N_4096,N_3901);
xor U4286 (N_4286,N_4098,N_4177);
nor U4287 (N_4287,N_4031,N_4173);
nand U4288 (N_4288,N_4196,N_4156);
or U4289 (N_4289,N_4162,N_4102);
nand U4290 (N_4290,N_3928,N_3918);
or U4291 (N_4291,N_3979,N_4161);
or U4292 (N_4292,N_3911,N_4149);
or U4293 (N_4293,N_4058,N_3936);
or U4294 (N_4294,N_4013,N_4129);
or U4295 (N_4295,N_4139,N_3948);
nor U4296 (N_4296,N_4079,N_3965);
and U4297 (N_4297,N_3905,N_4122);
or U4298 (N_4298,N_4123,N_4067);
or U4299 (N_4299,N_4192,N_4131);
nand U4300 (N_4300,N_4189,N_3930);
or U4301 (N_4301,N_4157,N_3986);
and U4302 (N_4302,N_4165,N_3991);
and U4303 (N_4303,N_3993,N_3907);
and U4304 (N_4304,N_4075,N_4106);
nor U4305 (N_4305,N_3978,N_4076);
nand U4306 (N_4306,N_4117,N_4014);
or U4307 (N_4307,N_4148,N_4005);
and U4308 (N_4308,N_4029,N_4186);
xor U4309 (N_4309,N_4052,N_4090);
xnor U4310 (N_4310,N_3962,N_4039);
and U4311 (N_4311,N_3990,N_3975);
or U4312 (N_4312,N_4049,N_4111);
or U4313 (N_4313,N_4066,N_4145);
and U4314 (N_4314,N_3973,N_4088);
nand U4315 (N_4315,N_3919,N_3971);
xor U4316 (N_4316,N_3945,N_4147);
nand U4317 (N_4317,N_3943,N_4064);
nor U4318 (N_4318,N_4114,N_4019);
or U4319 (N_4319,N_4071,N_4000);
or U4320 (N_4320,N_4101,N_4138);
xor U4321 (N_4321,N_4128,N_4027);
or U4322 (N_4322,N_4084,N_4176);
nand U4323 (N_4323,N_3910,N_3929);
or U4324 (N_4324,N_4130,N_4194);
xnor U4325 (N_4325,N_4178,N_4126);
xor U4326 (N_4326,N_4009,N_4181);
nand U4327 (N_4327,N_3959,N_3968);
nor U4328 (N_4328,N_4099,N_3924);
xor U4329 (N_4329,N_4146,N_4074);
nor U4330 (N_4330,N_4053,N_4022);
nand U4331 (N_4331,N_4116,N_3960);
nor U4332 (N_4332,N_4142,N_3923);
or U4333 (N_4333,N_4047,N_4004);
xnor U4334 (N_4334,N_3916,N_3985);
nor U4335 (N_4335,N_4179,N_3961);
nand U4336 (N_4336,N_4152,N_4044);
xor U4337 (N_4337,N_3944,N_3931);
and U4338 (N_4338,N_3949,N_3935);
nand U4339 (N_4339,N_4136,N_4118);
or U4340 (N_4340,N_4133,N_4151);
nand U4341 (N_4341,N_4113,N_4046);
xor U4342 (N_4342,N_4107,N_4072);
or U4343 (N_4343,N_4050,N_4093);
nand U4344 (N_4344,N_3933,N_4175);
and U4345 (N_4345,N_4030,N_4068);
nand U4346 (N_4346,N_3976,N_3995);
nand U4347 (N_4347,N_3902,N_3969);
or U4348 (N_4348,N_4191,N_4015);
nor U4349 (N_4349,N_4154,N_4140);
or U4350 (N_4350,N_3951,N_4150);
and U4351 (N_4351,N_4047,N_4189);
xnor U4352 (N_4352,N_3993,N_4083);
and U4353 (N_4353,N_3932,N_4088);
nand U4354 (N_4354,N_4084,N_3911);
xor U4355 (N_4355,N_4128,N_4169);
nor U4356 (N_4356,N_4143,N_4035);
or U4357 (N_4357,N_4106,N_4079);
or U4358 (N_4358,N_4181,N_4023);
nor U4359 (N_4359,N_4183,N_4084);
xnor U4360 (N_4360,N_3923,N_4097);
nor U4361 (N_4361,N_3913,N_4197);
and U4362 (N_4362,N_4089,N_4123);
nor U4363 (N_4363,N_4038,N_3972);
nand U4364 (N_4364,N_4061,N_4172);
and U4365 (N_4365,N_4105,N_3968);
or U4366 (N_4366,N_3970,N_4006);
nand U4367 (N_4367,N_3930,N_4123);
xor U4368 (N_4368,N_3964,N_4128);
xnor U4369 (N_4369,N_4176,N_4006);
and U4370 (N_4370,N_4191,N_4044);
nand U4371 (N_4371,N_3999,N_3964);
or U4372 (N_4372,N_4181,N_4152);
nand U4373 (N_4373,N_4053,N_4029);
nand U4374 (N_4374,N_4052,N_3930);
nand U4375 (N_4375,N_4055,N_3966);
nor U4376 (N_4376,N_3967,N_4091);
nand U4377 (N_4377,N_4092,N_4146);
or U4378 (N_4378,N_4070,N_4068);
or U4379 (N_4379,N_4090,N_3993);
and U4380 (N_4380,N_4116,N_3914);
xor U4381 (N_4381,N_4147,N_3967);
and U4382 (N_4382,N_4057,N_4177);
xnor U4383 (N_4383,N_4032,N_3902);
or U4384 (N_4384,N_3952,N_4180);
and U4385 (N_4385,N_4169,N_4197);
nand U4386 (N_4386,N_4127,N_3970);
nor U4387 (N_4387,N_4005,N_4115);
nor U4388 (N_4388,N_3934,N_3957);
and U4389 (N_4389,N_4190,N_3904);
nor U4390 (N_4390,N_3979,N_4071);
and U4391 (N_4391,N_4137,N_4167);
nor U4392 (N_4392,N_4160,N_4055);
and U4393 (N_4393,N_4182,N_4017);
or U4394 (N_4394,N_3934,N_4046);
or U4395 (N_4395,N_4180,N_4102);
or U4396 (N_4396,N_4013,N_3950);
xor U4397 (N_4397,N_4099,N_3978);
or U4398 (N_4398,N_3928,N_4000);
nand U4399 (N_4399,N_3983,N_3901);
and U4400 (N_4400,N_4074,N_4025);
xor U4401 (N_4401,N_3931,N_4140);
xor U4402 (N_4402,N_4130,N_4190);
nand U4403 (N_4403,N_4076,N_3917);
xor U4404 (N_4404,N_4120,N_3975);
nor U4405 (N_4405,N_4063,N_3951);
xnor U4406 (N_4406,N_3915,N_4096);
or U4407 (N_4407,N_3962,N_4072);
nand U4408 (N_4408,N_3907,N_4022);
nor U4409 (N_4409,N_3904,N_4056);
or U4410 (N_4410,N_4002,N_4196);
and U4411 (N_4411,N_4178,N_3927);
xnor U4412 (N_4412,N_4199,N_4057);
nand U4413 (N_4413,N_3922,N_4070);
xnor U4414 (N_4414,N_4188,N_3941);
xnor U4415 (N_4415,N_4007,N_4125);
nor U4416 (N_4416,N_3954,N_4055);
nand U4417 (N_4417,N_3983,N_4180);
xor U4418 (N_4418,N_3959,N_4146);
or U4419 (N_4419,N_4010,N_3924);
and U4420 (N_4420,N_4138,N_4146);
nand U4421 (N_4421,N_4121,N_3964);
nand U4422 (N_4422,N_3943,N_4060);
nor U4423 (N_4423,N_4119,N_4060);
nand U4424 (N_4424,N_4021,N_4107);
nand U4425 (N_4425,N_3941,N_3985);
nand U4426 (N_4426,N_3900,N_4045);
nand U4427 (N_4427,N_4165,N_4124);
nand U4428 (N_4428,N_4089,N_3945);
and U4429 (N_4429,N_4005,N_4053);
and U4430 (N_4430,N_3916,N_4157);
nand U4431 (N_4431,N_4075,N_4034);
nand U4432 (N_4432,N_4191,N_4070);
xor U4433 (N_4433,N_4193,N_4170);
nor U4434 (N_4434,N_4180,N_3972);
nor U4435 (N_4435,N_4030,N_4147);
nor U4436 (N_4436,N_4019,N_3931);
xnor U4437 (N_4437,N_3952,N_3949);
and U4438 (N_4438,N_3989,N_4037);
nor U4439 (N_4439,N_3923,N_4080);
nor U4440 (N_4440,N_4147,N_3994);
nand U4441 (N_4441,N_4189,N_3981);
nand U4442 (N_4442,N_4135,N_4140);
or U4443 (N_4443,N_4109,N_4199);
nand U4444 (N_4444,N_4018,N_4004);
nor U4445 (N_4445,N_4084,N_3936);
nor U4446 (N_4446,N_3908,N_3994);
or U4447 (N_4447,N_4180,N_3988);
nand U4448 (N_4448,N_4095,N_4111);
nor U4449 (N_4449,N_4164,N_4053);
nor U4450 (N_4450,N_4105,N_4115);
xnor U4451 (N_4451,N_4189,N_4049);
or U4452 (N_4452,N_4009,N_4100);
and U4453 (N_4453,N_4141,N_3970);
xnor U4454 (N_4454,N_4035,N_4109);
or U4455 (N_4455,N_4069,N_4182);
nor U4456 (N_4456,N_4064,N_4048);
nand U4457 (N_4457,N_4174,N_4185);
nor U4458 (N_4458,N_4069,N_4000);
xor U4459 (N_4459,N_3942,N_3978);
xor U4460 (N_4460,N_4018,N_4049);
or U4461 (N_4461,N_4054,N_3964);
xnor U4462 (N_4462,N_3929,N_4147);
or U4463 (N_4463,N_3986,N_4159);
and U4464 (N_4464,N_4073,N_3964);
xor U4465 (N_4465,N_4085,N_3966);
xnor U4466 (N_4466,N_4046,N_4029);
xnor U4467 (N_4467,N_4110,N_4089);
nor U4468 (N_4468,N_3929,N_3959);
nor U4469 (N_4469,N_4027,N_3941);
xor U4470 (N_4470,N_4184,N_3984);
xor U4471 (N_4471,N_3943,N_4054);
xnor U4472 (N_4472,N_4003,N_3961);
xnor U4473 (N_4473,N_4106,N_4033);
or U4474 (N_4474,N_3965,N_4017);
nand U4475 (N_4475,N_4135,N_3901);
and U4476 (N_4476,N_4089,N_3961);
or U4477 (N_4477,N_4091,N_4160);
xnor U4478 (N_4478,N_4030,N_3920);
nor U4479 (N_4479,N_4024,N_4027);
nor U4480 (N_4480,N_4148,N_4130);
nor U4481 (N_4481,N_3910,N_4070);
xnor U4482 (N_4482,N_4076,N_4002);
xor U4483 (N_4483,N_4134,N_3937);
xor U4484 (N_4484,N_3915,N_3980);
or U4485 (N_4485,N_4010,N_3900);
xnor U4486 (N_4486,N_4037,N_4027);
or U4487 (N_4487,N_4036,N_4115);
xor U4488 (N_4488,N_4072,N_4164);
nand U4489 (N_4489,N_4136,N_4001);
and U4490 (N_4490,N_4088,N_3998);
or U4491 (N_4491,N_3943,N_4059);
or U4492 (N_4492,N_4176,N_4127);
xnor U4493 (N_4493,N_3919,N_4072);
or U4494 (N_4494,N_4036,N_4080);
nand U4495 (N_4495,N_3994,N_3913);
nand U4496 (N_4496,N_3973,N_3965);
xor U4497 (N_4497,N_4141,N_3994);
and U4498 (N_4498,N_4026,N_4065);
nor U4499 (N_4499,N_4061,N_4049);
and U4500 (N_4500,N_4440,N_4260);
and U4501 (N_4501,N_4265,N_4415);
and U4502 (N_4502,N_4449,N_4295);
nand U4503 (N_4503,N_4427,N_4329);
and U4504 (N_4504,N_4497,N_4365);
xor U4505 (N_4505,N_4367,N_4202);
and U4506 (N_4506,N_4411,N_4481);
nand U4507 (N_4507,N_4320,N_4253);
xor U4508 (N_4508,N_4332,N_4483);
or U4509 (N_4509,N_4403,N_4257);
or U4510 (N_4510,N_4231,N_4454);
nand U4511 (N_4511,N_4331,N_4235);
or U4512 (N_4512,N_4315,N_4325);
and U4513 (N_4513,N_4416,N_4470);
xor U4514 (N_4514,N_4459,N_4418);
or U4515 (N_4515,N_4371,N_4254);
nor U4516 (N_4516,N_4467,N_4364);
nor U4517 (N_4517,N_4398,N_4323);
and U4518 (N_4518,N_4400,N_4296);
or U4519 (N_4519,N_4387,N_4232);
nor U4520 (N_4520,N_4443,N_4280);
xnor U4521 (N_4521,N_4362,N_4409);
nand U4522 (N_4522,N_4313,N_4351);
and U4523 (N_4523,N_4337,N_4247);
nand U4524 (N_4524,N_4203,N_4484);
xnor U4525 (N_4525,N_4300,N_4250);
or U4526 (N_4526,N_4356,N_4243);
and U4527 (N_4527,N_4264,N_4490);
xnor U4528 (N_4528,N_4368,N_4218);
nor U4529 (N_4529,N_4463,N_4432);
or U4530 (N_4530,N_4487,N_4405);
or U4531 (N_4531,N_4494,N_4468);
and U4532 (N_4532,N_4276,N_4294);
or U4533 (N_4533,N_4420,N_4486);
xor U4534 (N_4534,N_4471,N_4285);
nand U4535 (N_4535,N_4322,N_4397);
nor U4536 (N_4536,N_4346,N_4311);
nand U4537 (N_4537,N_4476,N_4386);
xnor U4538 (N_4538,N_4499,N_4248);
nor U4539 (N_4539,N_4357,N_4212);
or U4540 (N_4540,N_4225,N_4327);
xor U4541 (N_4541,N_4344,N_4431);
xor U4542 (N_4542,N_4422,N_4412);
and U4543 (N_4543,N_4413,N_4287);
nor U4544 (N_4544,N_4302,N_4338);
or U4545 (N_4545,N_4439,N_4293);
or U4546 (N_4546,N_4361,N_4414);
xnor U4547 (N_4547,N_4233,N_4430);
or U4548 (N_4548,N_4438,N_4474);
nand U4549 (N_4549,N_4259,N_4237);
xnor U4550 (N_4550,N_4215,N_4406);
xnor U4551 (N_4551,N_4230,N_4388);
nand U4552 (N_4552,N_4298,N_4282);
nor U4553 (N_4553,N_4214,N_4303);
and U4554 (N_4554,N_4429,N_4358);
xnor U4555 (N_4555,N_4348,N_4393);
or U4556 (N_4556,N_4426,N_4292);
or U4557 (N_4557,N_4316,N_4473);
or U4558 (N_4558,N_4442,N_4211);
xnor U4559 (N_4559,N_4434,N_4268);
nor U4560 (N_4560,N_4423,N_4223);
nand U4561 (N_4561,N_4339,N_4370);
nor U4562 (N_4562,N_4396,N_4301);
and U4563 (N_4563,N_4417,N_4226);
nor U4564 (N_4564,N_4465,N_4205);
nor U4565 (N_4565,N_4379,N_4290);
nor U4566 (N_4566,N_4381,N_4206);
nor U4567 (N_4567,N_4270,N_4385);
nor U4568 (N_4568,N_4217,N_4383);
or U4569 (N_4569,N_4389,N_4278);
or U4570 (N_4570,N_4275,N_4374);
nor U4571 (N_4571,N_4475,N_4450);
nor U4572 (N_4572,N_4466,N_4305);
or U4573 (N_4573,N_4283,N_4330);
nand U4574 (N_4574,N_4255,N_4221);
xor U4575 (N_4575,N_4343,N_4352);
nor U4576 (N_4576,N_4312,N_4273);
xnor U4577 (N_4577,N_4425,N_4266);
xor U4578 (N_4578,N_4355,N_4421);
or U4579 (N_4579,N_4261,N_4446);
and U4580 (N_4580,N_4216,N_4375);
or U4581 (N_4581,N_4314,N_4310);
xnor U4582 (N_4582,N_4469,N_4369);
nand U4583 (N_4583,N_4244,N_4492);
xnor U4584 (N_4584,N_4424,N_4213);
and U4585 (N_4585,N_4234,N_4324);
xnor U4586 (N_4586,N_4219,N_4384);
xnor U4587 (N_4587,N_4477,N_4391);
nand U4588 (N_4588,N_4222,N_4399);
nor U4589 (N_4589,N_4306,N_4460);
and U4590 (N_4590,N_4251,N_4491);
nand U4591 (N_4591,N_4263,N_4204);
nor U4592 (N_4592,N_4200,N_4286);
xnor U4593 (N_4593,N_4410,N_4291);
nor U4594 (N_4594,N_4373,N_4478);
nand U4595 (N_4595,N_4488,N_4239);
nor U4596 (N_4596,N_4453,N_4360);
nand U4597 (N_4597,N_4372,N_4359);
and U4598 (N_4598,N_4366,N_4240);
nand U4599 (N_4599,N_4493,N_4342);
or U4600 (N_4600,N_4267,N_4401);
or U4601 (N_4601,N_4209,N_4241);
nor U4602 (N_4602,N_4489,N_4318);
nand U4603 (N_4603,N_4402,N_4479);
nor U4604 (N_4604,N_4274,N_4377);
xor U4605 (N_4605,N_4363,N_4376);
or U4606 (N_4606,N_4228,N_4341);
nor U4607 (N_4607,N_4335,N_4269);
nor U4608 (N_4608,N_4350,N_4435);
and U4609 (N_4609,N_4307,N_4238);
and U4610 (N_4610,N_4245,N_4451);
xnor U4611 (N_4611,N_4256,N_4392);
nand U4612 (N_4612,N_4448,N_4437);
and U4613 (N_4613,N_4462,N_4229);
nor U4614 (N_4614,N_4224,N_4242);
and U4615 (N_4615,N_4317,N_4249);
nand U4616 (N_4616,N_4227,N_4445);
nor U4617 (N_4617,N_4408,N_4334);
or U4618 (N_4618,N_4279,N_4304);
and U4619 (N_4619,N_4433,N_4382);
nor U4620 (N_4620,N_4288,N_4452);
or U4621 (N_4621,N_4458,N_4395);
nor U4622 (N_4622,N_4210,N_4277);
nor U4623 (N_4623,N_4272,N_4281);
nor U4624 (N_4624,N_4353,N_4336);
xnor U4625 (N_4625,N_4419,N_4394);
xor U4626 (N_4626,N_4297,N_4326);
nand U4627 (N_4627,N_4252,N_4345);
and U4628 (N_4628,N_4461,N_4208);
nand U4629 (N_4629,N_4207,N_4495);
nand U4630 (N_4630,N_4407,N_4498);
xor U4631 (N_4631,N_4354,N_4404);
nor U4632 (N_4632,N_4308,N_4441);
nor U4633 (N_4633,N_4333,N_4378);
xor U4634 (N_4634,N_4444,N_4390);
nor U4635 (N_4635,N_4319,N_4428);
or U4636 (N_4636,N_4480,N_4455);
nor U4637 (N_4637,N_4347,N_4289);
xor U4638 (N_4638,N_4496,N_4284);
nand U4639 (N_4639,N_4246,N_4271);
nand U4640 (N_4640,N_4436,N_4220);
nand U4641 (N_4641,N_4236,N_4258);
and U4642 (N_4642,N_4299,N_4340);
or U4643 (N_4643,N_4464,N_4472);
and U4644 (N_4644,N_4349,N_4380);
and U4645 (N_4645,N_4457,N_4201);
nor U4646 (N_4646,N_4262,N_4447);
and U4647 (N_4647,N_4482,N_4456);
nor U4648 (N_4648,N_4321,N_4328);
xnor U4649 (N_4649,N_4309,N_4485);
nor U4650 (N_4650,N_4265,N_4250);
and U4651 (N_4651,N_4370,N_4396);
nand U4652 (N_4652,N_4314,N_4239);
or U4653 (N_4653,N_4381,N_4401);
nand U4654 (N_4654,N_4209,N_4473);
or U4655 (N_4655,N_4420,N_4241);
and U4656 (N_4656,N_4446,N_4426);
xor U4657 (N_4657,N_4400,N_4434);
nand U4658 (N_4658,N_4212,N_4289);
and U4659 (N_4659,N_4404,N_4229);
or U4660 (N_4660,N_4257,N_4376);
nand U4661 (N_4661,N_4375,N_4314);
and U4662 (N_4662,N_4234,N_4341);
nand U4663 (N_4663,N_4409,N_4491);
xor U4664 (N_4664,N_4494,N_4418);
or U4665 (N_4665,N_4413,N_4496);
xor U4666 (N_4666,N_4230,N_4203);
nand U4667 (N_4667,N_4301,N_4200);
nand U4668 (N_4668,N_4382,N_4263);
nor U4669 (N_4669,N_4237,N_4462);
nor U4670 (N_4670,N_4359,N_4225);
xnor U4671 (N_4671,N_4389,N_4221);
and U4672 (N_4672,N_4420,N_4350);
nor U4673 (N_4673,N_4313,N_4465);
xor U4674 (N_4674,N_4306,N_4483);
or U4675 (N_4675,N_4300,N_4401);
nor U4676 (N_4676,N_4424,N_4397);
xor U4677 (N_4677,N_4318,N_4471);
xor U4678 (N_4678,N_4282,N_4436);
and U4679 (N_4679,N_4344,N_4442);
nor U4680 (N_4680,N_4317,N_4371);
or U4681 (N_4681,N_4215,N_4210);
nor U4682 (N_4682,N_4233,N_4346);
and U4683 (N_4683,N_4362,N_4476);
nand U4684 (N_4684,N_4413,N_4400);
and U4685 (N_4685,N_4248,N_4396);
or U4686 (N_4686,N_4381,N_4287);
and U4687 (N_4687,N_4405,N_4307);
nand U4688 (N_4688,N_4293,N_4210);
xor U4689 (N_4689,N_4364,N_4495);
and U4690 (N_4690,N_4250,N_4395);
or U4691 (N_4691,N_4357,N_4435);
xor U4692 (N_4692,N_4305,N_4299);
nand U4693 (N_4693,N_4445,N_4281);
nor U4694 (N_4694,N_4334,N_4484);
xor U4695 (N_4695,N_4327,N_4322);
nor U4696 (N_4696,N_4345,N_4281);
nor U4697 (N_4697,N_4439,N_4415);
or U4698 (N_4698,N_4276,N_4495);
nand U4699 (N_4699,N_4208,N_4474);
nand U4700 (N_4700,N_4365,N_4296);
nor U4701 (N_4701,N_4246,N_4390);
or U4702 (N_4702,N_4428,N_4310);
nor U4703 (N_4703,N_4272,N_4287);
xnor U4704 (N_4704,N_4432,N_4351);
xnor U4705 (N_4705,N_4349,N_4272);
nor U4706 (N_4706,N_4359,N_4469);
and U4707 (N_4707,N_4331,N_4310);
nor U4708 (N_4708,N_4278,N_4269);
nor U4709 (N_4709,N_4399,N_4379);
nand U4710 (N_4710,N_4411,N_4470);
xor U4711 (N_4711,N_4488,N_4489);
and U4712 (N_4712,N_4417,N_4343);
or U4713 (N_4713,N_4267,N_4322);
and U4714 (N_4714,N_4233,N_4214);
nor U4715 (N_4715,N_4246,N_4430);
nor U4716 (N_4716,N_4462,N_4338);
xor U4717 (N_4717,N_4498,N_4351);
nor U4718 (N_4718,N_4211,N_4463);
xor U4719 (N_4719,N_4399,N_4338);
or U4720 (N_4720,N_4280,N_4334);
nand U4721 (N_4721,N_4401,N_4358);
nor U4722 (N_4722,N_4389,N_4355);
xnor U4723 (N_4723,N_4353,N_4375);
nor U4724 (N_4724,N_4202,N_4350);
nand U4725 (N_4725,N_4241,N_4404);
nand U4726 (N_4726,N_4311,N_4367);
nor U4727 (N_4727,N_4244,N_4368);
or U4728 (N_4728,N_4413,N_4318);
xor U4729 (N_4729,N_4226,N_4223);
xnor U4730 (N_4730,N_4496,N_4406);
and U4731 (N_4731,N_4425,N_4239);
nand U4732 (N_4732,N_4232,N_4419);
and U4733 (N_4733,N_4238,N_4356);
nor U4734 (N_4734,N_4207,N_4345);
xnor U4735 (N_4735,N_4219,N_4287);
and U4736 (N_4736,N_4245,N_4341);
and U4737 (N_4737,N_4309,N_4396);
nand U4738 (N_4738,N_4204,N_4499);
xor U4739 (N_4739,N_4441,N_4369);
nor U4740 (N_4740,N_4466,N_4259);
or U4741 (N_4741,N_4403,N_4416);
or U4742 (N_4742,N_4265,N_4258);
nor U4743 (N_4743,N_4403,N_4234);
xnor U4744 (N_4744,N_4478,N_4231);
and U4745 (N_4745,N_4276,N_4493);
or U4746 (N_4746,N_4342,N_4329);
and U4747 (N_4747,N_4230,N_4431);
and U4748 (N_4748,N_4277,N_4254);
nor U4749 (N_4749,N_4326,N_4490);
xnor U4750 (N_4750,N_4452,N_4379);
nor U4751 (N_4751,N_4298,N_4284);
or U4752 (N_4752,N_4327,N_4296);
and U4753 (N_4753,N_4405,N_4347);
nand U4754 (N_4754,N_4395,N_4373);
or U4755 (N_4755,N_4294,N_4481);
and U4756 (N_4756,N_4272,N_4480);
nor U4757 (N_4757,N_4438,N_4479);
nor U4758 (N_4758,N_4242,N_4390);
nor U4759 (N_4759,N_4404,N_4344);
nand U4760 (N_4760,N_4496,N_4410);
nand U4761 (N_4761,N_4367,N_4392);
or U4762 (N_4762,N_4362,N_4296);
xor U4763 (N_4763,N_4471,N_4380);
nor U4764 (N_4764,N_4221,N_4449);
or U4765 (N_4765,N_4429,N_4424);
or U4766 (N_4766,N_4410,N_4422);
or U4767 (N_4767,N_4355,N_4242);
nand U4768 (N_4768,N_4394,N_4364);
nand U4769 (N_4769,N_4336,N_4343);
nor U4770 (N_4770,N_4285,N_4442);
nand U4771 (N_4771,N_4396,N_4409);
xor U4772 (N_4772,N_4489,N_4345);
xor U4773 (N_4773,N_4449,N_4408);
xor U4774 (N_4774,N_4284,N_4432);
and U4775 (N_4775,N_4478,N_4292);
and U4776 (N_4776,N_4235,N_4460);
or U4777 (N_4777,N_4295,N_4248);
nand U4778 (N_4778,N_4463,N_4229);
nor U4779 (N_4779,N_4458,N_4424);
and U4780 (N_4780,N_4480,N_4413);
and U4781 (N_4781,N_4314,N_4225);
or U4782 (N_4782,N_4480,N_4357);
xor U4783 (N_4783,N_4439,N_4390);
nor U4784 (N_4784,N_4298,N_4280);
xor U4785 (N_4785,N_4337,N_4277);
and U4786 (N_4786,N_4273,N_4267);
nor U4787 (N_4787,N_4256,N_4283);
xnor U4788 (N_4788,N_4489,N_4413);
nand U4789 (N_4789,N_4359,N_4448);
or U4790 (N_4790,N_4495,N_4455);
nand U4791 (N_4791,N_4290,N_4473);
xnor U4792 (N_4792,N_4238,N_4295);
xnor U4793 (N_4793,N_4238,N_4288);
nand U4794 (N_4794,N_4322,N_4337);
nand U4795 (N_4795,N_4273,N_4406);
nor U4796 (N_4796,N_4363,N_4411);
nor U4797 (N_4797,N_4478,N_4356);
nand U4798 (N_4798,N_4400,N_4216);
and U4799 (N_4799,N_4384,N_4447);
nor U4800 (N_4800,N_4710,N_4587);
nand U4801 (N_4801,N_4607,N_4681);
nor U4802 (N_4802,N_4548,N_4533);
or U4803 (N_4803,N_4577,N_4591);
nand U4804 (N_4804,N_4702,N_4751);
and U4805 (N_4805,N_4638,N_4567);
nand U4806 (N_4806,N_4518,N_4568);
or U4807 (N_4807,N_4663,N_4620);
nand U4808 (N_4808,N_4783,N_4731);
nand U4809 (N_4809,N_4792,N_4606);
xnor U4810 (N_4810,N_4759,N_4537);
nor U4811 (N_4811,N_4570,N_4517);
nand U4812 (N_4812,N_4563,N_4747);
xnor U4813 (N_4813,N_4528,N_4791);
nor U4814 (N_4814,N_4616,N_4520);
nor U4815 (N_4815,N_4531,N_4544);
nor U4816 (N_4816,N_4772,N_4756);
nor U4817 (N_4817,N_4793,N_4505);
nand U4818 (N_4818,N_4562,N_4761);
or U4819 (N_4819,N_4569,N_4534);
or U4820 (N_4820,N_4704,N_4749);
or U4821 (N_4821,N_4526,N_4585);
xnor U4822 (N_4822,N_4615,N_4701);
xor U4823 (N_4823,N_4655,N_4629);
or U4824 (N_4824,N_4643,N_4797);
nand U4825 (N_4825,N_4672,N_4788);
nand U4826 (N_4826,N_4522,N_4546);
nor U4827 (N_4827,N_4547,N_4666);
and U4828 (N_4828,N_4727,N_4581);
nand U4829 (N_4829,N_4571,N_4769);
xnor U4830 (N_4830,N_4705,N_4694);
nor U4831 (N_4831,N_4765,N_4589);
and U4832 (N_4832,N_4550,N_4686);
nand U4833 (N_4833,N_4795,N_4778);
or U4834 (N_4834,N_4555,N_4665);
or U4835 (N_4835,N_4572,N_4541);
xnor U4836 (N_4836,N_4508,N_4594);
nand U4837 (N_4837,N_4636,N_4755);
and U4838 (N_4838,N_4692,N_4660);
or U4839 (N_4839,N_4733,N_4640);
and U4840 (N_4840,N_4651,N_4680);
and U4841 (N_4841,N_4623,N_4768);
nand U4842 (N_4842,N_4600,N_4584);
nor U4843 (N_4843,N_4646,N_4662);
xnor U4844 (N_4844,N_4762,N_4626);
nand U4845 (N_4845,N_4650,N_4599);
and U4846 (N_4846,N_4515,N_4529);
and U4847 (N_4847,N_4776,N_4763);
nor U4848 (N_4848,N_4743,N_4628);
xnor U4849 (N_4849,N_4794,N_4653);
or U4850 (N_4850,N_4746,N_4539);
and U4851 (N_4851,N_4545,N_4549);
xnor U4852 (N_4852,N_4595,N_4532);
and U4853 (N_4853,N_4516,N_4709);
nor U4854 (N_4854,N_4739,N_4698);
xnor U4855 (N_4855,N_4507,N_4513);
and U4856 (N_4856,N_4719,N_4784);
and U4857 (N_4857,N_4718,N_4503);
xor U4858 (N_4858,N_4566,N_4742);
and U4859 (N_4859,N_4675,N_4635);
and U4860 (N_4860,N_4699,N_4671);
or U4861 (N_4861,N_4676,N_4648);
nor U4862 (N_4862,N_4619,N_4559);
nor U4863 (N_4863,N_4734,N_4621);
nor U4864 (N_4864,N_4703,N_4735);
nor U4865 (N_4865,N_4542,N_4658);
and U4866 (N_4866,N_4752,N_4551);
or U4867 (N_4867,N_4576,N_4700);
or U4868 (N_4868,N_4780,N_4775);
or U4869 (N_4869,N_4717,N_4602);
or U4870 (N_4870,N_4707,N_4625);
nor U4871 (N_4871,N_4713,N_4682);
nor U4872 (N_4872,N_4564,N_4736);
nor U4873 (N_4873,N_4652,N_4524);
xor U4874 (N_4874,N_4732,N_4760);
nand U4875 (N_4875,N_4674,N_4512);
xor U4876 (N_4876,N_4668,N_4657);
nor U4877 (N_4877,N_4724,N_4538);
xor U4878 (N_4878,N_4501,N_4582);
nand U4879 (N_4879,N_4514,N_4553);
and U4880 (N_4880,N_4737,N_4504);
xnor U4881 (N_4881,N_4510,N_4774);
nor U4882 (N_4882,N_4575,N_4565);
nand U4883 (N_4883,N_4748,N_4716);
or U4884 (N_4884,N_4614,N_4767);
nand U4885 (N_4885,N_4624,N_4661);
nor U4886 (N_4886,N_4637,N_4771);
nor U4887 (N_4887,N_4678,N_4649);
and U4888 (N_4888,N_4593,N_4535);
and U4889 (N_4889,N_4723,N_4777);
and U4890 (N_4890,N_4521,N_4690);
xnor U4891 (N_4891,N_4779,N_4687);
xnor U4892 (N_4892,N_4622,N_4588);
xnor U4893 (N_4893,N_4645,N_4617);
and U4894 (N_4894,N_4740,N_4603);
xnor U4895 (N_4895,N_4509,N_4639);
xor U4896 (N_4896,N_4758,N_4711);
or U4897 (N_4897,N_4609,N_4722);
nor U4898 (N_4898,N_4506,N_4730);
or U4899 (N_4899,N_4706,N_4720);
xnor U4900 (N_4900,N_4691,N_4726);
nand U4901 (N_4901,N_4618,N_4738);
or U4902 (N_4902,N_4601,N_4789);
nand U4903 (N_4903,N_4592,N_4511);
or U4904 (N_4904,N_4627,N_4787);
xor U4905 (N_4905,N_4673,N_4502);
xnor U4906 (N_4906,N_4688,N_4561);
nor U4907 (N_4907,N_4525,N_4679);
nand U4908 (N_4908,N_4630,N_4697);
nor U4909 (N_4909,N_4741,N_4696);
xor U4910 (N_4910,N_4745,N_4764);
nor U4911 (N_4911,N_4770,N_4667);
xnor U4912 (N_4912,N_4611,N_4631);
and U4913 (N_4913,N_4790,N_4725);
nand U4914 (N_4914,N_4540,N_4560);
nand U4915 (N_4915,N_4766,N_4798);
and U4916 (N_4916,N_4586,N_4580);
nand U4917 (N_4917,N_4573,N_4659);
and U4918 (N_4918,N_4590,N_4664);
xor U4919 (N_4919,N_4574,N_4683);
or U4920 (N_4920,N_4557,N_4796);
xor U4921 (N_4921,N_4543,N_4632);
nor U4922 (N_4922,N_4527,N_4597);
or U4923 (N_4923,N_4695,N_4799);
nand U4924 (N_4924,N_4721,N_4744);
or U4925 (N_4925,N_4786,N_4536);
and U4926 (N_4926,N_4684,N_4583);
or U4927 (N_4927,N_4608,N_4754);
nand U4928 (N_4928,N_4728,N_4785);
nor U4929 (N_4929,N_4750,N_4523);
or U4930 (N_4930,N_4500,N_4579);
or U4931 (N_4931,N_4644,N_4782);
xor U4932 (N_4932,N_4712,N_4530);
nand U4933 (N_4933,N_4670,N_4604);
or U4934 (N_4934,N_4689,N_4610);
xnor U4935 (N_4935,N_4685,N_4654);
xnor U4936 (N_4936,N_4773,N_4598);
nand U4937 (N_4937,N_4641,N_4552);
xnor U4938 (N_4938,N_4729,N_4757);
nor U4939 (N_4939,N_4633,N_4613);
xnor U4940 (N_4940,N_4714,N_4656);
nor U4941 (N_4941,N_4647,N_4634);
nand U4942 (N_4942,N_4693,N_4715);
and U4943 (N_4943,N_4753,N_4558);
xor U4944 (N_4944,N_4642,N_4669);
nand U4945 (N_4945,N_4612,N_4677);
or U4946 (N_4946,N_4554,N_4519);
nor U4947 (N_4947,N_4596,N_4605);
or U4948 (N_4948,N_4578,N_4708);
and U4949 (N_4949,N_4781,N_4556);
or U4950 (N_4950,N_4760,N_4549);
or U4951 (N_4951,N_4687,N_4613);
and U4952 (N_4952,N_4684,N_4657);
nand U4953 (N_4953,N_4686,N_4551);
nand U4954 (N_4954,N_4632,N_4785);
or U4955 (N_4955,N_4601,N_4573);
nor U4956 (N_4956,N_4777,N_4525);
nand U4957 (N_4957,N_4768,N_4770);
and U4958 (N_4958,N_4578,N_4779);
nor U4959 (N_4959,N_4646,N_4571);
nand U4960 (N_4960,N_4564,N_4547);
nand U4961 (N_4961,N_4728,N_4749);
nand U4962 (N_4962,N_4661,N_4700);
xnor U4963 (N_4963,N_4771,N_4620);
nor U4964 (N_4964,N_4590,N_4651);
xor U4965 (N_4965,N_4515,N_4503);
or U4966 (N_4966,N_4702,N_4735);
xor U4967 (N_4967,N_4741,N_4738);
nor U4968 (N_4968,N_4647,N_4696);
nor U4969 (N_4969,N_4514,N_4678);
xor U4970 (N_4970,N_4653,N_4529);
nand U4971 (N_4971,N_4777,N_4570);
xnor U4972 (N_4972,N_4695,N_4614);
xnor U4973 (N_4973,N_4695,N_4598);
and U4974 (N_4974,N_4632,N_4731);
nand U4975 (N_4975,N_4699,N_4741);
nor U4976 (N_4976,N_4523,N_4743);
nor U4977 (N_4977,N_4775,N_4521);
or U4978 (N_4978,N_4749,N_4569);
xor U4979 (N_4979,N_4638,N_4626);
and U4980 (N_4980,N_4654,N_4785);
and U4981 (N_4981,N_4585,N_4659);
and U4982 (N_4982,N_4552,N_4687);
nor U4983 (N_4983,N_4525,N_4601);
nor U4984 (N_4984,N_4593,N_4564);
or U4985 (N_4985,N_4714,N_4596);
nand U4986 (N_4986,N_4601,N_4527);
nor U4987 (N_4987,N_4600,N_4528);
or U4988 (N_4988,N_4597,N_4718);
nand U4989 (N_4989,N_4750,N_4543);
nand U4990 (N_4990,N_4798,N_4764);
or U4991 (N_4991,N_4656,N_4617);
or U4992 (N_4992,N_4775,N_4582);
and U4993 (N_4993,N_4721,N_4539);
or U4994 (N_4994,N_4605,N_4512);
nand U4995 (N_4995,N_4679,N_4502);
xor U4996 (N_4996,N_4631,N_4639);
xnor U4997 (N_4997,N_4711,N_4681);
xnor U4998 (N_4998,N_4512,N_4739);
nor U4999 (N_4999,N_4572,N_4778);
xnor U5000 (N_5000,N_4789,N_4654);
xor U5001 (N_5001,N_4655,N_4625);
or U5002 (N_5002,N_4751,N_4740);
and U5003 (N_5003,N_4701,N_4790);
nor U5004 (N_5004,N_4514,N_4776);
and U5005 (N_5005,N_4602,N_4791);
nand U5006 (N_5006,N_4739,N_4610);
nor U5007 (N_5007,N_4775,N_4651);
and U5008 (N_5008,N_4570,N_4628);
or U5009 (N_5009,N_4518,N_4697);
nand U5010 (N_5010,N_4676,N_4737);
xnor U5011 (N_5011,N_4630,N_4773);
nor U5012 (N_5012,N_4562,N_4523);
nor U5013 (N_5013,N_4765,N_4629);
xnor U5014 (N_5014,N_4713,N_4762);
nand U5015 (N_5015,N_4600,N_4518);
xor U5016 (N_5016,N_4526,N_4684);
or U5017 (N_5017,N_4573,N_4641);
or U5018 (N_5018,N_4545,N_4749);
and U5019 (N_5019,N_4661,N_4752);
or U5020 (N_5020,N_4760,N_4632);
xor U5021 (N_5021,N_4691,N_4573);
xor U5022 (N_5022,N_4648,N_4554);
and U5023 (N_5023,N_4704,N_4667);
or U5024 (N_5024,N_4637,N_4798);
nand U5025 (N_5025,N_4697,N_4607);
nand U5026 (N_5026,N_4793,N_4767);
xnor U5027 (N_5027,N_4575,N_4770);
nor U5028 (N_5028,N_4765,N_4789);
xor U5029 (N_5029,N_4506,N_4625);
nand U5030 (N_5030,N_4612,N_4699);
and U5031 (N_5031,N_4511,N_4700);
and U5032 (N_5032,N_4579,N_4713);
and U5033 (N_5033,N_4732,N_4616);
nor U5034 (N_5034,N_4687,N_4617);
nor U5035 (N_5035,N_4767,N_4678);
nor U5036 (N_5036,N_4576,N_4549);
nor U5037 (N_5037,N_4687,N_4736);
xnor U5038 (N_5038,N_4660,N_4595);
nand U5039 (N_5039,N_4526,N_4757);
and U5040 (N_5040,N_4603,N_4705);
nand U5041 (N_5041,N_4509,N_4725);
and U5042 (N_5042,N_4683,N_4596);
and U5043 (N_5043,N_4796,N_4685);
or U5044 (N_5044,N_4603,N_4791);
or U5045 (N_5045,N_4639,N_4711);
and U5046 (N_5046,N_4687,N_4790);
nand U5047 (N_5047,N_4700,N_4600);
nor U5048 (N_5048,N_4775,N_4770);
nor U5049 (N_5049,N_4560,N_4799);
and U5050 (N_5050,N_4758,N_4619);
nor U5051 (N_5051,N_4688,N_4544);
nand U5052 (N_5052,N_4548,N_4772);
and U5053 (N_5053,N_4795,N_4690);
and U5054 (N_5054,N_4663,N_4758);
nand U5055 (N_5055,N_4509,N_4562);
and U5056 (N_5056,N_4517,N_4613);
or U5057 (N_5057,N_4616,N_4714);
or U5058 (N_5058,N_4708,N_4565);
nand U5059 (N_5059,N_4511,N_4712);
nor U5060 (N_5060,N_4536,N_4791);
or U5061 (N_5061,N_4591,N_4730);
xnor U5062 (N_5062,N_4687,N_4523);
nor U5063 (N_5063,N_4560,N_4667);
xor U5064 (N_5064,N_4705,N_4714);
and U5065 (N_5065,N_4764,N_4548);
xor U5066 (N_5066,N_4756,N_4752);
nand U5067 (N_5067,N_4717,N_4551);
or U5068 (N_5068,N_4725,N_4629);
nor U5069 (N_5069,N_4603,N_4780);
nand U5070 (N_5070,N_4639,N_4642);
nor U5071 (N_5071,N_4724,N_4587);
xnor U5072 (N_5072,N_4574,N_4566);
xor U5073 (N_5073,N_4601,N_4745);
xor U5074 (N_5074,N_4710,N_4767);
or U5075 (N_5075,N_4791,N_4700);
or U5076 (N_5076,N_4548,N_4771);
and U5077 (N_5077,N_4738,N_4597);
xor U5078 (N_5078,N_4623,N_4595);
nor U5079 (N_5079,N_4744,N_4686);
nand U5080 (N_5080,N_4735,N_4767);
or U5081 (N_5081,N_4759,N_4541);
and U5082 (N_5082,N_4543,N_4714);
nand U5083 (N_5083,N_4770,N_4681);
nand U5084 (N_5084,N_4571,N_4595);
xnor U5085 (N_5085,N_4618,N_4743);
nand U5086 (N_5086,N_4531,N_4612);
nand U5087 (N_5087,N_4708,N_4549);
and U5088 (N_5088,N_4530,N_4731);
or U5089 (N_5089,N_4505,N_4703);
or U5090 (N_5090,N_4792,N_4528);
xor U5091 (N_5091,N_4740,N_4647);
xnor U5092 (N_5092,N_4524,N_4727);
nor U5093 (N_5093,N_4640,N_4503);
or U5094 (N_5094,N_4738,N_4568);
and U5095 (N_5095,N_4753,N_4600);
or U5096 (N_5096,N_4536,N_4739);
and U5097 (N_5097,N_4618,N_4622);
nor U5098 (N_5098,N_4607,N_4775);
or U5099 (N_5099,N_4661,N_4586);
or U5100 (N_5100,N_5053,N_4934);
or U5101 (N_5101,N_5089,N_4950);
nand U5102 (N_5102,N_5095,N_5062);
nor U5103 (N_5103,N_4867,N_5022);
nand U5104 (N_5104,N_5086,N_4818);
xor U5105 (N_5105,N_4802,N_4894);
nor U5106 (N_5106,N_5085,N_5083);
and U5107 (N_5107,N_5060,N_5004);
nor U5108 (N_5108,N_4920,N_5021);
and U5109 (N_5109,N_5009,N_4907);
xor U5110 (N_5110,N_4979,N_4895);
and U5111 (N_5111,N_5065,N_4921);
xnor U5112 (N_5112,N_5034,N_5032);
nor U5113 (N_5113,N_4836,N_5033);
nor U5114 (N_5114,N_4838,N_5023);
nor U5115 (N_5115,N_4893,N_5002);
nand U5116 (N_5116,N_4885,N_4900);
and U5117 (N_5117,N_5097,N_4994);
or U5118 (N_5118,N_4884,N_5045);
nor U5119 (N_5119,N_5027,N_5000);
nor U5120 (N_5120,N_4957,N_4990);
or U5121 (N_5121,N_5092,N_4974);
or U5122 (N_5122,N_4846,N_4826);
nand U5123 (N_5123,N_5049,N_4830);
and U5124 (N_5124,N_4819,N_4806);
xnor U5125 (N_5125,N_4856,N_4828);
nor U5126 (N_5126,N_4824,N_4959);
nor U5127 (N_5127,N_4869,N_4993);
or U5128 (N_5128,N_4937,N_4804);
nand U5129 (N_5129,N_4968,N_4809);
and U5130 (N_5130,N_4963,N_5082);
or U5131 (N_5131,N_4919,N_4940);
or U5132 (N_5132,N_5016,N_4949);
or U5133 (N_5133,N_4999,N_5063);
nand U5134 (N_5134,N_5044,N_5019);
or U5135 (N_5135,N_4967,N_4803);
and U5136 (N_5136,N_4878,N_4813);
and U5137 (N_5137,N_5068,N_4850);
or U5138 (N_5138,N_4890,N_4834);
nand U5139 (N_5139,N_4989,N_5001);
xnor U5140 (N_5140,N_5061,N_4960);
or U5141 (N_5141,N_5037,N_4896);
nor U5142 (N_5142,N_4935,N_4945);
nor U5143 (N_5143,N_5028,N_5098);
nand U5144 (N_5144,N_4808,N_4975);
nand U5145 (N_5145,N_4970,N_4859);
nand U5146 (N_5146,N_5057,N_5025);
or U5147 (N_5147,N_4978,N_5003);
or U5148 (N_5148,N_4964,N_4868);
xnor U5149 (N_5149,N_4953,N_5052);
and U5150 (N_5150,N_4833,N_4936);
nand U5151 (N_5151,N_4906,N_5040);
xnor U5152 (N_5152,N_5073,N_5077);
nand U5153 (N_5153,N_4955,N_5013);
or U5154 (N_5154,N_4817,N_4944);
nand U5155 (N_5155,N_4841,N_4984);
nand U5156 (N_5156,N_5030,N_4837);
xor U5157 (N_5157,N_4961,N_4938);
or U5158 (N_5158,N_4962,N_5043);
and U5159 (N_5159,N_4827,N_4872);
nand U5160 (N_5160,N_4857,N_4845);
nand U5161 (N_5161,N_4849,N_5017);
or U5162 (N_5162,N_5054,N_4913);
nand U5163 (N_5163,N_5076,N_4998);
xor U5164 (N_5164,N_5014,N_5080);
or U5165 (N_5165,N_5048,N_5024);
nor U5166 (N_5166,N_5051,N_4946);
xnor U5167 (N_5167,N_4880,N_4996);
xnor U5168 (N_5168,N_4928,N_4914);
nor U5169 (N_5169,N_4892,N_4982);
nand U5170 (N_5170,N_4924,N_4917);
nor U5171 (N_5171,N_4882,N_4981);
and U5172 (N_5172,N_4911,N_4821);
xnor U5173 (N_5173,N_5041,N_4814);
nand U5174 (N_5174,N_4988,N_4898);
or U5175 (N_5175,N_4932,N_5078);
or U5176 (N_5176,N_4925,N_4948);
nor U5177 (N_5177,N_4939,N_5042);
or U5178 (N_5178,N_5020,N_4825);
and U5179 (N_5179,N_5059,N_4875);
or U5180 (N_5180,N_4983,N_4903);
nor U5181 (N_5181,N_4901,N_4865);
nand U5182 (N_5182,N_4943,N_4822);
nor U5183 (N_5183,N_5067,N_4816);
xor U5184 (N_5184,N_4972,N_4973);
or U5185 (N_5185,N_4874,N_4966);
and U5186 (N_5186,N_4855,N_5079);
nor U5187 (N_5187,N_5047,N_5055);
nor U5188 (N_5188,N_4941,N_4801);
or U5189 (N_5189,N_4860,N_4992);
nor U5190 (N_5190,N_4876,N_4862);
and U5191 (N_5191,N_4812,N_4969);
and U5192 (N_5192,N_5072,N_4887);
nand U5193 (N_5193,N_4861,N_5036);
nor U5194 (N_5194,N_4930,N_4976);
nand U5195 (N_5195,N_4977,N_5090);
xor U5196 (N_5196,N_5094,N_4954);
or U5197 (N_5197,N_5070,N_5026);
xor U5198 (N_5198,N_5091,N_4839);
nand U5199 (N_5199,N_5029,N_4870);
and U5200 (N_5200,N_4985,N_4971);
nand U5201 (N_5201,N_4915,N_4829);
nor U5202 (N_5202,N_5038,N_4888);
nand U5203 (N_5203,N_4986,N_4958);
or U5204 (N_5204,N_5046,N_4931);
nand U5205 (N_5205,N_4891,N_5007);
xnor U5206 (N_5206,N_4852,N_4922);
or U5207 (N_5207,N_4866,N_4899);
and U5208 (N_5208,N_5006,N_4987);
nor U5209 (N_5209,N_4897,N_4800);
nand U5210 (N_5210,N_4807,N_5035);
nand U5211 (N_5211,N_4811,N_5050);
nor U5212 (N_5212,N_4854,N_5064);
xor U5213 (N_5213,N_4835,N_4923);
nand U5214 (N_5214,N_4909,N_5093);
xnor U5215 (N_5215,N_4995,N_4951);
nor U5216 (N_5216,N_4805,N_4933);
and U5217 (N_5217,N_4810,N_4881);
nor U5218 (N_5218,N_4908,N_5075);
or U5219 (N_5219,N_5015,N_5088);
nor U5220 (N_5220,N_5011,N_4926);
or U5221 (N_5221,N_5099,N_4905);
nor U5222 (N_5222,N_5010,N_5056);
nand U5223 (N_5223,N_4873,N_5081);
xnor U5224 (N_5224,N_4952,N_4886);
or U5225 (N_5225,N_5005,N_5031);
nand U5226 (N_5226,N_4820,N_4847);
xor U5227 (N_5227,N_4844,N_5084);
or U5228 (N_5228,N_5008,N_4863);
nor U5229 (N_5229,N_4912,N_4956);
xnor U5230 (N_5230,N_4918,N_5074);
or U5231 (N_5231,N_4965,N_4879);
xor U5232 (N_5232,N_4997,N_4927);
nand U5233 (N_5233,N_5039,N_4904);
or U5234 (N_5234,N_4902,N_5012);
and U5235 (N_5235,N_5058,N_5096);
nand U5236 (N_5236,N_4815,N_4877);
xor U5237 (N_5237,N_4851,N_5071);
xnor U5238 (N_5238,N_4858,N_5018);
or U5239 (N_5239,N_5087,N_4843);
nor U5240 (N_5240,N_4929,N_4916);
nor U5241 (N_5241,N_4871,N_4864);
xor U5242 (N_5242,N_4853,N_4980);
nand U5243 (N_5243,N_4889,N_4942);
nor U5244 (N_5244,N_4840,N_4823);
nand U5245 (N_5245,N_5066,N_5069);
nand U5246 (N_5246,N_4910,N_4842);
and U5247 (N_5247,N_4848,N_4991);
and U5248 (N_5248,N_4832,N_4883);
nand U5249 (N_5249,N_4947,N_4831);
nor U5250 (N_5250,N_5005,N_5093);
and U5251 (N_5251,N_4964,N_4973);
xnor U5252 (N_5252,N_4887,N_4972);
or U5253 (N_5253,N_4873,N_4967);
xor U5254 (N_5254,N_4982,N_4922);
nand U5255 (N_5255,N_5033,N_5011);
nor U5256 (N_5256,N_4976,N_5085);
and U5257 (N_5257,N_5020,N_4946);
or U5258 (N_5258,N_4938,N_4948);
and U5259 (N_5259,N_5048,N_4889);
or U5260 (N_5260,N_4988,N_4814);
or U5261 (N_5261,N_5095,N_4847);
xnor U5262 (N_5262,N_5086,N_5011);
nor U5263 (N_5263,N_5029,N_4880);
xor U5264 (N_5264,N_5031,N_4866);
nor U5265 (N_5265,N_4979,N_4871);
or U5266 (N_5266,N_4949,N_5049);
or U5267 (N_5267,N_5082,N_5008);
nor U5268 (N_5268,N_4995,N_5063);
or U5269 (N_5269,N_5047,N_4883);
and U5270 (N_5270,N_4927,N_5065);
or U5271 (N_5271,N_5025,N_4994);
xnor U5272 (N_5272,N_5027,N_4850);
and U5273 (N_5273,N_5023,N_4933);
nand U5274 (N_5274,N_5085,N_4980);
nor U5275 (N_5275,N_5034,N_4909);
nand U5276 (N_5276,N_5058,N_4996);
nor U5277 (N_5277,N_4920,N_4997);
and U5278 (N_5278,N_4856,N_4811);
nand U5279 (N_5279,N_4942,N_4823);
and U5280 (N_5280,N_4901,N_4878);
nand U5281 (N_5281,N_4932,N_4982);
xnor U5282 (N_5282,N_4877,N_4961);
xor U5283 (N_5283,N_5008,N_4818);
and U5284 (N_5284,N_4841,N_5018);
nand U5285 (N_5285,N_4941,N_5060);
nor U5286 (N_5286,N_5026,N_5036);
or U5287 (N_5287,N_5041,N_4880);
or U5288 (N_5288,N_4826,N_4896);
nor U5289 (N_5289,N_4980,N_5015);
xor U5290 (N_5290,N_4963,N_5029);
nand U5291 (N_5291,N_4995,N_5021);
xor U5292 (N_5292,N_4812,N_4992);
nand U5293 (N_5293,N_4907,N_4872);
and U5294 (N_5294,N_5045,N_4906);
nand U5295 (N_5295,N_5041,N_5021);
nand U5296 (N_5296,N_5070,N_4965);
and U5297 (N_5297,N_4854,N_4972);
nor U5298 (N_5298,N_4859,N_4923);
or U5299 (N_5299,N_5086,N_4968);
nor U5300 (N_5300,N_5006,N_4895);
xor U5301 (N_5301,N_4942,N_4976);
xor U5302 (N_5302,N_5026,N_4956);
and U5303 (N_5303,N_5079,N_5036);
nand U5304 (N_5304,N_5050,N_5064);
nor U5305 (N_5305,N_4956,N_4913);
and U5306 (N_5306,N_4867,N_4957);
nor U5307 (N_5307,N_4976,N_4952);
or U5308 (N_5308,N_4837,N_4960);
xor U5309 (N_5309,N_5040,N_4810);
or U5310 (N_5310,N_4872,N_5096);
and U5311 (N_5311,N_4930,N_4830);
nand U5312 (N_5312,N_4877,N_4950);
nand U5313 (N_5313,N_4979,N_5041);
and U5314 (N_5314,N_4863,N_4904);
or U5315 (N_5315,N_4825,N_5004);
nor U5316 (N_5316,N_4878,N_5015);
nor U5317 (N_5317,N_5021,N_4948);
and U5318 (N_5318,N_4934,N_4852);
and U5319 (N_5319,N_4845,N_4937);
nor U5320 (N_5320,N_5027,N_4913);
xor U5321 (N_5321,N_5013,N_4892);
xor U5322 (N_5322,N_4890,N_4845);
xnor U5323 (N_5323,N_4888,N_5061);
and U5324 (N_5324,N_4968,N_4915);
nand U5325 (N_5325,N_5015,N_5099);
nor U5326 (N_5326,N_4973,N_4914);
nand U5327 (N_5327,N_5078,N_4827);
or U5328 (N_5328,N_4827,N_5093);
or U5329 (N_5329,N_5060,N_5098);
xnor U5330 (N_5330,N_5005,N_5079);
nand U5331 (N_5331,N_4960,N_5024);
or U5332 (N_5332,N_5061,N_4868);
xnor U5333 (N_5333,N_5071,N_4816);
or U5334 (N_5334,N_4950,N_4891);
and U5335 (N_5335,N_5087,N_4969);
and U5336 (N_5336,N_5079,N_4831);
nand U5337 (N_5337,N_4858,N_5043);
or U5338 (N_5338,N_4812,N_4873);
and U5339 (N_5339,N_4880,N_4975);
and U5340 (N_5340,N_5020,N_4925);
nand U5341 (N_5341,N_4989,N_4992);
or U5342 (N_5342,N_4885,N_4825);
nor U5343 (N_5343,N_4920,N_4892);
and U5344 (N_5344,N_4912,N_4918);
and U5345 (N_5345,N_4941,N_5088);
nand U5346 (N_5346,N_4863,N_5003);
or U5347 (N_5347,N_4934,N_5058);
nand U5348 (N_5348,N_4896,N_4892);
and U5349 (N_5349,N_4881,N_5043);
nor U5350 (N_5350,N_4964,N_4990);
and U5351 (N_5351,N_4886,N_4839);
nor U5352 (N_5352,N_4995,N_5098);
and U5353 (N_5353,N_5027,N_4985);
nor U5354 (N_5354,N_4969,N_4926);
nor U5355 (N_5355,N_5086,N_5098);
nand U5356 (N_5356,N_5072,N_4868);
xnor U5357 (N_5357,N_4916,N_5046);
xnor U5358 (N_5358,N_4934,N_4959);
nor U5359 (N_5359,N_4844,N_4846);
nand U5360 (N_5360,N_4964,N_4807);
nand U5361 (N_5361,N_4922,N_4826);
and U5362 (N_5362,N_4965,N_5071);
or U5363 (N_5363,N_4817,N_4953);
or U5364 (N_5364,N_5020,N_5046);
and U5365 (N_5365,N_5049,N_4980);
or U5366 (N_5366,N_4887,N_5029);
and U5367 (N_5367,N_4926,N_5054);
and U5368 (N_5368,N_5098,N_4916);
xnor U5369 (N_5369,N_4971,N_5075);
nor U5370 (N_5370,N_4929,N_4897);
xor U5371 (N_5371,N_4984,N_5037);
xnor U5372 (N_5372,N_4896,N_5051);
nand U5373 (N_5373,N_5098,N_4996);
nand U5374 (N_5374,N_5057,N_4880);
or U5375 (N_5375,N_4937,N_4958);
and U5376 (N_5376,N_5079,N_5073);
or U5377 (N_5377,N_4937,N_4933);
xor U5378 (N_5378,N_5002,N_5045);
and U5379 (N_5379,N_4876,N_4932);
nor U5380 (N_5380,N_4878,N_4994);
or U5381 (N_5381,N_4973,N_4818);
and U5382 (N_5382,N_5027,N_5059);
nor U5383 (N_5383,N_4905,N_5007);
nand U5384 (N_5384,N_4908,N_4936);
nor U5385 (N_5385,N_5024,N_4936);
xor U5386 (N_5386,N_4808,N_5091);
xnor U5387 (N_5387,N_5058,N_4931);
or U5388 (N_5388,N_4825,N_4919);
or U5389 (N_5389,N_4982,N_4965);
xnor U5390 (N_5390,N_4900,N_4913);
or U5391 (N_5391,N_4904,N_4807);
and U5392 (N_5392,N_4810,N_4858);
xnor U5393 (N_5393,N_5072,N_5041);
nand U5394 (N_5394,N_5076,N_4974);
or U5395 (N_5395,N_5043,N_4906);
or U5396 (N_5396,N_5081,N_4997);
xnor U5397 (N_5397,N_4828,N_5091);
and U5398 (N_5398,N_4842,N_4819);
or U5399 (N_5399,N_4935,N_5094);
nor U5400 (N_5400,N_5157,N_5345);
nand U5401 (N_5401,N_5287,N_5343);
xor U5402 (N_5402,N_5331,N_5192);
or U5403 (N_5403,N_5111,N_5377);
and U5404 (N_5404,N_5272,N_5254);
nor U5405 (N_5405,N_5125,N_5362);
and U5406 (N_5406,N_5222,N_5285);
nand U5407 (N_5407,N_5198,N_5102);
or U5408 (N_5408,N_5197,N_5283);
xnor U5409 (N_5409,N_5309,N_5239);
or U5410 (N_5410,N_5129,N_5316);
xnor U5411 (N_5411,N_5124,N_5349);
nor U5412 (N_5412,N_5258,N_5333);
xnor U5413 (N_5413,N_5325,N_5218);
and U5414 (N_5414,N_5302,N_5107);
xnor U5415 (N_5415,N_5312,N_5207);
xnor U5416 (N_5416,N_5127,N_5373);
or U5417 (N_5417,N_5137,N_5242);
xnor U5418 (N_5418,N_5162,N_5251);
nor U5419 (N_5419,N_5217,N_5147);
xor U5420 (N_5420,N_5255,N_5216);
and U5421 (N_5421,N_5173,N_5398);
nor U5422 (N_5422,N_5306,N_5115);
nand U5423 (N_5423,N_5353,N_5243);
and U5424 (N_5424,N_5322,N_5361);
nor U5425 (N_5425,N_5194,N_5152);
nand U5426 (N_5426,N_5391,N_5295);
nand U5427 (N_5427,N_5390,N_5387);
xnor U5428 (N_5428,N_5269,N_5143);
nor U5429 (N_5429,N_5342,N_5290);
or U5430 (N_5430,N_5165,N_5376);
nor U5431 (N_5431,N_5246,N_5153);
nor U5432 (N_5432,N_5378,N_5106);
xnor U5433 (N_5433,N_5151,N_5108);
nand U5434 (N_5434,N_5317,N_5277);
and U5435 (N_5435,N_5122,N_5100);
or U5436 (N_5436,N_5134,N_5148);
xor U5437 (N_5437,N_5381,N_5275);
and U5438 (N_5438,N_5367,N_5346);
nor U5439 (N_5439,N_5266,N_5365);
nor U5440 (N_5440,N_5109,N_5307);
nand U5441 (N_5441,N_5227,N_5232);
and U5442 (N_5442,N_5224,N_5288);
or U5443 (N_5443,N_5163,N_5399);
nor U5444 (N_5444,N_5313,N_5181);
xnor U5445 (N_5445,N_5369,N_5344);
nor U5446 (N_5446,N_5264,N_5187);
nand U5447 (N_5447,N_5291,N_5319);
nor U5448 (N_5448,N_5136,N_5237);
nand U5449 (N_5449,N_5328,N_5238);
nand U5450 (N_5450,N_5179,N_5171);
or U5451 (N_5451,N_5372,N_5248);
xor U5452 (N_5452,N_5204,N_5155);
xnor U5453 (N_5453,N_5395,N_5303);
or U5454 (N_5454,N_5371,N_5123);
nand U5455 (N_5455,N_5253,N_5357);
and U5456 (N_5456,N_5105,N_5249);
xor U5457 (N_5457,N_5396,N_5375);
and U5458 (N_5458,N_5265,N_5310);
and U5459 (N_5459,N_5347,N_5178);
or U5460 (N_5460,N_5300,N_5208);
or U5461 (N_5461,N_5268,N_5286);
and U5462 (N_5462,N_5104,N_5219);
or U5463 (N_5463,N_5182,N_5339);
nand U5464 (N_5464,N_5235,N_5386);
nor U5465 (N_5465,N_5281,N_5118);
and U5466 (N_5466,N_5128,N_5259);
xnor U5467 (N_5467,N_5220,N_5247);
nor U5468 (N_5468,N_5330,N_5233);
xor U5469 (N_5469,N_5358,N_5209);
nand U5470 (N_5470,N_5341,N_5210);
and U5471 (N_5471,N_5298,N_5267);
xnor U5472 (N_5472,N_5256,N_5245);
and U5473 (N_5473,N_5366,N_5379);
xor U5474 (N_5474,N_5324,N_5289);
xor U5475 (N_5475,N_5223,N_5314);
nor U5476 (N_5476,N_5190,N_5212);
xor U5477 (N_5477,N_5392,N_5160);
nand U5478 (N_5478,N_5299,N_5323);
xor U5479 (N_5479,N_5292,N_5282);
or U5480 (N_5480,N_5119,N_5229);
xor U5481 (N_5481,N_5241,N_5389);
or U5482 (N_5482,N_5294,N_5196);
xnor U5483 (N_5483,N_5296,N_5318);
or U5484 (N_5484,N_5188,N_5203);
and U5485 (N_5485,N_5360,N_5189);
xor U5486 (N_5486,N_5338,N_5103);
and U5487 (N_5487,N_5337,N_5174);
xor U5488 (N_5488,N_5270,N_5170);
xor U5489 (N_5489,N_5278,N_5380);
or U5490 (N_5490,N_5382,N_5262);
nor U5491 (N_5491,N_5110,N_5101);
nor U5492 (N_5492,N_5120,N_5113);
nor U5493 (N_5493,N_5321,N_5374);
and U5494 (N_5494,N_5225,N_5139);
or U5495 (N_5495,N_5240,N_5158);
and U5496 (N_5496,N_5274,N_5172);
nor U5497 (N_5497,N_5334,N_5132);
xor U5498 (N_5498,N_5284,N_5271);
nand U5499 (N_5499,N_5184,N_5116);
xnor U5500 (N_5500,N_5388,N_5159);
or U5501 (N_5501,N_5126,N_5363);
or U5502 (N_5502,N_5183,N_5231);
or U5503 (N_5503,N_5297,N_5193);
nand U5504 (N_5504,N_5351,N_5175);
xor U5505 (N_5505,N_5308,N_5234);
or U5506 (N_5506,N_5221,N_5146);
nor U5507 (N_5507,N_5154,N_5230);
xnor U5508 (N_5508,N_5121,N_5149);
and U5509 (N_5509,N_5244,N_5138);
nand U5510 (N_5510,N_5364,N_5140);
or U5511 (N_5511,N_5176,N_5327);
or U5512 (N_5512,N_5142,N_5383);
and U5513 (N_5513,N_5279,N_5191);
nand U5514 (N_5514,N_5356,N_5131);
nand U5515 (N_5515,N_5112,N_5293);
or U5516 (N_5516,N_5135,N_5156);
and U5517 (N_5517,N_5211,N_5200);
nor U5518 (N_5518,N_5384,N_5350);
or U5519 (N_5519,N_5167,N_5169);
and U5520 (N_5520,N_5332,N_5263);
or U5521 (N_5521,N_5228,N_5397);
nor U5522 (N_5522,N_5329,N_5186);
xnor U5523 (N_5523,N_5257,N_5168);
nor U5524 (N_5524,N_5311,N_5150);
or U5525 (N_5525,N_5304,N_5144);
xor U5526 (N_5526,N_5340,N_5335);
nor U5527 (N_5527,N_5276,N_5336);
nor U5528 (N_5528,N_5180,N_5315);
nand U5529 (N_5529,N_5355,N_5214);
nand U5530 (N_5530,N_5133,N_5260);
nand U5531 (N_5531,N_5385,N_5352);
nand U5532 (N_5532,N_5393,N_5305);
or U5533 (N_5533,N_5301,N_5199);
nand U5534 (N_5534,N_5145,N_5141);
xor U5535 (N_5535,N_5370,N_5368);
nor U5536 (N_5536,N_5280,N_5195);
xnor U5537 (N_5537,N_5226,N_5130);
nor U5538 (N_5538,N_5205,N_5161);
or U5539 (N_5539,N_5202,N_5215);
and U5540 (N_5540,N_5320,N_5348);
and U5541 (N_5541,N_5236,N_5185);
nor U5542 (N_5542,N_5261,N_5273);
or U5543 (N_5543,N_5177,N_5201);
nand U5544 (N_5544,N_5354,N_5164);
nor U5545 (N_5545,N_5114,N_5326);
nand U5546 (N_5546,N_5394,N_5250);
or U5547 (N_5547,N_5166,N_5359);
nand U5548 (N_5548,N_5117,N_5252);
and U5549 (N_5549,N_5206,N_5213);
nand U5550 (N_5550,N_5159,N_5392);
xnor U5551 (N_5551,N_5230,N_5155);
or U5552 (N_5552,N_5219,N_5284);
and U5553 (N_5553,N_5102,N_5338);
xor U5554 (N_5554,N_5174,N_5124);
and U5555 (N_5555,N_5361,N_5377);
nand U5556 (N_5556,N_5186,N_5143);
nand U5557 (N_5557,N_5347,N_5107);
nand U5558 (N_5558,N_5133,N_5262);
xor U5559 (N_5559,N_5330,N_5243);
nand U5560 (N_5560,N_5180,N_5201);
nor U5561 (N_5561,N_5179,N_5172);
and U5562 (N_5562,N_5271,N_5179);
xor U5563 (N_5563,N_5369,N_5355);
and U5564 (N_5564,N_5328,N_5185);
and U5565 (N_5565,N_5271,N_5137);
and U5566 (N_5566,N_5246,N_5289);
and U5567 (N_5567,N_5166,N_5280);
nand U5568 (N_5568,N_5297,N_5118);
nor U5569 (N_5569,N_5241,N_5166);
nor U5570 (N_5570,N_5355,N_5111);
and U5571 (N_5571,N_5202,N_5153);
or U5572 (N_5572,N_5239,N_5138);
and U5573 (N_5573,N_5364,N_5213);
nand U5574 (N_5574,N_5332,N_5338);
and U5575 (N_5575,N_5146,N_5388);
xnor U5576 (N_5576,N_5247,N_5194);
and U5577 (N_5577,N_5273,N_5370);
xor U5578 (N_5578,N_5340,N_5285);
xnor U5579 (N_5579,N_5119,N_5190);
nor U5580 (N_5580,N_5210,N_5218);
nand U5581 (N_5581,N_5193,N_5234);
or U5582 (N_5582,N_5197,N_5227);
and U5583 (N_5583,N_5371,N_5111);
or U5584 (N_5584,N_5357,N_5388);
nor U5585 (N_5585,N_5204,N_5394);
nor U5586 (N_5586,N_5127,N_5178);
and U5587 (N_5587,N_5310,N_5221);
nand U5588 (N_5588,N_5397,N_5282);
and U5589 (N_5589,N_5150,N_5310);
nor U5590 (N_5590,N_5252,N_5159);
nor U5591 (N_5591,N_5187,N_5285);
xnor U5592 (N_5592,N_5250,N_5379);
nor U5593 (N_5593,N_5319,N_5279);
xor U5594 (N_5594,N_5235,N_5237);
xor U5595 (N_5595,N_5169,N_5136);
xnor U5596 (N_5596,N_5137,N_5206);
nand U5597 (N_5597,N_5371,N_5181);
nor U5598 (N_5598,N_5131,N_5102);
xor U5599 (N_5599,N_5100,N_5161);
or U5600 (N_5600,N_5219,N_5341);
or U5601 (N_5601,N_5162,N_5349);
nor U5602 (N_5602,N_5282,N_5213);
xnor U5603 (N_5603,N_5350,N_5371);
nor U5604 (N_5604,N_5231,N_5125);
and U5605 (N_5605,N_5206,N_5320);
and U5606 (N_5606,N_5262,N_5193);
nand U5607 (N_5607,N_5218,N_5291);
xor U5608 (N_5608,N_5272,N_5268);
or U5609 (N_5609,N_5384,N_5190);
or U5610 (N_5610,N_5383,N_5318);
xor U5611 (N_5611,N_5342,N_5240);
and U5612 (N_5612,N_5226,N_5390);
xor U5613 (N_5613,N_5325,N_5367);
nand U5614 (N_5614,N_5281,N_5183);
or U5615 (N_5615,N_5344,N_5323);
or U5616 (N_5616,N_5148,N_5210);
or U5617 (N_5617,N_5370,N_5183);
and U5618 (N_5618,N_5282,N_5204);
xnor U5619 (N_5619,N_5204,N_5264);
nand U5620 (N_5620,N_5144,N_5375);
or U5621 (N_5621,N_5114,N_5190);
nor U5622 (N_5622,N_5202,N_5389);
or U5623 (N_5623,N_5273,N_5293);
nand U5624 (N_5624,N_5145,N_5282);
nor U5625 (N_5625,N_5124,N_5276);
and U5626 (N_5626,N_5117,N_5217);
xnor U5627 (N_5627,N_5359,N_5384);
and U5628 (N_5628,N_5158,N_5145);
xor U5629 (N_5629,N_5192,N_5319);
and U5630 (N_5630,N_5336,N_5106);
xnor U5631 (N_5631,N_5129,N_5163);
xor U5632 (N_5632,N_5104,N_5195);
nand U5633 (N_5633,N_5113,N_5109);
and U5634 (N_5634,N_5329,N_5118);
xnor U5635 (N_5635,N_5143,N_5220);
or U5636 (N_5636,N_5393,N_5216);
nor U5637 (N_5637,N_5184,N_5306);
and U5638 (N_5638,N_5283,N_5253);
xor U5639 (N_5639,N_5122,N_5161);
and U5640 (N_5640,N_5374,N_5205);
nand U5641 (N_5641,N_5145,N_5378);
nand U5642 (N_5642,N_5285,N_5168);
nor U5643 (N_5643,N_5392,N_5146);
or U5644 (N_5644,N_5344,N_5147);
and U5645 (N_5645,N_5187,N_5199);
or U5646 (N_5646,N_5297,N_5130);
xnor U5647 (N_5647,N_5383,N_5387);
nor U5648 (N_5648,N_5237,N_5218);
xor U5649 (N_5649,N_5334,N_5194);
nor U5650 (N_5650,N_5167,N_5187);
and U5651 (N_5651,N_5387,N_5284);
xnor U5652 (N_5652,N_5290,N_5362);
xnor U5653 (N_5653,N_5273,N_5191);
nand U5654 (N_5654,N_5155,N_5378);
or U5655 (N_5655,N_5251,N_5149);
or U5656 (N_5656,N_5218,N_5200);
xor U5657 (N_5657,N_5385,N_5253);
or U5658 (N_5658,N_5286,N_5262);
nor U5659 (N_5659,N_5167,N_5193);
or U5660 (N_5660,N_5311,N_5375);
or U5661 (N_5661,N_5386,N_5249);
and U5662 (N_5662,N_5261,N_5380);
nor U5663 (N_5663,N_5120,N_5142);
xor U5664 (N_5664,N_5213,N_5390);
nand U5665 (N_5665,N_5398,N_5236);
or U5666 (N_5666,N_5256,N_5136);
or U5667 (N_5667,N_5338,N_5344);
nor U5668 (N_5668,N_5173,N_5380);
xor U5669 (N_5669,N_5281,N_5115);
nand U5670 (N_5670,N_5356,N_5335);
and U5671 (N_5671,N_5177,N_5202);
nor U5672 (N_5672,N_5191,N_5221);
or U5673 (N_5673,N_5108,N_5111);
nand U5674 (N_5674,N_5349,N_5287);
or U5675 (N_5675,N_5330,N_5159);
nor U5676 (N_5676,N_5328,N_5250);
xor U5677 (N_5677,N_5100,N_5129);
nand U5678 (N_5678,N_5238,N_5388);
nand U5679 (N_5679,N_5208,N_5290);
and U5680 (N_5680,N_5354,N_5205);
nand U5681 (N_5681,N_5158,N_5217);
nor U5682 (N_5682,N_5239,N_5379);
and U5683 (N_5683,N_5208,N_5194);
nor U5684 (N_5684,N_5351,N_5259);
nand U5685 (N_5685,N_5250,N_5197);
nand U5686 (N_5686,N_5173,N_5121);
or U5687 (N_5687,N_5282,N_5160);
or U5688 (N_5688,N_5274,N_5202);
nor U5689 (N_5689,N_5320,N_5132);
or U5690 (N_5690,N_5197,N_5375);
and U5691 (N_5691,N_5108,N_5271);
and U5692 (N_5692,N_5253,N_5243);
nand U5693 (N_5693,N_5131,N_5190);
or U5694 (N_5694,N_5341,N_5183);
and U5695 (N_5695,N_5297,N_5156);
and U5696 (N_5696,N_5281,N_5119);
and U5697 (N_5697,N_5161,N_5322);
and U5698 (N_5698,N_5315,N_5185);
xor U5699 (N_5699,N_5250,N_5382);
and U5700 (N_5700,N_5630,N_5414);
and U5701 (N_5701,N_5596,N_5470);
and U5702 (N_5702,N_5586,N_5618);
nand U5703 (N_5703,N_5475,N_5445);
xor U5704 (N_5704,N_5581,N_5554);
or U5705 (N_5705,N_5698,N_5535);
and U5706 (N_5706,N_5430,N_5562);
xnor U5707 (N_5707,N_5664,N_5432);
or U5708 (N_5708,N_5602,N_5478);
nand U5709 (N_5709,N_5457,N_5696);
or U5710 (N_5710,N_5648,N_5532);
or U5711 (N_5711,N_5427,N_5472);
or U5712 (N_5712,N_5420,N_5659);
and U5713 (N_5713,N_5443,N_5568);
or U5714 (N_5714,N_5452,N_5636);
or U5715 (N_5715,N_5540,N_5592);
or U5716 (N_5716,N_5514,N_5507);
and U5717 (N_5717,N_5474,N_5661);
nor U5718 (N_5718,N_5519,N_5464);
or U5719 (N_5719,N_5666,N_5667);
xnor U5720 (N_5720,N_5597,N_5440);
xnor U5721 (N_5721,N_5439,N_5675);
or U5722 (N_5722,N_5516,N_5660);
and U5723 (N_5723,N_5561,N_5504);
nor U5724 (N_5724,N_5520,N_5541);
nor U5725 (N_5725,N_5578,N_5418);
or U5726 (N_5726,N_5685,N_5694);
nand U5727 (N_5727,N_5406,N_5575);
nor U5728 (N_5728,N_5650,N_5487);
nand U5729 (N_5729,N_5591,N_5436);
or U5730 (N_5730,N_5460,N_5466);
or U5731 (N_5731,N_5484,N_5405);
nand U5732 (N_5732,N_5428,N_5515);
nand U5733 (N_5733,N_5601,N_5438);
nor U5734 (N_5734,N_5673,N_5480);
or U5735 (N_5735,N_5419,N_5616);
and U5736 (N_5736,N_5593,N_5530);
nand U5737 (N_5737,N_5552,N_5412);
nor U5738 (N_5738,N_5579,N_5517);
nand U5739 (N_5739,N_5435,N_5413);
or U5740 (N_5740,N_5672,N_5501);
nand U5741 (N_5741,N_5537,N_5640);
nand U5742 (N_5742,N_5658,N_5547);
or U5743 (N_5743,N_5546,N_5599);
nor U5744 (N_5744,N_5437,N_5479);
nor U5745 (N_5745,N_5434,N_5500);
nor U5746 (N_5746,N_5495,N_5674);
and U5747 (N_5747,N_5473,N_5585);
or U5748 (N_5748,N_5598,N_5615);
or U5749 (N_5749,N_5691,N_5449);
or U5750 (N_5750,N_5619,N_5584);
xor U5751 (N_5751,N_5506,N_5489);
xor U5752 (N_5752,N_5624,N_5447);
nand U5753 (N_5753,N_5638,N_5695);
or U5754 (N_5754,N_5555,N_5632);
or U5755 (N_5755,N_5662,N_5684);
nor U5756 (N_5756,N_5682,N_5563);
nand U5757 (N_5757,N_5483,N_5402);
and U5758 (N_5758,N_5426,N_5494);
or U5759 (N_5759,N_5521,N_5486);
or U5760 (N_5760,N_5642,N_5560);
and U5761 (N_5761,N_5522,N_5551);
and U5762 (N_5762,N_5543,N_5463);
and U5763 (N_5763,N_5643,N_5482);
nor U5764 (N_5764,N_5416,N_5572);
nand U5765 (N_5765,N_5548,N_5512);
nor U5766 (N_5766,N_5467,N_5611);
or U5767 (N_5767,N_5655,N_5454);
nor U5768 (N_5768,N_5654,N_5692);
nand U5769 (N_5769,N_5431,N_5421);
nor U5770 (N_5770,N_5580,N_5549);
xor U5771 (N_5771,N_5669,N_5534);
nand U5772 (N_5772,N_5577,N_5441);
nand U5773 (N_5773,N_5641,N_5451);
nand U5774 (N_5774,N_5417,N_5678);
xor U5775 (N_5775,N_5576,N_5647);
nand U5776 (N_5776,N_5453,N_5404);
nor U5777 (N_5777,N_5415,N_5566);
nor U5778 (N_5778,N_5651,N_5536);
or U5779 (N_5779,N_5608,N_5653);
nand U5780 (N_5780,N_5595,N_5565);
nor U5781 (N_5781,N_5528,N_5679);
or U5782 (N_5782,N_5485,N_5557);
nor U5783 (N_5783,N_5491,N_5607);
and U5784 (N_5784,N_5677,N_5690);
xnor U5785 (N_5785,N_5687,N_5539);
or U5786 (N_5786,N_5542,N_5433);
or U5787 (N_5787,N_5456,N_5649);
and U5788 (N_5788,N_5644,N_5498);
or U5789 (N_5789,N_5424,N_5681);
nand U5790 (N_5790,N_5505,N_5408);
and U5791 (N_5791,N_5490,N_5465);
nand U5792 (N_5792,N_5497,N_5538);
and U5793 (N_5793,N_5623,N_5627);
and U5794 (N_5794,N_5468,N_5610);
nor U5795 (N_5795,N_5697,N_5544);
and U5796 (N_5796,N_5583,N_5587);
or U5797 (N_5797,N_5633,N_5693);
nor U5798 (N_5798,N_5604,N_5469);
and U5799 (N_5799,N_5476,N_5683);
nand U5800 (N_5800,N_5526,N_5639);
nor U5801 (N_5801,N_5422,N_5503);
nor U5802 (N_5802,N_5511,N_5645);
xor U5803 (N_5803,N_5410,N_5558);
xnor U5804 (N_5804,N_5588,N_5612);
nand U5805 (N_5805,N_5545,N_5510);
nor U5806 (N_5806,N_5411,N_5509);
and U5807 (N_5807,N_5614,N_5429);
or U5808 (N_5808,N_5670,N_5499);
nand U5809 (N_5809,N_5525,N_5622);
nand U5810 (N_5810,N_5613,N_5448);
and U5811 (N_5811,N_5527,N_5589);
nand U5812 (N_5812,N_5609,N_5524);
and U5813 (N_5813,N_5553,N_5686);
nor U5814 (N_5814,N_5400,N_5533);
and U5815 (N_5815,N_5458,N_5699);
and U5816 (N_5816,N_5564,N_5481);
and U5817 (N_5817,N_5676,N_5657);
nor U5818 (N_5818,N_5573,N_5455);
nand U5819 (N_5819,N_5603,N_5600);
xnor U5820 (N_5820,N_5409,N_5531);
nor U5821 (N_5821,N_5444,N_5594);
or U5822 (N_5822,N_5621,N_5629);
nand U5823 (N_5823,N_5571,N_5628);
or U5824 (N_5824,N_5462,N_5574);
and U5825 (N_5825,N_5656,N_5635);
nand U5826 (N_5826,N_5620,N_5668);
or U5827 (N_5827,N_5446,N_5634);
nand U5828 (N_5828,N_5529,N_5423);
or U5829 (N_5829,N_5582,N_5442);
nand U5830 (N_5830,N_5570,N_5663);
nand U5831 (N_5831,N_5496,N_5605);
or U5832 (N_5832,N_5477,N_5488);
xnor U5833 (N_5833,N_5646,N_5407);
nor U5834 (N_5834,N_5626,N_5567);
and U5835 (N_5835,N_5403,N_5606);
xor U5836 (N_5836,N_5556,N_5401);
or U5837 (N_5837,N_5523,N_5459);
nor U5838 (N_5838,N_5689,N_5508);
xnor U5839 (N_5839,N_5559,N_5569);
nand U5840 (N_5840,N_5471,N_5631);
nand U5841 (N_5841,N_5665,N_5637);
nand U5842 (N_5842,N_5518,N_5590);
xor U5843 (N_5843,N_5671,N_5492);
or U5844 (N_5844,N_5625,N_5450);
and U5845 (N_5845,N_5652,N_5688);
nand U5846 (N_5846,N_5425,N_5493);
nand U5847 (N_5847,N_5617,N_5502);
and U5848 (N_5848,N_5550,N_5513);
or U5849 (N_5849,N_5680,N_5461);
nand U5850 (N_5850,N_5624,N_5465);
and U5851 (N_5851,N_5595,N_5594);
xnor U5852 (N_5852,N_5449,N_5408);
and U5853 (N_5853,N_5417,N_5502);
nor U5854 (N_5854,N_5631,N_5402);
nor U5855 (N_5855,N_5698,N_5494);
xnor U5856 (N_5856,N_5519,N_5494);
nor U5857 (N_5857,N_5541,N_5675);
nand U5858 (N_5858,N_5527,N_5445);
or U5859 (N_5859,N_5512,N_5436);
xnor U5860 (N_5860,N_5675,N_5475);
nor U5861 (N_5861,N_5449,N_5498);
or U5862 (N_5862,N_5549,N_5656);
and U5863 (N_5863,N_5579,N_5538);
nor U5864 (N_5864,N_5531,N_5683);
nand U5865 (N_5865,N_5463,N_5560);
nor U5866 (N_5866,N_5446,N_5463);
nor U5867 (N_5867,N_5693,N_5492);
nor U5868 (N_5868,N_5522,N_5654);
nand U5869 (N_5869,N_5614,N_5470);
nor U5870 (N_5870,N_5699,N_5663);
xnor U5871 (N_5871,N_5654,N_5637);
and U5872 (N_5872,N_5592,N_5683);
nor U5873 (N_5873,N_5684,N_5494);
nor U5874 (N_5874,N_5590,N_5544);
xnor U5875 (N_5875,N_5696,N_5417);
xor U5876 (N_5876,N_5676,N_5546);
and U5877 (N_5877,N_5676,N_5493);
nand U5878 (N_5878,N_5580,N_5472);
xor U5879 (N_5879,N_5591,N_5471);
or U5880 (N_5880,N_5653,N_5582);
nor U5881 (N_5881,N_5495,N_5623);
nor U5882 (N_5882,N_5494,N_5606);
xnor U5883 (N_5883,N_5436,N_5534);
and U5884 (N_5884,N_5696,N_5615);
nor U5885 (N_5885,N_5691,N_5425);
and U5886 (N_5886,N_5597,N_5478);
nor U5887 (N_5887,N_5449,N_5456);
and U5888 (N_5888,N_5411,N_5467);
nor U5889 (N_5889,N_5454,N_5684);
or U5890 (N_5890,N_5411,N_5548);
nand U5891 (N_5891,N_5564,N_5407);
and U5892 (N_5892,N_5443,N_5636);
and U5893 (N_5893,N_5581,N_5681);
or U5894 (N_5894,N_5527,N_5432);
and U5895 (N_5895,N_5557,N_5436);
nor U5896 (N_5896,N_5631,N_5587);
nand U5897 (N_5897,N_5647,N_5609);
nor U5898 (N_5898,N_5444,N_5656);
nor U5899 (N_5899,N_5668,N_5496);
xor U5900 (N_5900,N_5409,N_5532);
and U5901 (N_5901,N_5403,N_5565);
and U5902 (N_5902,N_5417,N_5650);
nand U5903 (N_5903,N_5518,N_5636);
and U5904 (N_5904,N_5634,N_5500);
or U5905 (N_5905,N_5584,N_5410);
or U5906 (N_5906,N_5657,N_5425);
nor U5907 (N_5907,N_5459,N_5660);
and U5908 (N_5908,N_5587,N_5622);
or U5909 (N_5909,N_5648,N_5551);
and U5910 (N_5910,N_5628,N_5473);
nand U5911 (N_5911,N_5472,N_5561);
or U5912 (N_5912,N_5692,N_5403);
and U5913 (N_5913,N_5531,N_5652);
nor U5914 (N_5914,N_5672,N_5509);
or U5915 (N_5915,N_5599,N_5418);
nand U5916 (N_5916,N_5407,N_5563);
xor U5917 (N_5917,N_5661,N_5455);
nor U5918 (N_5918,N_5695,N_5529);
nand U5919 (N_5919,N_5431,N_5668);
or U5920 (N_5920,N_5449,N_5669);
nand U5921 (N_5921,N_5540,N_5651);
or U5922 (N_5922,N_5405,N_5516);
or U5923 (N_5923,N_5546,N_5470);
or U5924 (N_5924,N_5527,N_5639);
xnor U5925 (N_5925,N_5693,N_5515);
nor U5926 (N_5926,N_5639,N_5480);
or U5927 (N_5927,N_5444,N_5639);
nor U5928 (N_5928,N_5419,N_5639);
nand U5929 (N_5929,N_5574,N_5448);
and U5930 (N_5930,N_5681,N_5695);
and U5931 (N_5931,N_5634,N_5463);
or U5932 (N_5932,N_5417,N_5508);
and U5933 (N_5933,N_5446,N_5494);
xor U5934 (N_5934,N_5446,N_5626);
nand U5935 (N_5935,N_5457,N_5435);
nor U5936 (N_5936,N_5540,N_5578);
nor U5937 (N_5937,N_5491,N_5424);
xor U5938 (N_5938,N_5594,N_5403);
xor U5939 (N_5939,N_5457,N_5487);
xnor U5940 (N_5940,N_5581,N_5682);
nor U5941 (N_5941,N_5505,N_5413);
and U5942 (N_5942,N_5494,N_5670);
nand U5943 (N_5943,N_5679,N_5667);
nor U5944 (N_5944,N_5680,N_5594);
or U5945 (N_5945,N_5585,N_5440);
xor U5946 (N_5946,N_5579,N_5440);
nor U5947 (N_5947,N_5636,N_5431);
nand U5948 (N_5948,N_5633,N_5650);
or U5949 (N_5949,N_5672,N_5641);
nor U5950 (N_5950,N_5637,N_5412);
nor U5951 (N_5951,N_5421,N_5417);
nand U5952 (N_5952,N_5411,N_5451);
or U5953 (N_5953,N_5552,N_5635);
xor U5954 (N_5954,N_5445,N_5616);
or U5955 (N_5955,N_5663,N_5650);
nor U5956 (N_5956,N_5610,N_5440);
and U5957 (N_5957,N_5637,N_5594);
xor U5958 (N_5958,N_5673,N_5505);
xor U5959 (N_5959,N_5484,N_5602);
or U5960 (N_5960,N_5499,N_5422);
nor U5961 (N_5961,N_5534,N_5575);
nand U5962 (N_5962,N_5469,N_5628);
and U5963 (N_5963,N_5538,N_5429);
or U5964 (N_5964,N_5604,N_5635);
xor U5965 (N_5965,N_5449,N_5515);
or U5966 (N_5966,N_5588,N_5666);
or U5967 (N_5967,N_5401,N_5607);
nor U5968 (N_5968,N_5480,N_5643);
nand U5969 (N_5969,N_5660,N_5564);
xor U5970 (N_5970,N_5590,N_5565);
or U5971 (N_5971,N_5467,N_5691);
or U5972 (N_5972,N_5451,N_5672);
nor U5973 (N_5973,N_5458,N_5559);
and U5974 (N_5974,N_5631,N_5409);
nand U5975 (N_5975,N_5640,N_5637);
or U5976 (N_5976,N_5437,N_5529);
nor U5977 (N_5977,N_5414,N_5601);
xnor U5978 (N_5978,N_5431,N_5635);
nand U5979 (N_5979,N_5468,N_5572);
nand U5980 (N_5980,N_5686,N_5514);
or U5981 (N_5981,N_5603,N_5508);
or U5982 (N_5982,N_5557,N_5456);
nand U5983 (N_5983,N_5621,N_5667);
and U5984 (N_5984,N_5612,N_5486);
nand U5985 (N_5985,N_5558,N_5652);
or U5986 (N_5986,N_5523,N_5529);
xnor U5987 (N_5987,N_5533,N_5530);
and U5988 (N_5988,N_5555,N_5576);
xnor U5989 (N_5989,N_5674,N_5554);
xnor U5990 (N_5990,N_5588,N_5490);
nand U5991 (N_5991,N_5596,N_5639);
nand U5992 (N_5992,N_5623,N_5648);
nand U5993 (N_5993,N_5689,N_5680);
xor U5994 (N_5994,N_5512,N_5472);
and U5995 (N_5995,N_5586,N_5612);
or U5996 (N_5996,N_5424,N_5628);
nand U5997 (N_5997,N_5404,N_5427);
xor U5998 (N_5998,N_5560,N_5419);
nor U5999 (N_5999,N_5614,N_5643);
and U6000 (N_6000,N_5918,N_5922);
nor U6001 (N_6001,N_5977,N_5897);
nand U6002 (N_6002,N_5967,N_5966);
nor U6003 (N_6003,N_5742,N_5731);
and U6004 (N_6004,N_5991,N_5733);
and U6005 (N_6005,N_5750,N_5871);
or U6006 (N_6006,N_5719,N_5724);
nor U6007 (N_6007,N_5870,N_5956);
nand U6008 (N_6008,N_5976,N_5803);
or U6009 (N_6009,N_5720,N_5853);
or U6010 (N_6010,N_5906,N_5844);
and U6011 (N_6011,N_5867,N_5846);
xor U6012 (N_6012,N_5718,N_5944);
or U6013 (N_6013,N_5707,N_5861);
nor U6014 (N_6014,N_5789,N_5962);
or U6015 (N_6015,N_5968,N_5911);
or U6016 (N_6016,N_5704,N_5822);
nand U6017 (N_6017,N_5912,N_5886);
and U6018 (N_6018,N_5910,N_5808);
nor U6019 (N_6019,N_5751,N_5814);
nor U6020 (N_6020,N_5957,N_5998);
nor U6021 (N_6021,N_5915,N_5896);
nand U6022 (N_6022,N_5916,N_5826);
xor U6023 (N_6023,N_5869,N_5811);
nor U6024 (N_6024,N_5828,N_5947);
nor U6025 (N_6025,N_5908,N_5820);
or U6026 (N_6026,N_5900,N_5904);
xnor U6027 (N_6027,N_5955,N_5999);
and U6028 (N_6028,N_5934,N_5804);
and U6029 (N_6029,N_5798,N_5935);
nand U6030 (N_6030,N_5990,N_5891);
nand U6031 (N_6031,N_5772,N_5949);
nand U6032 (N_6032,N_5730,N_5920);
nor U6033 (N_6033,N_5997,N_5945);
nand U6034 (N_6034,N_5973,N_5903);
xnor U6035 (N_6035,N_5709,N_5778);
and U6036 (N_6036,N_5787,N_5817);
or U6037 (N_6037,N_5954,N_5721);
or U6038 (N_6038,N_5777,N_5836);
and U6039 (N_6039,N_5866,N_5980);
or U6040 (N_6040,N_5734,N_5879);
and U6041 (N_6041,N_5760,N_5880);
nand U6042 (N_6042,N_5986,N_5741);
and U6043 (N_6043,N_5958,N_5799);
nor U6044 (N_6044,N_5702,N_5763);
xor U6045 (N_6045,N_5797,N_5847);
nor U6046 (N_6046,N_5882,N_5941);
nor U6047 (N_6047,N_5907,N_5842);
and U6048 (N_6048,N_5786,N_5802);
nand U6049 (N_6049,N_5984,N_5963);
nand U6050 (N_6050,N_5863,N_5744);
xor U6051 (N_6051,N_5788,N_5855);
nand U6052 (N_6052,N_5746,N_5703);
nand U6053 (N_6053,N_5736,N_5767);
nand U6054 (N_6054,N_5994,N_5848);
and U6055 (N_6055,N_5969,N_5748);
nor U6056 (N_6056,N_5978,N_5854);
nand U6057 (N_6057,N_5840,N_5735);
or U6058 (N_6058,N_5876,N_5726);
or U6059 (N_6059,N_5852,N_5987);
and U6060 (N_6060,N_5776,N_5856);
nand U6061 (N_6061,N_5883,N_5830);
nand U6062 (N_6062,N_5850,N_5711);
xnor U6063 (N_6063,N_5796,N_5961);
xnor U6064 (N_6064,N_5924,N_5933);
or U6065 (N_6065,N_5706,N_5914);
nand U6066 (N_6066,N_5759,N_5909);
nor U6067 (N_6067,N_5927,N_5985);
and U6068 (N_6068,N_5732,N_5747);
nor U6069 (N_6069,N_5737,N_5781);
nand U6070 (N_6070,N_5783,N_5884);
nor U6071 (N_6071,N_5743,N_5723);
and U6072 (N_6072,N_5715,N_5810);
or U6073 (N_6073,N_5766,N_5975);
nor U6074 (N_6074,N_5819,N_5764);
or U6075 (N_6075,N_5902,N_5843);
nand U6076 (N_6076,N_5972,N_5713);
or U6077 (N_6077,N_5943,N_5923);
xnor U6078 (N_6078,N_5995,N_5881);
or U6079 (N_6079,N_5889,N_5717);
or U6080 (N_6080,N_5888,N_5942);
xnor U6081 (N_6081,N_5812,N_5992);
or U6082 (N_6082,N_5989,N_5762);
nor U6083 (N_6083,N_5859,N_5809);
nor U6084 (N_6084,N_5917,N_5971);
nor U6085 (N_6085,N_5834,N_5940);
and U6086 (N_6086,N_5710,N_5708);
and U6087 (N_6087,N_5983,N_5919);
xor U6088 (N_6088,N_5701,N_5851);
nor U6089 (N_6089,N_5700,N_5825);
nor U6090 (N_6090,N_5754,N_5800);
nand U6091 (N_6091,N_5905,N_5928);
or U6092 (N_6092,N_5784,N_5761);
and U6093 (N_6093,N_5832,N_5785);
nor U6094 (N_6094,N_5752,N_5727);
or U6095 (N_6095,N_5815,N_5716);
or U6096 (N_6096,N_5929,N_5779);
nand U6097 (N_6097,N_5837,N_5890);
nand U6098 (N_6098,N_5827,N_5770);
nor U6099 (N_6099,N_5887,N_5818);
or U6100 (N_6100,N_5996,N_5873);
or U6101 (N_6101,N_5892,N_5950);
xnor U6102 (N_6102,N_5790,N_5993);
xor U6103 (N_6103,N_5862,N_5740);
xor U6104 (N_6104,N_5801,N_5839);
nand U6105 (N_6105,N_5807,N_5959);
and U6106 (N_6106,N_5858,N_5951);
nor U6107 (N_6107,N_5757,N_5821);
nand U6108 (N_6108,N_5782,N_5816);
and U6109 (N_6109,N_5868,N_5780);
nand U6110 (N_6110,N_5965,N_5775);
xnor U6111 (N_6111,N_5712,N_5813);
and U6112 (N_6112,N_5758,N_5833);
xor U6113 (N_6113,N_5749,N_5974);
nor U6114 (N_6114,N_5936,N_5913);
nor U6115 (N_6115,N_5878,N_5769);
xor U6116 (N_6116,N_5792,N_5921);
or U6117 (N_6117,N_5795,N_5857);
xnor U6118 (N_6118,N_5806,N_5714);
nand U6119 (N_6119,N_5948,N_5753);
nor U6120 (N_6120,N_5960,N_5895);
nand U6121 (N_6121,N_5841,N_5885);
and U6122 (N_6122,N_5952,N_5953);
nand U6123 (N_6123,N_5745,N_5771);
or U6124 (N_6124,N_5937,N_5925);
nand U6125 (N_6125,N_5793,N_5926);
nor U6126 (N_6126,N_5875,N_5901);
nor U6127 (N_6127,N_5930,N_5725);
nor U6128 (N_6128,N_5738,N_5823);
nand U6129 (N_6129,N_5794,N_5835);
xnor U6130 (N_6130,N_5877,N_5774);
nor U6131 (N_6131,N_5729,N_5893);
and U6132 (N_6132,N_5860,N_5939);
or U6133 (N_6133,N_5845,N_5755);
and U6134 (N_6134,N_5831,N_5982);
xor U6135 (N_6135,N_5898,N_5946);
and U6136 (N_6136,N_5931,N_5938);
and U6137 (N_6137,N_5894,N_5849);
xnor U6138 (N_6138,N_5739,N_5768);
or U6139 (N_6139,N_5864,N_5872);
and U6140 (N_6140,N_5964,N_5970);
xnor U6141 (N_6141,N_5981,N_5865);
and U6142 (N_6142,N_5722,N_5874);
or U6143 (N_6143,N_5805,N_5932);
nand U6144 (N_6144,N_5791,N_5829);
xor U6145 (N_6145,N_5988,N_5838);
and U6146 (N_6146,N_5824,N_5705);
nand U6147 (N_6147,N_5979,N_5765);
or U6148 (N_6148,N_5773,N_5756);
nor U6149 (N_6149,N_5728,N_5899);
nand U6150 (N_6150,N_5895,N_5834);
xor U6151 (N_6151,N_5933,N_5706);
nor U6152 (N_6152,N_5963,N_5937);
xnor U6153 (N_6153,N_5924,N_5726);
nor U6154 (N_6154,N_5730,N_5831);
and U6155 (N_6155,N_5845,N_5992);
xor U6156 (N_6156,N_5893,N_5916);
xnor U6157 (N_6157,N_5978,N_5796);
xor U6158 (N_6158,N_5910,N_5921);
nor U6159 (N_6159,N_5875,N_5914);
and U6160 (N_6160,N_5877,N_5727);
nand U6161 (N_6161,N_5703,N_5858);
nand U6162 (N_6162,N_5965,N_5905);
xnor U6163 (N_6163,N_5734,N_5766);
or U6164 (N_6164,N_5919,N_5777);
xnor U6165 (N_6165,N_5803,N_5998);
nand U6166 (N_6166,N_5772,N_5757);
xor U6167 (N_6167,N_5833,N_5829);
xor U6168 (N_6168,N_5927,N_5945);
xnor U6169 (N_6169,N_5943,N_5973);
or U6170 (N_6170,N_5766,N_5982);
or U6171 (N_6171,N_5794,N_5743);
nand U6172 (N_6172,N_5761,N_5771);
nand U6173 (N_6173,N_5718,N_5787);
xnor U6174 (N_6174,N_5896,N_5729);
nand U6175 (N_6175,N_5920,N_5996);
xor U6176 (N_6176,N_5963,N_5749);
and U6177 (N_6177,N_5921,N_5712);
xnor U6178 (N_6178,N_5807,N_5914);
xor U6179 (N_6179,N_5815,N_5802);
or U6180 (N_6180,N_5990,N_5974);
nand U6181 (N_6181,N_5825,N_5910);
nor U6182 (N_6182,N_5779,N_5776);
xnor U6183 (N_6183,N_5958,N_5899);
xor U6184 (N_6184,N_5815,N_5705);
or U6185 (N_6185,N_5970,N_5855);
and U6186 (N_6186,N_5730,N_5781);
nand U6187 (N_6187,N_5939,N_5914);
or U6188 (N_6188,N_5704,N_5943);
nor U6189 (N_6189,N_5907,N_5823);
and U6190 (N_6190,N_5883,N_5863);
or U6191 (N_6191,N_5950,N_5807);
or U6192 (N_6192,N_5771,N_5982);
nand U6193 (N_6193,N_5897,N_5898);
or U6194 (N_6194,N_5914,N_5987);
nand U6195 (N_6195,N_5820,N_5994);
xnor U6196 (N_6196,N_5951,N_5796);
nor U6197 (N_6197,N_5926,N_5835);
and U6198 (N_6198,N_5848,N_5839);
nor U6199 (N_6199,N_5829,N_5742);
or U6200 (N_6200,N_5830,N_5832);
or U6201 (N_6201,N_5867,N_5925);
nor U6202 (N_6202,N_5963,N_5924);
and U6203 (N_6203,N_5884,N_5709);
nor U6204 (N_6204,N_5859,N_5944);
nand U6205 (N_6205,N_5982,N_5980);
nand U6206 (N_6206,N_5993,N_5729);
xnor U6207 (N_6207,N_5768,N_5810);
and U6208 (N_6208,N_5895,N_5757);
or U6209 (N_6209,N_5973,N_5832);
nand U6210 (N_6210,N_5939,N_5984);
nor U6211 (N_6211,N_5710,N_5954);
or U6212 (N_6212,N_5727,N_5821);
and U6213 (N_6213,N_5968,N_5945);
nand U6214 (N_6214,N_5863,N_5920);
xor U6215 (N_6215,N_5732,N_5750);
or U6216 (N_6216,N_5972,N_5848);
and U6217 (N_6217,N_5715,N_5990);
or U6218 (N_6218,N_5810,N_5970);
or U6219 (N_6219,N_5950,N_5840);
or U6220 (N_6220,N_5817,N_5960);
and U6221 (N_6221,N_5964,N_5840);
xor U6222 (N_6222,N_5909,N_5756);
and U6223 (N_6223,N_5913,N_5766);
or U6224 (N_6224,N_5887,N_5917);
nand U6225 (N_6225,N_5731,N_5779);
or U6226 (N_6226,N_5882,N_5997);
xor U6227 (N_6227,N_5881,N_5797);
and U6228 (N_6228,N_5713,N_5719);
or U6229 (N_6229,N_5858,N_5929);
nand U6230 (N_6230,N_5767,N_5785);
nor U6231 (N_6231,N_5753,N_5852);
and U6232 (N_6232,N_5790,N_5912);
nor U6233 (N_6233,N_5800,N_5958);
nand U6234 (N_6234,N_5769,N_5750);
xnor U6235 (N_6235,N_5971,N_5718);
or U6236 (N_6236,N_5864,N_5910);
and U6237 (N_6237,N_5785,N_5995);
or U6238 (N_6238,N_5746,N_5766);
nand U6239 (N_6239,N_5864,N_5891);
nand U6240 (N_6240,N_5841,N_5809);
and U6241 (N_6241,N_5977,N_5735);
xnor U6242 (N_6242,N_5820,N_5783);
nand U6243 (N_6243,N_5999,N_5943);
xor U6244 (N_6244,N_5931,N_5926);
and U6245 (N_6245,N_5901,N_5947);
xor U6246 (N_6246,N_5829,N_5949);
nand U6247 (N_6247,N_5847,N_5796);
xnor U6248 (N_6248,N_5940,N_5944);
or U6249 (N_6249,N_5818,N_5717);
or U6250 (N_6250,N_5798,N_5976);
nor U6251 (N_6251,N_5979,N_5764);
xor U6252 (N_6252,N_5939,N_5988);
and U6253 (N_6253,N_5959,N_5732);
nor U6254 (N_6254,N_5905,N_5948);
nor U6255 (N_6255,N_5720,N_5791);
nor U6256 (N_6256,N_5963,N_5753);
xor U6257 (N_6257,N_5848,N_5822);
xor U6258 (N_6258,N_5973,N_5960);
and U6259 (N_6259,N_5996,N_5830);
or U6260 (N_6260,N_5801,N_5758);
and U6261 (N_6261,N_5806,N_5798);
nand U6262 (N_6262,N_5836,N_5733);
nor U6263 (N_6263,N_5727,N_5950);
xnor U6264 (N_6264,N_5864,N_5814);
and U6265 (N_6265,N_5735,N_5839);
nand U6266 (N_6266,N_5836,N_5839);
or U6267 (N_6267,N_5973,N_5947);
and U6268 (N_6268,N_5872,N_5855);
nor U6269 (N_6269,N_5859,N_5946);
and U6270 (N_6270,N_5720,N_5926);
or U6271 (N_6271,N_5757,N_5867);
nand U6272 (N_6272,N_5808,N_5866);
or U6273 (N_6273,N_5956,N_5907);
nor U6274 (N_6274,N_5763,N_5736);
nand U6275 (N_6275,N_5852,N_5829);
nand U6276 (N_6276,N_5701,N_5792);
xnor U6277 (N_6277,N_5762,N_5963);
or U6278 (N_6278,N_5806,N_5744);
xnor U6279 (N_6279,N_5740,N_5720);
and U6280 (N_6280,N_5759,N_5745);
nor U6281 (N_6281,N_5952,N_5809);
nand U6282 (N_6282,N_5713,N_5773);
nor U6283 (N_6283,N_5995,N_5904);
xnor U6284 (N_6284,N_5903,N_5950);
and U6285 (N_6285,N_5934,N_5852);
nand U6286 (N_6286,N_5708,N_5936);
and U6287 (N_6287,N_5708,N_5867);
or U6288 (N_6288,N_5778,N_5956);
xor U6289 (N_6289,N_5705,N_5769);
and U6290 (N_6290,N_5878,N_5822);
xnor U6291 (N_6291,N_5863,N_5970);
xnor U6292 (N_6292,N_5895,N_5940);
and U6293 (N_6293,N_5777,N_5956);
nor U6294 (N_6294,N_5740,N_5902);
nor U6295 (N_6295,N_5735,N_5954);
xor U6296 (N_6296,N_5846,N_5939);
or U6297 (N_6297,N_5712,N_5909);
and U6298 (N_6298,N_5916,N_5926);
xor U6299 (N_6299,N_5917,N_5773);
nand U6300 (N_6300,N_6236,N_6271);
nand U6301 (N_6301,N_6109,N_6280);
nor U6302 (N_6302,N_6063,N_6249);
xnor U6303 (N_6303,N_6047,N_6279);
xor U6304 (N_6304,N_6146,N_6031);
or U6305 (N_6305,N_6144,N_6173);
nor U6306 (N_6306,N_6209,N_6093);
or U6307 (N_6307,N_6233,N_6101);
xnor U6308 (N_6308,N_6006,N_6065);
nor U6309 (N_6309,N_6077,N_6054);
or U6310 (N_6310,N_6180,N_6166);
xor U6311 (N_6311,N_6184,N_6020);
nand U6312 (N_6312,N_6099,N_6203);
xor U6313 (N_6313,N_6238,N_6145);
or U6314 (N_6314,N_6068,N_6148);
and U6315 (N_6315,N_6055,N_6149);
nor U6316 (N_6316,N_6086,N_6032);
nand U6317 (N_6317,N_6285,N_6001);
xor U6318 (N_6318,N_6261,N_6197);
nand U6319 (N_6319,N_6222,N_6038);
and U6320 (N_6320,N_6226,N_6023);
nand U6321 (N_6321,N_6100,N_6151);
nor U6322 (N_6322,N_6064,N_6143);
nand U6323 (N_6323,N_6281,N_6025);
nand U6324 (N_6324,N_6157,N_6074);
and U6325 (N_6325,N_6177,N_6220);
or U6326 (N_6326,N_6187,N_6258);
nand U6327 (N_6327,N_6162,N_6019);
xor U6328 (N_6328,N_6161,N_6034);
xor U6329 (N_6329,N_6275,N_6026);
nor U6330 (N_6330,N_6277,N_6259);
and U6331 (N_6331,N_6194,N_6278);
or U6332 (N_6332,N_6282,N_6060);
or U6333 (N_6333,N_6231,N_6293);
nand U6334 (N_6334,N_6090,N_6147);
xor U6335 (N_6335,N_6015,N_6295);
nor U6336 (N_6336,N_6056,N_6070);
and U6337 (N_6337,N_6171,N_6036);
or U6338 (N_6338,N_6136,N_6043);
nand U6339 (N_6339,N_6132,N_6103);
nor U6340 (N_6340,N_6199,N_6287);
xor U6341 (N_6341,N_6224,N_6154);
or U6342 (N_6342,N_6097,N_6254);
nor U6343 (N_6343,N_6170,N_6181);
xor U6344 (N_6344,N_6114,N_6130);
or U6345 (N_6345,N_6215,N_6158);
xor U6346 (N_6346,N_6299,N_6021);
nand U6347 (N_6347,N_6073,N_6276);
nor U6348 (N_6348,N_6094,N_6269);
or U6349 (N_6349,N_6118,N_6010);
nand U6350 (N_6350,N_6007,N_6121);
nand U6351 (N_6351,N_6018,N_6104);
nand U6352 (N_6352,N_6189,N_6223);
nand U6353 (N_6353,N_6046,N_6242);
xor U6354 (N_6354,N_6075,N_6252);
nand U6355 (N_6355,N_6084,N_6240);
xor U6356 (N_6356,N_6204,N_6017);
nor U6357 (N_6357,N_6079,N_6198);
nor U6358 (N_6358,N_6035,N_6080);
nor U6359 (N_6359,N_6078,N_6012);
xnor U6360 (N_6360,N_6102,N_6013);
xor U6361 (N_6361,N_6057,N_6095);
nand U6362 (N_6362,N_6241,N_6156);
nor U6363 (N_6363,N_6243,N_6152);
xor U6364 (N_6364,N_6288,N_6098);
nand U6365 (N_6365,N_6011,N_6027);
and U6366 (N_6366,N_6126,N_6244);
xnor U6367 (N_6367,N_6133,N_6140);
xor U6368 (N_6368,N_6196,N_6218);
and U6369 (N_6369,N_6270,N_6256);
nand U6370 (N_6370,N_6228,N_6273);
xnor U6371 (N_6371,N_6155,N_6202);
xor U6372 (N_6372,N_6264,N_6045);
nor U6373 (N_6373,N_6206,N_6009);
and U6374 (N_6374,N_6205,N_6120);
or U6375 (N_6375,N_6213,N_6179);
nand U6376 (N_6376,N_6106,N_6127);
xnor U6377 (N_6377,N_6150,N_6153);
or U6378 (N_6378,N_6211,N_6113);
and U6379 (N_6379,N_6245,N_6000);
or U6380 (N_6380,N_6044,N_6041);
or U6381 (N_6381,N_6297,N_6174);
nand U6382 (N_6382,N_6033,N_6076);
or U6383 (N_6383,N_6112,N_6286);
nand U6384 (N_6384,N_6030,N_6087);
xnor U6385 (N_6385,N_6111,N_6042);
nor U6386 (N_6386,N_6168,N_6028);
nand U6387 (N_6387,N_6039,N_6192);
and U6388 (N_6388,N_6003,N_6091);
xnor U6389 (N_6389,N_6283,N_6266);
xor U6390 (N_6390,N_6188,N_6227);
nand U6391 (N_6391,N_6260,N_6116);
nor U6392 (N_6392,N_6290,N_6235);
nor U6393 (N_6393,N_6124,N_6058);
nand U6394 (N_6394,N_6051,N_6200);
nor U6395 (N_6395,N_6085,N_6029);
xor U6396 (N_6396,N_6229,N_6050);
xor U6397 (N_6397,N_6014,N_6212);
and U6398 (N_6398,N_6214,N_6296);
or U6399 (N_6399,N_6004,N_6265);
nor U6400 (N_6400,N_6195,N_6160);
and U6401 (N_6401,N_6128,N_6217);
or U6402 (N_6402,N_6274,N_6272);
nand U6403 (N_6403,N_6268,N_6163);
nand U6404 (N_6404,N_6237,N_6037);
xor U6405 (N_6405,N_6239,N_6164);
nor U6406 (N_6406,N_6225,N_6040);
nor U6407 (N_6407,N_6096,N_6175);
nand U6408 (N_6408,N_6141,N_6002);
xnor U6409 (N_6409,N_6294,N_6176);
nor U6410 (N_6410,N_6210,N_6125);
and U6411 (N_6411,N_6230,N_6255);
nor U6412 (N_6412,N_6069,N_6066);
and U6413 (N_6413,N_6167,N_6083);
xor U6414 (N_6414,N_6016,N_6022);
xnor U6415 (N_6415,N_6247,N_6291);
nand U6416 (N_6416,N_6105,N_6088);
xnor U6417 (N_6417,N_6169,N_6191);
and U6418 (N_6418,N_6067,N_6089);
nor U6419 (N_6419,N_6072,N_6138);
nand U6420 (N_6420,N_6131,N_6071);
xnor U6421 (N_6421,N_6246,N_6123);
or U6422 (N_6422,N_6289,N_6221);
xor U6423 (N_6423,N_6119,N_6207);
and U6424 (N_6424,N_6298,N_6190);
xnor U6425 (N_6425,N_6159,N_6284);
nor U6426 (N_6426,N_6201,N_6219);
or U6427 (N_6427,N_6135,N_6062);
and U6428 (N_6428,N_6059,N_6024);
xor U6429 (N_6429,N_6251,N_6257);
and U6430 (N_6430,N_6232,N_6117);
nand U6431 (N_6431,N_6172,N_6139);
and U6432 (N_6432,N_6081,N_6137);
nand U6433 (N_6433,N_6108,N_6061);
nand U6434 (N_6434,N_6267,N_6092);
xnor U6435 (N_6435,N_6048,N_6193);
or U6436 (N_6436,N_6216,N_6253);
nor U6437 (N_6437,N_6122,N_6185);
xor U6438 (N_6438,N_6053,N_6005);
and U6439 (N_6439,N_6250,N_6234);
nand U6440 (N_6440,N_6134,N_6186);
nor U6441 (N_6441,N_6049,N_6129);
and U6442 (N_6442,N_6142,N_6182);
and U6443 (N_6443,N_6115,N_6165);
and U6444 (N_6444,N_6248,N_6082);
and U6445 (N_6445,N_6263,N_6262);
or U6446 (N_6446,N_6183,N_6052);
or U6447 (N_6447,N_6178,N_6292);
and U6448 (N_6448,N_6208,N_6107);
nor U6449 (N_6449,N_6008,N_6110);
xnor U6450 (N_6450,N_6208,N_6251);
and U6451 (N_6451,N_6004,N_6198);
and U6452 (N_6452,N_6122,N_6087);
xnor U6453 (N_6453,N_6154,N_6006);
or U6454 (N_6454,N_6129,N_6191);
and U6455 (N_6455,N_6120,N_6130);
nor U6456 (N_6456,N_6272,N_6184);
nand U6457 (N_6457,N_6073,N_6134);
nand U6458 (N_6458,N_6141,N_6275);
nand U6459 (N_6459,N_6152,N_6151);
or U6460 (N_6460,N_6187,N_6065);
or U6461 (N_6461,N_6059,N_6249);
xnor U6462 (N_6462,N_6190,N_6297);
or U6463 (N_6463,N_6070,N_6240);
and U6464 (N_6464,N_6164,N_6181);
nor U6465 (N_6465,N_6204,N_6010);
or U6466 (N_6466,N_6208,N_6239);
and U6467 (N_6467,N_6071,N_6238);
and U6468 (N_6468,N_6245,N_6121);
xor U6469 (N_6469,N_6117,N_6220);
nor U6470 (N_6470,N_6265,N_6155);
or U6471 (N_6471,N_6289,N_6065);
xnor U6472 (N_6472,N_6029,N_6170);
and U6473 (N_6473,N_6113,N_6060);
nor U6474 (N_6474,N_6161,N_6068);
xor U6475 (N_6475,N_6111,N_6197);
and U6476 (N_6476,N_6100,N_6072);
nor U6477 (N_6477,N_6172,N_6249);
or U6478 (N_6478,N_6132,N_6196);
and U6479 (N_6479,N_6008,N_6226);
nor U6480 (N_6480,N_6203,N_6069);
and U6481 (N_6481,N_6157,N_6289);
and U6482 (N_6482,N_6281,N_6022);
nand U6483 (N_6483,N_6086,N_6280);
nand U6484 (N_6484,N_6221,N_6136);
and U6485 (N_6485,N_6011,N_6067);
nor U6486 (N_6486,N_6292,N_6188);
nand U6487 (N_6487,N_6106,N_6089);
nand U6488 (N_6488,N_6260,N_6228);
nand U6489 (N_6489,N_6052,N_6090);
or U6490 (N_6490,N_6184,N_6181);
and U6491 (N_6491,N_6011,N_6074);
or U6492 (N_6492,N_6166,N_6061);
and U6493 (N_6493,N_6274,N_6018);
nor U6494 (N_6494,N_6262,N_6042);
xor U6495 (N_6495,N_6052,N_6295);
and U6496 (N_6496,N_6013,N_6154);
nand U6497 (N_6497,N_6267,N_6271);
nor U6498 (N_6498,N_6196,N_6020);
nand U6499 (N_6499,N_6148,N_6161);
or U6500 (N_6500,N_6142,N_6168);
nor U6501 (N_6501,N_6272,N_6221);
or U6502 (N_6502,N_6081,N_6098);
or U6503 (N_6503,N_6003,N_6225);
xnor U6504 (N_6504,N_6028,N_6119);
nand U6505 (N_6505,N_6284,N_6163);
and U6506 (N_6506,N_6107,N_6061);
xor U6507 (N_6507,N_6273,N_6155);
nor U6508 (N_6508,N_6128,N_6282);
xnor U6509 (N_6509,N_6102,N_6276);
nor U6510 (N_6510,N_6274,N_6235);
xor U6511 (N_6511,N_6261,N_6033);
xnor U6512 (N_6512,N_6166,N_6002);
nand U6513 (N_6513,N_6111,N_6020);
xor U6514 (N_6514,N_6299,N_6008);
nand U6515 (N_6515,N_6070,N_6140);
and U6516 (N_6516,N_6065,N_6113);
nor U6517 (N_6517,N_6014,N_6056);
nand U6518 (N_6518,N_6159,N_6021);
nor U6519 (N_6519,N_6050,N_6278);
xnor U6520 (N_6520,N_6171,N_6093);
and U6521 (N_6521,N_6136,N_6138);
nor U6522 (N_6522,N_6097,N_6246);
or U6523 (N_6523,N_6172,N_6259);
xor U6524 (N_6524,N_6111,N_6277);
or U6525 (N_6525,N_6097,N_6118);
nand U6526 (N_6526,N_6298,N_6202);
or U6527 (N_6527,N_6237,N_6209);
xor U6528 (N_6528,N_6046,N_6208);
and U6529 (N_6529,N_6246,N_6226);
xor U6530 (N_6530,N_6079,N_6255);
nor U6531 (N_6531,N_6028,N_6238);
or U6532 (N_6532,N_6011,N_6179);
nor U6533 (N_6533,N_6003,N_6066);
and U6534 (N_6534,N_6146,N_6137);
nor U6535 (N_6535,N_6068,N_6190);
and U6536 (N_6536,N_6233,N_6037);
xor U6537 (N_6537,N_6284,N_6286);
and U6538 (N_6538,N_6154,N_6144);
or U6539 (N_6539,N_6112,N_6089);
xnor U6540 (N_6540,N_6095,N_6237);
xnor U6541 (N_6541,N_6171,N_6232);
xor U6542 (N_6542,N_6198,N_6166);
nor U6543 (N_6543,N_6049,N_6115);
and U6544 (N_6544,N_6121,N_6091);
xnor U6545 (N_6545,N_6266,N_6052);
and U6546 (N_6546,N_6289,N_6151);
and U6547 (N_6547,N_6065,N_6084);
or U6548 (N_6548,N_6137,N_6240);
nor U6549 (N_6549,N_6113,N_6018);
nand U6550 (N_6550,N_6137,N_6272);
xor U6551 (N_6551,N_6151,N_6231);
or U6552 (N_6552,N_6153,N_6229);
nand U6553 (N_6553,N_6266,N_6028);
and U6554 (N_6554,N_6072,N_6262);
xnor U6555 (N_6555,N_6176,N_6070);
xnor U6556 (N_6556,N_6022,N_6160);
and U6557 (N_6557,N_6156,N_6164);
nand U6558 (N_6558,N_6001,N_6276);
nor U6559 (N_6559,N_6292,N_6130);
and U6560 (N_6560,N_6071,N_6007);
xnor U6561 (N_6561,N_6089,N_6278);
xor U6562 (N_6562,N_6120,N_6195);
xnor U6563 (N_6563,N_6150,N_6170);
nor U6564 (N_6564,N_6131,N_6169);
nor U6565 (N_6565,N_6155,N_6179);
nand U6566 (N_6566,N_6209,N_6133);
nand U6567 (N_6567,N_6221,N_6043);
and U6568 (N_6568,N_6148,N_6066);
or U6569 (N_6569,N_6134,N_6266);
or U6570 (N_6570,N_6167,N_6146);
nand U6571 (N_6571,N_6051,N_6292);
xor U6572 (N_6572,N_6141,N_6292);
xnor U6573 (N_6573,N_6240,N_6261);
and U6574 (N_6574,N_6214,N_6016);
nor U6575 (N_6575,N_6074,N_6127);
nand U6576 (N_6576,N_6064,N_6224);
xor U6577 (N_6577,N_6024,N_6254);
xnor U6578 (N_6578,N_6224,N_6087);
and U6579 (N_6579,N_6295,N_6182);
or U6580 (N_6580,N_6209,N_6020);
nand U6581 (N_6581,N_6085,N_6212);
xnor U6582 (N_6582,N_6087,N_6036);
xnor U6583 (N_6583,N_6082,N_6050);
or U6584 (N_6584,N_6141,N_6229);
nand U6585 (N_6585,N_6056,N_6120);
or U6586 (N_6586,N_6199,N_6190);
or U6587 (N_6587,N_6204,N_6261);
and U6588 (N_6588,N_6098,N_6210);
or U6589 (N_6589,N_6227,N_6264);
and U6590 (N_6590,N_6202,N_6080);
or U6591 (N_6591,N_6104,N_6048);
nor U6592 (N_6592,N_6220,N_6226);
nand U6593 (N_6593,N_6181,N_6176);
nor U6594 (N_6594,N_6218,N_6269);
or U6595 (N_6595,N_6166,N_6172);
xnor U6596 (N_6596,N_6238,N_6078);
xor U6597 (N_6597,N_6251,N_6016);
nor U6598 (N_6598,N_6264,N_6185);
nor U6599 (N_6599,N_6008,N_6138);
nand U6600 (N_6600,N_6551,N_6516);
or U6601 (N_6601,N_6333,N_6321);
nor U6602 (N_6602,N_6350,N_6398);
nor U6603 (N_6603,N_6420,N_6484);
nor U6604 (N_6604,N_6366,N_6590);
and U6605 (N_6605,N_6482,N_6523);
or U6606 (N_6606,N_6370,N_6494);
xnor U6607 (N_6607,N_6382,N_6446);
nand U6608 (N_6608,N_6584,N_6395);
and U6609 (N_6609,N_6381,N_6452);
and U6610 (N_6610,N_6463,N_6396);
nand U6611 (N_6611,N_6515,N_6388);
xnor U6612 (N_6612,N_6307,N_6409);
xor U6613 (N_6613,N_6471,N_6344);
xor U6614 (N_6614,N_6433,N_6392);
xnor U6615 (N_6615,N_6303,N_6456);
nand U6616 (N_6616,N_6541,N_6425);
or U6617 (N_6617,N_6459,N_6363);
xor U6618 (N_6618,N_6436,N_6449);
and U6619 (N_6619,N_6528,N_6427);
nand U6620 (N_6620,N_6473,N_6326);
nand U6621 (N_6621,N_6415,N_6592);
or U6622 (N_6622,N_6549,N_6499);
or U6623 (N_6623,N_6525,N_6569);
nand U6624 (N_6624,N_6393,N_6376);
and U6625 (N_6625,N_6531,N_6576);
xor U6626 (N_6626,N_6383,N_6357);
and U6627 (N_6627,N_6511,N_6588);
or U6628 (N_6628,N_6553,N_6422);
and U6629 (N_6629,N_6330,N_6517);
xnor U6630 (N_6630,N_6458,N_6340);
nand U6631 (N_6631,N_6390,N_6430);
nand U6632 (N_6632,N_6410,N_6416);
nand U6633 (N_6633,N_6597,N_6336);
xnor U6634 (N_6634,N_6571,N_6489);
xnor U6635 (N_6635,N_6419,N_6308);
nor U6636 (N_6636,N_6426,N_6478);
xnor U6637 (N_6637,N_6387,N_6341);
xor U6638 (N_6638,N_6552,N_6538);
nor U6639 (N_6639,N_6447,N_6497);
nor U6640 (N_6640,N_6580,N_6324);
nor U6641 (N_6641,N_6522,N_6506);
or U6642 (N_6642,N_6573,N_6323);
nand U6643 (N_6643,N_6359,N_6406);
xnor U6644 (N_6644,N_6556,N_6527);
xnor U6645 (N_6645,N_6502,N_6411);
nor U6646 (N_6646,N_6413,N_6306);
and U6647 (N_6647,N_6364,N_6334);
and U6648 (N_6648,N_6477,N_6487);
or U6649 (N_6649,N_6479,N_6582);
nand U6650 (N_6650,N_6310,N_6464);
and U6651 (N_6651,N_6399,N_6345);
or U6652 (N_6652,N_6378,N_6457);
and U6653 (N_6653,N_6567,N_6435);
xor U6654 (N_6654,N_6520,N_6309);
or U6655 (N_6655,N_6431,N_6314);
xnor U6656 (N_6656,N_6455,N_6480);
or U6657 (N_6657,N_6389,N_6402);
nand U6658 (N_6658,N_6300,N_6493);
and U6659 (N_6659,N_6587,N_6379);
xor U6660 (N_6660,N_6441,N_6562);
nor U6661 (N_6661,N_6377,N_6533);
or U6662 (N_6662,N_6346,N_6405);
nand U6663 (N_6663,N_6529,N_6437);
and U6664 (N_6664,N_6461,N_6512);
xnor U6665 (N_6665,N_6353,N_6375);
and U6666 (N_6666,N_6470,N_6347);
nor U6667 (N_6667,N_6380,N_6475);
and U6668 (N_6668,N_6579,N_6524);
xnor U6669 (N_6669,N_6554,N_6578);
xnor U6670 (N_6670,N_6443,N_6490);
and U6671 (N_6671,N_6591,N_6414);
nor U6672 (N_6672,N_6434,N_6439);
xor U6673 (N_6673,N_6474,N_6355);
nand U6674 (N_6674,N_6412,N_6599);
and U6675 (N_6675,N_6566,N_6574);
or U6676 (N_6676,N_6598,N_6327);
nor U6677 (N_6677,N_6561,N_6301);
nor U6678 (N_6678,N_6325,N_6544);
xnor U6679 (N_6679,N_6444,N_6338);
or U6680 (N_6680,N_6450,N_6401);
nor U6681 (N_6681,N_6408,N_6537);
or U6682 (N_6682,N_6467,N_6445);
and U6683 (N_6683,N_6486,N_6407);
nor U6684 (N_6684,N_6540,N_6384);
and U6685 (N_6685,N_6335,N_6558);
xor U6686 (N_6686,N_6348,N_6596);
nor U6687 (N_6687,N_6491,N_6351);
nor U6688 (N_6688,N_6429,N_6485);
xnor U6689 (N_6689,N_6440,N_6583);
nand U6690 (N_6690,N_6373,N_6460);
xor U6691 (N_6691,N_6318,N_6547);
or U6692 (N_6692,N_6371,N_6400);
nand U6693 (N_6693,N_6332,N_6313);
xnor U6694 (N_6694,N_6545,N_6394);
or U6695 (N_6695,N_6305,N_6386);
and U6696 (N_6696,N_6488,N_6331);
xnor U6697 (N_6697,N_6374,N_6403);
nand U6698 (N_6698,N_6481,N_6421);
nand U6699 (N_6699,N_6570,N_6385);
xor U6700 (N_6700,N_6543,N_6503);
nor U6701 (N_6701,N_6468,N_6311);
nor U6702 (N_6702,N_6526,N_6509);
nor U6703 (N_6703,N_6397,N_6352);
and U6704 (N_6704,N_6368,N_6535);
nand U6705 (N_6705,N_6572,N_6565);
nor U6706 (N_6706,N_6586,N_6342);
nor U6707 (N_6707,N_6304,N_6404);
nor U6708 (N_6708,N_6365,N_6563);
xnor U6709 (N_6709,N_6560,N_6536);
nand U6710 (N_6710,N_6557,N_6302);
or U6711 (N_6711,N_6507,N_6514);
nor U6712 (N_6712,N_6360,N_6519);
nand U6713 (N_6713,N_6589,N_6500);
nand U6714 (N_6714,N_6492,N_6339);
or U6715 (N_6715,N_6476,N_6498);
or U6716 (N_6716,N_6423,N_6513);
nand U6717 (N_6717,N_6518,N_6451);
nor U6718 (N_6718,N_6539,N_6372);
and U6719 (N_6719,N_6542,N_6510);
and U6720 (N_6720,N_6530,N_6532);
or U6721 (N_6721,N_6568,N_6564);
nor U6722 (N_6722,N_6593,N_6454);
xor U6723 (N_6723,N_6362,N_6391);
and U6724 (N_6724,N_6442,N_6462);
and U6725 (N_6725,N_6438,N_6521);
or U6726 (N_6726,N_6317,N_6483);
nor U6727 (N_6727,N_6428,N_6581);
nor U6728 (N_6728,N_6322,N_6417);
or U6729 (N_6729,N_6329,N_6496);
nor U6730 (N_6730,N_6555,N_6575);
or U6731 (N_6731,N_6534,N_6550);
nor U6732 (N_6732,N_6577,N_6343);
or U6733 (N_6733,N_6585,N_6337);
and U6734 (N_6734,N_6315,N_6548);
nor U6735 (N_6735,N_6369,N_6465);
nand U6736 (N_6736,N_6448,N_6504);
and U6737 (N_6737,N_6367,N_6319);
or U6738 (N_6738,N_6424,N_6469);
nand U6739 (N_6739,N_6418,N_6466);
or U6740 (N_6740,N_6349,N_6495);
nor U6741 (N_6741,N_6356,N_6546);
nor U6742 (N_6742,N_6594,N_6320);
and U6743 (N_6743,N_6508,N_6505);
and U6744 (N_6744,N_6595,N_6453);
or U6745 (N_6745,N_6472,N_6501);
and U6746 (N_6746,N_6316,N_6358);
nand U6747 (N_6747,N_6328,N_6354);
xor U6748 (N_6748,N_6361,N_6432);
xnor U6749 (N_6749,N_6559,N_6312);
or U6750 (N_6750,N_6593,N_6430);
nor U6751 (N_6751,N_6440,N_6449);
and U6752 (N_6752,N_6463,N_6339);
and U6753 (N_6753,N_6588,N_6310);
and U6754 (N_6754,N_6380,N_6576);
and U6755 (N_6755,N_6465,N_6356);
or U6756 (N_6756,N_6404,N_6421);
xnor U6757 (N_6757,N_6593,N_6563);
nand U6758 (N_6758,N_6593,N_6536);
nand U6759 (N_6759,N_6395,N_6322);
or U6760 (N_6760,N_6520,N_6408);
xnor U6761 (N_6761,N_6528,N_6470);
or U6762 (N_6762,N_6582,N_6572);
nor U6763 (N_6763,N_6437,N_6362);
or U6764 (N_6764,N_6404,N_6508);
or U6765 (N_6765,N_6365,N_6352);
nand U6766 (N_6766,N_6558,N_6595);
and U6767 (N_6767,N_6578,N_6362);
nor U6768 (N_6768,N_6318,N_6436);
or U6769 (N_6769,N_6355,N_6428);
xor U6770 (N_6770,N_6544,N_6345);
and U6771 (N_6771,N_6491,N_6550);
nor U6772 (N_6772,N_6578,N_6431);
and U6773 (N_6773,N_6571,N_6546);
and U6774 (N_6774,N_6351,N_6411);
nand U6775 (N_6775,N_6595,N_6593);
xnor U6776 (N_6776,N_6587,N_6476);
or U6777 (N_6777,N_6556,N_6590);
nand U6778 (N_6778,N_6392,N_6327);
xnor U6779 (N_6779,N_6534,N_6452);
nand U6780 (N_6780,N_6454,N_6515);
or U6781 (N_6781,N_6484,N_6352);
nand U6782 (N_6782,N_6543,N_6414);
and U6783 (N_6783,N_6390,N_6423);
nand U6784 (N_6784,N_6402,N_6411);
and U6785 (N_6785,N_6528,N_6327);
nor U6786 (N_6786,N_6534,N_6370);
nand U6787 (N_6787,N_6344,N_6508);
xnor U6788 (N_6788,N_6564,N_6475);
and U6789 (N_6789,N_6350,N_6393);
nand U6790 (N_6790,N_6314,N_6394);
or U6791 (N_6791,N_6485,N_6559);
nand U6792 (N_6792,N_6326,N_6511);
nor U6793 (N_6793,N_6310,N_6534);
and U6794 (N_6794,N_6518,N_6524);
nor U6795 (N_6795,N_6488,N_6376);
xor U6796 (N_6796,N_6460,N_6365);
and U6797 (N_6797,N_6553,N_6361);
and U6798 (N_6798,N_6356,N_6511);
nand U6799 (N_6799,N_6386,N_6395);
and U6800 (N_6800,N_6363,N_6493);
xnor U6801 (N_6801,N_6503,N_6564);
nand U6802 (N_6802,N_6386,N_6472);
or U6803 (N_6803,N_6310,N_6357);
nand U6804 (N_6804,N_6561,N_6418);
nand U6805 (N_6805,N_6449,N_6419);
or U6806 (N_6806,N_6558,N_6379);
xor U6807 (N_6807,N_6527,N_6406);
and U6808 (N_6808,N_6482,N_6408);
or U6809 (N_6809,N_6568,N_6355);
and U6810 (N_6810,N_6577,N_6365);
xnor U6811 (N_6811,N_6583,N_6594);
or U6812 (N_6812,N_6520,N_6436);
xnor U6813 (N_6813,N_6306,N_6353);
nand U6814 (N_6814,N_6444,N_6545);
nand U6815 (N_6815,N_6425,N_6553);
and U6816 (N_6816,N_6403,N_6472);
nand U6817 (N_6817,N_6400,N_6418);
nand U6818 (N_6818,N_6307,N_6513);
and U6819 (N_6819,N_6390,N_6547);
or U6820 (N_6820,N_6464,N_6481);
or U6821 (N_6821,N_6572,N_6301);
nor U6822 (N_6822,N_6381,N_6407);
nand U6823 (N_6823,N_6551,N_6519);
nand U6824 (N_6824,N_6375,N_6441);
nor U6825 (N_6825,N_6592,N_6541);
and U6826 (N_6826,N_6457,N_6515);
nor U6827 (N_6827,N_6508,N_6558);
or U6828 (N_6828,N_6597,N_6394);
and U6829 (N_6829,N_6455,N_6300);
nor U6830 (N_6830,N_6494,N_6590);
nand U6831 (N_6831,N_6324,N_6357);
xnor U6832 (N_6832,N_6355,N_6547);
nor U6833 (N_6833,N_6571,N_6460);
nor U6834 (N_6834,N_6374,N_6489);
and U6835 (N_6835,N_6514,N_6335);
nand U6836 (N_6836,N_6320,N_6490);
nor U6837 (N_6837,N_6402,N_6390);
and U6838 (N_6838,N_6475,N_6483);
nand U6839 (N_6839,N_6505,N_6409);
nand U6840 (N_6840,N_6488,N_6305);
nand U6841 (N_6841,N_6409,N_6319);
nor U6842 (N_6842,N_6402,N_6482);
nand U6843 (N_6843,N_6536,N_6314);
xnor U6844 (N_6844,N_6492,N_6407);
xor U6845 (N_6845,N_6588,N_6507);
nor U6846 (N_6846,N_6498,N_6470);
nor U6847 (N_6847,N_6395,N_6347);
nand U6848 (N_6848,N_6570,N_6516);
nand U6849 (N_6849,N_6488,N_6523);
nand U6850 (N_6850,N_6584,N_6530);
xor U6851 (N_6851,N_6431,N_6425);
nor U6852 (N_6852,N_6516,N_6445);
xor U6853 (N_6853,N_6327,N_6452);
xnor U6854 (N_6854,N_6503,N_6496);
and U6855 (N_6855,N_6559,N_6496);
nand U6856 (N_6856,N_6372,N_6358);
or U6857 (N_6857,N_6556,N_6558);
xor U6858 (N_6858,N_6544,N_6364);
and U6859 (N_6859,N_6385,N_6443);
or U6860 (N_6860,N_6544,N_6579);
and U6861 (N_6861,N_6501,N_6453);
nand U6862 (N_6862,N_6308,N_6445);
and U6863 (N_6863,N_6580,N_6552);
nor U6864 (N_6864,N_6493,N_6428);
nor U6865 (N_6865,N_6384,N_6450);
and U6866 (N_6866,N_6501,N_6328);
nand U6867 (N_6867,N_6407,N_6355);
or U6868 (N_6868,N_6373,N_6550);
xnor U6869 (N_6869,N_6370,N_6417);
and U6870 (N_6870,N_6597,N_6513);
or U6871 (N_6871,N_6305,N_6459);
xnor U6872 (N_6872,N_6560,N_6507);
or U6873 (N_6873,N_6352,N_6512);
nor U6874 (N_6874,N_6460,N_6368);
xor U6875 (N_6875,N_6412,N_6524);
xor U6876 (N_6876,N_6533,N_6531);
xor U6877 (N_6877,N_6468,N_6549);
nor U6878 (N_6878,N_6590,N_6333);
or U6879 (N_6879,N_6404,N_6378);
and U6880 (N_6880,N_6538,N_6303);
and U6881 (N_6881,N_6547,N_6571);
and U6882 (N_6882,N_6474,N_6592);
xor U6883 (N_6883,N_6324,N_6352);
xnor U6884 (N_6884,N_6595,N_6400);
nand U6885 (N_6885,N_6498,N_6306);
xnor U6886 (N_6886,N_6396,N_6465);
nor U6887 (N_6887,N_6327,N_6439);
nand U6888 (N_6888,N_6371,N_6422);
xnor U6889 (N_6889,N_6522,N_6345);
and U6890 (N_6890,N_6430,N_6597);
nor U6891 (N_6891,N_6326,N_6373);
nor U6892 (N_6892,N_6466,N_6591);
nor U6893 (N_6893,N_6456,N_6357);
nand U6894 (N_6894,N_6501,N_6512);
xnor U6895 (N_6895,N_6471,N_6546);
xor U6896 (N_6896,N_6337,N_6433);
and U6897 (N_6897,N_6497,N_6551);
nand U6898 (N_6898,N_6343,N_6553);
xor U6899 (N_6899,N_6516,N_6484);
nor U6900 (N_6900,N_6691,N_6820);
and U6901 (N_6901,N_6759,N_6608);
xnor U6902 (N_6902,N_6642,N_6626);
nor U6903 (N_6903,N_6693,N_6671);
nor U6904 (N_6904,N_6739,N_6833);
and U6905 (N_6905,N_6708,N_6782);
xor U6906 (N_6906,N_6712,N_6766);
nor U6907 (N_6907,N_6715,N_6618);
xnor U6908 (N_6908,N_6748,N_6772);
nor U6909 (N_6909,N_6711,N_6824);
nor U6910 (N_6910,N_6760,N_6605);
xor U6911 (N_6911,N_6835,N_6790);
nand U6912 (N_6912,N_6768,N_6873);
nor U6913 (N_6913,N_6675,N_6845);
xor U6914 (N_6914,N_6749,N_6807);
xor U6915 (N_6915,N_6789,N_6727);
nor U6916 (N_6916,N_6756,N_6813);
xor U6917 (N_6917,N_6705,N_6633);
xor U6918 (N_6918,N_6639,N_6850);
nand U6919 (N_6919,N_6791,N_6899);
and U6920 (N_6920,N_6604,N_6830);
or U6921 (N_6921,N_6855,N_6617);
xor U6922 (N_6922,N_6891,N_6754);
nand U6923 (N_6923,N_6848,N_6616);
and U6924 (N_6924,N_6630,N_6659);
nor U6925 (N_6925,N_6752,N_6796);
xnor U6926 (N_6926,N_6623,N_6722);
xnor U6927 (N_6927,N_6846,N_6731);
or U6928 (N_6928,N_6704,N_6734);
nor U6929 (N_6929,N_6612,N_6720);
nor U6930 (N_6930,N_6825,N_6888);
or U6931 (N_6931,N_6866,N_6613);
and U6932 (N_6932,N_6716,N_6742);
nor U6933 (N_6933,N_6680,N_6627);
or U6934 (N_6934,N_6672,N_6816);
nand U6935 (N_6935,N_6634,N_6829);
and U6936 (N_6936,N_6643,N_6859);
nor U6937 (N_6937,N_6834,N_6838);
xor U6938 (N_6938,N_6849,N_6883);
nor U6939 (N_6939,N_6644,N_6783);
xnor U6940 (N_6940,N_6778,N_6786);
and U6941 (N_6941,N_6890,N_6684);
and U6942 (N_6942,N_6867,N_6694);
xor U6943 (N_6943,N_6826,N_6682);
xor U6944 (N_6944,N_6851,N_6836);
nand U6945 (N_6945,N_6865,N_6841);
nor U6946 (N_6946,N_6886,N_6831);
xor U6947 (N_6947,N_6878,N_6755);
nand U6948 (N_6948,N_6858,N_6677);
xor U6949 (N_6949,N_6812,N_6687);
nand U6950 (N_6950,N_6713,N_6664);
and U6951 (N_6951,N_6800,N_6614);
and U6952 (N_6952,N_6674,N_6863);
or U6953 (N_6953,N_6894,N_6856);
nor U6954 (N_6954,N_6769,N_6655);
or U6955 (N_6955,N_6678,N_6663);
nand U6956 (N_6956,N_6828,N_6723);
nor U6957 (N_6957,N_6624,N_6683);
nor U6958 (N_6958,N_6628,N_6897);
nand U6959 (N_6959,N_6601,N_6870);
nor U6960 (N_6960,N_6681,N_6810);
and U6961 (N_6961,N_6893,N_6648);
nand U6962 (N_6962,N_6822,N_6788);
nor U6963 (N_6963,N_6762,N_6741);
and U6964 (N_6964,N_6780,N_6864);
nand U6965 (N_6965,N_6877,N_6717);
nand U6966 (N_6966,N_6821,N_6811);
and U6967 (N_6967,N_6736,N_6606);
or U6968 (N_6968,N_6666,N_6654);
and U6969 (N_6969,N_6844,N_6730);
nor U6970 (N_6970,N_6652,N_6869);
or U6971 (N_6971,N_6853,N_6765);
and U6972 (N_6972,N_6806,N_6771);
and U6973 (N_6973,N_6876,N_6898);
nand U6974 (N_6974,N_6697,N_6882);
nand U6975 (N_6975,N_6843,N_6615);
or U6976 (N_6976,N_6706,N_6745);
nor U6977 (N_6977,N_6602,N_6868);
nand U6978 (N_6978,N_6637,N_6784);
xor U6979 (N_6979,N_6874,N_6690);
and U6980 (N_6980,N_6857,N_6764);
xnor U6981 (N_6981,N_6719,N_6889);
nor U6982 (N_6982,N_6703,N_6647);
or U6983 (N_6983,N_6640,N_6885);
nand U6984 (N_6984,N_6662,N_6802);
nor U6985 (N_6985,N_6653,N_6793);
nand U6986 (N_6986,N_6718,N_6610);
or U6987 (N_6987,N_6732,N_6611);
nand U6988 (N_6988,N_6700,N_6747);
and U6989 (N_6989,N_6740,N_6638);
nor U6990 (N_6990,N_6636,N_6641);
nand U6991 (N_6991,N_6696,N_6798);
nor U6992 (N_6992,N_6896,N_6686);
or U6993 (N_6993,N_6862,N_6887);
and U6994 (N_6994,N_6805,N_6699);
nor U6995 (N_6995,N_6724,N_6629);
and U6996 (N_6996,N_6668,N_6702);
xor U6997 (N_6997,N_6679,N_6657);
and U6998 (N_6998,N_6767,N_6685);
xor U6999 (N_6999,N_6880,N_6854);
xor U7000 (N_7000,N_6650,N_6743);
nand U7001 (N_7001,N_6842,N_6799);
or U7002 (N_7002,N_6881,N_6701);
xor U7003 (N_7003,N_6603,N_6872);
nand U7004 (N_7004,N_6832,N_6660);
nand U7005 (N_7005,N_6775,N_6707);
nor U7006 (N_7006,N_6710,N_6669);
nand U7007 (N_7007,N_6620,N_6773);
and U7008 (N_7008,N_6794,N_6632);
nor U7009 (N_7009,N_6808,N_6779);
and U7010 (N_7010,N_6757,N_6744);
xnor U7011 (N_7011,N_6797,N_6688);
xor U7012 (N_7012,N_6665,N_6656);
xnor U7013 (N_7013,N_6667,N_6635);
nand U7014 (N_7014,N_6733,N_6792);
or U7015 (N_7015,N_6827,N_6692);
or U7016 (N_7016,N_6726,N_6737);
nor U7017 (N_7017,N_6884,N_6750);
or U7018 (N_7018,N_6709,N_6646);
nand U7019 (N_7019,N_6729,N_6631);
and U7020 (N_7020,N_6763,N_6621);
nand U7021 (N_7021,N_6676,N_6774);
nor U7022 (N_7022,N_6809,N_6761);
xor U7023 (N_7023,N_6728,N_6651);
or U7024 (N_7024,N_6819,N_6879);
nand U7025 (N_7025,N_6892,N_6847);
xor U7026 (N_7026,N_6817,N_6625);
nor U7027 (N_7027,N_6695,N_6785);
nor U7028 (N_7028,N_6746,N_6895);
xor U7029 (N_7029,N_6801,N_6776);
nand U7030 (N_7030,N_6804,N_6803);
or U7031 (N_7031,N_6751,N_6871);
xnor U7032 (N_7032,N_6649,N_6840);
nor U7033 (N_7033,N_6852,N_6725);
nor U7034 (N_7034,N_6714,N_6673);
xnor U7035 (N_7035,N_6670,N_6609);
nand U7036 (N_7036,N_6658,N_6600);
nor U7037 (N_7037,N_6622,N_6875);
nor U7038 (N_7038,N_6861,N_6738);
nand U7039 (N_7039,N_6607,N_6837);
nor U7040 (N_7040,N_6753,N_6619);
and U7041 (N_7041,N_6860,N_6689);
nand U7042 (N_7042,N_6770,N_6777);
and U7043 (N_7043,N_6818,N_6645);
nor U7044 (N_7044,N_6661,N_6815);
and U7045 (N_7045,N_6735,N_6787);
and U7046 (N_7046,N_6814,N_6839);
nand U7047 (N_7047,N_6758,N_6795);
and U7048 (N_7048,N_6721,N_6698);
nor U7049 (N_7049,N_6781,N_6823);
xor U7050 (N_7050,N_6704,N_6624);
xor U7051 (N_7051,N_6722,N_6834);
or U7052 (N_7052,N_6681,N_6661);
xnor U7053 (N_7053,N_6778,N_6862);
and U7054 (N_7054,N_6696,N_6609);
or U7055 (N_7055,N_6776,N_6839);
or U7056 (N_7056,N_6889,N_6766);
nor U7057 (N_7057,N_6745,N_6605);
or U7058 (N_7058,N_6754,N_6781);
or U7059 (N_7059,N_6635,N_6798);
and U7060 (N_7060,N_6695,N_6775);
nand U7061 (N_7061,N_6760,N_6884);
nor U7062 (N_7062,N_6617,N_6716);
nor U7063 (N_7063,N_6733,N_6837);
nand U7064 (N_7064,N_6806,N_6683);
or U7065 (N_7065,N_6828,N_6676);
or U7066 (N_7066,N_6646,N_6800);
or U7067 (N_7067,N_6842,N_6668);
nand U7068 (N_7068,N_6840,N_6796);
xnor U7069 (N_7069,N_6609,N_6851);
and U7070 (N_7070,N_6650,N_6800);
nand U7071 (N_7071,N_6631,N_6780);
or U7072 (N_7072,N_6633,N_6761);
and U7073 (N_7073,N_6879,N_6716);
xor U7074 (N_7074,N_6835,N_6648);
xor U7075 (N_7075,N_6685,N_6742);
nand U7076 (N_7076,N_6899,N_6717);
xor U7077 (N_7077,N_6895,N_6878);
and U7078 (N_7078,N_6811,N_6757);
and U7079 (N_7079,N_6852,N_6805);
nor U7080 (N_7080,N_6824,N_6788);
or U7081 (N_7081,N_6883,N_6808);
and U7082 (N_7082,N_6711,N_6753);
xnor U7083 (N_7083,N_6823,N_6614);
nand U7084 (N_7084,N_6670,N_6682);
nand U7085 (N_7085,N_6690,N_6811);
nand U7086 (N_7086,N_6853,N_6696);
or U7087 (N_7087,N_6743,N_6667);
and U7088 (N_7088,N_6717,N_6874);
xnor U7089 (N_7089,N_6704,N_6708);
nand U7090 (N_7090,N_6675,N_6684);
nor U7091 (N_7091,N_6610,N_6743);
or U7092 (N_7092,N_6669,N_6727);
or U7093 (N_7093,N_6745,N_6715);
nor U7094 (N_7094,N_6743,N_6805);
nor U7095 (N_7095,N_6866,N_6700);
xor U7096 (N_7096,N_6721,N_6668);
or U7097 (N_7097,N_6876,N_6754);
xor U7098 (N_7098,N_6660,N_6645);
nand U7099 (N_7099,N_6720,N_6771);
or U7100 (N_7100,N_6617,N_6794);
nand U7101 (N_7101,N_6747,N_6711);
nand U7102 (N_7102,N_6803,N_6828);
or U7103 (N_7103,N_6788,N_6838);
and U7104 (N_7104,N_6771,N_6792);
nand U7105 (N_7105,N_6853,N_6794);
and U7106 (N_7106,N_6889,N_6631);
or U7107 (N_7107,N_6887,N_6759);
or U7108 (N_7108,N_6838,N_6816);
xor U7109 (N_7109,N_6806,N_6622);
nand U7110 (N_7110,N_6770,N_6739);
xnor U7111 (N_7111,N_6747,N_6890);
and U7112 (N_7112,N_6810,N_6881);
and U7113 (N_7113,N_6657,N_6680);
and U7114 (N_7114,N_6779,N_6646);
nor U7115 (N_7115,N_6746,N_6871);
and U7116 (N_7116,N_6601,N_6769);
or U7117 (N_7117,N_6671,N_6811);
and U7118 (N_7118,N_6745,N_6827);
nand U7119 (N_7119,N_6676,N_6883);
nand U7120 (N_7120,N_6610,N_6628);
nand U7121 (N_7121,N_6636,N_6654);
nor U7122 (N_7122,N_6868,N_6774);
nand U7123 (N_7123,N_6689,N_6886);
or U7124 (N_7124,N_6658,N_6838);
nor U7125 (N_7125,N_6639,N_6710);
nand U7126 (N_7126,N_6834,N_6844);
nand U7127 (N_7127,N_6869,N_6657);
xnor U7128 (N_7128,N_6645,N_6621);
xor U7129 (N_7129,N_6878,N_6792);
and U7130 (N_7130,N_6842,N_6751);
xnor U7131 (N_7131,N_6623,N_6763);
xor U7132 (N_7132,N_6637,N_6817);
xor U7133 (N_7133,N_6694,N_6788);
xor U7134 (N_7134,N_6726,N_6832);
and U7135 (N_7135,N_6875,N_6860);
nand U7136 (N_7136,N_6603,N_6691);
nand U7137 (N_7137,N_6820,N_6891);
nor U7138 (N_7138,N_6865,N_6722);
nor U7139 (N_7139,N_6879,N_6817);
nand U7140 (N_7140,N_6889,N_6646);
xor U7141 (N_7141,N_6736,N_6845);
or U7142 (N_7142,N_6730,N_6709);
nand U7143 (N_7143,N_6868,N_6753);
nand U7144 (N_7144,N_6815,N_6790);
or U7145 (N_7145,N_6719,N_6876);
and U7146 (N_7146,N_6665,N_6851);
and U7147 (N_7147,N_6730,N_6659);
xnor U7148 (N_7148,N_6638,N_6853);
xor U7149 (N_7149,N_6771,N_6694);
or U7150 (N_7150,N_6846,N_6802);
nand U7151 (N_7151,N_6897,N_6834);
nand U7152 (N_7152,N_6721,N_6744);
xor U7153 (N_7153,N_6742,N_6654);
or U7154 (N_7154,N_6681,N_6811);
or U7155 (N_7155,N_6755,N_6712);
nand U7156 (N_7156,N_6632,N_6753);
or U7157 (N_7157,N_6821,N_6770);
nand U7158 (N_7158,N_6770,N_6757);
nand U7159 (N_7159,N_6665,N_6711);
or U7160 (N_7160,N_6799,N_6673);
and U7161 (N_7161,N_6767,N_6651);
nor U7162 (N_7162,N_6684,N_6616);
xor U7163 (N_7163,N_6646,N_6781);
xnor U7164 (N_7164,N_6848,N_6673);
and U7165 (N_7165,N_6725,N_6802);
or U7166 (N_7166,N_6866,N_6725);
nor U7167 (N_7167,N_6865,N_6657);
xnor U7168 (N_7168,N_6840,N_6613);
xnor U7169 (N_7169,N_6703,N_6668);
and U7170 (N_7170,N_6887,N_6811);
or U7171 (N_7171,N_6799,N_6890);
nor U7172 (N_7172,N_6765,N_6696);
nand U7173 (N_7173,N_6763,N_6606);
nand U7174 (N_7174,N_6761,N_6646);
or U7175 (N_7175,N_6658,N_6835);
nor U7176 (N_7176,N_6714,N_6629);
and U7177 (N_7177,N_6855,N_6761);
nand U7178 (N_7178,N_6892,N_6816);
nor U7179 (N_7179,N_6871,N_6771);
xor U7180 (N_7180,N_6849,N_6674);
and U7181 (N_7181,N_6658,N_6886);
or U7182 (N_7182,N_6676,N_6743);
and U7183 (N_7183,N_6762,N_6822);
xnor U7184 (N_7184,N_6690,N_6834);
and U7185 (N_7185,N_6826,N_6853);
nor U7186 (N_7186,N_6751,N_6639);
nor U7187 (N_7187,N_6840,N_6899);
and U7188 (N_7188,N_6845,N_6620);
nand U7189 (N_7189,N_6776,N_6826);
xnor U7190 (N_7190,N_6832,N_6851);
nor U7191 (N_7191,N_6745,N_6846);
and U7192 (N_7192,N_6711,N_6618);
or U7193 (N_7193,N_6806,N_6670);
or U7194 (N_7194,N_6606,N_6871);
nand U7195 (N_7195,N_6699,N_6678);
xnor U7196 (N_7196,N_6665,N_6864);
or U7197 (N_7197,N_6702,N_6849);
or U7198 (N_7198,N_6789,N_6759);
nand U7199 (N_7199,N_6609,N_6754);
or U7200 (N_7200,N_7066,N_7164);
or U7201 (N_7201,N_7138,N_6971);
and U7202 (N_7202,N_6955,N_7070);
and U7203 (N_7203,N_7150,N_7182);
nor U7204 (N_7204,N_7013,N_7012);
nand U7205 (N_7205,N_6927,N_6950);
xnor U7206 (N_7206,N_7133,N_6930);
or U7207 (N_7207,N_6965,N_7109);
and U7208 (N_7208,N_7049,N_7088);
nor U7209 (N_7209,N_6960,N_7082);
and U7210 (N_7210,N_7015,N_7187);
and U7211 (N_7211,N_6936,N_7031);
or U7212 (N_7212,N_7081,N_7148);
or U7213 (N_7213,N_7016,N_7160);
or U7214 (N_7214,N_6951,N_6948);
nor U7215 (N_7215,N_6975,N_7085);
nand U7216 (N_7216,N_7143,N_7137);
and U7217 (N_7217,N_7095,N_7147);
nand U7218 (N_7218,N_7196,N_7072);
nand U7219 (N_7219,N_7001,N_7041);
nor U7220 (N_7220,N_7043,N_7062);
xor U7221 (N_7221,N_6917,N_6920);
or U7222 (N_7222,N_6962,N_7184);
xor U7223 (N_7223,N_7018,N_7183);
and U7224 (N_7224,N_7136,N_6995);
and U7225 (N_7225,N_7122,N_7055);
nor U7226 (N_7226,N_6918,N_7107);
nor U7227 (N_7227,N_6925,N_7199);
nor U7228 (N_7228,N_7161,N_7142);
and U7229 (N_7229,N_6979,N_7071);
and U7230 (N_7230,N_7152,N_7195);
nand U7231 (N_7231,N_7141,N_6972);
and U7232 (N_7232,N_7039,N_7068);
nor U7233 (N_7233,N_6947,N_7017);
xor U7234 (N_7234,N_7144,N_6900);
nor U7235 (N_7235,N_6932,N_7140);
nand U7236 (N_7236,N_6988,N_6946);
or U7237 (N_7237,N_6953,N_6935);
and U7238 (N_7238,N_7076,N_7100);
nor U7239 (N_7239,N_7163,N_6957);
nand U7240 (N_7240,N_7084,N_6996);
xnor U7241 (N_7241,N_6929,N_7000);
or U7242 (N_7242,N_7063,N_7083);
nand U7243 (N_7243,N_7056,N_7194);
nor U7244 (N_7244,N_7158,N_7011);
or U7245 (N_7245,N_7179,N_7174);
or U7246 (N_7246,N_7098,N_7059);
nor U7247 (N_7247,N_7162,N_6912);
or U7248 (N_7248,N_7111,N_7053);
xnor U7249 (N_7249,N_6969,N_6949);
nor U7250 (N_7250,N_7112,N_7064);
or U7251 (N_7251,N_6991,N_6938);
nor U7252 (N_7252,N_7146,N_6924);
nor U7253 (N_7253,N_7159,N_7027);
nor U7254 (N_7254,N_7135,N_7009);
xor U7255 (N_7255,N_7114,N_6994);
or U7256 (N_7256,N_6937,N_7091);
or U7257 (N_7257,N_7010,N_6982);
xnor U7258 (N_7258,N_7155,N_6983);
nand U7259 (N_7259,N_7028,N_6944);
or U7260 (N_7260,N_7128,N_7169);
nand U7261 (N_7261,N_7089,N_7145);
and U7262 (N_7262,N_7004,N_7021);
or U7263 (N_7263,N_7119,N_7175);
xor U7264 (N_7264,N_6902,N_6976);
or U7265 (N_7265,N_7192,N_7022);
nand U7266 (N_7266,N_7047,N_7052);
and U7267 (N_7267,N_7156,N_7026);
xor U7268 (N_7268,N_6986,N_6963);
and U7269 (N_7269,N_6934,N_7077);
or U7270 (N_7270,N_7096,N_6999);
and U7271 (N_7271,N_7105,N_6942);
xnor U7272 (N_7272,N_7036,N_6973);
xor U7273 (N_7273,N_7067,N_6915);
nor U7274 (N_7274,N_7045,N_7178);
and U7275 (N_7275,N_6980,N_6968);
nand U7276 (N_7276,N_7153,N_6910);
nand U7277 (N_7277,N_6914,N_7037);
and U7278 (N_7278,N_7171,N_7108);
or U7279 (N_7279,N_7165,N_7177);
and U7280 (N_7280,N_7167,N_7097);
xor U7281 (N_7281,N_6911,N_6940);
xnor U7282 (N_7282,N_7181,N_6984);
or U7283 (N_7283,N_7005,N_7170);
xor U7284 (N_7284,N_7090,N_7166);
and U7285 (N_7285,N_6974,N_6959);
nor U7286 (N_7286,N_7030,N_6981);
nor U7287 (N_7287,N_7006,N_6989);
xor U7288 (N_7288,N_7121,N_7132);
nor U7289 (N_7289,N_7193,N_6958);
or U7290 (N_7290,N_7014,N_6954);
and U7291 (N_7291,N_7172,N_7032);
xor U7292 (N_7292,N_7117,N_7176);
nand U7293 (N_7293,N_6970,N_7131);
and U7294 (N_7294,N_7033,N_7024);
nand U7295 (N_7295,N_6907,N_6952);
or U7296 (N_7296,N_6926,N_6928);
nor U7297 (N_7297,N_7057,N_6939);
nand U7298 (N_7298,N_7106,N_7099);
nor U7299 (N_7299,N_7125,N_7087);
or U7300 (N_7300,N_6901,N_7025);
and U7301 (N_7301,N_6956,N_7020);
nand U7302 (N_7302,N_7129,N_7185);
xor U7303 (N_7303,N_7110,N_7134);
nand U7304 (N_7304,N_7127,N_7035);
nand U7305 (N_7305,N_7065,N_7054);
nand U7306 (N_7306,N_6985,N_7007);
and U7307 (N_7307,N_6916,N_7188);
and U7308 (N_7308,N_7046,N_7073);
nand U7309 (N_7309,N_7191,N_7115);
or U7310 (N_7310,N_7190,N_6922);
nor U7311 (N_7311,N_6966,N_7197);
or U7312 (N_7312,N_7189,N_7050);
and U7313 (N_7313,N_7002,N_7061);
nand U7314 (N_7314,N_6905,N_6997);
nand U7315 (N_7315,N_6992,N_7180);
xnor U7316 (N_7316,N_6961,N_7086);
or U7317 (N_7317,N_7044,N_7157);
xor U7318 (N_7318,N_7003,N_6945);
nor U7319 (N_7319,N_6906,N_6904);
and U7320 (N_7320,N_7079,N_6919);
nor U7321 (N_7321,N_7123,N_6943);
nor U7322 (N_7322,N_7186,N_7154);
and U7323 (N_7323,N_7104,N_6964);
nand U7324 (N_7324,N_7101,N_7023);
nor U7325 (N_7325,N_7019,N_6998);
or U7326 (N_7326,N_6967,N_7034);
nor U7327 (N_7327,N_7130,N_7069);
xnor U7328 (N_7328,N_6909,N_7149);
nand U7329 (N_7329,N_6903,N_7113);
xor U7330 (N_7330,N_6977,N_6987);
and U7331 (N_7331,N_7008,N_6933);
nand U7332 (N_7332,N_7040,N_6990);
nand U7333 (N_7333,N_7051,N_7118);
nand U7334 (N_7334,N_6978,N_7151);
nor U7335 (N_7335,N_6908,N_7173);
nand U7336 (N_7336,N_7078,N_7075);
nand U7337 (N_7337,N_7094,N_6931);
or U7338 (N_7338,N_6941,N_7103);
and U7339 (N_7339,N_6923,N_7060);
nand U7340 (N_7340,N_7080,N_7139);
xnor U7341 (N_7341,N_7120,N_7029);
nand U7342 (N_7342,N_6921,N_7038);
xnor U7343 (N_7343,N_7126,N_6913);
nand U7344 (N_7344,N_7116,N_7048);
or U7345 (N_7345,N_7058,N_7042);
and U7346 (N_7346,N_7093,N_7168);
nand U7347 (N_7347,N_7102,N_7074);
nor U7348 (N_7348,N_7092,N_7124);
nor U7349 (N_7349,N_6993,N_7198);
and U7350 (N_7350,N_7098,N_7108);
nor U7351 (N_7351,N_7182,N_7125);
and U7352 (N_7352,N_7117,N_7151);
nand U7353 (N_7353,N_6947,N_7106);
nor U7354 (N_7354,N_7115,N_7095);
or U7355 (N_7355,N_6969,N_7141);
xor U7356 (N_7356,N_7102,N_7046);
and U7357 (N_7357,N_7046,N_7004);
nand U7358 (N_7358,N_6954,N_7067);
or U7359 (N_7359,N_7169,N_6986);
nor U7360 (N_7360,N_7089,N_6934);
or U7361 (N_7361,N_7163,N_7031);
xor U7362 (N_7362,N_6979,N_7134);
and U7363 (N_7363,N_7106,N_7031);
nor U7364 (N_7364,N_7047,N_7046);
and U7365 (N_7365,N_6941,N_7095);
nor U7366 (N_7366,N_7035,N_7120);
and U7367 (N_7367,N_6948,N_7157);
xnor U7368 (N_7368,N_7145,N_7024);
and U7369 (N_7369,N_7100,N_7044);
or U7370 (N_7370,N_6950,N_7095);
or U7371 (N_7371,N_7064,N_6935);
nand U7372 (N_7372,N_7076,N_6950);
or U7373 (N_7373,N_7104,N_6977);
nor U7374 (N_7374,N_7028,N_7010);
and U7375 (N_7375,N_6933,N_6970);
xnor U7376 (N_7376,N_7139,N_7025);
xnor U7377 (N_7377,N_6965,N_6966);
xnor U7378 (N_7378,N_6922,N_7131);
nor U7379 (N_7379,N_7131,N_7030);
nor U7380 (N_7380,N_6970,N_7105);
or U7381 (N_7381,N_6944,N_7152);
and U7382 (N_7382,N_7169,N_7042);
nor U7383 (N_7383,N_7118,N_7064);
or U7384 (N_7384,N_7077,N_6932);
and U7385 (N_7385,N_6934,N_7061);
or U7386 (N_7386,N_7167,N_6971);
nand U7387 (N_7387,N_6910,N_6911);
and U7388 (N_7388,N_6971,N_7057);
xor U7389 (N_7389,N_7038,N_6940);
or U7390 (N_7390,N_7144,N_7141);
nand U7391 (N_7391,N_7133,N_7077);
xor U7392 (N_7392,N_7157,N_6992);
or U7393 (N_7393,N_7193,N_6990);
nor U7394 (N_7394,N_7120,N_7186);
or U7395 (N_7395,N_7144,N_6906);
and U7396 (N_7396,N_7146,N_7197);
nand U7397 (N_7397,N_7076,N_7031);
xor U7398 (N_7398,N_7154,N_7050);
or U7399 (N_7399,N_7184,N_7177);
xor U7400 (N_7400,N_7112,N_7086);
or U7401 (N_7401,N_7087,N_7044);
nand U7402 (N_7402,N_6934,N_7117);
xnor U7403 (N_7403,N_7023,N_7078);
xor U7404 (N_7404,N_6954,N_7123);
nor U7405 (N_7405,N_6947,N_6929);
and U7406 (N_7406,N_6965,N_6992);
nand U7407 (N_7407,N_7047,N_7149);
xnor U7408 (N_7408,N_7112,N_7084);
nand U7409 (N_7409,N_7030,N_7072);
nor U7410 (N_7410,N_7092,N_7003);
nor U7411 (N_7411,N_7037,N_6926);
or U7412 (N_7412,N_7044,N_7107);
and U7413 (N_7413,N_7127,N_7064);
and U7414 (N_7414,N_7071,N_7109);
xnor U7415 (N_7415,N_7019,N_7087);
nor U7416 (N_7416,N_7056,N_7041);
nand U7417 (N_7417,N_7007,N_6961);
or U7418 (N_7418,N_7115,N_6981);
xor U7419 (N_7419,N_6957,N_6915);
nand U7420 (N_7420,N_7003,N_7044);
nand U7421 (N_7421,N_7118,N_6979);
nor U7422 (N_7422,N_7078,N_7071);
nand U7423 (N_7423,N_7139,N_6995);
or U7424 (N_7424,N_7056,N_7148);
nand U7425 (N_7425,N_6942,N_6944);
and U7426 (N_7426,N_7158,N_6947);
nand U7427 (N_7427,N_6904,N_7021);
nand U7428 (N_7428,N_7034,N_7106);
xnor U7429 (N_7429,N_6919,N_7049);
nor U7430 (N_7430,N_7016,N_7039);
xnor U7431 (N_7431,N_7105,N_7182);
or U7432 (N_7432,N_7176,N_7155);
or U7433 (N_7433,N_7059,N_6971);
nand U7434 (N_7434,N_6937,N_7106);
and U7435 (N_7435,N_7116,N_7013);
nor U7436 (N_7436,N_6906,N_7184);
nand U7437 (N_7437,N_7057,N_7020);
xor U7438 (N_7438,N_7054,N_7007);
and U7439 (N_7439,N_7078,N_7150);
or U7440 (N_7440,N_6940,N_6918);
xnor U7441 (N_7441,N_6952,N_7083);
nand U7442 (N_7442,N_7062,N_6941);
or U7443 (N_7443,N_6927,N_7145);
or U7444 (N_7444,N_6986,N_6994);
xor U7445 (N_7445,N_7049,N_7013);
nand U7446 (N_7446,N_6979,N_7013);
or U7447 (N_7447,N_6959,N_7176);
xor U7448 (N_7448,N_7091,N_6990);
nor U7449 (N_7449,N_6984,N_7067);
xnor U7450 (N_7450,N_7009,N_6984);
nand U7451 (N_7451,N_6948,N_7093);
and U7452 (N_7452,N_7166,N_6914);
nand U7453 (N_7453,N_7020,N_7027);
nor U7454 (N_7454,N_7003,N_7014);
and U7455 (N_7455,N_6990,N_6914);
or U7456 (N_7456,N_7109,N_6920);
xnor U7457 (N_7457,N_7045,N_7100);
nor U7458 (N_7458,N_7036,N_7162);
nand U7459 (N_7459,N_7153,N_6902);
nor U7460 (N_7460,N_6972,N_7077);
xor U7461 (N_7461,N_6958,N_6991);
nand U7462 (N_7462,N_6986,N_6959);
xnor U7463 (N_7463,N_7120,N_6944);
or U7464 (N_7464,N_7002,N_7146);
and U7465 (N_7465,N_7135,N_7088);
and U7466 (N_7466,N_7132,N_7191);
nand U7467 (N_7467,N_7098,N_7069);
nand U7468 (N_7468,N_7195,N_6946);
nand U7469 (N_7469,N_6947,N_6982);
and U7470 (N_7470,N_7155,N_7008);
and U7471 (N_7471,N_6918,N_6904);
nor U7472 (N_7472,N_7196,N_7169);
and U7473 (N_7473,N_7104,N_7073);
xnor U7474 (N_7474,N_7050,N_6991);
or U7475 (N_7475,N_7194,N_7161);
nor U7476 (N_7476,N_6962,N_7105);
or U7477 (N_7477,N_7156,N_7115);
nand U7478 (N_7478,N_7073,N_7053);
nand U7479 (N_7479,N_6929,N_7082);
and U7480 (N_7480,N_6936,N_7044);
and U7481 (N_7481,N_7008,N_7107);
or U7482 (N_7482,N_7092,N_7138);
xnor U7483 (N_7483,N_7184,N_7123);
or U7484 (N_7484,N_6913,N_7030);
nor U7485 (N_7485,N_7177,N_6983);
xnor U7486 (N_7486,N_7054,N_7173);
nor U7487 (N_7487,N_7177,N_7099);
xnor U7488 (N_7488,N_7158,N_6989);
and U7489 (N_7489,N_7167,N_7127);
or U7490 (N_7490,N_7156,N_7197);
or U7491 (N_7491,N_6923,N_6948);
and U7492 (N_7492,N_7020,N_7078);
nor U7493 (N_7493,N_7169,N_7142);
nand U7494 (N_7494,N_7078,N_7096);
or U7495 (N_7495,N_7051,N_7155);
xnor U7496 (N_7496,N_7032,N_7175);
or U7497 (N_7497,N_7006,N_7020);
xnor U7498 (N_7498,N_6920,N_7090);
or U7499 (N_7499,N_7006,N_6996);
nand U7500 (N_7500,N_7204,N_7216);
nor U7501 (N_7501,N_7415,N_7213);
or U7502 (N_7502,N_7264,N_7481);
nand U7503 (N_7503,N_7348,N_7324);
xor U7504 (N_7504,N_7321,N_7482);
nor U7505 (N_7505,N_7443,N_7398);
or U7506 (N_7506,N_7233,N_7267);
nand U7507 (N_7507,N_7352,N_7360);
nor U7508 (N_7508,N_7230,N_7445);
nor U7509 (N_7509,N_7359,N_7364);
nand U7510 (N_7510,N_7435,N_7205);
nand U7511 (N_7511,N_7470,N_7257);
or U7512 (N_7512,N_7417,N_7382);
nand U7513 (N_7513,N_7355,N_7212);
nor U7514 (N_7514,N_7473,N_7336);
and U7515 (N_7515,N_7368,N_7312);
nor U7516 (N_7516,N_7416,N_7296);
or U7517 (N_7517,N_7349,N_7342);
xnor U7518 (N_7518,N_7392,N_7428);
xor U7519 (N_7519,N_7270,N_7381);
and U7520 (N_7520,N_7278,N_7406);
nand U7521 (N_7521,N_7479,N_7219);
nand U7522 (N_7522,N_7241,N_7492);
and U7523 (N_7523,N_7444,N_7434);
or U7524 (N_7524,N_7346,N_7301);
or U7525 (N_7525,N_7494,N_7248);
or U7526 (N_7526,N_7291,N_7283);
xor U7527 (N_7527,N_7439,N_7207);
and U7528 (N_7528,N_7497,N_7314);
nor U7529 (N_7529,N_7335,N_7455);
or U7530 (N_7530,N_7407,N_7351);
nand U7531 (N_7531,N_7225,N_7452);
xor U7532 (N_7532,N_7220,N_7269);
and U7533 (N_7533,N_7467,N_7401);
or U7534 (N_7534,N_7478,N_7440);
nand U7535 (N_7535,N_7320,N_7286);
nor U7536 (N_7536,N_7464,N_7474);
xor U7537 (N_7537,N_7246,N_7350);
or U7538 (N_7538,N_7400,N_7394);
nand U7539 (N_7539,N_7299,N_7463);
or U7540 (N_7540,N_7326,N_7268);
nor U7541 (N_7541,N_7211,N_7332);
nand U7542 (N_7542,N_7458,N_7449);
and U7543 (N_7543,N_7448,N_7423);
or U7544 (N_7544,N_7275,N_7472);
xor U7545 (N_7545,N_7466,N_7262);
or U7546 (N_7546,N_7384,N_7421);
nand U7547 (N_7547,N_7461,N_7403);
nor U7548 (N_7548,N_7387,N_7397);
and U7549 (N_7549,N_7243,N_7316);
or U7550 (N_7550,N_7453,N_7480);
xor U7551 (N_7551,N_7433,N_7311);
nand U7552 (N_7552,N_7234,N_7344);
nor U7553 (N_7553,N_7347,N_7222);
nand U7554 (N_7554,N_7391,N_7446);
xor U7555 (N_7555,N_7410,N_7411);
or U7556 (N_7556,N_7413,N_7253);
xor U7557 (N_7557,N_7318,N_7329);
xnor U7558 (N_7558,N_7343,N_7483);
and U7559 (N_7559,N_7367,N_7215);
xor U7560 (N_7560,N_7274,N_7208);
xor U7561 (N_7561,N_7288,N_7294);
or U7562 (N_7562,N_7227,N_7265);
xor U7563 (N_7563,N_7255,N_7424);
and U7564 (N_7564,N_7441,N_7425);
nand U7565 (N_7565,N_7371,N_7297);
nand U7566 (N_7566,N_7475,N_7366);
and U7567 (N_7567,N_7432,N_7457);
nand U7568 (N_7568,N_7447,N_7229);
nor U7569 (N_7569,N_7325,N_7237);
xor U7570 (N_7570,N_7361,N_7450);
xnor U7571 (N_7571,N_7295,N_7405);
xor U7572 (N_7572,N_7256,N_7362);
nor U7573 (N_7573,N_7385,N_7244);
nor U7574 (N_7574,N_7249,N_7322);
nor U7575 (N_7575,N_7284,N_7462);
or U7576 (N_7576,N_7380,N_7330);
or U7577 (N_7577,N_7307,N_7427);
or U7578 (N_7578,N_7389,N_7395);
xnor U7579 (N_7579,N_7372,N_7293);
nand U7580 (N_7580,N_7327,N_7402);
or U7581 (N_7581,N_7436,N_7370);
nand U7582 (N_7582,N_7471,N_7261);
nor U7583 (N_7583,N_7430,N_7390);
nand U7584 (N_7584,N_7438,N_7363);
nor U7585 (N_7585,N_7437,N_7309);
and U7586 (N_7586,N_7442,N_7236);
and U7587 (N_7587,N_7418,N_7328);
nand U7588 (N_7588,N_7337,N_7282);
nor U7589 (N_7589,N_7456,N_7218);
xor U7590 (N_7590,N_7254,N_7460);
and U7591 (N_7591,N_7409,N_7266);
nor U7592 (N_7592,N_7383,N_7221);
nor U7593 (N_7593,N_7200,N_7375);
nand U7594 (N_7594,N_7224,N_7228);
or U7595 (N_7595,N_7341,N_7426);
nor U7596 (N_7596,N_7491,N_7245);
xor U7597 (N_7597,N_7388,N_7276);
xnor U7598 (N_7598,N_7356,N_7468);
xnor U7599 (N_7599,N_7242,N_7223);
and U7600 (N_7600,N_7238,N_7280);
xor U7601 (N_7601,N_7313,N_7499);
and U7602 (N_7602,N_7232,N_7451);
nor U7603 (N_7603,N_7376,N_7374);
or U7604 (N_7604,N_7203,N_7323);
nor U7605 (N_7605,N_7305,N_7429);
nand U7606 (N_7606,N_7334,N_7226);
nand U7607 (N_7607,N_7214,N_7217);
nand U7608 (N_7608,N_7495,N_7490);
nor U7609 (N_7609,N_7298,N_7231);
or U7610 (N_7610,N_7292,N_7303);
nor U7611 (N_7611,N_7302,N_7210);
nor U7612 (N_7612,N_7431,N_7206);
and U7613 (N_7613,N_7252,N_7496);
nand U7614 (N_7614,N_7250,N_7202);
and U7615 (N_7615,N_7369,N_7289);
xor U7616 (N_7616,N_7251,N_7340);
or U7617 (N_7617,N_7279,N_7477);
and U7618 (N_7618,N_7285,N_7358);
or U7619 (N_7619,N_7393,N_7239);
or U7620 (N_7620,N_7454,N_7317);
and U7621 (N_7621,N_7396,N_7271);
or U7622 (N_7622,N_7408,N_7308);
nor U7623 (N_7623,N_7287,N_7290);
or U7624 (N_7624,N_7498,N_7319);
or U7625 (N_7625,N_7404,N_7306);
or U7626 (N_7626,N_7260,N_7488);
or U7627 (N_7627,N_7304,N_7459);
nand U7628 (N_7628,N_7414,N_7378);
xnor U7629 (N_7629,N_7331,N_7273);
nor U7630 (N_7630,N_7365,N_7399);
or U7631 (N_7631,N_7373,N_7333);
xor U7632 (N_7632,N_7485,N_7339);
and U7633 (N_7633,N_7486,N_7422);
and U7634 (N_7634,N_7353,N_7300);
nand U7635 (N_7635,N_7345,N_7386);
xnor U7636 (N_7636,N_7310,N_7209);
and U7637 (N_7637,N_7281,N_7419);
or U7638 (N_7638,N_7379,N_7420);
nor U7639 (N_7639,N_7263,N_7201);
and U7640 (N_7640,N_7258,N_7259);
xor U7641 (N_7641,N_7489,N_7465);
nor U7642 (N_7642,N_7476,N_7357);
nor U7643 (N_7643,N_7377,N_7493);
and U7644 (N_7644,N_7240,N_7469);
or U7645 (N_7645,N_7315,N_7338);
xor U7646 (N_7646,N_7235,N_7247);
or U7647 (N_7647,N_7412,N_7487);
nor U7648 (N_7648,N_7484,N_7272);
xnor U7649 (N_7649,N_7277,N_7354);
nand U7650 (N_7650,N_7296,N_7479);
nor U7651 (N_7651,N_7438,N_7269);
xnor U7652 (N_7652,N_7209,N_7265);
and U7653 (N_7653,N_7463,N_7284);
xor U7654 (N_7654,N_7320,N_7441);
and U7655 (N_7655,N_7455,N_7203);
or U7656 (N_7656,N_7228,N_7218);
xor U7657 (N_7657,N_7219,N_7271);
and U7658 (N_7658,N_7272,N_7357);
nand U7659 (N_7659,N_7281,N_7368);
xnor U7660 (N_7660,N_7427,N_7308);
nor U7661 (N_7661,N_7478,N_7242);
and U7662 (N_7662,N_7274,N_7229);
nor U7663 (N_7663,N_7437,N_7482);
nand U7664 (N_7664,N_7453,N_7398);
xnor U7665 (N_7665,N_7477,N_7479);
xor U7666 (N_7666,N_7357,N_7322);
xnor U7667 (N_7667,N_7317,N_7312);
nor U7668 (N_7668,N_7487,N_7498);
or U7669 (N_7669,N_7215,N_7457);
xor U7670 (N_7670,N_7216,N_7238);
nor U7671 (N_7671,N_7365,N_7466);
or U7672 (N_7672,N_7491,N_7401);
and U7673 (N_7673,N_7338,N_7340);
and U7674 (N_7674,N_7422,N_7207);
xnor U7675 (N_7675,N_7452,N_7434);
nor U7676 (N_7676,N_7219,N_7487);
and U7677 (N_7677,N_7431,N_7314);
or U7678 (N_7678,N_7420,N_7261);
and U7679 (N_7679,N_7367,N_7247);
and U7680 (N_7680,N_7471,N_7316);
nor U7681 (N_7681,N_7423,N_7306);
nor U7682 (N_7682,N_7416,N_7439);
or U7683 (N_7683,N_7498,N_7216);
nor U7684 (N_7684,N_7491,N_7246);
and U7685 (N_7685,N_7232,N_7273);
nor U7686 (N_7686,N_7448,N_7417);
nor U7687 (N_7687,N_7405,N_7360);
and U7688 (N_7688,N_7346,N_7379);
or U7689 (N_7689,N_7381,N_7401);
nor U7690 (N_7690,N_7392,N_7453);
nand U7691 (N_7691,N_7350,N_7318);
or U7692 (N_7692,N_7408,N_7311);
nand U7693 (N_7693,N_7292,N_7204);
xor U7694 (N_7694,N_7481,N_7388);
and U7695 (N_7695,N_7337,N_7256);
nand U7696 (N_7696,N_7406,N_7253);
or U7697 (N_7697,N_7232,N_7348);
nand U7698 (N_7698,N_7265,N_7404);
nor U7699 (N_7699,N_7476,N_7496);
and U7700 (N_7700,N_7357,N_7233);
or U7701 (N_7701,N_7367,N_7489);
nand U7702 (N_7702,N_7404,N_7323);
and U7703 (N_7703,N_7498,N_7326);
xor U7704 (N_7704,N_7285,N_7240);
nor U7705 (N_7705,N_7209,N_7255);
nand U7706 (N_7706,N_7392,N_7246);
xnor U7707 (N_7707,N_7214,N_7240);
xor U7708 (N_7708,N_7264,N_7497);
xnor U7709 (N_7709,N_7305,N_7251);
or U7710 (N_7710,N_7290,N_7390);
or U7711 (N_7711,N_7459,N_7402);
xor U7712 (N_7712,N_7332,N_7419);
nand U7713 (N_7713,N_7450,N_7433);
nand U7714 (N_7714,N_7253,N_7487);
xnor U7715 (N_7715,N_7288,N_7411);
xor U7716 (N_7716,N_7235,N_7292);
nor U7717 (N_7717,N_7464,N_7452);
xor U7718 (N_7718,N_7359,N_7319);
xnor U7719 (N_7719,N_7275,N_7252);
nand U7720 (N_7720,N_7359,N_7310);
and U7721 (N_7721,N_7441,N_7498);
or U7722 (N_7722,N_7275,N_7298);
nand U7723 (N_7723,N_7410,N_7481);
nand U7724 (N_7724,N_7296,N_7366);
nand U7725 (N_7725,N_7480,N_7435);
and U7726 (N_7726,N_7249,N_7492);
nor U7727 (N_7727,N_7212,N_7406);
or U7728 (N_7728,N_7415,N_7270);
nor U7729 (N_7729,N_7376,N_7281);
or U7730 (N_7730,N_7202,N_7205);
xnor U7731 (N_7731,N_7353,N_7410);
nor U7732 (N_7732,N_7291,N_7269);
nor U7733 (N_7733,N_7414,N_7244);
nor U7734 (N_7734,N_7415,N_7212);
and U7735 (N_7735,N_7415,N_7377);
or U7736 (N_7736,N_7365,N_7464);
xor U7737 (N_7737,N_7266,N_7230);
and U7738 (N_7738,N_7200,N_7266);
and U7739 (N_7739,N_7402,N_7332);
nor U7740 (N_7740,N_7314,N_7398);
nor U7741 (N_7741,N_7478,N_7348);
and U7742 (N_7742,N_7338,N_7375);
xnor U7743 (N_7743,N_7282,N_7407);
or U7744 (N_7744,N_7221,N_7404);
and U7745 (N_7745,N_7287,N_7369);
nand U7746 (N_7746,N_7284,N_7352);
nand U7747 (N_7747,N_7394,N_7309);
xor U7748 (N_7748,N_7241,N_7248);
or U7749 (N_7749,N_7353,N_7366);
or U7750 (N_7750,N_7201,N_7419);
or U7751 (N_7751,N_7206,N_7251);
nor U7752 (N_7752,N_7390,N_7409);
nand U7753 (N_7753,N_7246,N_7463);
or U7754 (N_7754,N_7499,N_7485);
nand U7755 (N_7755,N_7297,N_7357);
xnor U7756 (N_7756,N_7385,N_7261);
and U7757 (N_7757,N_7200,N_7440);
nand U7758 (N_7758,N_7423,N_7477);
or U7759 (N_7759,N_7484,N_7219);
and U7760 (N_7760,N_7304,N_7332);
nand U7761 (N_7761,N_7478,N_7295);
nand U7762 (N_7762,N_7243,N_7300);
or U7763 (N_7763,N_7489,N_7202);
and U7764 (N_7764,N_7338,N_7471);
and U7765 (N_7765,N_7218,N_7460);
nand U7766 (N_7766,N_7468,N_7218);
or U7767 (N_7767,N_7461,N_7204);
nor U7768 (N_7768,N_7431,N_7428);
xnor U7769 (N_7769,N_7243,N_7202);
nor U7770 (N_7770,N_7294,N_7230);
or U7771 (N_7771,N_7368,N_7389);
nand U7772 (N_7772,N_7333,N_7401);
nor U7773 (N_7773,N_7308,N_7434);
or U7774 (N_7774,N_7478,N_7256);
nor U7775 (N_7775,N_7468,N_7368);
and U7776 (N_7776,N_7352,N_7426);
or U7777 (N_7777,N_7401,N_7497);
or U7778 (N_7778,N_7316,N_7313);
nor U7779 (N_7779,N_7215,N_7404);
and U7780 (N_7780,N_7230,N_7429);
and U7781 (N_7781,N_7339,N_7343);
and U7782 (N_7782,N_7227,N_7279);
nand U7783 (N_7783,N_7261,N_7321);
nor U7784 (N_7784,N_7303,N_7224);
nor U7785 (N_7785,N_7339,N_7299);
or U7786 (N_7786,N_7332,N_7479);
nor U7787 (N_7787,N_7424,N_7267);
nor U7788 (N_7788,N_7383,N_7436);
nand U7789 (N_7789,N_7205,N_7326);
or U7790 (N_7790,N_7266,N_7436);
or U7791 (N_7791,N_7410,N_7380);
nor U7792 (N_7792,N_7229,N_7314);
and U7793 (N_7793,N_7414,N_7495);
and U7794 (N_7794,N_7334,N_7224);
or U7795 (N_7795,N_7323,N_7223);
nor U7796 (N_7796,N_7442,N_7344);
nand U7797 (N_7797,N_7482,N_7449);
nor U7798 (N_7798,N_7406,N_7312);
or U7799 (N_7799,N_7327,N_7246);
nand U7800 (N_7800,N_7658,N_7528);
and U7801 (N_7801,N_7695,N_7586);
nor U7802 (N_7802,N_7607,N_7591);
nor U7803 (N_7803,N_7652,N_7505);
nor U7804 (N_7804,N_7768,N_7545);
nand U7805 (N_7805,N_7654,N_7688);
and U7806 (N_7806,N_7677,N_7726);
xnor U7807 (N_7807,N_7585,N_7571);
nand U7808 (N_7808,N_7736,N_7553);
and U7809 (N_7809,N_7763,N_7567);
nor U7810 (N_7810,N_7708,N_7753);
and U7811 (N_7811,N_7539,N_7700);
nand U7812 (N_7812,N_7744,N_7582);
and U7813 (N_7813,N_7734,N_7631);
nand U7814 (N_7814,N_7541,N_7748);
or U7815 (N_7815,N_7699,N_7727);
xor U7816 (N_7816,N_7751,N_7657);
nand U7817 (N_7817,N_7504,N_7502);
or U7818 (N_7818,N_7540,N_7686);
nor U7819 (N_7819,N_7555,N_7612);
nor U7820 (N_7820,N_7756,N_7564);
xnor U7821 (N_7821,N_7627,N_7730);
and U7822 (N_7822,N_7630,N_7575);
xor U7823 (N_7823,N_7565,N_7617);
xnor U7824 (N_7824,N_7573,N_7587);
or U7825 (N_7825,N_7570,N_7723);
or U7826 (N_7826,N_7624,N_7637);
or U7827 (N_7827,N_7517,N_7603);
xor U7828 (N_7828,N_7622,N_7684);
nand U7829 (N_7829,N_7589,N_7534);
nor U7830 (N_7830,N_7619,N_7641);
nand U7831 (N_7831,N_7568,N_7712);
nor U7832 (N_7832,N_7635,N_7715);
xor U7833 (N_7833,N_7665,N_7507);
nand U7834 (N_7834,N_7662,N_7719);
and U7835 (N_7835,N_7560,N_7602);
xnor U7836 (N_7836,N_7610,N_7704);
nor U7837 (N_7837,N_7594,N_7551);
nand U7838 (N_7838,N_7669,N_7673);
or U7839 (N_7839,N_7664,N_7605);
and U7840 (N_7840,N_7767,N_7533);
xor U7841 (N_7841,N_7514,N_7724);
nand U7842 (N_7842,N_7638,N_7552);
and U7843 (N_7843,N_7739,N_7549);
or U7844 (N_7844,N_7584,N_7609);
or U7845 (N_7845,N_7762,N_7623);
nand U7846 (N_7846,N_7738,N_7659);
or U7847 (N_7847,N_7546,N_7765);
nand U7848 (N_7848,N_7663,N_7554);
nand U7849 (N_7849,N_7784,N_7590);
nor U7850 (N_7850,N_7707,N_7774);
xnor U7851 (N_7851,N_7548,N_7794);
or U7852 (N_7852,N_7697,N_7524);
or U7853 (N_7853,N_7769,N_7601);
and U7854 (N_7854,N_7614,N_7515);
xor U7855 (N_7855,N_7785,N_7773);
xor U7856 (N_7856,N_7574,N_7720);
and U7857 (N_7857,N_7562,N_7593);
nand U7858 (N_7858,N_7701,N_7639);
xnor U7859 (N_7859,N_7705,N_7579);
and U7860 (N_7860,N_7675,N_7692);
nand U7861 (N_7861,N_7625,N_7761);
xnor U7862 (N_7862,N_7752,N_7655);
and U7863 (N_7863,N_7728,N_7690);
nand U7864 (N_7864,N_7772,N_7796);
nand U7865 (N_7865,N_7522,N_7656);
and U7866 (N_7866,N_7759,N_7706);
xnor U7867 (N_7867,N_7710,N_7757);
nand U7868 (N_7868,N_7680,N_7709);
and U7869 (N_7869,N_7577,N_7501);
and U7870 (N_7870,N_7732,N_7521);
and U7871 (N_7871,N_7543,N_7640);
and U7872 (N_7872,N_7779,N_7559);
xnor U7873 (N_7873,N_7508,N_7535);
nand U7874 (N_7874,N_7671,N_7556);
and U7875 (N_7875,N_7745,N_7506);
or U7876 (N_7876,N_7681,N_7691);
nor U7877 (N_7877,N_7667,N_7511);
or U7878 (N_7878,N_7626,N_7679);
nand U7879 (N_7879,N_7721,N_7797);
nand U7880 (N_7880,N_7740,N_7725);
or U7881 (N_7881,N_7606,N_7520);
xnor U7882 (N_7882,N_7799,N_7592);
or U7883 (N_7883,N_7608,N_7743);
nor U7884 (N_7884,N_7718,N_7503);
xor U7885 (N_7885,N_7758,N_7683);
xor U7886 (N_7886,N_7621,N_7578);
nor U7887 (N_7887,N_7580,N_7531);
xor U7888 (N_7888,N_7500,N_7661);
and U7889 (N_7889,N_7597,N_7651);
xor U7890 (N_7890,N_7764,N_7616);
or U7891 (N_7891,N_7569,N_7563);
nand U7892 (N_7892,N_7791,N_7648);
and U7893 (N_7893,N_7643,N_7711);
nand U7894 (N_7894,N_7780,N_7537);
xor U7895 (N_7895,N_7509,N_7678);
nand U7896 (N_7896,N_7754,N_7512);
nand U7897 (N_7897,N_7600,N_7628);
nor U7898 (N_7898,N_7786,N_7733);
xnor U7899 (N_7899,N_7787,N_7523);
nand U7900 (N_7900,N_7530,N_7689);
nand U7901 (N_7901,N_7532,N_7583);
and U7902 (N_7902,N_7650,N_7510);
nor U7903 (N_7903,N_7790,N_7760);
xnor U7904 (N_7904,N_7777,N_7588);
xnor U7905 (N_7905,N_7750,N_7742);
xor U7906 (N_7906,N_7735,N_7703);
nand U7907 (N_7907,N_7649,N_7566);
or U7908 (N_7908,N_7518,N_7766);
nor U7909 (N_7909,N_7526,N_7698);
nor U7910 (N_7910,N_7629,N_7516);
and U7911 (N_7911,N_7618,N_7519);
and U7912 (N_7912,N_7694,N_7581);
or U7913 (N_7913,N_7666,N_7645);
nand U7914 (N_7914,N_7653,N_7778);
xnor U7915 (N_7915,N_7672,N_7731);
nor U7916 (N_7916,N_7741,N_7714);
xnor U7917 (N_7917,N_7550,N_7636);
and U7918 (N_7918,N_7749,N_7702);
and U7919 (N_7919,N_7644,N_7604);
xnor U7920 (N_7920,N_7722,N_7685);
nor U7921 (N_7921,N_7642,N_7632);
nor U7922 (N_7922,N_7538,N_7696);
nand U7923 (N_7923,N_7781,N_7668);
nor U7924 (N_7924,N_7674,N_7717);
and U7925 (N_7925,N_7634,N_7670);
nor U7926 (N_7926,N_7792,N_7798);
nand U7927 (N_7927,N_7687,N_7558);
nand U7928 (N_7928,N_7793,N_7783);
and U7929 (N_7929,N_7788,N_7789);
nor U7930 (N_7930,N_7755,N_7770);
nand U7931 (N_7931,N_7795,N_7572);
and U7932 (N_7932,N_7525,N_7747);
or U7933 (N_7933,N_7536,N_7529);
or U7934 (N_7934,N_7716,N_7682);
nor U7935 (N_7935,N_7633,N_7729);
and U7936 (N_7936,N_7782,N_7776);
xor U7937 (N_7937,N_7746,N_7542);
and U7938 (N_7938,N_7620,N_7646);
xor U7939 (N_7939,N_7775,N_7547);
and U7940 (N_7940,N_7576,N_7595);
and U7941 (N_7941,N_7557,N_7771);
or U7942 (N_7942,N_7596,N_7737);
and U7943 (N_7943,N_7599,N_7693);
and U7944 (N_7944,N_7676,N_7544);
or U7945 (N_7945,N_7611,N_7527);
nand U7946 (N_7946,N_7713,N_7615);
or U7947 (N_7947,N_7598,N_7660);
and U7948 (N_7948,N_7647,N_7561);
nor U7949 (N_7949,N_7613,N_7513);
and U7950 (N_7950,N_7616,N_7590);
or U7951 (N_7951,N_7517,N_7553);
xnor U7952 (N_7952,N_7564,N_7688);
nand U7953 (N_7953,N_7795,N_7666);
nand U7954 (N_7954,N_7605,N_7798);
nand U7955 (N_7955,N_7693,N_7668);
nand U7956 (N_7956,N_7717,N_7641);
nand U7957 (N_7957,N_7572,N_7604);
nand U7958 (N_7958,N_7693,N_7553);
nor U7959 (N_7959,N_7507,N_7721);
or U7960 (N_7960,N_7649,N_7646);
nand U7961 (N_7961,N_7613,N_7779);
nand U7962 (N_7962,N_7548,N_7739);
nand U7963 (N_7963,N_7793,N_7766);
xnor U7964 (N_7964,N_7610,N_7658);
xnor U7965 (N_7965,N_7787,N_7747);
nand U7966 (N_7966,N_7539,N_7548);
nor U7967 (N_7967,N_7798,N_7650);
or U7968 (N_7968,N_7539,N_7758);
and U7969 (N_7969,N_7611,N_7778);
nand U7970 (N_7970,N_7758,N_7767);
and U7971 (N_7971,N_7585,N_7647);
and U7972 (N_7972,N_7554,N_7551);
xor U7973 (N_7973,N_7635,N_7672);
xor U7974 (N_7974,N_7703,N_7626);
nand U7975 (N_7975,N_7615,N_7558);
xor U7976 (N_7976,N_7792,N_7583);
nand U7977 (N_7977,N_7748,N_7731);
xor U7978 (N_7978,N_7563,N_7667);
xor U7979 (N_7979,N_7783,N_7654);
nand U7980 (N_7980,N_7701,N_7605);
or U7981 (N_7981,N_7762,N_7525);
and U7982 (N_7982,N_7509,N_7599);
xnor U7983 (N_7983,N_7666,N_7698);
nand U7984 (N_7984,N_7615,N_7676);
and U7985 (N_7985,N_7767,N_7771);
nor U7986 (N_7986,N_7571,N_7747);
nor U7987 (N_7987,N_7627,N_7618);
xor U7988 (N_7988,N_7640,N_7741);
nor U7989 (N_7989,N_7561,N_7736);
xnor U7990 (N_7990,N_7538,N_7639);
nand U7991 (N_7991,N_7711,N_7722);
or U7992 (N_7992,N_7662,N_7591);
or U7993 (N_7993,N_7700,N_7659);
or U7994 (N_7994,N_7520,N_7668);
xnor U7995 (N_7995,N_7739,N_7715);
or U7996 (N_7996,N_7648,N_7516);
nand U7997 (N_7997,N_7613,N_7778);
nand U7998 (N_7998,N_7713,N_7500);
nor U7999 (N_7999,N_7752,N_7641);
xor U8000 (N_8000,N_7794,N_7694);
and U8001 (N_8001,N_7551,N_7753);
nand U8002 (N_8002,N_7614,N_7792);
xor U8003 (N_8003,N_7617,N_7721);
xor U8004 (N_8004,N_7557,N_7657);
nand U8005 (N_8005,N_7553,N_7762);
nor U8006 (N_8006,N_7768,N_7588);
and U8007 (N_8007,N_7671,N_7779);
xnor U8008 (N_8008,N_7660,N_7624);
and U8009 (N_8009,N_7662,N_7739);
nand U8010 (N_8010,N_7660,N_7683);
nor U8011 (N_8011,N_7676,N_7716);
and U8012 (N_8012,N_7676,N_7761);
or U8013 (N_8013,N_7565,N_7699);
nor U8014 (N_8014,N_7561,N_7650);
nand U8015 (N_8015,N_7582,N_7751);
nor U8016 (N_8016,N_7630,N_7544);
xor U8017 (N_8017,N_7649,N_7562);
nor U8018 (N_8018,N_7605,N_7662);
nand U8019 (N_8019,N_7648,N_7634);
or U8020 (N_8020,N_7635,N_7699);
or U8021 (N_8021,N_7517,N_7612);
and U8022 (N_8022,N_7742,N_7635);
xor U8023 (N_8023,N_7510,N_7627);
nand U8024 (N_8024,N_7684,N_7503);
xor U8025 (N_8025,N_7674,N_7579);
or U8026 (N_8026,N_7504,N_7696);
or U8027 (N_8027,N_7556,N_7635);
or U8028 (N_8028,N_7513,N_7666);
xnor U8029 (N_8029,N_7796,N_7513);
nand U8030 (N_8030,N_7725,N_7679);
or U8031 (N_8031,N_7593,N_7770);
and U8032 (N_8032,N_7731,N_7698);
xnor U8033 (N_8033,N_7743,N_7798);
nand U8034 (N_8034,N_7630,N_7747);
xnor U8035 (N_8035,N_7568,N_7547);
or U8036 (N_8036,N_7684,N_7728);
xor U8037 (N_8037,N_7559,N_7663);
xnor U8038 (N_8038,N_7774,N_7745);
xnor U8039 (N_8039,N_7505,N_7770);
or U8040 (N_8040,N_7793,N_7718);
and U8041 (N_8041,N_7660,N_7729);
and U8042 (N_8042,N_7749,N_7641);
nand U8043 (N_8043,N_7706,N_7627);
or U8044 (N_8044,N_7629,N_7759);
nand U8045 (N_8045,N_7692,N_7623);
nand U8046 (N_8046,N_7789,N_7696);
nor U8047 (N_8047,N_7583,N_7680);
nand U8048 (N_8048,N_7746,N_7591);
and U8049 (N_8049,N_7531,N_7576);
xor U8050 (N_8050,N_7525,N_7620);
nand U8051 (N_8051,N_7568,N_7609);
and U8052 (N_8052,N_7720,N_7686);
xnor U8053 (N_8053,N_7597,N_7630);
nand U8054 (N_8054,N_7595,N_7616);
nand U8055 (N_8055,N_7746,N_7709);
or U8056 (N_8056,N_7547,N_7736);
or U8057 (N_8057,N_7657,N_7586);
and U8058 (N_8058,N_7778,N_7629);
nor U8059 (N_8059,N_7657,N_7683);
and U8060 (N_8060,N_7795,N_7619);
and U8061 (N_8061,N_7674,N_7562);
nor U8062 (N_8062,N_7743,N_7689);
or U8063 (N_8063,N_7797,N_7656);
nor U8064 (N_8064,N_7786,N_7634);
xor U8065 (N_8065,N_7790,N_7606);
nor U8066 (N_8066,N_7742,N_7647);
and U8067 (N_8067,N_7506,N_7602);
and U8068 (N_8068,N_7669,N_7704);
nand U8069 (N_8069,N_7679,N_7757);
nor U8070 (N_8070,N_7681,N_7741);
nor U8071 (N_8071,N_7674,N_7651);
nand U8072 (N_8072,N_7503,N_7589);
nor U8073 (N_8073,N_7506,N_7608);
and U8074 (N_8074,N_7629,N_7628);
nand U8075 (N_8075,N_7751,N_7738);
and U8076 (N_8076,N_7743,N_7680);
or U8077 (N_8077,N_7780,N_7756);
and U8078 (N_8078,N_7791,N_7612);
nand U8079 (N_8079,N_7657,N_7503);
nor U8080 (N_8080,N_7590,N_7637);
nand U8081 (N_8081,N_7655,N_7556);
nand U8082 (N_8082,N_7660,N_7593);
xor U8083 (N_8083,N_7692,N_7662);
and U8084 (N_8084,N_7574,N_7791);
nor U8085 (N_8085,N_7736,N_7562);
nor U8086 (N_8086,N_7761,N_7750);
xnor U8087 (N_8087,N_7714,N_7736);
nor U8088 (N_8088,N_7740,N_7672);
nor U8089 (N_8089,N_7658,N_7766);
nand U8090 (N_8090,N_7516,N_7665);
or U8091 (N_8091,N_7563,N_7535);
xor U8092 (N_8092,N_7759,N_7724);
or U8093 (N_8093,N_7589,N_7736);
and U8094 (N_8094,N_7546,N_7684);
nand U8095 (N_8095,N_7757,N_7611);
or U8096 (N_8096,N_7506,N_7634);
and U8097 (N_8097,N_7585,N_7740);
nor U8098 (N_8098,N_7666,N_7769);
nand U8099 (N_8099,N_7678,N_7669);
or U8100 (N_8100,N_7920,N_7837);
nor U8101 (N_8101,N_8030,N_7975);
nand U8102 (N_8102,N_7972,N_7953);
or U8103 (N_8103,N_8071,N_8023);
xnor U8104 (N_8104,N_8099,N_7808);
nand U8105 (N_8105,N_8064,N_7862);
xnor U8106 (N_8106,N_7985,N_7951);
and U8107 (N_8107,N_8011,N_7906);
nand U8108 (N_8108,N_7804,N_8024);
nor U8109 (N_8109,N_7934,N_7829);
or U8110 (N_8110,N_8012,N_7960);
and U8111 (N_8111,N_7959,N_8045);
nand U8112 (N_8112,N_7852,N_7921);
xnor U8113 (N_8113,N_7999,N_8083);
or U8114 (N_8114,N_7922,N_8016);
nand U8115 (N_8115,N_7832,N_7865);
nand U8116 (N_8116,N_8032,N_8027);
xnor U8117 (N_8117,N_7807,N_7944);
and U8118 (N_8118,N_7954,N_7942);
xor U8119 (N_8119,N_7900,N_7925);
or U8120 (N_8120,N_8098,N_7966);
and U8121 (N_8121,N_7809,N_8088);
nor U8122 (N_8122,N_7991,N_8072);
xnor U8123 (N_8123,N_7806,N_7812);
and U8124 (N_8124,N_8006,N_7903);
nor U8125 (N_8125,N_8082,N_7969);
or U8126 (N_8126,N_7819,N_8003);
xor U8127 (N_8127,N_8002,N_8075);
nor U8128 (N_8128,N_7945,N_8037);
and U8129 (N_8129,N_7820,N_7823);
nand U8130 (N_8130,N_7917,N_8080);
or U8131 (N_8131,N_8035,N_7965);
and U8132 (N_8132,N_7834,N_8068);
nand U8133 (N_8133,N_8093,N_7963);
or U8134 (N_8134,N_7818,N_7802);
nor U8135 (N_8135,N_7997,N_7898);
nand U8136 (N_8136,N_8010,N_7842);
and U8137 (N_8137,N_8020,N_7870);
nor U8138 (N_8138,N_7844,N_7957);
or U8139 (N_8139,N_7872,N_7964);
xnor U8140 (N_8140,N_8033,N_7861);
xnor U8141 (N_8141,N_7995,N_8074);
and U8142 (N_8142,N_8041,N_7986);
xnor U8143 (N_8143,N_7883,N_7811);
nand U8144 (N_8144,N_7878,N_8013);
and U8145 (N_8145,N_7912,N_7801);
nor U8146 (N_8146,N_7843,N_7989);
xnor U8147 (N_8147,N_7887,N_7800);
nand U8148 (N_8148,N_7825,N_8061);
nor U8149 (N_8149,N_8065,N_8029);
nor U8150 (N_8150,N_8092,N_7919);
or U8151 (N_8151,N_7810,N_7877);
and U8152 (N_8152,N_7824,N_7909);
xnor U8153 (N_8153,N_8044,N_7876);
or U8154 (N_8154,N_7893,N_7853);
nand U8155 (N_8155,N_7827,N_7952);
or U8156 (N_8156,N_7973,N_7902);
or U8157 (N_8157,N_8095,N_7979);
nand U8158 (N_8158,N_7981,N_8039);
nor U8159 (N_8159,N_7990,N_7894);
nand U8160 (N_8160,N_7857,N_7996);
xor U8161 (N_8161,N_7927,N_7897);
or U8162 (N_8162,N_7821,N_7935);
or U8163 (N_8163,N_7856,N_7830);
or U8164 (N_8164,N_8026,N_8091);
xnor U8165 (N_8165,N_7905,N_7841);
xnor U8166 (N_8166,N_7815,N_8081);
xor U8167 (N_8167,N_7982,N_7978);
nand U8168 (N_8168,N_7845,N_7923);
and U8169 (N_8169,N_7936,N_7863);
xnor U8170 (N_8170,N_7881,N_8056);
xnor U8171 (N_8171,N_7871,N_7974);
nand U8172 (N_8172,N_7911,N_7910);
xor U8173 (N_8173,N_7892,N_8040);
and U8174 (N_8174,N_8051,N_7896);
or U8175 (N_8175,N_7992,N_7926);
xnor U8176 (N_8176,N_8007,N_7846);
nand U8177 (N_8177,N_8000,N_8058);
xnor U8178 (N_8178,N_8097,N_8019);
nor U8179 (N_8179,N_7895,N_8015);
and U8180 (N_8180,N_7924,N_7987);
xor U8181 (N_8181,N_7867,N_7828);
and U8182 (N_8182,N_7943,N_8014);
and U8183 (N_8183,N_7941,N_7918);
nor U8184 (N_8184,N_8052,N_7994);
nor U8185 (N_8185,N_8070,N_8085);
and U8186 (N_8186,N_7822,N_8005);
xnor U8187 (N_8187,N_7940,N_8084);
and U8188 (N_8188,N_7984,N_7916);
nand U8189 (N_8189,N_7998,N_8046);
nor U8190 (N_8190,N_7826,N_7805);
or U8191 (N_8191,N_7850,N_8059);
nor U8192 (N_8192,N_7955,N_8018);
and U8193 (N_8193,N_8009,N_7962);
or U8194 (N_8194,N_8022,N_7946);
xnor U8195 (N_8195,N_7888,N_8049);
nor U8196 (N_8196,N_7977,N_7901);
or U8197 (N_8197,N_7884,N_7869);
nor U8198 (N_8198,N_7933,N_8008);
xor U8199 (N_8199,N_8063,N_7913);
and U8200 (N_8200,N_8054,N_8057);
or U8201 (N_8201,N_7835,N_8086);
or U8202 (N_8202,N_8055,N_7950);
nor U8203 (N_8203,N_7885,N_7814);
and U8204 (N_8204,N_7854,N_7851);
or U8205 (N_8205,N_7980,N_8043);
and U8206 (N_8206,N_7803,N_7931);
and U8207 (N_8207,N_7873,N_8094);
nor U8208 (N_8208,N_7847,N_7891);
xor U8209 (N_8209,N_7929,N_8060);
and U8210 (N_8210,N_7938,N_8076);
or U8211 (N_8211,N_7840,N_8001);
and U8212 (N_8212,N_7988,N_7839);
and U8213 (N_8213,N_7813,N_8062);
nand U8214 (N_8214,N_7848,N_7855);
nor U8215 (N_8215,N_7879,N_7949);
or U8216 (N_8216,N_7915,N_7874);
xnor U8217 (N_8217,N_7866,N_7968);
and U8218 (N_8218,N_7961,N_7907);
nand U8219 (N_8219,N_8050,N_7833);
nor U8220 (N_8220,N_7817,N_7947);
or U8221 (N_8221,N_7904,N_7875);
nand U8222 (N_8222,N_8038,N_7889);
nor U8223 (N_8223,N_8047,N_8067);
and U8224 (N_8224,N_7868,N_8079);
or U8225 (N_8225,N_8028,N_8017);
nor U8226 (N_8226,N_7958,N_7993);
or U8227 (N_8227,N_8066,N_7976);
nor U8228 (N_8228,N_8036,N_7908);
nor U8229 (N_8229,N_7983,N_7948);
or U8230 (N_8230,N_7928,N_7886);
nor U8231 (N_8231,N_7939,N_7932);
nand U8232 (N_8232,N_7849,N_7882);
xnor U8233 (N_8233,N_8021,N_8077);
xor U8234 (N_8234,N_7831,N_8031);
or U8235 (N_8235,N_8096,N_7971);
nor U8236 (N_8236,N_8090,N_8034);
and U8237 (N_8237,N_7880,N_7890);
nand U8238 (N_8238,N_7899,N_7914);
or U8239 (N_8239,N_8025,N_8087);
nand U8240 (N_8240,N_7967,N_7930);
nor U8241 (N_8241,N_7838,N_7860);
nor U8242 (N_8242,N_7937,N_7970);
nand U8243 (N_8243,N_8042,N_7858);
nor U8244 (N_8244,N_7859,N_7836);
xnor U8245 (N_8245,N_8053,N_8078);
xnor U8246 (N_8246,N_7864,N_8069);
or U8247 (N_8247,N_7956,N_8048);
nand U8248 (N_8248,N_8089,N_8004);
or U8249 (N_8249,N_8073,N_7816);
xnor U8250 (N_8250,N_7809,N_8034);
and U8251 (N_8251,N_7969,N_7822);
and U8252 (N_8252,N_7838,N_7954);
nand U8253 (N_8253,N_7937,N_8017);
nor U8254 (N_8254,N_8053,N_8075);
nand U8255 (N_8255,N_8037,N_8028);
and U8256 (N_8256,N_7922,N_7838);
nand U8257 (N_8257,N_7977,N_7898);
nand U8258 (N_8258,N_7853,N_7993);
nand U8259 (N_8259,N_8023,N_7928);
nand U8260 (N_8260,N_7994,N_7896);
nor U8261 (N_8261,N_7902,N_8008);
nor U8262 (N_8262,N_8061,N_8097);
xnor U8263 (N_8263,N_7847,N_7954);
nor U8264 (N_8264,N_7835,N_7953);
or U8265 (N_8265,N_7823,N_7937);
xnor U8266 (N_8266,N_8010,N_7936);
nand U8267 (N_8267,N_7906,N_7874);
or U8268 (N_8268,N_8063,N_7807);
or U8269 (N_8269,N_8016,N_7834);
xnor U8270 (N_8270,N_7891,N_8040);
xnor U8271 (N_8271,N_8040,N_7934);
nand U8272 (N_8272,N_7923,N_7906);
or U8273 (N_8273,N_8066,N_7929);
nand U8274 (N_8274,N_7856,N_7917);
and U8275 (N_8275,N_7930,N_7999);
xnor U8276 (N_8276,N_7904,N_8045);
or U8277 (N_8277,N_8036,N_7812);
and U8278 (N_8278,N_7945,N_8073);
nand U8279 (N_8279,N_8012,N_7818);
and U8280 (N_8280,N_7920,N_7877);
nand U8281 (N_8281,N_7813,N_7822);
xnor U8282 (N_8282,N_7864,N_8011);
nand U8283 (N_8283,N_7805,N_8009);
or U8284 (N_8284,N_8020,N_7951);
and U8285 (N_8285,N_7830,N_7872);
and U8286 (N_8286,N_7989,N_8093);
or U8287 (N_8287,N_7849,N_8010);
nand U8288 (N_8288,N_8091,N_8037);
and U8289 (N_8289,N_8073,N_7967);
xor U8290 (N_8290,N_7842,N_7937);
nand U8291 (N_8291,N_7902,N_7932);
xor U8292 (N_8292,N_8077,N_8063);
or U8293 (N_8293,N_8080,N_8015);
and U8294 (N_8294,N_8003,N_8007);
nand U8295 (N_8295,N_7865,N_7956);
and U8296 (N_8296,N_7888,N_8022);
nor U8297 (N_8297,N_7990,N_7806);
and U8298 (N_8298,N_7831,N_7958);
nand U8299 (N_8299,N_7934,N_7816);
nand U8300 (N_8300,N_8013,N_8059);
and U8301 (N_8301,N_7881,N_7933);
xnor U8302 (N_8302,N_7927,N_7815);
nand U8303 (N_8303,N_7921,N_7968);
or U8304 (N_8304,N_8055,N_7912);
and U8305 (N_8305,N_8060,N_8096);
nor U8306 (N_8306,N_7962,N_7971);
xor U8307 (N_8307,N_8068,N_8012);
nor U8308 (N_8308,N_8080,N_7832);
nand U8309 (N_8309,N_7997,N_8077);
nor U8310 (N_8310,N_8047,N_8007);
nor U8311 (N_8311,N_7988,N_7929);
nand U8312 (N_8312,N_7971,N_8061);
nand U8313 (N_8313,N_7992,N_7889);
nand U8314 (N_8314,N_7890,N_7963);
nand U8315 (N_8315,N_7894,N_8093);
nand U8316 (N_8316,N_8066,N_7844);
or U8317 (N_8317,N_8002,N_7982);
nand U8318 (N_8318,N_7995,N_7845);
nand U8319 (N_8319,N_7825,N_7939);
or U8320 (N_8320,N_7960,N_7952);
nand U8321 (N_8321,N_8056,N_7807);
or U8322 (N_8322,N_7823,N_8030);
nand U8323 (N_8323,N_8003,N_7991);
nor U8324 (N_8324,N_8078,N_7922);
and U8325 (N_8325,N_7846,N_8008);
or U8326 (N_8326,N_8011,N_8031);
or U8327 (N_8327,N_7980,N_7825);
xnor U8328 (N_8328,N_7886,N_8046);
nand U8329 (N_8329,N_8075,N_7878);
and U8330 (N_8330,N_7808,N_7975);
nor U8331 (N_8331,N_7977,N_7864);
xnor U8332 (N_8332,N_8081,N_7976);
nor U8333 (N_8333,N_7992,N_7942);
nand U8334 (N_8334,N_7924,N_8084);
and U8335 (N_8335,N_8002,N_7829);
nand U8336 (N_8336,N_7825,N_8086);
nor U8337 (N_8337,N_7937,N_7854);
or U8338 (N_8338,N_7911,N_7942);
and U8339 (N_8339,N_8056,N_7913);
xnor U8340 (N_8340,N_7979,N_7959);
nand U8341 (N_8341,N_7822,N_7889);
xor U8342 (N_8342,N_8098,N_7930);
nand U8343 (N_8343,N_8029,N_7983);
nand U8344 (N_8344,N_7999,N_8051);
nand U8345 (N_8345,N_8060,N_7868);
xor U8346 (N_8346,N_7920,N_8001);
nand U8347 (N_8347,N_7967,N_7952);
nand U8348 (N_8348,N_7975,N_7846);
and U8349 (N_8349,N_8030,N_7847);
or U8350 (N_8350,N_8005,N_7853);
nand U8351 (N_8351,N_7900,N_7837);
nor U8352 (N_8352,N_8050,N_7995);
or U8353 (N_8353,N_7945,N_7888);
nand U8354 (N_8354,N_7892,N_7897);
xor U8355 (N_8355,N_7811,N_8006);
xor U8356 (N_8356,N_8072,N_8035);
nand U8357 (N_8357,N_7974,N_7853);
and U8358 (N_8358,N_7949,N_8091);
or U8359 (N_8359,N_8068,N_7801);
xor U8360 (N_8360,N_7846,N_7852);
or U8361 (N_8361,N_7992,N_8020);
xnor U8362 (N_8362,N_8021,N_7937);
nor U8363 (N_8363,N_7814,N_7996);
and U8364 (N_8364,N_7804,N_8097);
and U8365 (N_8365,N_7885,N_7939);
nand U8366 (N_8366,N_8008,N_7929);
or U8367 (N_8367,N_7809,N_7906);
nor U8368 (N_8368,N_7949,N_7952);
and U8369 (N_8369,N_7975,N_7845);
xor U8370 (N_8370,N_7859,N_7909);
or U8371 (N_8371,N_7890,N_8059);
and U8372 (N_8372,N_7818,N_7991);
xor U8373 (N_8373,N_8006,N_7929);
xor U8374 (N_8374,N_7931,N_7937);
nand U8375 (N_8375,N_7847,N_7888);
nand U8376 (N_8376,N_8018,N_7988);
xnor U8377 (N_8377,N_8094,N_7884);
nand U8378 (N_8378,N_7823,N_7876);
xnor U8379 (N_8379,N_8066,N_8037);
nand U8380 (N_8380,N_7895,N_8057);
xor U8381 (N_8381,N_7959,N_7845);
xnor U8382 (N_8382,N_7991,N_7812);
nand U8383 (N_8383,N_7943,N_8044);
xnor U8384 (N_8384,N_7895,N_7991);
or U8385 (N_8385,N_7975,N_7979);
nand U8386 (N_8386,N_7903,N_7910);
nand U8387 (N_8387,N_8033,N_8005);
xnor U8388 (N_8388,N_7974,N_7822);
nand U8389 (N_8389,N_7854,N_7837);
nor U8390 (N_8390,N_8070,N_7853);
xor U8391 (N_8391,N_7994,N_8085);
xnor U8392 (N_8392,N_8068,N_7996);
nand U8393 (N_8393,N_8090,N_7982);
and U8394 (N_8394,N_7891,N_7864);
and U8395 (N_8395,N_7912,N_7940);
or U8396 (N_8396,N_7978,N_8025);
nor U8397 (N_8397,N_7907,N_7954);
or U8398 (N_8398,N_8074,N_7889);
nand U8399 (N_8399,N_8029,N_7890);
xor U8400 (N_8400,N_8286,N_8346);
xor U8401 (N_8401,N_8239,N_8368);
xnor U8402 (N_8402,N_8102,N_8390);
nand U8403 (N_8403,N_8397,N_8183);
nand U8404 (N_8404,N_8240,N_8379);
or U8405 (N_8405,N_8225,N_8280);
or U8406 (N_8406,N_8350,N_8103);
nand U8407 (N_8407,N_8215,N_8101);
nand U8408 (N_8408,N_8333,N_8169);
nand U8409 (N_8409,N_8195,N_8224);
nor U8410 (N_8410,N_8115,N_8209);
nand U8411 (N_8411,N_8228,N_8185);
xor U8412 (N_8412,N_8159,N_8151);
nand U8413 (N_8413,N_8315,N_8398);
and U8414 (N_8414,N_8150,N_8389);
nand U8415 (N_8415,N_8275,N_8129);
and U8416 (N_8416,N_8313,N_8160);
nand U8417 (N_8417,N_8383,N_8367);
or U8418 (N_8418,N_8120,N_8170);
nor U8419 (N_8419,N_8235,N_8393);
nor U8420 (N_8420,N_8245,N_8107);
or U8421 (N_8421,N_8381,N_8281);
xor U8422 (N_8422,N_8362,N_8136);
nand U8423 (N_8423,N_8269,N_8283);
and U8424 (N_8424,N_8312,N_8143);
and U8425 (N_8425,N_8144,N_8382);
nor U8426 (N_8426,N_8268,N_8249);
and U8427 (N_8427,N_8250,N_8207);
and U8428 (N_8428,N_8260,N_8234);
nor U8429 (N_8429,N_8306,N_8282);
nand U8430 (N_8430,N_8329,N_8272);
nand U8431 (N_8431,N_8292,N_8366);
nor U8432 (N_8432,N_8158,N_8387);
nor U8433 (N_8433,N_8267,N_8347);
xor U8434 (N_8434,N_8331,N_8104);
and U8435 (N_8435,N_8203,N_8376);
or U8436 (N_8436,N_8246,N_8307);
or U8437 (N_8437,N_8348,N_8192);
or U8438 (N_8438,N_8277,N_8180);
xnor U8439 (N_8439,N_8298,N_8221);
nor U8440 (N_8440,N_8175,N_8201);
xnor U8441 (N_8441,N_8178,N_8237);
or U8442 (N_8442,N_8188,N_8165);
xnor U8443 (N_8443,N_8352,N_8243);
nand U8444 (N_8444,N_8375,N_8179);
and U8445 (N_8445,N_8216,N_8285);
xor U8446 (N_8446,N_8155,N_8141);
or U8447 (N_8447,N_8344,N_8276);
and U8448 (N_8448,N_8238,N_8130);
nand U8449 (N_8449,N_8223,N_8162);
nor U8450 (N_8450,N_8318,N_8324);
nor U8451 (N_8451,N_8258,N_8374);
nand U8452 (N_8452,N_8135,N_8380);
nor U8453 (N_8453,N_8392,N_8241);
xor U8454 (N_8454,N_8154,N_8290);
or U8455 (N_8455,N_8229,N_8113);
nand U8456 (N_8456,N_8386,N_8127);
nand U8457 (N_8457,N_8371,N_8369);
nand U8458 (N_8458,N_8217,N_8328);
xnor U8459 (N_8459,N_8182,N_8213);
and U8460 (N_8460,N_8364,N_8167);
xor U8461 (N_8461,N_8138,N_8373);
nor U8462 (N_8462,N_8247,N_8124);
nor U8463 (N_8463,N_8140,N_8126);
xnor U8464 (N_8464,N_8142,N_8322);
nand U8465 (N_8465,N_8230,N_8314);
or U8466 (N_8466,N_8190,N_8289);
or U8467 (N_8467,N_8174,N_8134);
nand U8468 (N_8468,N_8214,N_8219);
nand U8469 (N_8469,N_8359,N_8173);
xnor U8470 (N_8470,N_8163,N_8197);
nand U8471 (N_8471,N_8334,N_8222);
and U8472 (N_8472,N_8394,N_8252);
xor U8473 (N_8473,N_8122,N_8205);
xor U8474 (N_8474,N_8321,N_8261);
or U8475 (N_8475,N_8399,N_8264);
nor U8476 (N_8476,N_8156,N_8161);
xor U8477 (N_8477,N_8149,N_8337);
or U8478 (N_8478,N_8172,N_8273);
xor U8479 (N_8479,N_8262,N_8147);
nand U8480 (N_8480,N_8356,N_8365);
xor U8481 (N_8481,N_8302,N_8152);
nor U8482 (N_8482,N_8291,N_8327);
nor U8483 (N_8483,N_8300,N_8297);
xor U8484 (N_8484,N_8330,N_8168);
xnor U8485 (N_8485,N_8299,N_8351);
nand U8486 (N_8486,N_8384,N_8372);
xor U8487 (N_8487,N_8184,N_8319);
nand U8488 (N_8488,N_8339,N_8320);
xor U8489 (N_8489,N_8106,N_8231);
or U8490 (N_8490,N_8284,N_8370);
or U8491 (N_8491,N_8293,N_8354);
nor U8492 (N_8492,N_8308,N_8257);
nand U8493 (N_8493,N_8187,N_8202);
and U8494 (N_8494,N_8131,N_8388);
and U8495 (N_8495,N_8316,N_8193);
nand U8496 (N_8496,N_8226,N_8125);
nand U8497 (N_8497,N_8349,N_8164);
xor U8498 (N_8498,N_8326,N_8189);
or U8499 (N_8499,N_8204,N_8177);
nor U8500 (N_8500,N_8119,N_8391);
or U8501 (N_8501,N_8117,N_8153);
xnor U8502 (N_8502,N_8353,N_8111);
or U8503 (N_8503,N_8311,N_8199);
and U8504 (N_8504,N_8363,N_8305);
and U8505 (N_8505,N_8256,N_8211);
nor U8506 (N_8506,N_8358,N_8146);
xor U8507 (N_8507,N_8342,N_8212);
nor U8508 (N_8508,N_8139,N_8196);
and U8509 (N_8509,N_8378,N_8294);
nor U8510 (N_8510,N_8251,N_8287);
nor U8511 (N_8511,N_8310,N_8116);
nor U8512 (N_8512,N_8198,N_8145);
xor U8513 (N_8513,N_8360,N_8309);
xor U8514 (N_8514,N_8206,N_8227);
nand U8515 (N_8515,N_8244,N_8114);
nor U8516 (N_8516,N_8176,N_8171);
nand U8517 (N_8517,N_8236,N_8385);
nor U8518 (N_8518,N_8323,N_8301);
nor U8519 (N_8519,N_8361,N_8259);
and U8520 (N_8520,N_8181,N_8110);
nor U8521 (N_8521,N_8242,N_8295);
nand U8522 (N_8522,N_8137,N_8266);
or U8523 (N_8523,N_8233,N_8132);
and U8524 (N_8524,N_8274,N_8166);
nor U8525 (N_8525,N_8303,N_8105);
nor U8526 (N_8526,N_8271,N_8288);
xor U8527 (N_8527,N_8296,N_8255);
nor U8528 (N_8528,N_8232,N_8335);
or U8529 (N_8529,N_8148,N_8338);
and U8530 (N_8530,N_8263,N_8109);
or U8531 (N_8531,N_8340,N_8194);
xor U8532 (N_8532,N_8157,N_8200);
nor U8533 (N_8533,N_8121,N_8278);
xor U8534 (N_8534,N_8112,N_8128);
or U8535 (N_8535,N_8218,N_8220);
or U8536 (N_8536,N_8317,N_8304);
nor U8537 (N_8537,N_8100,N_8123);
nand U8538 (N_8538,N_8265,N_8253);
nand U8539 (N_8539,N_8254,N_8325);
and U8540 (N_8540,N_8341,N_8377);
and U8541 (N_8541,N_8355,N_8270);
or U8542 (N_8542,N_8118,N_8248);
nor U8543 (N_8543,N_8332,N_8108);
xor U8544 (N_8544,N_8133,N_8186);
and U8545 (N_8545,N_8396,N_8336);
xnor U8546 (N_8546,N_8357,N_8191);
nand U8547 (N_8547,N_8210,N_8343);
or U8548 (N_8548,N_8395,N_8208);
and U8549 (N_8549,N_8345,N_8279);
nor U8550 (N_8550,N_8132,N_8161);
nor U8551 (N_8551,N_8213,N_8341);
and U8552 (N_8552,N_8246,N_8292);
or U8553 (N_8553,N_8141,N_8329);
xor U8554 (N_8554,N_8322,N_8325);
nand U8555 (N_8555,N_8321,N_8243);
nor U8556 (N_8556,N_8259,N_8368);
nand U8557 (N_8557,N_8135,N_8132);
nor U8558 (N_8558,N_8190,N_8158);
or U8559 (N_8559,N_8185,N_8125);
nor U8560 (N_8560,N_8374,N_8395);
xnor U8561 (N_8561,N_8324,N_8326);
and U8562 (N_8562,N_8339,N_8198);
or U8563 (N_8563,N_8353,N_8143);
nor U8564 (N_8564,N_8260,N_8276);
xnor U8565 (N_8565,N_8270,N_8227);
or U8566 (N_8566,N_8310,N_8395);
or U8567 (N_8567,N_8305,N_8252);
xnor U8568 (N_8568,N_8317,N_8216);
or U8569 (N_8569,N_8146,N_8279);
and U8570 (N_8570,N_8147,N_8142);
nand U8571 (N_8571,N_8142,N_8100);
nor U8572 (N_8572,N_8143,N_8205);
xor U8573 (N_8573,N_8219,N_8231);
xnor U8574 (N_8574,N_8136,N_8397);
or U8575 (N_8575,N_8331,N_8360);
and U8576 (N_8576,N_8294,N_8239);
nand U8577 (N_8577,N_8114,N_8130);
nand U8578 (N_8578,N_8392,N_8317);
nand U8579 (N_8579,N_8248,N_8279);
nand U8580 (N_8580,N_8374,N_8238);
nor U8581 (N_8581,N_8181,N_8330);
nand U8582 (N_8582,N_8140,N_8330);
nor U8583 (N_8583,N_8331,N_8338);
nor U8584 (N_8584,N_8301,N_8132);
xor U8585 (N_8585,N_8150,N_8139);
xnor U8586 (N_8586,N_8376,N_8250);
nor U8587 (N_8587,N_8278,N_8107);
or U8588 (N_8588,N_8129,N_8321);
nor U8589 (N_8589,N_8184,N_8131);
nor U8590 (N_8590,N_8334,N_8279);
and U8591 (N_8591,N_8150,N_8205);
or U8592 (N_8592,N_8392,N_8211);
xnor U8593 (N_8593,N_8306,N_8397);
and U8594 (N_8594,N_8128,N_8195);
and U8595 (N_8595,N_8389,N_8393);
nor U8596 (N_8596,N_8272,N_8104);
xnor U8597 (N_8597,N_8175,N_8189);
nor U8598 (N_8598,N_8277,N_8338);
xor U8599 (N_8599,N_8374,N_8334);
or U8600 (N_8600,N_8216,N_8153);
xnor U8601 (N_8601,N_8296,N_8314);
nor U8602 (N_8602,N_8236,N_8117);
nand U8603 (N_8603,N_8256,N_8360);
nor U8604 (N_8604,N_8100,N_8232);
nand U8605 (N_8605,N_8340,N_8319);
xor U8606 (N_8606,N_8147,N_8320);
nand U8607 (N_8607,N_8118,N_8323);
or U8608 (N_8608,N_8302,N_8142);
nor U8609 (N_8609,N_8240,N_8220);
and U8610 (N_8610,N_8200,N_8211);
or U8611 (N_8611,N_8274,N_8295);
and U8612 (N_8612,N_8245,N_8367);
and U8613 (N_8613,N_8108,N_8207);
nand U8614 (N_8614,N_8377,N_8314);
nand U8615 (N_8615,N_8104,N_8108);
nor U8616 (N_8616,N_8345,N_8207);
and U8617 (N_8617,N_8273,N_8146);
nor U8618 (N_8618,N_8184,N_8378);
nand U8619 (N_8619,N_8269,N_8342);
xnor U8620 (N_8620,N_8360,N_8189);
and U8621 (N_8621,N_8252,N_8237);
xor U8622 (N_8622,N_8379,N_8349);
nor U8623 (N_8623,N_8336,N_8303);
nand U8624 (N_8624,N_8142,N_8160);
nand U8625 (N_8625,N_8312,N_8166);
and U8626 (N_8626,N_8213,N_8131);
and U8627 (N_8627,N_8124,N_8257);
nor U8628 (N_8628,N_8219,N_8225);
nor U8629 (N_8629,N_8168,N_8159);
or U8630 (N_8630,N_8113,N_8239);
or U8631 (N_8631,N_8188,N_8142);
nor U8632 (N_8632,N_8274,N_8329);
nand U8633 (N_8633,N_8214,N_8340);
xnor U8634 (N_8634,N_8288,N_8254);
nand U8635 (N_8635,N_8124,N_8113);
nand U8636 (N_8636,N_8139,N_8282);
xor U8637 (N_8637,N_8326,N_8242);
xnor U8638 (N_8638,N_8343,N_8368);
and U8639 (N_8639,N_8298,N_8213);
nand U8640 (N_8640,N_8341,N_8203);
nand U8641 (N_8641,N_8366,N_8399);
nand U8642 (N_8642,N_8286,N_8347);
xor U8643 (N_8643,N_8277,N_8385);
or U8644 (N_8644,N_8190,N_8392);
or U8645 (N_8645,N_8261,N_8371);
nand U8646 (N_8646,N_8220,N_8239);
nor U8647 (N_8647,N_8105,N_8204);
or U8648 (N_8648,N_8135,N_8264);
or U8649 (N_8649,N_8101,N_8103);
and U8650 (N_8650,N_8291,N_8279);
nor U8651 (N_8651,N_8207,N_8142);
and U8652 (N_8652,N_8139,N_8285);
xnor U8653 (N_8653,N_8287,N_8310);
nor U8654 (N_8654,N_8282,N_8252);
nor U8655 (N_8655,N_8344,N_8256);
nor U8656 (N_8656,N_8144,N_8125);
nand U8657 (N_8657,N_8196,N_8385);
xor U8658 (N_8658,N_8381,N_8244);
and U8659 (N_8659,N_8124,N_8366);
nand U8660 (N_8660,N_8249,N_8156);
nor U8661 (N_8661,N_8251,N_8277);
xor U8662 (N_8662,N_8154,N_8258);
and U8663 (N_8663,N_8353,N_8320);
or U8664 (N_8664,N_8222,N_8385);
xor U8665 (N_8665,N_8257,N_8106);
nand U8666 (N_8666,N_8122,N_8319);
or U8667 (N_8667,N_8287,N_8323);
xnor U8668 (N_8668,N_8110,N_8240);
xor U8669 (N_8669,N_8271,N_8228);
nand U8670 (N_8670,N_8222,N_8354);
and U8671 (N_8671,N_8395,N_8134);
and U8672 (N_8672,N_8119,N_8220);
nand U8673 (N_8673,N_8302,N_8248);
xnor U8674 (N_8674,N_8256,N_8266);
xnor U8675 (N_8675,N_8101,N_8356);
and U8676 (N_8676,N_8167,N_8365);
xor U8677 (N_8677,N_8276,N_8180);
nand U8678 (N_8678,N_8286,N_8205);
nor U8679 (N_8679,N_8245,N_8282);
nand U8680 (N_8680,N_8268,N_8341);
nor U8681 (N_8681,N_8164,N_8141);
nand U8682 (N_8682,N_8347,N_8240);
and U8683 (N_8683,N_8210,N_8345);
or U8684 (N_8684,N_8347,N_8256);
xor U8685 (N_8685,N_8170,N_8335);
nand U8686 (N_8686,N_8239,N_8329);
nand U8687 (N_8687,N_8276,N_8104);
nand U8688 (N_8688,N_8286,N_8297);
nand U8689 (N_8689,N_8225,N_8109);
nor U8690 (N_8690,N_8317,N_8203);
nand U8691 (N_8691,N_8306,N_8371);
and U8692 (N_8692,N_8296,N_8394);
or U8693 (N_8693,N_8125,N_8259);
and U8694 (N_8694,N_8224,N_8187);
and U8695 (N_8695,N_8118,N_8396);
or U8696 (N_8696,N_8390,N_8203);
xnor U8697 (N_8697,N_8103,N_8235);
and U8698 (N_8698,N_8149,N_8235);
xor U8699 (N_8699,N_8394,N_8223);
or U8700 (N_8700,N_8698,N_8587);
xor U8701 (N_8701,N_8582,N_8466);
xnor U8702 (N_8702,N_8670,N_8584);
and U8703 (N_8703,N_8435,N_8617);
or U8704 (N_8704,N_8609,N_8694);
xnor U8705 (N_8705,N_8431,N_8636);
xor U8706 (N_8706,N_8571,N_8403);
nor U8707 (N_8707,N_8622,N_8551);
and U8708 (N_8708,N_8643,N_8432);
nor U8709 (N_8709,N_8409,N_8592);
xor U8710 (N_8710,N_8553,N_8594);
nand U8711 (N_8711,N_8413,N_8494);
and U8712 (N_8712,N_8442,N_8591);
and U8713 (N_8713,N_8642,N_8569);
xnor U8714 (N_8714,N_8401,N_8681);
xnor U8715 (N_8715,N_8597,N_8545);
or U8716 (N_8716,N_8464,N_8461);
and U8717 (N_8717,N_8679,N_8665);
xor U8718 (N_8718,N_8512,N_8497);
or U8719 (N_8719,N_8596,N_8533);
xnor U8720 (N_8720,N_8502,N_8635);
and U8721 (N_8721,N_8486,N_8619);
xor U8722 (N_8722,N_8680,N_8568);
or U8723 (N_8723,N_8580,N_8540);
or U8724 (N_8724,N_8601,N_8405);
or U8725 (N_8725,N_8437,N_8542);
xnor U8726 (N_8726,N_8653,N_8657);
nor U8727 (N_8727,N_8566,N_8589);
or U8728 (N_8728,N_8570,N_8599);
xnor U8729 (N_8729,N_8523,N_8633);
xor U8730 (N_8730,N_8581,N_8530);
nand U8731 (N_8731,N_8450,N_8526);
or U8732 (N_8732,N_8691,N_8645);
nor U8733 (N_8733,N_8620,N_8534);
xnor U8734 (N_8734,N_8663,N_8419);
or U8735 (N_8735,N_8406,N_8471);
or U8736 (N_8736,N_8425,N_8404);
nand U8737 (N_8737,N_8561,N_8506);
nor U8738 (N_8738,N_8448,N_8460);
or U8739 (N_8739,N_8400,N_8456);
xor U8740 (N_8740,N_8529,N_8675);
or U8741 (N_8741,N_8402,N_8490);
nor U8742 (N_8742,N_8430,N_8600);
nor U8743 (N_8743,N_8583,N_8588);
and U8744 (N_8744,N_8557,N_8647);
and U8745 (N_8745,N_8614,N_8493);
nand U8746 (N_8746,N_8624,N_8519);
xor U8747 (N_8747,N_8436,N_8669);
and U8748 (N_8748,N_8682,N_8412);
xnor U8749 (N_8749,N_8503,N_8631);
xnor U8750 (N_8750,N_8517,N_8524);
nor U8751 (N_8751,N_8516,N_8666);
xor U8752 (N_8752,N_8485,N_8625);
xnor U8753 (N_8753,N_8439,N_8472);
xor U8754 (N_8754,N_8480,N_8550);
or U8755 (N_8755,N_8573,N_8626);
or U8756 (N_8756,N_8611,N_8606);
or U8757 (N_8757,N_8556,N_8613);
nand U8758 (N_8758,N_8664,N_8408);
and U8759 (N_8759,N_8515,N_8661);
nand U8760 (N_8760,N_8513,N_8484);
nor U8761 (N_8761,N_8504,N_8543);
and U8762 (N_8762,N_8446,N_8465);
xnor U8763 (N_8763,N_8659,N_8415);
xnor U8764 (N_8764,N_8638,N_8567);
or U8765 (N_8765,N_8541,N_8438);
nor U8766 (N_8766,N_8654,N_8443);
xor U8767 (N_8767,N_8574,N_8693);
or U8768 (N_8768,N_8518,N_8469);
nand U8769 (N_8769,N_8632,N_8414);
nand U8770 (N_8770,N_8467,N_8454);
nand U8771 (N_8771,N_8558,N_8668);
nor U8772 (N_8772,N_8605,N_8699);
nand U8773 (N_8773,N_8423,N_8552);
nor U8774 (N_8774,N_8627,N_8487);
or U8775 (N_8775,N_8420,N_8473);
and U8776 (N_8776,N_8585,N_8528);
nor U8777 (N_8777,N_8685,N_8562);
nand U8778 (N_8778,N_8629,N_8683);
xnor U8779 (N_8779,N_8482,N_8410);
or U8780 (N_8780,N_8433,N_8416);
or U8781 (N_8781,N_8579,N_8697);
nand U8782 (N_8782,N_8559,N_8563);
and U8783 (N_8783,N_8521,N_8538);
nor U8784 (N_8784,N_8445,N_8544);
xnor U8785 (N_8785,N_8610,N_8689);
xnor U8786 (N_8786,N_8692,N_8508);
or U8787 (N_8787,N_8648,N_8674);
or U8788 (N_8788,N_8531,N_8656);
nand U8789 (N_8789,N_8628,N_8429);
or U8790 (N_8790,N_8673,N_8586);
nand U8791 (N_8791,N_8441,N_8608);
and U8792 (N_8792,N_8476,N_8478);
and U8793 (N_8793,N_8652,N_8474);
xor U8794 (N_8794,N_8695,N_8499);
xnor U8795 (N_8795,N_8554,N_8462);
or U8796 (N_8796,N_8444,N_8676);
nand U8797 (N_8797,N_8547,N_8488);
nor U8798 (N_8798,N_8495,N_8549);
xor U8799 (N_8799,N_8483,N_8560);
or U8800 (N_8800,N_8593,N_8578);
xor U8801 (N_8801,N_8576,N_8535);
nor U8802 (N_8802,N_8424,N_8667);
nand U8803 (N_8803,N_8640,N_8427);
xor U8804 (N_8804,N_8658,N_8696);
or U8805 (N_8805,N_8615,N_8477);
and U8806 (N_8806,N_8595,N_8520);
or U8807 (N_8807,N_8489,N_8447);
nand U8808 (N_8808,N_8537,N_8407);
and U8809 (N_8809,N_8525,N_8422);
xor U8810 (N_8810,N_8514,N_8565);
and U8811 (N_8811,N_8655,N_8603);
and U8812 (N_8812,N_8660,N_8649);
nor U8813 (N_8813,N_8548,N_8644);
nand U8814 (N_8814,N_8688,N_8527);
and U8815 (N_8815,N_8498,N_8479);
nor U8816 (N_8816,N_8492,N_8532);
nor U8817 (N_8817,N_8481,N_8510);
or U8818 (N_8818,N_8612,N_8598);
nand U8819 (N_8819,N_8616,N_8505);
xnor U8820 (N_8820,N_8539,N_8451);
nand U8821 (N_8821,N_8496,N_8421);
nor U8822 (N_8822,N_8623,N_8639);
xor U8823 (N_8823,N_8672,N_8677);
xor U8824 (N_8824,N_8511,N_8470);
or U8825 (N_8825,N_8468,N_8646);
and U8826 (N_8826,N_8453,N_8452);
xor U8827 (N_8827,N_8684,N_8536);
xnor U8828 (N_8828,N_8455,N_8417);
or U8829 (N_8829,N_8418,N_8671);
and U8830 (N_8830,N_8428,N_8440);
xor U8831 (N_8831,N_8463,N_8564);
and U8832 (N_8832,N_8411,N_8491);
and U8833 (N_8833,N_8662,N_8577);
nor U8834 (N_8834,N_8590,N_8507);
xnor U8835 (N_8835,N_8522,N_8449);
nand U8836 (N_8836,N_8457,N_8637);
nor U8837 (N_8837,N_8607,N_8687);
xor U8838 (N_8838,N_8475,N_8500);
and U8839 (N_8839,N_8634,N_8690);
or U8840 (N_8840,N_8602,N_8621);
and U8841 (N_8841,N_8546,N_8575);
and U8842 (N_8842,N_8501,N_8458);
nand U8843 (N_8843,N_8604,N_8686);
xor U8844 (N_8844,N_8678,N_8509);
nand U8845 (N_8845,N_8555,N_8459);
and U8846 (N_8846,N_8618,N_8630);
nor U8847 (N_8847,N_8426,N_8434);
or U8848 (N_8848,N_8650,N_8651);
nand U8849 (N_8849,N_8641,N_8572);
nor U8850 (N_8850,N_8672,N_8459);
or U8851 (N_8851,N_8449,N_8410);
xnor U8852 (N_8852,N_8639,N_8503);
nor U8853 (N_8853,N_8687,N_8677);
nand U8854 (N_8854,N_8462,N_8542);
nand U8855 (N_8855,N_8535,N_8575);
xor U8856 (N_8856,N_8647,N_8411);
nor U8857 (N_8857,N_8506,N_8493);
and U8858 (N_8858,N_8420,N_8651);
or U8859 (N_8859,N_8675,N_8679);
nand U8860 (N_8860,N_8434,N_8458);
nor U8861 (N_8861,N_8541,N_8448);
nor U8862 (N_8862,N_8544,N_8639);
or U8863 (N_8863,N_8574,N_8486);
xnor U8864 (N_8864,N_8502,N_8536);
or U8865 (N_8865,N_8482,N_8670);
or U8866 (N_8866,N_8547,N_8575);
nor U8867 (N_8867,N_8660,N_8585);
nor U8868 (N_8868,N_8575,N_8657);
or U8869 (N_8869,N_8538,N_8486);
or U8870 (N_8870,N_8548,N_8650);
and U8871 (N_8871,N_8600,N_8632);
xor U8872 (N_8872,N_8485,N_8670);
and U8873 (N_8873,N_8585,N_8517);
nor U8874 (N_8874,N_8600,N_8417);
xnor U8875 (N_8875,N_8583,N_8692);
and U8876 (N_8876,N_8450,N_8676);
and U8877 (N_8877,N_8589,N_8536);
or U8878 (N_8878,N_8413,N_8572);
nand U8879 (N_8879,N_8496,N_8671);
xor U8880 (N_8880,N_8420,N_8639);
nor U8881 (N_8881,N_8623,N_8650);
and U8882 (N_8882,N_8681,N_8547);
or U8883 (N_8883,N_8657,N_8688);
or U8884 (N_8884,N_8664,N_8435);
xor U8885 (N_8885,N_8434,N_8460);
xor U8886 (N_8886,N_8586,N_8562);
nor U8887 (N_8887,N_8572,N_8685);
xor U8888 (N_8888,N_8674,N_8676);
and U8889 (N_8889,N_8665,N_8514);
and U8890 (N_8890,N_8556,N_8422);
xor U8891 (N_8891,N_8577,N_8561);
and U8892 (N_8892,N_8581,N_8578);
or U8893 (N_8893,N_8436,N_8481);
nor U8894 (N_8894,N_8625,N_8593);
and U8895 (N_8895,N_8601,N_8567);
and U8896 (N_8896,N_8549,N_8527);
or U8897 (N_8897,N_8458,N_8599);
nor U8898 (N_8898,N_8521,N_8658);
nand U8899 (N_8899,N_8518,N_8622);
xnor U8900 (N_8900,N_8537,N_8699);
nand U8901 (N_8901,N_8490,N_8612);
xor U8902 (N_8902,N_8693,N_8508);
xnor U8903 (N_8903,N_8689,N_8428);
and U8904 (N_8904,N_8415,N_8566);
or U8905 (N_8905,N_8584,N_8431);
nand U8906 (N_8906,N_8424,N_8656);
or U8907 (N_8907,N_8622,N_8661);
nand U8908 (N_8908,N_8400,N_8484);
and U8909 (N_8909,N_8658,N_8672);
xor U8910 (N_8910,N_8405,N_8445);
or U8911 (N_8911,N_8607,N_8544);
or U8912 (N_8912,N_8415,N_8649);
nand U8913 (N_8913,N_8497,N_8586);
nand U8914 (N_8914,N_8685,N_8662);
and U8915 (N_8915,N_8629,N_8561);
nor U8916 (N_8916,N_8407,N_8636);
and U8917 (N_8917,N_8426,N_8653);
nor U8918 (N_8918,N_8539,N_8512);
nor U8919 (N_8919,N_8461,N_8652);
nor U8920 (N_8920,N_8407,N_8410);
nor U8921 (N_8921,N_8625,N_8536);
nand U8922 (N_8922,N_8419,N_8405);
nand U8923 (N_8923,N_8676,N_8572);
or U8924 (N_8924,N_8582,N_8621);
xnor U8925 (N_8925,N_8613,N_8590);
nor U8926 (N_8926,N_8428,N_8452);
nor U8927 (N_8927,N_8609,N_8683);
nand U8928 (N_8928,N_8523,N_8681);
nand U8929 (N_8929,N_8505,N_8450);
nand U8930 (N_8930,N_8649,N_8400);
and U8931 (N_8931,N_8545,N_8424);
xnor U8932 (N_8932,N_8546,N_8537);
and U8933 (N_8933,N_8532,N_8693);
nand U8934 (N_8934,N_8455,N_8570);
nor U8935 (N_8935,N_8432,N_8695);
or U8936 (N_8936,N_8647,N_8579);
nand U8937 (N_8937,N_8629,N_8648);
nand U8938 (N_8938,N_8670,N_8629);
nor U8939 (N_8939,N_8518,N_8530);
and U8940 (N_8940,N_8528,N_8423);
or U8941 (N_8941,N_8635,N_8689);
xnor U8942 (N_8942,N_8602,N_8430);
or U8943 (N_8943,N_8411,N_8695);
or U8944 (N_8944,N_8528,N_8653);
nor U8945 (N_8945,N_8628,N_8418);
nor U8946 (N_8946,N_8523,N_8619);
xor U8947 (N_8947,N_8502,N_8668);
or U8948 (N_8948,N_8443,N_8431);
and U8949 (N_8949,N_8423,N_8629);
xnor U8950 (N_8950,N_8542,N_8521);
nand U8951 (N_8951,N_8646,N_8580);
nor U8952 (N_8952,N_8641,N_8445);
xnor U8953 (N_8953,N_8621,N_8508);
xor U8954 (N_8954,N_8583,N_8425);
nand U8955 (N_8955,N_8619,N_8477);
xnor U8956 (N_8956,N_8509,N_8699);
or U8957 (N_8957,N_8528,N_8480);
and U8958 (N_8958,N_8470,N_8668);
nand U8959 (N_8959,N_8541,N_8593);
and U8960 (N_8960,N_8655,N_8431);
nand U8961 (N_8961,N_8661,N_8555);
xor U8962 (N_8962,N_8667,N_8543);
and U8963 (N_8963,N_8445,N_8566);
nand U8964 (N_8964,N_8562,N_8502);
xnor U8965 (N_8965,N_8572,N_8404);
xnor U8966 (N_8966,N_8595,N_8508);
nand U8967 (N_8967,N_8611,N_8547);
and U8968 (N_8968,N_8651,N_8640);
and U8969 (N_8969,N_8512,N_8679);
or U8970 (N_8970,N_8435,N_8422);
nand U8971 (N_8971,N_8501,N_8670);
xor U8972 (N_8972,N_8538,N_8670);
and U8973 (N_8973,N_8406,N_8470);
nor U8974 (N_8974,N_8624,N_8541);
xnor U8975 (N_8975,N_8687,N_8494);
nor U8976 (N_8976,N_8516,N_8621);
nor U8977 (N_8977,N_8509,N_8416);
and U8978 (N_8978,N_8462,N_8533);
nor U8979 (N_8979,N_8475,N_8617);
nor U8980 (N_8980,N_8417,N_8658);
and U8981 (N_8981,N_8618,N_8535);
nand U8982 (N_8982,N_8475,N_8597);
nor U8983 (N_8983,N_8604,N_8465);
and U8984 (N_8984,N_8690,N_8498);
xor U8985 (N_8985,N_8612,N_8463);
nand U8986 (N_8986,N_8581,N_8402);
or U8987 (N_8987,N_8558,N_8594);
nor U8988 (N_8988,N_8528,N_8556);
or U8989 (N_8989,N_8643,N_8493);
xor U8990 (N_8990,N_8615,N_8487);
xor U8991 (N_8991,N_8604,N_8555);
nor U8992 (N_8992,N_8589,N_8672);
or U8993 (N_8993,N_8683,N_8506);
xor U8994 (N_8994,N_8479,N_8544);
nor U8995 (N_8995,N_8477,N_8691);
or U8996 (N_8996,N_8634,N_8513);
nand U8997 (N_8997,N_8490,N_8558);
xor U8998 (N_8998,N_8542,N_8492);
nand U8999 (N_8999,N_8545,N_8684);
nand U9000 (N_9000,N_8976,N_8826);
xnor U9001 (N_9001,N_8978,N_8831);
or U9002 (N_9002,N_8992,N_8825);
xor U9003 (N_9003,N_8941,N_8870);
or U9004 (N_9004,N_8944,N_8799);
xor U9005 (N_9005,N_8769,N_8847);
nand U9006 (N_9006,N_8701,N_8962);
and U9007 (N_9007,N_8951,N_8706);
or U9008 (N_9008,N_8998,N_8728);
and U9009 (N_9009,N_8982,N_8904);
or U9010 (N_9010,N_8788,N_8913);
nand U9011 (N_9011,N_8990,N_8731);
xor U9012 (N_9012,N_8873,N_8861);
or U9013 (N_9013,N_8919,N_8794);
or U9014 (N_9014,N_8848,N_8757);
nor U9015 (N_9015,N_8778,N_8797);
and U9016 (N_9016,N_8755,N_8866);
and U9017 (N_9017,N_8879,N_8885);
and U9018 (N_9018,N_8751,N_8928);
nand U9019 (N_9019,N_8878,N_8897);
xor U9020 (N_9020,N_8853,N_8971);
nand U9021 (N_9021,N_8760,N_8958);
or U9022 (N_9022,N_8785,N_8790);
or U9023 (N_9023,N_8752,N_8834);
nand U9024 (N_9024,N_8929,N_8812);
or U9025 (N_9025,N_8918,N_8827);
and U9026 (N_9026,N_8773,N_8874);
or U9027 (N_9027,N_8739,N_8732);
nor U9028 (N_9028,N_8758,N_8965);
xor U9029 (N_9029,N_8750,N_8767);
nor U9030 (N_9030,N_8914,N_8796);
or U9031 (N_9031,N_8930,N_8849);
xnor U9032 (N_9032,N_8940,N_8815);
and U9033 (N_9033,N_8884,N_8725);
nor U9034 (N_9034,N_8991,N_8880);
nor U9035 (N_9035,N_8737,N_8886);
or U9036 (N_9036,N_8933,N_8912);
nand U9037 (N_9037,N_8721,N_8926);
or U9038 (N_9038,N_8865,N_8939);
xnor U9039 (N_9039,N_8882,N_8810);
and U9040 (N_9040,N_8840,N_8860);
nor U9041 (N_9041,N_8856,N_8993);
xnor U9042 (N_9042,N_8868,N_8804);
and U9043 (N_9043,N_8822,N_8942);
and U9044 (N_9044,N_8768,N_8871);
xnor U9045 (N_9045,N_8771,N_8744);
or U9046 (N_9046,N_8859,N_8902);
nand U9047 (N_9047,N_8846,N_8700);
xnor U9048 (N_9048,N_8872,N_8945);
xnor U9049 (N_9049,N_8759,N_8782);
nor U9050 (N_9050,N_8809,N_8988);
or U9051 (N_9051,N_8890,N_8843);
nor U9052 (N_9052,N_8828,N_8775);
nand U9053 (N_9053,N_8844,N_8922);
xnor U9054 (N_9054,N_8858,N_8772);
nand U9055 (N_9055,N_8749,N_8915);
or U9056 (N_9056,N_8854,N_8889);
nand U9057 (N_9057,N_8800,N_8895);
and U9058 (N_9058,N_8711,N_8949);
nor U9059 (N_9059,N_8805,N_8841);
and U9060 (N_9060,N_8961,N_8702);
nand U9061 (N_9061,N_8981,N_8832);
and U9062 (N_9062,N_8999,N_8932);
and U9063 (N_9063,N_8989,N_8776);
xor U9064 (N_9064,N_8983,N_8712);
and U9065 (N_9065,N_8845,N_8898);
nand U9066 (N_9066,N_8713,N_8803);
nor U9067 (N_9067,N_8789,N_8837);
nor U9068 (N_9068,N_8955,N_8753);
xnor U9069 (N_9069,N_8984,N_8892);
nor U9070 (N_9070,N_8927,N_8781);
nor U9071 (N_9071,N_8817,N_8907);
nor U9072 (N_9072,N_8975,N_8742);
or U9073 (N_9073,N_8777,N_8814);
xnor U9074 (N_9074,N_8977,N_8908);
xnor U9075 (N_9075,N_8823,N_8877);
nor U9076 (N_9076,N_8808,N_8906);
and U9077 (N_9077,N_8801,N_8936);
and U9078 (N_9078,N_8792,N_8935);
and U9079 (N_9079,N_8964,N_8952);
xnor U9080 (N_9080,N_8748,N_8899);
or U9081 (N_9081,N_8957,N_8900);
or U9082 (N_9082,N_8787,N_8722);
nand U9083 (N_9083,N_8791,N_8770);
xor U9084 (N_9084,N_8724,N_8887);
or U9085 (N_9085,N_8920,N_8723);
and U9086 (N_9086,N_8802,N_8973);
and U9087 (N_9087,N_8714,N_8811);
and U9088 (N_9088,N_8716,N_8979);
xnor U9089 (N_9089,N_8762,N_8705);
and U9090 (N_9090,N_8719,N_8851);
and U9091 (N_9091,N_8855,N_8783);
nor U9092 (N_9092,N_8876,N_8972);
or U9093 (N_9093,N_8974,N_8996);
nand U9094 (N_9094,N_8745,N_8730);
and U9095 (N_9095,N_8960,N_8896);
nor U9096 (N_9096,N_8763,N_8818);
xnor U9097 (N_9097,N_8881,N_8747);
and U9098 (N_9098,N_8894,N_8765);
xnor U9099 (N_9099,N_8925,N_8954);
and U9100 (N_9100,N_8830,N_8901);
xnor U9101 (N_9101,N_8917,N_8970);
and U9102 (N_9102,N_8921,N_8909);
xor U9103 (N_9103,N_8756,N_8829);
nand U9104 (N_9104,N_8888,N_8764);
or U9105 (N_9105,N_8986,N_8980);
and U9106 (N_9106,N_8835,N_8806);
nand U9107 (N_9107,N_8891,N_8820);
nor U9108 (N_9108,N_8703,N_8867);
or U9109 (N_9109,N_8943,N_8816);
and U9110 (N_9110,N_8948,N_8916);
xnor U9111 (N_9111,N_8985,N_8953);
nand U9112 (N_9112,N_8937,N_8761);
nor U9113 (N_9113,N_8807,N_8946);
nor U9114 (N_9114,N_8735,N_8824);
xnor U9115 (N_9115,N_8708,N_8821);
and U9116 (N_9116,N_8741,N_8774);
xor U9117 (N_9117,N_8710,N_8995);
xnor U9118 (N_9118,N_8836,N_8717);
and U9119 (N_9119,N_8963,N_8766);
nand U9120 (N_9120,N_8947,N_8910);
and U9121 (N_9121,N_8709,N_8715);
and U9122 (N_9122,N_8734,N_8743);
nor U9123 (N_9123,N_8833,N_8875);
xor U9124 (N_9124,N_8869,N_8862);
nor U9125 (N_9125,N_8720,N_8819);
nor U9126 (N_9126,N_8726,N_8852);
or U9127 (N_9127,N_8924,N_8704);
and U9128 (N_9128,N_8883,N_8969);
or U9129 (N_9129,N_8779,N_8718);
xor U9130 (N_9130,N_8754,N_8793);
and U9131 (N_9131,N_8903,N_8997);
nand U9132 (N_9132,N_8950,N_8729);
and U9133 (N_9133,N_8780,N_8707);
nor U9134 (N_9134,N_8798,N_8967);
xor U9135 (N_9135,N_8850,N_8738);
xnor U9136 (N_9136,N_8733,N_8842);
xor U9137 (N_9137,N_8893,N_8736);
or U9138 (N_9138,N_8923,N_8864);
and U9139 (N_9139,N_8911,N_8740);
or U9140 (N_9140,N_8968,N_8795);
nand U9141 (N_9141,N_8857,N_8863);
and U9142 (N_9142,N_8931,N_8938);
nand U9143 (N_9143,N_8934,N_8839);
nand U9144 (N_9144,N_8966,N_8813);
and U9145 (N_9145,N_8784,N_8786);
and U9146 (N_9146,N_8959,N_8838);
nand U9147 (N_9147,N_8746,N_8905);
and U9148 (N_9148,N_8727,N_8987);
nor U9149 (N_9149,N_8956,N_8994);
nor U9150 (N_9150,N_8706,N_8782);
xnor U9151 (N_9151,N_8985,N_8911);
and U9152 (N_9152,N_8714,N_8874);
nor U9153 (N_9153,N_8974,N_8965);
xor U9154 (N_9154,N_8971,N_8856);
or U9155 (N_9155,N_8978,N_8913);
xnor U9156 (N_9156,N_8888,N_8912);
and U9157 (N_9157,N_8909,N_8719);
or U9158 (N_9158,N_8718,N_8969);
or U9159 (N_9159,N_8702,N_8794);
or U9160 (N_9160,N_8798,N_8879);
nand U9161 (N_9161,N_8900,N_8941);
nor U9162 (N_9162,N_8854,N_8855);
xnor U9163 (N_9163,N_8914,N_8961);
xnor U9164 (N_9164,N_8953,N_8819);
and U9165 (N_9165,N_8709,N_8953);
nand U9166 (N_9166,N_8895,N_8837);
nor U9167 (N_9167,N_8770,N_8972);
nor U9168 (N_9168,N_8910,N_8950);
or U9169 (N_9169,N_8830,N_8903);
nor U9170 (N_9170,N_8958,N_8896);
and U9171 (N_9171,N_8876,N_8862);
xor U9172 (N_9172,N_8737,N_8797);
or U9173 (N_9173,N_8878,N_8984);
nand U9174 (N_9174,N_8756,N_8743);
nand U9175 (N_9175,N_8935,N_8896);
and U9176 (N_9176,N_8932,N_8916);
nand U9177 (N_9177,N_8997,N_8782);
nor U9178 (N_9178,N_8814,N_8711);
and U9179 (N_9179,N_8746,N_8774);
nand U9180 (N_9180,N_8894,N_8790);
nor U9181 (N_9181,N_8843,N_8834);
and U9182 (N_9182,N_8820,N_8850);
and U9183 (N_9183,N_8958,N_8869);
and U9184 (N_9184,N_8767,N_8871);
and U9185 (N_9185,N_8771,N_8710);
and U9186 (N_9186,N_8972,N_8983);
or U9187 (N_9187,N_8948,N_8991);
xor U9188 (N_9188,N_8756,N_8769);
xor U9189 (N_9189,N_8929,N_8933);
nor U9190 (N_9190,N_8793,N_8836);
or U9191 (N_9191,N_8976,N_8943);
nand U9192 (N_9192,N_8734,N_8735);
nand U9193 (N_9193,N_8902,N_8839);
xor U9194 (N_9194,N_8968,N_8719);
nand U9195 (N_9195,N_8970,N_8841);
xnor U9196 (N_9196,N_8718,N_8795);
xnor U9197 (N_9197,N_8848,N_8989);
nor U9198 (N_9198,N_8920,N_8963);
or U9199 (N_9199,N_8874,N_8883);
or U9200 (N_9200,N_8810,N_8851);
or U9201 (N_9201,N_8855,N_8989);
nor U9202 (N_9202,N_8863,N_8898);
and U9203 (N_9203,N_8894,N_8810);
nor U9204 (N_9204,N_8998,N_8911);
and U9205 (N_9205,N_8714,N_8840);
nand U9206 (N_9206,N_8846,N_8950);
nor U9207 (N_9207,N_8764,N_8886);
nand U9208 (N_9208,N_8766,N_8868);
or U9209 (N_9209,N_8849,N_8826);
nand U9210 (N_9210,N_8771,N_8740);
and U9211 (N_9211,N_8948,N_8703);
xnor U9212 (N_9212,N_8908,N_8811);
nand U9213 (N_9213,N_8719,N_8810);
xor U9214 (N_9214,N_8731,N_8701);
and U9215 (N_9215,N_8944,N_8858);
xnor U9216 (N_9216,N_8939,N_8925);
xnor U9217 (N_9217,N_8745,N_8939);
nor U9218 (N_9218,N_8928,N_8888);
and U9219 (N_9219,N_8855,N_8952);
or U9220 (N_9220,N_8739,N_8711);
and U9221 (N_9221,N_8870,N_8960);
and U9222 (N_9222,N_8991,N_8796);
nor U9223 (N_9223,N_8761,N_8820);
or U9224 (N_9224,N_8878,N_8802);
and U9225 (N_9225,N_8978,N_8869);
nor U9226 (N_9226,N_8895,N_8865);
xor U9227 (N_9227,N_8944,N_8996);
or U9228 (N_9228,N_8823,N_8734);
nor U9229 (N_9229,N_8765,N_8817);
or U9230 (N_9230,N_8726,N_8729);
nand U9231 (N_9231,N_8999,N_8785);
or U9232 (N_9232,N_8898,N_8878);
nor U9233 (N_9233,N_8996,N_8882);
nand U9234 (N_9234,N_8804,N_8819);
or U9235 (N_9235,N_8978,N_8917);
nor U9236 (N_9236,N_8747,N_8890);
and U9237 (N_9237,N_8740,N_8916);
xnor U9238 (N_9238,N_8746,N_8732);
nand U9239 (N_9239,N_8989,N_8741);
and U9240 (N_9240,N_8851,N_8925);
xor U9241 (N_9241,N_8917,N_8868);
nor U9242 (N_9242,N_8765,N_8726);
and U9243 (N_9243,N_8766,N_8896);
xor U9244 (N_9244,N_8962,N_8963);
and U9245 (N_9245,N_8995,N_8806);
and U9246 (N_9246,N_8760,N_8711);
and U9247 (N_9247,N_8875,N_8883);
nor U9248 (N_9248,N_8712,N_8810);
or U9249 (N_9249,N_8706,N_8922);
and U9250 (N_9250,N_8795,N_8766);
nand U9251 (N_9251,N_8916,N_8793);
or U9252 (N_9252,N_8710,N_8884);
and U9253 (N_9253,N_8850,N_8716);
or U9254 (N_9254,N_8996,N_8777);
or U9255 (N_9255,N_8849,N_8932);
nand U9256 (N_9256,N_8750,N_8783);
and U9257 (N_9257,N_8977,N_8808);
and U9258 (N_9258,N_8831,N_8784);
nor U9259 (N_9259,N_8972,N_8950);
nand U9260 (N_9260,N_8956,N_8735);
or U9261 (N_9261,N_8717,N_8949);
or U9262 (N_9262,N_8730,N_8778);
or U9263 (N_9263,N_8826,N_8788);
nor U9264 (N_9264,N_8806,N_8879);
xor U9265 (N_9265,N_8790,N_8806);
or U9266 (N_9266,N_8966,N_8998);
or U9267 (N_9267,N_8796,N_8894);
nor U9268 (N_9268,N_8875,N_8784);
nand U9269 (N_9269,N_8759,N_8979);
and U9270 (N_9270,N_8784,N_8897);
xnor U9271 (N_9271,N_8902,N_8810);
xnor U9272 (N_9272,N_8701,N_8914);
nor U9273 (N_9273,N_8755,N_8977);
xor U9274 (N_9274,N_8840,N_8969);
and U9275 (N_9275,N_8773,N_8736);
nand U9276 (N_9276,N_8826,N_8830);
nor U9277 (N_9277,N_8909,N_8775);
or U9278 (N_9278,N_8780,N_8852);
nand U9279 (N_9279,N_8987,N_8806);
nor U9280 (N_9280,N_8973,N_8719);
xor U9281 (N_9281,N_8719,N_8938);
xor U9282 (N_9282,N_8832,N_8867);
nand U9283 (N_9283,N_8838,N_8958);
nor U9284 (N_9284,N_8939,N_8862);
or U9285 (N_9285,N_8913,N_8805);
and U9286 (N_9286,N_8843,N_8759);
or U9287 (N_9287,N_8737,N_8833);
xor U9288 (N_9288,N_8739,N_8759);
nor U9289 (N_9289,N_8724,N_8973);
nand U9290 (N_9290,N_8804,N_8908);
or U9291 (N_9291,N_8799,N_8972);
nor U9292 (N_9292,N_8879,N_8762);
xnor U9293 (N_9293,N_8707,N_8988);
xor U9294 (N_9294,N_8962,N_8739);
xnor U9295 (N_9295,N_8766,N_8840);
and U9296 (N_9296,N_8956,N_8808);
or U9297 (N_9297,N_8986,N_8728);
or U9298 (N_9298,N_8961,N_8718);
and U9299 (N_9299,N_8790,N_8864);
xor U9300 (N_9300,N_9161,N_9002);
xnor U9301 (N_9301,N_9063,N_9170);
and U9302 (N_9302,N_9009,N_9249);
or U9303 (N_9303,N_9213,N_9155);
nand U9304 (N_9304,N_9199,N_9119);
and U9305 (N_9305,N_9087,N_9089);
xnor U9306 (N_9306,N_9299,N_9158);
nand U9307 (N_9307,N_9215,N_9172);
xnor U9308 (N_9308,N_9032,N_9135);
or U9309 (N_9309,N_9064,N_9188);
and U9310 (N_9310,N_9148,N_9140);
nand U9311 (N_9311,N_9198,N_9273);
or U9312 (N_9312,N_9005,N_9131);
xor U9313 (N_9313,N_9256,N_9132);
xnor U9314 (N_9314,N_9151,N_9159);
or U9315 (N_9315,N_9065,N_9124);
and U9316 (N_9316,N_9157,N_9189);
nand U9317 (N_9317,N_9239,N_9283);
or U9318 (N_9318,N_9066,N_9056);
nor U9319 (N_9319,N_9220,N_9041);
nand U9320 (N_9320,N_9125,N_9275);
or U9321 (N_9321,N_9204,N_9060);
xor U9322 (N_9322,N_9141,N_9106);
xor U9323 (N_9323,N_9208,N_9218);
nand U9324 (N_9324,N_9296,N_9271);
or U9325 (N_9325,N_9209,N_9137);
and U9326 (N_9326,N_9045,N_9284);
xor U9327 (N_9327,N_9238,N_9136);
nand U9328 (N_9328,N_9112,N_9186);
or U9329 (N_9329,N_9200,N_9234);
or U9330 (N_9330,N_9242,N_9297);
or U9331 (N_9331,N_9054,N_9241);
nor U9332 (N_9332,N_9171,N_9192);
and U9333 (N_9333,N_9079,N_9026);
nand U9334 (N_9334,N_9232,N_9012);
xor U9335 (N_9335,N_9122,N_9103);
nand U9336 (N_9336,N_9235,N_9202);
or U9337 (N_9337,N_9207,N_9255);
nor U9338 (N_9338,N_9134,N_9016);
or U9339 (N_9339,N_9127,N_9197);
and U9340 (N_9340,N_9211,N_9260);
xnor U9341 (N_9341,N_9093,N_9014);
xor U9342 (N_9342,N_9034,N_9258);
nor U9343 (N_9343,N_9274,N_9084);
nand U9344 (N_9344,N_9292,N_9270);
and U9345 (N_9345,N_9115,N_9289);
or U9346 (N_9346,N_9264,N_9081);
nand U9347 (N_9347,N_9191,N_9225);
nand U9348 (N_9348,N_9048,N_9219);
and U9349 (N_9349,N_9183,N_9287);
xor U9350 (N_9350,N_9050,N_9227);
and U9351 (N_9351,N_9248,N_9099);
nand U9352 (N_9352,N_9243,N_9096);
xor U9353 (N_9353,N_9195,N_9182);
nor U9354 (N_9354,N_9261,N_9246);
nor U9355 (N_9355,N_9001,N_9163);
or U9356 (N_9356,N_9116,N_9031);
or U9357 (N_9357,N_9082,N_9147);
or U9358 (N_9358,N_9053,N_9166);
nand U9359 (N_9359,N_9250,N_9169);
nand U9360 (N_9360,N_9080,N_9088);
nor U9361 (N_9361,N_9092,N_9117);
nand U9362 (N_9362,N_9259,N_9187);
or U9363 (N_9363,N_9173,N_9111);
xnor U9364 (N_9364,N_9201,N_9049);
or U9365 (N_9365,N_9291,N_9196);
and U9366 (N_9366,N_9128,N_9279);
or U9367 (N_9367,N_9216,N_9105);
nor U9368 (N_9368,N_9098,N_9221);
nand U9369 (N_9369,N_9152,N_9280);
and U9370 (N_9370,N_9007,N_9162);
xnor U9371 (N_9371,N_9078,N_9013);
xor U9372 (N_9372,N_9091,N_9118);
and U9373 (N_9373,N_9214,N_9018);
and U9374 (N_9374,N_9010,N_9236);
and U9375 (N_9375,N_9203,N_9095);
or U9376 (N_9376,N_9130,N_9229);
nor U9377 (N_9377,N_9101,N_9073);
and U9378 (N_9378,N_9126,N_9177);
or U9379 (N_9379,N_9019,N_9046);
xor U9380 (N_9380,N_9193,N_9061);
or U9381 (N_9381,N_9097,N_9164);
xnor U9382 (N_9382,N_9022,N_9024);
nand U9383 (N_9383,N_9160,N_9100);
xnor U9384 (N_9384,N_9083,N_9120);
nand U9385 (N_9385,N_9020,N_9138);
and U9386 (N_9386,N_9068,N_9194);
nand U9387 (N_9387,N_9278,N_9206);
nor U9388 (N_9388,N_9165,N_9039);
nand U9389 (N_9389,N_9205,N_9228);
or U9390 (N_9390,N_9210,N_9003);
nor U9391 (N_9391,N_9000,N_9181);
xor U9392 (N_9392,N_9075,N_9174);
nor U9393 (N_9393,N_9047,N_9244);
nor U9394 (N_9394,N_9070,N_9176);
and U9395 (N_9395,N_9040,N_9231);
xnor U9396 (N_9396,N_9042,N_9153);
nand U9397 (N_9397,N_9129,N_9276);
and U9398 (N_9398,N_9245,N_9133);
nor U9399 (N_9399,N_9038,N_9017);
or U9400 (N_9400,N_9104,N_9254);
nor U9401 (N_9401,N_9036,N_9121);
xnor U9402 (N_9402,N_9108,N_9077);
nor U9403 (N_9403,N_9033,N_9251);
nand U9404 (N_9404,N_9051,N_9025);
xor U9405 (N_9405,N_9027,N_9156);
nor U9406 (N_9406,N_9142,N_9268);
or U9407 (N_9407,N_9110,N_9015);
and U9408 (N_9408,N_9272,N_9069);
or U9409 (N_9409,N_9233,N_9217);
nand U9410 (N_9410,N_9072,N_9146);
and U9411 (N_9411,N_9178,N_9113);
nand U9412 (N_9412,N_9269,N_9223);
nor U9413 (N_9413,N_9085,N_9253);
xor U9414 (N_9414,N_9257,N_9109);
or U9415 (N_9415,N_9175,N_9102);
nor U9416 (N_9416,N_9185,N_9252);
or U9417 (N_9417,N_9154,N_9190);
or U9418 (N_9418,N_9037,N_9028);
or U9419 (N_9419,N_9030,N_9298);
xor U9420 (N_9420,N_9145,N_9267);
nor U9421 (N_9421,N_9035,N_9044);
or U9422 (N_9422,N_9011,N_9179);
nor U9423 (N_9423,N_9230,N_9139);
nand U9424 (N_9424,N_9074,N_9094);
or U9425 (N_9425,N_9076,N_9168);
nor U9426 (N_9426,N_9237,N_9023);
and U9427 (N_9427,N_9290,N_9281);
and U9428 (N_9428,N_9240,N_9006);
nand U9429 (N_9429,N_9285,N_9150);
xor U9430 (N_9430,N_9057,N_9288);
or U9431 (N_9431,N_9167,N_9004);
xnor U9432 (N_9432,N_9262,N_9266);
or U9433 (N_9433,N_9282,N_9059);
xor U9434 (N_9434,N_9029,N_9071);
or U9435 (N_9435,N_9224,N_9184);
nor U9436 (N_9436,N_9058,N_9021);
and U9437 (N_9437,N_9090,N_9294);
and U9438 (N_9438,N_9295,N_9212);
nor U9439 (N_9439,N_9247,N_9143);
xor U9440 (N_9440,N_9055,N_9222);
nor U9441 (N_9441,N_9277,N_9149);
nor U9442 (N_9442,N_9226,N_9008);
nor U9443 (N_9443,N_9144,N_9114);
xor U9444 (N_9444,N_9180,N_9265);
xor U9445 (N_9445,N_9062,N_9086);
nor U9446 (N_9446,N_9043,N_9067);
nand U9447 (N_9447,N_9263,N_9107);
nor U9448 (N_9448,N_9052,N_9286);
nor U9449 (N_9449,N_9123,N_9293);
and U9450 (N_9450,N_9279,N_9275);
nor U9451 (N_9451,N_9236,N_9090);
nand U9452 (N_9452,N_9290,N_9129);
nand U9453 (N_9453,N_9213,N_9160);
nor U9454 (N_9454,N_9278,N_9031);
nor U9455 (N_9455,N_9226,N_9157);
or U9456 (N_9456,N_9181,N_9054);
and U9457 (N_9457,N_9265,N_9198);
xnor U9458 (N_9458,N_9080,N_9172);
or U9459 (N_9459,N_9060,N_9158);
and U9460 (N_9460,N_9008,N_9235);
and U9461 (N_9461,N_9139,N_9218);
nand U9462 (N_9462,N_9129,N_9173);
or U9463 (N_9463,N_9227,N_9248);
and U9464 (N_9464,N_9183,N_9219);
nor U9465 (N_9465,N_9294,N_9116);
and U9466 (N_9466,N_9245,N_9093);
and U9467 (N_9467,N_9036,N_9279);
xnor U9468 (N_9468,N_9254,N_9227);
nor U9469 (N_9469,N_9135,N_9231);
or U9470 (N_9470,N_9044,N_9019);
or U9471 (N_9471,N_9104,N_9142);
nand U9472 (N_9472,N_9239,N_9023);
xor U9473 (N_9473,N_9166,N_9018);
xnor U9474 (N_9474,N_9045,N_9078);
nor U9475 (N_9475,N_9234,N_9101);
nor U9476 (N_9476,N_9065,N_9057);
and U9477 (N_9477,N_9187,N_9224);
xor U9478 (N_9478,N_9186,N_9048);
and U9479 (N_9479,N_9014,N_9274);
nor U9480 (N_9480,N_9116,N_9150);
nor U9481 (N_9481,N_9192,N_9233);
nand U9482 (N_9482,N_9201,N_9279);
and U9483 (N_9483,N_9258,N_9288);
or U9484 (N_9484,N_9125,N_9069);
nor U9485 (N_9485,N_9248,N_9068);
or U9486 (N_9486,N_9039,N_9164);
nor U9487 (N_9487,N_9139,N_9172);
xor U9488 (N_9488,N_9250,N_9144);
xor U9489 (N_9489,N_9001,N_9201);
nor U9490 (N_9490,N_9144,N_9207);
or U9491 (N_9491,N_9240,N_9071);
xor U9492 (N_9492,N_9113,N_9159);
nor U9493 (N_9493,N_9049,N_9070);
xor U9494 (N_9494,N_9199,N_9220);
nand U9495 (N_9495,N_9237,N_9095);
nand U9496 (N_9496,N_9133,N_9257);
nor U9497 (N_9497,N_9294,N_9298);
nor U9498 (N_9498,N_9289,N_9000);
nor U9499 (N_9499,N_9019,N_9255);
nand U9500 (N_9500,N_9207,N_9093);
nor U9501 (N_9501,N_9179,N_9240);
xnor U9502 (N_9502,N_9200,N_9221);
nor U9503 (N_9503,N_9198,N_9148);
nand U9504 (N_9504,N_9174,N_9057);
or U9505 (N_9505,N_9134,N_9084);
nand U9506 (N_9506,N_9050,N_9140);
and U9507 (N_9507,N_9276,N_9055);
nand U9508 (N_9508,N_9208,N_9061);
or U9509 (N_9509,N_9037,N_9000);
xnor U9510 (N_9510,N_9110,N_9279);
nor U9511 (N_9511,N_9147,N_9205);
and U9512 (N_9512,N_9151,N_9055);
nand U9513 (N_9513,N_9252,N_9223);
xor U9514 (N_9514,N_9059,N_9145);
nand U9515 (N_9515,N_9261,N_9126);
xnor U9516 (N_9516,N_9093,N_9160);
or U9517 (N_9517,N_9090,N_9003);
and U9518 (N_9518,N_9128,N_9280);
nor U9519 (N_9519,N_9008,N_9149);
nand U9520 (N_9520,N_9151,N_9007);
nor U9521 (N_9521,N_9271,N_9149);
nor U9522 (N_9522,N_9059,N_9104);
or U9523 (N_9523,N_9182,N_9119);
or U9524 (N_9524,N_9116,N_9202);
nor U9525 (N_9525,N_9287,N_9053);
or U9526 (N_9526,N_9058,N_9281);
and U9527 (N_9527,N_9158,N_9217);
or U9528 (N_9528,N_9134,N_9151);
and U9529 (N_9529,N_9183,N_9048);
nor U9530 (N_9530,N_9200,N_9223);
nor U9531 (N_9531,N_9150,N_9230);
or U9532 (N_9532,N_9046,N_9276);
nor U9533 (N_9533,N_9255,N_9036);
nor U9534 (N_9534,N_9234,N_9057);
nor U9535 (N_9535,N_9234,N_9072);
nor U9536 (N_9536,N_9245,N_9019);
nor U9537 (N_9537,N_9068,N_9266);
nand U9538 (N_9538,N_9020,N_9063);
xnor U9539 (N_9539,N_9102,N_9053);
nand U9540 (N_9540,N_9242,N_9052);
xor U9541 (N_9541,N_9127,N_9240);
or U9542 (N_9542,N_9287,N_9012);
xor U9543 (N_9543,N_9083,N_9172);
nand U9544 (N_9544,N_9006,N_9252);
nand U9545 (N_9545,N_9019,N_9027);
or U9546 (N_9546,N_9048,N_9090);
or U9547 (N_9547,N_9204,N_9008);
or U9548 (N_9548,N_9072,N_9175);
nand U9549 (N_9549,N_9115,N_9145);
xor U9550 (N_9550,N_9240,N_9187);
xnor U9551 (N_9551,N_9204,N_9023);
nor U9552 (N_9552,N_9062,N_9053);
or U9553 (N_9553,N_9200,N_9027);
nor U9554 (N_9554,N_9172,N_9073);
and U9555 (N_9555,N_9227,N_9190);
and U9556 (N_9556,N_9186,N_9129);
or U9557 (N_9557,N_9100,N_9233);
xnor U9558 (N_9558,N_9101,N_9261);
xor U9559 (N_9559,N_9108,N_9290);
xnor U9560 (N_9560,N_9043,N_9177);
xnor U9561 (N_9561,N_9272,N_9164);
nand U9562 (N_9562,N_9093,N_9299);
nand U9563 (N_9563,N_9262,N_9257);
nor U9564 (N_9564,N_9176,N_9253);
xor U9565 (N_9565,N_9141,N_9161);
nand U9566 (N_9566,N_9281,N_9232);
nand U9567 (N_9567,N_9147,N_9284);
nor U9568 (N_9568,N_9202,N_9064);
nand U9569 (N_9569,N_9138,N_9128);
nand U9570 (N_9570,N_9051,N_9289);
or U9571 (N_9571,N_9137,N_9242);
xor U9572 (N_9572,N_9070,N_9254);
and U9573 (N_9573,N_9268,N_9201);
xnor U9574 (N_9574,N_9146,N_9174);
and U9575 (N_9575,N_9176,N_9285);
nor U9576 (N_9576,N_9060,N_9057);
nor U9577 (N_9577,N_9137,N_9153);
and U9578 (N_9578,N_9217,N_9059);
or U9579 (N_9579,N_9150,N_9090);
nor U9580 (N_9580,N_9132,N_9172);
nand U9581 (N_9581,N_9166,N_9179);
and U9582 (N_9582,N_9180,N_9272);
xnor U9583 (N_9583,N_9147,N_9165);
nor U9584 (N_9584,N_9149,N_9124);
or U9585 (N_9585,N_9027,N_9211);
xnor U9586 (N_9586,N_9056,N_9115);
nor U9587 (N_9587,N_9050,N_9186);
nand U9588 (N_9588,N_9183,N_9189);
or U9589 (N_9589,N_9057,N_9163);
nand U9590 (N_9590,N_9043,N_9159);
nor U9591 (N_9591,N_9217,N_9281);
or U9592 (N_9592,N_9007,N_9050);
xor U9593 (N_9593,N_9273,N_9279);
xor U9594 (N_9594,N_9096,N_9144);
xor U9595 (N_9595,N_9197,N_9047);
nand U9596 (N_9596,N_9259,N_9082);
nand U9597 (N_9597,N_9173,N_9238);
and U9598 (N_9598,N_9015,N_9274);
or U9599 (N_9599,N_9115,N_9000);
nand U9600 (N_9600,N_9377,N_9473);
or U9601 (N_9601,N_9302,N_9443);
nor U9602 (N_9602,N_9332,N_9487);
xnor U9603 (N_9603,N_9540,N_9499);
nor U9604 (N_9604,N_9305,N_9368);
xor U9605 (N_9605,N_9543,N_9406);
nand U9606 (N_9606,N_9585,N_9347);
and U9607 (N_9607,N_9574,N_9433);
xnor U9608 (N_9608,N_9388,N_9333);
nand U9609 (N_9609,N_9599,N_9519);
or U9610 (N_9610,N_9355,N_9399);
nand U9611 (N_9611,N_9530,N_9568);
nand U9612 (N_9612,N_9589,N_9515);
or U9613 (N_9613,N_9314,N_9549);
xnor U9614 (N_9614,N_9538,N_9509);
nor U9615 (N_9615,N_9490,N_9358);
or U9616 (N_9616,N_9409,N_9430);
nand U9617 (N_9617,N_9576,N_9571);
or U9618 (N_9618,N_9553,N_9348);
or U9619 (N_9619,N_9491,N_9466);
and U9620 (N_9620,N_9437,N_9391);
or U9621 (N_9621,N_9455,N_9337);
xnor U9622 (N_9622,N_9563,N_9582);
xnor U9623 (N_9623,N_9431,N_9457);
xnor U9624 (N_9624,N_9422,N_9590);
nor U9625 (N_9625,N_9322,N_9504);
or U9626 (N_9626,N_9480,N_9415);
or U9627 (N_9627,N_9561,N_9407);
or U9628 (N_9628,N_9526,N_9463);
and U9629 (N_9629,N_9336,N_9313);
nand U9630 (N_9630,N_9343,N_9339);
and U9631 (N_9631,N_9379,N_9566);
nor U9632 (N_9632,N_9350,N_9303);
nand U9633 (N_9633,N_9570,N_9334);
and U9634 (N_9634,N_9465,N_9342);
or U9635 (N_9635,N_9307,N_9488);
or U9636 (N_9636,N_9572,N_9482);
nor U9637 (N_9637,N_9500,N_9469);
nor U9638 (N_9638,N_9554,N_9479);
nor U9639 (N_9639,N_9395,N_9414);
nand U9640 (N_9640,N_9575,N_9529);
and U9641 (N_9641,N_9468,N_9360);
or U9642 (N_9642,N_9310,N_9592);
and U9643 (N_9643,N_9489,N_9412);
or U9644 (N_9644,N_9404,N_9581);
or U9645 (N_9645,N_9435,N_9387);
nand U9646 (N_9646,N_9375,N_9595);
nand U9647 (N_9647,N_9361,N_9386);
and U9648 (N_9648,N_9493,N_9579);
and U9649 (N_9649,N_9472,N_9384);
xor U9650 (N_9650,N_9506,N_9486);
and U9651 (N_9651,N_9382,N_9419);
or U9652 (N_9652,N_9418,N_9319);
xor U9653 (N_9653,N_9309,N_9359);
nor U9654 (N_9654,N_9567,N_9555);
xnor U9655 (N_9655,N_9328,N_9356);
nor U9656 (N_9656,N_9536,N_9380);
and U9657 (N_9657,N_9312,N_9428);
nor U9658 (N_9658,N_9338,N_9373);
nand U9659 (N_9659,N_9442,N_9496);
nor U9660 (N_9660,N_9531,N_9545);
or U9661 (N_9661,N_9454,N_9459);
xor U9662 (N_9662,N_9453,N_9548);
or U9663 (N_9663,N_9357,N_9478);
nor U9664 (N_9664,N_9335,N_9432);
or U9665 (N_9665,N_9315,N_9485);
and U9666 (N_9666,N_9370,N_9378);
xor U9667 (N_9667,N_9346,N_9522);
nand U9668 (N_9668,N_9492,N_9362);
and U9669 (N_9669,N_9341,N_9318);
and U9670 (N_9670,N_9525,N_9301);
xor U9671 (N_9671,N_9327,N_9573);
xnor U9672 (N_9672,N_9476,N_9441);
nor U9673 (N_9673,N_9446,N_9507);
nand U9674 (N_9674,N_9401,N_9405);
xnor U9675 (N_9675,N_9411,N_9367);
or U9676 (N_9676,N_9546,N_9474);
nor U9677 (N_9677,N_9577,N_9400);
xnor U9678 (N_9678,N_9593,N_9300);
nor U9679 (N_9679,N_9340,N_9591);
or U9680 (N_9680,N_9528,N_9539);
and U9681 (N_9681,N_9532,N_9452);
and U9682 (N_9682,N_9512,N_9505);
or U9683 (N_9683,N_9304,N_9330);
nor U9684 (N_9684,N_9521,N_9436);
and U9685 (N_9685,N_9434,N_9510);
nor U9686 (N_9686,N_9502,N_9456);
nand U9687 (N_9687,N_9320,N_9393);
or U9688 (N_9688,N_9578,N_9584);
and U9689 (N_9689,N_9494,N_9326);
nor U9690 (N_9690,N_9403,N_9503);
nand U9691 (N_9691,N_9547,N_9583);
and U9692 (N_9692,N_9523,N_9475);
and U9693 (N_9693,N_9449,N_9402);
and U9694 (N_9694,N_9349,N_9481);
xnor U9695 (N_9695,N_9438,N_9383);
and U9696 (N_9696,N_9381,N_9439);
nand U9697 (N_9697,N_9324,N_9596);
and U9698 (N_9698,N_9413,N_9535);
or U9699 (N_9699,N_9483,N_9417);
xnor U9700 (N_9700,N_9564,N_9559);
nand U9701 (N_9701,N_9464,N_9560);
nor U9702 (N_9702,N_9524,N_9440);
xnor U9703 (N_9703,N_9558,N_9448);
xor U9704 (N_9704,N_9467,N_9408);
xor U9705 (N_9705,N_9533,N_9534);
nor U9706 (N_9706,N_9508,N_9557);
nand U9707 (N_9707,N_9562,N_9484);
nand U9708 (N_9708,N_9598,N_9372);
nand U9709 (N_9709,N_9353,N_9451);
or U9710 (N_9710,N_9323,N_9477);
and U9711 (N_9711,N_9364,N_9392);
and U9712 (N_9712,N_9369,N_9351);
nor U9713 (N_9713,N_9321,N_9552);
and U9714 (N_9714,N_9447,N_9420);
or U9715 (N_9715,N_9462,N_9498);
and U9716 (N_9716,N_9354,N_9421);
and U9717 (N_9717,N_9363,N_9471);
nand U9718 (N_9718,N_9365,N_9565);
or U9719 (N_9719,N_9513,N_9556);
nor U9720 (N_9720,N_9345,N_9344);
nor U9721 (N_9721,N_9308,N_9423);
or U9722 (N_9722,N_9394,N_9325);
or U9723 (N_9723,N_9317,N_9410);
and U9724 (N_9724,N_9374,N_9416);
or U9725 (N_9725,N_9517,N_9429);
or U9726 (N_9726,N_9569,N_9425);
or U9727 (N_9727,N_9397,N_9588);
and U9728 (N_9728,N_9514,N_9376);
nor U9729 (N_9729,N_9461,N_9389);
nand U9730 (N_9730,N_9501,N_9424);
nor U9731 (N_9731,N_9470,N_9390);
or U9732 (N_9732,N_9580,N_9366);
or U9733 (N_9733,N_9371,N_9311);
nand U9734 (N_9734,N_9597,N_9396);
nand U9735 (N_9735,N_9551,N_9520);
nand U9736 (N_9736,N_9427,N_9398);
nor U9737 (N_9737,N_9586,N_9306);
and U9738 (N_9738,N_9587,N_9426);
or U9739 (N_9739,N_9542,N_9444);
nand U9740 (N_9740,N_9550,N_9495);
nand U9741 (N_9741,N_9594,N_9331);
nor U9742 (N_9742,N_9445,N_9385);
nor U9743 (N_9743,N_9458,N_9460);
or U9744 (N_9744,N_9497,N_9518);
and U9745 (N_9745,N_9527,N_9544);
or U9746 (N_9746,N_9511,N_9316);
nor U9747 (N_9747,N_9450,N_9352);
xor U9748 (N_9748,N_9541,N_9329);
or U9749 (N_9749,N_9537,N_9516);
and U9750 (N_9750,N_9563,N_9595);
xor U9751 (N_9751,N_9362,N_9491);
and U9752 (N_9752,N_9348,N_9349);
nor U9753 (N_9753,N_9582,N_9357);
nor U9754 (N_9754,N_9330,N_9433);
xnor U9755 (N_9755,N_9500,N_9379);
nand U9756 (N_9756,N_9413,N_9443);
and U9757 (N_9757,N_9406,N_9410);
nor U9758 (N_9758,N_9333,N_9498);
nor U9759 (N_9759,N_9337,N_9565);
and U9760 (N_9760,N_9354,N_9395);
xnor U9761 (N_9761,N_9453,N_9483);
nor U9762 (N_9762,N_9379,N_9504);
and U9763 (N_9763,N_9538,N_9361);
xor U9764 (N_9764,N_9422,N_9466);
nor U9765 (N_9765,N_9314,N_9564);
xnor U9766 (N_9766,N_9363,N_9313);
xnor U9767 (N_9767,N_9512,N_9388);
nor U9768 (N_9768,N_9390,N_9374);
xnor U9769 (N_9769,N_9462,N_9511);
or U9770 (N_9770,N_9450,N_9302);
nor U9771 (N_9771,N_9403,N_9480);
nor U9772 (N_9772,N_9520,N_9594);
or U9773 (N_9773,N_9542,N_9490);
nor U9774 (N_9774,N_9379,N_9442);
nor U9775 (N_9775,N_9515,N_9330);
xnor U9776 (N_9776,N_9332,N_9562);
or U9777 (N_9777,N_9477,N_9409);
xor U9778 (N_9778,N_9400,N_9319);
nand U9779 (N_9779,N_9329,N_9449);
nand U9780 (N_9780,N_9400,N_9362);
and U9781 (N_9781,N_9548,N_9434);
or U9782 (N_9782,N_9498,N_9325);
and U9783 (N_9783,N_9327,N_9537);
and U9784 (N_9784,N_9399,N_9553);
xor U9785 (N_9785,N_9405,N_9335);
xnor U9786 (N_9786,N_9444,N_9504);
xnor U9787 (N_9787,N_9308,N_9465);
and U9788 (N_9788,N_9342,N_9365);
or U9789 (N_9789,N_9485,N_9423);
or U9790 (N_9790,N_9391,N_9420);
and U9791 (N_9791,N_9552,N_9467);
xor U9792 (N_9792,N_9359,N_9454);
nor U9793 (N_9793,N_9586,N_9465);
nor U9794 (N_9794,N_9508,N_9439);
or U9795 (N_9795,N_9500,N_9400);
nand U9796 (N_9796,N_9582,N_9488);
or U9797 (N_9797,N_9459,N_9496);
and U9798 (N_9798,N_9351,N_9587);
xor U9799 (N_9799,N_9516,N_9587);
nor U9800 (N_9800,N_9313,N_9302);
and U9801 (N_9801,N_9433,N_9415);
nand U9802 (N_9802,N_9539,N_9546);
and U9803 (N_9803,N_9564,N_9441);
and U9804 (N_9804,N_9436,N_9450);
nand U9805 (N_9805,N_9533,N_9423);
xor U9806 (N_9806,N_9454,N_9394);
nor U9807 (N_9807,N_9365,N_9555);
nand U9808 (N_9808,N_9558,N_9338);
or U9809 (N_9809,N_9311,N_9472);
nor U9810 (N_9810,N_9332,N_9375);
nand U9811 (N_9811,N_9519,N_9553);
and U9812 (N_9812,N_9494,N_9397);
nor U9813 (N_9813,N_9307,N_9535);
or U9814 (N_9814,N_9437,N_9483);
or U9815 (N_9815,N_9563,N_9456);
or U9816 (N_9816,N_9363,N_9482);
or U9817 (N_9817,N_9412,N_9541);
or U9818 (N_9818,N_9516,N_9573);
nand U9819 (N_9819,N_9400,N_9456);
xnor U9820 (N_9820,N_9537,N_9444);
xnor U9821 (N_9821,N_9472,N_9416);
nand U9822 (N_9822,N_9481,N_9344);
xor U9823 (N_9823,N_9345,N_9337);
nand U9824 (N_9824,N_9519,N_9592);
xnor U9825 (N_9825,N_9485,N_9345);
or U9826 (N_9826,N_9426,N_9374);
or U9827 (N_9827,N_9301,N_9530);
nor U9828 (N_9828,N_9391,N_9523);
nor U9829 (N_9829,N_9587,N_9576);
or U9830 (N_9830,N_9378,N_9328);
nor U9831 (N_9831,N_9372,N_9440);
and U9832 (N_9832,N_9598,N_9446);
nor U9833 (N_9833,N_9383,N_9414);
or U9834 (N_9834,N_9313,N_9331);
and U9835 (N_9835,N_9306,N_9533);
xnor U9836 (N_9836,N_9516,N_9320);
or U9837 (N_9837,N_9488,N_9381);
nor U9838 (N_9838,N_9318,N_9378);
xor U9839 (N_9839,N_9349,N_9594);
xnor U9840 (N_9840,N_9437,N_9349);
and U9841 (N_9841,N_9369,N_9334);
and U9842 (N_9842,N_9389,N_9525);
nor U9843 (N_9843,N_9473,N_9517);
or U9844 (N_9844,N_9519,N_9305);
nand U9845 (N_9845,N_9374,N_9542);
nor U9846 (N_9846,N_9574,N_9410);
or U9847 (N_9847,N_9398,N_9311);
nand U9848 (N_9848,N_9416,N_9585);
and U9849 (N_9849,N_9312,N_9378);
and U9850 (N_9850,N_9428,N_9557);
nor U9851 (N_9851,N_9476,N_9416);
nor U9852 (N_9852,N_9508,N_9468);
xnor U9853 (N_9853,N_9386,N_9330);
and U9854 (N_9854,N_9477,N_9560);
and U9855 (N_9855,N_9478,N_9387);
nand U9856 (N_9856,N_9334,N_9396);
nor U9857 (N_9857,N_9505,N_9573);
and U9858 (N_9858,N_9464,N_9382);
and U9859 (N_9859,N_9583,N_9559);
nor U9860 (N_9860,N_9513,N_9516);
nor U9861 (N_9861,N_9421,N_9394);
and U9862 (N_9862,N_9402,N_9420);
xor U9863 (N_9863,N_9570,N_9598);
and U9864 (N_9864,N_9329,N_9495);
or U9865 (N_9865,N_9391,N_9379);
and U9866 (N_9866,N_9567,N_9326);
nand U9867 (N_9867,N_9593,N_9597);
nor U9868 (N_9868,N_9548,N_9501);
nor U9869 (N_9869,N_9545,N_9580);
nor U9870 (N_9870,N_9373,N_9349);
nand U9871 (N_9871,N_9425,N_9308);
nor U9872 (N_9872,N_9466,N_9312);
xor U9873 (N_9873,N_9475,N_9591);
and U9874 (N_9874,N_9579,N_9431);
or U9875 (N_9875,N_9396,N_9585);
nor U9876 (N_9876,N_9405,N_9339);
xor U9877 (N_9877,N_9361,N_9413);
and U9878 (N_9878,N_9433,N_9591);
or U9879 (N_9879,N_9545,N_9342);
nand U9880 (N_9880,N_9311,N_9532);
and U9881 (N_9881,N_9408,N_9539);
nor U9882 (N_9882,N_9353,N_9490);
nor U9883 (N_9883,N_9547,N_9322);
and U9884 (N_9884,N_9302,N_9354);
xnor U9885 (N_9885,N_9423,N_9419);
or U9886 (N_9886,N_9518,N_9413);
nor U9887 (N_9887,N_9552,N_9477);
xor U9888 (N_9888,N_9492,N_9385);
nand U9889 (N_9889,N_9400,N_9315);
xor U9890 (N_9890,N_9490,N_9540);
nand U9891 (N_9891,N_9420,N_9466);
and U9892 (N_9892,N_9329,N_9526);
and U9893 (N_9893,N_9300,N_9421);
or U9894 (N_9894,N_9587,N_9524);
nor U9895 (N_9895,N_9435,N_9348);
or U9896 (N_9896,N_9414,N_9546);
or U9897 (N_9897,N_9497,N_9367);
nand U9898 (N_9898,N_9357,N_9483);
nor U9899 (N_9899,N_9565,N_9305);
or U9900 (N_9900,N_9803,N_9667);
nor U9901 (N_9901,N_9778,N_9899);
xnor U9902 (N_9902,N_9807,N_9631);
nand U9903 (N_9903,N_9616,N_9830);
and U9904 (N_9904,N_9756,N_9892);
and U9905 (N_9905,N_9619,N_9841);
nand U9906 (N_9906,N_9896,N_9883);
or U9907 (N_9907,N_9638,N_9708);
nor U9908 (N_9908,N_9767,N_9663);
nor U9909 (N_9909,N_9664,N_9866);
nand U9910 (N_9910,N_9763,N_9820);
nor U9911 (N_9911,N_9831,N_9683);
xor U9912 (N_9912,N_9810,N_9688);
and U9913 (N_9913,N_9797,N_9684);
xnor U9914 (N_9914,N_9709,N_9702);
and U9915 (N_9915,N_9698,N_9605);
xnor U9916 (N_9916,N_9718,N_9855);
nor U9917 (N_9917,N_9791,N_9719);
xor U9918 (N_9918,N_9827,N_9865);
nand U9919 (N_9919,N_9736,N_9644);
or U9920 (N_9920,N_9660,N_9705);
nor U9921 (N_9921,N_9732,N_9861);
nor U9922 (N_9922,N_9801,N_9781);
nor U9923 (N_9923,N_9824,N_9700);
xnor U9924 (N_9924,N_9670,N_9628);
or U9925 (N_9925,N_9601,N_9787);
and U9926 (N_9926,N_9617,N_9838);
nand U9927 (N_9927,N_9757,N_9868);
xor U9928 (N_9928,N_9615,N_9706);
nand U9929 (N_9929,N_9761,N_9893);
nand U9930 (N_9930,N_9730,N_9879);
nor U9931 (N_9931,N_9654,N_9877);
nand U9932 (N_9932,N_9720,N_9884);
xor U9933 (N_9933,N_9834,N_9607);
nor U9934 (N_9934,N_9612,N_9783);
nor U9935 (N_9935,N_9737,N_9898);
nor U9936 (N_9936,N_9739,N_9669);
or U9937 (N_9937,N_9673,N_9792);
nand U9938 (N_9938,N_9755,N_9740);
and U9939 (N_9939,N_9859,N_9746);
nand U9940 (N_9940,N_9864,N_9817);
nand U9941 (N_9941,N_9774,N_9636);
or U9942 (N_9942,N_9657,N_9687);
and U9943 (N_9943,N_9871,N_9745);
nand U9944 (N_9944,N_9742,N_9848);
or U9945 (N_9945,N_9776,N_9637);
nand U9946 (N_9946,N_9710,N_9693);
nand U9947 (N_9947,N_9701,N_9875);
or U9948 (N_9948,N_9729,N_9680);
nor U9949 (N_9949,N_9852,N_9895);
nand U9950 (N_9950,N_9651,N_9798);
or U9951 (N_9951,N_9695,N_9675);
and U9952 (N_9952,N_9629,N_9794);
xor U9953 (N_9953,N_9823,N_9854);
and U9954 (N_9954,N_9788,N_9839);
nand U9955 (N_9955,N_9816,N_9885);
nand U9956 (N_9956,N_9785,N_9840);
or U9957 (N_9957,N_9608,N_9773);
xor U9958 (N_9958,N_9799,N_9843);
xnor U9959 (N_9959,N_9743,N_9822);
or U9960 (N_9960,N_9818,N_9749);
nand U9961 (N_9961,N_9647,N_9775);
nand U9962 (N_9962,N_9751,N_9815);
nand U9963 (N_9963,N_9727,N_9639);
nor U9964 (N_9964,N_9829,N_9672);
and U9965 (N_9965,N_9626,N_9766);
nand U9966 (N_9966,N_9836,N_9802);
nor U9967 (N_9967,N_9635,N_9860);
nand U9968 (N_9968,N_9658,N_9741);
nor U9969 (N_9969,N_9849,N_9624);
xnor U9970 (N_9970,N_9845,N_9846);
nand U9971 (N_9971,N_9808,N_9665);
xor U9972 (N_9972,N_9640,N_9691);
and U9973 (N_9973,N_9677,N_9867);
nor U9974 (N_9974,N_9880,N_9876);
or U9975 (N_9975,N_9645,N_9887);
and U9976 (N_9976,N_9717,N_9721);
xnor U9977 (N_9977,N_9873,N_9796);
nand U9978 (N_9978,N_9851,N_9704);
nor U9979 (N_9979,N_9857,N_9770);
nand U9980 (N_9980,N_9800,N_9678);
xnor U9981 (N_9981,N_9835,N_9814);
or U9982 (N_9982,N_9881,N_9804);
or U9983 (N_9983,N_9622,N_9768);
or U9984 (N_9984,N_9703,N_9837);
or U9985 (N_9985,N_9809,N_9692);
or U9986 (N_9986,N_9805,N_9643);
nor U9987 (N_9987,N_9627,N_9652);
xor U9988 (N_9988,N_9689,N_9784);
nor U9989 (N_9989,N_9646,N_9681);
or U9990 (N_9990,N_9793,N_9878);
nand U9991 (N_9991,N_9610,N_9782);
nor U9992 (N_9992,N_9850,N_9754);
nand U9993 (N_9993,N_9641,N_9869);
nor U9994 (N_9994,N_9603,N_9762);
nand U9995 (N_9995,N_9716,N_9712);
or U9996 (N_9996,N_9630,N_9733);
and U9997 (N_9997,N_9696,N_9890);
and U9998 (N_9998,N_9750,N_9600);
xor U9999 (N_9999,N_9725,N_9602);
or U10000 (N_10000,N_9795,N_9694);
xor U10001 (N_10001,N_9889,N_9894);
nand U10002 (N_10002,N_9697,N_9772);
nand U10003 (N_10003,N_9613,N_9790);
nor U10004 (N_10004,N_9886,N_9847);
nand U10005 (N_10005,N_9711,N_9726);
xor U10006 (N_10006,N_9786,N_9806);
and U10007 (N_10007,N_9633,N_9819);
xor U10008 (N_10008,N_9826,N_9874);
nand U10009 (N_10009,N_9780,N_9611);
xor U10010 (N_10010,N_9833,N_9655);
nor U10011 (N_10011,N_9666,N_9744);
and U10012 (N_10012,N_9648,N_9724);
xnor U10013 (N_10013,N_9862,N_9812);
xnor U10014 (N_10014,N_9623,N_9858);
nor U10015 (N_10015,N_9759,N_9625);
nand U10016 (N_10016,N_9609,N_9882);
nand U10017 (N_10017,N_9738,N_9752);
xnor U10018 (N_10018,N_9606,N_9811);
nor U10019 (N_10019,N_9722,N_9813);
nand U10020 (N_10020,N_9735,N_9789);
nor U10021 (N_10021,N_9671,N_9656);
or U10022 (N_10022,N_9604,N_9614);
nor U10023 (N_10023,N_9707,N_9821);
nand U10024 (N_10024,N_9753,N_9779);
xor U10025 (N_10025,N_9621,N_9828);
nor U10026 (N_10026,N_9897,N_9699);
or U10027 (N_10027,N_9714,N_9825);
nand U10028 (N_10028,N_9760,N_9679);
and U10029 (N_10029,N_9734,N_9674);
nor U10030 (N_10030,N_9662,N_9765);
nor U10031 (N_10031,N_9856,N_9891);
or U10032 (N_10032,N_9642,N_9769);
nor U10033 (N_10033,N_9650,N_9853);
or U10034 (N_10034,N_9676,N_9888);
nor U10035 (N_10035,N_9872,N_9863);
and U10036 (N_10036,N_9668,N_9842);
nand U10037 (N_10037,N_9685,N_9686);
nand U10038 (N_10038,N_9682,N_9713);
and U10039 (N_10039,N_9832,N_9747);
xor U10040 (N_10040,N_9748,N_9731);
nor U10041 (N_10041,N_9618,N_9715);
xnor U10042 (N_10042,N_9690,N_9653);
or U10043 (N_10043,N_9661,N_9659);
nand U10044 (N_10044,N_9764,N_9771);
or U10045 (N_10045,N_9620,N_9723);
xor U10046 (N_10046,N_9728,N_9777);
or U10047 (N_10047,N_9870,N_9844);
nand U10048 (N_10048,N_9634,N_9632);
nor U10049 (N_10049,N_9758,N_9649);
nor U10050 (N_10050,N_9723,N_9784);
nand U10051 (N_10051,N_9825,N_9785);
and U10052 (N_10052,N_9620,N_9887);
or U10053 (N_10053,N_9619,N_9804);
nor U10054 (N_10054,N_9784,N_9827);
nand U10055 (N_10055,N_9730,N_9790);
nand U10056 (N_10056,N_9706,N_9666);
nor U10057 (N_10057,N_9619,N_9807);
or U10058 (N_10058,N_9686,N_9605);
nand U10059 (N_10059,N_9886,N_9633);
and U10060 (N_10060,N_9601,N_9766);
xor U10061 (N_10061,N_9726,N_9738);
or U10062 (N_10062,N_9792,N_9629);
nand U10063 (N_10063,N_9892,N_9776);
or U10064 (N_10064,N_9743,N_9884);
xor U10065 (N_10065,N_9776,N_9875);
nor U10066 (N_10066,N_9733,N_9646);
nor U10067 (N_10067,N_9765,N_9852);
or U10068 (N_10068,N_9638,N_9687);
nand U10069 (N_10069,N_9738,N_9716);
nand U10070 (N_10070,N_9812,N_9754);
or U10071 (N_10071,N_9613,N_9741);
nand U10072 (N_10072,N_9849,N_9820);
and U10073 (N_10073,N_9776,N_9680);
nand U10074 (N_10074,N_9795,N_9887);
and U10075 (N_10075,N_9844,N_9858);
nor U10076 (N_10076,N_9775,N_9756);
xnor U10077 (N_10077,N_9709,N_9758);
or U10078 (N_10078,N_9684,N_9740);
nand U10079 (N_10079,N_9607,N_9792);
and U10080 (N_10080,N_9668,N_9822);
nor U10081 (N_10081,N_9797,N_9830);
and U10082 (N_10082,N_9756,N_9835);
or U10083 (N_10083,N_9854,N_9841);
and U10084 (N_10084,N_9629,N_9782);
or U10085 (N_10085,N_9742,N_9702);
xnor U10086 (N_10086,N_9755,N_9750);
nand U10087 (N_10087,N_9856,N_9635);
and U10088 (N_10088,N_9687,N_9815);
nor U10089 (N_10089,N_9739,N_9699);
nand U10090 (N_10090,N_9632,N_9654);
or U10091 (N_10091,N_9827,N_9860);
xor U10092 (N_10092,N_9875,N_9755);
or U10093 (N_10093,N_9785,N_9853);
and U10094 (N_10094,N_9613,N_9660);
nand U10095 (N_10095,N_9757,N_9670);
or U10096 (N_10096,N_9787,N_9863);
or U10097 (N_10097,N_9687,N_9748);
xnor U10098 (N_10098,N_9690,N_9891);
and U10099 (N_10099,N_9831,N_9895);
xor U10100 (N_10100,N_9672,N_9741);
nor U10101 (N_10101,N_9784,N_9856);
nor U10102 (N_10102,N_9836,N_9677);
nand U10103 (N_10103,N_9737,N_9658);
or U10104 (N_10104,N_9899,N_9770);
xor U10105 (N_10105,N_9622,N_9869);
and U10106 (N_10106,N_9873,N_9766);
nor U10107 (N_10107,N_9858,N_9689);
nor U10108 (N_10108,N_9614,N_9859);
nor U10109 (N_10109,N_9822,N_9630);
nor U10110 (N_10110,N_9873,N_9783);
or U10111 (N_10111,N_9678,N_9735);
or U10112 (N_10112,N_9810,N_9833);
nor U10113 (N_10113,N_9730,N_9750);
xor U10114 (N_10114,N_9651,N_9743);
xnor U10115 (N_10115,N_9638,N_9603);
and U10116 (N_10116,N_9668,N_9869);
xnor U10117 (N_10117,N_9635,N_9885);
nand U10118 (N_10118,N_9789,N_9690);
nor U10119 (N_10119,N_9687,N_9720);
nand U10120 (N_10120,N_9633,N_9729);
and U10121 (N_10121,N_9737,N_9741);
xor U10122 (N_10122,N_9738,N_9813);
nand U10123 (N_10123,N_9822,N_9614);
and U10124 (N_10124,N_9827,N_9619);
and U10125 (N_10125,N_9659,N_9882);
xnor U10126 (N_10126,N_9765,N_9812);
nand U10127 (N_10127,N_9734,N_9666);
nor U10128 (N_10128,N_9731,N_9698);
or U10129 (N_10129,N_9660,N_9717);
nand U10130 (N_10130,N_9645,N_9805);
xor U10131 (N_10131,N_9668,N_9744);
and U10132 (N_10132,N_9782,N_9739);
or U10133 (N_10133,N_9812,N_9734);
nand U10134 (N_10134,N_9637,N_9621);
or U10135 (N_10135,N_9758,N_9745);
or U10136 (N_10136,N_9658,N_9612);
nand U10137 (N_10137,N_9781,N_9793);
and U10138 (N_10138,N_9637,N_9773);
and U10139 (N_10139,N_9898,N_9767);
nand U10140 (N_10140,N_9720,N_9698);
or U10141 (N_10141,N_9678,N_9629);
xor U10142 (N_10142,N_9864,N_9826);
and U10143 (N_10143,N_9856,N_9652);
and U10144 (N_10144,N_9655,N_9696);
xnor U10145 (N_10145,N_9744,N_9754);
or U10146 (N_10146,N_9679,N_9759);
and U10147 (N_10147,N_9730,N_9717);
nand U10148 (N_10148,N_9619,N_9894);
nand U10149 (N_10149,N_9778,N_9662);
or U10150 (N_10150,N_9730,N_9662);
nand U10151 (N_10151,N_9676,N_9724);
nand U10152 (N_10152,N_9767,N_9697);
xor U10153 (N_10153,N_9803,N_9793);
and U10154 (N_10154,N_9699,N_9876);
or U10155 (N_10155,N_9799,N_9618);
xor U10156 (N_10156,N_9819,N_9681);
and U10157 (N_10157,N_9857,N_9874);
and U10158 (N_10158,N_9743,N_9726);
and U10159 (N_10159,N_9655,N_9703);
nand U10160 (N_10160,N_9618,N_9635);
or U10161 (N_10161,N_9878,N_9845);
nor U10162 (N_10162,N_9792,N_9668);
nand U10163 (N_10163,N_9754,N_9644);
nor U10164 (N_10164,N_9699,N_9848);
nor U10165 (N_10165,N_9637,N_9742);
or U10166 (N_10166,N_9798,N_9827);
xnor U10167 (N_10167,N_9640,N_9769);
and U10168 (N_10168,N_9760,N_9670);
and U10169 (N_10169,N_9700,N_9765);
and U10170 (N_10170,N_9724,N_9675);
or U10171 (N_10171,N_9631,N_9866);
xnor U10172 (N_10172,N_9859,N_9637);
and U10173 (N_10173,N_9836,N_9600);
or U10174 (N_10174,N_9895,N_9635);
nand U10175 (N_10175,N_9696,N_9782);
nand U10176 (N_10176,N_9725,N_9777);
nor U10177 (N_10177,N_9892,N_9651);
nand U10178 (N_10178,N_9776,N_9817);
nor U10179 (N_10179,N_9651,N_9628);
or U10180 (N_10180,N_9755,N_9672);
xnor U10181 (N_10181,N_9695,N_9858);
nor U10182 (N_10182,N_9746,N_9651);
nor U10183 (N_10183,N_9707,N_9651);
nand U10184 (N_10184,N_9713,N_9661);
and U10185 (N_10185,N_9733,N_9784);
xor U10186 (N_10186,N_9868,N_9890);
xor U10187 (N_10187,N_9750,N_9663);
nor U10188 (N_10188,N_9618,N_9837);
or U10189 (N_10189,N_9877,N_9785);
or U10190 (N_10190,N_9718,N_9842);
xor U10191 (N_10191,N_9783,N_9632);
xor U10192 (N_10192,N_9800,N_9639);
or U10193 (N_10193,N_9683,N_9623);
or U10194 (N_10194,N_9819,N_9703);
and U10195 (N_10195,N_9775,N_9621);
nor U10196 (N_10196,N_9755,N_9730);
xor U10197 (N_10197,N_9742,N_9789);
xor U10198 (N_10198,N_9690,N_9797);
xnor U10199 (N_10199,N_9709,N_9615);
and U10200 (N_10200,N_10154,N_10020);
nand U10201 (N_10201,N_10142,N_10104);
nor U10202 (N_10202,N_9948,N_10110);
and U10203 (N_10203,N_10064,N_10146);
nor U10204 (N_10204,N_9944,N_10148);
nor U10205 (N_10205,N_10084,N_10103);
nand U10206 (N_10206,N_10065,N_9985);
or U10207 (N_10207,N_9953,N_10163);
nor U10208 (N_10208,N_10074,N_10185);
nand U10209 (N_10209,N_10151,N_10112);
or U10210 (N_10210,N_9901,N_10013);
or U10211 (N_10211,N_9938,N_10097);
or U10212 (N_10212,N_9980,N_9950);
and U10213 (N_10213,N_9979,N_9919);
xnor U10214 (N_10214,N_9930,N_10001);
and U10215 (N_10215,N_10149,N_9968);
xor U10216 (N_10216,N_10088,N_10028);
or U10217 (N_10217,N_10113,N_9957);
nor U10218 (N_10218,N_10130,N_10127);
nand U10219 (N_10219,N_10161,N_10137);
and U10220 (N_10220,N_9940,N_9971);
nand U10221 (N_10221,N_9970,N_10165);
or U10222 (N_10222,N_10176,N_10026);
xor U10223 (N_10223,N_9990,N_10140);
nor U10224 (N_10224,N_10045,N_10136);
and U10225 (N_10225,N_10105,N_10187);
or U10226 (N_10226,N_10119,N_10059);
nor U10227 (N_10227,N_9956,N_10016);
xor U10228 (N_10228,N_10082,N_10094);
nor U10229 (N_10229,N_10174,N_9952);
and U10230 (N_10230,N_9947,N_10175);
xnor U10231 (N_10231,N_10156,N_9965);
nand U10232 (N_10232,N_10051,N_9914);
nand U10233 (N_10233,N_9967,N_10124);
nand U10234 (N_10234,N_10086,N_10170);
nor U10235 (N_10235,N_9935,N_10005);
and U10236 (N_10236,N_10193,N_9933);
and U10237 (N_10237,N_10181,N_10116);
xor U10238 (N_10238,N_10197,N_9966);
and U10239 (N_10239,N_10056,N_10095);
nor U10240 (N_10240,N_10004,N_9912);
nor U10241 (N_10241,N_9991,N_9988);
nor U10242 (N_10242,N_10077,N_10031);
xnor U10243 (N_10243,N_9923,N_9982);
nand U10244 (N_10244,N_10007,N_9928);
xor U10245 (N_10245,N_10164,N_9993);
and U10246 (N_10246,N_10192,N_10035);
and U10247 (N_10247,N_10123,N_10171);
or U10248 (N_10248,N_9904,N_9902);
nor U10249 (N_10249,N_9961,N_10017);
or U10250 (N_10250,N_10108,N_10180);
and U10251 (N_10251,N_10195,N_9984);
nor U10252 (N_10252,N_10043,N_10138);
xor U10253 (N_10253,N_10050,N_9976);
nor U10254 (N_10254,N_10129,N_10060);
nor U10255 (N_10255,N_10145,N_9945);
and U10256 (N_10256,N_10033,N_9921);
nor U10257 (N_10257,N_10141,N_9954);
and U10258 (N_10258,N_10184,N_10081);
nor U10259 (N_10259,N_9908,N_9931);
nand U10260 (N_10260,N_10040,N_10090);
xnor U10261 (N_10261,N_10032,N_10076);
nor U10262 (N_10262,N_10179,N_10134);
nand U10263 (N_10263,N_10055,N_10014);
and U10264 (N_10264,N_10049,N_10018);
xnor U10265 (N_10265,N_10096,N_10121);
nand U10266 (N_10266,N_10169,N_10027);
nor U10267 (N_10267,N_9946,N_10071);
or U10268 (N_10268,N_10011,N_10101);
nor U10269 (N_10269,N_10102,N_9918);
or U10270 (N_10270,N_10126,N_10075);
nor U10271 (N_10271,N_9973,N_9911);
nand U10272 (N_10272,N_10162,N_10067);
and U10273 (N_10273,N_10186,N_10003);
or U10274 (N_10274,N_10167,N_10015);
or U10275 (N_10275,N_10131,N_9998);
and U10276 (N_10276,N_10109,N_10012);
and U10277 (N_10277,N_9958,N_9920);
nand U10278 (N_10278,N_9924,N_9964);
xnor U10279 (N_10279,N_10029,N_10182);
nor U10280 (N_10280,N_10139,N_10155);
nand U10281 (N_10281,N_9977,N_9989);
nor U10282 (N_10282,N_10062,N_9959);
nor U10283 (N_10283,N_10052,N_10099);
nand U10284 (N_10284,N_9929,N_10010);
and U10285 (N_10285,N_10189,N_10147);
nand U10286 (N_10286,N_10019,N_10114);
xor U10287 (N_10287,N_10006,N_9974);
nor U10288 (N_10288,N_10191,N_10152);
or U10289 (N_10289,N_9969,N_9934);
nor U10290 (N_10290,N_10039,N_9906);
xor U10291 (N_10291,N_10117,N_9915);
and U10292 (N_10292,N_10072,N_9926);
nor U10293 (N_10293,N_10150,N_9986);
nand U10294 (N_10294,N_9905,N_10022);
nor U10295 (N_10295,N_9900,N_10034);
xor U10296 (N_10296,N_10091,N_9999);
nor U10297 (N_10297,N_9925,N_10070);
nor U10298 (N_10298,N_10115,N_10128);
xnor U10299 (N_10299,N_10118,N_10196);
or U10300 (N_10300,N_10135,N_10068);
nor U10301 (N_10301,N_10009,N_10038);
xnor U10302 (N_10302,N_10120,N_10044);
or U10303 (N_10303,N_9992,N_10073);
or U10304 (N_10304,N_10160,N_10093);
nor U10305 (N_10305,N_10002,N_10143);
nor U10306 (N_10306,N_10172,N_10063);
or U10307 (N_10307,N_9962,N_9907);
and U10308 (N_10308,N_9997,N_10085);
xor U10309 (N_10309,N_10080,N_9972);
or U10310 (N_10310,N_10106,N_9917);
and U10311 (N_10311,N_10157,N_10199);
or U10312 (N_10312,N_10153,N_10057);
and U10313 (N_10313,N_9936,N_9981);
or U10314 (N_10314,N_9951,N_10132);
nand U10315 (N_10315,N_9994,N_9913);
nor U10316 (N_10316,N_10061,N_10048);
or U10317 (N_10317,N_10083,N_10079);
xnor U10318 (N_10318,N_10078,N_10058);
xnor U10319 (N_10319,N_10036,N_10133);
or U10320 (N_10320,N_10025,N_10066);
nor U10321 (N_10321,N_9978,N_9903);
or U10322 (N_10322,N_9955,N_10030);
nand U10323 (N_10323,N_10168,N_10166);
nor U10324 (N_10324,N_10125,N_10144);
and U10325 (N_10325,N_9983,N_10178);
nor U10326 (N_10326,N_10177,N_9941);
and U10327 (N_10327,N_9942,N_10107);
or U10328 (N_10328,N_10111,N_9987);
nor U10329 (N_10329,N_9995,N_10188);
xor U10330 (N_10330,N_10000,N_10098);
xnor U10331 (N_10331,N_10087,N_9932);
or U10332 (N_10332,N_10092,N_10069);
and U10333 (N_10333,N_10190,N_10089);
xnor U10334 (N_10334,N_9975,N_9927);
xor U10335 (N_10335,N_10122,N_10159);
xnor U10336 (N_10336,N_9937,N_10100);
or U10337 (N_10337,N_10053,N_10173);
and U10338 (N_10338,N_9909,N_9996);
nor U10339 (N_10339,N_9949,N_10041);
or U10340 (N_10340,N_10046,N_10158);
xor U10341 (N_10341,N_9960,N_10194);
or U10342 (N_10342,N_10047,N_10198);
nand U10343 (N_10343,N_10037,N_9910);
or U10344 (N_10344,N_10008,N_9963);
and U10345 (N_10345,N_10021,N_9939);
nand U10346 (N_10346,N_10042,N_10024);
or U10347 (N_10347,N_9922,N_10023);
or U10348 (N_10348,N_10054,N_10183);
or U10349 (N_10349,N_9916,N_9943);
and U10350 (N_10350,N_10085,N_10095);
nor U10351 (N_10351,N_10007,N_10188);
xnor U10352 (N_10352,N_9965,N_10008);
nor U10353 (N_10353,N_10135,N_10150);
or U10354 (N_10354,N_10094,N_10199);
and U10355 (N_10355,N_10081,N_9926);
and U10356 (N_10356,N_10049,N_10166);
and U10357 (N_10357,N_10151,N_10170);
or U10358 (N_10358,N_10185,N_10059);
nor U10359 (N_10359,N_10151,N_10187);
or U10360 (N_10360,N_10066,N_9988);
and U10361 (N_10361,N_10173,N_10088);
and U10362 (N_10362,N_9921,N_10041);
and U10363 (N_10363,N_10129,N_10059);
xor U10364 (N_10364,N_9904,N_9913);
nand U10365 (N_10365,N_10162,N_10135);
nor U10366 (N_10366,N_10032,N_10010);
or U10367 (N_10367,N_10167,N_9926);
nand U10368 (N_10368,N_10087,N_10052);
or U10369 (N_10369,N_10159,N_10187);
and U10370 (N_10370,N_10041,N_10034);
and U10371 (N_10371,N_10077,N_10012);
and U10372 (N_10372,N_10194,N_10065);
xnor U10373 (N_10373,N_10037,N_9944);
xor U10374 (N_10374,N_10196,N_10141);
nand U10375 (N_10375,N_9919,N_10048);
and U10376 (N_10376,N_10148,N_10160);
nor U10377 (N_10377,N_9920,N_9937);
nor U10378 (N_10378,N_9939,N_9946);
or U10379 (N_10379,N_10035,N_10117);
xor U10380 (N_10380,N_10024,N_10160);
nor U10381 (N_10381,N_9943,N_9934);
xnor U10382 (N_10382,N_9985,N_10019);
or U10383 (N_10383,N_9921,N_10162);
or U10384 (N_10384,N_9947,N_10031);
xnor U10385 (N_10385,N_10081,N_9924);
nand U10386 (N_10386,N_10152,N_10098);
nand U10387 (N_10387,N_10058,N_10041);
or U10388 (N_10388,N_10056,N_10100);
or U10389 (N_10389,N_9954,N_10195);
xnor U10390 (N_10390,N_10182,N_9984);
and U10391 (N_10391,N_10174,N_10111);
and U10392 (N_10392,N_9932,N_10068);
or U10393 (N_10393,N_9952,N_10158);
and U10394 (N_10394,N_10157,N_9938);
and U10395 (N_10395,N_10117,N_10107);
nor U10396 (N_10396,N_10020,N_10194);
and U10397 (N_10397,N_9974,N_10130);
nor U10398 (N_10398,N_10117,N_10013);
or U10399 (N_10399,N_10091,N_9990);
and U10400 (N_10400,N_9970,N_9917);
nor U10401 (N_10401,N_9930,N_10165);
and U10402 (N_10402,N_9966,N_9903);
or U10403 (N_10403,N_10049,N_10185);
nor U10404 (N_10404,N_10181,N_10148);
or U10405 (N_10405,N_9990,N_10172);
xor U10406 (N_10406,N_10020,N_10123);
and U10407 (N_10407,N_10114,N_10194);
nor U10408 (N_10408,N_10172,N_9935);
xnor U10409 (N_10409,N_9979,N_10095);
nand U10410 (N_10410,N_9978,N_10197);
and U10411 (N_10411,N_10087,N_9995);
nand U10412 (N_10412,N_10182,N_10027);
or U10413 (N_10413,N_10170,N_10147);
or U10414 (N_10414,N_10036,N_10027);
or U10415 (N_10415,N_9927,N_10127);
or U10416 (N_10416,N_9970,N_10008);
and U10417 (N_10417,N_10047,N_9986);
nand U10418 (N_10418,N_10096,N_10060);
nor U10419 (N_10419,N_9962,N_10047);
xnor U10420 (N_10420,N_10062,N_9979);
or U10421 (N_10421,N_10067,N_10122);
and U10422 (N_10422,N_10069,N_10060);
or U10423 (N_10423,N_9954,N_10160);
xor U10424 (N_10424,N_10187,N_10077);
or U10425 (N_10425,N_10185,N_10168);
nand U10426 (N_10426,N_10124,N_9936);
xnor U10427 (N_10427,N_10197,N_10055);
xnor U10428 (N_10428,N_10070,N_10041);
or U10429 (N_10429,N_9919,N_10127);
and U10430 (N_10430,N_9995,N_10036);
or U10431 (N_10431,N_10120,N_9962);
and U10432 (N_10432,N_10193,N_10107);
or U10433 (N_10433,N_10061,N_9924);
xor U10434 (N_10434,N_9948,N_10112);
nor U10435 (N_10435,N_9969,N_10138);
or U10436 (N_10436,N_9948,N_10082);
xor U10437 (N_10437,N_10109,N_9942);
or U10438 (N_10438,N_9941,N_10027);
nand U10439 (N_10439,N_10031,N_10143);
or U10440 (N_10440,N_10115,N_10109);
nand U10441 (N_10441,N_10040,N_10116);
nor U10442 (N_10442,N_9960,N_10147);
nor U10443 (N_10443,N_10051,N_10149);
xnor U10444 (N_10444,N_10041,N_10028);
xnor U10445 (N_10445,N_10177,N_9907);
nor U10446 (N_10446,N_10143,N_10012);
and U10447 (N_10447,N_9904,N_10012);
or U10448 (N_10448,N_9941,N_10119);
xnor U10449 (N_10449,N_10126,N_10033);
or U10450 (N_10450,N_10142,N_10111);
and U10451 (N_10451,N_10189,N_9926);
nand U10452 (N_10452,N_10070,N_9970);
nor U10453 (N_10453,N_10108,N_10114);
and U10454 (N_10454,N_10136,N_10060);
or U10455 (N_10455,N_9949,N_10016);
xnor U10456 (N_10456,N_9940,N_10093);
nand U10457 (N_10457,N_10083,N_10130);
and U10458 (N_10458,N_9998,N_10138);
xor U10459 (N_10459,N_9970,N_10186);
nand U10460 (N_10460,N_10122,N_9906);
nand U10461 (N_10461,N_10111,N_9994);
or U10462 (N_10462,N_9943,N_10188);
or U10463 (N_10463,N_10108,N_9949);
and U10464 (N_10464,N_10155,N_9950);
and U10465 (N_10465,N_9998,N_10159);
nand U10466 (N_10466,N_9924,N_9995);
xor U10467 (N_10467,N_10123,N_9950);
or U10468 (N_10468,N_9975,N_10031);
or U10469 (N_10469,N_10074,N_10006);
nand U10470 (N_10470,N_9984,N_9942);
nand U10471 (N_10471,N_10029,N_10006);
and U10472 (N_10472,N_10105,N_10182);
xnor U10473 (N_10473,N_10116,N_10102);
and U10474 (N_10474,N_10154,N_9905);
and U10475 (N_10475,N_9921,N_10145);
nor U10476 (N_10476,N_10006,N_9997);
nor U10477 (N_10477,N_10093,N_10001);
or U10478 (N_10478,N_9920,N_9991);
nor U10479 (N_10479,N_9938,N_9957);
nor U10480 (N_10480,N_10140,N_9973);
xor U10481 (N_10481,N_9964,N_10018);
nand U10482 (N_10482,N_10149,N_9980);
xnor U10483 (N_10483,N_10046,N_10189);
nor U10484 (N_10484,N_10014,N_10088);
and U10485 (N_10485,N_10088,N_9960);
xor U10486 (N_10486,N_10121,N_10072);
or U10487 (N_10487,N_10069,N_9970);
nor U10488 (N_10488,N_10066,N_10057);
and U10489 (N_10489,N_10007,N_9976);
or U10490 (N_10490,N_10199,N_10017);
xor U10491 (N_10491,N_9906,N_10037);
xnor U10492 (N_10492,N_9903,N_9915);
or U10493 (N_10493,N_10166,N_10106);
nor U10494 (N_10494,N_10061,N_10042);
nor U10495 (N_10495,N_10022,N_9913);
and U10496 (N_10496,N_9960,N_9959);
nand U10497 (N_10497,N_9921,N_10067);
and U10498 (N_10498,N_10133,N_10181);
xor U10499 (N_10499,N_10151,N_10018);
or U10500 (N_10500,N_10393,N_10262);
nor U10501 (N_10501,N_10499,N_10396);
or U10502 (N_10502,N_10244,N_10338);
nand U10503 (N_10503,N_10240,N_10237);
nand U10504 (N_10504,N_10346,N_10308);
or U10505 (N_10505,N_10249,N_10284);
nand U10506 (N_10506,N_10459,N_10213);
or U10507 (N_10507,N_10397,N_10443);
nor U10508 (N_10508,N_10370,N_10353);
xor U10509 (N_10509,N_10405,N_10328);
nand U10510 (N_10510,N_10285,N_10255);
or U10511 (N_10511,N_10301,N_10371);
xnor U10512 (N_10512,N_10481,N_10463);
or U10513 (N_10513,N_10433,N_10462);
nand U10514 (N_10514,N_10254,N_10354);
nor U10515 (N_10515,N_10402,N_10283);
nor U10516 (N_10516,N_10485,N_10434);
nor U10517 (N_10517,N_10467,N_10343);
or U10518 (N_10518,N_10468,N_10281);
nand U10519 (N_10519,N_10436,N_10289);
nand U10520 (N_10520,N_10426,N_10300);
or U10521 (N_10521,N_10440,N_10329);
nor U10522 (N_10522,N_10486,N_10480);
or U10523 (N_10523,N_10239,N_10482);
and U10524 (N_10524,N_10216,N_10245);
nor U10525 (N_10525,N_10274,N_10364);
or U10526 (N_10526,N_10407,N_10327);
xor U10527 (N_10527,N_10309,N_10496);
or U10528 (N_10528,N_10305,N_10429);
nand U10529 (N_10529,N_10418,N_10363);
and U10530 (N_10530,N_10386,N_10493);
nand U10531 (N_10531,N_10413,N_10264);
nor U10532 (N_10532,N_10470,N_10401);
or U10533 (N_10533,N_10252,N_10372);
and U10534 (N_10534,N_10414,N_10207);
xnor U10535 (N_10535,N_10212,N_10415);
xnor U10536 (N_10536,N_10447,N_10204);
nand U10537 (N_10537,N_10474,N_10458);
nor U10538 (N_10538,N_10484,N_10417);
nand U10539 (N_10539,N_10427,N_10286);
or U10540 (N_10540,N_10491,N_10473);
nor U10541 (N_10541,N_10333,N_10208);
and U10542 (N_10542,N_10444,N_10241);
nor U10543 (N_10543,N_10307,N_10389);
xor U10544 (N_10544,N_10369,N_10258);
nor U10545 (N_10545,N_10478,N_10276);
and U10546 (N_10546,N_10288,N_10223);
or U10547 (N_10547,N_10411,N_10339);
nor U10548 (N_10548,N_10416,N_10391);
or U10549 (N_10549,N_10383,N_10382);
xor U10550 (N_10550,N_10206,N_10457);
xnor U10551 (N_10551,N_10430,N_10437);
xor U10552 (N_10552,N_10366,N_10290);
xnor U10553 (N_10553,N_10466,N_10282);
nand U10554 (N_10554,N_10228,N_10344);
xor U10555 (N_10555,N_10351,N_10326);
xor U10556 (N_10556,N_10266,N_10292);
xor U10557 (N_10557,N_10475,N_10464);
or U10558 (N_10558,N_10422,N_10250);
nor U10559 (N_10559,N_10247,N_10439);
or U10560 (N_10560,N_10201,N_10404);
xnor U10561 (N_10561,N_10242,N_10409);
nor U10562 (N_10562,N_10445,N_10441);
nand U10563 (N_10563,N_10345,N_10248);
nor U10564 (N_10564,N_10321,N_10337);
xnor U10565 (N_10565,N_10373,N_10267);
or U10566 (N_10566,N_10403,N_10296);
nor U10567 (N_10567,N_10279,N_10498);
or U10568 (N_10568,N_10243,N_10231);
xor U10569 (N_10569,N_10356,N_10320);
nand U10570 (N_10570,N_10280,N_10450);
nor U10571 (N_10571,N_10315,N_10492);
or U10572 (N_10572,N_10361,N_10472);
nand U10573 (N_10573,N_10358,N_10215);
or U10574 (N_10574,N_10375,N_10259);
nor U10575 (N_10575,N_10374,N_10420);
nand U10576 (N_10576,N_10214,N_10256);
nand U10577 (N_10577,N_10218,N_10360);
and U10578 (N_10578,N_10203,N_10224);
nand U10579 (N_10579,N_10298,N_10236);
nor U10580 (N_10580,N_10271,N_10350);
nand U10581 (N_10581,N_10477,N_10421);
xor U10582 (N_10582,N_10225,N_10385);
nor U10583 (N_10583,N_10387,N_10270);
xnor U10584 (N_10584,N_10340,N_10273);
nand U10585 (N_10585,N_10209,N_10419);
nand U10586 (N_10586,N_10332,N_10287);
and U10587 (N_10587,N_10390,N_10490);
nor U10588 (N_10588,N_10408,N_10448);
nand U10589 (N_10589,N_10451,N_10489);
or U10590 (N_10590,N_10494,N_10318);
nor U10591 (N_10591,N_10347,N_10362);
xnor U10592 (N_10592,N_10355,N_10342);
nor U10593 (N_10593,N_10455,N_10306);
nand U10594 (N_10594,N_10263,N_10211);
nand U10595 (N_10595,N_10428,N_10476);
or U10596 (N_10596,N_10469,N_10400);
and U10597 (N_10597,N_10221,N_10226);
nand U10598 (N_10598,N_10435,N_10222);
xnor U10599 (N_10599,N_10446,N_10323);
nand U10600 (N_10600,N_10299,N_10322);
xnor U10601 (N_10601,N_10379,N_10234);
xor U10602 (N_10602,N_10257,N_10495);
xnor U10603 (N_10603,N_10202,N_10265);
nor U10604 (N_10604,N_10330,N_10497);
nor U10605 (N_10605,N_10210,N_10291);
or U10606 (N_10606,N_10260,N_10406);
nor U10607 (N_10607,N_10479,N_10232);
nand U10608 (N_10608,N_10378,N_10335);
xnor U10609 (N_10609,N_10314,N_10410);
and U10610 (N_10610,N_10269,N_10423);
nor U10611 (N_10611,N_10357,N_10461);
and U10612 (N_10612,N_10376,N_10398);
and U10613 (N_10613,N_10293,N_10365);
nand U10614 (N_10614,N_10487,N_10384);
or U10615 (N_10615,N_10253,N_10238);
xor U10616 (N_10616,N_10304,N_10229);
xnor U10617 (N_10617,N_10460,N_10277);
and U10618 (N_10618,N_10275,N_10454);
nand U10619 (N_10619,N_10431,N_10261);
nor U10620 (N_10620,N_10456,N_10392);
or U10621 (N_10621,N_10325,N_10368);
xnor U10622 (N_10622,N_10294,N_10453);
and U10623 (N_10623,N_10311,N_10395);
and U10624 (N_10624,N_10488,N_10295);
or U10625 (N_10625,N_10278,N_10432);
xnor U10626 (N_10626,N_10452,N_10465);
xor U10627 (N_10627,N_10230,N_10425);
xnor U10628 (N_10628,N_10367,N_10272);
or U10629 (N_10629,N_10303,N_10377);
or U10630 (N_10630,N_10227,N_10297);
nand U10631 (N_10631,N_10233,N_10341);
nor U10632 (N_10632,N_10235,N_10246);
or U10633 (N_10633,N_10217,N_10310);
nand U10634 (N_10634,N_10302,N_10394);
xor U10635 (N_10635,N_10331,N_10359);
xor U10636 (N_10636,N_10334,N_10349);
xnor U10637 (N_10637,N_10336,N_10442);
xnor U10638 (N_10638,N_10205,N_10319);
nor U10639 (N_10639,N_10348,N_10324);
and U10640 (N_10640,N_10399,N_10219);
nand U10641 (N_10641,N_10380,N_10449);
and U10642 (N_10642,N_10381,N_10313);
nor U10643 (N_10643,N_10352,N_10412);
or U10644 (N_10644,N_10424,N_10268);
nor U10645 (N_10645,N_10317,N_10251);
xor U10646 (N_10646,N_10438,N_10200);
or U10647 (N_10647,N_10312,N_10483);
nand U10648 (N_10648,N_10471,N_10220);
or U10649 (N_10649,N_10388,N_10316);
nand U10650 (N_10650,N_10361,N_10282);
nand U10651 (N_10651,N_10276,N_10311);
nand U10652 (N_10652,N_10264,N_10306);
xnor U10653 (N_10653,N_10274,N_10341);
nor U10654 (N_10654,N_10434,N_10442);
nand U10655 (N_10655,N_10291,N_10275);
or U10656 (N_10656,N_10352,N_10200);
nand U10657 (N_10657,N_10460,N_10429);
nor U10658 (N_10658,N_10444,N_10276);
xnor U10659 (N_10659,N_10284,N_10248);
nor U10660 (N_10660,N_10390,N_10303);
nand U10661 (N_10661,N_10281,N_10435);
and U10662 (N_10662,N_10446,N_10245);
nor U10663 (N_10663,N_10354,N_10255);
and U10664 (N_10664,N_10345,N_10276);
nand U10665 (N_10665,N_10485,N_10222);
nor U10666 (N_10666,N_10300,N_10369);
xor U10667 (N_10667,N_10441,N_10284);
and U10668 (N_10668,N_10385,N_10458);
nand U10669 (N_10669,N_10365,N_10360);
xor U10670 (N_10670,N_10250,N_10316);
nand U10671 (N_10671,N_10447,N_10296);
xnor U10672 (N_10672,N_10311,N_10388);
and U10673 (N_10673,N_10433,N_10367);
or U10674 (N_10674,N_10257,N_10497);
xor U10675 (N_10675,N_10210,N_10399);
nand U10676 (N_10676,N_10401,N_10255);
nand U10677 (N_10677,N_10215,N_10362);
and U10678 (N_10678,N_10306,N_10332);
nand U10679 (N_10679,N_10479,N_10215);
xor U10680 (N_10680,N_10255,N_10470);
or U10681 (N_10681,N_10480,N_10381);
and U10682 (N_10682,N_10411,N_10456);
nor U10683 (N_10683,N_10470,N_10318);
xnor U10684 (N_10684,N_10396,N_10477);
nor U10685 (N_10685,N_10271,N_10459);
and U10686 (N_10686,N_10238,N_10381);
and U10687 (N_10687,N_10257,N_10354);
xor U10688 (N_10688,N_10342,N_10260);
and U10689 (N_10689,N_10324,N_10250);
or U10690 (N_10690,N_10243,N_10387);
nor U10691 (N_10691,N_10341,N_10259);
xor U10692 (N_10692,N_10306,N_10441);
and U10693 (N_10693,N_10372,N_10358);
nand U10694 (N_10694,N_10316,N_10335);
nor U10695 (N_10695,N_10348,N_10386);
or U10696 (N_10696,N_10421,N_10431);
nor U10697 (N_10697,N_10263,N_10322);
or U10698 (N_10698,N_10448,N_10411);
nand U10699 (N_10699,N_10479,N_10368);
xnor U10700 (N_10700,N_10408,N_10372);
and U10701 (N_10701,N_10224,N_10216);
nand U10702 (N_10702,N_10223,N_10266);
and U10703 (N_10703,N_10486,N_10256);
or U10704 (N_10704,N_10300,N_10317);
nand U10705 (N_10705,N_10499,N_10425);
xnor U10706 (N_10706,N_10390,N_10386);
xnor U10707 (N_10707,N_10494,N_10371);
and U10708 (N_10708,N_10381,N_10252);
or U10709 (N_10709,N_10439,N_10245);
nand U10710 (N_10710,N_10255,N_10389);
nor U10711 (N_10711,N_10262,N_10288);
xor U10712 (N_10712,N_10405,N_10287);
or U10713 (N_10713,N_10270,N_10302);
nor U10714 (N_10714,N_10494,N_10277);
xnor U10715 (N_10715,N_10248,N_10312);
and U10716 (N_10716,N_10255,N_10393);
xor U10717 (N_10717,N_10366,N_10226);
nand U10718 (N_10718,N_10358,N_10416);
xnor U10719 (N_10719,N_10476,N_10239);
nor U10720 (N_10720,N_10421,N_10405);
xor U10721 (N_10721,N_10228,N_10436);
xor U10722 (N_10722,N_10335,N_10416);
or U10723 (N_10723,N_10280,N_10268);
or U10724 (N_10724,N_10364,N_10213);
xor U10725 (N_10725,N_10223,N_10331);
nand U10726 (N_10726,N_10459,N_10240);
or U10727 (N_10727,N_10224,N_10271);
and U10728 (N_10728,N_10348,N_10457);
nor U10729 (N_10729,N_10395,N_10296);
or U10730 (N_10730,N_10411,N_10419);
xnor U10731 (N_10731,N_10385,N_10368);
or U10732 (N_10732,N_10485,N_10318);
or U10733 (N_10733,N_10408,N_10273);
xnor U10734 (N_10734,N_10356,N_10215);
or U10735 (N_10735,N_10420,N_10412);
xor U10736 (N_10736,N_10266,N_10293);
and U10737 (N_10737,N_10445,N_10336);
nor U10738 (N_10738,N_10490,N_10474);
nand U10739 (N_10739,N_10275,N_10403);
or U10740 (N_10740,N_10249,N_10245);
nand U10741 (N_10741,N_10363,N_10467);
nor U10742 (N_10742,N_10445,N_10313);
or U10743 (N_10743,N_10445,N_10478);
nand U10744 (N_10744,N_10408,N_10462);
or U10745 (N_10745,N_10354,N_10280);
xnor U10746 (N_10746,N_10263,N_10452);
or U10747 (N_10747,N_10376,N_10382);
or U10748 (N_10748,N_10208,N_10327);
nor U10749 (N_10749,N_10343,N_10423);
and U10750 (N_10750,N_10480,N_10459);
and U10751 (N_10751,N_10388,N_10486);
nor U10752 (N_10752,N_10316,N_10487);
nor U10753 (N_10753,N_10398,N_10247);
and U10754 (N_10754,N_10397,N_10309);
nand U10755 (N_10755,N_10354,N_10430);
xor U10756 (N_10756,N_10354,N_10328);
nor U10757 (N_10757,N_10305,N_10203);
or U10758 (N_10758,N_10357,N_10314);
and U10759 (N_10759,N_10384,N_10294);
xnor U10760 (N_10760,N_10232,N_10259);
nand U10761 (N_10761,N_10498,N_10251);
or U10762 (N_10762,N_10239,N_10481);
or U10763 (N_10763,N_10431,N_10308);
nor U10764 (N_10764,N_10294,N_10457);
and U10765 (N_10765,N_10307,N_10415);
or U10766 (N_10766,N_10406,N_10369);
or U10767 (N_10767,N_10321,N_10450);
or U10768 (N_10768,N_10462,N_10444);
or U10769 (N_10769,N_10470,N_10420);
or U10770 (N_10770,N_10475,N_10335);
and U10771 (N_10771,N_10318,N_10211);
or U10772 (N_10772,N_10486,N_10317);
xor U10773 (N_10773,N_10232,N_10271);
nand U10774 (N_10774,N_10289,N_10452);
or U10775 (N_10775,N_10477,N_10320);
nor U10776 (N_10776,N_10242,N_10222);
nor U10777 (N_10777,N_10390,N_10424);
and U10778 (N_10778,N_10456,N_10426);
nor U10779 (N_10779,N_10330,N_10291);
xor U10780 (N_10780,N_10389,N_10454);
nor U10781 (N_10781,N_10317,N_10432);
or U10782 (N_10782,N_10493,N_10400);
nor U10783 (N_10783,N_10290,N_10394);
nor U10784 (N_10784,N_10276,N_10474);
nand U10785 (N_10785,N_10305,N_10254);
nor U10786 (N_10786,N_10449,N_10492);
or U10787 (N_10787,N_10389,N_10487);
nor U10788 (N_10788,N_10223,N_10415);
nand U10789 (N_10789,N_10407,N_10479);
and U10790 (N_10790,N_10416,N_10301);
or U10791 (N_10791,N_10387,N_10424);
nor U10792 (N_10792,N_10369,N_10403);
or U10793 (N_10793,N_10213,N_10405);
nor U10794 (N_10794,N_10410,N_10307);
xor U10795 (N_10795,N_10281,N_10396);
xor U10796 (N_10796,N_10395,N_10378);
nand U10797 (N_10797,N_10478,N_10332);
xnor U10798 (N_10798,N_10327,N_10436);
and U10799 (N_10799,N_10200,N_10356);
and U10800 (N_10800,N_10709,N_10586);
or U10801 (N_10801,N_10769,N_10549);
or U10802 (N_10802,N_10619,N_10640);
xor U10803 (N_10803,N_10780,N_10734);
nand U10804 (N_10804,N_10599,N_10721);
or U10805 (N_10805,N_10545,N_10691);
nand U10806 (N_10806,N_10704,N_10714);
and U10807 (N_10807,N_10560,N_10661);
xor U10808 (N_10808,N_10713,N_10783);
or U10809 (N_10809,N_10637,N_10509);
or U10810 (N_10810,N_10767,N_10508);
xor U10811 (N_10811,N_10676,N_10500);
nand U10812 (N_10812,N_10528,N_10542);
nand U10813 (N_10813,N_10700,N_10649);
or U10814 (N_10814,N_10644,N_10642);
and U10815 (N_10815,N_10554,N_10611);
nand U10816 (N_10816,N_10543,N_10752);
or U10817 (N_10817,N_10510,N_10565);
xnor U10818 (N_10818,N_10635,N_10712);
or U10819 (N_10819,N_10658,N_10774);
nand U10820 (N_10820,N_10773,N_10553);
xnor U10821 (N_10821,N_10681,N_10502);
or U10822 (N_10822,N_10732,N_10777);
nand U10823 (N_10823,N_10756,N_10630);
xor U10824 (N_10824,N_10778,N_10701);
xnor U10825 (N_10825,N_10536,N_10548);
nand U10826 (N_10826,N_10601,N_10561);
or U10827 (N_10827,N_10753,N_10538);
nor U10828 (N_10828,N_10740,N_10585);
and U10829 (N_10829,N_10574,N_10795);
xor U10830 (N_10830,N_10657,N_10575);
nand U10831 (N_10831,N_10641,N_10720);
xnor U10832 (N_10832,N_10763,N_10648);
nand U10833 (N_10833,N_10787,N_10547);
xnor U10834 (N_10834,N_10782,N_10789);
and U10835 (N_10835,N_10512,N_10504);
and U10836 (N_10836,N_10555,N_10647);
or U10837 (N_10837,N_10743,N_10730);
and U10838 (N_10838,N_10604,N_10583);
or U10839 (N_10839,N_10516,N_10715);
or U10840 (N_10840,N_10632,N_10692);
nand U10841 (N_10841,N_10653,N_10564);
and U10842 (N_10842,N_10551,N_10592);
nor U10843 (N_10843,N_10639,N_10530);
or U10844 (N_10844,N_10505,N_10615);
xnor U10845 (N_10845,N_10742,N_10697);
nor U10846 (N_10846,N_10638,N_10607);
or U10847 (N_10847,N_10750,N_10762);
nor U10848 (N_10848,N_10798,N_10673);
nand U10849 (N_10849,N_10520,N_10797);
xor U10850 (N_10850,N_10580,N_10758);
or U10851 (N_10851,N_10522,N_10771);
nor U10852 (N_10852,N_10534,N_10723);
nor U10853 (N_10853,N_10693,N_10682);
nand U10854 (N_10854,N_10563,N_10550);
nand U10855 (N_10855,N_10728,N_10727);
and U10856 (N_10856,N_10594,N_10775);
xor U10857 (N_10857,N_10633,N_10610);
nand U10858 (N_10858,N_10518,N_10786);
and U10859 (N_10859,N_10790,N_10757);
or U10860 (N_10860,N_10539,N_10659);
and U10861 (N_10861,N_10595,N_10687);
nand U10862 (N_10862,N_10625,N_10537);
or U10863 (N_10863,N_10627,N_10646);
nor U10864 (N_10864,N_10710,N_10770);
and U10865 (N_10865,N_10568,N_10576);
xor U10866 (N_10866,N_10589,N_10624);
nand U10867 (N_10867,N_10572,N_10737);
nor U10868 (N_10868,N_10702,N_10579);
and U10869 (N_10869,N_10501,N_10540);
or U10870 (N_10870,N_10722,N_10747);
nor U10871 (N_10871,N_10717,N_10794);
and U10872 (N_10872,N_10552,N_10707);
nand U10873 (N_10873,N_10581,N_10695);
nand U10874 (N_10874,N_10684,N_10598);
or U10875 (N_10875,N_10514,N_10706);
and U10876 (N_10876,N_10655,N_10622);
nand U10877 (N_10877,N_10577,N_10716);
nor U10878 (N_10878,N_10525,N_10760);
or U10879 (N_10879,N_10678,N_10602);
nor U10880 (N_10880,N_10652,N_10672);
xor U10881 (N_10881,N_10733,N_10650);
nand U10882 (N_10882,N_10524,N_10685);
nor U10883 (N_10883,N_10614,N_10683);
and U10884 (N_10884,N_10527,N_10541);
or U10885 (N_10885,N_10664,N_10507);
and U10886 (N_10886,N_10779,N_10784);
or U10887 (N_10887,N_10671,N_10620);
and U10888 (N_10888,N_10725,N_10674);
nand U10889 (N_10889,N_10590,N_10670);
xor U10890 (N_10890,N_10596,N_10544);
and U10891 (N_10891,N_10517,N_10739);
or U10892 (N_10892,N_10677,N_10591);
and U10893 (N_10893,N_10593,N_10785);
or U10894 (N_10894,N_10588,N_10751);
nand U10895 (N_10895,N_10662,N_10791);
xor U10896 (N_10896,N_10645,N_10711);
nor U10897 (N_10897,N_10506,N_10689);
xor U10898 (N_10898,N_10634,N_10562);
and U10899 (N_10899,N_10666,N_10643);
nor U10900 (N_10900,N_10754,N_10718);
and U10901 (N_10901,N_10533,N_10587);
xor U10902 (N_10902,N_10513,N_10799);
or U10903 (N_10903,N_10667,N_10546);
or U10904 (N_10904,N_10665,N_10705);
xor U10905 (N_10905,N_10621,N_10663);
and U10906 (N_10906,N_10567,N_10738);
nand U10907 (N_10907,N_10571,N_10557);
nand U10908 (N_10908,N_10680,N_10613);
and U10909 (N_10909,N_10793,N_10746);
xor U10910 (N_10910,N_10675,N_10526);
and U10911 (N_10911,N_10612,N_10556);
nor U10912 (N_10912,N_10729,N_10569);
nand U10913 (N_10913,N_10566,N_10616);
and U10914 (N_10914,N_10690,N_10660);
and U10915 (N_10915,N_10759,N_10741);
or U10916 (N_10916,N_10605,N_10656);
xnor U10917 (N_10917,N_10558,N_10606);
nand U10918 (N_10918,N_10573,N_10523);
xor U10919 (N_10919,N_10511,N_10519);
nand U10920 (N_10920,N_10531,N_10559);
xnor U10921 (N_10921,N_10532,N_10629);
nor U10922 (N_10922,N_10608,N_10651);
and U10923 (N_10923,N_10669,N_10582);
xor U10924 (N_10924,N_10600,N_10766);
or U10925 (N_10925,N_10529,N_10626);
nor U10926 (N_10926,N_10748,N_10584);
xor U10927 (N_10927,N_10696,N_10628);
xnor U10928 (N_10928,N_10761,N_10631);
or U10929 (N_10929,N_10668,N_10578);
and U10930 (N_10930,N_10736,N_10617);
nand U10931 (N_10931,N_10788,N_10654);
nand U10932 (N_10932,N_10535,N_10724);
and U10933 (N_10933,N_10686,N_10623);
nor U10934 (N_10934,N_10749,N_10688);
or U10935 (N_10935,N_10521,N_10776);
and U10936 (N_10936,N_10744,N_10679);
nand U10937 (N_10937,N_10597,N_10694);
nand U10938 (N_10938,N_10731,N_10609);
or U10939 (N_10939,N_10796,N_10603);
nor U10940 (N_10940,N_10636,N_10726);
and U10941 (N_10941,N_10735,N_10503);
xor U10942 (N_10942,N_10745,N_10515);
or U10943 (N_10943,N_10570,N_10768);
and U10944 (N_10944,N_10781,N_10755);
xor U10945 (N_10945,N_10698,N_10792);
and U10946 (N_10946,N_10772,N_10699);
and U10947 (N_10947,N_10618,N_10765);
or U10948 (N_10948,N_10708,N_10703);
and U10949 (N_10949,N_10764,N_10719);
and U10950 (N_10950,N_10530,N_10697);
xor U10951 (N_10951,N_10604,N_10590);
xnor U10952 (N_10952,N_10762,N_10720);
xor U10953 (N_10953,N_10776,N_10782);
or U10954 (N_10954,N_10787,N_10662);
nand U10955 (N_10955,N_10623,N_10531);
xor U10956 (N_10956,N_10638,N_10640);
nand U10957 (N_10957,N_10642,N_10796);
and U10958 (N_10958,N_10562,N_10556);
nor U10959 (N_10959,N_10550,N_10580);
or U10960 (N_10960,N_10537,N_10536);
nor U10961 (N_10961,N_10530,N_10573);
or U10962 (N_10962,N_10579,N_10605);
or U10963 (N_10963,N_10709,N_10636);
xnor U10964 (N_10964,N_10775,N_10602);
xnor U10965 (N_10965,N_10515,N_10507);
nor U10966 (N_10966,N_10721,N_10546);
xor U10967 (N_10967,N_10553,N_10734);
or U10968 (N_10968,N_10574,N_10643);
and U10969 (N_10969,N_10728,N_10714);
and U10970 (N_10970,N_10601,N_10757);
or U10971 (N_10971,N_10520,N_10700);
and U10972 (N_10972,N_10717,N_10560);
nor U10973 (N_10973,N_10687,N_10579);
nor U10974 (N_10974,N_10545,N_10788);
and U10975 (N_10975,N_10725,N_10710);
and U10976 (N_10976,N_10759,N_10786);
and U10977 (N_10977,N_10766,N_10570);
or U10978 (N_10978,N_10574,N_10763);
xor U10979 (N_10979,N_10640,N_10613);
nand U10980 (N_10980,N_10726,N_10590);
and U10981 (N_10981,N_10767,N_10504);
or U10982 (N_10982,N_10529,N_10722);
nand U10983 (N_10983,N_10669,N_10704);
nand U10984 (N_10984,N_10536,N_10720);
or U10985 (N_10985,N_10634,N_10794);
nor U10986 (N_10986,N_10799,N_10666);
nor U10987 (N_10987,N_10529,N_10750);
nand U10988 (N_10988,N_10748,N_10696);
nand U10989 (N_10989,N_10510,N_10521);
or U10990 (N_10990,N_10705,N_10546);
nand U10991 (N_10991,N_10671,N_10512);
xor U10992 (N_10992,N_10663,N_10660);
nand U10993 (N_10993,N_10594,N_10549);
nor U10994 (N_10994,N_10775,N_10794);
xnor U10995 (N_10995,N_10610,N_10590);
nor U10996 (N_10996,N_10548,N_10557);
xnor U10997 (N_10997,N_10692,N_10528);
nor U10998 (N_10998,N_10582,N_10616);
and U10999 (N_10999,N_10516,N_10583);
nand U11000 (N_11000,N_10776,N_10740);
nor U11001 (N_11001,N_10555,N_10546);
xnor U11002 (N_11002,N_10641,N_10631);
nor U11003 (N_11003,N_10733,N_10726);
nor U11004 (N_11004,N_10595,N_10501);
nand U11005 (N_11005,N_10646,N_10503);
xnor U11006 (N_11006,N_10676,N_10518);
xor U11007 (N_11007,N_10669,N_10628);
nand U11008 (N_11008,N_10672,N_10761);
or U11009 (N_11009,N_10757,N_10719);
xor U11010 (N_11010,N_10726,N_10763);
xor U11011 (N_11011,N_10657,N_10757);
nand U11012 (N_11012,N_10642,N_10578);
and U11013 (N_11013,N_10646,N_10500);
and U11014 (N_11014,N_10527,N_10757);
and U11015 (N_11015,N_10661,N_10598);
and U11016 (N_11016,N_10778,N_10616);
nand U11017 (N_11017,N_10618,N_10592);
or U11018 (N_11018,N_10730,N_10685);
or U11019 (N_11019,N_10738,N_10704);
or U11020 (N_11020,N_10520,N_10667);
and U11021 (N_11021,N_10704,N_10640);
or U11022 (N_11022,N_10600,N_10585);
or U11023 (N_11023,N_10795,N_10684);
or U11024 (N_11024,N_10705,N_10603);
nand U11025 (N_11025,N_10764,N_10608);
or U11026 (N_11026,N_10525,N_10722);
xor U11027 (N_11027,N_10685,N_10643);
and U11028 (N_11028,N_10695,N_10508);
xor U11029 (N_11029,N_10506,N_10738);
or U11030 (N_11030,N_10616,N_10764);
or U11031 (N_11031,N_10633,N_10736);
and U11032 (N_11032,N_10729,N_10741);
or U11033 (N_11033,N_10695,N_10596);
or U11034 (N_11034,N_10527,N_10730);
xor U11035 (N_11035,N_10736,N_10503);
xnor U11036 (N_11036,N_10608,N_10679);
nand U11037 (N_11037,N_10786,N_10791);
nand U11038 (N_11038,N_10712,N_10748);
or U11039 (N_11039,N_10606,N_10695);
xnor U11040 (N_11040,N_10725,N_10650);
or U11041 (N_11041,N_10797,N_10608);
xor U11042 (N_11042,N_10715,N_10770);
xnor U11043 (N_11043,N_10785,N_10523);
nand U11044 (N_11044,N_10676,N_10768);
nand U11045 (N_11045,N_10623,N_10657);
xor U11046 (N_11046,N_10660,N_10528);
and U11047 (N_11047,N_10668,N_10728);
or U11048 (N_11048,N_10649,N_10568);
xor U11049 (N_11049,N_10728,N_10627);
or U11050 (N_11050,N_10637,N_10679);
and U11051 (N_11051,N_10777,N_10755);
and U11052 (N_11052,N_10733,N_10768);
and U11053 (N_11053,N_10672,N_10595);
nand U11054 (N_11054,N_10666,N_10554);
nand U11055 (N_11055,N_10578,N_10639);
or U11056 (N_11056,N_10675,N_10741);
nand U11057 (N_11057,N_10539,N_10731);
xnor U11058 (N_11058,N_10557,N_10758);
nor U11059 (N_11059,N_10576,N_10782);
and U11060 (N_11060,N_10749,N_10689);
nand U11061 (N_11061,N_10668,N_10607);
nor U11062 (N_11062,N_10697,N_10582);
and U11063 (N_11063,N_10534,N_10548);
xor U11064 (N_11064,N_10758,N_10790);
and U11065 (N_11065,N_10525,N_10748);
nand U11066 (N_11066,N_10737,N_10670);
nor U11067 (N_11067,N_10540,N_10577);
nand U11068 (N_11068,N_10537,N_10591);
nand U11069 (N_11069,N_10690,N_10758);
or U11070 (N_11070,N_10547,N_10641);
and U11071 (N_11071,N_10725,N_10724);
xor U11072 (N_11072,N_10748,N_10608);
or U11073 (N_11073,N_10528,N_10597);
and U11074 (N_11074,N_10677,N_10588);
or U11075 (N_11075,N_10571,N_10696);
xnor U11076 (N_11076,N_10580,N_10703);
or U11077 (N_11077,N_10603,N_10555);
nor U11078 (N_11078,N_10728,N_10567);
xnor U11079 (N_11079,N_10628,N_10645);
xor U11080 (N_11080,N_10743,N_10591);
xor U11081 (N_11081,N_10641,N_10639);
and U11082 (N_11082,N_10550,N_10734);
and U11083 (N_11083,N_10765,N_10790);
or U11084 (N_11084,N_10601,N_10739);
or U11085 (N_11085,N_10693,N_10602);
and U11086 (N_11086,N_10542,N_10640);
or U11087 (N_11087,N_10726,N_10626);
xnor U11088 (N_11088,N_10784,N_10670);
nand U11089 (N_11089,N_10600,N_10573);
or U11090 (N_11090,N_10740,N_10524);
nor U11091 (N_11091,N_10601,N_10655);
nand U11092 (N_11092,N_10544,N_10524);
nor U11093 (N_11093,N_10508,N_10612);
and U11094 (N_11094,N_10569,N_10718);
nor U11095 (N_11095,N_10569,N_10781);
or U11096 (N_11096,N_10624,N_10712);
or U11097 (N_11097,N_10665,N_10565);
or U11098 (N_11098,N_10733,N_10626);
nor U11099 (N_11099,N_10700,N_10678);
nor U11100 (N_11100,N_10971,N_10932);
nand U11101 (N_11101,N_10814,N_10910);
and U11102 (N_11102,N_11097,N_11063);
or U11103 (N_11103,N_10874,N_11051);
or U11104 (N_11104,N_10886,N_10850);
nand U11105 (N_11105,N_11012,N_11060);
or U11106 (N_11106,N_11062,N_11045);
or U11107 (N_11107,N_10859,N_10863);
or U11108 (N_11108,N_11087,N_10849);
xnor U11109 (N_11109,N_10963,N_10846);
or U11110 (N_11110,N_10804,N_10908);
and U11111 (N_11111,N_10950,N_11072);
or U11112 (N_11112,N_10817,N_10939);
and U11113 (N_11113,N_10969,N_11073);
xnor U11114 (N_11114,N_10848,N_11078);
nor U11115 (N_11115,N_11093,N_11009);
xnor U11116 (N_11116,N_11085,N_10942);
xor U11117 (N_11117,N_10845,N_10857);
and U11118 (N_11118,N_10919,N_10974);
xor U11119 (N_11119,N_11084,N_10955);
xnor U11120 (N_11120,N_10821,N_10875);
nor U11121 (N_11121,N_11025,N_10914);
and U11122 (N_11122,N_10809,N_10866);
nand U11123 (N_11123,N_11017,N_10871);
nor U11124 (N_11124,N_10880,N_11043);
xor U11125 (N_11125,N_10893,N_10927);
xnor U11126 (N_11126,N_10807,N_10881);
nor U11127 (N_11127,N_11040,N_10847);
nor U11128 (N_11128,N_10929,N_10991);
nor U11129 (N_11129,N_10907,N_11094);
or U11130 (N_11130,N_10812,N_11034);
nand U11131 (N_11131,N_10889,N_10968);
or U11132 (N_11132,N_11048,N_10964);
and U11133 (N_11133,N_10916,N_10933);
or U11134 (N_11134,N_10873,N_11029);
nand U11135 (N_11135,N_10987,N_10926);
xnor U11136 (N_11136,N_10900,N_10958);
nand U11137 (N_11137,N_10860,N_10839);
nor U11138 (N_11138,N_10823,N_10913);
and U11139 (N_11139,N_11075,N_11019);
xnor U11140 (N_11140,N_11077,N_11064);
or U11141 (N_11141,N_10962,N_10878);
nand U11142 (N_11142,N_10975,N_10903);
nand U11143 (N_11143,N_11057,N_10803);
xnor U11144 (N_11144,N_10992,N_11038);
xnor U11145 (N_11145,N_10935,N_11053);
and U11146 (N_11146,N_10851,N_11020);
xnor U11147 (N_11147,N_11023,N_11055);
nor U11148 (N_11148,N_10905,N_11056);
nor U11149 (N_11149,N_11018,N_10834);
nor U11150 (N_11150,N_10966,N_10830);
nand U11151 (N_11151,N_10802,N_10855);
xnor U11152 (N_11152,N_10922,N_10887);
and U11153 (N_11153,N_11016,N_10923);
and U11154 (N_11154,N_11036,N_11052);
nor U11155 (N_11155,N_10832,N_10999);
nand U11156 (N_11156,N_10957,N_10843);
xnor U11157 (N_11157,N_11079,N_10810);
nor U11158 (N_11158,N_10808,N_10983);
or U11159 (N_11159,N_11008,N_10998);
and U11160 (N_11160,N_10972,N_10824);
nor U11161 (N_11161,N_10853,N_10976);
nand U11162 (N_11162,N_11059,N_11033);
xnor U11163 (N_11163,N_11004,N_10961);
and U11164 (N_11164,N_10829,N_10858);
xor U11165 (N_11165,N_11089,N_10938);
nand U11166 (N_11166,N_11065,N_10937);
xor U11167 (N_11167,N_10985,N_10979);
and U11168 (N_11168,N_10915,N_11046);
or U11169 (N_11169,N_11042,N_10925);
xnor U11170 (N_11170,N_11006,N_11026);
nor U11171 (N_11171,N_10854,N_10896);
xor U11172 (N_11172,N_10838,N_10864);
nor U11173 (N_11173,N_11047,N_10970);
nand U11174 (N_11174,N_10898,N_10884);
and U11175 (N_11175,N_10986,N_11090);
and U11176 (N_11176,N_11031,N_10841);
and U11177 (N_11177,N_10870,N_10902);
nor U11178 (N_11178,N_10947,N_10988);
nor U11179 (N_11179,N_11070,N_11082);
xor U11180 (N_11180,N_10941,N_10813);
nor U11181 (N_11181,N_10872,N_10953);
nor U11182 (N_11182,N_10917,N_10894);
and U11183 (N_11183,N_10982,N_10949);
and U11184 (N_11184,N_10836,N_11010);
xor U11185 (N_11185,N_11099,N_10944);
or U11186 (N_11186,N_11005,N_11068);
or U11187 (N_11187,N_10811,N_10945);
nor U11188 (N_11188,N_11069,N_10997);
nor U11189 (N_11189,N_11081,N_10951);
nand U11190 (N_11190,N_10948,N_10888);
and U11191 (N_11191,N_10954,N_11091);
or U11192 (N_11192,N_11028,N_11088);
and U11193 (N_11193,N_10995,N_11024);
nor U11194 (N_11194,N_10924,N_11032);
xnor U11195 (N_11195,N_11066,N_10862);
and U11196 (N_11196,N_11086,N_11071);
and U11197 (N_11197,N_11002,N_10852);
xor U11198 (N_11198,N_10879,N_11067);
and U11199 (N_11199,N_10911,N_10885);
and U11200 (N_11200,N_10904,N_10967);
nand U11201 (N_11201,N_10956,N_10993);
nand U11202 (N_11202,N_11030,N_10909);
and U11203 (N_11203,N_10895,N_11080);
and U11204 (N_11204,N_10816,N_10869);
nor U11205 (N_11205,N_11011,N_11054);
nor U11206 (N_11206,N_10901,N_10861);
or U11207 (N_11207,N_10936,N_10877);
and U11208 (N_11208,N_10826,N_10996);
nor U11209 (N_11209,N_10876,N_11015);
or U11210 (N_11210,N_10825,N_10994);
nand U11211 (N_11211,N_10952,N_10981);
nor U11212 (N_11212,N_10844,N_10892);
xnor U11213 (N_11213,N_11022,N_10805);
or U11214 (N_11214,N_10882,N_11061);
and U11215 (N_11215,N_10899,N_11039);
and U11216 (N_11216,N_10801,N_11037);
nor U11217 (N_11217,N_10918,N_10868);
nand U11218 (N_11218,N_11058,N_10833);
nor U11219 (N_11219,N_11035,N_10906);
nand U11220 (N_11220,N_11049,N_10842);
nand U11221 (N_11221,N_10928,N_11074);
nand U11222 (N_11222,N_10930,N_10965);
or U11223 (N_11223,N_11041,N_11044);
nand U11224 (N_11224,N_10921,N_10912);
nor U11225 (N_11225,N_10943,N_10989);
nor U11226 (N_11226,N_11083,N_10818);
or U11227 (N_11227,N_11013,N_10897);
or U11228 (N_11228,N_10827,N_10822);
or U11229 (N_11229,N_10973,N_10840);
and U11230 (N_11230,N_10837,N_10977);
nor U11231 (N_11231,N_10831,N_10934);
nor U11232 (N_11232,N_10883,N_11076);
nand U11233 (N_11233,N_11096,N_10806);
nand U11234 (N_11234,N_10890,N_10867);
nand U11235 (N_11235,N_10946,N_10980);
xnor U11236 (N_11236,N_11050,N_10891);
xor U11237 (N_11237,N_10984,N_11095);
nand U11238 (N_11238,N_10920,N_10865);
nor U11239 (N_11239,N_10940,N_11014);
nand U11240 (N_11240,N_11027,N_10978);
nand U11241 (N_11241,N_10820,N_10856);
nor U11242 (N_11242,N_10800,N_10815);
nor U11243 (N_11243,N_11021,N_10819);
and U11244 (N_11244,N_11000,N_10960);
and U11245 (N_11245,N_10828,N_10931);
or U11246 (N_11246,N_11098,N_11003);
nor U11247 (N_11247,N_11001,N_10959);
xnor U11248 (N_11248,N_11007,N_10835);
nand U11249 (N_11249,N_11092,N_10990);
xor U11250 (N_11250,N_10992,N_11007);
and U11251 (N_11251,N_10936,N_11016);
nor U11252 (N_11252,N_10838,N_11060);
xor U11253 (N_11253,N_11044,N_10906);
xnor U11254 (N_11254,N_10817,N_10944);
or U11255 (N_11255,N_10837,N_11095);
and U11256 (N_11256,N_10992,N_10887);
nor U11257 (N_11257,N_10919,N_10972);
and U11258 (N_11258,N_10833,N_10827);
and U11259 (N_11259,N_11020,N_10822);
nor U11260 (N_11260,N_10805,N_10828);
and U11261 (N_11261,N_10996,N_10976);
xnor U11262 (N_11262,N_10886,N_10892);
xor U11263 (N_11263,N_10920,N_10826);
nand U11264 (N_11264,N_11069,N_11038);
or U11265 (N_11265,N_11038,N_11045);
and U11266 (N_11266,N_11092,N_10810);
or U11267 (N_11267,N_10913,N_11058);
xnor U11268 (N_11268,N_11062,N_11033);
or U11269 (N_11269,N_10998,N_11007);
nor U11270 (N_11270,N_10839,N_10904);
nand U11271 (N_11271,N_10847,N_10928);
or U11272 (N_11272,N_10963,N_10933);
xor U11273 (N_11273,N_11084,N_11082);
or U11274 (N_11274,N_10906,N_10934);
nand U11275 (N_11275,N_10840,N_11022);
xor U11276 (N_11276,N_10806,N_10915);
xnor U11277 (N_11277,N_10889,N_10944);
nand U11278 (N_11278,N_10952,N_11048);
and U11279 (N_11279,N_11061,N_10809);
nor U11280 (N_11280,N_10859,N_11071);
and U11281 (N_11281,N_11071,N_10887);
and U11282 (N_11282,N_11095,N_10898);
and U11283 (N_11283,N_11066,N_11080);
xor U11284 (N_11284,N_11092,N_10862);
and U11285 (N_11285,N_11072,N_10902);
and U11286 (N_11286,N_10940,N_10805);
xor U11287 (N_11287,N_11047,N_10807);
nand U11288 (N_11288,N_10866,N_10886);
xor U11289 (N_11289,N_10871,N_10819);
nand U11290 (N_11290,N_11001,N_10926);
and U11291 (N_11291,N_10918,N_10962);
or U11292 (N_11292,N_10956,N_10995);
and U11293 (N_11293,N_11044,N_10828);
and U11294 (N_11294,N_10816,N_11032);
nor U11295 (N_11295,N_10958,N_10905);
and U11296 (N_11296,N_10898,N_11055);
or U11297 (N_11297,N_10858,N_11000);
nor U11298 (N_11298,N_10898,N_11030);
and U11299 (N_11299,N_10930,N_10887);
or U11300 (N_11300,N_10879,N_10981);
xor U11301 (N_11301,N_10999,N_10857);
and U11302 (N_11302,N_10829,N_10918);
nand U11303 (N_11303,N_10887,N_10929);
and U11304 (N_11304,N_10903,N_10828);
or U11305 (N_11305,N_11087,N_10817);
or U11306 (N_11306,N_10905,N_10914);
or U11307 (N_11307,N_10994,N_10971);
and U11308 (N_11308,N_10827,N_11037);
or U11309 (N_11309,N_11097,N_10938);
or U11310 (N_11310,N_10939,N_11045);
nand U11311 (N_11311,N_10902,N_11091);
or U11312 (N_11312,N_11093,N_10851);
nand U11313 (N_11313,N_11046,N_10818);
and U11314 (N_11314,N_10956,N_10942);
xor U11315 (N_11315,N_10859,N_10800);
xor U11316 (N_11316,N_10991,N_11053);
nor U11317 (N_11317,N_11036,N_10882);
nor U11318 (N_11318,N_10989,N_11082);
or U11319 (N_11319,N_10941,N_10949);
or U11320 (N_11320,N_11084,N_10837);
nand U11321 (N_11321,N_10920,N_11003);
or U11322 (N_11322,N_10932,N_10921);
and U11323 (N_11323,N_11097,N_10925);
nand U11324 (N_11324,N_10997,N_10831);
or U11325 (N_11325,N_10821,N_11056);
nand U11326 (N_11326,N_10898,N_11065);
or U11327 (N_11327,N_10979,N_10927);
and U11328 (N_11328,N_11031,N_11070);
nand U11329 (N_11329,N_11055,N_11016);
and U11330 (N_11330,N_10814,N_10856);
and U11331 (N_11331,N_11030,N_10836);
nand U11332 (N_11332,N_10843,N_10844);
or U11333 (N_11333,N_10808,N_10800);
and U11334 (N_11334,N_11087,N_11042);
and U11335 (N_11335,N_11057,N_10900);
nor U11336 (N_11336,N_10998,N_10912);
nand U11337 (N_11337,N_10805,N_11025);
or U11338 (N_11338,N_10920,N_11033);
xor U11339 (N_11339,N_11089,N_11081);
or U11340 (N_11340,N_10904,N_11069);
or U11341 (N_11341,N_11072,N_11052);
xnor U11342 (N_11342,N_11014,N_10894);
xor U11343 (N_11343,N_10866,N_10995);
nand U11344 (N_11344,N_10808,N_10866);
or U11345 (N_11345,N_10993,N_11071);
and U11346 (N_11346,N_11076,N_10841);
nand U11347 (N_11347,N_10830,N_11061);
or U11348 (N_11348,N_11091,N_11094);
and U11349 (N_11349,N_10930,N_10949);
or U11350 (N_11350,N_10845,N_10930);
nand U11351 (N_11351,N_10942,N_10981);
nand U11352 (N_11352,N_11075,N_11054);
nand U11353 (N_11353,N_10901,N_10864);
or U11354 (N_11354,N_10820,N_10874);
nor U11355 (N_11355,N_10934,N_10851);
xnor U11356 (N_11356,N_10853,N_10925);
and U11357 (N_11357,N_10954,N_10886);
or U11358 (N_11358,N_10873,N_11025);
xor U11359 (N_11359,N_11011,N_10828);
or U11360 (N_11360,N_10896,N_11029);
nand U11361 (N_11361,N_11017,N_10839);
nor U11362 (N_11362,N_10909,N_10862);
and U11363 (N_11363,N_10883,N_11027);
nor U11364 (N_11364,N_11020,N_11010);
and U11365 (N_11365,N_10892,N_10993);
and U11366 (N_11366,N_10991,N_11068);
nor U11367 (N_11367,N_10801,N_10927);
and U11368 (N_11368,N_10893,N_10928);
nor U11369 (N_11369,N_11008,N_10823);
or U11370 (N_11370,N_11086,N_11041);
nor U11371 (N_11371,N_11028,N_10973);
nor U11372 (N_11372,N_11066,N_10933);
xnor U11373 (N_11373,N_10998,N_10820);
nor U11374 (N_11374,N_11029,N_10909);
nor U11375 (N_11375,N_11092,N_11039);
nand U11376 (N_11376,N_11085,N_11047);
nor U11377 (N_11377,N_10918,N_10933);
xnor U11378 (N_11378,N_11046,N_10946);
xor U11379 (N_11379,N_10865,N_10849);
nand U11380 (N_11380,N_10929,N_10821);
xor U11381 (N_11381,N_11079,N_10942);
nor U11382 (N_11382,N_11006,N_11046);
xnor U11383 (N_11383,N_11047,N_11003);
and U11384 (N_11384,N_10879,N_10822);
xnor U11385 (N_11385,N_10875,N_10822);
nand U11386 (N_11386,N_11029,N_10908);
xor U11387 (N_11387,N_10815,N_11073);
nor U11388 (N_11388,N_10975,N_10864);
nor U11389 (N_11389,N_10979,N_10948);
xnor U11390 (N_11390,N_11045,N_11081);
nand U11391 (N_11391,N_10930,N_10829);
and U11392 (N_11392,N_10823,N_10970);
and U11393 (N_11393,N_10971,N_11095);
or U11394 (N_11394,N_10958,N_11009);
nor U11395 (N_11395,N_11053,N_10947);
nand U11396 (N_11396,N_10894,N_11047);
or U11397 (N_11397,N_10978,N_11004);
nand U11398 (N_11398,N_11071,N_10873);
and U11399 (N_11399,N_10807,N_10813);
or U11400 (N_11400,N_11202,N_11311);
or U11401 (N_11401,N_11115,N_11239);
nand U11402 (N_11402,N_11133,N_11357);
or U11403 (N_11403,N_11255,N_11237);
nor U11404 (N_11404,N_11379,N_11360);
and U11405 (N_11405,N_11376,N_11352);
and U11406 (N_11406,N_11129,N_11214);
and U11407 (N_11407,N_11331,N_11354);
nand U11408 (N_11408,N_11396,N_11264);
xnor U11409 (N_11409,N_11278,N_11162);
nand U11410 (N_11410,N_11218,N_11228);
nor U11411 (N_11411,N_11235,N_11119);
xor U11412 (N_11412,N_11150,N_11367);
and U11413 (N_11413,N_11280,N_11224);
nand U11414 (N_11414,N_11275,N_11193);
nor U11415 (N_11415,N_11299,N_11212);
nand U11416 (N_11416,N_11206,N_11344);
and U11417 (N_11417,N_11222,N_11223);
nand U11418 (N_11418,N_11363,N_11211);
and U11419 (N_11419,N_11110,N_11329);
xnor U11420 (N_11420,N_11347,N_11371);
xnor U11421 (N_11421,N_11192,N_11167);
nand U11422 (N_11422,N_11317,N_11144);
or U11423 (N_11423,N_11159,N_11180);
xor U11424 (N_11424,N_11301,N_11216);
or U11425 (N_11425,N_11321,N_11345);
xnor U11426 (N_11426,N_11173,N_11296);
and U11427 (N_11427,N_11274,N_11226);
and U11428 (N_11428,N_11297,N_11334);
nand U11429 (N_11429,N_11377,N_11199);
nand U11430 (N_11430,N_11298,N_11335);
xor U11431 (N_11431,N_11361,N_11149);
xor U11432 (N_11432,N_11349,N_11389);
or U11433 (N_11433,N_11249,N_11147);
nor U11434 (N_11434,N_11247,N_11324);
xnor U11435 (N_11435,N_11251,N_11305);
nor U11436 (N_11436,N_11289,N_11156);
nor U11437 (N_11437,N_11260,N_11244);
or U11438 (N_11438,N_11262,N_11269);
and U11439 (N_11439,N_11383,N_11388);
nor U11440 (N_11440,N_11165,N_11241);
or U11441 (N_11441,N_11328,N_11179);
nor U11442 (N_11442,N_11395,N_11210);
or U11443 (N_11443,N_11151,N_11337);
and U11444 (N_11444,N_11390,N_11384);
nor U11445 (N_11445,N_11185,N_11368);
xor U11446 (N_11446,N_11341,N_11233);
nor U11447 (N_11447,N_11333,N_11309);
and U11448 (N_11448,N_11172,N_11370);
xor U11449 (N_11449,N_11327,N_11303);
nand U11450 (N_11450,N_11141,N_11200);
nor U11451 (N_11451,N_11380,N_11254);
xnor U11452 (N_11452,N_11136,N_11177);
nand U11453 (N_11453,N_11188,N_11300);
nand U11454 (N_11454,N_11304,N_11163);
xor U11455 (N_11455,N_11117,N_11273);
or U11456 (N_11456,N_11293,N_11288);
or U11457 (N_11457,N_11307,N_11325);
nand U11458 (N_11458,N_11291,N_11148);
and U11459 (N_11459,N_11339,N_11381);
nand U11460 (N_11460,N_11205,N_11330);
nand U11461 (N_11461,N_11127,N_11178);
and U11462 (N_11462,N_11124,N_11375);
xnor U11463 (N_11463,N_11242,N_11153);
and U11464 (N_11464,N_11365,N_11318);
xnor U11465 (N_11465,N_11314,N_11362);
nand U11466 (N_11466,N_11181,N_11104);
or U11467 (N_11467,N_11230,N_11310);
nor U11468 (N_11468,N_11257,N_11234);
nor U11469 (N_11469,N_11350,N_11154);
xnor U11470 (N_11470,N_11109,N_11290);
and U11471 (N_11471,N_11171,N_11392);
xor U11472 (N_11472,N_11100,N_11277);
nand U11473 (N_11473,N_11338,N_11146);
nor U11474 (N_11474,N_11279,N_11252);
and U11475 (N_11475,N_11320,N_11123);
and U11476 (N_11476,N_11221,N_11281);
nor U11477 (N_11477,N_11316,N_11143);
and U11478 (N_11478,N_11217,N_11322);
nand U11479 (N_11479,N_11258,N_11256);
nand U11480 (N_11480,N_11356,N_11283);
nor U11481 (N_11481,N_11139,N_11243);
nor U11482 (N_11482,N_11116,N_11261);
and U11483 (N_11483,N_11391,N_11340);
xor U11484 (N_11484,N_11213,N_11346);
nand U11485 (N_11485,N_11203,N_11229);
or U11486 (N_11486,N_11306,N_11267);
nand U11487 (N_11487,N_11385,N_11209);
or U11488 (N_11488,N_11236,N_11176);
nand U11489 (N_11489,N_11186,N_11155);
xor U11490 (N_11490,N_11245,N_11366);
nor U11491 (N_11491,N_11166,N_11250);
or U11492 (N_11492,N_11198,N_11382);
or U11493 (N_11493,N_11120,N_11272);
nand U11494 (N_11494,N_11358,N_11302);
nand U11495 (N_11495,N_11187,N_11138);
nor U11496 (N_11496,N_11204,N_11332);
or U11497 (N_11497,N_11207,N_11152);
nand U11498 (N_11498,N_11263,N_11348);
or U11499 (N_11499,N_11369,N_11259);
nand U11500 (N_11500,N_11323,N_11268);
nor U11501 (N_11501,N_11215,N_11292);
nor U11502 (N_11502,N_11169,N_11351);
and U11503 (N_11503,N_11287,N_11378);
and U11504 (N_11504,N_11353,N_11208);
or U11505 (N_11505,N_11227,N_11394);
or U11506 (N_11506,N_11113,N_11220);
and U11507 (N_11507,N_11364,N_11219);
xor U11508 (N_11508,N_11276,N_11231);
xnor U11509 (N_11509,N_11355,N_11114);
nor U11510 (N_11510,N_11160,N_11194);
nand U11511 (N_11511,N_11336,N_11112);
and U11512 (N_11512,N_11266,N_11373);
nand U11513 (N_11513,N_11102,N_11111);
nor U11514 (N_11514,N_11387,N_11196);
or U11515 (N_11515,N_11270,N_11158);
or U11516 (N_11516,N_11175,N_11145);
xnor U11517 (N_11517,N_11106,N_11126);
and U11518 (N_11518,N_11319,N_11182);
and U11519 (N_11519,N_11399,N_11170);
and U11520 (N_11520,N_11295,N_11343);
and U11521 (N_11521,N_11372,N_11359);
or U11522 (N_11522,N_11191,N_11134);
and U11523 (N_11523,N_11118,N_11137);
nor U11524 (N_11524,N_11253,N_11131);
nor U11525 (N_11525,N_11313,N_11184);
or U11526 (N_11526,N_11232,N_11168);
nor U11527 (N_11527,N_11386,N_11140);
xnor U11528 (N_11528,N_11315,N_11286);
nor U11529 (N_11529,N_11125,N_11308);
and U11530 (N_11530,N_11122,N_11183);
nor U11531 (N_11531,N_11284,N_11132);
or U11532 (N_11532,N_11130,N_11271);
or U11533 (N_11533,N_11135,N_11107);
nand U11534 (N_11534,N_11121,N_11312);
nand U11535 (N_11535,N_11265,N_11374);
or U11536 (N_11536,N_11174,N_11195);
nor U11537 (N_11537,N_11240,N_11164);
and U11538 (N_11538,N_11398,N_11103);
or U11539 (N_11539,N_11225,N_11157);
or U11540 (N_11540,N_11201,N_11128);
and U11541 (N_11541,N_11397,N_11190);
and U11542 (N_11542,N_11142,N_11285);
or U11543 (N_11543,N_11342,N_11108);
or U11544 (N_11544,N_11105,N_11326);
nor U11545 (N_11545,N_11161,N_11238);
nand U11546 (N_11546,N_11248,N_11101);
xnor U11547 (N_11547,N_11189,N_11246);
nor U11548 (N_11548,N_11197,N_11393);
nor U11549 (N_11549,N_11294,N_11282);
xnor U11550 (N_11550,N_11115,N_11357);
nor U11551 (N_11551,N_11195,N_11370);
or U11552 (N_11552,N_11350,N_11335);
nor U11553 (N_11553,N_11284,N_11224);
xnor U11554 (N_11554,N_11337,N_11192);
nor U11555 (N_11555,N_11325,N_11261);
nand U11556 (N_11556,N_11137,N_11329);
nand U11557 (N_11557,N_11388,N_11157);
and U11558 (N_11558,N_11373,N_11273);
or U11559 (N_11559,N_11384,N_11259);
or U11560 (N_11560,N_11152,N_11235);
and U11561 (N_11561,N_11212,N_11187);
nor U11562 (N_11562,N_11299,N_11174);
xor U11563 (N_11563,N_11195,N_11347);
nor U11564 (N_11564,N_11337,N_11302);
or U11565 (N_11565,N_11161,N_11222);
nor U11566 (N_11566,N_11279,N_11308);
nor U11567 (N_11567,N_11350,N_11362);
and U11568 (N_11568,N_11187,N_11145);
xor U11569 (N_11569,N_11282,N_11215);
xnor U11570 (N_11570,N_11166,N_11313);
and U11571 (N_11571,N_11185,N_11257);
nand U11572 (N_11572,N_11303,N_11266);
nor U11573 (N_11573,N_11320,N_11363);
and U11574 (N_11574,N_11245,N_11254);
or U11575 (N_11575,N_11244,N_11237);
xnor U11576 (N_11576,N_11273,N_11153);
nor U11577 (N_11577,N_11191,N_11158);
xnor U11578 (N_11578,N_11343,N_11294);
xnor U11579 (N_11579,N_11363,N_11384);
nor U11580 (N_11580,N_11138,N_11111);
nor U11581 (N_11581,N_11206,N_11277);
or U11582 (N_11582,N_11224,N_11150);
and U11583 (N_11583,N_11122,N_11222);
nand U11584 (N_11584,N_11217,N_11131);
nand U11585 (N_11585,N_11106,N_11327);
or U11586 (N_11586,N_11332,N_11252);
or U11587 (N_11587,N_11155,N_11383);
and U11588 (N_11588,N_11293,N_11325);
nor U11589 (N_11589,N_11338,N_11128);
xnor U11590 (N_11590,N_11180,N_11364);
nand U11591 (N_11591,N_11259,N_11173);
nand U11592 (N_11592,N_11391,N_11318);
or U11593 (N_11593,N_11140,N_11190);
nor U11594 (N_11594,N_11137,N_11283);
and U11595 (N_11595,N_11172,N_11146);
and U11596 (N_11596,N_11177,N_11293);
nor U11597 (N_11597,N_11384,N_11221);
and U11598 (N_11598,N_11298,N_11230);
nand U11599 (N_11599,N_11326,N_11168);
nand U11600 (N_11600,N_11292,N_11212);
nand U11601 (N_11601,N_11351,N_11146);
and U11602 (N_11602,N_11171,N_11305);
xnor U11603 (N_11603,N_11214,N_11154);
nand U11604 (N_11604,N_11344,N_11233);
or U11605 (N_11605,N_11161,N_11227);
nor U11606 (N_11606,N_11332,N_11180);
nand U11607 (N_11607,N_11381,N_11223);
or U11608 (N_11608,N_11143,N_11361);
or U11609 (N_11609,N_11126,N_11375);
nor U11610 (N_11610,N_11161,N_11339);
xnor U11611 (N_11611,N_11357,N_11240);
nand U11612 (N_11612,N_11192,N_11306);
and U11613 (N_11613,N_11330,N_11371);
nor U11614 (N_11614,N_11306,N_11242);
nand U11615 (N_11615,N_11224,N_11182);
nor U11616 (N_11616,N_11335,N_11347);
xor U11617 (N_11617,N_11323,N_11172);
nand U11618 (N_11618,N_11149,N_11303);
nor U11619 (N_11619,N_11308,N_11215);
nor U11620 (N_11620,N_11387,N_11333);
or U11621 (N_11621,N_11325,N_11146);
or U11622 (N_11622,N_11195,N_11385);
nand U11623 (N_11623,N_11283,N_11348);
and U11624 (N_11624,N_11201,N_11320);
or U11625 (N_11625,N_11157,N_11360);
and U11626 (N_11626,N_11297,N_11328);
nor U11627 (N_11627,N_11116,N_11159);
and U11628 (N_11628,N_11168,N_11234);
nor U11629 (N_11629,N_11258,N_11371);
or U11630 (N_11630,N_11302,N_11243);
and U11631 (N_11631,N_11223,N_11117);
nor U11632 (N_11632,N_11298,N_11393);
nor U11633 (N_11633,N_11380,N_11374);
nand U11634 (N_11634,N_11335,N_11328);
nand U11635 (N_11635,N_11272,N_11188);
nor U11636 (N_11636,N_11276,N_11299);
nor U11637 (N_11637,N_11339,N_11327);
and U11638 (N_11638,N_11152,N_11358);
nor U11639 (N_11639,N_11363,N_11144);
or U11640 (N_11640,N_11104,N_11215);
or U11641 (N_11641,N_11148,N_11379);
nor U11642 (N_11642,N_11180,N_11120);
xor U11643 (N_11643,N_11158,N_11239);
and U11644 (N_11644,N_11324,N_11311);
xnor U11645 (N_11645,N_11151,N_11284);
xnor U11646 (N_11646,N_11388,N_11372);
or U11647 (N_11647,N_11248,N_11350);
nor U11648 (N_11648,N_11227,N_11179);
or U11649 (N_11649,N_11304,N_11148);
xnor U11650 (N_11650,N_11284,N_11352);
and U11651 (N_11651,N_11384,N_11105);
xnor U11652 (N_11652,N_11250,N_11120);
and U11653 (N_11653,N_11272,N_11275);
xnor U11654 (N_11654,N_11140,N_11215);
or U11655 (N_11655,N_11357,N_11337);
nand U11656 (N_11656,N_11280,N_11331);
nand U11657 (N_11657,N_11389,N_11314);
xor U11658 (N_11658,N_11106,N_11103);
or U11659 (N_11659,N_11235,N_11250);
or U11660 (N_11660,N_11101,N_11137);
nand U11661 (N_11661,N_11144,N_11264);
xor U11662 (N_11662,N_11198,N_11385);
and U11663 (N_11663,N_11347,N_11209);
or U11664 (N_11664,N_11318,N_11173);
xnor U11665 (N_11665,N_11341,N_11327);
xor U11666 (N_11666,N_11333,N_11265);
and U11667 (N_11667,N_11187,N_11303);
and U11668 (N_11668,N_11277,N_11339);
nand U11669 (N_11669,N_11125,N_11325);
nor U11670 (N_11670,N_11129,N_11242);
nor U11671 (N_11671,N_11345,N_11270);
and U11672 (N_11672,N_11388,N_11293);
nand U11673 (N_11673,N_11284,N_11104);
nor U11674 (N_11674,N_11246,N_11152);
nand U11675 (N_11675,N_11328,N_11207);
and U11676 (N_11676,N_11168,N_11186);
xor U11677 (N_11677,N_11247,N_11314);
nand U11678 (N_11678,N_11314,N_11377);
nor U11679 (N_11679,N_11148,N_11320);
nor U11680 (N_11680,N_11245,N_11246);
and U11681 (N_11681,N_11107,N_11352);
or U11682 (N_11682,N_11320,N_11215);
nor U11683 (N_11683,N_11235,N_11291);
nand U11684 (N_11684,N_11357,N_11287);
and U11685 (N_11685,N_11174,N_11162);
xnor U11686 (N_11686,N_11256,N_11244);
nor U11687 (N_11687,N_11206,N_11266);
or U11688 (N_11688,N_11373,N_11295);
or U11689 (N_11689,N_11180,N_11150);
and U11690 (N_11690,N_11220,N_11326);
or U11691 (N_11691,N_11235,N_11309);
and U11692 (N_11692,N_11327,N_11306);
or U11693 (N_11693,N_11151,N_11253);
and U11694 (N_11694,N_11267,N_11216);
xor U11695 (N_11695,N_11160,N_11238);
or U11696 (N_11696,N_11368,N_11314);
xor U11697 (N_11697,N_11155,N_11245);
nand U11698 (N_11698,N_11219,N_11144);
or U11699 (N_11699,N_11373,N_11121);
and U11700 (N_11700,N_11445,N_11584);
nand U11701 (N_11701,N_11545,N_11461);
xor U11702 (N_11702,N_11480,N_11441);
or U11703 (N_11703,N_11623,N_11589);
or U11704 (N_11704,N_11609,N_11427);
or U11705 (N_11705,N_11476,N_11411);
nand U11706 (N_11706,N_11534,N_11674);
nor U11707 (N_11707,N_11574,N_11661);
and U11708 (N_11708,N_11501,N_11564);
nand U11709 (N_11709,N_11648,N_11526);
and U11710 (N_11710,N_11512,N_11601);
or U11711 (N_11711,N_11525,N_11503);
or U11712 (N_11712,N_11467,N_11506);
nand U11713 (N_11713,N_11695,N_11687);
nor U11714 (N_11714,N_11621,N_11537);
nor U11715 (N_11715,N_11699,N_11667);
xor U11716 (N_11716,N_11577,N_11624);
xor U11717 (N_11717,N_11400,N_11446);
or U11718 (N_11718,N_11529,N_11531);
nand U11719 (N_11719,N_11613,N_11603);
nand U11720 (N_11720,N_11638,N_11421);
nor U11721 (N_11721,N_11485,N_11418);
or U11722 (N_11722,N_11471,N_11554);
nor U11723 (N_11723,N_11659,N_11604);
nand U11724 (N_11724,N_11678,N_11553);
nand U11725 (N_11725,N_11488,N_11495);
xor U11726 (N_11726,N_11555,N_11653);
nor U11727 (N_11727,N_11548,N_11683);
or U11728 (N_11728,N_11403,N_11449);
and U11729 (N_11729,N_11662,N_11406);
nor U11730 (N_11730,N_11426,N_11658);
nor U11731 (N_11731,N_11516,N_11669);
xor U11732 (N_11732,N_11620,N_11673);
nor U11733 (N_11733,N_11686,N_11644);
nor U11734 (N_11734,N_11505,N_11413);
or U11735 (N_11735,N_11663,N_11514);
and U11736 (N_11736,N_11435,N_11697);
and U11737 (N_11737,N_11568,N_11448);
and U11738 (N_11738,N_11544,N_11469);
nand U11739 (N_11739,N_11551,N_11596);
or U11740 (N_11740,N_11600,N_11415);
nor U11741 (N_11741,N_11556,N_11493);
nor U11742 (N_11742,N_11492,N_11575);
xor U11743 (N_11743,N_11528,N_11407);
and U11744 (N_11744,N_11549,N_11414);
and U11745 (N_11745,N_11566,N_11474);
nand U11746 (N_11746,N_11666,N_11557);
nor U11747 (N_11747,N_11677,N_11571);
nor U11748 (N_11748,N_11422,N_11473);
nor U11749 (N_11749,N_11558,N_11573);
nor U11750 (N_11750,N_11481,N_11434);
nand U11751 (N_11751,N_11521,N_11567);
nor U11752 (N_11752,N_11684,N_11465);
nand U11753 (N_11753,N_11626,N_11572);
nor U11754 (N_11754,N_11513,N_11420);
or U11755 (N_11755,N_11694,N_11616);
or U11756 (N_11756,N_11450,N_11424);
xnor U11757 (N_11757,N_11691,N_11504);
nor U11758 (N_11758,N_11483,N_11486);
nor U11759 (N_11759,N_11496,N_11565);
and U11760 (N_11760,N_11649,N_11645);
nand U11761 (N_11761,N_11560,N_11462);
nor U11762 (N_11762,N_11665,N_11404);
or U11763 (N_11763,N_11583,N_11543);
or U11764 (N_11764,N_11619,N_11588);
xnor U11765 (N_11765,N_11425,N_11618);
or U11766 (N_11766,N_11532,N_11670);
nand U11767 (N_11767,N_11508,N_11438);
xnor U11768 (N_11768,N_11671,N_11439);
or U11769 (N_11769,N_11550,N_11442);
nand U11770 (N_11770,N_11472,N_11651);
or U11771 (N_11771,N_11646,N_11402);
or U11772 (N_11772,N_11656,N_11436);
xnor U11773 (N_11773,N_11541,N_11538);
nor U11774 (N_11774,N_11685,N_11672);
nor U11775 (N_11775,N_11459,N_11614);
nand U11776 (N_11776,N_11535,N_11497);
and U11777 (N_11777,N_11615,N_11410);
or U11778 (N_11778,N_11692,N_11668);
or U11779 (N_11779,N_11546,N_11429);
or U11780 (N_11780,N_11636,N_11679);
or U11781 (N_11781,N_11579,N_11494);
and U11782 (N_11782,N_11428,N_11696);
xor U11783 (N_11783,N_11511,N_11432);
or U11784 (N_11784,N_11515,N_11605);
nand U11785 (N_11785,N_11581,N_11641);
and U11786 (N_11786,N_11660,N_11466);
nand U11787 (N_11787,N_11519,N_11527);
xor U11788 (N_11788,N_11591,N_11444);
xor U11789 (N_11789,N_11417,N_11639);
xnor U11790 (N_11790,N_11454,N_11552);
and U11791 (N_11791,N_11587,N_11455);
nor U11792 (N_11792,N_11468,N_11416);
nor U11793 (N_11793,N_11632,N_11437);
nor U11794 (N_11794,N_11491,N_11509);
nor U11795 (N_11795,N_11419,N_11561);
and U11796 (N_11796,N_11606,N_11570);
nand U11797 (N_11797,N_11690,N_11478);
and U11798 (N_11798,N_11681,N_11682);
and U11799 (N_11799,N_11460,N_11592);
xnor U11800 (N_11800,N_11507,N_11676);
nor U11801 (N_11801,N_11647,N_11423);
xnor U11802 (N_11802,N_11458,N_11586);
or U11803 (N_11803,N_11582,N_11562);
or U11804 (N_11804,N_11482,N_11447);
and U11805 (N_11805,N_11542,N_11593);
and U11806 (N_11806,N_11457,N_11530);
or U11807 (N_11807,N_11499,N_11675);
and U11808 (N_11808,N_11405,N_11452);
nand U11809 (N_11809,N_11520,N_11634);
or U11810 (N_11810,N_11522,N_11650);
nor U11811 (N_11811,N_11433,N_11498);
nand U11812 (N_11812,N_11479,N_11612);
nor U11813 (N_11813,N_11633,N_11559);
nand U11814 (N_11814,N_11536,N_11635);
xor U11815 (N_11815,N_11451,N_11500);
nand U11816 (N_11816,N_11401,N_11540);
xnor U11817 (N_11817,N_11431,N_11409);
and U11818 (N_11818,N_11608,N_11533);
nand U11819 (N_11819,N_11477,N_11578);
or U11820 (N_11820,N_11599,N_11598);
and U11821 (N_11821,N_11689,N_11664);
and U11822 (N_11822,N_11524,N_11518);
or U11823 (N_11823,N_11517,N_11680);
nand U11824 (N_11824,N_11617,N_11652);
nand U11825 (N_11825,N_11640,N_11563);
nor U11826 (N_11826,N_11487,N_11569);
nand U11827 (N_11827,N_11622,N_11456);
and U11828 (N_11828,N_11627,N_11408);
and U11829 (N_11829,N_11688,N_11611);
and U11830 (N_11830,N_11484,N_11585);
nand U11831 (N_11831,N_11643,N_11607);
nand U11832 (N_11832,N_11594,N_11654);
nor U11833 (N_11833,N_11631,N_11657);
nand U11834 (N_11834,N_11597,N_11595);
nand U11835 (N_11835,N_11630,N_11625);
nand U11836 (N_11836,N_11453,N_11539);
nand U11837 (N_11837,N_11637,N_11602);
and U11838 (N_11838,N_11464,N_11475);
and U11839 (N_11839,N_11489,N_11698);
xnor U11840 (N_11840,N_11440,N_11430);
and U11841 (N_11841,N_11523,N_11629);
nand U11842 (N_11842,N_11628,N_11510);
nor U11843 (N_11843,N_11576,N_11502);
xnor U11844 (N_11844,N_11443,N_11470);
and U11845 (N_11845,N_11580,N_11547);
or U11846 (N_11846,N_11463,N_11642);
xnor U11847 (N_11847,N_11610,N_11590);
xor U11848 (N_11848,N_11655,N_11412);
xor U11849 (N_11849,N_11693,N_11490);
nor U11850 (N_11850,N_11422,N_11526);
xnor U11851 (N_11851,N_11628,N_11447);
and U11852 (N_11852,N_11502,N_11526);
xnor U11853 (N_11853,N_11592,N_11487);
xnor U11854 (N_11854,N_11592,N_11434);
xor U11855 (N_11855,N_11596,N_11457);
nor U11856 (N_11856,N_11611,N_11683);
xnor U11857 (N_11857,N_11620,N_11479);
or U11858 (N_11858,N_11430,N_11453);
nand U11859 (N_11859,N_11675,N_11588);
or U11860 (N_11860,N_11689,N_11547);
and U11861 (N_11861,N_11519,N_11435);
nand U11862 (N_11862,N_11643,N_11496);
xnor U11863 (N_11863,N_11508,N_11658);
nand U11864 (N_11864,N_11585,N_11539);
or U11865 (N_11865,N_11489,N_11585);
nand U11866 (N_11866,N_11453,N_11630);
nand U11867 (N_11867,N_11687,N_11513);
nor U11868 (N_11868,N_11431,N_11593);
and U11869 (N_11869,N_11553,N_11597);
nor U11870 (N_11870,N_11449,N_11567);
or U11871 (N_11871,N_11469,N_11508);
and U11872 (N_11872,N_11600,N_11643);
xor U11873 (N_11873,N_11566,N_11502);
and U11874 (N_11874,N_11573,N_11562);
nand U11875 (N_11875,N_11652,N_11484);
or U11876 (N_11876,N_11511,N_11460);
and U11877 (N_11877,N_11485,N_11555);
nor U11878 (N_11878,N_11485,N_11524);
nand U11879 (N_11879,N_11455,N_11610);
nand U11880 (N_11880,N_11516,N_11553);
nand U11881 (N_11881,N_11583,N_11472);
or U11882 (N_11882,N_11680,N_11646);
nor U11883 (N_11883,N_11611,N_11433);
nand U11884 (N_11884,N_11561,N_11540);
and U11885 (N_11885,N_11421,N_11576);
xor U11886 (N_11886,N_11418,N_11599);
nor U11887 (N_11887,N_11658,N_11522);
or U11888 (N_11888,N_11495,N_11595);
nor U11889 (N_11889,N_11641,N_11430);
nor U11890 (N_11890,N_11671,N_11689);
and U11891 (N_11891,N_11495,N_11683);
nand U11892 (N_11892,N_11409,N_11454);
and U11893 (N_11893,N_11421,N_11500);
nor U11894 (N_11894,N_11676,N_11608);
xnor U11895 (N_11895,N_11655,N_11612);
nand U11896 (N_11896,N_11517,N_11420);
and U11897 (N_11897,N_11500,N_11620);
and U11898 (N_11898,N_11603,N_11591);
xnor U11899 (N_11899,N_11571,N_11667);
or U11900 (N_11900,N_11676,N_11510);
or U11901 (N_11901,N_11525,N_11557);
or U11902 (N_11902,N_11647,N_11654);
and U11903 (N_11903,N_11448,N_11566);
and U11904 (N_11904,N_11546,N_11569);
nor U11905 (N_11905,N_11640,N_11448);
xor U11906 (N_11906,N_11461,N_11406);
or U11907 (N_11907,N_11568,N_11454);
and U11908 (N_11908,N_11609,N_11432);
xnor U11909 (N_11909,N_11421,N_11699);
nand U11910 (N_11910,N_11639,N_11513);
nand U11911 (N_11911,N_11428,N_11567);
or U11912 (N_11912,N_11681,N_11450);
nor U11913 (N_11913,N_11566,N_11458);
nand U11914 (N_11914,N_11585,N_11572);
and U11915 (N_11915,N_11634,N_11667);
or U11916 (N_11916,N_11456,N_11669);
and U11917 (N_11917,N_11531,N_11588);
nor U11918 (N_11918,N_11542,N_11508);
nand U11919 (N_11919,N_11683,N_11599);
nor U11920 (N_11920,N_11644,N_11508);
nor U11921 (N_11921,N_11632,N_11602);
nor U11922 (N_11922,N_11460,N_11496);
or U11923 (N_11923,N_11550,N_11498);
or U11924 (N_11924,N_11498,N_11451);
nor U11925 (N_11925,N_11427,N_11607);
or U11926 (N_11926,N_11516,N_11687);
xor U11927 (N_11927,N_11402,N_11696);
xnor U11928 (N_11928,N_11451,N_11506);
or U11929 (N_11929,N_11526,N_11641);
xnor U11930 (N_11930,N_11673,N_11529);
nor U11931 (N_11931,N_11639,N_11543);
nand U11932 (N_11932,N_11545,N_11490);
nor U11933 (N_11933,N_11610,N_11574);
xnor U11934 (N_11934,N_11600,N_11632);
nor U11935 (N_11935,N_11614,N_11603);
nand U11936 (N_11936,N_11487,N_11407);
or U11937 (N_11937,N_11468,N_11419);
or U11938 (N_11938,N_11699,N_11698);
nand U11939 (N_11939,N_11580,N_11503);
nand U11940 (N_11940,N_11487,N_11615);
and U11941 (N_11941,N_11451,N_11649);
xnor U11942 (N_11942,N_11538,N_11525);
and U11943 (N_11943,N_11560,N_11499);
xor U11944 (N_11944,N_11552,N_11492);
or U11945 (N_11945,N_11447,N_11476);
nor U11946 (N_11946,N_11652,N_11513);
nand U11947 (N_11947,N_11408,N_11480);
or U11948 (N_11948,N_11520,N_11424);
and U11949 (N_11949,N_11504,N_11483);
nand U11950 (N_11950,N_11654,N_11438);
nand U11951 (N_11951,N_11664,N_11514);
nand U11952 (N_11952,N_11661,N_11405);
nor U11953 (N_11953,N_11664,N_11412);
nor U11954 (N_11954,N_11535,N_11613);
nand U11955 (N_11955,N_11447,N_11473);
xnor U11956 (N_11956,N_11527,N_11687);
and U11957 (N_11957,N_11567,N_11459);
xnor U11958 (N_11958,N_11590,N_11501);
or U11959 (N_11959,N_11538,N_11423);
xnor U11960 (N_11960,N_11452,N_11471);
and U11961 (N_11961,N_11597,N_11698);
or U11962 (N_11962,N_11643,N_11687);
nand U11963 (N_11963,N_11496,N_11425);
xnor U11964 (N_11964,N_11494,N_11578);
and U11965 (N_11965,N_11446,N_11591);
xor U11966 (N_11966,N_11581,N_11443);
nor U11967 (N_11967,N_11685,N_11588);
nand U11968 (N_11968,N_11602,N_11696);
xor U11969 (N_11969,N_11665,N_11629);
xor U11970 (N_11970,N_11509,N_11485);
or U11971 (N_11971,N_11597,N_11530);
xor U11972 (N_11972,N_11460,N_11615);
and U11973 (N_11973,N_11421,N_11503);
nand U11974 (N_11974,N_11487,N_11434);
or U11975 (N_11975,N_11433,N_11666);
and U11976 (N_11976,N_11451,N_11499);
or U11977 (N_11977,N_11426,N_11407);
nand U11978 (N_11978,N_11503,N_11645);
nand U11979 (N_11979,N_11566,N_11407);
xor U11980 (N_11980,N_11547,N_11595);
nor U11981 (N_11981,N_11475,N_11459);
and U11982 (N_11982,N_11635,N_11419);
nand U11983 (N_11983,N_11581,N_11457);
nor U11984 (N_11984,N_11696,N_11657);
or U11985 (N_11985,N_11605,N_11670);
nor U11986 (N_11986,N_11585,N_11475);
and U11987 (N_11987,N_11501,N_11534);
and U11988 (N_11988,N_11699,N_11597);
nor U11989 (N_11989,N_11520,N_11443);
nand U11990 (N_11990,N_11575,N_11657);
nand U11991 (N_11991,N_11688,N_11580);
xnor U11992 (N_11992,N_11574,N_11593);
xnor U11993 (N_11993,N_11667,N_11418);
nand U11994 (N_11994,N_11409,N_11576);
or U11995 (N_11995,N_11499,N_11647);
xor U11996 (N_11996,N_11462,N_11403);
or U11997 (N_11997,N_11447,N_11655);
xnor U11998 (N_11998,N_11578,N_11420);
nand U11999 (N_11999,N_11561,N_11571);
nand U12000 (N_12000,N_11951,N_11767);
xnor U12001 (N_12001,N_11955,N_11858);
and U12002 (N_12002,N_11877,N_11717);
or U12003 (N_12003,N_11935,N_11946);
and U12004 (N_12004,N_11974,N_11711);
nand U12005 (N_12005,N_11792,N_11906);
nand U12006 (N_12006,N_11850,N_11771);
xnor U12007 (N_12007,N_11794,N_11878);
nor U12008 (N_12008,N_11710,N_11800);
nand U12009 (N_12009,N_11954,N_11762);
nand U12010 (N_12010,N_11876,N_11927);
nand U12011 (N_12011,N_11857,N_11803);
or U12012 (N_12012,N_11772,N_11962);
nand U12013 (N_12013,N_11854,N_11789);
xnor U12014 (N_12014,N_11702,N_11731);
nor U12015 (N_12015,N_11719,N_11766);
xnor U12016 (N_12016,N_11920,N_11916);
and U12017 (N_12017,N_11904,N_11832);
nand U12018 (N_12018,N_11883,N_11795);
nand U12019 (N_12019,N_11793,N_11805);
and U12020 (N_12020,N_11897,N_11868);
xor U12021 (N_12021,N_11776,N_11949);
nand U12022 (N_12022,N_11888,N_11703);
nor U12023 (N_12023,N_11864,N_11853);
nand U12024 (N_12024,N_11727,N_11957);
nand U12025 (N_12025,N_11783,N_11918);
nor U12026 (N_12026,N_11737,N_11742);
and U12027 (N_12027,N_11726,N_11700);
xor U12028 (N_12028,N_11915,N_11882);
and U12029 (N_12029,N_11929,N_11934);
xnor U12030 (N_12030,N_11744,N_11980);
nor U12031 (N_12031,N_11900,N_11937);
nor U12032 (N_12032,N_11981,N_11777);
or U12033 (N_12033,N_11720,N_11826);
nor U12034 (N_12034,N_11985,N_11862);
nand U12035 (N_12035,N_11791,N_11829);
or U12036 (N_12036,N_11865,N_11938);
nand U12037 (N_12037,N_11716,N_11709);
nor U12038 (N_12038,N_11899,N_11966);
and U12039 (N_12039,N_11705,N_11936);
nand U12040 (N_12040,N_11848,N_11815);
nand U12041 (N_12041,N_11713,N_11953);
nand U12042 (N_12042,N_11843,N_11714);
nor U12043 (N_12043,N_11841,N_11820);
xor U12044 (N_12044,N_11851,N_11859);
or U12045 (N_12045,N_11991,N_11738);
nand U12046 (N_12046,N_11707,N_11736);
nand U12047 (N_12047,N_11788,N_11779);
and U12048 (N_12048,N_11952,N_11922);
or U12049 (N_12049,N_11890,N_11961);
nor U12050 (N_12050,N_11875,N_11901);
or U12051 (N_12051,N_11976,N_11804);
and U12052 (N_12052,N_11913,N_11842);
or U12053 (N_12053,N_11839,N_11836);
nand U12054 (N_12054,N_11960,N_11894);
nor U12055 (N_12055,N_11723,N_11830);
or U12056 (N_12056,N_11739,N_11802);
or U12057 (N_12057,N_11796,N_11898);
or U12058 (N_12058,N_11847,N_11846);
nor U12059 (N_12059,N_11818,N_11910);
or U12060 (N_12060,N_11874,N_11751);
and U12061 (N_12061,N_11835,N_11940);
xor U12062 (N_12062,N_11970,N_11828);
nor U12063 (N_12063,N_11799,N_11807);
xnor U12064 (N_12064,N_11909,N_11964);
nor U12065 (N_12065,N_11860,N_11867);
or U12066 (N_12066,N_11824,N_11706);
nand U12067 (N_12067,N_11749,N_11768);
nand U12068 (N_12068,N_11784,N_11813);
xnor U12069 (N_12069,N_11994,N_11903);
nand U12070 (N_12070,N_11765,N_11973);
nand U12071 (N_12071,N_11925,N_11780);
nor U12072 (N_12072,N_11914,N_11945);
or U12073 (N_12073,N_11701,N_11978);
and U12074 (N_12074,N_11947,N_11752);
and U12075 (N_12075,N_11745,N_11919);
nor U12076 (N_12076,N_11756,N_11785);
or U12077 (N_12077,N_11969,N_11834);
or U12078 (N_12078,N_11782,N_11984);
or U12079 (N_12079,N_11956,N_11753);
and U12080 (N_12080,N_11993,N_11798);
and U12081 (N_12081,N_11942,N_11856);
or U12082 (N_12082,N_11764,N_11972);
xnor U12083 (N_12083,N_11725,N_11816);
xor U12084 (N_12084,N_11928,N_11755);
nand U12085 (N_12085,N_11950,N_11741);
nor U12086 (N_12086,N_11790,N_11965);
nand U12087 (N_12087,N_11730,N_11735);
and U12088 (N_12088,N_11704,N_11775);
nor U12089 (N_12089,N_11822,N_11891);
nor U12090 (N_12090,N_11724,N_11941);
xnor U12091 (N_12091,N_11733,N_11747);
nand U12092 (N_12092,N_11852,N_11886);
xnor U12093 (N_12093,N_11971,N_11827);
xnor U12094 (N_12094,N_11748,N_11825);
xnor U12095 (N_12095,N_11884,N_11734);
and U12096 (N_12096,N_11721,N_11769);
nand U12097 (N_12097,N_11931,N_11786);
nand U12098 (N_12098,N_11917,N_11778);
and U12099 (N_12099,N_11926,N_11740);
nor U12100 (N_12100,N_11712,N_11902);
nand U12101 (N_12101,N_11872,N_11750);
or U12102 (N_12102,N_11995,N_11943);
and U12103 (N_12103,N_11811,N_11773);
xnor U12104 (N_12104,N_11932,N_11758);
nand U12105 (N_12105,N_11990,N_11895);
xor U12106 (N_12106,N_11999,N_11787);
nor U12107 (N_12107,N_11761,N_11968);
nor U12108 (N_12108,N_11743,N_11781);
xnor U12109 (N_12109,N_11992,N_11959);
and U12110 (N_12110,N_11814,N_11746);
or U12111 (N_12111,N_11849,N_11963);
nand U12112 (N_12112,N_11808,N_11844);
nor U12113 (N_12113,N_11908,N_11715);
or U12114 (N_12114,N_11921,N_11838);
and U12115 (N_12115,N_11997,N_11810);
nand U12116 (N_12116,N_11806,N_11879);
xor U12117 (N_12117,N_11923,N_11885);
and U12118 (N_12118,N_11754,N_11729);
xnor U12119 (N_12119,N_11907,N_11939);
xor U12120 (N_12120,N_11770,N_11889);
xnor U12121 (N_12121,N_11801,N_11975);
xnor U12122 (N_12122,N_11870,N_11866);
or U12123 (N_12123,N_11863,N_11967);
and U12124 (N_12124,N_11905,N_11983);
xor U12125 (N_12125,N_11979,N_11924);
and U12126 (N_12126,N_11958,N_11809);
nand U12127 (N_12127,N_11933,N_11873);
nand U12128 (N_12128,N_11759,N_11817);
nor U12129 (N_12129,N_11812,N_11998);
nand U12130 (N_12130,N_11861,N_11912);
and U12131 (N_12131,N_11989,N_11948);
and U12132 (N_12132,N_11887,N_11821);
xnor U12133 (N_12133,N_11797,N_11977);
nand U12134 (N_12134,N_11869,N_11837);
and U12135 (N_12135,N_11757,N_11732);
and U12136 (N_12136,N_11881,N_11930);
or U12137 (N_12137,N_11763,N_11855);
or U12138 (N_12138,N_11986,N_11774);
or U12139 (N_12139,N_11988,N_11987);
and U12140 (N_12140,N_11845,N_11893);
xnor U12141 (N_12141,N_11728,N_11831);
and U12142 (N_12142,N_11722,N_11823);
nand U12143 (N_12143,N_11911,N_11871);
nor U12144 (N_12144,N_11944,N_11760);
nand U12145 (N_12145,N_11833,N_11718);
nor U12146 (N_12146,N_11892,N_11840);
and U12147 (N_12147,N_11819,N_11896);
or U12148 (N_12148,N_11996,N_11880);
or U12149 (N_12149,N_11982,N_11708);
or U12150 (N_12150,N_11914,N_11787);
and U12151 (N_12151,N_11859,N_11834);
or U12152 (N_12152,N_11920,N_11799);
xnor U12153 (N_12153,N_11956,N_11992);
or U12154 (N_12154,N_11804,N_11880);
or U12155 (N_12155,N_11737,N_11736);
or U12156 (N_12156,N_11712,N_11972);
xnor U12157 (N_12157,N_11900,N_11911);
nor U12158 (N_12158,N_11778,N_11837);
nand U12159 (N_12159,N_11762,N_11749);
xnor U12160 (N_12160,N_11914,N_11724);
nor U12161 (N_12161,N_11728,N_11936);
nand U12162 (N_12162,N_11911,N_11748);
xnor U12163 (N_12163,N_11868,N_11984);
nand U12164 (N_12164,N_11871,N_11807);
or U12165 (N_12165,N_11918,N_11909);
and U12166 (N_12166,N_11948,N_11962);
and U12167 (N_12167,N_11747,N_11738);
xnor U12168 (N_12168,N_11911,N_11805);
nor U12169 (N_12169,N_11781,N_11716);
xor U12170 (N_12170,N_11974,N_11912);
nor U12171 (N_12171,N_11915,N_11872);
nand U12172 (N_12172,N_11720,N_11800);
nand U12173 (N_12173,N_11950,N_11793);
nand U12174 (N_12174,N_11936,N_11976);
or U12175 (N_12175,N_11976,N_11811);
nor U12176 (N_12176,N_11848,N_11808);
xor U12177 (N_12177,N_11979,N_11814);
or U12178 (N_12178,N_11730,N_11806);
and U12179 (N_12179,N_11712,N_11988);
xor U12180 (N_12180,N_11899,N_11943);
nand U12181 (N_12181,N_11897,N_11964);
nor U12182 (N_12182,N_11776,N_11713);
nor U12183 (N_12183,N_11994,N_11792);
nor U12184 (N_12184,N_11915,N_11897);
nand U12185 (N_12185,N_11983,N_11779);
nor U12186 (N_12186,N_11774,N_11981);
nor U12187 (N_12187,N_11908,N_11799);
or U12188 (N_12188,N_11972,N_11776);
nand U12189 (N_12189,N_11820,N_11809);
or U12190 (N_12190,N_11771,N_11999);
and U12191 (N_12191,N_11848,N_11798);
nand U12192 (N_12192,N_11961,N_11829);
nor U12193 (N_12193,N_11811,N_11987);
xor U12194 (N_12194,N_11998,N_11983);
and U12195 (N_12195,N_11975,N_11943);
xor U12196 (N_12196,N_11935,N_11900);
nand U12197 (N_12197,N_11930,N_11794);
and U12198 (N_12198,N_11803,N_11917);
nand U12199 (N_12199,N_11980,N_11747);
xor U12200 (N_12200,N_11814,N_11737);
and U12201 (N_12201,N_11730,N_11981);
and U12202 (N_12202,N_11731,N_11931);
xnor U12203 (N_12203,N_11728,N_11839);
nand U12204 (N_12204,N_11953,N_11765);
or U12205 (N_12205,N_11816,N_11945);
or U12206 (N_12206,N_11710,N_11876);
and U12207 (N_12207,N_11885,N_11765);
or U12208 (N_12208,N_11761,N_11792);
nand U12209 (N_12209,N_11944,N_11748);
xor U12210 (N_12210,N_11802,N_11782);
or U12211 (N_12211,N_11947,N_11704);
or U12212 (N_12212,N_11957,N_11811);
nand U12213 (N_12213,N_11945,N_11747);
and U12214 (N_12214,N_11895,N_11957);
and U12215 (N_12215,N_11712,N_11741);
xnor U12216 (N_12216,N_11750,N_11925);
or U12217 (N_12217,N_11761,N_11953);
or U12218 (N_12218,N_11814,N_11751);
or U12219 (N_12219,N_11914,N_11960);
nor U12220 (N_12220,N_11946,N_11840);
nand U12221 (N_12221,N_11962,N_11888);
nor U12222 (N_12222,N_11723,N_11858);
xor U12223 (N_12223,N_11774,N_11742);
and U12224 (N_12224,N_11907,N_11828);
xor U12225 (N_12225,N_11963,N_11749);
and U12226 (N_12226,N_11949,N_11800);
xnor U12227 (N_12227,N_11995,N_11753);
or U12228 (N_12228,N_11708,N_11913);
xor U12229 (N_12229,N_11967,N_11929);
or U12230 (N_12230,N_11951,N_11968);
nor U12231 (N_12231,N_11793,N_11829);
or U12232 (N_12232,N_11768,N_11829);
nor U12233 (N_12233,N_11963,N_11716);
nor U12234 (N_12234,N_11754,N_11853);
nor U12235 (N_12235,N_11934,N_11764);
or U12236 (N_12236,N_11719,N_11931);
or U12237 (N_12237,N_11932,N_11754);
nor U12238 (N_12238,N_11734,N_11887);
xor U12239 (N_12239,N_11811,N_11783);
xnor U12240 (N_12240,N_11881,N_11910);
and U12241 (N_12241,N_11870,N_11858);
nand U12242 (N_12242,N_11797,N_11826);
and U12243 (N_12243,N_11976,N_11803);
or U12244 (N_12244,N_11932,N_11767);
or U12245 (N_12245,N_11804,N_11771);
nand U12246 (N_12246,N_11757,N_11926);
and U12247 (N_12247,N_11903,N_11841);
nand U12248 (N_12248,N_11993,N_11947);
xor U12249 (N_12249,N_11777,N_11859);
nand U12250 (N_12250,N_11829,N_11813);
and U12251 (N_12251,N_11863,N_11768);
and U12252 (N_12252,N_11748,N_11939);
xnor U12253 (N_12253,N_11714,N_11766);
xor U12254 (N_12254,N_11988,N_11963);
and U12255 (N_12255,N_11879,N_11716);
nor U12256 (N_12256,N_11891,N_11817);
and U12257 (N_12257,N_11820,N_11935);
nor U12258 (N_12258,N_11852,N_11773);
nor U12259 (N_12259,N_11991,N_11710);
nor U12260 (N_12260,N_11965,N_11910);
and U12261 (N_12261,N_11883,N_11835);
nor U12262 (N_12262,N_11954,N_11967);
nor U12263 (N_12263,N_11938,N_11795);
and U12264 (N_12264,N_11967,N_11808);
nor U12265 (N_12265,N_11760,N_11796);
or U12266 (N_12266,N_11842,N_11808);
and U12267 (N_12267,N_11801,N_11700);
nor U12268 (N_12268,N_11959,N_11957);
and U12269 (N_12269,N_11910,N_11769);
and U12270 (N_12270,N_11970,N_11976);
and U12271 (N_12271,N_11762,N_11982);
nor U12272 (N_12272,N_11801,N_11925);
or U12273 (N_12273,N_11914,N_11743);
and U12274 (N_12274,N_11712,N_11938);
nor U12275 (N_12275,N_11791,N_11902);
and U12276 (N_12276,N_11812,N_11954);
and U12277 (N_12277,N_11957,N_11786);
xnor U12278 (N_12278,N_11757,N_11736);
and U12279 (N_12279,N_11807,N_11765);
nand U12280 (N_12280,N_11835,N_11724);
or U12281 (N_12281,N_11877,N_11979);
nor U12282 (N_12282,N_11746,N_11820);
and U12283 (N_12283,N_11855,N_11919);
nor U12284 (N_12284,N_11717,N_11753);
and U12285 (N_12285,N_11925,N_11716);
and U12286 (N_12286,N_11946,N_11842);
xor U12287 (N_12287,N_11849,N_11855);
and U12288 (N_12288,N_11816,N_11873);
nor U12289 (N_12289,N_11972,N_11763);
nand U12290 (N_12290,N_11843,N_11984);
xnor U12291 (N_12291,N_11997,N_11790);
nand U12292 (N_12292,N_11940,N_11802);
xnor U12293 (N_12293,N_11925,N_11826);
and U12294 (N_12294,N_11782,N_11765);
and U12295 (N_12295,N_11970,N_11765);
xor U12296 (N_12296,N_11811,N_11861);
xnor U12297 (N_12297,N_11937,N_11813);
nand U12298 (N_12298,N_11983,N_11786);
xor U12299 (N_12299,N_11824,N_11744);
nand U12300 (N_12300,N_12286,N_12056);
or U12301 (N_12301,N_12219,N_12237);
xnor U12302 (N_12302,N_12039,N_12227);
and U12303 (N_12303,N_12203,N_12125);
nor U12304 (N_12304,N_12263,N_12111);
xnor U12305 (N_12305,N_12045,N_12254);
or U12306 (N_12306,N_12072,N_12006);
xor U12307 (N_12307,N_12060,N_12257);
xnor U12308 (N_12308,N_12226,N_12032);
xor U12309 (N_12309,N_12174,N_12143);
nand U12310 (N_12310,N_12275,N_12061);
xnor U12311 (N_12311,N_12102,N_12183);
xor U12312 (N_12312,N_12068,N_12293);
nand U12313 (N_12313,N_12224,N_12059);
and U12314 (N_12314,N_12242,N_12245);
or U12315 (N_12315,N_12049,N_12262);
xnor U12316 (N_12316,N_12236,N_12172);
xnor U12317 (N_12317,N_12155,N_12292);
and U12318 (N_12318,N_12101,N_12199);
and U12319 (N_12319,N_12050,N_12162);
and U12320 (N_12320,N_12122,N_12089);
nand U12321 (N_12321,N_12184,N_12063);
nor U12322 (N_12322,N_12109,N_12233);
nor U12323 (N_12323,N_12285,N_12255);
xnor U12324 (N_12324,N_12094,N_12142);
or U12325 (N_12325,N_12280,N_12106);
or U12326 (N_12326,N_12071,N_12114);
nand U12327 (N_12327,N_12211,N_12024);
xor U12328 (N_12328,N_12279,N_12260);
nand U12329 (N_12329,N_12189,N_12154);
or U12330 (N_12330,N_12197,N_12112);
nand U12331 (N_12331,N_12244,N_12126);
nand U12332 (N_12332,N_12267,N_12241);
nor U12333 (N_12333,N_12149,N_12099);
nand U12334 (N_12334,N_12261,N_12046);
nor U12335 (N_12335,N_12041,N_12167);
and U12336 (N_12336,N_12287,N_12164);
nor U12337 (N_12337,N_12277,N_12294);
xor U12338 (N_12338,N_12284,N_12290);
and U12339 (N_12339,N_12163,N_12210);
nand U12340 (N_12340,N_12234,N_12034);
nand U12341 (N_12341,N_12066,N_12259);
nor U12342 (N_12342,N_12201,N_12077);
or U12343 (N_12343,N_12216,N_12198);
or U12344 (N_12344,N_12202,N_12170);
and U12345 (N_12345,N_12080,N_12095);
xor U12346 (N_12346,N_12073,N_12282);
nor U12347 (N_12347,N_12187,N_12186);
xor U12348 (N_12348,N_12135,N_12212);
or U12349 (N_12349,N_12036,N_12270);
and U12350 (N_12350,N_12214,N_12087);
or U12351 (N_12351,N_12192,N_12191);
and U12352 (N_12352,N_12140,N_12157);
and U12353 (N_12353,N_12204,N_12030);
xnor U12354 (N_12354,N_12119,N_12220);
nand U12355 (N_12355,N_12173,N_12289);
xor U12356 (N_12356,N_12141,N_12139);
nand U12357 (N_12357,N_12103,N_12064);
and U12358 (N_12358,N_12079,N_12252);
xnor U12359 (N_12359,N_12124,N_12017);
or U12360 (N_12360,N_12190,N_12269);
or U12361 (N_12361,N_12169,N_12021);
or U12362 (N_12362,N_12042,N_12028);
nand U12363 (N_12363,N_12092,N_12193);
and U12364 (N_12364,N_12007,N_12108);
or U12365 (N_12365,N_12001,N_12008);
or U12366 (N_12366,N_12247,N_12020);
nor U12367 (N_12367,N_12129,N_12098);
nor U12368 (N_12368,N_12067,N_12209);
or U12369 (N_12369,N_12240,N_12011);
xor U12370 (N_12370,N_12206,N_12086);
xnor U12371 (N_12371,N_12037,N_12018);
xor U12372 (N_12372,N_12096,N_12274);
nand U12373 (N_12373,N_12022,N_12268);
and U12374 (N_12374,N_12065,N_12205);
nand U12375 (N_12375,N_12168,N_12136);
xor U12376 (N_12376,N_12035,N_12093);
or U12377 (N_12377,N_12179,N_12070);
or U12378 (N_12378,N_12053,N_12027);
or U12379 (N_12379,N_12180,N_12055);
xnor U12380 (N_12380,N_12014,N_12273);
nor U12381 (N_12381,N_12009,N_12264);
and U12382 (N_12382,N_12058,N_12196);
nand U12383 (N_12383,N_12047,N_12171);
or U12384 (N_12384,N_12177,N_12083);
nand U12385 (N_12385,N_12150,N_12250);
and U12386 (N_12386,N_12117,N_12110);
nor U12387 (N_12387,N_12074,N_12105);
xnor U12388 (N_12388,N_12249,N_12299);
and U12389 (N_12389,N_12276,N_12288);
nor U12390 (N_12390,N_12272,N_12145);
and U12391 (N_12391,N_12005,N_12075);
nor U12392 (N_12392,N_12128,N_12256);
and U12393 (N_12393,N_12104,N_12218);
nand U12394 (N_12394,N_12081,N_12091);
or U12395 (N_12395,N_12148,N_12243);
nor U12396 (N_12396,N_12121,N_12231);
and U12397 (N_12397,N_12000,N_12085);
nand U12398 (N_12398,N_12152,N_12107);
or U12399 (N_12399,N_12076,N_12217);
and U12400 (N_12400,N_12160,N_12084);
nor U12401 (N_12401,N_12161,N_12131);
xor U12402 (N_12402,N_12040,N_12246);
nor U12403 (N_12403,N_12012,N_12281);
nor U12404 (N_12404,N_12115,N_12052);
or U12405 (N_12405,N_12166,N_12178);
nand U12406 (N_12406,N_12175,N_12044);
and U12407 (N_12407,N_12134,N_12090);
or U12408 (N_12408,N_12144,N_12238);
or U12409 (N_12409,N_12004,N_12116);
nand U12410 (N_12410,N_12147,N_12026);
nand U12411 (N_12411,N_12297,N_12043);
nand U12412 (N_12412,N_12151,N_12278);
or U12413 (N_12413,N_12132,N_12031);
xnor U12414 (N_12414,N_12158,N_12133);
nor U12415 (N_12415,N_12230,N_12010);
nor U12416 (N_12416,N_12195,N_12228);
or U12417 (N_12417,N_12113,N_12146);
nor U12418 (N_12418,N_12069,N_12025);
or U12419 (N_12419,N_12265,N_12251);
or U12420 (N_12420,N_12295,N_12221);
or U12421 (N_12421,N_12038,N_12029);
or U12422 (N_12422,N_12078,N_12291);
and U12423 (N_12423,N_12153,N_12023);
and U12424 (N_12424,N_12100,N_12182);
nor U12425 (N_12425,N_12003,N_12054);
nor U12426 (N_12426,N_12120,N_12225);
nor U12427 (N_12427,N_12222,N_12013);
nor U12428 (N_12428,N_12130,N_12207);
nor U12429 (N_12429,N_12271,N_12019);
and U12430 (N_12430,N_12235,N_12016);
or U12431 (N_12431,N_12159,N_12239);
and U12432 (N_12432,N_12127,N_12015);
and U12433 (N_12433,N_12223,N_12208);
nor U12434 (N_12434,N_12194,N_12097);
or U12435 (N_12435,N_12057,N_12229);
and U12436 (N_12436,N_12298,N_12051);
xnor U12437 (N_12437,N_12176,N_12200);
xnor U12438 (N_12438,N_12266,N_12156);
nor U12439 (N_12439,N_12296,N_12123);
nand U12440 (N_12440,N_12033,N_12248);
nand U12441 (N_12441,N_12213,N_12062);
and U12442 (N_12442,N_12082,N_12048);
xor U12443 (N_12443,N_12253,N_12188);
nand U12444 (N_12444,N_12215,N_12185);
and U12445 (N_12445,N_12258,N_12118);
or U12446 (N_12446,N_12232,N_12088);
nand U12447 (N_12447,N_12165,N_12181);
or U12448 (N_12448,N_12002,N_12138);
and U12449 (N_12449,N_12283,N_12137);
nand U12450 (N_12450,N_12285,N_12170);
nand U12451 (N_12451,N_12039,N_12031);
nor U12452 (N_12452,N_12119,N_12250);
nor U12453 (N_12453,N_12035,N_12084);
nor U12454 (N_12454,N_12143,N_12057);
nor U12455 (N_12455,N_12006,N_12251);
xor U12456 (N_12456,N_12009,N_12113);
nand U12457 (N_12457,N_12195,N_12008);
nor U12458 (N_12458,N_12033,N_12127);
nand U12459 (N_12459,N_12173,N_12074);
nor U12460 (N_12460,N_12190,N_12143);
nor U12461 (N_12461,N_12134,N_12112);
and U12462 (N_12462,N_12269,N_12129);
nand U12463 (N_12463,N_12126,N_12145);
xnor U12464 (N_12464,N_12045,N_12178);
and U12465 (N_12465,N_12044,N_12031);
or U12466 (N_12466,N_12201,N_12117);
and U12467 (N_12467,N_12103,N_12194);
xor U12468 (N_12468,N_12218,N_12063);
or U12469 (N_12469,N_12046,N_12175);
xor U12470 (N_12470,N_12062,N_12154);
nor U12471 (N_12471,N_12235,N_12112);
and U12472 (N_12472,N_12053,N_12183);
and U12473 (N_12473,N_12079,N_12247);
or U12474 (N_12474,N_12040,N_12019);
nand U12475 (N_12475,N_12226,N_12060);
xor U12476 (N_12476,N_12184,N_12259);
xor U12477 (N_12477,N_12087,N_12191);
and U12478 (N_12478,N_12047,N_12206);
or U12479 (N_12479,N_12128,N_12125);
nand U12480 (N_12480,N_12027,N_12168);
nor U12481 (N_12481,N_12043,N_12254);
and U12482 (N_12482,N_12032,N_12074);
or U12483 (N_12483,N_12276,N_12019);
and U12484 (N_12484,N_12146,N_12243);
nand U12485 (N_12485,N_12246,N_12045);
xnor U12486 (N_12486,N_12262,N_12098);
and U12487 (N_12487,N_12226,N_12205);
xnor U12488 (N_12488,N_12191,N_12214);
nor U12489 (N_12489,N_12051,N_12014);
nor U12490 (N_12490,N_12287,N_12212);
or U12491 (N_12491,N_12103,N_12216);
and U12492 (N_12492,N_12027,N_12175);
xor U12493 (N_12493,N_12103,N_12137);
and U12494 (N_12494,N_12005,N_12196);
or U12495 (N_12495,N_12241,N_12200);
nand U12496 (N_12496,N_12036,N_12047);
or U12497 (N_12497,N_12013,N_12148);
nor U12498 (N_12498,N_12253,N_12238);
and U12499 (N_12499,N_12027,N_12031);
xor U12500 (N_12500,N_12046,N_12070);
or U12501 (N_12501,N_12048,N_12074);
nand U12502 (N_12502,N_12259,N_12062);
xnor U12503 (N_12503,N_12054,N_12260);
nor U12504 (N_12504,N_12031,N_12054);
or U12505 (N_12505,N_12232,N_12287);
nor U12506 (N_12506,N_12232,N_12242);
and U12507 (N_12507,N_12033,N_12189);
xnor U12508 (N_12508,N_12223,N_12159);
and U12509 (N_12509,N_12257,N_12172);
nor U12510 (N_12510,N_12002,N_12036);
and U12511 (N_12511,N_12023,N_12043);
nand U12512 (N_12512,N_12054,N_12191);
nor U12513 (N_12513,N_12233,N_12281);
xnor U12514 (N_12514,N_12013,N_12144);
xnor U12515 (N_12515,N_12045,N_12063);
or U12516 (N_12516,N_12299,N_12285);
nor U12517 (N_12517,N_12062,N_12294);
or U12518 (N_12518,N_12017,N_12184);
nand U12519 (N_12519,N_12229,N_12161);
or U12520 (N_12520,N_12186,N_12013);
nand U12521 (N_12521,N_12081,N_12065);
nor U12522 (N_12522,N_12049,N_12203);
or U12523 (N_12523,N_12111,N_12298);
nor U12524 (N_12524,N_12120,N_12228);
xnor U12525 (N_12525,N_12248,N_12080);
xor U12526 (N_12526,N_12276,N_12065);
nor U12527 (N_12527,N_12241,N_12111);
nor U12528 (N_12528,N_12193,N_12015);
nor U12529 (N_12529,N_12210,N_12172);
nor U12530 (N_12530,N_12298,N_12032);
and U12531 (N_12531,N_12012,N_12114);
nand U12532 (N_12532,N_12283,N_12133);
nand U12533 (N_12533,N_12250,N_12006);
nor U12534 (N_12534,N_12144,N_12224);
xor U12535 (N_12535,N_12089,N_12195);
nand U12536 (N_12536,N_12107,N_12163);
nor U12537 (N_12537,N_12129,N_12108);
nand U12538 (N_12538,N_12223,N_12232);
nand U12539 (N_12539,N_12109,N_12225);
or U12540 (N_12540,N_12014,N_12297);
nor U12541 (N_12541,N_12035,N_12094);
nor U12542 (N_12542,N_12088,N_12084);
nand U12543 (N_12543,N_12250,N_12111);
nor U12544 (N_12544,N_12192,N_12032);
and U12545 (N_12545,N_12096,N_12224);
nor U12546 (N_12546,N_12264,N_12058);
nor U12547 (N_12547,N_12074,N_12296);
or U12548 (N_12548,N_12182,N_12147);
nor U12549 (N_12549,N_12161,N_12091);
nor U12550 (N_12550,N_12044,N_12254);
nor U12551 (N_12551,N_12095,N_12245);
xor U12552 (N_12552,N_12122,N_12267);
nand U12553 (N_12553,N_12262,N_12014);
nand U12554 (N_12554,N_12092,N_12100);
or U12555 (N_12555,N_12119,N_12078);
and U12556 (N_12556,N_12241,N_12185);
and U12557 (N_12557,N_12145,N_12013);
or U12558 (N_12558,N_12049,N_12283);
nor U12559 (N_12559,N_12097,N_12091);
or U12560 (N_12560,N_12208,N_12220);
or U12561 (N_12561,N_12292,N_12050);
xnor U12562 (N_12562,N_12030,N_12055);
xnor U12563 (N_12563,N_12159,N_12061);
xor U12564 (N_12564,N_12101,N_12184);
xnor U12565 (N_12565,N_12181,N_12044);
nor U12566 (N_12566,N_12031,N_12176);
nand U12567 (N_12567,N_12146,N_12142);
xor U12568 (N_12568,N_12074,N_12208);
or U12569 (N_12569,N_12252,N_12099);
or U12570 (N_12570,N_12222,N_12245);
xor U12571 (N_12571,N_12125,N_12085);
nor U12572 (N_12572,N_12203,N_12207);
and U12573 (N_12573,N_12009,N_12122);
or U12574 (N_12574,N_12121,N_12061);
xnor U12575 (N_12575,N_12211,N_12087);
xnor U12576 (N_12576,N_12030,N_12291);
nor U12577 (N_12577,N_12200,N_12033);
or U12578 (N_12578,N_12295,N_12056);
xor U12579 (N_12579,N_12161,N_12200);
nand U12580 (N_12580,N_12155,N_12296);
or U12581 (N_12581,N_12284,N_12074);
or U12582 (N_12582,N_12175,N_12262);
and U12583 (N_12583,N_12016,N_12294);
or U12584 (N_12584,N_12190,N_12098);
and U12585 (N_12585,N_12048,N_12249);
nand U12586 (N_12586,N_12190,N_12205);
and U12587 (N_12587,N_12061,N_12108);
and U12588 (N_12588,N_12027,N_12043);
nand U12589 (N_12589,N_12025,N_12030);
or U12590 (N_12590,N_12015,N_12123);
xnor U12591 (N_12591,N_12232,N_12258);
nor U12592 (N_12592,N_12223,N_12019);
xnor U12593 (N_12593,N_12149,N_12027);
and U12594 (N_12594,N_12163,N_12058);
and U12595 (N_12595,N_12223,N_12295);
nor U12596 (N_12596,N_12041,N_12263);
or U12597 (N_12597,N_12251,N_12196);
and U12598 (N_12598,N_12280,N_12052);
nor U12599 (N_12599,N_12181,N_12225);
or U12600 (N_12600,N_12460,N_12578);
or U12601 (N_12601,N_12502,N_12495);
xor U12602 (N_12602,N_12565,N_12331);
or U12603 (N_12603,N_12351,N_12568);
nand U12604 (N_12604,N_12396,N_12592);
nor U12605 (N_12605,N_12473,N_12304);
and U12606 (N_12606,N_12507,N_12597);
nand U12607 (N_12607,N_12463,N_12591);
or U12608 (N_12608,N_12374,N_12394);
xnor U12609 (N_12609,N_12350,N_12328);
or U12610 (N_12610,N_12343,N_12488);
or U12611 (N_12611,N_12531,N_12423);
nand U12612 (N_12612,N_12588,N_12530);
or U12613 (N_12613,N_12528,N_12490);
xor U12614 (N_12614,N_12389,N_12334);
xor U12615 (N_12615,N_12519,N_12478);
or U12616 (N_12616,N_12563,N_12527);
xor U12617 (N_12617,N_12403,N_12566);
xnor U12618 (N_12618,N_12518,N_12479);
xnor U12619 (N_12619,N_12316,N_12310);
nand U12620 (N_12620,N_12366,N_12329);
and U12621 (N_12621,N_12554,N_12431);
nor U12622 (N_12622,N_12562,N_12544);
and U12623 (N_12623,N_12494,N_12582);
xor U12624 (N_12624,N_12577,N_12349);
xor U12625 (N_12625,N_12451,N_12429);
nor U12626 (N_12626,N_12355,N_12556);
and U12627 (N_12627,N_12443,N_12402);
nor U12628 (N_12628,N_12560,N_12324);
xnor U12629 (N_12629,N_12462,N_12322);
nor U12630 (N_12630,N_12342,N_12599);
xor U12631 (N_12631,N_12552,N_12598);
xor U12632 (N_12632,N_12520,N_12533);
nor U12633 (N_12633,N_12506,N_12487);
nand U12634 (N_12634,N_12433,N_12421);
nand U12635 (N_12635,N_12492,N_12541);
or U12636 (N_12636,N_12486,N_12457);
and U12637 (N_12637,N_12575,N_12307);
nand U12638 (N_12638,N_12428,N_12344);
or U12639 (N_12639,N_12424,N_12373);
or U12640 (N_12640,N_12557,N_12455);
or U12641 (N_12641,N_12559,N_12441);
xnor U12642 (N_12642,N_12318,N_12500);
and U12643 (N_12643,N_12364,N_12372);
nand U12644 (N_12644,N_12311,N_12337);
xor U12645 (N_12645,N_12300,N_12580);
nand U12646 (N_12646,N_12320,N_12529);
and U12647 (N_12647,N_12362,N_12303);
and U12648 (N_12648,N_12489,N_12589);
xnor U12649 (N_12649,N_12471,N_12392);
nor U12650 (N_12650,N_12442,N_12384);
and U12651 (N_12651,N_12315,N_12590);
and U12652 (N_12652,N_12425,N_12593);
and U12653 (N_12653,N_12321,N_12436);
xor U12654 (N_12654,N_12444,N_12543);
and U12655 (N_12655,N_12369,N_12553);
or U12656 (N_12656,N_12569,N_12395);
or U12657 (N_12657,N_12417,N_12409);
nor U12658 (N_12658,N_12503,N_12522);
nand U12659 (N_12659,N_12330,N_12539);
xor U12660 (N_12660,N_12356,N_12536);
xnor U12661 (N_12661,N_12561,N_12537);
and U12662 (N_12662,N_12549,N_12352);
nor U12663 (N_12663,N_12341,N_12439);
xor U12664 (N_12664,N_12564,N_12516);
nand U12665 (N_12665,N_12491,N_12447);
nand U12666 (N_12666,N_12474,N_12584);
and U12667 (N_12667,N_12432,N_12523);
or U12668 (N_12668,N_12435,N_12312);
xnor U12669 (N_12669,N_12482,N_12466);
or U12670 (N_12670,N_12416,N_12378);
xnor U12671 (N_12671,N_12586,N_12326);
nor U12672 (N_12672,N_12576,N_12302);
and U12673 (N_12673,N_12480,N_12357);
xor U12674 (N_12674,N_12380,N_12393);
or U12675 (N_12675,N_12524,N_12540);
nor U12676 (N_12676,N_12420,N_12390);
nand U12677 (N_12677,N_12314,N_12477);
nor U12678 (N_12678,N_12510,N_12313);
nor U12679 (N_12679,N_12496,N_12358);
and U12680 (N_12680,N_12332,N_12365);
and U12681 (N_12681,N_12407,N_12335);
nor U12682 (N_12682,N_12572,N_12458);
nor U12683 (N_12683,N_12382,N_12521);
or U12684 (N_12684,N_12448,N_12469);
or U12685 (N_12685,N_12596,N_12381);
nand U12686 (N_12686,N_12360,N_12585);
xor U12687 (N_12687,N_12445,N_12414);
and U12688 (N_12688,N_12309,N_12472);
and U12689 (N_12689,N_12450,N_12499);
or U12690 (N_12690,N_12422,N_12485);
nand U12691 (N_12691,N_12498,N_12579);
xor U12692 (N_12692,N_12319,N_12308);
xor U12693 (N_12693,N_12323,N_12570);
nand U12694 (N_12694,N_12456,N_12400);
and U12695 (N_12695,N_12345,N_12508);
xnor U12696 (N_12696,N_12548,N_12468);
xnor U12697 (N_12697,N_12449,N_12375);
nand U12698 (N_12698,N_12410,N_12464);
nor U12699 (N_12699,N_12391,N_12419);
or U12700 (N_12700,N_12571,N_12383);
and U12701 (N_12701,N_12301,N_12574);
xor U12702 (N_12702,N_12504,N_12434);
and U12703 (N_12703,N_12340,N_12534);
nand U12704 (N_12704,N_12339,N_12333);
nand U12705 (N_12705,N_12336,N_12399);
and U12706 (N_12706,N_12346,N_12317);
or U12707 (N_12707,N_12446,N_12470);
and U12708 (N_12708,N_12412,N_12397);
nand U12709 (N_12709,N_12515,N_12595);
nor U12710 (N_12710,N_12501,N_12567);
and U12711 (N_12711,N_12532,N_12376);
nand U12712 (N_12712,N_12481,N_12587);
nand U12713 (N_12713,N_12546,N_12388);
and U12714 (N_12714,N_12368,N_12493);
or U12715 (N_12715,N_12367,N_12370);
nor U12716 (N_12716,N_12483,N_12535);
xnor U12717 (N_12717,N_12514,N_12411);
nor U12718 (N_12718,N_12359,N_12551);
nor U12719 (N_12719,N_12379,N_12452);
xor U12720 (N_12720,N_12550,N_12467);
nor U12721 (N_12721,N_12581,N_12413);
nand U12722 (N_12722,N_12525,N_12459);
or U12723 (N_12723,N_12348,N_12338);
xnor U12724 (N_12724,N_12377,N_12347);
nand U12725 (N_12725,N_12484,N_12371);
or U12726 (N_12726,N_12461,N_12545);
and U12727 (N_12727,N_12387,N_12542);
nor U12728 (N_12728,N_12361,N_12398);
nor U12729 (N_12729,N_12426,N_12511);
or U12730 (N_12730,N_12306,N_12354);
or U12731 (N_12731,N_12430,N_12555);
nor U12732 (N_12732,N_12512,N_12427);
or U12733 (N_12733,N_12408,N_12405);
xnor U12734 (N_12734,N_12415,N_12517);
nor U12735 (N_12735,N_12418,N_12453);
and U12736 (N_12736,N_12386,N_12475);
and U12737 (N_12737,N_12547,N_12558);
xor U12738 (N_12738,N_12465,N_12476);
and U12739 (N_12739,N_12538,N_12509);
nand U12740 (N_12740,N_12454,N_12325);
and U12741 (N_12741,N_12573,N_12513);
xor U12742 (N_12742,N_12406,N_12438);
and U12743 (N_12743,N_12404,N_12497);
nor U12744 (N_12744,N_12363,N_12594);
nor U12745 (N_12745,N_12505,N_12583);
nor U12746 (N_12746,N_12327,N_12385);
or U12747 (N_12747,N_12353,N_12437);
or U12748 (N_12748,N_12401,N_12440);
xor U12749 (N_12749,N_12526,N_12305);
or U12750 (N_12750,N_12422,N_12539);
or U12751 (N_12751,N_12513,N_12440);
or U12752 (N_12752,N_12530,N_12514);
xor U12753 (N_12753,N_12323,N_12517);
and U12754 (N_12754,N_12391,N_12463);
nor U12755 (N_12755,N_12372,N_12517);
or U12756 (N_12756,N_12460,N_12494);
or U12757 (N_12757,N_12562,N_12411);
or U12758 (N_12758,N_12510,N_12356);
nand U12759 (N_12759,N_12302,N_12507);
xnor U12760 (N_12760,N_12484,N_12467);
xnor U12761 (N_12761,N_12556,N_12331);
nor U12762 (N_12762,N_12364,N_12481);
and U12763 (N_12763,N_12569,N_12383);
and U12764 (N_12764,N_12572,N_12526);
or U12765 (N_12765,N_12529,N_12339);
xor U12766 (N_12766,N_12595,N_12305);
xor U12767 (N_12767,N_12537,N_12457);
nand U12768 (N_12768,N_12506,N_12305);
and U12769 (N_12769,N_12338,N_12565);
nand U12770 (N_12770,N_12359,N_12399);
xnor U12771 (N_12771,N_12365,N_12432);
xor U12772 (N_12772,N_12571,N_12355);
xnor U12773 (N_12773,N_12440,N_12553);
or U12774 (N_12774,N_12577,N_12531);
nor U12775 (N_12775,N_12481,N_12334);
and U12776 (N_12776,N_12380,N_12356);
and U12777 (N_12777,N_12457,N_12563);
and U12778 (N_12778,N_12313,N_12466);
nor U12779 (N_12779,N_12593,N_12563);
and U12780 (N_12780,N_12587,N_12397);
nand U12781 (N_12781,N_12561,N_12403);
nand U12782 (N_12782,N_12381,N_12375);
or U12783 (N_12783,N_12350,N_12404);
xnor U12784 (N_12784,N_12318,N_12457);
or U12785 (N_12785,N_12424,N_12440);
nor U12786 (N_12786,N_12349,N_12338);
or U12787 (N_12787,N_12311,N_12417);
or U12788 (N_12788,N_12386,N_12452);
nand U12789 (N_12789,N_12517,N_12398);
or U12790 (N_12790,N_12347,N_12594);
xnor U12791 (N_12791,N_12391,N_12339);
and U12792 (N_12792,N_12344,N_12424);
nand U12793 (N_12793,N_12583,N_12598);
xor U12794 (N_12794,N_12477,N_12548);
or U12795 (N_12795,N_12586,N_12450);
nor U12796 (N_12796,N_12445,N_12384);
xor U12797 (N_12797,N_12596,N_12556);
nand U12798 (N_12798,N_12379,N_12329);
xnor U12799 (N_12799,N_12393,N_12318);
xor U12800 (N_12800,N_12322,N_12564);
nand U12801 (N_12801,N_12594,N_12338);
xnor U12802 (N_12802,N_12304,N_12391);
xor U12803 (N_12803,N_12459,N_12564);
and U12804 (N_12804,N_12570,N_12465);
and U12805 (N_12805,N_12531,N_12441);
nor U12806 (N_12806,N_12405,N_12407);
nor U12807 (N_12807,N_12519,N_12470);
or U12808 (N_12808,N_12449,N_12417);
nand U12809 (N_12809,N_12557,N_12499);
and U12810 (N_12810,N_12500,N_12389);
nand U12811 (N_12811,N_12586,N_12466);
and U12812 (N_12812,N_12397,N_12414);
nor U12813 (N_12813,N_12448,N_12309);
nor U12814 (N_12814,N_12592,N_12424);
xor U12815 (N_12815,N_12305,N_12323);
nor U12816 (N_12816,N_12492,N_12342);
nor U12817 (N_12817,N_12436,N_12589);
xnor U12818 (N_12818,N_12300,N_12386);
and U12819 (N_12819,N_12306,N_12364);
xnor U12820 (N_12820,N_12443,N_12430);
nor U12821 (N_12821,N_12334,N_12538);
xor U12822 (N_12822,N_12462,N_12498);
and U12823 (N_12823,N_12330,N_12449);
nor U12824 (N_12824,N_12395,N_12530);
xor U12825 (N_12825,N_12454,N_12587);
xor U12826 (N_12826,N_12565,N_12342);
nor U12827 (N_12827,N_12342,N_12463);
xor U12828 (N_12828,N_12540,N_12375);
nand U12829 (N_12829,N_12314,N_12560);
or U12830 (N_12830,N_12562,N_12550);
and U12831 (N_12831,N_12349,N_12393);
or U12832 (N_12832,N_12399,N_12515);
or U12833 (N_12833,N_12535,N_12580);
xnor U12834 (N_12834,N_12542,N_12572);
nor U12835 (N_12835,N_12476,N_12544);
xnor U12836 (N_12836,N_12392,N_12326);
nor U12837 (N_12837,N_12307,N_12402);
nand U12838 (N_12838,N_12403,N_12434);
xnor U12839 (N_12839,N_12335,N_12504);
nand U12840 (N_12840,N_12330,N_12424);
and U12841 (N_12841,N_12494,N_12416);
and U12842 (N_12842,N_12346,N_12476);
nor U12843 (N_12843,N_12465,N_12359);
and U12844 (N_12844,N_12522,N_12329);
and U12845 (N_12845,N_12491,N_12357);
nor U12846 (N_12846,N_12528,N_12585);
or U12847 (N_12847,N_12569,N_12370);
or U12848 (N_12848,N_12332,N_12481);
or U12849 (N_12849,N_12371,N_12482);
xnor U12850 (N_12850,N_12530,N_12354);
nor U12851 (N_12851,N_12361,N_12451);
and U12852 (N_12852,N_12496,N_12304);
or U12853 (N_12853,N_12597,N_12588);
nor U12854 (N_12854,N_12422,N_12438);
nor U12855 (N_12855,N_12573,N_12380);
or U12856 (N_12856,N_12589,N_12432);
nand U12857 (N_12857,N_12571,N_12468);
or U12858 (N_12858,N_12322,N_12405);
nor U12859 (N_12859,N_12339,N_12386);
nand U12860 (N_12860,N_12583,N_12386);
and U12861 (N_12861,N_12474,N_12568);
and U12862 (N_12862,N_12528,N_12365);
or U12863 (N_12863,N_12546,N_12596);
nand U12864 (N_12864,N_12512,N_12383);
or U12865 (N_12865,N_12488,N_12550);
nor U12866 (N_12866,N_12472,N_12462);
xor U12867 (N_12867,N_12364,N_12444);
and U12868 (N_12868,N_12303,N_12490);
or U12869 (N_12869,N_12524,N_12470);
nand U12870 (N_12870,N_12575,N_12550);
and U12871 (N_12871,N_12318,N_12409);
xor U12872 (N_12872,N_12377,N_12461);
xnor U12873 (N_12873,N_12328,N_12446);
and U12874 (N_12874,N_12323,N_12397);
nor U12875 (N_12875,N_12564,N_12339);
and U12876 (N_12876,N_12559,N_12440);
or U12877 (N_12877,N_12525,N_12408);
or U12878 (N_12878,N_12562,N_12525);
xnor U12879 (N_12879,N_12469,N_12377);
nor U12880 (N_12880,N_12586,N_12402);
or U12881 (N_12881,N_12400,N_12503);
or U12882 (N_12882,N_12521,N_12563);
xnor U12883 (N_12883,N_12516,N_12462);
and U12884 (N_12884,N_12362,N_12342);
nor U12885 (N_12885,N_12571,N_12447);
and U12886 (N_12886,N_12516,N_12409);
or U12887 (N_12887,N_12468,N_12330);
nand U12888 (N_12888,N_12550,N_12582);
xor U12889 (N_12889,N_12387,N_12337);
or U12890 (N_12890,N_12350,N_12353);
and U12891 (N_12891,N_12537,N_12463);
nor U12892 (N_12892,N_12392,N_12421);
nor U12893 (N_12893,N_12518,N_12549);
nand U12894 (N_12894,N_12320,N_12503);
and U12895 (N_12895,N_12392,N_12515);
nor U12896 (N_12896,N_12570,N_12300);
xnor U12897 (N_12897,N_12363,N_12538);
or U12898 (N_12898,N_12389,N_12393);
xnor U12899 (N_12899,N_12482,N_12593);
nor U12900 (N_12900,N_12868,N_12676);
nand U12901 (N_12901,N_12734,N_12839);
xnor U12902 (N_12902,N_12895,N_12763);
or U12903 (N_12903,N_12606,N_12664);
nand U12904 (N_12904,N_12767,N_12883);
xnor U12905 (N_12905,N_12702,N_12741);
and U12906 (N_12906,N_12844,N_12604);
nand U12907 (N_12907,N_12771,N_12810);
xnor U12908 (N_12908,N_12808,N_12815);
or U12909 (N_12909,N_12758,N_12634);
nand U12910 (N_12910,N_12750,N_12677);
or U12911 (N_12911,N_12625,N_12826);
and U12912 (N_12912,N_12878,N_12827);
nor U12913 (N_12913,N_12695,N_12730);
and U12914 (N_12914,N_12719,N_12890);
or U12915 (N_12915,N_12757,N_12683);
or U12916 (N_12916,N_12887,N_12748);
nand U12917 (N_12917,N_12862,N_12843);
or U12918 (N_12918,N_12655,N_12718);
and U12919 (N_12919,N_12877,N_12837);
xnor U12920 (N_12920,N_12651,N_12638);
and U12921 (N_12921,N_12674,N_12832);
nor U12922 (N_12922,N_12770,N_12640);
nand U12923 (N_12923,N_12735,N_12654);
nand U12924 (N_12924,N_12687,N_12737);
xor U12925 (N_12925,N_12834,N_12622);
or U12926 (N_12926,N_12681,N_12786);
nand U12927 (N_12927,N_12699,N_12792);
and U12928 (N_12928,N_12742,N_12873);
xor U12929 (N_12929,N_12715,N_12891);
xnor U12930 (N_12930,N_12639,N_12870);
nor U12931 (N_12931,N_12635,N_12644);
and U12932 (N_12932,N_12805,N_12628);
and U12933 (N_12933,N_12807,N_12614);
nand U12934 (N_12934,N_12835,N_12813);
or U12935 (N_12935,N_12793,N_12896);
nor U12936 (N_12936,N_12766,N_12860);
nand U12937 (N_12937,N_12636,N_12866);
and U12938 (N_12938,N_12684,N_12712);
nor U12939 (N_12939,N_12814,N_12739);
nand U12940 (N_12940,N_12812,N_12892);
xor U12941 (N_12941,N_12851,N_12672);
nand U12942 (N_12942,N_12776,N_12705);
and U12943 (N_12943,N_12772,N_12693);
or U12944 (N_12944,N_12852,N_12652);
nor U12945 (N_12945,N_12609,N_12624);
xnor U12946 (N_12946,N_12875,N_12889);
xnor U12947 (N_12947,N_12759,N_12617);
nor U12948 (N_12948,N_12662,N_12673);
or U12949 (N_12949,N_12897,N_12898);
nand U12950 (N_12950,N_12736,N_12857);
nand U12951 (N_12951,N_12721,N_12820);
xnor U12952 (N_12952,N_12818,N_12893);
nor U12953 (N_12953,N_12782,N_12828);
xnor U12954 (N_12954,N_12605,N_12738);
and U12955 (N_12955,N_12823,N_12854);
nor U12956 (N_12956,N_12803,N_12637);
xnor U12957 (N_12957,N_12732,N_12894);
or U12958 (N_12958,N_12841,N_12795);
xnor U12959 (N_12959,N_12885,N_12765);
and U12960 (N_12960,N_12751,N_12899);
xnor U12961 (N_12961,N_12879,N_12615);
or U12962 (N_12962,N_12755,N_12709);
xor U12963 (N_12963,N_12847,N_12733);
or U12964 (N_12964,N_12831,N_12849);
xnor U12965 (N_12965,N_12608,N_12711);
nor U12966 (N_12966,N_12799,N_12886);
or U12967 (N_12967,N_12881,N_12858);
nand U12968 (N_12968,N_12783,N_12788);
nand U12969 (N_12969,N_12830,N_12773);
xor U12970 (N_12970,N_12645,N_12717);
or U12971 (N_12971,N_12657,N_12884);
and U12972 (N_12972,N_12630,N_12665);
nor U12973 (N_12973,N_12871,N_12669);
or U12974 (N_12974,N_12679,N_12760);
xor U12975 (N_12975,N_12747,N_12840);
or U12976 (N_12976,N_12731,N_12667);
or U12977 (N_12977,N_12714,N_12789);
and U12978 (N_12978,N_12701,N_12725);
xnor U12979 (N_12979,N_12685,N_12698);
or U12980 (N_12980,N_12728,N_12631);
nor U12981 (N_12981,N_12829,N_12680);
xor U12982 (N_12982,N_12727,N_12646);
or U12983 (N_12983,N_12817,N_12845);
or U12984 (N_12984,N_12692,N_12762);
and U12985 (N_12985,N_12797,N_12846);
nor U12986 (N_12986,N_12769,N_12650);
xor U12987 (N_12987,N_12686,N_12867);
nand U12988 (N_12988,N_12602,N_12864);
nand U12989 (N_12989,N_12855,N_12798);
or U12990 (N_12990,N_12777,N_12743);
nand U12991 (N_12991,N_12821,N_12729);
or U12992 (N_12992,N_12791,N_12740);
nand U12993 (N_12993,N_12675,N_12648);
xnor U12994 (N_12994,N_12724,N_12666);
nor U12995 (N_12995,N_12613,N_12611);
and U12996 (N_12996,N_12643,N_12874);
nand U12997 (N_12997,N_12656,N_12787);
and U12998 (N_12998,N_12706,N_12663);
xor U12999 (N_12999,N_12612,N_12811);
nand U13000 (N_13000,N_12670,N_12802);
nand U13001 (N_13001,N_12688,N_12745);
nor U13002 (N_13002,N_12775,N_12690);
and U13003 (N_13003,N_12647,N_12618);
and U13004 (N_13004,N_12689,N_12801);
nor U13005 (N_13005,N_12761,N_12861);
nand U13006 (N_13006,N_12649,N_12865);
and U13007 (N_13007,N_12754,N_12658);
or U13008 (N_13008,N_12704,N_12691);
nor U13009 (N_13009,N_12784,N_12809);
nor U13010 (N_13010,N_12707,N_12619);
nor U13011 (N_13011,N_12842,N_12816);
xor U13012 (N_13012,N_12627,N_12876);
nand U13013 (N_13013,N_12856,N_12682);
and U13014 (N_13014,N_12642,N_12882);
or U13015 (N_13015,N_12744,N_12779);
xor U13016 (N_13016,N_12603,N_12700);
nand U13017 (N_13017,N_12697,N_12632);
xor U13018 (N_13018,N_12781,N_12749);
xor U13019 (N_13019,N_12872,N_12696);
nor U13020 (N_13020,N_12824,N_12853);
nor U13021 (N_13021,N_12804,N_12653);
nand U13022 (N_13022,N_12780,N_12796);
nor U13023 (N_13023,N_12785,N_12800);
xor U13024 (N_13024,N_12678,N_12610);
nor U13025 (N_13025,N_12659,N_12756);
or U13026 (N_13026,N_12778,N_12620);
xor U13027 (N_13027,N_12713,N_12825);
nand U13028 (N_13028,N_12600,N_12623);
nor U13029 (N_13029,N_12607,N_12671);
or U13030 (N_13030,N_12621,N_12752);
nand U13031 (N_13031,N_12641,N_12774);
or U13032 (N_13032,N_12661,N_12888);
or U13033 (N_13033,N_12694,N_12716);
and U13034 (N_13034,N_12819,N_12629);
and U13035 (N_13035,N_12822,N_12722);
and U13036 (N_13036,N_12616,N_12601);
nor U13037 (N_13037,N_12848,N_12708);
or U13038 (N_13038,N_12806,N_12746);
nand U13039 (N_13039,N_12794,N_12833);
and U13040 (N_13040,N_12626,N_12723);
xor U13041 (N_13041,N_12768,N_12863);
and U13042 (N_13042,N_12660,N_12859);
xor U13043 (N_13043,N_12869,N_12633);
nand U13044 (N_13044,N_12753,N_12710);
xnor U13045 (N_13045,N_12764,N_12880);
xnor U13046 (N_13046,N_12720,N_12850);
nand U13047 (N_13047,N_12790,N_12838);
nor U13048 (N_13048,N_12726,N_12703);
or U13049 (N_13049,N_12668,N_12836);
or U13050 (N_13050,N_12829,N_12840);
nand U13051 (N_13051,N_12832,N_12689);
nand U13052 (N_13052,N_12613,N_12892);
xnor U13053 (N_13053,N_12717,N_12780);
nand U13054 (N_13054,N_12761,N_12664);
or U13055 (N_13055,N_12871,N_12891);
xor U13056 (N_13056,N_12801,N_12819);
nand U13057 (N_13057,N_12851,N_12626);
or U13058 (N_13058,N_12723,N_12770);
nor U13059 (N_13059,N_12683,N_12833);
nand U13060 (N_13060,N_12891,N_12625);
nor U13061 (N_13061,N_12785,N_12741);
and U13062 (N_13062,N_12888,N_12653);
xnor U13063 (N_13063,N_12865,N_12682);
xor U13064 (N_13064,N_12705,N_12806);
and U13065 (N_13065,N_12787,N_12799);
xor U13066 (N_13066,N_12753,N_12749);
nor U13067 (N_13067,N_12732,N_12812);
or U13068 (N_13068,N_12814,N_12721);
nand U13069 (N_13069,N_12644,N_12674);
or U13070 (N_13070,N_12753,N_12662);
and U13071 (N_13071,N_12765,N_12650);
nor U13072 (N_13072,N_12885,N_12619);
nand U13073 (N_13073,N_12789,N_12837);
xor U13074 (N_13074,N_12733,N_12625);
and U13075 (N_13075,N_12842,N_12673);
nor U13076 (N_13076,N_12666,N_12628);
or U13077 (N_13077,N_12842,N_12603);
and U13078 (N_13078,N_12755,N_12607);
nand U13079 (N_13079,N_12604,N_12804);
xor U13080 (N_13080,N_12708,N_12723);
nor U13081 (N_13081,N_12726,N_12780);
and U13082 (N_13082,N_12677,N_12640);
or U13083 (N_13083,N_12717,N_12653);
nand U13084 (N_13084,N_12751,N_12605);
or U13085 (N_13085,N_12896,N_12691);
nand U13086 (N_13086,N_12682,N_12840);
nor U13087 (N_13087,N_12855,N_12864);
and U13088 (N_13088,N_12762,N_12760);
nor U13089 (N_13089,N_12647,N_12761);
xnor U13090 (N_13090,N_12626,N_12771);
nor U13091 (N_13091,N_12841,N_12826);
or U13092 (N_13092,N_12781,N_12802);
xnor U13093 (N_13093,N_12733,N_12679);
and U13094 (N_13094,N_12756,N_12794);
nor U13095 (N_13095,N_12821,N_12662);
nand U13096 (N_13096,N_12847,N_12827);
nand U13097 (N_13097,N_12888,N_12890);
or U13098 (N_13098,N_12898,N_12835);
xnor U13099 (N_13099,N_12694,N_12603);
and U13100 (N_13100,N_12695,N_12622);
nor U13101 (N_13101,N_12763,N_12684);
and U13102 (N_13102,N_12800,N_12624);
or U13103 (N_13103,N_12845,N_12848);
xnor U13104 (N_13104,N_12671,N_12674);
or U13105 (N_13105,N_12614,N_12659);
or U13106 (N_13106,N_12763,N_12841);
nor U13107 (N_13107,N_12876,N_12863);
nor U13108 (N_13108,N_12603,N_12887);
or U13109 (N_13109,N_12631,N_12833);
or U13110 (N_13110,N_12786,N_12853);
xnor U13111 (N_13111,N_12628,N_12643);
nor U13112 (N_13112,N_12892,N_12618);
and U13113 (N_13113,N_12658,N_12872);
xor U13114 (N_13114,N_12700,N_12655);
and U13115 (N_13115,N_12845,N_12766);
nand U13116 (N_13116,N_12676,N_12629);
and U13117 (N_13117,N_12834,N_12647);
xor U13118 (N_13118,N_12735,N_12844);
and U13119 (N_13119,N_12784,N_12695);
nand U13120 (N_13120,N_12684,N_12893);
nor U13121 (N_13121,N_12643,N_12641);
xnor U13122 (N_13122,N_12607,N_12650);
or U13123 (N_13123,N_12615,N_12792);
and U13124 (N_13124,N_12830,N_12840);
nand U13125 (N_13125,N_12646,N_12821);
nor U13126 (N_13126,N_12740,N_12674);
nand U13127 (N_13127,N_12757,N_12660);
or U13128 (N_13128,N_12722,N_12687);
xor U13129 (N_13129,N_12899,N_12698);
xnor U13130 (N_13130,N_12649,N_12860);
nand U13131 (N_13131,N_12890,N_12617);
nor U13132 (N_13132,N_12721,N_12770);
nand U13133 (N_13133,N_12796,N_12790);
xnor U13134 (N_13134,N_12848,N_12800);
and U13135 (N_13135,N_12803,N_12619);
nor U13136 (N_13136,N_12843,N_12616);
or U13137 (N_13137,N_12705,N_12652);
nand U13138 (N_13138,N_12740,N_12783);
nand U13139 (N_13139,N_12794,N_12777);
or U13140 (N_13140,N_12684,N_12771);
xor U13141 (N_13141,N_12725,N_12871);
or U13142 (N_13142,N_12735,N_12838);
and U13143 (N_13143,N_12665,N_12685);
and U13144 (N_13144,N_12712,N_12656);
and U13145 (N_13145,N_12823,N_12646);
nand U13146 (N_13146,N_12882,N_12705);
nor U13147 (N_13147,N_12793,N_12622);
or U13148 (N_13148,N_12892,N_12667);
xnor U13149 (N_13149,N_12782,N_12834);
and U13150 (N_13150,N_12773,N_12860);
xnor U13151 (N_13151,N_12860,N_12737);
nor U13152 (N_13152,N_12782,N_12826);
or U13153 (N_13153,N_12627,N_12607);
nand U13154 (N_13154,N_12665,N_12731);
nand U13155 (N_13155,N_12609,N_12629);
and U13156 (N_13156,N_12802,N_12849);
or U13157 (N_13157,N_12845,N_12687);
xnor U13158 (N_13158,N_12894,N_12836);
nor U13159 (N_13159,N_12794,N_12868);
or U13160 (N_13160,N_12808,N_12749);
xnor U13161 (N_13161,N_12777,N_12671);
and U13162 (N_13162,N_12653,N_12845);
and U13163 (N_13163,N_12649,N_12844);
and U13164 (N_13164,N_12719,N_12837);
xor U13165 (N_13165,N_12830,N_12831);
nor U13166 (N_13166,N_12777,N_12773);
nand U13167 (N_13167,N_12643,N_12801);
and U13168 (N_13168,N_12738,N_12891);
and U13169 (N_13169,N_12713,N_12758);
xor U13170 (N_13170,N_12648,N_12680);
and U13171 (N_13171,N_12674,N_12845);
nor U13172 (N_13172,N_12603,N_12831);
nand U13173 (N_13173,N_12807,N_12824);
xnor U13174 (N_13174,N_12775,N_12785);
xor U13175 (N_13175,N_12678,N_12853);
nand U13176 (N_13176,N_12849,N_12755);
nor U13177 (N_13177,N_12796,N_12838);
and U13178 (N_13178,N_12763,N_12752);
and U13179 (N_13179,N_12817,N_12735);
xor U13180 (N_13180,N_12615,N_12818);
nor U13181 (N_13181,N_12660,N_12635);
nand U13182 (N_13182,N_12833,N_12734);
nand U13183 (N_13183,N_12688,N_12687);
xnor U13184 (N_13184,N_12820,N_12699);
or U13185 (N_13185,N_12776,N_12701);
and U13186 (N_13186,N_12650,N_12696);
nor U13187 (N_13187,N_12651,N_12893);
nor U13188 (N_13188,N_12855,N_12677);
xnor U13189 (N_13189,N_12879,N_12799);
nor U13190 (N_13190,N_12866,N_12600);
or U13191 (N_13191,N_12831,N_12696);
nand U13192 (N_13192,N_12678,N_12601);
xor U13193 (N_13193,N_12771,N_12601);
and U13194 (N_13194,N_12821,N_12701);
or U13195 (N_13195,N_12831,N_12882);
or U13196 (N_13196,N_12692,N_12821);
nand U13197 (N_13197,N_12782,N_12680);
nor U13198 (N_13198,N_12762,N_12844);
xnor U13199 (N_13199,N_12886,N_12887);
or U13200 (N_13200,N_13115,N_12977);
nand U13201 (N_13201,N_13157,N_12968);
nand U13202 (N_13202,N_12998,N_12909);
or U13203 (N_13203,N_12984,N_13196);
nor U13204 (N_13204,N_13160,N_12925);
and U13205 (N_13205,N_13088,N_13132);
and U13206 (N_13206,N_13097,N_13043);
and U13207 (N_13207,N_12985,N_13144);
xnor U13208 (N_13208,N_13016,N_13029);
or U13209 (N_13209,N_12976,N_13106);
xor U13210 (N_13210,N_13104,N_12945);
and U13211 (N_13211,N_13102,N_13165);
nand U13212 (N_13212,N_13071,N_13151);
xor U13213 (N_13213,N_13079,N_13128);
nor U13214 (N_13214,N_13078,N_13024);
and U13215 (N_13215,N_13152,N_13061);
or U13216 (N_13216,N_12927,N_13176);
or U13217 (N_13217,N_13073,N_12922);
nor U13218 (N_13218,N_13085,N_12926);
or U13219 (N_13219,N_13008,N_13181);
nand U13220 (N_13220,N_12939,N_13080);
and U13221 (N_13221,N_13040,N_13191);
and U13222 (N_13222,N_13118,N_13103);
and U13223 (N_13223,N_13095,N_12983);
and U13224 (N_13224,N_12938,N_12914);
and U13225 (N_13225,N_12924,N_13094);
xor U13226 (N_13226,N_12917,N_12932);
nand U13227 (N_13227,N_13048,N_13018);
and U13228 (N_13228,N_13058,N_13142);
nand U13229 (N_13229,N_12934,N_12996);
xor U13230 (N_13230,N_13098,N_13154);
and U13231 (N_13231,N_13017,N_13036);
nor U13232 (N_13232,N_13039,N_13133);
nor U13233 (N_13233,N_12979,N_13167);
xnor U13234 (N_13234,N_13141,N_13113);
or U13235 (N_13235,N_13198,N_13112);
xnor U13236 (N_13236,N_12966,N_13170);
or U13237 (N_13237,N_12967,N_12929);
nor U13238 (N_13238,N_13188,N_13059);
nor U13239 (N_13239,N_13091,N_13035);
nand U13240 (N_13240,N_13013,N_13052);
nand U13241 (N_13241,N_13114,N_12959);
xor U13242 (N_13242,N_12990,N_13003);
nor U13243 (N_13243,N_13044,N_12915);
and U13244 (N_13244,N_12957,N_13068);
or U13245 (N_13245,N_13140,N_12908);
nand U13246 (N_13246,N_12992,N_13183);
or U13247 (N_13247,N_13143,N_13051);
xor U13248 (N_13248,N_13014,N_12961);
and U13249 (N_13249,N_13186,N_13137);
xnor U13250 (N_13250,N_12958,N_13185);
and U13251 (N_13251,N_13010,N_12988);
nor U13252 (N_13252,N_12950,N_13194);
and U13253 (N_13253,N_13006,N_12964);
or U13254 (N_13254,N_12991,N_12952);
nand U13255 (N_13255,N_13177,N_13193);
or U13256 (N_13256,N_13020,N_13138);
nand U13257 (N_13257,N_12910,N_13145);
or U13258 (N_13258,N_13045,N_13129);
xnor U13259 (N_13259,N_13049,N_13082);
xnor U13260 (N_13260,N_12993,N_13083);
xor U13261 (N_13261,N_13108,N_12982);
and U13262 (N_13262,N_13002,N_12975);
and U13263 (N_13263,N_13107,N_13175);
nand U13264 (N_13264,N_13099,N_13166);
and U13265 (N_13265,N_13077,N_13011);
and U13266 (N_13266,N_13069,N_13093);
xnor U13267 (N_13267,N_13120,N_13111);
and U13268 (N_13268,N_13123,N_13060);
or U13269 (N_13269,N_13007,N_13197);
nand U13270 (N_13270,N_12974,N_13171);
xor U13271 (N_13271,N_13047,N_12916);
and U13272 (N_13272,N_13053,N_12956);
and U13273 (N_13273,N_12944,N_13086);
nand U13274 (N_13274,N_13195,N_13130);
or U13275 (N_13275,N_13055,N_13146);
nand U13276 (N_13276,N_13122,N_13127);
nand U13277 (N_13277,N_12971,N_13169);
nand U13278 (N_13278,N_12965,N_13147);
and U13279 (N_13279,N_13156,N_12943);
or U13280 (N_13280,N_13066,N_12987);
xnor U13281 (N_13281,N_12940,N_13182);
nor U13282 (N_13282,N_13134,N_13121);
xnor U13283 (N_13283,N_12913,N_13090);
nor U13284 (N_13284,N_13075,N_13004);
nor U13285 (N_13285,N_12907,N_13050);
xor U13286 (N_13286,N_12921,N_12994);
nand U13287 (N_13287,N_13153,N_13084);
xor U13288 (N_13288,N_13119,N_13030);
xor U13289 (N_13289,N_13189,N_12960);
nor U13290 (N_13290,N_13125,N_12933);
and U13291 (N_13291,N_13184,N_12936);
and U13292 (N_13292,N_13056,N_13089);
nor U13293 (N_13293,N_13131,N_13032);
nor U13294 (N_13294,N_12912,N_13038);
and U13295 (N_13295,N_13064,N_13046);
nand U13296 (N_13296,N_12973,N_13022);
nor U13297 (N_13297,N_13174,N_13101);
nor U13298 (N_13298,N_13162,N_12948);
and U13299 (N_13299,N_12949,N_12920);
xor U13300 (N_13300,N_12995,N_12904);
xnor U13301 (N_13301,N_12947,N_13117);
nor U13302 (N_13302,N_13173,N_12986);
xor U13303 (N_13303,N_12906,N_13023);
or U13304 (N_13304,N_13081,N_13179);
and U13305 (N_13305,N_13105,N_13092);
nand U13306 (N_13306,N_12905,N_13062);
nand U13307 (N_13307,N_12963,N_13057);
nand U13308 (N_13308,N_13042,N_13116);
nor U13309 (N_13309,N_12942,N_13087);
or U13310 (N_13310,N_13109,N_13168);
or U13311 (N_13311,N_13031,N_13028);
nand U13312 (N_13312,N_13012,N_12946);
and U13313 (N_13313,N_13158,N_13126);
and U13314 (N_13314,N_13074,N_13001);
xor U13315 (N_13315,N_13159,N_12918);
xnor U13316 (N_13316,N_13025,N_13065);
and U13317 (N_13317,N_13190,N_12941);
or U13318 (N_13318,N_12980,N_13192);
nor U13319 (N_13319,N_12937,N_12972);
and U13320 (N_13320,N_12969,N_12951);
or U13321 (N_13321,N_13135,N_12970);
or U13322 (N_13322,N_13005,N_13139);
or U13323 (N_13323,N_13199,N_12978);
or U13324 (N_13324,N_12928,N_13019);
and U13325 (N_13325,N_13033,N_13072);
xnor U13326 (N_13326,N_12900,N_13124);
or U13327 (N_13327,N_13009,N_13096);
nand U13328 (N_13328,N_12981,N_13150);
xor U13329 (N_13329,N_12911,N_13155);
nor U13330 (N_13330,N_13172,N_13187);
nor U13331 (N_13331,N_13148,N_12930);
and U13332 (N_13332,N_13161,N_13026);
nand U13333 (N_13333,N_12919,N_13178);
and U13334 (N_13334,N_13027,N_13067);
xnor U13335 (N_13335,N_12962,N_13076);
xor U13336 (N_13336,N_13021,N_13034);
or U13337 (N_13337,N_12903,N_13180);
xnor U13338 (N_13338,N_12955,N_13164);
nand U13339 (N_13339,N_13163,N_13100);
and U13340 (N_13340,N_13136,N_12931);
nand U13341 (N_13341,N_13054,N_13070);
xor U13342 (N_13342,N_12902,N_13149);
or U13343 (N_13343,N_12901,N_13110);
or U13344 (N_13344,N_12989,N_12953);
and U13345 (N_13345,N_13041,N_12923);
nor U13346 (N_13346,N_12935,N_13015);
nand U13347 (N_13347,N_13000,N_12999);
nor U13348 (N_13348,N_12997,N_12954);
and U13349 (N_13349,N_13037,N_13063);
nor U13350 (N_13350,N_12976,N_12931);
xor U13351 (N_13351,N_13181,N_13082);
nand U13352 (N_13352,N_12933,N_13101);
nand U13353 (N_13353,N_12971,N_13174);
or U13354 (N_13354,N_12982,N_13192);
nand U13355 (N_13355,N_13109,N_13079);
or U13356 (N_13356,N_12987,N_12957);
or U13357 (N_13357,N_12947,N_12989);
nor U13358 (N_13358,N_13051,N_13000);
xor U13359 (N_13359,N_13123,N_13190);
xnor U13360 (N_13360,N_13179,N_13033);
and U13361 (N_13361,N_13188,N_13100);
nor U13362 (N_13362,N_13090,N_13093);
nand U13363 (N_13363,N_13001,N_12926);
xor U13364 (N_13364,N_13109,N_13162);
and U13365 (N_13365,N_13105,N_13115);
nor U13366 (N_13366,N_12947,N_12942);
xor U13367 (N_13367,N_13078,N_13094);
or U13368 (N_13368,N_13059,N_13083);
or U13369 (N_13369,N_13085,N_13024);
nor U13370 (N_13370,N_12974,N_13164);
xor U13371 (N_13371,N_13149,N_12966);
and U13372 (N_13372,N_13185,N_13099);
and U13373 (N_13373,N_13193,N_12907);
and U13374 (N_13374,N_13109,N_12952);
nor U13375 (N_13375,N_13180,N_12950);
nand U13376 (N_13376,N_12936,N_12932);
nor U13377 (N_13377,N_13079,N_12938);
nand U13378 (N_13378,N_13166,N_13028);
and U13379 (N_13379,N_13030,N_13078);
nand U13380 (N_13380,N_13171,N_13154);
or U13381 (N_13381,N_13187,N_12950);
and U13382 (N_13382,N_13125,N_13176);
nand U13383 (N_13383,N_12999,N_13101);
nand U13384 (N_13384,N_12986,N_13143);
nor U13385 (N_13385,N_13044,N_12913);
and U13386 (N_13386,N_13161,N_13031);
nor U13387 (N_13387,N_12916,N_12967);
or U13388 (N_13388,N_13163,N_12921);
and U13389 (N_13389,N_13174,N_13084);
nor U13390 (N_13390,N_12931,N_13059);
nand U13391 (N_13391,N_13137,N_13144);
xnor U13392 (N_13392,N_13071,N_12951);
xor U13393 (N_13393,N_12905,N_13171);
and U13394 (N_13394,N_12954,N_13132);
and U13395 (N_13395,N_13066,N_13184);
and U13396 (N_13396,N_12968,N_13015);
xor U13397 (N_13397,N_12977,N_12980);
and U13398 (N_13398,N_13036,N_12976);
xnor U13399 (N_13399,N_13001,N_13014);
and U13400 (N_13400,N_12952,N_12989);
nor U13401 (N_13401,N_13185,N_12952);
nor U13402 (N_13402,N_13083,N_12927);
nor U13403 (N_13403,N_13124,N_13159);
or U13404 (N_13404,N_13043,N_13120);
and U13405 (N_13405,N_13160,N_12953);
nand U13406 (N_13406,N_12916,N_13000);
or U13407 (N_13407,N_13132,N_13145);
and U13408 (N_13408,N_13047,N_12980);
nand U13409 (N_13409,N_13039,N_13008);
and U13410 (N_13410,N_12912,N_13071);
and U13411 (N_13411,N_13179,N_13171);
or U13412 (N_13412,N_12919,N_13049);
xor U13413 (N_13413,N_13022,N_13054);
and U13414 (N_13414,N_12962,N_12912);
nor U13415 (N_13415,N_13176,N_13050);
or U13416 (N_13416,N_13101,N_13065);
and U13417 (N_13417,N_12906,N_13058);
nand U13418 (N_13418,N_12914,N_12940);
and U13419 (N_13419,N_13191,N_12915);
nor U13420 (N_13420,N_13050,N_13177);
xnor U13421 (N_13421,N_13169,N_12938);
xor U13422 (N_13422,N_13160,N_13058);
nor U13423 (N_13423,N_12982,N_13006);
xor U13424 (N_13424,N_13193,N_13143);
or U13425 (N_13425,N_13141,N_13019);
and U13426 (N_13426,N_12986,N_13149);
nand U13427 (N_13427,N_13099,N_13123);
nand U13428 (N_13428,N_13007,N_13103);
nor U13429 (N_13429,N_13092,N_12931);
xor U13430 (N_13430,N_13080,N_12955);
and U13431 (N_13431,N_13058,N_12909);
nand U13432 (N_13432,N_13143,N_13039);
xor U13433 (N_13433,N_12954,N_13068);
nor U13434 (N_13434,N_12974,N_13119);
and U13435 (N_13435,N_13164,N_13049);
or U13436 (N_13436,N_13098,N_13120);
and U13437 (N_13437,N_12954,N_13131);
or U13438 (N_13438,N_13041,N_12971);
and U13439 (N_13439,N_12918,N_12980);
nor U13440 (N_13440,N_13151,N_13070);
and U13441 (N_13441,N_13002,N_13007);
nand U13442 (N_13442,N_12995,N_13044);
nand U13443 (N_13443,N_13085,N_13071);
or U13444 (N_13444,N_13039,N_12905);
xor U13445 (N_13445,N_13153,N_13106);
or U13446 (N_13446,N_13193,N_13008);
xor U13447 (N_13447,N_12932,N_13007);
or U13448 (N_13448,N_13099,N_12908);
nor U13449 (N_13449,N_12907,N_13027);
and U13450 (N_13450,N_13002,N_13031);
nand U13451 (N_13451,N_13030,N_12931);
and U13452 (N_13452,N_12922,N_13008);
or U13453 (N_13453,N_12964,N_12950);
or U13454 (N_13454,N_13168,N_13113);
or U13455 (N_13455,N_13111,N_13094);
nand U13456 (N_13456,N_12988,N_13118);
xnor U13457 (N_13457,N_13117,N_13069);
nor U13458 (N_13458,N_13150,N_12998);
nor U13459 (N_13459,N_13157,N_13006);
or U13460 (N_13460,N_12943,N_13059);
or U13461 (N_13461,N_12909,N_13083);
and U13462 (N_13462,N_12972,N_13193);
nor U13463 (N_13463,N_13028,N_12919);
nor U13464 (N_13464,N_13074,N_13030);
nand U13465 (N_13465,N_13199,N_13153);
or U13466 (N_13466,N_12938,N_13070);
xnor U13467 (N_13467,N_12985,N_13078);
nand U13468 (N_13468,N_13010,N_13075);
nor U13469 (N_13469,N_13129,N_12962);
and U13470 (N_13470,N_13182,N_13168);
xor U13471 (N_13471,N_12950,N_12919);
and U13472 (N_13472,N_13153,N_13177);
xor U13473 (N_13473,N_12938,N_13194);
and U13474 (N_13474,N_12943,N_13128);
nor U13475 (N_13475,N_13001,N_13067);
nor U13476 (N_13476,N_13050,N_12911);
nor U13477 (N_13477,N_12985,N_13159);
and U13478 (N_13478,N_12966,N_12963);
nand U13479 (N_13479,N_13082,N_12912);
xnor U13480 (N_13480,N_13111,N_13096);
nor U13481 (N_13481,N_13015,N_13130);
nor U13482 (N_13482,N_13119,N_12938);
xor U13483 (N_13483,N_13123,N_13026);
nand U13484 (N_13484,N_12982,N_13157);
xnor U13485 (N_13485,N_13036,N_12988);
or U13486 (N_13486,N_12987,N_12941);
and U13487 (N_13487,N_13170,N_13196);
nand U13488 (N_13488,N_12921,N_13015);
nor U13489 (N_13489,N_13084,N_13184);
xnor U13490 (N_13490,N_13122,N_13076);
xnor U13491 (N_13491,N_12989,N_13084);
or U13492 (N_13492,N_13085,N_13033);
xor U13493 (N_13493,N_12950,N_13016);
and U13494 (N_13494,N_13053,N_13014);
nand U13495 (N_13495,N_13180,N_13015);
xor U13496 (N_13496,N_13136,N_13100);
xor U13497 (N_13497,N_13002,N_12933);
and U13498 (N_13498,N_13056,N_13035);
and U13499 (N_13499,N_12926,N_12962);
and U13500 (N_13500,N_13491,N_13466);
and U13501 (N_13501,N_13394,N_13340);
and U13502 (N_13502,N_13276,N_13312);
or U13503 (N_13503,N_13332,N_13495);
and U13504 (N_13504,N_13341,N_13271);
nor U13505 (N_13505,N_13446,N_13259);
nand U13506 (N_13506,N_13263,N_13286);
nand U13507 (N_13507,N_13464,N_13447);
nor U13508 (N_13508,N_13435,N_13236);
and U13509 (N_13509,N_13377,N_13265);
xor U13510 (N_13510,N_13389,N_13357);
xnor U13511 (N_13511,N_13454,N_13399);
or U13512 (N_13512,N_13224,N_13436);
nand U13513 (N_13513,N_13392,N_13362);
nand U13514 (N_13514,N_13343,N_13477);
nor U13515 (N_13515,N_13405,N_13244);
nand U13516 (N_13516,N_13470,N_13300);
and U13517 (N_13517,N_13327,N_13472);
xor U13518 (N_13518,N_13234,N_13202);
nor U13519 (N_13519,N_13274,N_13431);
nor U13520 (N_13520,N_13251,N_13297);
and U13521 (N_13521,N_13277,N_13320);
nand U13522 (N_13522,N_13324,N_13359);
or U13523 (N_13523,N_13473,N_13413);
nand U13524 (N_13524,N_13424,N_13308);
xor U13525 (N_13525,N_13273,N_13299);
nand U13526 (N_13526,N_13368,N_13289);
nand U13527 (N_13527,N_13246,N_13262);
or U13528 (N_13528,N_13203,N_13385);
nand U13529 (N_13529,N_13328,N_13344);
xor U13530 (N_13530,N_13498,N_13449);
and U13531 (N_13531,N_13302,N_13411);
nor U13532 (N_13532,N_13426,N_13205);
xnor U13533 (N_13533,N_13369,N_13442);
nor U13534 (N_13534,N_13418,N_13230);
nor U13535 (N_13535,N_13420,N_13462);
or U13536 (N_13536,N_13363,N_13346);
or U13537 (N_13537,N_13206,N_13295);
nor U13538 (N_13538,N_13417,N_13459);
and U13539 (N_13539,N_13401,N_13255);
xnor U13540 (N_13540,N_13314,N_13358);
or U13541 (N_13541,N_13301,N_13348);
nand U13542 (N_13542,N_13266,N_13267);
nand U13543 (N_13543,N_13400,N_13335);
nor U13544 (N_13544,N_13425,N_13269);
and U13545 (N_13545,N_13317,N_13445);
nand U13546 (N_13546,N_13298,N_13351);
nand U13547 (N_13547,N_13311,N_13256);
nor U13548 (N_13548,N_13408,N_13252);
or U13549 (N_13549,N_13290,N_13370);
nand U13550 (N_13550,N_13235,N_13434);
and U13551 (N_13551,N_13282,N_13221);
xnor U13552 (N_13552,N_13333,N_13427);
or U13553 (N_13553,N_13430,N_13478);
nand U13554 (N_13554,N_13339,N_13275);
and U13555 (N_13555,N_13248,N_13390);
nand U13556 (N_13556,N_13443,N_13467);
xnor U13557 (N_13557,N_13294,N_13291);
and U13558 (N_13558,N_13437,N_13219);
xnor U13559 (N_13559,N_13372,N_13450);
nor U13560 (N_13560,N_13229,N_13485);
xnor U13561 (N_13561,N_13233,N_13260);
nor U13562 (N_13562,N_13376,N_13241);
xor U13563 (N_13563,N_13322,N_13240);
nand U13564 (N_13564,N_13326,N_13371);
and U13565 (N_13565,N_13220,N_13336);
or U13566 (N_13566,N_13393,N_13432);
xnor U13567 (N_13567,N_13379,N_13404);
xor U13568 (N_13568,N_13249,N_13475);
nand U13569 (N_13569,N_13448,N_13319);
xor U13570 (N_13570,N_13486,N_13208);
nand U13571 (N_13571,N_13451,N_13396);
nand U13572 (N_13572,N_13409,N_13497);
nand U13573 (N_13573,N_13288,N_13216);
xnor U13574 (N_13574,N_13223,N_13360);
nand U13575 (N_13575,N_13496,N_13334);
nor U13576 (N_13576,N_13460,N_13330);
and U13577 (N_13577,N_13323,N_13452);
or U13578 (N_13578,N_13225,N_13471);
nand U13579 (N_13579,N_13321,N_13361);
or U13580 (N_13580,N_13428,N_13226);
or U13581 (N_13581,N_13272,N_13488);
xnor U13582 (N_13582,N_13227,N_13374);
xnor U13583 (N_13583,N_13398,N_13479);
xnor U13584 (N_13584,N_13438,N_13316);
nand U13585 (N_13585,N_13354,N_13421);
nor U13586 (N_13586,N_13211,N_13453);
nand U13587 (N_13587,N_13373,N_13474);
nand U13588 (N_13588,N_13490,N_13352);
nand U13589 (N_13589,N_13313,N_13456);
nor U13590 (N_13590,N_13366,N_13455);
and U13591 (N_13591,N_13440,N_13414);
nor U13592 (N_13592,N_13304,N_13231);
nand U13593 (N_13593,N_13461,N_13315);
xor U13594 (N_13594,N_13342,N_13247);
and U13595 (N_13595,N_13481,N_13367);
or U13596 (N_13596,N_13381,N_13364);
and U13597 (N_13597,N_13469,N_13388);
and U13598 (N_13598,N_13303,N_13292);
nor U13599 (N_13599,N_13412,N_13283);
xnor U13600 (N_13600,N_13356,N_13329);
or U13601 (N_13601,N_13204,N_13207);
nor U13602 (N_13602,N_13402,N_13476);
nor U13603 (N_13603,N_13457,N_13391);
xnor U13604 (N_13604,N_13397,N_13383);
nor U13605 (N_13605,N_13243,N_13242);
and U13606 (N_13606,N_13492,N_13213);
or U13607 (N_13607,N_13380,N_13296);
nor U13608 (N_13608,N_13209,N_13258);
nand U13609 (N_13609,N_13279,N_13254);
and U13610 (N_13610,N_13250,N_13386);
nor U13611 (N_13611,N_13423,N_13214);
xor U13612 (N_13612,N_13284,N_13419);
nand U13613 (N_13613,N_13465,N_13444);
xor U13614 (N_13614,N_13433,N_13422);
xnor U13615 (N_13615,N_13309,N_13499);
and U13616 (N_13616,N_13487,N_13305);
or U13617 (N_13617,N_13349,N_13350);
nor U13618 (N_13618,N_13280,N_13384);
nand U13619 (N_13619,N_13382,N_13238);
nor U13620 (N_13620,N_13337,N_13318);
nand U13621 (N_13621,N_13458,N_13468);
nand U13622 (N_13622,N_13403,N_13257);
nor U13623 (N_13623,N_13201,N_13217);
nor U13624 (N_13624,N_13375,N_13228);
nor U13625 (N_13625,N_13489,N_13463);
and U13626 (N_13626,N_13493,N_13239);
and U13627 (N_13627,N_13484,N_13415);
xnor U13628 (N_13628,N_13325,N_13215);
or U13629 (N_13629,N_13441,N_13338);
xnor U13630 (N_13630,N_13261,N_13416);
nand U13631 (N_13631,N_13483,N_13218);
nand U13632 (N_13632,N_13307,N_13245);
or U13633 (N_13633,N_13378,N_13494);
or U13634 (N_13634,N_13480,N_13264);
xnor U13635 (N_13635,N_13306,N_13310);
xnor U13636 (N_13636,N_13395,N_13407);
xor U13637 (N_13637,N_13347,N_13268);
nand U13638 (N_13638,N_13253,N_13355);
nand U13639 (N_13639,N_13212,N_13410);
xnor U13640 (N_13640,N_13237,N_13210);
and U13641 (N_13641,N_13331,N_13365);
nand U13642 (N_13642,N_13285,N_13270);
or U13643 (N_13643,N_13353,N_13439);
nor U13644 (N_13644,N_13406,N_13278);
nor U13645 (N_13645,N_13429,N_13287);
nor U13646 (N_13646,N_13293,N_13482);
xor U13647 (N_13647,N_13200,N_13222);
xor U13648 (N_13648,N_13345,N_13387);
nor U13649 (N_13649,N_13281,N_13232);
nor U13650 (N_13650,N_13206,N_13371);
xnor U13651 (N_13651,N_13401,N_13370);
xor U13652 (N_13652,N_13273,N_13395);
or U13653 (N_13653,N_13455,N_13419);
and U13654 (N_13654,N_13426,N_13365);
or U13655 (N_13655,N_13354,N_13280);
nor U13656 (N_13656,N_13496,N_13306);
nand U13657 (N_13657,N_13420,N_13366);
and U13658 (N_13658,N_13273,N_13264);
nor U13659 (N_13659,N_13238,N_13277);
or U13660 (N_13660,N_13460,N_13375);
nand U13661 (N_13661,N_13360,N_13402);
and U13662 (N_13662,N_13352,N_13438);
xor U13663 (N_13663,N_13494,N_13355);
and U13664 (N_13664,N_13385,N_13324);
xnor U13665 (N_13665,N_13322,N_13491);
and U13666 (N_13666,N_13485,N_13409);
and U13667 (N_13667,N_13394,N_13297);
and U13668 (N_13668,N_13397,N_13476);
and U13669 (N_13669,N_13236,N_13372);
xnor U13670 (N_13670,N_13466,N_13264);
nand U13671 (N_13671,N_13360,N_13226);
xnor U13672 (N_13672,N_13224,N_13378);
and U13673 (N_13673,N_13342,N_13224);
nor U13674 (N_13674,N_13437,N_13245);
nor U13675 (N_13675,N_13409,N_13490);
and U13676 (N_13676,N_13395,N_13461);
and U13677 (N_13677,N_13251,N_13372);
xor U13678 (N_13678,N_13495,N_13337);
or U13679 (N_13679,N_13216,N_13298);
or U13680 (N_13680,N_13351,N_13257);
xnor U13681 (N_13681,N_13363,N_13310);
xnor U13682 (N_13682,N_13393,N_13323);
nor U13683 (N_13683,N_13391,N_13369);
nand U13684 (N_13684,N_13416,N_13484);
nor U13685 (N_13685,N_13442,N_13428);
xnor U13686 (N_13686,N_13350,N_13342);
or U13687 (N_13687,N_13241,N_13242);
nor U13688 (N_13688,N_13491,N_13370);
and U13689 (N_13689,N_13308,N_13258);
nor U13690 (N_13690,N_13354,N_13406);
or U13691 (N_13691,N_13265,N_13394);
nand U13692 (N_13692,N_13208,N_13299);
nand U13693 (N_13693,N_13268,N_13304);
or U13694 (N_13694,N_13368,N_13284);
nand U13695 (N_13695,N_13276,N_13316);
nand U13696 (N_13696,N_13491,N_13337);
nand U13697 (N_13697,N_13330,N_13356);
xnor U13698 (N_13698,N_13459,N_13482);
xor U13699 (N_13699,N_13485,N_13414);
nor U13700 (N_13700,N_13492,N_13314);
nor U13701 (N_13701,N_13443,N_13250);
and U13702 (N_13702,N_13418,N_13464);
nand U13703 (N_13703,N_13408,N_13346);
or U13704 (N_13704,N_13320,N_13348);
nand U13705 (N_13705,N_13428,N_13330);
or U13706 (N_13706,N_13333,N_13477);
and U13707 (N_13707,N_13365,N_13385);
and U13708 (N_13708,N_13287,N_13265);
xnor U13709 (N_13709,N_13278,N_13408);
nand U13710 (N_13710,N_13419,N_13285);
nor U13711 (N_13711,N_13266,N_13292);
nand U13712 (N_13712,N_13323,N_13233);
nand U13713 (N_13713,N_13283,N_13233);
nand U13714 (N_13714,N_13457,N_13386);
and U13715 (N_13715,N_13221,N_13294);
xor U13716 (N_13716,N_13495,N_13467);
and U13717 (N_13717,N_13496,N_13386);
nor U13718 (N_13718,N_13331,N_13421);
nor U13719 (N_13719,N_13263,N_13280);
nand U13720 (N_13720,N_13370,N_13482);
and U13721 (N_13721,N_13446,N_13495);
and U13722 (N_13722,N_13203,N_13472);
or U13723 (N_13723,N_13386,N_13479);
nand U13724 (N_13724,N_13392,N_13486);
or U13725 (N_13725,N_13247,N_13253);
xnor U13726 (N_13726,N_13234,N_13472);
and U13727 (N_13727,N_13382,N_13231);
nand U13728 (N_13728,N_13409,N_13262);
nor U13729 (N_13729,N_13399,N_13483);
xnor U13730 (N_13730,N_13405,N_13398);
and U13731 (N_13731,N_13410,N_13446);
xor U13732 (N_13732,N_13398,N_13335);
or U13733 (N_13733,N_13287,N_13349);
xnor U13734 (N_13734,N_13352,N_13351);
or U13735 (N_13735,N_13200,N_13381);
and U13736 (N_13736,N_13380,N_13389);
and U13737 (N_13737,N_13404,N_13450);
nor U13738 (N_13738,N_13242,N_13233);
xnor U13739 (N_13739,N_13255,N_13311);
or U13740 (N_13740,N_13478,N_13339);
and U13741 (N_13741,N_13473,N_13202);
nand U13742 (N_13742,N_13255,N_13461);
nand U13743 (N_13743,N_13418,N_13318);
xor U13744 (N_13744,N_13205,N_13327);
nand U13745 (N_13745,N_13440,N_13352);
and U13746 (N_13746,N_13358,N_13437);
nand U13747 (N_13747,N_13226,N_13367);
nand U13748 (N_13748,N_13397,N_13212);
xnor U13749 (N_13749,N_13398,N_13212);
nor U13750 (N_13750,N_13346,N_13389);
xnor U13751 (N_13751,N_13390,N_13291);
and U13752 (N_13752,N_13294,N_13364);
and U13753 (N_13753,N_13266,N_13367);
or U13754 (N_13754,N_13353,N_13304);
nor U13755 (N_13755,N_13375,N_13382);
or U13756 (N_13756,N_13202,N_13350);
nor U13757 (N_13757,N_13401,N_13493);
and U13758 (N_13758,N_13375,N_13365);
xor U13759 (N_13759,N_13437,N_13289);
xor U13760 (N_13760,N_13488,N_13348);
nand U13761 (N_13761,N_13210,N_13436);
xor U13762 (N_13762,N_13423,N_13230);
xor U13763 (N_13763,N_13260,N_13301);
nor U13764 (N_13764,N_13312,N_13252);
or U13765 (N_13765,N_13447,N_13352);
nor U13766 (N_13766,N_13322,N_13263);
nand U13767 (N_13767,N_13333,N_13280);
xnor U13768 (N_13768,N_13274,N_13454);
and U13769 (N_13769,N_13465,N_13342);
nand U13770 (N_13770,N_13311,N_13383);
or U13771 (N_13771,N_13292,N_13264);
and U13772 (N_13772,N_13498,N_13344);
nor U13773 (N_13773,N_13303,N_13409);
xor U13774 (N_13774,N_13200,N_13393);
or U13775 (N_13775,N_13492,N_13266);
and U13776 (N_13776,N_13331,N_13322);
and U13777 (N_13777,N_13310,N_13447);
nand U13778 (N_13778,N_13397,N_13409);
and U13779 (N_13779,N_13497,N_13218);
xnor U13780 (N_13780,N_13260,N_13461);
and U13781 (N_13781,N_13470,N_13337);
nand U13782 (N_13782,N_13305,N_13321);
and U13783 (N_13783,N_13309,N_13410);
xnor U13784 (N_13784,N_13348,N_13290);
nand U13785 (N_13785,N_13412,N_13275);
xnor U13786 (N_13786,N_13435,N_13418);
and U13787 (N_13787,N_13373,N_13394);
or U13788 (N_13788,N_13448,N_13330);
nor U13789 (N_13789,N_13453,N_13492);
nand U13790 (N_13790,N_13216,N_13494);
xnor U13791 (N_13791,N_13273,N_13239);
nand U13792 (N_13792,N_13262,N_13202);
nand U13793 (N_13793,N_13394,N_13241);
nor U13794 (N_13794,N_13383,N_13394);
nor U13795 (N_13795,N_13318,N_13209);
nor U13796 (N_13796,N_13366,N_13338);
or U13797 (N_13797,N_13353,N_13256);
nand U13798 (N_13798,N_13470,N_13359);
nor U13799 (N_13799,N_13407,N_13263);
and U13800 (N_13800,N_13512,N_13704);
nor U13801 (N_13801,N_13665,N_13672);
nand U13802 (N_13802,N_13646,N_13670);
xor U13803 (N_13803,N_13707,N_13727);
nand U13804 (N_13804,N_13630,N_13615);
or U13805 (N_13805,N_13641,N_13793);
and U13806 (N_13806,N_13504,N_13509);
and U13807 (N_13807,N_13576,N_13786);
nor U13808 (N_13808,N_13533,N_13739);
xnor U13809 (N_13809,N_13703,N_13575);
and U13810 (N_13810,N_13563,N_13668);
nor U13811 (N_13811,N_13626,N_13518);
and U13812 (N_13812,N_13769,N_13729);
nand U13813 (N_13813,N_13607,N_13652);
nand U13814 (N_13814,N_13708,N_13523);
and U13815 (N_13815,N_13642,N_13647);
and U13816 (N_13816,N_13751,N_13578);
nand U13817 (N_13817,N_13543,N_13595);
nand U13818 (N_13818,N_13745,N_13763);
xor U13819 (N_13819,N_13757,N_13795);
and U13820 (N_13820,N_13591,N_13606);
nor U13821 (N_13821,N_13726,N_13722);
and U13822 (N_13822,N_13621,N_13577);
nand U13823 (N_13823,N_13560,N_13515);
and U13824 (N_13824,N_13691,N_13545);
nor U13825 (N_13825,N_13564,N_13603);
or U13826 (N_13826,N_13746,N_13624);
and U13827 (N_13827,N_13737,N_13747);
nand U13828 (N_13828,N_13549,N_13594);
or U13829 (N_13829,N_13659,N_13649);
and U13830 (N_13830,N_13787,N_13521);
nand U13831 (N_13831,N_13532,N_13669);
xor U13832 (N_13832,N_13799,N_13548);
nand U13833 (N_13833,N_13540,N_13681);
nor U13834 (N_13834,N_13655,N_13536);
and U13835 (N_13835,N_13710,N_13782);
nor U13836 (N_13836,N_13752,N_13709);
or U13837 (N_13837,N_13645,N_13663);
nand U13838 (N_13838,N_13590,N_13565);
and U13839 (N_13839,N_13559,N_13654);
nor U13840 (N_13840,N_13785,N_13612);
and U13841 (N_13841,N_13776,N_13625);
or U13842 (N_13842,N_13748,N_13608);
xor U13843 (N_13843,N_13721,N_13713);
nand U13844 (N_13844,N_13679,N_13740);
nor U13845 (N_13845,N_13601,N_13653);
or U13846 (N_13846,N_13728,N_13667);
nand U13847 (N_13847,N_13586,N_13724);
nor U13848 (N_13848,N_13566,N_13730);
or U13849 (N_13849,N_13584,N_13770);
nand U13850 (N_13850,N_13680,N_13749);
nand U13851 (N_13851,N_13597,N_13609);
or U13852 (N_13852,N_13592,N_13706);
nor U13853 (N_13853,N_13554,N_13750);
nand U13854 (N_13854,N_13682,N_13526);
or U13855 (N_13855,N_13767,N_13535);
or U13856 (N_13856,N_13735,N_13598);
xor U13857 (N_13857,N_13501,N_13517);
and U13858 (N_13858,N_13503,N_13781);
or U13859 (N_13859,N_13695,N_13705);
nor U13860 (N_13860,N_13761,N_13677);
and U13861 (N_13861,N_13676,N_13502);
or U13862 (N_13862,N_13760,N_13620);
nor U13863 (N_13863,N_13696,N_13765);
or U13864 (N_13864,N_13604,N_13519);
xnor U13865 (N_13865,N_13513,N_13500);
and U13866 (N_13866,N_13797,N_13508);
xnor U13867 (N_13867,N_13700,N_13694);
or U13868 (N_13868,N_13666,N_13628);
xnor U13869 (N_13869,N_13798,N_13585);
nor U13870 (N_13870,N_13611,N_13553);
xnor U13871 (N_13871,N_13675,N_13617);
nand U13872 (N_13872,N_13725,N_13651);
xnor U13873 (N_13873,N_13744,N_13593);
xor U13874 (N_13874,N_13683,N_13734);
nor U13875 (N_13875,N_13759,N_13661);
or U13876 (N_13876,N_13531,N_13562);
nor U13877 (N_13877,N_13511,N_13534);
and U13878 (N_13878,N_13627,N_13778);
or U13879 (N_13879,N_13633,N_13580);
xor U13880 (N_13880,N_13567,N_13688);
xnor U13881 (N_13881,N_13522,N_13678);
or U13882 (N_13882,N_13643,N_13636);
and U13883 (N_13883,N_13557,N_13600);
and U13884 (N_13884,N_13736,N_13768);
and U13885 (N_13885,N_13637,N_13648);
xor U13886 (N_13886,N_13605,N_13658);
and U13887 (N_13887,N_13715,N_13650);
or U13888 (N_13888,N_13506,N_13690);
and U13889 (N_13889,N_13790,N_13719);
nor U13890 (N_13890,N_13572,N_13570);
nor U13891 (N_13891,N_13568,N_13716);
or U13892 (N_13892,N_13689,N_13635);
nand U13893 (N_13893,N_13662,N_13552);
and U13894 (N_13894,N_13796,N_13547);
nand U13895 (N_13895,N_13610,N_13783);
or U13896 (N_13896,N_13530,N_13520);
nand U13897 (N_13897,N_13777,N_13656);
xor U13898 (N_13898,N_13774,N_13673);
nand U13899 (N_13899,N_13657,N_13743);
nand U13900 (N_13900,N_13556,N_13525);
nor U13901 (N_13901,N_13784,N_13514);
nor U13902 (N_13902,N_13773,N_13766);
xor U13903 (N_13903,N_13771,N_13583);
and U13904 (N_13904,N_13596,N_13634);
and U13905 (N_13905,N_13714,N_13664);
nor U13906 (N_13906,N_13619,N_13640);
and U13907 (N_13907,N_13622,N_13685);
xor U13908 (N_13908,N_13632,N_13623);
and U13909 (N_13909,N_13550,N_13582);
nor U13910 (N_13910,N_13794,N_13711);
and U13911 (N_13911,N_13764,N_13701);
xor U13912 (N_13912,N_13602,N_13697);
xnor U13913 (N_13913,N_13779,N_13754);
and U13914 (N_13914,N_13524,N_13758);
and U13915 (N_13915,N_13720,N_13756);
nor U13916 (N_13916,N_13588,N_13712);
and U13917 (N_13917,N_13546,N_13762);
and U13918 (N_13918,N_13528,N_13573);
or U13919 (N_13919,N_13780,N_13698);
or U13920 (N_13920,N_13741,N_13537);
or U13921 (N_13921,N_13732,N_13529);
or U13922 (N_13922,N_13516,N_13693);
nand U13923 (N_13923,N_13558,N_13718);
xor U13924 (N_13924,N_13731,N_13733);
xor U13925 (N_13925,N_13723,N_13541);
nor U13926 (N_13926,N_13687,N_13671);
or U13927 (N_13927,N_13772,N_13589);
or U13928 (N_13928,N_13755,N_13544);
or U13929 (N_13929,N_13738,N_13539);
or U13930 (N_13930,N_13613,N_13789);
nor U13931 (N_13931,N_13644,N_13692);
or U13932 (N_13932,N_13555,N_13579);
or U13933 (N_13933,N_13791,N_13792);
or U13934 (N_13934,N_13569,N_13614);
and U13935 (N_13935,N_13631,N_13542);
or U13936 (N_13936,N_13616,N_13551);
nand U13937 (N_13937,N_13581,N_13639);
or U13938 (N_13938,N_13629,N_13505);
or U13939 (N_13939,N_13660,N_13753);
and U13940 (N_13940,N_13686,N_13618);
xor U13941 (N_13941,N_13538,N_13574);
nor U13942 (N_13942,N_13702,N_13775);
or U13943 (N_13943,N_13507,N_13527);
xor U13944 (N_13944,N_13587,N_13717);
and U13945 (N_13945,N_13699,N_13684);
nor U13946 (N_13946,N_13510,N_13638);
and U13947 (N_13947,N_13561,N_13599);
nand U13948 (N_13948,N_13742,N_13571);
xor U13949 (N_13949,N_13674,N_13788);
nand U13950 (N_13950,N_13546,N_13589);
or U13951 (N_13951,N_13611,N_13765);
nand U13952 (N_13952,N_13781,N_13707);
nand U13953 (N_13953,N_13631,N_13643);
nand U13954 (N_13954,N_13535,N_13608);
nor U13955 (N_13955,N_13586,N_13552);
nand U13956 (N_13956,N_13662,N_13562);
xnor U13957 (N_13957,N_13545,N_13517);
xor U13958 (N_13958,N_13671,N_13759);
nor U13959 (N_13959,N_13675,N_13793);
xnor U13960 (N_13960,N_13740,N_13669);
nand U13961 (N_13961,N_13636,N_13529);
or U13962 (N_13962,N_13762,N_13645);
or U13963 (N_13963,N_13590,N_13690);
xor U13964 (N_13964,N_13563,N_13656);
nor U13965 (N_13965,N_13720,N_13545);
and U13966 (N_13966,N_13577,N_13664);
xor U13967 (N_13967,N_13536,N_13654);
nand U13968 (N_13968,N_13655,N_13743);
nor U13969 (N_13969,N_13611,N_13506);
and U13970 (N_13970,N_13550,N_13549);
or U13971 (N_13971,N_13508,N_13795);
xor U13972 (N_13972,N_13744,N_13620);
and U13973 (N_13973,N_13551,N_13620);
nor U13974 (N_13974,N_13525,N_13785);
and U13975 (N_13975,N_13601,N_13535);
nand U13976 (N_13976,N_13591,N_13757);
xnor U13977 (N_13977,N_13693,N_13690);
nor U13978 (N_13978,N_13571,N_13754);
nand U13979 (N_13979,N_13519,N_13674);
xor U13980 (N_13980,N_13736,N_13632);
nor U13981 (N_13981,N_13713,N_13550);
or U13982 (N_13982,N_13711,N_13636);
nor U13983 (N_13983,N_13739,N_13700);
nand U13984 (N_13984,N_13761,N_13779);
and U13985 (N_13985,N_13676,N_13645);
xor U13986 (N_13986,N_13710,N_13502);
and U13987 (N_13987,N_13516,N_13792);
nand U13988 (N_13988,N_13573,N_13742);
xnor U13989 (N_13989,N_13609,N_13507);
xnor U13990 (N_13990,N_13653,N_13521);
nor U13991 (N_13991,N_13525,N_13682);
xor U13992 (N_13992,N_13768,N_13683);
and U13993 (N_13993,N_13734,N_13535);
and U13994 (N_13994,N_13505,N_13785);
and U13995 (N_13995,N_13799,N_13601);
or U13996 (N_13996,N_13501,N_13562);
nand U13997 (N_13997,N_13620,N_13781);
or U13998 (N_13998,N_13598,N_13745);
nor U13999 (N_13999,N_13765,N_13724);
xnor U14000 (N_14000,N_13739,N_13527);
and U14001 (N_14001,N_13776,N_13736);
and U14002 (N_14002,N_13504,N_13642);
nand U14003 (N_14003,N_13645,N_13621);
nor U14004 (N_14004,N_13560,N_13655);
and U14005 (N_14005,N_13764,N_13577);
nand U14006 (N_14006,N_13669,N_13528);
xnor U14007 (N_14007,N_13769,N_13611);
nand U14008 (N_14008,N_13751,N_13612);
and U14009 (N_14009,N_13648,N_13642);
nand U14010 (N_14010,N_13593,N_13641);
and U14011 (N_14011,N_13536,N_13669);
or U14012 (N_14012,N_13745,N_13567);
xnor U14013 (N_14013,N_13517,N_13796);
and U14014 (N_14014,N_13637,N_13508);
xnor U14015 (N_14015,N_13722,N_13524);
or U14016 (N_14016,N_13628,N_13760);
nor U14017 (N_14017,N_13583,N_13522);
nor U14018 (N_14018,N_13544,N_13789);
nand U14019 (N_14019,N_13505,N_13660);
nand U14020 (N_14020,N_13513,N_13618);
or U14021 (N_14021,N_13766,N_13613);
or U14022 (N_14022,N_13777,N_13598);
or U14023 (N_14023,N_13638,N_13684);
and U14024 (N_14024,N_13616,N_13569);
nand U14025 (N_14025,N_13535,N_13580);
xnor U14026 (N_14026,N_13678,N_13782);
nand U14027 (N_14027,N_13509,N_13620);
or U14028 (N_14028,N_13623,N_13629);
and U14029 (N_14029,N_13537,N_13740);
nand U14030 (N_14030,N_13543,N_13650);
nor U14031 (N_14031,N_13763,N_13556);
xor U14032 (N_14032,N_13525,N_13702);
or U14033 (N_14033,N_13595,N_13565);
and U14034 (N_14034,N_13602,N_13634);
and U14035 (N_14035,N_13695,N_13749);
xnor U14036 (N_14036,N_13761,N_13634);
or U14037 (N_14037,N_13661,N_13627);
xnor U14038 (N_14038,N_13724,N_13773);
nand U14039 (N_14039,N_13786,N_13584);
nand U14040 (N_14040,N_13789,N_13552);
nor U14041 (N_14041,N_13544,N_13635);
nor U14042 (N_14042,N_13502,N_13605);
nand U14043 (N_14043,N_13793,N_13795);
or U14044 (N_14044,N_13720,N_13762);
xnor U14045 (N_14045,N_13762,N_13514);
and U14046 (N_14046,N_13781,N_13525);
or U14047 (N_14047,N_13795,N_13585);
and U14048 (N_14048,N_13793,N_13757);
xor U14049 (N_14049,N_13517,N_13779);
nor U14050 (N_14050,N_13736,N_13592);
and U14051 (N_14051,N_13646,N_13655);
nor U14052 (N_14052,N_13659,N_13545);
nor U14053 (N_14053,N_13708,N_13543);
xnor U14054 (N_14054,N_13653,N_13511);
or U14055 (N_14055,N_13666,N_13522);
nand U14056 (N_14056,N_13583,N_13534);
or U14057 (N_14057,N_13738,N_13542);
and U14058 (N_14058,N_13537,N_13714);
or U14059 (N_14059,N_13615,N_13593);
nor U14060 (N_14060,N_13593,N_13787);
and U14061 (N_14061,N_13757,N_13799);
nand U14062 (N_14062,N_13648,N_13541);
and U14063 (N_14063,N_13550,N_13534);
or U14064 (N_14064,N_13732,N_13565);
xnor U14065 (N_14065,N_13726,N_13535);
nand U14066 (N_14066,N_13659,N_13507);
nor U14067 (N_14067,N_13624,N_13737);
or U14068 (N_14068,N_13591,N_13645);
nor U14069 (N_14069,N_13722,N_13634);
nand U14070 (N_14070,N_13562,N_13693);
xor U14071 (N_14071,N_13518,N_13630);
nor U14072 (N_14072,N_13613,N_13501);
xor U14073 (N_14073,N_13502,N_13718);
nand U14074 (N_14074,N_13563,N_13776);
and U14075 (N_14075,N_13670,N_13583);
nor U14076 (N_14076,N_13558,N_13527);
or U14077 (N_14077,N_13790,N_13692);
nor U14078 (N_14078,N_13615,N_13737);
or U14079 (N_14079,N_13509,N_13687);
nor U14080 (N_14080,N_13621,N_13617);
nor U14081 (N_14081,N_13685,N_13770);
and U14082 (N_14082,N_13770,N_13690);
and U14083 (N_14083,N_13719,N_13723);
nor U14084 (N_14084,N_13511,N_13509);
nand U14085 (N_14085,N_13597,N_13660);
xor U14086 (N_14086,N_13775,N_13779);
xor U14087 (N_14087,N_13745,N_13622);
and U14088 (N_14088,N_13796,N_13785);
nand U14089 (N_14089,N_13506,N_13722);
xor U14090 (N_14090,N_13721,N_13705);
nor U14091 (N_14091,N_13547,N_13552);
nor U14092 (N_14092,N_13794,N_13686);
and U14093 (N_14093,N_13761,N_13722);
nand U14094 (N_14094,N_13548,N_13715);
xnor U14095 (N_14095,N_13781,N_13565);
nand U14096 (N_14096,N_13602,N_13519);
and U14097 (N_14097,N_13590,N_13595);
nand U14098 (N_14098,N_13568,N_13534);
and U14099 (N_14099,N_13730,N_13661);
and U14100 (N_14100,N_13828,N_13864);
and U14101 (N_14101,N_14017,N_13913);
and U14102 (N_14102,N_13836,N_13943);
and U14103 (N_14103,N_13955,N_13965);
nor U14104 (N_14104,N_13893,N_13963);
nand U14105 (N_14105,N_13876,N_13996);
or U14106 (N_14106,N_13928,N_14056);
nor U14107 (N_14107,N_13948,N_13842);
xnor U14108 (N_14108,N_14014,N_14057);
or U14109 (N_14109,N_14088,N_13950);
nand U14110 (N_14110,N_14035,N_14095);
or U14111 (N_14111,N_13824,N_14062);
and U14112 (N_14112,N_13885,N_13802);
or U14113 (N_14113,N_14010,N_13917);
nor U14114 (N_14114,N_14066,N_14071);
nand U14115 (N_14115,N_13947,N_13961);
or U14116 (N_14116,N_13859,N_13811);
xor U14117 (N_14117,N_13863,N_14027);
or U14118 (N_14118,N_14031,N_13887);
nor U14119 (N_14119,N_14079,N_13967);
nand U14120 (N_14120,N_14093,N_14016);
xnor U14121 (N_14121,N_14084,N_14067);
and U14122 (N_14122,N_13998,N_13982);
nand U14123 (N_14123,N_13924,N_13820);
xnor U14124 (N_14124,N_14051,N_13976);
or U14125 (N_14125,N_13986,N_13891);
xor U14126 (N_14126,N_14006,N_13946);
nor U14127 (N_14127,N_14078,N_13980);
nand U14128 (N_14128,N_13894,N_14099);
xnor U14129 (N_14129,N_14007,N_14075);
nor U14130 (N_14130,N_14040,N_13892);
or U14131 (N_14131,N_14030,N_13845);
and U14132 (N_14132,N_13973,N_13971);
xor U14133 (N_14133,N_14072,N_13869);
or U14134 (N_14134,N_13997,N_13911);
nand U14135 (N_14135,N_13930,N_13933);
nor U14136 (N_14136,N_13932,N_13877);
and U14137 (N_14137,N_13860,N_13839);
or U14138 (N_14138,N_13992,N_13935);
nor U14139 (N_14139,N_13847,N_13871);
or U14140 (N_14140,N_13926,N_14073);
and U14141 (N_14141,N_13964,N_13919);
xor U14142 (N_14142,N_14024,N_13931);
nand U14143 (N_14143,N_13800,N_13814);
nand U14144 (N_14144,N_14052,N_13835);
xnor U14145 (N_14145,N_13848,N_13858);
nand U14146 (N_14146,N_13880,N_13874);
nor U14147 (N_14147,N_14025,N_13881);
nand U14148 (N_14148,N_13957,N_13870);
or U14149 (N_14149,N_14008,N_13900);
nor U14150 (N_14150,N_13896,N_13807);
xor U14151 (N_14151,N_13938,N_14022);
nor U14152 (N_14152,N_13993,N_13805);
and U14153 (N_14153,N_13899,N_14068);
or U14154 (N_14154,N_13868,N_13903);
nand U14155 (N_14155,N_13939,N_13974);
and U14156 (N_14156,N_13921,N_14003);
and U14157 (N_14157,N_13825,N_14080);
and U14158 (N_14158,N_13987,N_13873);
nor U14159 (N_14159,N_13856,N_13831);
and U14160 (N_14160,N_13975,N_14055);
nand U14161 (N_14161,N_13968,N_13949);
nor U14162 (N_14162,N_14038,N_13951);
or U14163 (N_14163,N_13834,N_14076);
and U14164 (N_14164,N_13819,N_14091);
nand U14165 (N_14165,N_13907,N_13806);
or U14166 (N_14166,N_13940,N_14023);
or U14167 (N_14167,N_13840,N_13843);
xor U14168 (N_14168,N_13808,N_14042);
nand U14169 (N_14169,N_13956,N_13920);
nand U14170 (N_14170,N_13875,N_13882);
nor U14171 (N_14171,N_13857,N_14096);
or U14172 (N_14172,N_13945,N_13905);
or U14173 (N_14173,N_13815,N_14061);
or U14174 (N_14174,N_13898,N_13929);
nor U14175 (N_14175,N_14060,N_14029);
nor U14176 (N_14176,N_14009,N_14020);
and U14177 (N_14177,N_13809,N_13988);
and U14178 (N_14178,N_13852,N_14034);
and U14179 (N_14179,N_14049,N_13972);
nand U14180 (N_14180,N_13959,N_14069);
or U14181 (N_14181,N_13983,N_14089);
nand U14182 (N_14182,N_14000,N_13902);
nor U14183 (N_14183,N_13867,N_13906);
nand U14184 (N_14184,N_13995,N_13994);
nor U14185 (N_14185,N_14043,N_13884);
xnor U14186 (N_14186,N_13878,N_14026);
nand U14187 (N_14187,N_14081,N_13944);
or U14188 (N_14188,N_13927,N_14033);
nand U14189 (N_14189,N_13901,N_13810);
nor U14190 (N_14190,N_13801,N_13883);
or U14191 (N_14191,N_14044,N_13990);
and U14192 (N_14192,N_13912,N_13841);
and U14193 (N_14193,N_13851,N_13979);
xor U14194 (N_14194,N_13952,N_13826);
or U14195 (N_14195,N_13984,N_13999);
or U14196 (N_14196,N_14059,N_14082);
nor U14197 (N_14197,N_13832,N_13897);
and U14198 (N_14198,N_13960,N_14021);
xnor U14199 (N_14199,N_14064,N_13886);
and U14200 (N_14200,N_14013,N_14015);
or U14201 (N_14201,N_13889,N_14085);
and U14202 (N_14202,N_13895,N_13844);
xor U14203 (N_14203,N_14087,N_14039);
nor U14204 (N_14204,N_13991,N_14094);
xor U14205 (N_14205,N_13890,N_14053);
xor U14206 (N_14206,N_14065,N_13977);
nand U14207 (N_14207,N_13914,N_14050);
xnor U14208 (N_14208,N_13925,N_14077);
nand U14209 (N_14209,N_14092,N_13812);
xor U14210 (N_14210,N_13915,N_13837);
or U14211 (N_14211,N_13942,N_13846);
xor U14212 (N_14212,N_14090,N_13849);
xnor U14213 (N_14213,N_14048,N_14001);
or U14214 (N_14214,N_14012,N_13855);
xor U14215 (N_14215,N_13888,N_14086);
and U14216 (N_14216,N_13953,N_14028);
nor U14217 (N_14217,N_14058,N_13962);
or U14218 (N_14218,N_13827,N_13818);
and U14219 (N_14219,N_14011,N_13937);
nor U14220 (N_14220,N_14037,N_13934);
or U14221 (N_14221,N_13923,N_13908);
nand U14222 (N_14222,N_13804,N_13866);
nand U14223 (N_14223,N_14074,N_13861);
nand U14224 (N_14224,N_13916,N_14083);
nand U14225 (N_14225,N_14041,N_13922);
nor U14226 (N_14226,N_13941,N_14070);
or U14227 (N_14227,N_13803,N_13872);
nand U14228 (N_14228,N_14032,N_13978);
nor U14229 (N_14229,N_13904,N_14005);
nand U14230 (N_14230,N_13969,N_13817);
and U14231 (N_14231,N_13829,N_13854);
or U14232 (N_14232,N_14018,N_13966);
and U14233 (N_14233,N_14036,N_13909);
nand U14234 (N_14234,N_13862,N_13936);
or U14235 (N_14235,N_13985,N_14046);
nor U14236 (N_14236,N_14047,N_14002);
and U14237 (N_14237,N_13970,N_14063);
xnor U14238 (N_14238,N_13879,N_13958);
xnor U14239 (N_14239,N_13823,N_14097);
xor U14240 (N_14240,N_13865,N_14054);
nor U14241 (N_14241,N_13813,N_13954);
nor U14242 (N_14242,N_13816,N_14004);
and U14243 (N_14243,N_14098,N_13822);
and U14244 (N_14244,N_13989,N_13853);
xnor U14245 (N_14245,N_13821,N_14045);
nand U14246 (N_14246,N_14019,N_13830);
or U14247 (N_14247,N_13833,N_13838);
nor U14248 (N_14248,N_13910,N_13918);
nor U14249 (N_14249,N_13850,N_13981);
nor U14250 (N_14250,N_13996,N_13802);
and U14251 (N_14251,N_14054,N_14041);
nand U14252 (N_14252,N_13809,N_14052);
nand U14253 (N_14253,N_13934,N_13900);
nor U14254 (N_14254,N_13983,N_13868);
nor U14255 (N_14255,N_13886,N_14018);
xor U14256 (N_14256,N_13818,N_13831);
nand U14257 (N_14257,N_13926,N_14026);
nor U14258 (N_14258,N_13871,N_13996);
nand U14259 (N_14259,N_14032,N_13990);
nor U14260 (N_14260,N_13823,N_13812);
xnor U14261 (N_14261,N_13956,N_14066);
nor U14262 (N_14262,N_14088,N_13835);
or U14263 (N_14263,N_14037,N_13915);
nand U14264 (N_14264,N_13948,N_13972);
nand U14265 (N_14265,N_13950,N_14089);
and U14266 (N_14266,N_13958,N_14074);
nor U14267 (N_14267,N_14053,N_14031);
or U14268 (N_14268,N_13881,N_14091);
and U14269 (N_14269,N_14070,N_13897);
or U14270 (N_14270,N_14023,N_13893);
nor U14271 (N_14271,N_14002,N_14012);
nand U14272 (N_14272,N_13980,N_14019);
or U14273 (N_14273,N_13895,N_13933);
nor U14274 (N_14274,N_13982,N_13885);
nand U14275 (N_14275,N_13855,N_14013);
xnor U14276 (N_14276,N_14065,N_13995);
xor U14277 (N_14277,N_13905,N_13980);
and U14278 (N_14278,N_13975,N_13943);
nor U14279 (N_14279,N_13948,N_14055);
xor U14280 (N_14280,N_13926,N_13800);
nor U14281 (N_14281,N_14034,N_13945);
nand U14282 (N_14282,N_13841,N_13831);
and U14283 (N_14283,N_13887,N_13824);
or U14284 (N_14284,N_13918,N_13863);
or U14285 (N_14285,N_14063,N_14044);
nor U14286 (N_14286,N_13840,N_13846);
or U14287 (N_14287,N_13916,N_13950);
or U14288 (N_14288,N_13805,N_13939);
or U14289 (N_14289,N_13880,N_13972);
and U14290 (N_14290,N_13867,N_13920);
nand U14291 (N_14291,N_13858,N_14015);
and U14292 (N_14292,N_13826,N_14014);
xnor U14293 (N_14293,N_13906,N_13818);
xnor U14294 (N_14294,N_13862,N_13988);
and U14295 (N_14295,N_14097,N_14006);
and U14296 (N_14296,N_13842,N_14021);
and U14297 (N_14297,N_13834,N_13929);
or U14298 (N_14298,N_13940,N_14039);
nand U14299 (N_14299,N_14020,N_13854);
and U14300 (N_14300,N_13924,N_14016);
or U14301 (N_14301,N_14093,N_13813);
or U14302 (N_14302,N_14089,N_13859);
xor U14303 (N_14303,N_14017,N_14019);
nor U14304 (N_14304,N_13885,N_13993);
nor U14305 (N_14305,N_13963,N_13804);
xnor U14306 (N_14306,N_13905,N_13851);
xnor U14307 (N_14307,N_14046,N_13873);
nand U14308 (N_14308,N_13830,N_13822);
nand U14309 (N_14309,N_13945,N_14039);
and U14310 (N_14310,N_13980,N_14039);
and U14311 (N_14311,N_13894,N_13971);
and U14312 (N_14312,N_13949,N_14059);
and U14313 (N_14313,N_14077,N_14090);
nor U14314 (N_14314,N_13870,N_13994);
nor U14315 (N_14315,N_13929,N_13947);
or U14316 (N_14316,N_14057,N_13882);
nor U14317 (N_14317,N_13978,N_13872);
nand U14318 (N_14318,N_13810,N_14093);
or U14319 (N_14319,N_14027,N_13987);
nor U14320 (N_14320,N_14031,N_13932);
xor U14321 (N_14321,N_13930,N_14063);
or U14322 (N_14322,N_14062,N_14095);
nand U14323 (N_14323,N_13869,N_14020);
or U14324 (N_14324,N_14014,N_13947);
nand U14325 (N_14325,N_13807,N_14048);
and U14326 (N_14326,N_13825,N_14081);
and U14327 (N_14327,N_13971,N_14060);
xnor U14328 (N_14328,N_14076,N_13964);
and U14329 (N_14329,N_13915,N_14075);
and U14330 (N_14330,N_13839,N_13861);
or U14331 (N_14331,N_13954,N_14077);
nor U14332 (N_14332,N_14054,N_13907);
nor U14333 (N_14333,N_13855,N_14064);
xnor U14334 (N_14334,N_13940,N_14053);
or U14335 (N_14335,N_13989,N_13804);
and U14336 (N_14336,N_14069,N_14062);
and U14337 (N_14337,N_13886,N_13922);
and U14338 (N_14338,N_13886,N_13966);
nand U14339 (N_14339,N_13802,N_14072);
or U14340 (N_14340,N_14019,N_13867);
and U14341 (N_14341,N_13966,N_13847);
and U14342 (N_14342,N_13916,N_14043);
nand U14343 (N_14343,N_13834,N_13996);
xor U14344 (N_14344,N_13939,N_14083);
nand U14345 (N_14345,N_13905,N_13918);
xnor U14346 (N_14346,N_13826,N_13889);
nor U14347 (N_14347,N_13813,N_14039);
or U14348 (N_14348,N_13861,N_13993);
and U14349 (N_14349,N_14044,N_14003);
nor U14350 (N_14350,N_13999,N_13935);
nor U14351 (N_14351,N_13808,N_13828);
nand U14352 (N_14352,N_14048,N_13859);
nor U14353 (N_14353,N_13819,N_14016);
xor U14354 (N_14354,N_13867,N_13973);
or U14355 (N_14355,N_14076,N_13950);
or U14356 (N_14356,N_13855,N_14066);
and U14357 (N_14357,N_13881,N_13926);
nand U14358 (N_14358,N_14022,N_13994);
or U14359 (N_14359,N_13870,N_13979);
nor U14360 (N_14360,N_13969,N_14057);
xor U14361 (N_14361,N_14060,N_13898);
nand U14362 (N_14362,N_13918,N_14067);
nand U14363 (N_14363,N_14058,N_13886);
nor U14364 (N_14364,N_14053,N_14080);
and U14365 (N_14365,N_13915,N_13921);
nor U14366 (N_14366,N_13895,N_13952);
nand U14367 (N_14367,N_13871,N_13803);
and U14368 (N_14368,N_14097,N_14026);
nand U14369 (N_14369,N_13923,N_13828);
or U14370 (N_14370,N_13805,N_13900);
nor U14371 (N_14371,N_13883,N_13938);
or U14372 (N_14372,N_13806,N_14062);
xnor U14373 (N_14373,N_14084,N_13831);
or U14374 (N_14374,N_13809,N_13826);
nand U14375 (N_14375,N_14078,N_13815);
or U14376 (N_14376,N_14099,N_13908);
or U14377 (N_14377,N_13993,N_13811);
xor U14378 (N_14378,N_13906,N_14051);
nand U14379 (N_14379,N_13814,N_13813);
nand U14380 (N_14380,N_14041,N_14049);
and U14381 (N_14381,N_13918,N_13877);
nand U14382 (N_14382,N_13975,N_13867);
nand U14383 (N_14383,N_14000,N_13935);
and U14384 (N_14384,N_14078,N_13881);
xor U14385 (N_14385,N_13924,N_13929);
nand U14386 (N_14386,N_14093,N_13829);
nand U14387 (N_14387,N_13924,N_14089);
nor U14388 (N_14388,N_13803,N_13873);
nand U14389 (N_14389,N_13872,N_13983);
xor U14390 (N_14390,N_14059,N_14043);
and U14391 (N_14391,N_13928,N_14008);
nor U14392 (N_14392,N_13975,N_13973);
or U14393 (N_14393,N_13930,N_13833);
and U14394 (N_14394,N_13965,N_13896);
xor U14395 (N_14395,N_13803,N_13943);
nor U14396 (N_14396,N_14089,N_14072);
nand U14397 (N_14397,N_13997,N_13953);
and U14398 (N_14398,N_13983,N_14065);
or U14399 (N_14399,N_13982,N_13856);
nor U14400 (N_14400,N_14143,N_14360);
nand U14401 (N_14401,N_14135,N_14123);
or U14402 (N_14402,N_14285,N_14374);
xnor U14403 (N_14403,N_14392,N_14241);
nand U14404 (N_14404,N_14362,N_14179);
or U14405 (N_14405,N_14152,N_14365);
xnor U14406 (N_14406,N_14363,N_14265);
nand U14407 (N_14407,N_14234,N_14187);
nor U14408 (N_14408,N_14289,N_14367);
or U14409 (N_14409,N_14314,N_14346);
and U14410 (N_14410,N_14116,N_14120);
nor U14411 (N_14411,N_14303,N_14221);
nor U14412 (N_14412,N_14100,N_14337);
xnor U14413 (N_14413,N_14262,N_14345);
and U14414 (N_14414,N_14249,N_14259);
and U14415 (N_14415,N_14390,N_14385);
and U14416 (N_14416,N_14292,N_14293);
xnor U14417 (N_14417,N_14266,N_14319);
or U14418 (N_14418,N_14202,N_14258);
nand U14419 (N_14419,N_14338,N_14284);
or U14420 (N_14420,N_14190,N_14255);
and U14421 (N_14421,N_14272,N_14307);
and U14422 (N_14422,N_14324,N_14162);
or U14423 (N_14423,N_14302,N_14192);
and U14424 (N_14424,N_14119,N_14368);
and U14425 (N_14425,N_14348,N_14250);
or U14426 (N_14426,N_14261,N_14147);
nor U14427 (N_14427,N_14208,N_14167);
nor U14428 (N_14428,N_14201,N_14229);
xnor U14429 (N_14429,N_14125,N_14163);
nand U14430 (N_14430,N_14198,N_14386);
nand U14431 (N_14431,N_14211,N_14233);
or U14432 (N_14432,N_14355,N_14347);
and U14433 (N_14433,N_14160,N_14349);
and U14434 (N_14434,N_14205,N_14173);
nor U14435 (N_14435,N_14137,N_14180);
xor U14436 (N_14436,N_14296,N_14339);
xor U14437 (N_14437,N_14376,N_14109);
or U14438 (N_14438,N_14220,N_14188);
and U14439 (N_14439,N_14395,N_14256);
or U14440 (N_14440,N_14216,N_14246);
nand U14441 (N_14441,N_14257,N_14154);
and U14442 (N_14442,N_14354,N_14223);
and U14443 (N_14443,N_14364,N_14254);
nor U14444 (N_14444,N_14297,N_14281);
nand U14445 (N_14445,N_14271,N_14113);
and U14446 (N_14446,N_14157,N_14299);
nand U14447 (N_14447,N_14264,N_14184);
xor U14448 (N_14448,N_14286,N_14305);
or U14449 (N_14449,N_14115,N_14290);
and U14450 (N_14450,N_14231,N_14225);
or U14451 (N_14451,N_14183,N_14164);
or U14452 (N_14452,N_14182,N_14169);
nor U14453 (N_14453,N_14295,N_14334);
and U14454 (N_14454,N_14253,N_14107);
nand U14455 (N_14455,N_14146,N_14325);
nor U14456 (N_14456,N_14318,N_14101);
and U14457 (N_14457,N_14260,N_14326);
nor U14458 (N_14458,N_14341,N_14359);
or U14459 (N_14459,N_14383,N_14219);
or U14460 (N_14460,N_14239,N_14194);
and U14461 (N_14461,N_14232,N_14397);
or U14462 (N_14462,N_14248,N_14186);
nand U14463 (N_14463,N_14171,N_14230);
nand U14464 (N_14464,N_14158,N_14329);
or U14465 (N_14465,N_14235,N_14370);
nor U14466 (N_14466,N_14149,N_14283);
xor U14467 (N_14467,N_14270,N_14336);
nand U14468 (N_14468,N_14322,N_14134);
nand U14469 (N_14469,N_14291,N_14206);
or U14470 (N_14470,N_14122,N_14207);
nor U14471 (N_14471,N_14380,N_14298);
nand U14472 (N_14472,N_14199,N_14128);
nor U14473 (N_14473,N_14103,N_14369);
nor U14474 (N_14474,N_14398,N_14175);
nor U14475 (N_14475,N_14333,N_14251);
xnor U14476 (N_14476,N_14300,N_14170);
and U14477 (N_14477,N_14165,N_14312);
nand U14478 (N_14478,N_14166,N_14138);
nand U14479 (N_14479,N_14274,N_14309);
nor U14480 (N_14480,N_14130,N_14153);
nor U14481 (N_14481,N_14136,N_14176);
and U14482 (N_14482,N_14335,N_14382);
nor U14483 (N_14483,N_14150,N_14228);
or U14484 (N_14484,N_14287,N_14222);
or U14485 (N_14485,N_14155,N_14151);
nor U14486 (N_14486,N_14379,N_14321);
and U14487 (N_14487,N_14213,N_14244);
and U14488 (N_14488,N_14375,N_14301);
nand U14489 (N_14489,N_14310,N_14140);
and U14490 (N_14490,N_14350,N_14294);
xor U14491 (N_14491,N_14282,N_14328);
and U14492 (N_14492,N_14217,N_14315);
xor U14493 (N_14493,N_14185,N_14373);
nor U14494 (N_14494,N_14378,N_14394);
nand U14495 (N_14495,N_14276,N_14215);
and U14496 (N_14496,N_14145,N_14269);
xnor U14497 (N_14497,N_14108,N_14132);
xor U14498 (N_14498,N_14237,N_14126);
and U14499 (N_14499,N_14131,N_14288);
and U14500 (N_14500,N_14263,N_14124);
nor U14501 (N_14501,N_14238,N_14267);
nor U14502 (N_14502,N_14332,N_14242);
xnor U14503 (N_14503,N_14142,N_14371);
and U14504 (N_14504,N_14189,N_14195);
and U14505 (N_14505,N_14224,N_14227);
nand U14506 (N_14506,N_14327,N_14177);
nand U14507 (N_14507,N_14148,N_14156);
or U14508 (N_14508,N_14247,N_14133);
nor U14509 (N_14509,N_14313,N_14245);
xnor U14510 (N_14510,N_14353,N_14352);
xnor U14511 (N_14511,N_14112,N_14323);
nor U14512 (N_14512,N_14320,N_14279);
nand U14513 (N_14513,N_14317,N_14191);
xor U14514 (N_14514,N_14114,N_14174);
nand U14515 (N_14515,N_14280,N_14344);
xnor U14516 (N_14516,N_14311,N_14366);
or U14517 (N_14517,N_14172,N_14278);
nand U14518 (N_14518,N_14340,N_14393);
and U14519 (N_14519,N_14168,N_14388);
nand U14520 (N_14520,N_14372,N_14252);
or U14521 (N_14521,N_14361,N_14391);
or U14522 (N_14522,N_14141,N_14331);
xor U14523 (N_14523,N_14356,N_14193);
or U14524 (N_14524,N_14197,N_14273);
nor U14525 (N_14525,N_14387,N_14357);
or U14526 (N_14526,N_14304,N_14226);
and U14527 (N_14527,N_14330,N_14209);
and U14528 (N_14528,N_14343,N_14178);
and U14529 (N_14529,N_14342,N_14161);
or U14530 (N_14530,N_14127,N_14275);
xor U14531 (N_14531,N_14316,N_14139);
xor U14532 (N_14532,N_14159,N_14117);
nor U14533 (N_14533,N_14243,N_14218);
and U14534 (N_14534,N_14214,N_14236);
nand U14535 (N_14535,N_14110,N_14210);
or U14536 (N_14536,N_14308,N_14358);
nand U14537 (N_14537,N_14200,N_14129);
nand U14538 (N_14538,N_14268,N_14203);
and U14539 (N_14539,N_14204,N_14181);
xor U14540 (N_14540,N_14306,N_14389);
nand U14541 (N_14541,N_14118,N_14399);
nor U14542 (N_14542,N_14196,N_14104);
nand U14543 (N_14543,N_14381,N_14240);
and U14544 (N_14544,N_14144,N_14396);
nand U14545 (N_14545,N_14102,N_14105);
nand U14546 (N_14546,N_14111,N_14121);
nor U14547 (N_14547,N_14384,N_14106);
nor U14548 (N_14548,N_14212,N_14277);
or U14549 (N_14549,N_14377,N_14351);
nand U14550 (N_14550,N_14330,N_14135);
nand U14551 (N_14551,N_14230,N_14303);
and U14552 (N_14552,N_14318,N_14159);
and U14553 (N_14553,N_14139,N_14165);
nand U14554 (N_14554,N_14260,N_14295);
nand U14555 (N_14555,N_14216,N_14238);
or U14556 (N_14556,N_14226,N_14219);
xnor U14557 (N_14557,N_14238,N_14378);
xor U14558 (N_14558,N_14190,N_14195);
xor U14559 (N_14559,N_14349,N_14203);
xor U14560 (N_14560,N_14305,N_14115);
nor U14561 (N_14561,N_14190,N_14122);
nand U14562 (N_14562,N_14281,N_14102);
and U14563 (N_14563,N_14304,N_14368);
xnor U14564 (N_14564,N_14276,N_14290);
nor U14565 (N_14565,N_14339,N_14154);
and U14566 (N_14566,N_14304,N_14216);
nand U14567 (N_14567,N_14275,N_14316);
xor U14568 (N_14568,N_14228,N_14158);
and U14569 (N_14569,N_14157,N_14273);
nand U14570 (N_14570,N_14261,N_14139);
nand U14571 (N_14571,N_14275,N_14167);
nand U14572 (N_14572,N_14223,N_14197);
and U14573 (N_14573,N_14178,N_14225);
xor U14574 (N_14574,N_14216,N_14166);
and U14575 (N_14575,N_14169,N_14268);
nand U14576 (N_14576,N_14237,N_14324);
or U14577 (N_14577,N_14324,N_14298);
nand U14578 (N_14578,N_14172,N_14227);
and U14579 (N_14579,N_14174,N_14185);
or U14580 (N_14580,N_14234,N_14358);
or U14581 (N_14581,N_14231,N_14139);
or U14582 (N_14582,N_14150,N_14278);
nand U14583 (N_14583,N_14387,N_14113);
or U14584 (N_14584,N_14396,N_14127);
and U14585 (N_14585,N_14152,N_14338);
or U14586 (N_14586,N_14268,N_14386);
or U14587 (N_14587,N_14236,N_14286);
and U14588 (N_14588,N_14104,N_14371);
and U14589 (N_14589,N_14222,N_14268);
xor U14590 (N_14590,N_14277,N_14182);
nand U14591 (N_14591,N_14242,N_14324);
and U14592 (N_14592,N_14372,N_14246);
or U14593 (N_14593,N_14280,N_14236);
and U14594 (N_14594,N_14249,N_14140);
nor U14595 (N_14595,N_14255,N_14318);
or U14596 (N_14596,N_14246,N_14203);
nand U14597 (N_14597,N_14135,N_14312);
or U14598 (N_14598,N_14266,N_14185);
xnor U14599 (N_14599,N_14353,N_14241);
nand U14600 (N_14600,N_14187,N_14243);
or U14601 (N_14601,N_14182,N_14151);
nand U14602 (N_14602,N_14306,N_14396);
or U14603 (N_14603,N_14248,N_14334);
xor U14604 (N_14604,N_14132,N_14321);
nand U14605 (N_14605,N_14305,N_14291);
xnor U14606 (N_14606,N_14286,N_14218);
xnor U14607 (N_14607,N_14182,N_14354);
or U14608 (N_14608,N_14322,N_14186);
xnor U14609 (N_14609,N_14373,N_14194);
and U14610 (N_14610,N_14174,N_14389);
nand U14611 (N_14611,N_14334,N_14136);
or U14612 (N_14612,N_14284,N_14348);
nand U14613 (N_14613,N_14169,N_14132);
or U14614 (N_14614,N_14246,N_14155);
nand U14615 (N_14615,N_14133,N_14105);
nand U14616 (N_14616,N_14124,N_14284);
nand U14617 (N_14617,N_14161,N_14245);
nand U14618 (N_14618,N_14220,N_14145);
and U14619 (N_14619,N_14218,N_14374);
nor U14620 (N_14620,N_14323,N_14307);
and U14621 (N_14621,N_14304,N_14374);
and U14622 (N_14622,N_14132,N_14278);
nand U14623 (N_14623,N_14295,N_14278);
xnor U14624 (N_14624,N_14316,N_14174);
xor U14625 (N_14625,N_14350,N_14101);
and U14626 (N_14626,N_14328,N_14198);
and U14627 (N_14627,N_14135,N_14239);
nor U14628 (N_14628,N_14164,N_14218);
and U14629 (N_14629,N_14369,N_14361);
nand U14630 (N_14630,N_14358,N_14118);
or U14631 (N_14631,N_14206,N_14392);
or U14632 (N_14632,N_14239,N_14341);
and U14633 (N_14633,N_14354,N_14119);
xnor U14634 (N_14634,N_14243,N_14288);
and U14635 (N_14635,N_14166,N_14380);
nand U14636 (N_14636,N_14128,N_14353);
nor U14637 (N_14637,N_14302,N_14118);
xor U14638 (N_14638,N_14294,N_14278);
xor U14639 (N_14639,N_14397,N_14385);
nor U14640 (N_14640,N_14344,N_14309);
nand U14641 (N_14641,N_14340,N_14327);
nor U14642 (N_14642,N_14258,N_14396);
and U14643 (N_14643,N_14102,N_14219);
or U14644 (N_14644,N_14172,N_14346);
and U14645 (N_14645,N_14184,N_14277);
xnor U14646 (N_14646,N_14206,N_14255);
nand U14647 (N_14647,N_14345,N_14113);
nor U14648 (N_14648,N_14337,N_14282);
or U14649 (N_14649,N_14376,N_14282);
xor U14650 (N_14650,N_14303,N_14279);
nand U14651 (N_14651,N_14146,N_14366);
and U14652 (N_14652,N_14124,N_14241);
xnor U14653 (N_14653,N_14117,N_14384);
nand U14654 (N_14654,N_14233,N_14128);
or U14655 (N_14655,N_14301,N_14290);
nor U14656 (N_14656,N_14154,N_14337);
xnor U14657 (N_14657,N_14342,N_14252);
or U14658 (N_14658,N_14103,N_14322);
nor U14659 (N_14659,N_14165,N_14366);
or U14660 (N_14660,N_14199,N_14365);
or U14661 (N_14661,N_14151,N_14272);
and U14662 (N_14662,N_14136,N_14140);
nand U14663 (N_14663,N_14177,N_14150);
nand U14664 (N_14664,N_14193,N_14218);
and U14665 (N_14665,N_14107,N_14362);
nand U14666 (N_14666,N_14279,N_14105);
nand U14667 (N_14667,N_14225,N_14343);
nor U14668 (N_14668,N_14358,N_14388);
or U14669 (N_14669,N_14166,N_14100);
nand U14670 (N_14670,N_14197,N_14131);
and U14671 (N_14671,N_14173,N_14381);
nand U14672 (N_14672,N_14280,N_14389);
and U14673 (N_14673,N_14345,N_14147);
nand U14674 (N_14674,N_14347,N_14262);
or U14675 (N_14675,N_14279,N_14273);
or U14676 (N_14676,N_14370,N_14251);
or U14677 (N_14677,N_14268,N_14397);
and U14678 (N_14678,N_14121,N_14208);
nor U14679 (N_14679,N_14187,N_14295);
and U14680 (N_14680,N_14343,N_14243);
and U14681 (N_14681,N_14134,N_14123);
or U14682 (N_14682,N_14239,N_14168);
and U14683 (N_14683,N_14239,N_14184);
nor U14684 (N_14684,N_14396,N_14261);
nand U14685 (N_14685,N_14235,N_14220);
and U14686 (N_14686,N_14188,N_14399);
nor U14687 (N_14687,N_14293,N_14230);
nor U14688 (N_14688,N_14276,N_14319);
nand U14689 (N_14689,N_14364,N_14295);
or U14690 (N_14690,N_14124,N_14314);
xor U14691 (N_14691,N_14206,N_14369);
and U14692 (N_14692,N_14265,N_14262);
nor U14693 (N_14693,N_14216,N_14229);
and U14694 (N_14694,N_14173,N_14184);
or U14695 (N_14695,N_14232,N_14105);
nand U14696 (N_14696,N_14152,N_14130);
or U14697 (N_14697,N_14171,N_14379);
nand U14698 (N_14698,N_14180,N_14151);
xor U14699 (N_14699,N_14316,N_14322);
or U14700 (N_14700,N_14536,N_14663);
nand U14701 (N_14701,N_14693,N_14467);
nand U14702 (N_14702,N_14562,N_14649);
xor U14703 (N_14703,N_14610,N_14516);
or U14704 (N_14704,N_14637,N_14688);
or U14705 (N_14705,N_14561,N_14483);
nor U14706 (N_14706,N_14560,N_14667);
nand U14707 (N_14707,N_14611,N_14548);
nor U14708 (N_14708,N_14640,N_14435);
nor U14709 (N_14709,N_14574,N_14503);
or U14710 (N_14710,N_14659,N_14591);
nor U14711 (N_14711,N_14567,N_14454);
xnor U14712 (N_14712,N_14669,N_14477);
nand U14713 (N_14713,N_14513,N_14534);
or U14714 (N_14714,N_14401,N_14546);
nand U14715 (N_14715,N_14554,N_14539);
xnor U14716 (N_14716,N_14438,N_14564);
nor U14717 (N_14717,N_14422,N_14457);
nor U14718 (N_14718,N_14645,N_14405);
xor U14719 (N_14719,N_14577,N_14638);
nand U14720 (N_14720,N_14585,N_14698);
and U14721 (N_14721,N_14506,N_14650);
or U14722 (N_14722,N_14631,N_14686);
and U14723 (N_14723,N_14586,N_14528);
or U14724 (N_14724,N_14432,N_14572);
xnor U14725 (N_14725,N_14589,N_14532);
and U14726 (N_14726,N_14699,N_14488);
xnor U14727 (N_14727,N_14529,N_14458);
xor U14728 (N_14728,N_14406,N_14696);
and U14729 (N_14729,N_14552,N_14630);
nor U14730 (N_14730,N_14617,N_14531);
or U14731 (N_14731,N_14607,N_14485);
xor U14732 (N_14732,N_14523,N_14648);
xor U14733 (N_14733,N_14451,N_14547);
and U14734 (N_14734,N_14445,N_14495);
or U14735 (N_14735,N_14521,N_14537);
or U14736 (N_14736,N_14456,N_14480);
and U14737 (N_14737,N_14424,N_14605);
nand U14738 (N_14738,N_14555,N_14608);
nand U14739 (N_14739,N_14573,N_14520);
nor U14740 (N_14740,N_14690,N_14471);
and U14741 (N_14741,N_14668,N_14543);
xnor U14742 (N_14742,N_14412,N_14671);
and U14743 (N_14743,N_14404,N_14440);
nand U14744 (N_14744,N_14525,N_14545);
nor U14745 (N_14745,N_14580,N_14499);
xnor U14746 (N_14746,N_14428,N_14450);
or U14747 (N_14747,N_14694,N_14455);
and U14748 (N_14748,N_14655,N_14524);
nor U14749 (N_14749,N_14647,N_14675);
nand U14750 (N_14750,N_14615,N_14402);
or U14751 (N_14751,N_14502,N_14578);
nand U14752 (N_14752,N_14446,N_14596);
xor U14753 (N_14753,N_14621,N_14594);
or U14754 (N_14754,N_14590,N_14491);
and U14755 (N_14755,N_14481,N_14409);
xor U14756 (N_14756,N_14571,N_14504);
nand U14757 (N_14757,N_14408,N_14598);
nand U14758 (N_14758,N_14421,N_14437);
and U14759 (N_14759,N_14508,N_14470);
nor U14760 (N_14760,N_14544,N_14665);
or U14761 (N_14761,N_14417,N_14678);
nand U14762 (N_14762,N_14601,N_14697);
nor U14763 (N_14763,N_14622,N_14558);
and U14764 (N_14764,N_14430,N_14484);
and U14765 (N_14765,N_14627,N_14416);
nand U14766 (N_14766,N_14489,N_14660);
and U14767 (N_14767,N_14468,N_14582);
xor U14768 (N_14768,N_14498,N_14514);
xor U14769 (N_14769,N_14509,N_14486);
nor U14770 (N_14770,N_14602,N_14618);
xor U14771 (N_14771,N_14633,N_14670);
nand U14772 (N_14772,N_14527,N_14629);
and U14773 (N_14773,N_14654,N_14542);
nand U14774 (N_14774,N_14653,N_14579);
nand U14775 (N_14775,N_14526,N_14676);
nor U14776 (N_14776,N_14614,N_14553);
nor U14777 (N_14777,N_14419,N_14666);
nand U14778 (N_14778,N_14403,N_14415);
nor U14779 (N_14779,N_14444,N_14613);
or U14780 (N_14780,N_14680,N_14501);
and U14781 (N_14781,N_14448,N_14691);
and U14782 (N_14782,N_14535,N_14626);
nand U14783 (N_14783,N_14664,N_14533);
xor U14784 (N_14784,N_14541,N_14550);
and U14785 (N_14785,N_14496,N_14677);
nor U14786 (N_14786,N_14681,N_14494);
nor U14787 (N_14787,N_14563,N_14593);
and U14788 (N_14788,N_14619,N_14518);
and U14789 (N_14789,N_14413,N_14685);
or U14790 (N_14790,N_14587,N_14497);
nand U14791 (N_14791,N_14616,N_14466);
or U14792 (N_14792,N_14682,N_14657);
and U14793 (N_14793,N_14420,N_14464);
xnor U14794 (N_14794,N_14559,N_14433);
and U14795 (N_14795,N_14628,N_14434);
xnor U14796 (N_14796,N_14549,N_14636);
nand U14797 (N_14797,N_14538,N_14427);
and U14798 (N_14798,N_14505,N_14436);
and U14799 (N_14799,N_14687,N_14476);
and U14800 (N_14800,N_14465,N_14646);
nand U14801 (N_14801,N_14620,N_14644);
or U14802 (N_14802,N_14673,N_14684);
or U14803 (N_14803,N_14661,N_14418);
xor U14804 (N_14804,N_14500,N_14439);
or U14805 (N_14805,N_14592,N_14597);
nor U14806 (N_14806,N_14426,N_14606);
xnor U14807 (N_14807,N_14584,N_14568);
or U14808 (N_14808,N_14530,N_14623);
or U14809 (N_14809,N_14447,N_14425);
xor U14810 (N_14810,N_14557,N_14429);
nor U14811 (N_14811,N_14570,N_14609);
nand U14812 (N_14812,N_14603,N_14656);
nand U14813 (N_14813,N_14431,N_14479);
xnor U14814 (N_14814,N_14423,N_14474);
and U14815 (N_14815,N_14460,N_14566);
or U14816 (N_14816,N_14461,N_14487);
xor U14817 (N_14817,N_14452,N_14695);
nand U14818 (N_14818,N_14674,N_14463);
and U14819 (N_14819,N_14689,N_14642);
and U14820 (N_14820,N_14473,N_14510);
nand U14821 (N_14821,N_14595,N_14443);
and U14822 (N_14822,N_14540,N_14569);
and U14823 (N_14823,N_14639,N_14490);
nand U14824 (N_14824,N_14400,N_14459);
nor U14825 (N_14825,N_14641,N_14512);
nor U14826 (N_14826,N_14411,N_14515);
xnor U14827 (N_14827,N_14634,N_14462);
xor U14828 (N_14828,N_14492,N_14517);
or U14829 (N_14829,N_14672,N_14556);
xnor U14830 (N_14830,N_14522,N_14679);
nor U14831 (N_14831,N_14441,N_14600);
nand U14832 (N_14832,N_14511,N_14565);
and U14833 (N_14833,N_14414,N_14472);
xnor U14834 (N_14834,N_14442,N_14612);
nand U14835 (N_14835,N_14652,N_14581);
nand U14836 (N_14836,N_14453,N_14482);
and U14837 (N_14837,N_14692,N_14588);
xnor U14838 (N_14838,N_14683,N_14469);
xor U14839 (N_14839,N_14599,N_14662);
xor U14840 (N_14840,N_14632,N_14625);
or U14841 (N_14841,N_14583,N_14478);
or U14842 (N_14842,N_14551,N_14493);
nand U14843 (N_14843,N_14575,N_14643);
or U14844 (N_14844,N_14604,N_14475);
or U14845 (N_14845,N_14651,N_14507);
nand U14846 (N_14846,N_14624,N_14635);
nand U14847 (N_14847,N_14449,N_14410);
or U14848 (N_14848,N_14519,N_14407);
xor U14849 (N_14849,N_14576,N_14658);
nand U14850 (N_14850,N_14648,N_14627);
nor U14851 (N_14851,N_14406,N_14639);
and U14852 (N_14852,N_14614,N_14416);
or U14853 (N_14853,N_14463,N_14695);
and U14854 (N_14854,N_14437,N_14419);
xnor U14855 (N_14855,N_14617,N_14408);
nor U14856 (N_14856,N_14589,N_14594);
nor U14857 (N_14857,N_14506,N_14575);
or U14858 (N_14858,N_14673,N_14412);
xor U14859 (N_14859,N_14524,N_14641);
or U14860 (N_14860,N_14580,N_14670);
xnor U14861 (N_14861,N_14520,N_14448);
xnor U14862 (N_14862,N_14555,N_14460);
xor U14863 (N_14863,N_14515,N_14683);
xnor U14864 (N_14864,N_14424,N_14697);
or U14865 (N_14865,N_14527,N_14619);
and U14866 (N_14866,N_14628,N_14570);
nand U14867 (N_14867,N_14680,N_14440);
xnor U14868 (N_14868,N_14648,N_14492);
nor U14869 (N_14869,N_14458,N_14673);
or U14870 (N_14870,N_14502,N_14616);
or U14871 (N_14871,N_14681,N_14540);
or U14872 (N_14872,N_14589,N_14420);
nand U14873 (N_14873,N_14460,N_14539);
or U14874 (N_14874,N_14439,N_14446);
xnor U14875 (N_14875,N_14693,N_14660);
nand U14876 (N_14876,N_14562,N_14442);
and U14877 (N_14877,N_14501,N_14539);
xor U14878 (N_14878,N_14672,N_14683);
or U14879 (N_14879,N_14559,N_14486);
or U14880 (N_14880,N_14524,N_14491);
nand U14881 (N_14881,N_14577,N_14686);
nand U14882 (N_14882,N_14410,N_14521);
xor U14883 (N_14883,N_14523,N_14690);
xor U14884 (N_14884,N_14511,N_14623);
xnor U14885 (N_14885,N_14675,N_14407);
xor U14886 (N_14886,N_14646,N_14482);
nor U14887 (N_14887,N_14567,N_14496);
and U14888 (N_14888,N_14460,N_14590);
or U14889 (N_14889,N_14666,N_14630);
nand U14890 (N_14890,N_14619,N_14551);
nor U14891 (N_14891,N_14629,N_14550);
nor U14892 (N_14892,N_14691,N_14401);
nor U14893 (N_14893,N_14468,N_14490);
and U14894 (N_14894,N_14525,N_14678);
xnor U14895 (N_14895,N_14519,N_14485);
xnor U14896 (N_14896,N_14448,N_14619);
nand U14897 (N_14897,N_14510,N_14533);
and U14898 (N_14898,N_14692,N_14543);
nand U14899 (N_14899,N_14423,N_14524);
or U14900 (N_14900,N_14523,N_14662);
nor U14901 (N_14901,N_14462,N_14588);
xor U14902 (N_14902,N_14580,N_14532);
xnor U14903 (N_14903,N_14572,N_14676);
nor U14904 (N_14904,N_14616,N_14665);
or U14905 (N_14905,N_14510,N_14580);
and U14906 (N_14906,N_14693,N_14592);
nand U14907 (N_14907,N_14414,N_14592);
xnor U14908 (N_14908,N_14619,N_14627);
xnor U14909 (N_14909,N_14513,N_14673);
or U14910 (N_14910,N_14646,N_14540);
nand U14911 (N_14911,N_14638,N_14440);
nor U14912 (N_14912,N_14459,N_14594);
xnor U14913 (N_14913,N_14475,N_14653);
nor U14914 (N_14914,N_14480,N_14458);
xor U14915 (N_14915,N_14529,N_14596);
nor U14916 (N_14916,N_14498,N_14416);
nand U14917 (N_14917,N_14546,N_14499);
xnor U14918 (N_14918,N_14668,N_14675);
nor U14919 (N_14919,N_14660,N_14400);
or U14920 (N_14920,N_14622,N_14668);
xor U14921 (N_14921,N_14412,N_14574);
xnor U14922 (N_14922,N_14580,N_14482);
and U14923 (N_14923,N_14518,N_14558);
nor U14924 (N_14924,N_14528,N_14409);
or U14925 (N_14925,N_14434,N_14649);
nor U14926 (N_14926,N_14468,N_14646);
nor U14927 (N_14927,N_14589,N_14533);
nand U14928 (N_14928,N_14590,N_14674);
xor U14929 (N_14929,N_14450,N_14531);
nor U14930 (N_14930,N_14642,N_14425);
and U14931 (N_14931,N_14454,N_14472);
xor U14932 (N_14932,N_14595,N_14408);
and U14933 (N_14933,N_14588,N_14672);
xnor U14934 (N_14934,N_14649,N_14690);
or U14935 (N_14935,N_14481,N_14510);
or U14936 (N_14936,N_14488,N_14591);
nor U14937 (N_14937,N_14627,N_14555);
and U14938 (N_14938,N_14544,N_14588);
nand U14939 (N_14939,N_14445,N_14438);
nor U14940 (N_14940,N_14554,N_14551);
or U14941 (N_14941,N_14573,N_14481);
and U14942 (N_14942,N_14690,N_14634);
or U14943 (N_14943,N_14524,N_14649);
xnor U14944 (N_14944,N_14665,N_14663);
nor U14945 (N_14945,N_14656,N_14412);
and U14946 (N_14946,N_14614,N_14401);
nor U14947 (N_14947,N_14404,N_14510);
nand U14948 (N_14948,N_14677,N_14573);
xor U14949 (N_14949,N_14689,N_14514);
or U14950 (N_14950,N_14520,N_14550);
nand U14951 (N_14951,N_14504,N_14468);
or U14952 (N_14952,N_14451,N_14457);
nor U14953 (N_14953,N_14577,N_14651);
or U14954 (N_14954,N_14433,N_14430);
xnor U14955 (N_14955,N_14520,N_14685);
xor U14956 (N_14956,N_14612,N_14628);
and U14957 (N_14957,N_14435,N_14483);
xnor U14958 (N_14958,N_14414,N_14682);
nand U14959 (N_14959,N_14579,N_14465);
or U14960 (N_14960,N_14531,N_14457);
xor U14961 (N_14961,N_14409,N_14607);
nor U14962 (N_14962,N_14580,N_14572);
or U14963 (N_14963,N_14621,N_14659);
xnor U14964 (N_14964,N_14556,N_14652);
and U14965 (N_14965,N_14439,N_14657);
nand U14966 (N_14966,N_14446,N_14637);
nor U14967 (N_14967,N_14552,N_14696);
or U14968 (N_14968,N_14502,N_14457);
nor U14969 (N_14969,N_14606,N_14446);
or U14970 (N_14970,N_14691,N_14661);
and U14971 (N_14971,N_14426,N_14697);
nand U14972 (N_14972,N_14644,N_14633);
or U14973 (N_14973,N_14650,N_14545);
or U14974 (N_14974,N_14578,N_14637);
or U14975 (N_14975,N_14689,N_14660);
nor U14976 (N_14976,N_14645,N_14672);
nand U14977 (N_14977,N_14652,N_14501);
nand U14978 (N_14978,N_14699,N_14688);
or U14979 (N_14979,N_14514,N_14672);
or U14980 (N_14980,N_14647,N_14470);
and U14981 (N_14981,N_14695,N_14477);
and U14982 (N_14982,N_14410,N_14484);
or U14983 (N_14983,N_14661,N_14414);
and U14984 (N_14984,N_14476,N_14560);
nor U14985 (N_14985,N_14587,N_14457);
xnor U14986 (N_14986,N_14421,N_14470);
nor U14987 (N_14987,N_14682,N_14667);
nor U14988 (N_14988,N_14491,N_14679);
or U14989 (N_14989,N_14404,N_14548);
or U14990 (N_14990,N_14654,N_14552);
nand U14991 (N_14991,N_14459,N_14694);
xor U14992 (N_14992,N_14663,N_14637);
nor U14993 (N_14993,N_14459,N_14500);
nor U14994 (N_14994,N_14602,N_14682);
nor U14995 (N_14995,N_14460,N_14521);
nor U14996 (N_14996,N_14669,N_14529);
nand U14997 (N_14997,N_14627,N_14666);
nor U14998 (N_14998,N_14653,N_14422);
or U14999 (N_14999,N_14660,N_14471);
xnor UO_0 (O_0,N_14753,N_14715);
or UO_1 (O_1,N_14772,N_14947);
xor UO_2 (O_2,N_14730,N_14802);
nand UO_3 (O_3,N_14971,N_14993);
or UO_4 (O_4,N_14756,N_14892);
xor UO_5 (O_5,N_14758,N_14981);
nand UO_6 (O_6,N_14765,N_14934);
and UO_7 (O_7,N_14776,N_14903);
xor UO_8 (O_8,N_14705,N_14725);
nand UO_9 (O_9,N_14915,N_14724);
nand UO_10 (O_10,N_14840,N_14959);
nand UO_11 (O_11,N_14931,N_14864);
xnor UO_12 (O_12,N_14976,N_14963);
xnor UO_13 (O_13,N_14737,N_14755);
nor UO_14 (O_14,N_14708,N_14711);
and UO_15 (O_15,N_14768,N_14996);
nor UO_16 (O_16,N_14799,N_14906);
and UO_17 (O_17,N_14707,N_14740);
nor UO_18 (O_18,N_14932,N_14913);
xnor UO_19 (O_19,N_14872,N_14783);
xnor UO_20 (O_20,N_14822,N_14773);
or UO_21 (O_21,N_14882,N_14865);
and UO_22 (O_22,N_14806,N_14972);
and UO_23 (O_23,N_14874,N_14710);
nand UO_24 (O_24,N_14851,N_14798);
or UO_25 (O_25,N_14780,N_14941);
and UO_26 (O_26,N_14835,N_14933);
and UO_27 (O_27,N_14803,N_14842);
or UO_28 (O_28,N_14742,N_14973);
xor UO_29 (O_29,N_14916,N_14739);
nor UO_30 (O_30,N_14831,N_14863);
nor UO_31 (O_31,N_14791,N_14829);
and UO_32 (O_32,N_14837,N_14958);
xnor UO_33 (O_33,N_14808,N_14718);
nand UO_34 (O_34,N_14997,N_14905);
and UO_35 (O_35,N_14890,N_14969);
xnor UO_36 (O_36,N_14950,N_14716);
nand UO_37 (O_37,N_14746,N_14704);
and UO_38 (O_38,N_14952,N_14879);
and UO_39 (O_39,N_14717,N_14878);
nor UO_40 (O_40,N_14982,N_14804);
xor UO_41 (O_41,N_14914,N_14989);
or UO_42 (O_42,N_14848,N_14935);
nor UO_43 (O_43,N_14771,N_14819);
or UO_44 (O_44,N_14713,N_14985);
xor UO_45 (O_45,N_14857,N_14841);
and UO_46 (O_46,N_14861,N_14850);
or UO_47 (O_47,N_14991,N_14908);
nor UO_48 (O_48,N_14774,N_14983);
nand UO_49 (O_49,N_14902,N_14794);
or UO_50 (O_50,N_14800,N_14889);
nand UO_51 (O_51,N_14787,N_14812);
nor UO_52 (O_52,N_14723,N_14712);
or UO_53 (O_53,N_14979,N_14883);
or UO_54 (O_54,N_14929,N_14719);
nand UO_55 (O_55,N_14786,N_14960);
nor UO_56 (O_56,N_14954,N_14899);
nand UO_57 (O_57,N_14990,N_14834);
nor UO_58 (O_58,N_14894,N_14792);
xor UO_59 (O_59,N_14956,N_14923);
nand UO_60 (O_60,N_14757,N_14778);
or UO_61 (O_61,N_14828,N_14824);
or UO_62 (O_62,N_14953,N_14825);
nand UO_63 (O_63,N_14978,N_14826);
and UO_64 (O_64,N_14820,N_14832);
nor UO_65 (O_65,N_14980,N_14839);
xnor UO_66 (O_66,N_14790,N_14846);
nor UO_67 (O_67,N_14745,N_14927);
and UO_68 (O_68,N_14880,N_14873);
nand UO_69 (O_69,N_14911,N_14801);
xnor UO_70 (O_70,N_14856,N_14734);
nand UO_71 (O_71,N_14948,N_14944);
or UO_72 (O_72,N_14962,N_14917);
nand UO_73 (O_73,N_14830,N_14898);
xor UO_74 (O_74,N_14827,N_14881);
nor UO_75 (O_75,N_14924,N_14862);
and UO_76 (O_76,N_14930,N_14887);
and UO_77 (O_77,N_14775,N_14749);
and UO_78 (O_78,N_14919,N_14918);
or UO_79 (O_79,N_14759,N_14974);
nor UO_80 (O_80,N_14900,N_14965);
nor UO_81 (O_81,N_14984,N_14867);
nor UO_82 (O_82,N_14833,N_14714);
xnor UO_83 (O_83,N_14823,N_14738);
xor UO_84 (O_84,N_14907,N_14999);
xor UO_85 (O_85,N_14781,N_14858);
and UO_86 (O_86,N_14943,N_14946);
xnor UO_87 (O_87,N_14849,N_14870);
nand UO_88 (O_88,N_14987,N_14809);
or UO_89 (O_89,N_14843,N_14855);
xor UO_90 (O_90,N_14945,N_14810);
nor UO_91 (O_91,N_14942,N_14975);
nor UO_92 (O_92,N_14788,N_14817);
nor UO_93 (O_93,N_14928,N_14821);
xor UO_94 (O_94,N_14847,N_14875);
or UO_95 (O_95,N_14949,N_14744);
or UO_96 (O_96,N_14729,N_14709);
nor UO_97 (O_97,N_14761,N_14920);
nand UO_98 (O_98,N_14702,N_14995);
and UO_99 (O_99,N_14896,N_14937);
nor UO_100 (O_100,N_14836,N_14726);
xor UO_101 (O_101,N_14754,N_14922);
nor UO_102 (O_102,N_14992,N_14910);
xor UO_103 (O_103,N_14779,N_14904);
nand UO_104 (O_104,N_14891,N_14877);
and UO_105 (O_105,N_14720,N_14795);
xor UO_106 (O_106,N_14764,N_14722);
and UO_107 (O_107,N_14784,N_14860);
and UO_108 (O_108,N_14813,N_14763);
and UO_109 (O_109,N_14752,N_14853);
or UO_110 (O_110,N_14706,N_14951);
xor UO_111 (O_111,N_14701,N_14811);
and UO_112 (O_112,N_14888,N_14789);
xnor UO_113 (O_113,N_14727,N_14814);
nor UO_114 (O_114,N_14782,N_14748);
nor UO_115 (O_115,N_14869,N_14807);
and UO_116 (O_116,N_14735,N_14751);
and UO_117 (O_117,N_14838,N_14762);
nor UO_118 (O_118,N_14921,N_14741);
xnor UO_119 (O_119,N_14925,N_14961);
and UO_120 (O_120,N_14747,N_14866);
and UO_121 (O_121,N_14939,N_14893);
xnor UO_122 (O_122,N_14700,N_14728);
nand UO_123 (O_123,N_14721,N_14964);
nand UO_124 (O_124,N_14977,N_14743);
and UO_125 (O_125,N_14912,N_14970);
nand UO_126 (O_126,N_14868,N_14777);
and UO_127 (O_127,N_14793,N_14998);
nand UO_128 (O_128,N_14968,N_14854);
nand UO_129 (O_129,N_14816,N_14940);
and UO_130 (O_130,N_14845,N_14884);
or UO_131 (O_131,N_14769,N_14936);
and UO_132 (O_132,N_14703,N_14897);
or UO_133 (O_133,N_14967,N_14760);
nand UO_134 (O_134,N_14926,N_14994);
xnor UO_135 (O_135,N_14750,N_14886);
nor UO_136 (O_136,N_14957,N_14733);
nand UO_137 (O_137,N_14859,N_14909);
nand UO_138 (O_138,N_14732,N_14901);
and UO_139 (O_139,N_14785,N_14895);
xnor UO_140 (O_140,N_14966,N_14986);
nor UO_141 (O_141,N_14815,N_14955);
nand UO_142 (O_142,N_14885,N_14766);
xnor UO_143 (O_143,N_14736,N_14852);
and UO_144 (O_144,N_14871,N_14770);
and UO_145 (O_145,N_14797,N_14844);
and UO_146 (O_146,N_14988,N_14796);
xnor UO_147 (O_147,N_14767,N_14805);
or UO_148 (O_148,N_14731,N_14938);
and UO_149 (O_149,N_14876,N_14818);
nand UO_150 (O_150,N_14929,N_14836);
nor UO_151 (O_151,N_14965,N_14749);
and UO_152 (O_152,N_14768,N_14997);
nor UO_153 (O_153,N_14969,N_14727);
nand UO_154 (O_154,N_14817,N_14759);
or UO_155 (O_155,N_14898,N_14909);
nor UO_156 (O_156,N_14966,N_14772);
nor UO_157 (O_157,N_14870,N_14791);
xnor UO_158 (O_158,N_14765,N_14894);
or UO_159 (O_159,N_14776,N_14751);
nand UO_160 (O_160,N_14830,N_14783);
and UO_161 (O_161,N_14881,N_14722);
xnor UO_162 (O_162,N_14756,N_14786);
nor UO_163 (O_163,N_14754,N_14817);
nand UO_164 (O_164,N_14880,N_14751);
or UO_165 (O_165,N_14925,N_14759);
xnor UO_166 (O_166,N_14978,N_14842);
or UO_167 (O_167,N_14879,N_14999);
or UO_168 (O_168,N_14866,N_14778);
or UO_169 (O_169,N_14826,N_14957);
or UO_170 (O_170,N_14859,N_14817);
or UO_171 (O_171,N_14989,N_14867);
xor UO_172 (O_172,N_14799,N_14893);
or UO_173 (O_173,N_14833,N_14772);
nor UO_174 (O_174,N_14993,N_14952);
nor UO_175 (O_175,N_14940,N_14885);
nand UO_176 (O_176,N_14752,N_14827);
nand UO_177 (O_177,N_14901,N_14965);
nor UO_178 (O_178,N_14755,N_14817);
and UO_179 (O_179,N_14959,N_14859);
xor UO_180 (O_180,N_14867,N_14710);
xor UO_181 (O_181,N_14836,N_14710);
nor UO_182 (O_182,N_14831,N_14772);
xor UO_183 (O_183,N_14871,N_14702);
or UO_184 (O_184,N_14762,N_14912);
nand UO_185 (O_185,N_14731,N_14988);
xor UO_186 (O_186,N_14991,N_14726);
nand UO_187 (O_187,N_14951,N_14742);
and UO_188 (O_188,N_14717,N_14744);
nand UO_189 (O_189,N_14935,N_14902);
nor UO_190 (O_190,N_14971,N_14884);
xnor UO_191 (O_191,N_14702,N_14902);
xor UO_192 (O_192,N_14881,N_14724);
nand UO_193 (O_193,N_14899,N_14913);
xnor UO_194 (O_194,N_14764,N_14705);
xor UO_195 (O_195,N_14881,N_14789);
or UO_196 (O_196,N_14703,N_14828);
nor UO_197 (O_197,N_14923,N_14725);
and UO_198 (O_198,N_14862,N_14799);
nor UO_199 (O_199,N_14928,N_14892);
nand UO_200 (O_200,N_14724,N_14986);
nor UO_201 (O_201,N_14897,N_14957);
xnor UO_202 (O_202,N_14802,N_14954);
nand UO_203 (O_203,N_14869,N_14936);
or UO_204 (O_204,N_14883,N_14882);
or UO_205 (O_205,N_14794,N_14939);
xnor UO_206 (O_206,N_14752,N_14766);
nand UO_207 (O_207,N_14731,N_14715);
nor UO_208 (O_208,N_14861,N_14749);
or UO_209 (O_209,N_14886,N_14870);
xnor UO_210 (O_210,N_14757,N_14998);
and UO_211 (O_211,N_14751,N_14872);
nand UO_212 (O_212,N_14914,N_14738);
nor UO_213 (O_213,N_14701,N_14741);
nand UO_214 (O_214,N_14902,N_14900);
and UO_215 (O_215,N_14780,N_14770);
or UO_216 (O_216,N_14962,N_14944);
xnor UO_217 (O_217,N_14779,N_14906);
and UO_218 (O_218,N_14856,N_14798);
and UO_219 (O_219,N_14864,N_14995);
and UO_220 (O_220,N_14888,N_14998);
or UO_221 (O_221,N_14715,N_14943);
or UO_222 (O_222,N_14763,N_14725);
and UO_223 (O_223,N_14957,N_14744);
and UO_224 (O_224,N_14742,N_14972);
and UO_225 (O_225,N_14718,N_14738);
nand UO_226 (O_226,N_14917,N_14711);
and UO_227 (O_227,N_14909,N_14733);
nor UO_228 (O_228,N_14921,N_14903);
nand UO_229 (O_229,N_14898,N_14827);
and UO_230 (O_230,N_14940,N_14763);
nand UO_231 (O_231,N_14788,N_14915);
or UO_232 (O_232,N_14837,N_14878);
xnor UO_233 (O_233,N_14951,N_14899);
nand UO_234 (O_234,N_14899,N_14750);
and UO_235 (O_235,N_14796,N_14832);
xnor UO_236 (O_236,N_14764,N_14961);
or UO_237 (O_237,N_14933,N_14801);
nand UO_238 (O_238,N_14896,N_14753);
nand UO_239 (O_239,N_14891,N_14929);
xor UO_240 (O_240,N_14766,N_14822);
xor UO_241 (O_241,N_14716,N_14702);
and UO_242 (O_242,N_14777,N_14948);
nand UO_243 (O_243,N_14981,N_14850);
nor UO_244 (O_244,N_14808,N_14939);
or UO_245 (O_245,N_14856,N_14703);
xor UO_246 (O_246,N_14814,N_14867);
nand UO_247 (O_247,N_14953,N_14799);
or UO_248 (O_248,N_14706,N_14852);
nand UO_249 (O_249,N_14946,N_14983);
or UO_250 (O_250,N_14740,N_14927);
nor UO_251 (O_251,N_14864,N_14830);
nor UO_252 (O_252,N_14719,N_14875);
nor UO_253 (O_253,N_14938,N_14932);
nor UO_254 (O_254,N_14980,N_14948);
nand UO_255 (O_255,N_14792,N_14992);
or UO_256 (O_256,N_14970,N_14776);
nor UO_257 (O_257,N_14895,N_14900);
or UO_258 (O_258,N_14932,N_14720);
nor UO_259 (O_259,N_14853,N_14830);
xnor UO_260 (O_260,N_14879,N_14980);
nand UO_261 (O_261,N_14910,N_14763);
nor UO_262 (O_262,N_14997,N_14868);
xnor UO_263 (O_263,N_14775,N_14846);
xor UO_264 (O_264,N_14810,N_14979);
nand UO_265 (O_265,N_14857,N_14820);
xor UO_266 (O_266,N_14924,N_14779);
xnor UO_267 (O_267,N_14871,N_14815);
xor UO_268 (O_268,N_14879,N_14814);
xnor UO_269 (O_269,N_14736,N_14988);
nand UO_270 (O_270,N_14896,N_14810);
and UO_271 (O_271,N_14980,N_14714);
nand UO_272 (O_272,N_14762,N_14768);
or UO_273 (O_273,N_14818,N_14845);
or UO_274 (O_274,N_14853,N_14832);
and UO_275 (O_275,N_14964,N_14815);
nor UO_276 (O_276,N_14951,N_14715);
xnor UO_277 (O_277,N_14816,N_14910);
xnor UO_278 (O_278,N_14855,N_14929);
and UO_279 (O_279,N_14986,N_14781);
nand UO_280 (O_280,N_14735,N_14829);
nor UO_281 (O_281,N_14990,N_14711);
nand UO_282 (O_282,N_14926,N_14787);
nand UO_283 (O_283,N_14958,N_14729);
xnor UO_284 (O_284,N_14740,N_14892);
or UO_285 (O_285,N_14796,N_14803);
or UO_286 (O_286,N_14714,N_14929);
xnor UO_287 (O_287,N_14765,N_14799);
nand UO_288 (O_288,N_14878,N_14702);
nand UO_289 (O_289,N_14760,N_14719);
nor UO_290 (O_290,N_14986,N_14985);
xnor UO_291 (O_291,N_14851,N_14980);
and UO_292 (O_292,N_14864,N_14726);
nand UO_293 (O_293,N_14836,N_14807);
xor UO_294 (O_294,N_14901,N_14912);
or UO_295 (O_295,N_14823,N_14880);
or UO_296 (O_296,N_14825,N_14815);
or UO_297 (O_297,N_14769,N_14840);
or UO_298 (O_298,N_14726,N_14975);
nand UO_299 (O_299,N_14827,N_14968);
nor UO_300 (O_300,N_14938,N_14904);
or UO_301 (O_301,N_14867,N_14929);
xnor UO_302 (O_302,N_14908,N_14923);
and UO_303 (O_303,N_14946,N_14937);
nor UO_304 (O_304,N_14953,N_14891);
or UO_305 (O_305,N_14851,N_14895);
xnor UO_306 (O_306,N_14869,N_14772);
nand UO_307 (O_307,N_14835,N_14737);
and UO_308 (O_308,N_14845,N_14979);
nand UO_309 (O_309,N_14707,N_14772);
or UO_310 (O_310,N_14977,N_14869);
nor UO_311 (O_311,N_14718,N_14858);
nand UO_312 (O_312,N_14865,N_14898);
nand UO_313 (O_313,N_14910,N_14972);
nand UO_314 (O_314,N_14924,N_14793);
nand UO_315 (O_315,N_14847,N_14811);
or UO_316 (O_316,N_14855,N_14999);
or UO_317 (O_317,N_14870,N_14892);
or UO_318 (O_318,N_14932,N_14725);
or UO_319 (O_319,N_14777,N_14831);
nor UO_320 (O_320,N_14717,N_14805);
xor UO_321 (O_321,N_14844,N_14788);
or UO_322 (O_322,N_14777,N_14908);
nor UO_323 (O_323,N_14906,N_14875);
xor UO_324 (O_324,N_14978,N_14969);
and UO_325 (O_325,N_14736,N_14761);
and UO_326 (O_326,N_14769,N_14782);
nand UO_327 (O_327,N_14907,N_14988);
nand UO_328 (O_328,N_14853,N_14781);
or UO_329 (O_329,N_14902,N_14759);
nor UO_330 (O_330,N_14808,N_14817);
nor UO_331 (O_331,N_14993,N_14787);
nand UO_332 (O_332,N_14802,N_14868);
or UO_333 (O_333,N_14842,N_14775);
or UO_334 (O_334,N_14849,N_14757);
nor UO_335 (O_335,N_14741,N_14869);
nand UO_336 (O_336,N_14803,N_14786);
nand UO_337 (O_337,N_14773,N_14790);
or UO_338 (O_338,N_14885,N_14712);
xor UO_339 (O_339,N_14943,N_14739);
xnor UO_340 (O_340,N_14750,N_14961);
or UO_341 (O_341,N_14832,N_14790);
xor UO_342 (O_342,N_14874,N_14867);
xnor UO_343 (O_343,N_14730,N_14772);
xnor UO_344 (O_344,N_14959,N_14719);
and UO_345 (O_345,N_14767,N_14713);
nand UO_346 (O_346,N_14996,N_14753);
xor UO_347 (O_347,N_14863,N_14956);
nand UO_348 (O_348,N_14891,N_14713);
nor UO_349 (O_349,N_14973,N_14832);
nor UO_350 (O_350,N_14754,N_14877);
nor UO_351 (O_351,N_14757,N_14846);
or UO_352 (O_352,N_14753,N_14945);
and UO_353 (O_353,N_14898,N_14922);
nor UO_354 (O_354,N_14959,N_14858);
xnor UO_355 (O_355,N_14774,N_14925);
xor UO_356 (O_356,N_14834,N_14932);
and UO_357 (O_357,N_14835,N_14941);
nor UO_358 (O_358,N_14722,N_14889);
xor UO_359 (O_359,N_14705,N_14758);
xor UO_360 (O_360,N_14826,N_14800);
and UO_361 (O_361,N_14787,N_14775);
and UO_362 (O_362,N_14847,N_14805);
nor UO_363 (O_363,N_14936,N_14891);
or UO_364 (O_364,N_14747,N_14915);
nand UO_365 (O_365,N_14959,N_14870);
nor UO_366 (O_366,N_14837,N_14747);
nand UO_367 (O_367,N_14776,N_14924);
xor UO_368 (O_368,N_14927,N_14706);
and UO_369 (O_369,N_14891,N_14910);
or UO_370 (O_370,N_14926,N_14789);
nand UO_371 (O_371,N_14851,N_14716);
or UO_372 (O_372,N_14719,N_14954);
nand UO_373 (O_373,N_14913,N_14883);
xor UO_374 (O_374,N_14821,N_14721);
nor UO_375 (O_375,N_14807,N_14984);
nand UO_376 (O_376,N_14964,N_14974);
nand UO_377 (O_377,N_14706,N_14963);
nand UO_378 (O_378,N_14738,N_14917);
nand UO_379 (O_379,N_14883,N_14811);
and UO_380 (O_380,N_14795,N_14747);
xor UO_381 (O_381,N_14794,N_14957);
and UO_382 (O_382,N_14924,N_14811);
nor UO_383 (O_383,N_14881,N_14898);
or UO_384 (O_384,N_14949,N_14978);
xnor UO_385 (O_385,N_14959,N_14876);
and UO_386 (O_386,N_14748,N_14815);
nand UO_387 (O_387,N_14722,N_14820);
or UO_388 (O_388,N_14971,N_14867);
nand UO_389 (O_389,N_14987,N_14988);
xor UO_390 (O_390,N_14831,N_14729);
and UO_391 (O_391,N_14863,N_14747);
and UO_392 (O_392,N_14889,N_14934);
or UO_393 (O_393,N_14760,N_14780);
nor UO_394 (O_394,N_14719,N_14825);
nor UO_395 (O_395,N_14862,N_14752);
and UO_396 (O_396,N_14881,N_14763);
or UO_397 (O_397,N_14795,N_14758);
and UO_398 (O_398,N_14757,N_14925);
xor UO_399 (O_399,N_14852,N_14949);
nor UO_400 (O_400,N_14847,N_14822);
xor UO_401 (O_401,N_14849,N_14958);
xnor UO_402 (O_402,N_14749,N_14764);
and UO_403 (O_403,N_14714,N_14880);
nor UO_404 (O_404,N_14987,N_14921);
and UO_405 (O_405,N_14990,N_14995);
nor UO_406 (O_406,N_14900,N_14817);
nor UO_407 (O_407,N_14778,N_14726);
nor UO_408 (O_408,N_14837,N_14737);
nor UO_409 (O_409,N_14984,N_14912);
nor UO_410 (O_410,N_14786,N_14843);
xor UO_411 (O_411,N_14812,N_14882);
and UO_412 (O_412,N_14805,N_14949);
nor UO_413 (O_413,N_14985,N_14780);
or UO_414 (O_414,N_14999,N_14871);
and UO_415 (O_415,N_14972,N_14892);
xnor UO_416 (O_416,N_14729,N_14875);
nor UO_417 (O_417,N_14987,N_14994);
nor UO_418 (O_418,N_14822,N_14865);
nor UO_419 (O_419,N_14739,N_14767);
and UO_420 (O_420,N_14888,N_14922);
and UO_421 (O_421,N_14980,N_14987);
nand UO_422 (O_422,N_14935,N_14932);
or UO_423 (O_423,N_14762,N_14754);
nand UO_424 (O_424,N_14853,N_14759);
nand UO_425 (O_425,N_14993,N_14843);
xnor UO_426 (O_426,N_14815,N_14706);
nor UO_427 (O_427,N_14708,N_14760);
xnor UO_428 (O_428,N_14864,N_14891);
and UO_429 (O_429,N_14865,N_14989);
nor UO_430 (O_430,N_14738,N_14869);
xnor UO_431 (O_431,N_14883,N_14784);
and UO_432 (O_432,N_14759,N_14890);
xnor UO_433 (O_433,N_14845,N_14928);
xor UO_434 (O_434,N_14759,N_14947);
xor UO_435 (O_435,N_14972,N_14948);
nand UO_436 (O_436,N_14930,N_14990);
and UO_437 (O_437,N_14908,N_14956);
xnor UO_438 (O_438,N_14759,N_14745);
nand UO_439 (O_439,N_14778,N_14889);
xor UO_440 (O_440,N_14754,N_14806);
or UO_441 (O_441,N_14704,N_14957);
or UO_442 (O_442,N_14926,N_14793);
nand UO_443 (O_443,N_14955,N_14974);
nand UO_444 (O_444,N_14712,N_14904);
xor UO_445 (O_445,N_14921,N_14705);
xor UO_446 (O_446,N_14973,N_14951);
nand UO_447 (O_447,N_14845,N_14703);
or UO_448 (O_448,N_14760,N_14776);
xor UO_449 (O_449,N_14962,N_14721);
nand UO_450 (O_450,N_14713,N_14703);
xnor UO_451 (O_451,N_14830,N_14837);
nand UO_452 (O_452,N_14852,N_14899);
xor UO_453 (O_453,N_14943,N_14766);
nand UO_454 (O_454,N_14781,N_14832);
nor UO_455 (O_455,N_14889,N_14835);
nor UO_456 (O_456,N_14905,N_14763);
or UO_457 (O_457,N_14757,N_14801);
and UO_458 (O_458,N_14759,N_14798);
nor UO_459 (O_459,N_14812,N_14820);
nor UO_460 (O_460,N_14751,N_14949);
or UO_461 (O_461,N_14937,N_14809);
xor UO_462 (O_462,N_14937,N_14709);
nor UO_463 (O_463,N_14918,N_14860);
and UO_464 (O_464,N_14949,N_14787);
nor UO_465 (O_465,N_14702,N_14928);
xor UO_466 (O_466,N_14707,N_14832);
xor UO_467 (O_467,N_14771,N_14986);
nor UO_468 (O_468,N_14851,N_14897);
nand UO_469 (O_469,N_14804,N_14820);
nand UO_470 (O_470,N_14837,N_14782);
nor UO_471 (O_471,N_14803,N_14715);
and UO_472 (O_472,N_14703,N_14872);
nand UO_473 (O_473,N_14857,N_14715);
xor UO_474 (O_474,N_14956,N_14828);
xnor UO_475 (O_475,N_14838,N_14936);
xnor UO_476 (O_476,N_14956,N_14798);
or UO_477 (O_477,N_14949,N_14867);
and UO_478 (O_478,N_14937,N_14825);
nor UO_479 (O_479,N_14901,N_14930);
or UO_480 (O_480,N_14770,N_14838);
nor UO_481 (O_481,N_14853,N_14847);
nor UO_482 (O_482,N_14784,N_14787);
xor UO_483 (O_483,N_14784,N_14949);
or UO_484 (O_484,N_14914,N_14841);
nor UO_485 (O_485,N_14869,N_14792);
or UO_486 (O_486,N_14791,N_14780);
xnor UO_487 (O_487,N_14927,N_14888);
and UO_488 (O_488,N_14900,N_14898);
nor UO_489 (O_489,N_14833,N_14781);
and UO_490 (O_490,N_14882,N_14778);
nand UO_491 (O_491,N_14701,N_14732);
or UO_492 (O_492,N_14898,N_14994);
xnor UO_493 (O_493,N_14736,N_14804);
nor UO_494 (O_494,N_14886,N_14986);
or UO_495 (O_495,N_14904,N_14968);
and UO_496 (O_496,N_14771,N_14827);
nand UO_497 (O_497,N_14763,N_14846);
nand UO_498 (O_498,N_14941,N_14777);
or UO_499 (O_499,N_14753,N_14778);
and UO_500 (O_500,N_14789,N_14808);
nor UO_501 (O_501,N_14955,N_14777);
nand UO_502 (O_502,N_14898,N_14783);
and UO_503 (O_503,N_14751,N_14989);
nor UO_504 (O_504,N_14955,N_14830);
nand UO_505 (O_505,N_14843,N_14890);
xnor UO_506 (O_506,N_14715,N_14908);
nor UO_507 (O_507,N_14839,N_14996);
nand UO_508 (O_508,N_14982,N_14818);
nor UO_509 (O_509,N_14918,N_14758);
and UO_510 (O_510,N_14869,N_14710);
xor UO_511 (O_511,N_14831,N_14846);
nor UO_512 (O_512,N_14721,N_14803);
nor UO_513 (O_513,N_14923,N_14967);
xnor UO_514 (O_514,N_14971,N_14776);
or UO_515 (O_515,N_14869,N_14824);
or UO_516 (O_516,N_14933,N_14934);
or UO_517 (O_517,N_14791,N_14960);
nor UO_518 (O_518,N_14940,N_14907);
nor UO_519 (O_519,N_14917,N_14967);
xor UO_520 (O_520,N_14820,N_14991);
nand UO_521 (O_521,N_14890,N_14902);
or UO_522 (O_522,N_14803,N_14802);
and UO_523 (O_523,N_14822,N_14844);
nand UO_524 (O_524,N_14874,N_14836);
or UO_525 (O_525,N_14745,N_14895);
and UO_526 (O_526,N_14817,N_14965);
or UO_527 (O_527,N_14932,N_14793);
or UO_528 (O_528,N_14911,N_14920);
or UO_529 (O_529,N_14907,N_14983);
nor UO_530 (O_530,N_14805,N_14798);
xor UO_531 (O_531,N_14881,N_14948);
xnor UO_532 (O_532,N_14969,N_14875);
nor UO_533 (O_533,N_14750,N_14716);
or UO_534 (O_534,N_14918,N_14916);
or UO_535 (O_535,N_14772,N_14967);
or UO_536 (O_536,N_14914,N_14876);
or UO_537 (O_537,N_14790,N_14874);
xnor UO_538 (O_538,N_14844,N_14842);
and UO_539 (O_539,N_14931,N_14854);
nand UO_540 (O_540,N_14881,N_14762);
nor UO_541 (O_541,N_14796,N_14718);
xnor UO_542 (O_542,N_14784,N_14999);
nor UO_543 (O_543,N_14858,N_14845);
or UO_544 (O_544,N_14804,N_14971);
xnor UO_545 (O_545,N_14734,N_14719);
nand UO_546 (O_546,N_14793,N_14730);
nand UO_547 (O_547,N_14752,N_14843);
and UO_548 (O_548,N_14729,N_14949);
nor UO_549 (O_549,N_14953,N_14967);
nand UO_550 (O_550,N_14961,N_14810);
nand UO_551 (O_551,N_14950,N_14799);
and UO_552 (O_552,N_14830,N_14961);
or UO_553 (O_553,N_14777,N_14715);
or UO_554 (O_554,N_14764,N_14896);
nand UO_555 (O_555,N_14776,N_14758);
or UO_556 (O_556,N_14987,N_14900);
xnor UO_557 (O_557,N_14902,N_14833);
or UO_558 (O_558,N_14931,N_14882);
xnor UO_559 (O_559,N_14802,N_14761);
xor UO_560 (O_560,N_14792,N_14860);
and UO_561 (O_561,N_14902,N_14924);
xnor UO_562 (O_562,N_14921,N_14792);
nor UO_563 (O_563,N_14752,N_14848);
and UO_564 (O_564,N_14991,N_14719);
xor UO_565 (O_565,N_14801,N_14722);
or UO_566 (O_566,N_14923,N_14802);
or UO_567 (O_567,N_14960,N_14875);
nor UO_568 (O_568,N_14708,N_14870);
and UO_569 (O_569,N_14774,N_14867);
nor UO_570 (O_570,N_14745,N_14718);
and UO_571 (O_571,N_14705,N_14722);
or UO_572 (O_572,N_14876,N_14946);
or UO_573 (O_573,N_14963,N_14727);
nand UO_574 (O_574,N_14929,N_14772);
or UO_575 (O_575,N_14749,N_14860);
and UO_576 (O_576,N_14790,N_14836);
xor UO_577 (O_577,N_14968,N_14924);
nand UO_578 (O_578,N_14916,N_14919);
or UO_579 (O_579,N_14849,N_14919);
xnor UO_580 (O_580,N_14796,N_14841);
and UO_581 (O_581,N_14714,N_14976);
xor UO_582 (O_582,N_14853,N_14913);
nand UO_583 (O_583,N_14952,N_14925);
nor UO_584 (O_584,N_14963,N_14957);
nand UO_585 (O_585,N_14757,N_14800);
nand UO_586 (O_586,N_14984,N_14702);
or UO_587 (O_587,N_14847,N_14828);
nand UO_588 (O_588,N_14825,N_14847);
or UO_589 (O_589,N_14772,N_14839);
or UO_590 (O_590,N_14945,N_14783);
xnor UO_591 (O_591,N_14993,N_14857);
or UO_592 (O_592,N_14827,N_14914);
or UO_593 (O_593,N_14874,N_14995);
nand UO_594 (O_594,N_14878,N_14751);
xnor UO_595 (O_595,N_14726,N_14894);
xnor UO_596 (O_596,N_14758,N_14751);
xor UO_597 (O_597,N_14860,N_14808);
nor UO_598 (O_598,N_14764,N_14700);
or UO_599 (O_599,N_14725,N_14846);
nand UO_600 (O_600,N_14753,N_14772);
xnor UO_601 (O_601,N_14752,N_14929);
nand UO_602 (O_602,N_14999,N_14708);
and UO_603 (O_603,N_14856,N_14877);
nor UO_604 (O_604,N_14802,N_14793);
or UO_605 (O_605,N_14926,N_14740);
nor UO_606 (O_606,N_14923,N_14867);
or UO_607 (O_607,N_14791,N_14987);
or UO_608 (O_608,N_14763,N_14850);
or UO_609 (O_609,N_14908,N_14769);
nor UO_610 (O_610,N_14971,N_14874);
xor UO_611 (O_611,N_14962,N_14754);
xnor UO_612 (O_612,N_14720,N_14702);
or UO_613 (O_613,N_14830,N_14944);
nand UO_614 (O_614,N_14820,N_14968);
or UO_615 (O_615,N_14767,N_14730);
xor UO_616 (O_616,N_14895,N_14905);
nor UO_617 (O_617,N_14917,N_14861);
and UO_618 (O_618,N_14995,N_14903);
nand UO_619 (O_619,N_14959,N_14931);
nand UO_620 (O_620,N_14771,N_14804);
nand UO_621 (O_621,N_14946,N_14733);
or UO_622 (O_622,N_14783,N_14916);
nand UO_623 (O_623,N_14705,N_14805);
nor UO_624 (O_624,N_14950,N_14826);
or UO_625 (O_625,N_14966,N_14780);
and UO_626 (O_626,N_14894,N_14897);
or UO_627 (O_627,N_14999,N_14997);
xnor UO_628 (O_628,N_14863,N_14964);
xnor UO_629 (O_629,N_14950,N_14798);
or UO_630 (O_630,N_14711,N_14740);
xor UO_631 (O_631,N_14787,N_14761);
nand UO_632 (O_632,N_14822,N_14743);
or UO_633 (O_633,N_14718,N_14960);
and UO_634 (O_634,N_14814,N_14856);
nor UO_635 (O_635,N_14927,N_14774);
or UO_636 (O_636,N_14804,N_14824);
or UO_637 (O_637,N_14990,N_14745);
and UO_638 (O_638,N_14703,N_14782);
nand UO_639 (O_639,N_14797,N_14888);
or UO_640 (O_640,N_14740,N_14918);
nand UO_641 (O_641,N_14793,N_14717);
xnor UO_642 (O_642,N_14701,N_14904);
xor UO_643 (O_643,N_14930,N_14902);
or UO_644 (O_644,N_14902,N_14745);
nand UO_645 (O_645,N_14947,N_14822);
nand UO_646 (O_646,N_14731,N_14728);
xnor UO_647 (O_647,N_14776,N_14761);
and UO_648 (O_648,N_14982,N_14701);
xor UO_649 (O_649,N_14918,N_14830);
nand UO_650 (O_650,N_14830,N_14785);
and UO_651 (O_651,N_14771,N_14783);
nand UO_652 (O_652,N_14838,N_14758);
nand UO_653 (O_653,N_14713,N_14778);
nand UO_654 (O_654,N_14883,N_14859);
and UO_655 (O_655,N_14764,N_14995);
or UO_656 (O_656,N_14844,N_14780);
xnor UO_657 (O_657,N_14724,N_14813);
nand UO_658 (O_658,N_14731,N_14930);
or UO_659 (O_659,N_14718,N_14845);
nand UO_660 (O_660,N_14965,N_14806);
and UO_661 (O_661,N_14861,N_14950);
or UO_662 (O_662,N_14988,N_14784);
nor UO_663 (O_663,N_14752,N_14841);
xor UO_664 (O_664,N_14903,N_14802);
nand UO_665 (O_665,N_14705,N_14897);
nand UO_666 (O_666,N_14952,N_14838);
or UO_667 (O_667,N_14814,N_14852);
nand UO_668 (O_668,N_14961,N_14880);
or UO_669 (O_669,N_14951,N_14771);
xnor UO_670 (O_670,N_14999,N_14705);
nor UO_671 (O_671,N_14982,N_14795);
and UO_672 (O_672,N_14755,N_14938);
nor UO_673 (O_673,N_14941,N_14914);
nand UO_674 (O_674,N_14906,N_14762);
xor UO_675 (O_675,N_14766,N_14772);
nor UO_676 (O_676,N_14804,N_14843);
xor UO_677 (O_677,N_14911,N_14953);
nand UO_678 (O_678,N_14796,N_14914);
and UO_679 (O_679,N_14861,N_14938);
or UO_680 (O_680,N_14985,N_14944);
and UO_681 (O_681,N_14827,N_14769);
nand UO_682 (O_682,N_14728,N_14858);
nand UO_683 (O_683,N_14722,N_14836);
xor UO_684 (O_684,N_14796,N_14905);
nand UO_685 (O_685,N_14736,N_14872);
and UO_686 (O_686,N_14980,N_14810);
and UO_687 (O_687,N_14960,N_14899);
and UO_688 (O_688,N_14815,N_14838);
nor UO_689 (O_689,N_14819,N_14865);
or UO_690 (O_690,N_14740,N_14787);
and UO_691 (O_691,N_14991,N_14858);
or UO_692 (O_692,N_14792,N_14732);
nor UO_693 (O_693,N_14873,N_14927);
xnor UO_694 (O_694,N_14795,N_14752);
nor UO_695 (O_695,N_14857,N_14972);
nand UO_696 (O_696,N_14938,N_14703);
nand UO_697 (O_697,N_14730,N_14710);
or UO_698 (O_698,N_14749,N_14721);
and UO_699 (O_699,N_14701,N_14840);
nor UO_700 (O_700,N_14784,N_14866);
and UO_701 (O_701,N_14711,N_14808);
nand UO_702 (O_702,N_14942,N_14841);
xnor UO_703 (O_703,N_14898,N_14805);
and UO_704 (O_704,N_14985,N_14935);
nand UO_705 (O_705,N_14875,N_14790);
nor UO_706 (O_706,N_14934,N_14929);
nand UO_707 (O_707,N_14802,N_14762);
or UO_708 (O_708,N_14946,N_14803);
xor UO_709 (O_709,N_14981,N_14769);
and UO_710 (O_710,N_14722,N_14726);
and UO_711 (O_711,N_14845,N_14743);
or UO_712 (O_712,N_14782,N_14932);
xor UO_713 (O_713,N_14940,N_14903);
and UO_714 (O_714,N_14822,N_14912);
or UO_715 (O_715,N_14818,N_14897);
nand UO_716 (O_716,N_14897,N_14939);
nand UO_717 (O_717,N_14849,N_14949);
or UO_718 (O_718,N_14774,N_14817);
nand UO_719 (O_719,N_14929,N_14989);
and UO_720 (O_720,N_14937,N_14978);
and UO_721 (O_721,N_14774,N_14960);
and UO_722 (O_722,N_14797,N_14979);
nor UO_723 (O_723,N_14766,N_14798);
and UO_724 (O_724,N_14925,N_14881);
and UO_725 (O_725,N_14988,N_14709);
and UO_726 (O_726,N_14940,N_14843);
nor UO_727 (O_727,N_14805,N_14727);
nand UO_728 (O_728,N_14867,N_14910);
nor UO_729 (O_729,N_14910,N_14739);
and UO_730 (O_730,N_14768,N_14704);
and UO_731 (O_731,N_14836,N_14972);
nand UO_732 (O_732,N_14787,N_14731);
or UO_733 (O_733,N_14831,N_14870);
nor UO_734 (O_734,N_14719,N_14771);
and UO_735 (O_735,N_14819,N_14904);
nand UO_736 (O_736,N_14864,N_14967);
nor UO_737 (O_737,N_14802,N_14772);
nand UO_738 (O_738,N_14753,N_14933);
xor UO_739 (O_739,N_14707,N_14953);
xnor UO_740 (O_740,N_14776,N_14734);
and UO_741 (O_741,N_14718,N_14860);
nor UO_742 (O_742,N_14906,N_14719);
nor UO_743 (O_743,N_14709,N_14985);
and UO_744 (O_744,N_14723,N_14962);
or UO_745 (O_745,N_14805,N_14766);
xor UO_746 (O_746,N_14946,N_14738);
nor UO_747 (O_747,N_14724,N_14925);
and UO_748 (O_748,N_14786,N_14789);
nand UO_749 (O_749,N_14795,N_14915);
xnor UO_750 (O_750,N_14938,N_14720);
nand UO_751 (O_751,N_14968,N_14776);
xnor UO_752 (O_752,N_14969,N_14928);
or UO_753 (O_753,N_14860,N_14804);
nand UO_754 (O_754,N_14930,N_14926);
nor UO_755 (O_755,N_14879,N_14947);
nand UO_756 (O_756,N_14982,N_14940);
nand UO_757 (O_757,N_14903,N_14853);
nor UO_758 (O_758,N_14727,N_14831);
xor UO_759 (O_759,N_14861,N_14916);
nand UO_760 (O_760,N_14901,N_14703);
nor UO_761 (O_761,N_14720,N_14731);
or UO_762 (O_762,N_14947,N_14942);
nor UO_763 (O_763,N_14847,N_14738);
and UO_764 (O_764,N_14936,N_14972);
nor UO_765 (O_765,N_14712,N_14887);
nor UO_766 (O_766,N_14788,N_14702);
xnor UO_767 (O_767,N_14933,N_14841);
nor UO_768 (O_768,N_14748,N_14978);
xor UO_769 (O_769,N_14876,N_14960);
nor UO_770 (O_770,N_14882,N_14962);
xnor UO_771 (O_771,N_14895,N_14790);
xor UO_772 (O_772,N_14750,N_14732);
nand UO_773 (O_773,N_14750,N_14908);
nand UO_774 (O_774,N_14868,N_14873);
or UO_775 (O_775,N_14927,N_14945);
xor UO_776 (O_776,N_14896,N_14828);
and UO_777 (O_777,N_14841,N_14734);
xnor UO_778 (O_778,N_14952,N_14932);
xor UO_779 (O_779,N_14959,N_14852);
xnor UO_780 (O_780,N_14871,N_14957);
xor UO_781 (O_781,N_14948,N_14707);
xnor UO_782 (O_782,N_14835,N_14736);
nand UO_783 (O_783,N_14759,N_14791);
nor UO_784 (O_784,N_14910,N_14885);
nand UO_785 (O_785,N_14938,N_14798);
nand UO_786 (O_786,N_14741,N_14713);
and UO_787 (O_787,N_14771,N_14935);
nor UO_788 (O_788,N_14899,N_14971);
nor UO_789 (O_789,N_14843,N_14772);
or UO_790 (O_790,N_14905,N_14897);
and UO_791 (O_791,N_14793,N_14864);
nand UO_792 (O_792,N_14773,N_14802);
xnor UO_793 (O_793,N_14923,N_14918);
nand UO_794 (O_794,N_14975,N_14947);
xnor UO_795 (O_795,N_14898,N_14983);
xnor UO_796 (O_796,N_14710,N_14797);
nor UO_797 (O_797,N_14986,N_14833);
nor UO_798 (O_798,N_14876,N_14925);
nand UO_799 (O_799,N_14972,N_14874);
or UO_800 (O_800,N_14761,N_14719);
nor UO_801 (O_801,N_14820,N_14974);
xnor UO_802 (O_802,N_14919,N_14983);
nor UO_803 (O_803,N_14854,N_14950);
and UO_804 (O_804,N_14748,N_14892);
and UO_805 (O_805,N_14910,N_14824);
or UO_806 (O_806,N_14990,N_14978);
and UO_807 (O_807,N_14976,N_14982);
and UO_808 (O_808,N_14823,N_14928);
nand UO_809 (O_809,N_14797,N_14786);
and UO_810 (O_810,N_14713,N_14919);
nor UO_811 (O_811,N_14911,N_14851);
nor UO_812 (O_812,N_14962,N_14743);
or UO_813 (O_813,N_14803,N_14966);
xnor UO_814 (O_814,N_14765,N_14701);
nor UO_815 (O_815,N_14796,N_14759);
or UO_816 (O_816,N_14712,N_14902);
xor UO_817 (O_817,N_14768,N_14754);
nand UO_818 (O_818,N_14997,N_14756);
xor UO_819 (O_819,N_14930,N_14795);
and UO_820 (O_820,N_14998,N_14799);
and UO_821 (O_821,N_14736,N_14896);
nor UO_822 (O_822,N_14956,N_14937);
and UO_823 (O_823,N_14743,N_14839);
and UO_824 (O_824,N_14828,N_14909);
and UO_825 (O_825,N_14948,N_14918);
xnor UO_826 (O_826,N_14717,N_14970);
and UO_827 (O_827,N_14953,N_14918);
nor UO_828 (O_828,N_14964,N_14700);
and UO_829 (O_829,N_14948,N_14867);
or UO_830 (O_830,N_14913,N_14838);
and UO_831 (O_831,N_14705,N_14743);
or UO_832 (O_832,N_14748,N_14979);
nor UO_833 (O_833,N_14938,N_14734);
xor UO_834 (O_834,N_14973,N_14929);
and UO_835 (O_835,N_14753,N_14727);
and UO_836 (O_836,N_14966,N_14727);
and UO_837 (O_837,N_14966,N_14769);
nor UO_838 (O_838,N_14906,N_14776);
and UO_839 (O_839,N_14894,N_14945);
nand UO_840 (O_840,N_14837,N_14891);
nand UO_841 (O_841,N_14843,N_14975);
nand UO_842 (O_842,N_14995,N_14997);
or UO_843 (O_843,N_14968,N_14921);
xor UO_844 (O_844,N_14730,N_14963);
and UO_845 (O_845,N_14866,N_14889);
or UO_846 (O_846,N_14962,N_14750);
xnor UO_847 (O_847,N_14979,N_14902);
and UO_848 (O_848,N_14924,N_14916);
or UO_849 (O_849,N_14782,N_14760);
or UO_850 (O_850,N_14762,N_14710);
xor UO_851 (O_851,N_14746,N_14818);
xnor UO_852 (O_852,N_14938,N_14936);
or UO_853 (O_853,N_14975,N_14961);
nand UO_854 (O_854,N_14868,N_14707);
and UO_855 (O_855,N_14722,N_14937);
nor UO_856 (O_856,N_14825,N_14814);
xor UO_857 (O_857,N_14816,N_14703);
nor UO_858 (O_858,N_14895,N_14997);
or UO_859 (O_859,N_14876,N_14821);
nor UO_860 (O_860,N_14780,N_14928);
nor UO_861 (O_861,N_14887,N_14935);
nor UO_862 (O_862,N_14957,N_14853);
nand UO_863 (O_863,N_14882,N_14707);
xor UO_864 (O_864,N_14846,N_14785);
xor UO_865 (O_865,N_14757,N_14728);
nor UO_866 (O_866,N_14915,N_14735);
xnor UO_867 (O_867,N_14983,N_14834);
or UO_868 (O_868,N_14913,N_14807);
xnor UO_869 (O_869,N_14771,N_14736);
nand UO_870 (O_870,N_14964,N_14811);
nor UO_871 (O_871,N_14751,N_14993);
and UO_872 (O_872,N_14976,N_14964);
and UO_873 (O_873,N_14818,N_14927);
or UO_874 (O_874,N_14909,N_14822);
or UO_875 (O_875,N_14999,N_14810);
nand UO_876 (O_876,N_14759,N_14708);
and UO_877 (O_877,N_14997,N_14927);
nand UO_878 (O_878,N_14858,N_14741);
and UO_879 (O_879,N_14921,N_14994);
xor UO_880 (O_880,N_14703,N_14911);
nand UO_881 (O_881,N_14892,N_14766);
or UO_882 (O_882,N_14815,N_14850);
and UO_883 (O_883,N_14775,N_14947);
nand UO_884 (O_884,N_14770,N_14934);
nor UO_885 (O_885,N_14903,N_14855);
and UO_886 (O_886,N_14970,N_14816);
and UO_887 (O_887,N_14955,N_14972);
and UO_888 (O_888,N_14939,N_14852);
and UO_889 (O_889,N_14751,N_14916);
nand UO_890 (O_890,N_14982,N_14914);
nor UO_891 (O_891,N_14952,N_14953);
nor UO_892 (O_892,N_14805,N_14827);
or UO_893 (O_893,N_14864,N_14949);
nand UO_894 (O_894,N_14897,N_14826);
nand UO_895 (O_895,N_14820,N_14953);
and UO_896 (O_896,N_14844,N_14968);
nand UO_897 (O_897,N_14822,N_14975);
nor UO_898 (O_898,N_14993,N_14722);
xor UO_899 (O_899,N_14825,N_14727);
nor UO_900 (O_900,N_14708,N_14810);
xnor UO_901 (O_901,N_14849,N_14703);
or UO_902 (O_902,N_14711,N_14852);
and UO_903 (O_903,N_14767,N_14871);
xnor UO_904 (O_904,N_14872,N_14981);
xnor UO_905 (O_905,N_14807,N_14828);
nor UO_906 (O_906,N_14798,N_14866);
nor UO_907 (O_907,N_14718,N_14852);
xnor UO_908 (O_908,N_14743,N_14778);
nor UO_909 (O_909,N_14989,N_14843);
nor UO_910 (O_910,N_14761,N_14814);
and UO_911 (O_911,N_14861,N_14988);
or UO_912 (O_912,N_14766,N_14706);
nand UO_913 (O_913,N_14724,N_14818);
nor UO_914 (O_914,N_14953,N_14758);
xor UO_915 (O_915,N_14800,N_14772);
nand UO_916 (O_916,N_14743,N_14980);
xor UO_917 (O_917,N_14958,N_14779);
or UO_918 (O_918,N_14912,N_14733);
xnor UO_919 (O_919,N_14837,N_14745);
nand UO_920 (O_920,N_14939,N_14740);
or UO_921 (O_921,N_14962,N_14714);
xor UO_922 (O_922,N_14832,N_14885);
nand UO_923 (O_923,N_14997,N_14812);
nand UO_924 (O_924,N_14727,N_14768);
or UO_925 (O_925,N_14875,N_14805);
xnor UO_926 (O_926,N_14974,N_14787);
nand UO_927 (O_927,N_14788,N_14876);
xnor UO_928 (O_928,N_14934,N_14802);
xnor UO_929 (O_929,N_14970,N_14860);
or UO_930 (O_930,N_14909,N_14840);
nand UO_931 (O_931,N_14984,N_14858);
or UO_932 (O_932,N_14876,N_14822);
or UO_933 (O_933,N_14705,N_14753);
xnor UO_934 (O_934,N_14805,N_14761);
xnor UO_935 (O_935,N_14713,N_14731);
xnor UO_936 (O_936,N_14810,N_14954);
and UO_937 (O_937,N_14956,N_14921);
xor UO_938 (O_938,N_14951,N_14819);
nor UO_939 (O_939,N_14913,N_14945);
or UO_940 (O_940,N_14812,N_14868);
or UO_941 (O_941,N_14762,N_14750);
nor UO_942 (O_942,N_14937,N_14725);
xnor UO_943 (O_943,N_14885,N_14736);
and UO_944 (O_944,N_14729,N_14783);
nand UO_945 (O_945,N_14807,N_14716);
or UO_946 (O_946,N_14736,N_14802);
nor UO_947 (O_947,N_14825,N_14846);
nor UO_948 (O_948,N_14741,N_14829);
and UO_949 (O_949,N_14923,N_14807);
and UO_950 (O_950,N_14911,N_14946);
nand UO_951 (O_951,N_14768,N_14971);
xnor UO_952 (O_952,N_14826,N_14941);
xor UO_953 (O_953,N_14943,N_14935);
or UO_954 (O_954,N_14738,N_14834);
and UO_955 (O_955,N_14893,N_14855);
or UO_956 (O_956,N_14797,N_14855);
and UO_957 (O_957,N_14884,N_14753);
nor UO_958 (O_958,N_14803,N_14896);
xor UO_959 (O_959,N_14707,N_14785);
and UO_960 (O_960,N_14813,N_14959);
xnor UO_961 (O_961,N_14716,N_14908);
nand UO_962 (O_962,N_14885,N_14884);
xor UO_963 (O_963,N_14779,N_14957);
nand UO_964 (O_964,N_14912,N_14950);
nor UO_965 (O_965,N_14764,N_14853);
nand UO_966 (O_966,N_14854,N_14732);
xnor UO_967 (O_967,N_14996,N_14743);
nand UO_968 (O_968,N_14922,N_14934);
nand UO_969 (O_969,N_14731,N_14809);
nor UO_970 (O_970,N_14969,N_14737);
nand UO_971 (O_971,N_14755,N_14874);
and UO_972 (O_972,N_14758,N_14962);
nor UO_973 (O_973,N_14701,N_14992);
and UO_974 (O_974,N_14902,N_14736);
and UO_975 (O_975,N_14885,N_14709);
and UO_976 (O_976,N_14883,N_14999);
and UO_977 (O_977,N_14816,N_14716);
nand UO_978 (O_978,N_14778,N_14764);
nor UO_979 (O_979,N_14909,N_14813);
or UO_980 (O_980,N_14991,N_14904);
nor UO_981 (O_981,N_14959,N_14936);
and UO_982 (O_982,N_14750,N_14770);
or UO_983 (O_983,N_14779,N_14848);
nor UO_984 (O_984,N_14946,N_14700);
xnor UO_985 (O_985,N_14993,N_14854);
and UO_986 (O_986,N_14731,N_14905);
or UO_987 (O_987,N_14997,N_14744);
nand UO_988 (O_988,N_14877,N_14828);
xor UO_989 (O_989,N_14704,N_14713);
xor UO_990 (O_990,N_14917,N_14907);
xnor UO_991 (O_991,N_14736,N_14746);
nor UO_992 (O_992,N_14896,N_14904);
nand UO_993 (O_993,N_14806,N_14803);
nor UO_994 (O_994,N_14816,N_14883);
or UO_995 (O_995,N_14895,N_14814);
nand UO_996 (O_996,N_14911,N_14857);
or UO_997 (O_997,N_14780,N_14877);
nor UO_998 (O_998,N_14719,N_14794);
or UO_999 (O_999,N_14850,N_14883);
xor UO_1000 (O_1000,N_14738,N_14769);
nor UO_1001 (O_1001,N_14798,N_14918);
and UO_1002 (O_1002,N_14734,N_14779);
nor UO_1003 (O_1003,N_14849,N_14981);
nand UO_1004 (O_1004,N_14710,N_14917);
or UO_1005 (O_1005,N_14700,N_14820);
nand UO_1006 (O_1006,N_14814,N_14758);
or UO_1007 (O_1007,N_14716,N_14758);
nor UO_1008 (O_1008,N_14956,N_14704);
nand UO_1009 (O_1009,N_14932,N_14839);
nor UO_1010 (O_1010,N_14833,N_14964);
nand UO_1011 (O_1011,N_14961,N_14978);
nand UO_1012 (O_1012,N_14754,N_14737);
xor UO_1013 (O_1013,N_14780,N_14718);
or UO_1014 (O_1014,N_14870,N_14852);
nand UO_1015 (O_1015,N_14836,N_14905);
and UO_1016 (O_1016,N_14849,N_14712);
and UO_1017 (O_1017,N_14820,N_14980);
or UO_1018 (O_1018,N_14974,N_14775);
and UO_1019 (O_1019,N_14791,N_14939);
xor UO_1020 (O_1020,N_14779,N_14926);
nand UO_1021 (O_1021,N_14760,N_14951);
or UO_1022 (O_1022,N_14927,N_14970);
xnor UO_1023 (O_1023,N_14937,N_14847);
nand UO_1024 (O_1024,N_14774,N_14823);
xnor UO_1025 (O_1025,N_14884,N_14880);
nor UO_1026 (O_1026,N_14730,N_14876);
xor UO_1027 (O_1027,N_14957,N_14758);
or UO_1028 (O_1028,N_14843,N_14951);
or UO_1029 (O_1029,N_14738,N_14942);
or UO_1030 (O_1030,N_14804,N_14901);
nand UO_1031 (O_1031,N_14919,N_14770);
nor UO_1032 (O_1032,N_14959,N_14984);
xnor UO_1033 (O_1033,N_14960,N_14994);
xnor UO_1034 (O_1034,N_14953,N_14956);
xnor UO_1035 (O_1035,N_14832,N_14810);
nand UO_1036 (O_1036,N_14889,N_14906);
nand UO_1037 (O_1037,N_14803,N_14730);
and UO_1038 (O_1038,N_14971,N_14931);
or UO_1039 (O_1039,N_14816,N_14874);
nor UO_1040 (O_1040,N_14897,N_14739);
or UO_1041 (O_1041,N_14904,N_14885);
nor UO_1042 (O_1042,N_14821,N_14732);
nor UO_1043 (O_1043,N_14891,N_14893);
xor UO_1044 (O_1044,N_14835,N_14873);
nand UO_1045 (O_1045,N_14787,N_14962);
and UO_1046 (O_1046,N_14898,N_14725);
and UO_1047 (O_1047,N_14910,N_14975);
nor UO_1048 (O_1048,N_14828,N_14771);
xor UO_1049 (O_1049,N_14875,N_14796);
nand UO_1050 (O_1050,N_14871,N_14963);
and UO_1051 (O_1051,N_14758,N_14857);
and UO_1052 (O_1052,N_14966,N_14980);
nor UO_1053 (O_1053,N_14853,N_14990);
nor UO_1054 (O_1054,N_14898,N_14893);
xor UO_1055 (O_1055,N_14735,N_14935);
nor UO_1056 (O_1056,N_14889,N_14785);
nand UO_1057 (O_1057,N_14793,N_14983);
xor UO_1058 (O_1058,N_14996,N_14971);
xor UO_1059 (O_1059,N_14901,N_14798);
xor UO_1060 (O_1060,N_14717,N_14896);
xor UO_1061 (O_1061,N_14843,N_14892);
or UO_1062 (O_1062,N_14837,N_14842);
nor UO_1063 (O_1063,N_14991,N_14880);
nand UO_1064 (O_1064,N_14896,N_14856);
nor UO_1065 (O_1065,N_14742,N_14996);
and UO_1066 (O_1066,N_14942,N_14728);
xor UO_1067 (O_1067,N_14855,N_14700);
or UO_1068 (O_1068,N_14791,N_14903);
or UO_1069 (O_1069,N_14963,N_14781);
nor UO_1070 (O_1070,N_14736,N_14990);
xnor UO_1071 (O_1071,N_14943,N_14941);
and UO_1072 (O_1072,N_14897,N_14719);
and UO_1073 (O_1073,N_14990,N_14744);
and UO_1074 (O_1074,N_14714,N_14708);
and UO_1075 (O_1075,N_14865,N_14911);
xor UO_1076 (O_1076,N_14886,N_14814);
or UO_1077 (O_1077,N_14929,N_14963);
nand UO_1078 (O_1078,N_14782,N_14989);
nand UO_1079 (O_1079,N_14804,N_14807);
xor UO_1080 (O_1080,N_14874,N_14890);
or UO_1081 (O_1081,N_14911,N_14881);
nor UO_1082 (O_1082,N_14732,N_14791);
nor UO_1083 (O_1083,N_14747,N_14814);
or UO_1084 (O_1084,N_14981,N_14960);
nand UO_1085 (O_1085,N_14990,N_14810);
xnor UO_1086 (O_1086,N_14718,N_14969);
nand UO_1087 (O_1087,N_14771,N_14918);
or UO_1088 (O_1088,N_14790,N_14902);
nand UO_1089 (O_1089,N_14805,N_14974);
nand UO_1090 (O_1090,N_14787,N_14785);
nand UO_1091 (O_1091,N_14735,N_14761);
xnor UO_1092 (O_1092,N_14809,N_14995);
nand UO_1093 (O_1093,N_14889,N_14710);
or UO_1094 (O_1094,N_14885,N_14815);
nand UO_1095 (O_1095,N_14819,N_14850);
or UO_1096 (O_1096,N_14845,N_14844);
nand UO_1097 (O_1097,N_14862,N_14952);
and UO_1098 (O_1098,N_14893,N_14923);
and UO_1099 (O_1099,N_14988,N_14967);
nor UO_1100 (O_1100,N_14790,N_14823);
or UO_1101 (O_1101,N_14864,N_14797);
nor UO_1102 (O_1102,N_14931,N_14732);
nand UO_1103 (O_1103,N_14726,N_14700);
nor UO_1104 (O_1104,N_14872,N_14737);
xnor UO_1105 (O_1105,N_14937,N_14968);
and UO_1106 (O_1106,N_14781,N_14869);
and UO_1107 (O_1107,N_14805,N_14874);
or UO_1108 (O_1108,N_14969,N_14745);
nor UO_1109 (O_1109,N_14904,N_14866);
nand UO_1110 (O_1110,N_14830,N_14923);
xnor UO_1111 (O_1111,N_14892,N_14932);
or UO_1112 (O_1112,N_14902,N_14887);
xor UO_1113 (O_1113,N_14759,N_14741);
and UO_1114 (O_1114,N_14882,N_14765);
nand UO_1115 (O_1115,N_14883,N_14734);
xnor UO_1116 (O_1116,N_14878,N_14852);
xnor UO_1117 (O_1117,N_14844,N_14964);
or UO_1118 (O_1118,N_14898,N_14978);
and UO_1119 (O_1119,N_14947,N_14731);
nand UO_1120 (O_1120,N_14952,N_14789);
or UO_1121 (O_1121,N_14987,N_14903);
nor UO_1122 (O_1122,N_14897,N_14718);
nor UO_1123 (O_1123,N_14833,N_14913);
nor UO_1124 (O_1124,N_14715,N_14814);
nand UO_1125 (O_1125,N_14870,N_14949);
or UO_1126 (O_1126,N_14731,N_14767);
xor UO_1127 (O_1127,N_14947,N_14914);
or UO_1128 (O_1128,N_14905,N_14736);
or UO_1129 (O_1129,N_14981,N_14873);
nor UO_1130 (O_1130,N_14904,N_14782);
nand UO_1131 (O_1131,N_14866,N_14933);
xor UO_1132 (O_1132,N_14872,N_14994);
xor UO_1133 (O_1133,N_14970,N_14993);
nand UO_1134 (O_1134,N_14806,N_14737);
or UO_1135 (O_1135,N_14993,N_14712);
xor UO_1136 (O_1136,N_14721,N_14923);
xnor UO_1137 (O_1137,N_14937,N_14767);
or UO_1138 (O_1138,N_14874,N_14839);
or UO_1139 (O_1139,N_14843,N_14702);
xnor UO_1140 (O_1140,N_14846,N_14868);
and UO_1141 (O_1141,N_14895,N_14964);
nand UO_1142 (O_1142,N_14723,N_14904);
and UO_1143 (O_1143,N_14991,N_14867);
nand UO_1144 (O_1144,N_14812,N_14979);
nand UO_1145 (O_1145,N_14736,N_14806);
xnor UO_1146 (O_1146,N_14823,N_14732);
or UO_1147 (O_1147,N_14734,N_14989);
xnor UO_1148 (O_1148,N_14767,N_14881);
xnor UO_1149 (O_1149,N_14795,N_14751);
nor UO_1150 (O_1150,N_14775,N_14967);
or UO_1151 (O_1151,N_14835,N_14716);
or UO_1152 (O_1152,N_14809,N_14900);
and UO_1153 (O_1153,N_14831,N_14817);
or UO_1154 (O_1154,N_14865,N_14774);
and UO_1155 (O_1155,N_14779,N_14746);
nor UO_1156 (O_1156,N_14796,N_14726);
xor UO_1157 (O_1157,N_14747,N_14812);
and UO_1158 (O_1158,N_14813,N_14951);
xor UO_1159 (O_1159,N_14870,N_14830);
and UO_1160 (O_1160,N_14775,N_14907);
nor UO_1161 (O_1161,N_14966,N_14929);
nand UO_1162 (O_1162,N_14981,N_14738);
and UO_1163 (O_1163,N_14858,N_14755);
and UO_1164 (O_1164,N_14950,N_14745);
xor UO_1165 (O_1165,N_14954,N_14952);
or UO_1166 (O_1166,N_14829,N_14828);
nand UO_1167 (O_1167,N_14799,N_14912);
xnor UO_1168 (O_1168,N_14763,N_14862);
nand UO_1169 (O_1169,N_14737,N_14880);
or UO_1170 (O_1170,N_14901,N_14976);
xor UO_1171 (O_1171,N_14860,N_14717);
nand UO_1172 (O_1172,N_14773,N_14799);
xnor UO_1173 (O_1173,N_14732,N_14871);
or UO_1174 (O_1174,N_14724,N_14710);
or UO_1175 (O_1175,N_14908,N_14935);
nand UO_1176 (O_1176,N_14886,N_14734);
nand UO_1177 (O_1177,N_14749,N_14900);
nor UO_1178 (O_1178,N_14914,N_14975);
and UO_1179 (O_1179,N_14985,N_14925);
or UO_1180 (O_1180,N_14981,N_14728);
and UO_1181 (O_1181,N_14747,N_14743);
nand UO_1182 (O_1182,N_14916,N_14943);
or UO_1183 (O_1183,N_14847,N_14855);
nor UO_1184 (O_1184,N_14807,N_14728);
nor UO_1185 (O_1185,N_14887,N_14812);
xnor UO_1186 (O_1186,N_14873,N_14945);
and UO_1187 (O_1187,N_14892,N_14906);
and UO_1188 (O_1188,N_14900,N_14804);
xor UO_1189 (O_1189,N_14726,N_14767);
or UO_1190 (O_1190,N_14969,N_14889);
xor UO_1191 (O_1191,N_14861,N_14994);
nand UO_1192 (O_1192,N_14797,N_14723);
xnor UO_1193 (O_1193,N_14862,N_14700);
xor UO_1194 (O_1194,N_14888,N_14838);
nor UO_1195 (O_1195,N_14950,N_14975);
or UO_1196 (O_1196,N_14793,N_14906);
or UO_1197 (O_1197,N_14902,N_14982);
nor UO_1198 (O_1198,N_14883,N_14729);
or UO_1199 (O_1199,N_14937,N_14726);
nor UO_1200 (O_1200,N_14836,N_14815);
xor UO_1201 (O_1201,N_14755,N_14816);
nand UO_1202 (O_1202,N_14827,N_14866);
nand UO_1203 (O_1203,N_14959,N_14734);
nor UO_1204 (O_1204,N_14727,N_14874);
and UO_1205 (O_1205,N_14766,N_14923);
nor UO_1206 (O_1206,N_14731,N_14920);
and UO_1207 (O_1207,N_14736,N_14963);
xor UO_1208 (O_1208,N_14960,N_14949);
or UO_1209 (O_1209,N_14881,N_14765);
or UO_1210 (O_1210,N_14754,N_14712);
and UO_1211 (O_1211,N_14851,N_14823);
and UO_1212 (O_1212,N_14715,N_14917);
xnor UO_1213 (O_1213,N_14803,N_14856);
nand UO_1214 (O_1214,N_14971,N_14858);
or UO_1215 (O_1215,N_14871,N_14925);
and UO_1216 (O_1216,N_14933,N_14911);
nor UO_1217 (O_1217,N_14895,N_14983);
nand UO_1218 (O_1218,N_14866,N_14999);
nand UO_1219 (O_1219,N_14799,N_14980);
xor UO_1220 (O_1220,N_14764,N_14889);
or UO_1221 (O_1221,N_14848,N_14893);
or UO_1222 (O_1222,N_14914,N_14834);
and UO_1223 (O_1223,N_14823,N_14831);
and UO_1224 (O_1224,N_14938,N_14924);
nor UO_1225 (O_1225,N_14933,N_14992);
or UO_1226 (O_1226,N_14943,N_14869);
and UO_1227 (O_1227,N_14783,N_14866);
or UO_1228 (O_1228,N_14884,N_14800);
nand UO_1229 (O_1229,N_14887,N_14931);
or UO_1230 (O_1230,N_14865,N_14717);
or UO_1231 (O_1231,N_14960,N_14700);
nand UO_1232 (O_1232,N_14946,N_14822);
and UO_1233 (O_1233,N_14799,N_14861);
or UO_1234 (O_1234,N_14781,N_14803);
nand UO_1235 (O_1235,N_14806,N_14894);
or UO_1236 (O_1236,N_14971,N_14895);
nor UO_1237 (O_1237,N_14726,N_14900);
nor UO_1238 (O_1238,N_14936,N_14990);
and UO_1239 (O_1239,N_14726,N_14908);
xor UO_1240 (O_1240,N_14920,N_14852);
nand UO_1241 (O_1241,N_14743,N_14978);
nor UO_1242 (O_1242,N_14959,N_14737);
nor UO_1243 (O_1243,N_14841,N_14902);
or UO_1244 (O_1244,N_14832,N_14894);
nand UO_1245 (O_1245,N_14790,N_14712);
and UO_1246 (O_1246,N_14987,N_14703);
or UO_1247 (O_1247,N_14784,N_14900);
xor UO_1248 (O_1248,N_14970,N_14742);
nand UO_1249 (O_1249,N_14993,N_14834);
nand UO_1250 (O_1250,N_14808,N_14810);
xor UO_1251 (O_1251,N_14979,N_14760);
nand UO_1252 (O_1252,N_14771,N_14718);
nand UO_1253 (O_1253,N_14953,N_14717);
xnor UO_1254 (O_1254,N_14901,N_14909);
nand UO_1255 (O_1255,N_14734,N_14965);
or UO_1256 (O_1256,N_14713,N_14856);
nor UO_1257 (O_1257,N_14912,N_14715);
nand UO_1258 (O_1258,N_14823,N_14947);
xor UO_1259 (O_1259,N_14971,N_14887);
nor UO_1260 (O_1260,N_14965,N_14867);
nand UO_1261 (O_1261,N_14824,N_14736);
nand UO_1262 (O_1262,N_14924,N_14866);
nand UO_1263 (O_1263,N_14968,N_14797);
nand UO_1264 (O_1264,N_14747,N_14926);
nand UO_1265 (O_1265,N_14717,N_14763);
xnor UO_1266 (O_1266,N_14857,N_14831);
or UO_1267 (O_1267,N_14915,N_14869);
nand UO_1268 (O_1268,N_14827,N_14784);
or UO_1269 (O_1269,N_14973,N_14700);
nand UO_1270 (O_1270,N_14744,N_14821);
and UO_1271 (O_1271,N_14716,N_14820);
nor UO_1272 (O_1272,N_14855,N_14995);
and UO_1273 (O_1273,N_14756,N_14824);
nor UO_1274 (O_1274,N_14856,N_14815);
xor UO_1275 (O_1275,N_14838,N_14951);
and UO_1276 (O_1276,N_14926,N_14749);
or UO_1277 (O_1277,N_14718,N_14705);
nor UO_1278 (O_1278,N_14762,N_14771);
xor UO_1279 (O_1279,N_14712,N_14991);
or UO_1280 (O_1280,N_14956,N_14751);
nand UO_1281 (O_1281,N_14907,N_14732);
nand UO_1282 (O_1282,N_14805,N_14708);
nor UO_1283 (O_1283,N_14805,N_14760);
nand UO_1284 (O_1284,N_14724,N_14911);
and UO_1285 (O_1285,N_14965,N_14969);
or UO_1286 (O_1286,N_14844,N_14838);
nand UO_1287 (O_1287,N_14896,N_14923);
xor UO_1288 (O_1288,N_14934,N_14950);
xnor UO_1289 (O_1289,N_14931,N_14968);
nand UO_1290 (O_1290,N_14704,N_14701);
or UO_1291 (O_1291,N_14748,N_14901);
xnor UO_1292 (O_1292,N_14918,N_14709);
nor UO_1293 (O_1293,N_14836,N_14944);
and UO_1294 (O_1294,N_14935,N_14742);
or UO_1295 (O_1295,N_14737,N_14832);
or UO_1296 (O_1296,N_14964,N_14807);
and UO_1297 (O_1297,N_14763,N_14922);
nand UO_1298 (O_1298,N_14915,N_14810);
nand UO_1299 (O_1299,N_14955,N_14778);
nor UO_1300 (O_1300,N_14984,N_14722);
and UO_1301 (O_1301,N_14885,N_14897);
or UO_1302 (O_1302,N_14748,N_14957);
nor UO_1303 (O_1303,N_14856,N_14987);
nand UO_1304 (O_1304,N_14752,N_14811);
nand UO_1305 (O_1305,N_14937,N_14739);
nand UO_1306 (O_1306,N_14829,N_14845);
nand UO_1307 (O_1307,N_14922,N_14751);
nand UO_1308 (O_1308,N_14975,N_14953);
nor UO_1309 (O_1309,N_14885,N_14789);
and UO_1310 (O_1310,N_14742,N_14737);
and UO_1311 (O_1311,N_14996,N_14876);
nor UO_1312 (O_1312,N_14856,N_14967);
nor UO_1313 (O_1313,N_14741,N_14765);
nor UO_1314 (O_1314,N_14976,N_14926);
xnor UO_1315 (O_1315,N_14918,N_14831);
or UO_1316 (O_1316,N_14706,N_14902);
nor UO_1317 (O_1317,N_14886,N_14764);
and UO_1318 (O_1318,N_14923,N_14795);
xor UO_1319 (O_1319,N_14893,N_14824);
or UO_1320 (O_1320,N_14964,N_14883);
and UO_1321 (O_1321,N_14964,N_14825);
and UO_1322 (O_1322,N_14876,N_14809);
xnor UO_1323 (O_1323,N_14779,N_14869);
xnor UO_1324 (O_1324,N_14882,N_14897);
nor UO_1325 (O_1325,N_14894,N_14879);
nor UO_1326 (O_1326,N_14890,N_14993);
nor UO_1327 (O_1327,N_14744,N_14740);
or UO_1328 (O_1328,N_14712,N_14814);
and UO_1329 (O_1329,N_14873,N_14890);
nand UO_1330 (O_1330,N_14835,N_14932);
nor UO_1331 (O_1331,N_14764,N_14845);
nand UO_1332 (O_1332,N_14854,N_14821);
xnor UO_1333 (O_1333,N_14961,N_14738);
nor UO_1334 (O_1334,N_14829,N_14911);
or UO_1335 (O_1335,N_14841,N_14992);
nand UO_1336 (O_1336,N_14816,N_14877);
or UO_1337 (O_1337,N_14736,N_14900);
xnor UO_1338 (O_1338,N_14994,N_14922);
and UO_1339 (O_1339,N_14933,N_14781);
and UO_1340 (O_1340,N_14999,N_14930);
nor UO_1341 (O_1341,N_14934,N_14961);
nand UO_1342 (O_1342,N_14836,N_14760);
and UO_1343 (O_1343,N_14764,N_14835);
or UO_1344 (O_1344,N_14800,N_14945);
nand UO_1345 (O_1345,N_14984,N_14721);
or UO_1346 (O_1346,N_14846,N_14709);
xor UO_1347 (O_1347,N_14770,N_14998);
and UO_1348 (O_1348,N_14976,N_14826);
nand UO_1349 (O_1349,N_14933,N_14959);
nand UO_1350 (O_1350,N_14780,N_14772);
and UO_1351 (O_1351,N_14914,N_14971);
and UO_1352 (O_1352,N_14854,N_14976);
and UO_1353 (O_1353,N_14717,N_14831);
nand UO_1354 (O_1354,N_14941,N_14957);
or UO_1355 (O_1355,N_14815,N_14707);
xor UO_1356 (O_1356,N_14870,N_14828);
and UO_1357 (O_1357,N_14965,N_14752);
nor UO_1358 (O_1358,N_14701,N_14872);
and UO_1359 (O_1359,N_14915,N_14734);
or UO_1360 (O_1360,N_14893,N_14867);
or UO_1361 (O_1361,N_14902,N_14801);
nand UO_1362 (O_1362,N_14758,N_14908);
nand UO_1363 (O_1363,N_14778,N_14730);
xnor UO_1364 (O_1364,N_14721,N_14762);
nand UO_1365 (O_1365,N_14985,N_14962);
nor UO_1366 (O_1366,N_14999,N_14704);
nand UO_1367 (O_1367,N_14803,N_14886);
or UO_1368 (O_1368,N_14913,N_14995);
and UO_1369 (O_1369,N_14892,N_14761);
and UO_1370 (O_1370,N_14895,N_14704);
nor UO_1371 (O_1371,N_14961,N_14779);
nor UO_1372 (O_1372,N_14940,N_14892);
or UO_1373 (O_1373,N_14811,N_14878);
or UO_1374 (O_1374,N_14741,N_14793);
or UO_1375 (O_1375,N_14811,N_14750);
nand UO_1376 (O_1376,N_14785,N_14802);
nand UO_1377 (O_1377,N_14874,N_14885);
xor UO_1378 (O_1378,N_14980,N_14709);
nor UO_1379 (O_1379,N_14917,N_14723);
and UO_1380 (O_1380,N_14840,N_14890);
nor UO_1381 (O_1381,N_14920,N_14953);
nor UO_1382 (O_1382,N_14934,N_14869);
and UO_1383 (O_1383,N_14821,N_14912);
nor UO_1384 (O_1384,N_14940,N_14815);
nand UO_1385 (O_1385,N_14822,N_14779);
xor UO_1386 (O_1386,N_14935,N_14892);
xor UO_1387 (O_1387,N_14990,N_14882);
and UO_1388 (O_1388,N_14903,N_14833);
xor UO_1389 (O_1389,N_14702,N_14856);
xnor UO_1390 (O_1390,N_14883,N_14996);
and UO_1391 (O_1391,N_14936,N_14881);
nand UO_1392 (O_1392,N_14964,N_14719);
nor UO_1393 (O_1393,N_14994,N_14746);
or UO_1394 (O_1394,N_14954,N_14790);
and UO_1395 (O_1395,N_14724,N_14840);
and UO_1396 (O_1396,N_14722,N_14711);
nand UO_1397 (O_1397,N_14911,N_14896);
nand UO_1398 (O_1398,N_14961,N_14927);
xnor UO_1399 (O_1399,N_14874,N_14759);
nand UO_1400 (O_1400,N_14706,N_14717);
nor UO_1401 (O_1401,N_14817,N_14728);
xor UO_1402 (O_1402,N_14881,N_14906);
or UO_1403 (O_1403,N_14819,N_14726);
xor UO_1404 (O_1404,N_14853,N_14904);
or UO_1405 (O_1405,N_14763,N_14864);
and UO_1406 (O_1406,N_14821,N_14718);
nand UO_1407 (O_1407,N_14743,N_14913);
nor UO_1408 (O_1408,N_14912,N_14745);
nor UO_1409 (O_1409,N_14792,N_14969);
nand UO_1410 (O_1410,N_14890,N_14711);
and UO_1411 (O_1411,N_14818,N_14866);
nor UO_1412 (O_1412,N_14793,N_14999);
or UO_1413 (O_1413,N_14792,N_14723);
xnor UO_1414 (O_1414,N_14848,N_14908);
xnor UO_1415 (O_1415,N_14745,N_14983);
nand UO_1416 (O_1416,N_14777,N_14749);
nor UO_1417 (O_1417,N_14725,N_14890);
nor UO_1418 (O_1418,N_14932,N_14840);
xor UO_1419 (O_1419,N_14896,N_14745);
nand UO_1420 (O_1420,N_14872,N_14885);
nor UO_1421 (O_1421,N_14946,N_14804);
nand UO_1422 (O_1422,N_14765,N_14873);
or UO_1423 (O_1423,N_14778,N_14785);
xor UO_1424 (O_1424,N_14959,N_14714);
nand UO_1425 (O_1425,N_14905,N_14920);
xnor UO_1426 (O_1426,N_14956,N_14849);
nand UO_1427 (O_1427,N_14883,N_14716);
and UO_1428 (O_1428,N_14806,N_14997);
xnor UO_1429 (O_1429,N_14764,N_14794);
or UO_1430 (O_1430,N_14920,N_14824);
nand UO_1431 (O_1431,N_14766,N_14759);
xor UO_1432 (O_1432,N_14749,N_14853);
and UO_1433 (O_1433,N_14952,N_14740);
or UO_1434 (O_1434,N_14781,N_14932);
and UO_1435 (O_1435,N_14779,N_14854);
or UO_1436 (O_1436,N_14954,N_14753);
and UO_1437 (O_1437,N_14861,N_14852);
nand UO_1438 (O_1438,N_14990,N_14706);
and UO_1439 (O_1439,N_14854,N_14951);
nor UO_1440 (O_1440,N_14882,N_14847);
and UO_1441 (O_1441,N_14933,N_14736);
xor UO_1442 (O_1442,N_14901,N_14995);
xnor UO_1443 (O_1443,N_14752,N_14968);
and UO_1444 (O_1444,N_14787,N_14739);
nand UO_1445 (O_1445,N_14925,N_14755);
nor UO_1446 (O_1446,N_14745,N_14945);
xor UO_1447 (O_1447,N_14860,N_14961);
and UO_1448 (O_1448,N_14890,N_14742);
nand UO_1449 (O_1449,N_14838,N_14764);
or UO_1450 (O_1450,N_14924,N_14827);
and UO_1451 (O_1451,N_14836,N_14731);
xnor UO_1452 (O_1452,N_14707,N_14720);
or UO_1453 (O_1453,N_14755,N_14722);
and UO_1454 (O_1454,N_14915,N_14748);
or UO_1455 (O_1455,N_14898,N_14987);
and UO_1456 (O_1456,N_14871,N_14786);
nor UO_1457 (O_1457,N_14903,N_14974);
xnor UO_1458 (O_1458,N_14942,N_14746);
nand UO_1459 (O_1459,N_14750,N_14900);
xor UO_1460 (O_1460,N_14906,N_14962);
nor UO_1461 (O_1461,N_14999,N_14726);
nand UO_1462 (O_1462,N_14912,N_14856);
and UO_1463 (O_1463,N_14862,N_14971);
nand UO_1464 (O_1464,N_14931,N_14860);
nand UO_1465 (O_1465,N_14701,N_14755);
nor UO_1466 (O_1466,N_14959,N_14926);
nand UO_1467 (O_1467,N_14734,N_14980);
xor UO_1468 (O_1468,N_14745,N_14768);
and UO_1469 (O_1469,N_14834,N_14955);
and UO_1470 (O_1470,N_14928,N_14718);
xor UO_1471 (O_1471,N_14947,N_14734);
and UO_1472 (O_1472,N_14789,N_14843);
nor UO_1473 (O_1473,N_14885,N_14739);
or UO_1474 (O_1474,N_14930,N_14855);
and UO_1475 (O_1475,N_14779,N_14847);
xnor UO_1476 (O_1476,N_14920,N_14806);
nor UO_1477 (O_1477,N_14971,N_14756);
nor UO_1478 (O_1478,N_14710,N_14941);
and UO_1479 (O_1479,N_14985,N_14822);
xnor UO_1480 (O_1480,N_14877,N_14897);
nor UO_1481 (O_1481,N_14812,N_14950);
nor UO_1482 (O_1482,N_14998,N_14979);
nor UO_1483 (O_1483,N_14918,N_14908);
xor UO_1484 (O_1484,N_14803,N_14881);
and UO_1485 (O_1485,N_14786,N_14830);
and UO_1486 (O_1486,N_14719,N_14818);
nand UO_1487 (O_1487,N_14795,N_14732);
or UO_1488 (O_1488,N_14721,N_14705);
xor UO_1489 (O_1489,N_14744,N_14836);
nand UO_1490 (O_1490,N_14849,N_14977);
nand UO_1491 (O_1491,N_14729,N_14952);
and UO_1492 (O_1492,N_14794,N_14782);
or UO_1493 (O_1493,N_14979,N_14780);
xor UO_1494 (O_1494,N_14815,N_14711);
or UO_1495 (O_1495,N_14966,N_14722);
nor UO_1496 (O_1496,N_14801,N_14843);
nor UO_1497 (O_1497,N_14906,N_14941);
xnor UO_1498 (O_1498,N_14719,N_14725);
or UO_1499 (O_1499,N_14994,N_14774);
nand UO_1500 (O_1500,N_14809,N_14931);
xor UO_1501 (O_1501,N_14770,N_14884);
nand UO_1502 (O_1502,N_14936,N_14798);
xnor UO_1503 (O_1503,N_14757,N_14919);
xor UO_1504 (O_1504,N_14788,N_14759);
and UO_1505 (O_1505,N_14901,N_14762);
nand UO_1506 (O_1506,N_14937,N_14729);
xor UO_1507 (O_1507,N_14763,N_14882);
nand UO_1508 (O_1508,N_14824,N_14812);
and UO_1509 (O_1509,N_14895,N_14871);
xor UO_1510 (O_1510,N_14912,N_14731);
nand UO_1511 (O_1511,N_14971,N_14873);
or UO_1512 (O_1512,N_14776,N_14736);
nand UO_1513 (O_1513,N_14748,N_14886);
nor UO_1514 (O_1514,N_14932,N_14770);
and UO_1515 (O_1515,N_14719,N_14955);
nand UO_1516 (O_1516,N_14972,N_14746);
and UO_1517 (O_1517,N_14931,N_14806);
or UO_1518 (O_1518,N_14929,N_14809);
nand UO_1519 (O_1519,N_14908,N_14724);
nor UO_1520 (O_1520,N_14948,N_14873);
and UO_1521 (O_1521,N_14820,N_14717);
and UO_1522 (O_1522,N_14895,N_14712);
xnor UO_1523 (O_1523,N_14908,N_14957);
nand UO_1524 (O_1524,N_14906,N_14710);
nand UO_1525 (O_1525,N_14765,N_14989);
or UO_1526 (O_1526,N_14783,N_14812);
xnor UO_1527 (O_1527,N_14931,N_14925);
nand UO_1528 (O_1528,N_14957,N_14942);
or UO_1529 (O_1529,N_14919,N_14900);
nor UO_1530 (O_1530,N_14791,N_14793);
or UO_1531 (O_1531,N_14904,N_14736);
nand UO_1532 (O_1532,N_14796,N_14919);
nand UO_1533 (O_1533,N_14912,N_14729);
nand UO_1534 (O_1534,N_14924,N_14828);
nand UO_1535 (O_1535,N_14824,N_14793);
xor UO_1536 (O_1536,N_14889,N_14749);
or UO_1537 (O_1537,N_14737,N_14948);
nor UO_1538 (O_1538,N_14835,N_14885);
nand UO_1539 (O_1539,N_14851,N_14924);
xor UO_1540 (O_1540,N_14996,N_14882);
nand UO_1541 (O_1541,N_14727,N_14950);
and UO_1542 (O_1542,N_14953,N_14723);
and UO_1543 (O_1543,N_14855,N_14904);
xnor UO_1544 (O_1544,N_14828,N_14722);
and UO_1545 (O_1545,N_14855,N_14980);
xnor UO_1546 (O_1546,N_14833,N_14816);
nor UO_1547 (O_1547,N_14930,N_14945);
nand UO_1548 (O_1548,N_14954,N_14870);
nor UO_1549 (O_1549,N_14747,N_14983);
nand UO_1550 (O_1550,N_14982,N_14916);
xnor UO_1551 (O_1551,N_14747,N_14703);
nor UO_1552 (O_1552,N_14817,N_14870);
nand UO_1553 (O_1553,N_14965,N_14897);
or UO_1554 (O_1554,N_14713,N_14886);
nand UO_1555 (O_1555,N_14835,N_14907);
xor UO_1556 (O_1556,N_14861,N_14897);
nor UO_1557 (O_1557,N_14965,N_14784);
xor UO_1558 (O_1558,N_14845,N_14874);
or UO_1559 (O_1559,N_14952,N_14734);
nand UO_1560 (O_1560,N_14764,N_14904);
nor UO_1561 (O_1561,N_14862,N_14961);
nand UO_1562 (O_1562,N_14773,N_14769);
and UO_1563 (O_1563,N_14842,N_14857);
nor UO_1564 (O_1564,N_14798,N_14760);
or UO_1565 (O_1565,N_14743,N_14734);
nand UO_1566 (O_1566,N_14727,N_14832);
nand UO_1567 (O_1567,N_14983,N_14902);
nor UO_1568 (O_1568,N_14773,N_14928);
and UO_1569 (O_1569,N_14988,N_14978);
or UO_1570 (O_1570,N_14958,N_14858);
xnor UO_1571 (O_1571,N_14907,N_14719);
or UO_1572 (O_1572,N_14997,N_14720);
nor UO_1573 (O_1573,N_14719,N_14971);
nor UO_1574 (O_1574,N_14846,N_14793);
nand UO_1575 (O_1575,N_14881,N_14875);
nand UO_1576 (O_1576,N_14980,N_14705);
nand UO_1577 (O_1577,N_14908,N_14946);
or UO_1578 (O_1578,N_14936,N_14943);
nand UO_1579 (O_1579,N_14781,N_14782);
or UO_1580 (O_1580,N_14987,N_14708);
nand UO_1581 (O_1581,N_14704,N_14752);
nor UO_1582 (O_1582,N_14727,N_14886);
or UO_1583 (O_1583,N_14788,N_14778);
and UO_1584 (O_1584,N_14852,N_14725);
or UO_1585 (O_1585,N_14961,N_14843);
xnor UO_1586 (O_1586,N_14938,N_14850);
and UO_1587 (O_1587,N_14923,N_14882);
nand UO_1588 (O_1588,N_14957,N_14969);
xor UO_1589 (O_1589,N_14960,N_14715);
nor UO_1590 (O_1590,N_14824,N_14877);
and UO_1591 (O_1591,N_14765,N_14888);
and UO_1592 (O_1592,N_14888,N_14905);
xnor UO_1593 (O_1593,N_14736,N_14726);
nand UO_1594 (O_1594,N_14977,N_14946);
xor UO_1595 (O_1595,N_14793,N_14790);
xnor UO_1596 (O_1596,N_14842,N_14754);
and UO_1597 (O_1597,N_14836,N_14879);
xor UO_1598 (O_1598,N_14905,N_14717);
xor UO_1599 (O_1599,N_14969,N_14887);
and UO_1600 (O_1600,N_14965,N_14796);
nand UO_1601 (O_1601,N_14954,N_14922);
nor UO_1602 (O_1602,N_14704,N_14969);
or UO_1603 (O_1603,N_14749,N_14922);
nor UO_1604 (O_1604,N_14850,N_14998);
or UO_1605 (O_1605,N_14960,N_14862);
nand UO_1606 (O_1606,N_14965,N_14943);
xnor UO_1607 (O_1607,N_14909,N_14764);
nor UO_1608 (O_1608,N_14893,N_14731);
and UO_1609 (O_1609,N_14899,N_14762);
nor UO_1610 (O_1610,N_14718,N_14865);
xnor UO_1611 (O_1611,N_14709,N_14714);
nand UO_1612 (O_1612,N_14934,N_14736);
or UO_1613 (O_1613,N_14894,N_14803);
nand UO_1614 (O_1614,N_14880,N_14876);
or UO_1615 (O_1615,N_14921,N_14871);
xor UO_1616 (O_1616,N_14785,N_14825);
or UO_1617 (O_1617,N_14723,N_14853);
and UO_1618 (O_1618,N_14787,N_14970);
xor UO_1619 (O_1619,N_14947,N_14730);
nand UO_1620 (O_1620,N_14952,N_14905);
nand UO_1621 (O_1621,N_14742,N_14709);
nand UO_1622 (O_1622,N_14844,N_14933);
nand UO_1623 (O_1623,N_14755,N_14774);
nand UO_1624 (O_1624,N_14731,N_14958);
xnor UO_1625 (O_1625,N_14819,N_14979);
nand UO_1626 (O_1626,N_14859,N_14811);
or UO_1627 (O_1627,N_14785,N_14816);
or UO_1628 (O_1628,N_14824,N_14757);
nand UO_1629 (O_1629,N_14798,N_14788);
xor UO_1630 (O_1630,N_14783,N_14849);
nor UO_1631 (O_1631,N_14865,N_14723);
nor UO_1632 (O_1632,N_14865,N_14827);
nand UO_1633 (O_1633,N_14791,N_14883);
nor UO_1634 (O_1634,N_14703,N_14895);
or UO_1635 (O_1635,N_14852,N_14853);
xnor UO_1636 (O_1636,N_14998,N_14841);
nand UO_1637 (O_1637,N_14728,N_14759);
xnor UO_1638 (O_1638,N_14813,N_14727);
nor UO_1639 (O_1639,N_14809,N_14952);
nand UO_1640 (O_1640,N_14774,N_14970);
or UO_1641 (O_1641,N_14748,N_14899);
xnor UO_1642 (O_1642,N_14903,N_14935);
or UO_1643 (O_1643,N_14874,N_14775);
or UO_1644 (O_1644,N_14848,N_14709);
nand UO_1645 (O_1645,N_14817,N_14752);
nor UO_1646 (O_1646,N_14854,N_14769);
and UO_1647 (O_1647,N_14807,N_14845);
and UO_1648 (O_1648,N_14742,N_14766);
nor UO_1649 (O_1649,N_14887,N_14979);
or UO_1650 (O_1650,N_14905,N_14921);
nor UO_1651 (O_1651,N_14710,N_14920);
and UO_1652 (O_1652,N_14854,N_14864);
nor UO_1653 (O_1653,N_14758,N_14986);
xnor UO_1654 (O_1654,N_14837,N_14818);
nor UO_1655 (O_1655,N_14891,N_14753);
xor UO_1656 (O_1656,N_14864,N_14738);
nor UO_1657 (O_1657,N_14863,N_14979);
or UO_1658 (O_1658,N_14787,N_14941);
xnor UO_1659 (O_1659,N_14746,N_14850);
nor UO_1660 (O_1660,N_14775,N_14857);
or UO_1661 (O_1661,N_14984,N_14872);
xor UO_1662 (O_1662,N_14756,N_14866);
or UO_1663 (O_1663,N_14717,N_14797);
and UO_1664 (O_1664,N_14881,N_14730);
nor UO_1665 (O_1665,N_14789,N_14791);
and UO_1666 (O_1666,N_14799,N_14889);
xor UO_1667 (O_1667,N_14766,N_14925);
xnor UO_1668 (O_1668,N_14944,N_14935);
or UO_1669 (O_1669,N_14931,N_14716);
or UO_1670 (O_1670,N_14728,N_14770);
nand UO_1671 (O_1671,N_14766,N_14843);
xnor UO_1672 (O_1672,N_14933,N_14975);
and UO_1673 (O_1673,N_14887,N_14724);
xnor UO_1674 (O_1674,N_14729,N_14728);
and UO_1675 (O_1675,N_14984,N_14941);
and UO_1676 (O_1676,N_14907,N_14861);
and UO_1677 (O_1677,N_14716,N_14795);
xnor UO_1678 (O_1678,N_14975,N_14913);
xor UO_1679 (O_1679,N_14702,N_14724);
and UO_1680 (O_1680,N_14999,N_14943);
and UO_1681 (O_1681,N_14775,N_14773);
xnor UO_1682 (O_1682,N_14810,N_14819);
nand UO_1683 (O_1683,N_14814,N_14875);
and UO_1684 (O_1684,N_14928,N_14988);
nor UO_1685 (O_1685,N_14711,N_14803);
or UO_1686 (O_1686,N_14921,N_14975);
nand UO_1687 (O_1687,N_14934,N_14942);
xnor UO_1688 (O_1688,N_14732,N_14957);
and UO_1689 (O_1689,N_14840,N_14924);
or UO_1690 (O_1690,N_14798,N_14841);
xor UO_1691 (O_1691,N_14865,N_14834);
xor UO_1692 (O_1692,N_14946,N_14860);
nand UO_1693 (O_1693,N_14961,N_14842);
xor UO_1694 (O_1694,N_14967,N_14950);
nor UO_1695 (O_1695,N_14830,N_14795);
and UO_1696 (O_1696,N_14967,N_14938);
and UO_1697 (O_1697,N_14968,N_14994);
nor UO_1698 (O_1698,N_14927,N_14775);
xnor UO_1699 (O_1699,N_14843,N_14753);
nand UO_1700 (O_1700,N_14781,N_14780);
or UO_1701 (O_1701,N_14704,N_14983);
nor UO_1702 (O_1702,N_14882,N_14868);
xnor UO_1703 (O_1703,N_14799,N_14840);
nor UO_1704 (O_1704,N_14948,N_14763);
or UO_1705 (O_1705,N_14970,N_14973);
and UO_1706 (O_1706,N_14811,N_14987);
and UO_1707 (O_1707,N_14910,N_14955);
xnor UO_1708 (O_1708,N_14713,N_14750);
and UO_1709 (O_1709,N_14963,N_14881);
nor UO_1710 (O_1710,N_14926,N_14897);
nor UO_1711 (O_1711,N_14983,N_14918);
nor UO_1712 (O_1712,N_14768,N_14785);
xnor UO_1713 (O_1713,N_14806,N_14986);
and UO_1714 (O_1714,N_14779,N_14751);
xor UO_1715 (O_1715,N_14744,N_14925);
xnor UO_1716 (O_1716,N_14750,N_14767);
and UO_1717 (O_1717,N_14893,N_14761);
nor UO_1718 (O_1718,N_14703,N_14880);
xor UO_1719 (O_1719,N_14903,N_14709);
and UO_1720 (O_1720,N_14750,N_14801);
nor UO_1721 (O_1721,N_14778,N_14931);
nand UO_1722 (O_1722,N_14881,N_14708);
nor UO_1723 (O_1723,N_14856,N_14989);
xor UO_1724 (O_1724,N_14702,N_14904);
nor UO_1725 (O_1725,N_14785,N_14858);
xnor UO_1726 (O_1726,N_14935,N_14933);
nor UO_1727 (O_1727,N_14704,N_14919);
xnor UO_1728 (O_1728,N_14963,N_14813);
nand UO_1729 (O_1729,N_14866,N_14906);
and UO_1730 (O_1730,N_14851,N_14781);
nor UO_1731 (O_1731,N_14963,N_14705);
nand UO_1732 (O_1732,N_14921,N_14818);
and UO_1733 (O_1733,N_14741,N_14994);
or UO_1734 (O_1734,N_14939,N_14954);
nand UO_1735 (O_1735,N_14717,N_14914);
or UO_1736 (O_1736,N_14999,N_14893);
xor UO_1737 (O_1737,N_14796,N_14716);
nor UO_1738 (O_1738,N_14825,N_14898);
and UO_1739 (O_1739,N_14850,N_14865);
nand UO_1740 (O_1740,N_14854,N_14764);
or UO_1741 (O_1741,N_14931,N_14842);
nor UO_1742 (O_1742,N_14918,N_14856);
xor UO_1743 (O_1743,N_14796,N_14865);
or UO_1744 (O_1744,N_14806,N_14715);
nor UO_1745 (O_1745,N_14970,N_14916);
or UO_1746 (O_1746,N_14906,N_14940);
and UO_1747 (O_1747,N_14967,N_14959);
nand UO_1748 (O_1748,N_14752,N_14908);
or UO_1749 (O_1749,N_14757,N_14953);
nand UO_1750 (O_1750,N_14823,N_14713);
nor UO_1751 (O_1751,N_14909,N_14878);
xor UO_1752 (O_1752,N_14904,N_14719);
nor UO_1753 (O_1753,N_14704,N_14954);
nor UO_1754 (O_1754,N_14893,N_14920);
or UO_1755 (O_1755,N_14707,N_14767);
nand UO_1756 (O_1756,N_14784,N_14709);
nor UO_1757 (O_1757,N_14745,N_14797);
and UO_1758 (O_1758,N_14965,N_14961);
and UO_1759 (O_1759,N_14976,N_14701);
and UO_1760 (O_1760,N_14847,N_14992);
xnor UO_1761 (O_1761,N_14943,N_14985);
nand UO_1762 (O_1762,N_14706,N_14909);
nand UO_1763 (O_1763,N_14834,N_14971);
or UO_1764 (O_1764,N_14807,N_14754);
or UO_1765 (O_1765,N_14836,N_14730);
nor UO_1766 (O_1766,N_14720,N_14937);
or UO_1767 (O_1767,N_14972,N_14752);
xnor UO_1768 (O_1768,N_14724,N_14791);
and UO_1769 (O_1769,N_14911,N_14763);
nand UO_1770 (O_1770,N_14766,N_14802);
nand UO_1771 (O_1771,N_14765,N_14734);
or UO_1772 (O_1772,N_14712,N_14874);
nor UO_1773 (O_1773,N_14866,N_14819);
and UO_1774 (O_1774,N_14712,N_14968);
and UO_1775 (O_1775,N_14754,N_14917);
nor UO_1776 (O_1776,N_14746,N_14788);
and UO_1777 (O_1777,N_14758,N_14898);
xor UO_1778 (O_1778,N_14887,N_14766);
or UO_1779 (O_1779,N_14940,N_14913);
nand UO_1780 (O_1780,N_14730,N_14939);
nand UO_1781 (O_1781,N_14883,N_14966);
nand UO_1782 (O_1782,N_14836,N_14761);
or UO_1783 (O_1783,N_14779,N_14960);
or UO_1784 (O_1784,N_14804,N_14895);
and UO_1785 (O_1785,N_14830,N_14801);
nor UO_1786 (O_1786,N_14713,N_14879);
nand UO_1787 (O_1787,N_14706,N_14759);
and UO_1788 (O_1788,N_14881,N_14817);
xnor UO_1789 (O_1789,N_14841,N_14769);
xor UO_1790 (O_1790,N_14966,N_14750);
nand UO_1791 (O_1791,N_14964,N_14999);
nor UO_1792 (O_1792,N_14760,N_14845);
nor UO_1793 (O_1793,N_14714,N_14824);
nor UO_1794 (O_1794,N_14998,N_14981);
nor UO_1795 (O_1795,N_14788,N_14704);
and UO_1796 (O_1796,N_14830,N_14726);
xor UO_1797 (O_1797,N_14967,N_14876);
nand UO_1798 (O_1798,N_14883,N_14890);
nor UO_1799 (O_1799,N_14923,N_14931);
and UO_1800 (O_1800,N_14767,N_14943);
nand UO_1801 (O_1801,N_14705,N_14823);
nor UO_1802 (O_1802,N_14801,N_14965);
or UO_1803 (O_1803,N_14810,N_14809);
xor UO_1804 (O_1804,N_14858,N_14868);
and UO_1805 (O_1805,N_14740,N_14764);
and UO_1806 (O_1806,N_14939,N_14756);
nand UO_1807 (O_1807,N_14774,N_14843);
xor UO_1808 (O_1808,N_14787,N_14905);
nand UO_1809 (O_1809,N_14910,N_14707);
or UO_1810 (O_1810,N_14841,N_14729);
nand UO_1811 (O_1811,N_14821,N_14702);
nand UO_1812 (O_1812,N_14746,N_14890);
and UO_1813 (O_1813,N_14805,N_14881);
or UO_1814 (O_1814,N_14765,N_14939);
and UO_1815 (O_1815,N_14775,N_14722);
nor UO_1816 (O_1816,N_14899,N_14861);
or UO_1817 (O_1817,N_14928,N_14957);
nor UO_1818 (O_1818,N_14877,N_14984);
nor UO_1819 (O_1819,N_14786,N_14997);
xnor UO_1820 (O_1820,N_14719,N_14963);
nor UO_1821 (O_1821,N_14714,N_14829);
nor UO_1822 (O_1822,N_14866,N_14883);
and UO_1823 (O_1823,N_14994,N_14967);
or UO_1824 (O_1824,N_14771,N_14802);
and UO_1825 (O_1825,N_14751,N_14896);
nor UO_1826 (O_1826,N_14908,N_14794);
xor UO_1827 (O_1827,N_14783,N_14750);
nand UO_1828 (O_1828,N_14831,N_14805);
or UO_1829 (O_1829,N_14814,N_14869);
nor UO_1830 (O_1830,N_14991,N_14717);
nor UO_1831 (O_1831,N_14964,N_14746);
and UO_1832 (O_1832,N_14816,N_14802);
nand UO_1833 (O_1833,N_14851,N_14959);
nor UO_1834 (O_1834,N_14914,N_14839);
nor UO_1835 (O_1835,N_14771,N_14887);
or UO_1836 (O_1836,N_14962,N_14851);
nor UO_1837 (O_1837,N_14979,N_14909);
xnor UO_1838 (O_1838,N_14963,N_14913);
nor UO_1839 (O_1839,N_14898,N_14950);
nand UO_1840 (O_1840,N_14962,N_14742);
xor UO_1841 (O_1841,N_14857,N_14799);
or UO_1842 (O_1842,N_14870,N_14737);
nor UO_1843 (O_1843,N_14838,N_14968);
nand UO_1844 (O_1844,N_14984,N_14706);
nor UO_1845 (O_1845,N_14961,N_14919);
or UO_1846 (O_1846,N_14969,N_14898);
nand UO_1847 (O_1847,N_14768,N_14786);
nor UO_1848 (O_1848,N_14790,N_14818);
nand UO_1849 (O_1849,N_14860,N_14865);
or UO_1850 (O_1850,N_14912,N_14928);
or UO_1851 (O_1851,N_14816,N_14784);
or UO_1852 (O_1852,N_14890,N_14871);
nand UO_1853 (O_1853,N_14940,N_14886);
or UO_1854 (O_1854,N_14923,N_14943);
nor UO_1855 (O_1855,N_14993,N_14979);
or UO_1856 (O_1856,N_14820,N_14964);
or UO_1857 (O_1857,N_14949,N_14951);
and UO_1858 (O_1858,N_14932,N_14791);
xnor UO_1859 (O_1859,N_14916,N_14802);
or UO_1860 (O_1860,N_14757,N_14902);
nor UO_1861 (O_1861,N_14980,N_14906);
xnor UO_1862 (O_1862,N_14925,N_14883);
and UO_1863 (O_1863,N_14936,N_14853);
nor UO_1864 (O_1864,N_14833,N_14815);
nor UO_1865 (O_1865,N_14824,N_14930);
nand UO_1866 (O_1866,N_14912,N_14777);
xnor UO_1867 (O_1867,N_14819,N_14701);
nor UO_1868 (O_1868,N_14887,N_14977);
nand UO_1869 (O_1869,N_14891,N_14726);
or UO_1870 (O_1870,N_14964,N_14767);
nand UO_1871 (O_1871,N_14731,N_14842);
and UO_1872 (O_1872,N_14886,N_14709);
and UO_1873 (O_1873,N_14922,N_14854);
or UO_1874 (O_1874,N_14824,N_14908);
and UO_1875 (O_1875,N_14882,N_14844);
and UO_1876 (O_1876,N_14946,N_14787);
or UO_1877 (O_1877,N_14825,N_14986);
xor UO_1878 (O_1878,N_14939,N_14847);
nor UO_1879 (O_1879,N_14710,N_14982);
xnor UO_1880 (O_1880,N_14869,N_14963);
nor UO_1881 (O_1881,N_14837,N_14934);
xor UO_1882 (O_1882,N_14744,N_14928);
xnor UO_1883 (O_1883,N_14745,N_14841);
or UO_1884 (O_1884,N_14995,N_14710);
and UO_1885 (O_1885,N_14934,N_14813);
or UO_1886 (O_1886,N_14749,N_14894);
xnor UO_1887 (O_1887,N_14709,N_14806);
and UO_1888 (O_1888,N_14745,N_14726);
and UO_1889 (O_1889,N_14892,N_14730);
xnor UO_1890 (O_1890,N_14780,N_14900);
xnor UO_1891 (O_1891,N_14828,N_14881);
xnor UO_1892 (O_1892,N_14916,N_14866);
and UO_1893 (O_1893,N_14710,N_14871);
nor UO_1894 (O_1894,N_14808,N_14930);
nand UO_1895 (O_1895,N_14868,N_14865);
xor UO_1896 (O_1896,N_14940,N_14812);
xor UO_1897 (O_1897,N_14836,N_14748);
nor UO_1898 (O_1898,N_14835,N_14773);
or UO_1899 (O_1899,N_14755,N_14726);
or UO_1900 (O_1900,N_14894,N_14737);
nor UO_1901 (O_1901,N_14939,N_14737);
xnor UO_1902 (O_1902,N_14802,N_14896);
xor UO_1903 (O_1903,N_14952,N_14894);
or UO_1904 (O_1904,N_14740,N_14784);
xnor UO_1905 (O_1905,N_14870,N_14725);
and UO_1906 (O_1906,N_14979,N_14807);
and UO_1907 (O_1907,N_14788,N_14889);
nor UO_1908 (O_1908,N_14806,N_14942);
or UO_1909 (O_1909,N_14722,N_14749);
and UO_1910 (O_1910,N_14967,N_14799);
and UO_1911 (O_1911,N_14989,N_14985);
nor UO_1912 (O_1912,N_14811,N_14723);
or UO_1913 (O_1913,N_14976,N_14822);
nor UO_1914 (O_1914,N_14850,N_14703);
nor UO_1915 (O_1915,N_14922,N_14914);
and UO_1916 (O_1916,N_14742,N_14801);
or UO_1917 (O_1917,N_14812,N_14942);
and UO_1918 (O_1918,N_14930,N_14951);
nor UO_1919 (O_1919,N_14828,N_14891);
and UO_1920 (O_1920,N_14953,N_14768);
nand UO_1921 (O_1921,N_14821,N_14948);
nor UO_1922 (O_1922,N_14964,N_14720);
nor UO_1923 (O_1923,N_14935,N_14833);
xor UO_1924 (O_1924,N_14963,N_14816);
and UO_1925 (O_1925,N_14883,N_14808);
or UO_1926 (O_1926,N_14997,N_14802);
or UO_1927 (O_1927,N_14944,N_14955);
or UO_1928 (O_1928,N_14770,N_14869);
nor UO_1929 (O_1929,N_14895,N_14805);
nor UO_1930 (O_1930,N_14741,N_14838);
or UO_1931 (O_1931,N_14997,N_14763);
xnor UO_1932 (O_1932,N_14742,N_14783);
and UO_1933 (O_1933,N_14850,N_14963);
xor UO_1934 (O_1934,N_14812,N_14768);
xnor UO_1935 (O_1935,N_14991,N_14725);
or UO_1936 (O_1936,N_14788,N_14727);
xnor UO_1937 (O_1937,N_14723,N_14824);
nand UO_1938 (O_1938,N_14841,N_14896);
nand UO_1939 (O_1939,N_14944,N_14718);
xor UO_1940 (O_1940,N_14741,N_14706);
or UO_1941 (O_1941,N_14702,N_14804);
and UO_1942 (O_1942,N_14960,N_14753);
and UO_1943 (O_1943,N_14945,N_14942);
xor UO_1944 (O_1944,N_14908,N_14979);
xnor UO_1945 (O_1945,N_14862,N_14853);
nor UO_1946 (O_1946,N_14962,N_14716);
and UO_1947 (O_1947,N_14717,N_14702);
nand UO_1948 (O_1948,N_14802,N_14960);
xor UO_1949 (O_1949,N_14768,N_14822);
nand UO_1950 (O_1950,N_14841,N_14948);
nand UO_1951 (O_1951,N_14910,N_14713);
nor UO_1952 (O_1952,N_14972,N_14727);
xor UO_1953 (O_1953,N_14856,N_14947);
and UO_1954 (O_1954,N_14939,N_14943);
or UO_1955 (O_1955,N_14948,N_14703);
nor UO_1956 (O_1956,N_14788,N_14848);
or UO_1957 (O_1957,N_14911,N_14708);
nand UO_1958 (O_1958,N_14708,N_14947);
nand UO_1959 (O_1959,N_14824,N_14975);
and UO_1960 (O_1960,N_14895,N_14996);
and UO_1961 (O_1961,N_14881,N_14719);
nor UO_1962 (O_1962,N_14859,N_14890);
nand UO_1963 (O_1963,N_14822,N_14804);
nand UO_1964 (O_1964,N_14987,N_14738);
or UO_1965 (O_1965,N_14778,N_14834);
or UO_1966 (O_1966,N_14968,N_14965);
nor UO_1967 (O_1967,N_14808,N_14779);
xnor UO_1968 (O_1968,N_14866,N_14776);
and UO_1969 (O_1969,N_14724,N_14939);
nor UO_1970 (O_1970,N_14890,N_14807);
nor UO_1971 (O_1971,N_14969,N_14926);
nor UO_1972 (O_1972,N_14948,N_14897);
and UO_1973 (O_1973,N_14736,N_14906);
or UO_1974 (O_1974,N_14812,N_14976);
nand UO_1975 (O_1975,N_14985,N_14764);
or UO_1976 (O_1976,N_14835,N_14976);
nand UO_1977 (O_1977,N_14851,N_14715);
and UO_1978 (O_1978,N_14765,N_14849);
or UO_1979 (O_1979,N_14886,N_14702);
and UO_1980 (O_1980,N_14876,N_14952);
nor UO_1981 (O_1981,N_14966,N_14744);
nand UO_1982 (O_1982,N_14710,N_14980);
nand UO_1983 (O_1983,N_14810,N_14958);
xor UO_1984 (O_1984,N_14995,N_14946);
or UO_1985 (O_1985,N_14883,N_14910);
nor UO_1986 (O_1986,N_14805,N_14740);
nand UO_1987 (O_1987,N_14981,N_14751);
nor UO_1988 (O_1988,N_14964,N_14944);
and UO_1989 (O_1989,N_14768,N_14807);
or UO_1990 (O_1990,N_14963,N_14915);
and UO_1991 (O_1991,N_14849,N_14889);
xor UO_1992 (O_1992,N_14904,N_14876);
nand UO_1993 (O_1993,N_14890,N_14767);
or UO_1994 (O_1994,N_14972,N_14780);
nand UO_1995 (O_1995,N_14920,N_14892);
nand UO_1996 (O_1996,N_14814,N_14897);
nor UO_1997 (O_1997,N_14889,N_14791);
xnor UO_1998 (O_1998,N_14909,N_14995);
and UO_1999 (O_1999,N_14732,N_14846);
endmodule