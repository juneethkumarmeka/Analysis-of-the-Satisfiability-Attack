module basic_500_3000_500_4_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_19,In_464);
nor U1 (N_1,In_114,In_34);
and U2 (N_2,In_460,In_363);
nand U3 (N_3,In_60,In_158);
nor U4 (N_4,In_32,In_52);
and U5 (N_5,In_488,In_246);
nor U6 (N_6,In_344,In_226);
or U7 (N_7,In_35,In_339);
nor U8 (N_8,In_210,In_200);
or U9 (N_9,In_404,In_175);
and U10 (N_10,In_438,In_316);
xor U11 (N_11,In_391,In_94);
nor U12 (N_12,In_69,In_231);
and U13 (N_13,In_66,In_394);
nor U14 (N_14,In_287,In_173);
nor U15 (N_15,In_365,In_112);
or U16 (N_16,In_352,In_4);
nor U17 (N_17,In_25,In_189);
or U18 (N_18,In_197,In_380);
nand U19 (N_19,In_355,In_169);
and U20 (N_20,In_468,In_240);
or U21 (N_21,In_9,In_342);
or U22 (N_22,In_259,In_469);
nor U23 (N_23,In_194,In_149);
nor U24 (N_24,In_164,In_284);
nor U25 (N_25,In_178,In_136);
or U26 (N_26,In_38,In_470);
or U27 (N_27,In_228,In_386);
and U28 (N_28,In_309,In_249);
or U29 (N_29,In_459,In_304);
and U30 (N_30,In_268,In_426);
nor U31 (N_31,In_446,In_491);
nor U32 (N_32,In_87,In_224);
and U33 (N_33,In_241,In_92);
and U34 (N_34,In_98,In_239);
nand U35 (N_35,In_418,In_190);
nand U36 (N_36,In_367,In_95);
and U37 (N_37,In_408,In_429);
nand U38 (N_38,In_8,In_440);
nor U39 (N_39,In_67,In_122);
or U40 (N_40,In_117,In_337);
xor U41 (N_41,In_91,In_78);
or U42 (N_42,In_320,In_46);
and U43 (N_43,In_144,In_244);
nand U44 (N_44,In_218,In_456);
and U45 (N_45,In_319,In_230);
nand U46 (N_46,In_195,In_314);
xor U47 (N_47,In_0,In_192);
nor U48 (N_48,In_214,In_444);
or U49 (N_49,In_286,In_261);
nand U50 (N_50,In_274,In_361);
or U51 (N_51,In_97,In_484);
nor U52 (N_52,In_420,In_250);
nand U53 (N_53,In_366,In_223);
nor U54 (N_54,In_166,In_351);
or U55 (N_55,In_74,In_350);
and U56 (N_56,In_42,In_400);
nand U57 (N_57,In_237,In_119);
and U58 (N_58,In_248,In_265);
or U59 (N_59,In_70,In_81);
nor U60 (N_60,In_152,In_292);
and U61 (N_61,In_13,In_49);
and U62 (N_62,In_354,In_102);
and U63 (N_63,In_289,In_76);
and U64 (N_64,In_346,In_306);
nor U65 (N_65,In_439,In_121);
nand U66 (N_66,In_61,In_315);
or U67 (N_67,In_196,In_308);
nand U68 (N_68,In_193,In_495);
nor U69 (N_69,In_353,In_130);
nor U70 (N_70,In_311,In_139);
or U71 (N_71,In_419,In_123);
nand U72 (N_72,In_243,In_232);
and U73 (N_73,In_43,In_465);
nand U74 (N_74,In_103,In_160);
and U75 (N_75,In_312,In_211);
nor U76 (N_76,In_82,In_148);
or U77 (N_77,In_180,In_23);
nand U78 (N_78,In_168,In_37);
nand U79 (N_79,In_402,In_176);
and U80 (N_80,In_267,In_137);
or U81 (N_81,In_397,In_55);
nand U82 (N_82,In_405,In_255);
and U83 (N_83,In_179,In_454);
nand U84 (N_84,In_296,In_343);
nand U85 (N_85,In_452,In_475);
nor U86 (N_86,In_15,In_22);
nand U87 (N_87,In_104,In_39);
or U88 (N_88,In_428,In_409);
or U89 (N_89,In_480,In_234);
nand U90 (N_90,In_172,In_323);
or U91 (N_91,In_256,In_263);
nor U92 (N_92,In_5,In_435);
and U93 (N_93,In_448,In_299);
and U94 (N_94,In_421,In_340);
nor U95 (N_95,In_151,In_177);
nor U96 (N_96,In_254,In_145);
and U97 (N_97,In_257,In_411);
nor U98 (N_98,In_235,In_389);
and U99 (N_99,In_202,In_467);
and U100 (N_100,In_31,In_364);
or U101 (N_101,In_75,In_424);
nand U102 (N_102,In_154,In_203);
or U103 (N_103,In_146,In_71);
or U104 (N_104,In_163,In_381);
nand U105 (N_105,In_310,In_115);
nand U106 (N_106,In_253,In_415);
or U107 (N_107,In_159,In_291);
nand U108 (N_108,In_118,In_184);
nand U109 (N_109,In_251,In_450);
or U110 (N_110,In_165,In_479);
and U111 (N_111,In_417,In_264);
and U112 (N_112,In_79,In_282);
or U113 (N_113,In_345,In_432);
and U114 (N_114,In_157,In_116);
nor U115 (N_115,In_212,In_276);
nor U116 (N_116,In_124,In_161);
nand U117 (N_117,In_490,In_16);
nor U118 (N_118,In_455,In_478);
or U119 (N_119,In_131,In_412);
nor U120 (N_120,In_225,In_398);
and U121 (N_121,In_278,In_209);
and U122 (N_122,In_474,In_390);
xnor U123 (N_123,In_403,In_477);
nand U124 (N_124,In_392,In_462);
nor U125 (N_125,In_50,In_324);
nand U126 (N_126,In_167,In_44);
nor U127 (N_127,In_476,In_199);
nor U128 (N_128,In_285,In_187);
nand U129 (N_129,In_373,In_301);
or U130 (N_130,In_499,In_105);
or U131 (N_131,In_185,In_442);
nor U132 (N_132,In_96,In_362);
or U133 (N_133,In_280,In_383);
nand U134 (N_134,In_7,In_325);
nor U135 (N_135,In_86,In_422);
or U136 (N_136,In_28,In_85);
xor U137 (N_137,In_84,In_29);
nor U138 (N_138,In_229,In_247);
nor U139 (N_139,In_242,In_57);
nand U140 (N_140,In_300,In_191);
or U141 (N_141,In_425,In_277);
nor U142 (N_142,In_6,In_3);
or U143 (N_143,In_334,In_335);
and U144 (N_144,In_414,In_64);
and U145 (N_145,In_332,In_447);
or U146 (N_146,In_449,In_407);
and U147 (N_147,In_17,In_215);
and U148 (N_148,In_483,In_376);
and U149 (N_149,In_378,In_321);
xor U150 (N_150,In_134,In_36);
and U151 (N_151,In_107,In_431);
and U152 (N_152,In_140,In_341);
nor U153 (N_153,In_150,In_328);
and U154 (N_154,In_106,In_377);
and U155 (N_155,In_359,In_100);
or U156 (N_156,In_348,In_399);
and U157 (N_157,In_436,In_283);
or U158 (N_158,In_497,In_443);
and U159 (N_159,In_153,In_80);
and U160 (N_160,In_138,In_269);
nand U161 (N_161,In_492,In_24);
and U162 (N_162,In_385,In_368);
and U163 (N_163,In_260,In_349);
nor U164 (N_164,In_427,In_481);
and U165 (N_165,In_207,In_88);
nand U166 (N_166,In_494,In_305);
nor U167 (N_167,In_54,In_382);
nor U168 (N_168,In_132,In_441);
and U169 (N_169,In_1,In_208);
or U170 (N_170,In_93,In_496);
xnor U171 (N_171,In_222,In_182);
and U172 (N_172,In_198,In_206);
and U173 (N_173,In_338,In_77);
nor U174 (N_174,In_135,In_220);
nand U175 (N_175,In_293,In_11);
nand U176 (N_176,In_10,In_143);
nand U177 (N_177,In_72,In_453);
nand U178 (N_178,In_47,In_374);
or U179 (N_179,In_487,In_90);
and U180 (N_180,In_410,In_99);
nand U181 (N_181,In_273,In_384);
and U182 (N_182,In_110,In_489);
or U183 (N_183,In_233,In_396);
or U184 (N_184,In_14,In_120);
nor U185 (N_185,In_245,In_387);
or U186 (N_186,In_473,In_188);
nand U187 (N_187,In_295,In_451);
and U188 (N_188,In_485,In_329);
and U189 (N_189,In_457,In_371);
or U190 (N_190,In_471,In_358);
or U191 (N_191,In_434,In_51);
nand U192 (N_192,In_171,In_347);
nand U193 (N_193,In_27,In_430);
nor U194 (N_194,In_73,In_333);
nor U195 (N_195,In_461,In_181);
or U196 (N_196,In_318,In_109);
nor U197 (N_197,In_302,In_375);
or U198 (N_198,In_2,In_423);
and U199 (N_199,In_40,In_186);
and U200 (N_200,In_317,In_258);
nand U201 (N_201,In_463,In_356);
xnor U202 (N_202,In_58,In_327);
or U203 (N_203,In_482,In_65);
or U204 (N_204,In_413,In_238);
nand U205 (N_205,In_205,In_156);
nor U206 (N_206,In_155,In_108);
or U207 (N_207,In_113,In_59);
xor U208 (N_208,In_307,In_204);
nor U209 (N_209,In_458,In_128);
and U210 (N_210,In_252,In_227);
nand U211 (N_211,In_20,In_326);
nand U212 (N_212,In_21,In_288);
and U213 (N_213,In_162,In_48);
nor U214 (N_214,In_393,In_217);
nor U215 (N_215,In_336,In_221);
nand U216 (N_216,In_26,In_493);
and U217 (N_217,In_379,In_89);
or U218 (N_218,In_33,In_313);
and U219 (N_219,In_416,In_216);
nand U220 (N_220,In_433,In_56);
nand U221 (N_221,In_262,In_236);
nor U222 (N_222,In_360,In_30);
nand U223 (N_223,In_18,In_445);
nand U224 (N_224,In_127,In_303);
and U225 (N_225,In_281,In_101);
nand U226 (N_226,In_272,In_466);
or U227 (N_227,In_322,In_388);
and U228 (N_228,In_174,In_290);
nand U229 (N_229,In_68,In_498);
or U230 (N_230,In_486,In_62);
and U231 (N_231,In_406,In_142);
or U232 (N_232,In_331,In_45);
or U233 (N_233,In_12,In_63);
nand U234 (N_234,In_294,In_370);
nor U235 (N_235,In_369,In_275);
nand U236 (N_236,In_401,In_297);
or U237 (N_237,In_472,In_141);
or U238 (N_238,In_83,In_213);
nand U239 (N_239,In_129,In_266);
nor U240 (N_240,In_170,In_330);
and U241 (N_241,In_279,In_53);
or U242 (N_242,In_271,In_111);
nand U243 (N_243,In_201,In_298);
nor U244 (N_244,In_125,In_437);
xor U245 (N_245,In_41,In_126);
and U246 (N_246,In_372,In_183);
and U247 (N_247,In_357,In_270);
nor U248 (N_248,In_147,In_133);
xor U249 (N_249,In_395,In_219);
or U250 (N_250,In_484,In_379);
nand U251 (N_251,In_397,In_121);
nand U252 (N_252,In_425,In_371);
and U253 (N_253,In_246,In_194);
nand U254 (N_254,In_489,In_417);
nand U255 (N_255,In_294,In_398);
or U256 (N_256,In_447,In_29);
nand U257 (N_257,In_160,In_389);
nor U258 (N_258,In_60,In_226);
or U259 (N_259,In_94,In_392);
nand U260 (N_260,In_111,In_166);
nand U261 (N_261,In_463,In_80);
or U262 (N_262,In_441,In_22);
or U263 (N_263,In_355,In_398);
nor U264 (N_264,In_270,In_191);
and U265 (N_265,In_46,In_377);
nor U266 (N_266,In_14,In_110);
and U267 (N_267,In_477,In_338);
or U268 (N_268,In_196,In_134);
nand U269 (N_269,In_106,In_368);
and U270 (N_270,In_175,In_489);
and U271 (N_271,In_297,In_443);
or U272 (N_272,In_140,In_141);
or U273 (N_273,In_479,In_176);
and U274 (N_274,In_323,In_366);
nand U275 (N_275,In_484,In_457);
nor U276 (N_276,In_67,In_354);
and U277 (N_277,In_72,In_470);
nand U278 (N_278,In_128,In_481);
nor U279 (N_279,In_192,In_455);
nor U280 (N_280,In_281,In_62);
nand U281 (N_281,In_380,In_376);
nor U282 (N_282,In_242,In_87);
nand U283 (N_283,In_82,In_427);
nor U284 (N_284,In_62,In_5);
or U285 (N_285,In_277,In_438);
or U286 (N_286,In_201,In_303);
nand U287 (N_287,In_457,In_34);
or U288 (N_288,In_358,In_287);
or U289 (N_289,In_450,In_71);
nand U290 (N_290,In_70,In_117);
nor U291 (N_291,In_238,In_304);
or U292 (N_292,In_496,In_55);
and U293 (N_293,In_346,In_11);
xnor U294 (N_294,In_118,In_359);
nand U295 (N_295,In_202,In_296);
and U296 (N_296,In_263,In_269);
or U297 (N_297,In_282,In_71);
nand U298 (N_298,In_44,In_293);
nor U299 (N_299,In_148,In_177);
nor U300 (N_300,In_178,In_311);
or U301 (N_301,In_31,In_151);
nand U302 (N_302,In_303,In_111);
nand U303 (N_303,In_396,In_53);
nor U304 (N_304,In_376,In_400);
or U305 (N_305,In_139,In_135);
nor U306 (N_306,In_354,In_170);
nor U307 (N_307,In_210,In_353);
and U308 (N_308,In_206,In_93);
or U309 (N_309,In_129,In_137);
nor U310 (N_310,In_350,In_327);
and U311 (N_311,In_198,In_414);
nand U312 (N_312,In_150,In_132);
or U313 (N_313,In_119,In_453);
or U314 (N_314,In_378,In_299);
nor U315 (N_315,In_74,In_406);
and U316 (N_316,In_54,In_100);
and U317 (N_317,In_241,In_65);
and U318 (N_318,In_60,In_222);
and U319 (N_319,In_115,In_356);
nand U320 (N_320,In_40,In_284);
nand U321 (N_321,In_381,In_458);
and U322 (N_322,In_480,In_49);
nor U323 (N_323,In_190,In_440);
nand U324 (N_324,In_358,In_131);
nand U325 (N_325,In_318,In_433);
and U326 (N_326,In_241,In_199);
nor U327 (N_327,In_140,In_396);
or U328 (N_328,In_381,In_277);
or U329 (N_329,In_496,In_295);
nor U330 (N_330,In_458,In_372);
nor U331 (N_331,In_346,In_261);
or U332 (N_332,In_0,In_468);
or U333 (N_333,In_467,In_338);
and U334 (N_334,In_190,In_335);
or U335 (N_335,In_279,In_142);
nor U336 (N_336,In_467,In_264);
or U337 (N_337,In_222,In_361);
and U338 (N_338,In_188,In_161);
or U339 (N_339,In_20,In_231);
nor U340 (N_340,In_50,In_58);
and U341 (N_341,In_81,In_46);
or U342 (N_342,In_340,In_30);
nor U343 (N_343,In_122,In_172);
nand U344 (N_344,In_457,In_188);
and U345 (N_345,In_436,In_177);
and U346 (N_346,In_153,In_4);
nor U347 (N_347,In_438,In_247);
nor U348 (N_348,In_333,In_308);
and U349 (N_349,In_23,In_108);
or U350 (N_350,In_226,In_455);
or U351 (N_351,In_410,In_403);
nor U352 (N_352,In_447,In_149);
and U353 (N_353,In_168,In_273);
nor U354 (N_354,In_189,In_279);
nand U355 (N_355,In_208,In_293);
and U356 (N_356,In_290,In_63);
nor U357 (N_357,In_355,In_209);
or U358 (N_358,In_289,In_452);
xor U359 (N_359,In_483,In_251);
or U360 (N_360,In_260,In_156);
nand U361 (N_361,In_430,In_489);
and U362 (N_362,In_337,In_389);
or U363 (N_363,In_167,In_73);
nand U364 (N_364,In_403,In_439);
or U365 (N_365,In_2,In_185);
and U366 (N_366,In_413,In_0);
nand U367 (N_367,In_247,In_78);
or U368 (N_368,In_219,In_60);
nand U369 (N_369,In_493,In_488);
or U370 (N_370,In_51,In_15);
and U371 (N_371,In_430,In_484);
nor U372 (N_372,In_314,In_55);
nand U373 (N_373,In_352,In_51);
and U374 (N_374,In_26,In_37);
or U375 (N_375,In_370,In_86);
and U376 (N_376,In_69,In_402);
nand U377 (N_377,In_73,In_484);
nand U378 (N_378,In_161,In_261);
nand U379 (N_379,In_288,In_246);
and U380 (N_380,In_341,In_230);
nor U381 (N_381,In_384,In_95);
xor U382 (N_382,In_184,In_228);
nor U383 (N_383,In_236,In_167);
and U384 (N_384,In_401,In_126);
and U385 (N_385,In_202,In_355);
or U386 (N_386,In_450,In_310);
nand U387 (N_387,In_284,In_309);
or U388 (N_388,In_333,In_381);
and U389 (N_389,In_215,In_273);
xor U390 (N_390,In_321,In_371);
or U391 (N_391,In_369,In_435);
nor U392 (N_392,In_453,In_14);
or U393 (N_393,In_256,In_449);
nor U394 (N_394,In_127,In_408);
or U395 (N_395,In_418,In_489);
or U396 (N_396,In_251,In_48);
and U397 (N_397,In_487,In_123);
nand U398 (N_398,In_309,In_310);
nor U399 (N_399,In_473,In_403);
or U400 (N_400,In_84,In_269);
and U401 (N_401,In_234,In_393);
nand U402 (N_402,In_205,In_70);
nor U403 (N_403,In_462,In_266);
and U404 (N_404,In_460,In_331);
nand U405 (N_405,In_412,In_490);
and U406 (N_406,In_298,In_110);
or U407 (N_407,In_407,In_46);
or U408 (N_408,In_72,In_368);
nand U409 (N_409,In_184,In_48);
nand U410 (N_410,In_425,In_140);
nor U411 (N_411,In_254,In_131);
or U412 (N_412,In_245,In_79);
nand U413 (N_413,In_453,In_448);
nand U414 (N_414,In_128,In_424);
nand U415 (N_415,In_96,In_353);
or U416 (N_416,In_86,In_335);
nand U417 (N_417,In_55,In_394);
nor U418 (N_418,In_375,In_389);
nor U419 (N_419,In_275,In_477);
nor U420 (N_420,In_470,In_348);
or U421 (N_421,In_493,In_180);
nor U422 (N_422,In_253,In_457);
nand U423 (N_423,In_251,In_458);
and U424 (N_424,In_382,In_159);
nor U425 (N_425,In_126,In_240);
or U426 (N_426,In_439,In_91);
nor U427 (N_427,In_328,In_45);
and U428 (N_428,In_407,In_488);
and U429 (N_429,In_337,In_91);
and U430 (N_430,In_10,In_211);
nand U431 (N_431,In_113,In_159);
nand U432 (N_432,In_353,In_341);
or U433 (N_433,In_22,In_48);
and U434 (N_434,In_121,In_142);
nor U435 (N_435,In_289,In_260);
nor U436 (N_436,In_362,In_480);
and U437 (N_437,In_437,In_171);
xor U438 (N_438,In_324,In_128);
nand U439 (N_439,In_145,In_132);
or U440 (N_440,In_277,In_184);
nand U441 (N_441,In_130,In_338);
or U442 (N_442,In_276,In_335);
nor U443 (N_443,In_2,In_248);
nor U444 (N_444,In_203,In_88);
or U445 (N_445,In_87,In_9);
or U446 (N_446,In_156,In_34);
or U447 (N_447,In_216,In_162);
or U448 (N_448,In_152,In_154);
nor U449 (N_449,In_41,In_238);
nor U450 (N_450,In_281,In_127);
nand U451 (N_451,In_370,In_216);
nand U452 (N_452,In_418,In_189);
nand U453 (N_453,In_369,In_30);
nand U454 (N_454,In_63,In_13);
and U455 (N_455,In_190,In_128);
or U456 (N_456,In_377,In_411);
nand U457 (N_457,In_370,In_318);
nand U458 (N_458,In_387,In_115);
or U459 (N_459,In_330,In_294);
or U460 (N_460,In_344,In_498);
and U461 (N_461,In_174,In_30);
and U462 (N_462,In_266,In_28);
and U463 (N_463,In_79,In_301);
nor U464 (N_464,In_205,In_319);
nor U465 (N_465,In_147,In_187);
nor U466 (N_466,In_399,In_485);
or U467 (N_467,In_101,In_347);
nand U468 (N_468,In_397,In_402);
or U469 (N_469,In_88,In_216);
and U470 (N_470,In_31,In_370);
or U471 (N_471,In_487,In_430);
nor U472 (N_472,In_84,In_358);
nor U473 (N_473,In_77,In_12);
and U474 (N_474,In_312,In_90);
and U475 (N_475,In_251,In_489);
nor U476 (N_476,In_118,In_20);
nor U477 (N_477,In_496,In_118);
or U478 (N_478,In_429,In_245);
and U479 (N_479,In_295,In_227);
and U480 (N_480,In_200,In_365);
nand U481 (N_481,In_178,In_397);
xnor U482 (N_482,In_28,In_219);
and U483 (N_483,In_22,In_284);
and U484 (N_484,In_161,In_100);
nand U485 (N_485,In_280,In_176);
or U486 (N_486,In_86,In_80);
nor U487 (N_487,In_469,In_360);
nand U488 (N_488,In_232,In_449);
or U489 (N_489,In_266,In_283);
and U490 (N_490,In_25,In_487);
nor U491 (N_491,In_131,In_101);
nor U492 (N_492,In_57,In_234);
nand U493 (N_493,In_416,In_212);
and U494 (N_494,In_249,In_173);
and U495 (N_495,In_387,In_409);
nor U496 (N_496,In_414,In_33);
or U497 (N_497,In_297,In_369);
nand U498 (N_498,In_91,In_343);
and U499 (N_499,In_435,In_89);
and U500 (N_500,In_496,In_422);
nor U501 (N_501,In_274,In_212);
nor U502 (N_502,In_397,In_257);
or U503 (N_503,In_402,In_14);
and U504 (N_504,In_332,In_476);
or U505 (N_505,In_333,In_103);
and U506 (N_506,In_248,In_432);
nor U507 (N_507,In_133,In_200);
nor U508 (N_508,In_423,In_113);
and U509 (N_509,In_155,In_408);
nand U510 (N_510,In_499,In_91);
nand U511 (N_511,In_304,In_297);
nand U512 (N_512,In_224,In_494);
or U513 (N_513,In_410,In_383);
and U514 (N_514,In_428,In_172);
nand U515 (N_515,In_362,In_499);
nand U516 (N_516,In_134,In_309);
nor U517 (N_517,In_240,In_402);
nor U518 (N_518,In_288,In_175);
nor U519 (N_519,In_7,In_2);
or U520 (N_520,In_304,In_187);
nor U521 (N_521,In_94,In_67);
or U522 (N_522,In_292,In_164);
nor U523 (N_523,In_356,In_462);
and U524 (N_524,In_193,In_405);
nand U525 (N_525,In_136,In_312);
or U526 (N_526,In_99,In_349);
nor U527 (N_527,In_442,In_363);
and U528 (N_528,In_157,In_481);
nor U529 (N_529,In_365,In_52);
xnor U530 (N_530,In_7,In_165);
or U531 (N_531,In_87,In_83);
nor U532 (N_532,In_280,In_91);
nor U533 (N_533,In_171,In_224);
nand U534 (N_534,In_192,In_31);
or U535 (N_535,In_216,In_191);
or U536 (N_536,In_112,In_124);
nand U537 (N_537,In_441,In_188);
nand U538 (N_538,In_116,In_75);
nand U539 (N_539,In_63,In_415);
nor U540 (N_540,In_5,In_271);
or U541 (N_541,In_213,In_372);
nor U542 (N_542,In_333,In_281);
and U543 (N_543,In_276,In_309);
and U544 (N_544,In_332,In_446);
or U545 (N_545,In_105,In_289);
nand U546 (N_546,In_169,In_407);
or U547 (N_547,In_332,In_105);
nand U548 (N_548,In_391,In_409);
and U549 (N_549,In_429,In_283);
nand U550 (N_550,In_73,In_181);
and U551 (N_551,In_23,In_365);
nor U552 (N_552,In_214,In_28);
and U553 (N_553,In_414,In_61);
or U554 (N_554,In_96,In_316);
nor U555 (N_555,In_163,In_72);
or U556 (N_556,In_396,In_408);
nand U557 (N_557,In_113,In_425);
nand U558 (N_558,In_107,In_184);
and U559 (N_559,In_137,In_197);
or U560 (N_560,In_211,In_435);
nor U561 (N_561,In_93,In_387);
or U562 (N_562,In_278,In_220);
nor U563 (N_563,In_324,In_331);
and U564 (N_564,In_473,In_36);
nand U565 (N_565,In_247,In_175);
xor U566 (N_566,In_450,In_199);
and U567 (N_567,In_307,In_6);
nand U568 (N_568,In_81,In_236);
or U569 (N_569,In_229,In_467);
nor U570 (N_570,In_236,In_51);
nand U571 (N_571,In_202,In_119);
nand U572 (N_572,In_28,In_42);
nand U573 (N_573,In_498,In_386);
nand U574 (N_574,In_125,In_348);
nand U575 (N_575,In_364,In_321);
nand U576 (N_576,In_55,In_9);
nand U577 (N_577,In_471,In_199);
nand U578 (N_578,In_219,In_189);
or U579 (N_579,In_58,In_242);
nand U580 (N_580,In_207,In_497);
or U581 (N_581,In_337,In_130);
nor U582 (N_582,In_83,In_465);
nor U583 (N_583,In_112,In_405);
and U584 (N_584,In_33,In_329);
nor U585 (N_585,In_266,In_79);
nand U586 (N_586,In_150,In_28);
and U587 (N_587,In_421,In_19);
and U588 (N_588,In_455,In_124);
nor U589 (N_589,In_456,In_410);
or U590 (N_590,In_476,In_149);
and U591 (N_591,In_146,In_13);
or U592 (N_592,In_355,In_350);
nor U593 (N_593,In_85,In_223);
and U594 (N_594,In_259,In_253);
or U595 (N_595,In_79,In_485);
nor U596 (N_596,In_359,In_474);
xnor U597 (N_597,In_153,In_202);
nand U598 (N_598,In_492,In_384);
and U599 (N_599,In_168,In_295);
nor U600 (N_600,In_395,In_224);
nor U601 (N_601,In_461,In_81);
nand U602 (N_602,In_204,In_150);
and U603 (N_603,In_40,In_26);
nand U604 (N_604,In_167,In_59);
or U605 (N_605,In_237,In_291);
nand U606 (N_606,In_498,In_346);
or U607 (N_607,In_274,In_265);
nand U608 (N_608,In_437,In_38);
or U609 (N_609,In_292,In_151);
nand U610 (N_610,In_70,In_455);
and U611 (N_611,In_264,In_307);
and U612 (N_612,In_105,In_473);
or U613 (N_613,In_37,In_12);
or U614 (N_614,In_484,In_150);
nand U615 (N_615,In_487,In_265);
nand U616 (N_616,In_97,In_498);
and U617 (N_617,In_420,In_454);
or U618 (N_618,In_330,In_122);
and U619 (N_619,In_105,In_389);
or U620 (N_620,In_444,In_485);
or U621 (N_621,In_195,In_463);
and U622 (N_622,In_461,In_170);
nand U623 (N_623,In_499,In_224);
nand U624 (N_624,In_156,In_219);
or U625 (N_625,In_366,In_276);
nand U626 (N_626,In_338,In_263);
and U627 (N_627,In_182,In_343);
and U628 (N_628,In_190,In_216);
and U629 (N_629,In_471,In_208);
or U630 (N_630,In_490,In_227);
xnor U631 (N_631,In_404,In_457);
and U632 (N_632,In_227,In_189);
or U633 (N_633,In_75,In_328);
or U634 (N_634,In_94,In_356);
nor U635 (N_635,In_89,In_42);
nor U636 (N_636,In_50,In_18);
nand U637 (N_637,In_16,In_342);
or U638 (N_638,In_451,In_57);
nor U639 (N_639,In_177,In_17);
nand U640 (N_640,In_165,In_312);
or U641 (N_641,In_308,In_96);
and U642 (N_642,In_225,In_113);
nor U643 (N_643,In_22,In_46);
and U644 (N_644,In_344,In_398);
or U645 (N_645,In_476,In_146);
nor U646 (N_646,In_115,In_251);
nor U647 (N_647,In_76,In_416);
and U648 (N_648,In_38,In_403);
and U649 (N_649,In_169,In_387);
nand U650 (N_650,In_492,In_382);
nand U651 (N_651,In_379,In_241);
and U652 (N_652,In_327,In_464);
or U653 (N_653,In_185,In_100);
nand U654 (N_654,In_488,In_193);
nor U655 (N_655,In_285,In_308);
nand U656 (N_656,In_66,In_246);
nor U657 (N_657,In_51,In_351);
nand U658 (N_658,In_146,In_233);
nor U659 (N_659,In_94,In_71);
and U660 (N_660,In_10,In_161);
nor U661 (N_661,In_258,In_496);
and U662 (N_662,In_217,In_436);
and U663 (N_663,In_421,In_307);
nor U664 (N_664,In_2,In_223);
nand U665 (N_665,In_237,In_402);
and U666 (N_666,In_57,In_146);
nor U667 (N_667,In_458,In_385);
and U668 (N_668,In_165,In_55);
nor U669 (N_669,In_292,In_312);
and U670 (N_670,In_252,In_51);
and U671 (N_671,In_61,In_185);
nand U672 (N_672,In_126,In_35);
nand U673 (N_673,In_164,In_260);
and U674 (N_674,In_262,In_487);
or U675 (N_675,In_451,In_357);
and U676 (N_676,In_40,In_444);
or U677 (N_677,In_343,In_183);
nor U678 (N_678,In_497,In_333);
nor U679 (N_679,In_171,In_276);
and U680 (N_680,In_463,In_414);
and U681 (N_681,In_261,In_469);
or U682 (N_682,In_490,In_67);
nor U683 (N_683,In_100,In_268);
nand U684 (N_684,In_386,In_384);
or U685 (N_685,In_128,In_422);
nor U686 (N_686,In_93,In_113);
nor U687 (N_687,In_303,In_468);
and U688 (N_688,In_225,In_301);
nor U689 (N_689,In_465,In_239);
and U690 (N_690,In_126,In_402);
nand U691 (N_691,In_308,In_41);
and U692 (N_692,In_140,In_169);
and U693 (N_693,In_337,In_446);
or U694 (N_694,In_444,In_277);
nor U695 (N_695,In_78,In_342);
or U696 (N_696,In_29,In_31);
nand U697 (N_697,In_231,In_92);
nor U698 (N_698,In_248,In_217);
and U699 (N_699,In_478,In_357);
nor U700 (N_700,In_331,In_210);
and U701 (N_701,In_301,In_281);
and U702 (N_702,In_20,In_91);
and U703 (N_703,In_22,In_39);
nand U704 (N_704,In_388,In_206);
and U705 (N_705,In_129,In_483);
nand U706 (N_706,In_287,In_372);
and U707 (N_707,In_323,In_429);
nand U708 (N_708,In_178,In_422);
nand U709 (N_709,In_216,In_229);
and U710 (N_710,In_123,In_121);
nor U711 (N_711,In_61,In_301);
or U712 (N_712,In_170,In_22);
nand U713 (N_713,In_305,In_84);
nand U714 (N_714,In_427,In_320);
nor U715 (N_715,In_308,In_401);
nor U716 (N_716,In_490,In_251);
and U717 (N_717,In_360,In_94);
or U718 (N_718,In_370,In_234);
or U719 (N_719,In_492,In_214);
or U720 (N_720,In_119,In_380);
and U721 (N_721,In_310,In_273);
or U722 (N_722,In_298,In_166);
and U723 (N_723,In_152,In_184);
nand U724 (N_724,In_366,In_3);
nor U725 (N_725,In_95,In_17);
nand U726 (N_726,In_224,In_27);
nor U727 (N_727,In_70,In_236);
nor U728 (N_728,In_128,In_480);
nor U729 (N_729,In_322,In_84);
nand U730 (N_730,In_368,In_184);
and U731 (N_731,In_358,In_162);
nor U732 (N_732,In_27,In_456);
or U733 (N_733,In_85,In_253);
xnor U734 (N_734,In_162,In_147);
and U735 (N_735,In_347,In_373);
nand U736 (N_736,In_477,In_355);
nand U737 (N_737,In_329,In_295);
nand U738 (N_738,In_236,In_404);
nand U739 (N_739,In_262,In_202);
or U740 (N_740,In_210,In_341);
nor U741 (N_741,In_202,In_272);
nand U742 (N_742,In_176,In_358);
and U743 (N_743,In_407,In_224);
or U744 (N_744,In_146,In_164);
or U745 (N_745,In_458,In_195);
nor U746 (N_746,In_67,In_120);
nor U747 (N_747,In_182,In_248);
nand U748 (N_748,In_21,In_428);
or U749 (N_749,In_104,In_178);
and U750 (N_750,N_39,N_662);
or U751 (N_751,N_627,N_618);
nor U752 (N_752,N_561,N_238);
or U753 (N_753,N_182,N_147);
nand U754 (N_754,N_52,N_732);
nand U755 (N_755,N_491,N_582);
and U756 (N_756,N_635,N_684);
and U757 (N_757,N_176,N_544);
nor U758 (N_758,N_432,N_434);
nor U759 (N_759,N_549,N_510);
nor U760 (N_760,N_509,N_112);
nand U761 (N_761,N_563,N_343);
or U762 (N_762,N_153,N_49);
and U763 (N_763,N_78,N_605);
or U764 (N_764,N_553,N_589);
nand U765 (N_765,N_195,N_728);
nor U766 (N_766,N_671,N_127);
nor U767 (N_767,N_460,N_314);
and U768 (N_768,N_722,N_174);
or U769 (N_769,N_739,N_641);
or U770 (N_770,N_375,N_276);
nand U771 (N_771,N_397,N_642);
nand U772 (N_772,N_436,N_424);
nand U773 (N_773,N_22,N_337);
and U774 (N_774,N_443,N_185);
and U775 (N_775,N_304,N_20);
or U776 (N_776,N_154,N_242);
nand U777 (N_777,N_298,N_344);
and U778 (N_778,N_137,N_483);
nand U779 (N_779,N_535,N_548);
and U780 (N_780,N_707,N_656);
or U781 (N_781,N_53,N_416);
nor U782 (N_782,N_437,N_226);
nor U783 (N_783,N_514,N_96);
and U784 (N_784,N_305,N_248);
nand U785 (N_785,N_19,N_172);
and U786 (N_786,N_178,N_719);
nor U787 (N_787,N_27,N_396);
or U788 (N_788,N_482,N_426);
nor U789 (N_789,N_80,N_152);
xor U790 (N_790,N_513,N_651);
nor U791 (N_791,N_478,N_158);
nor U792 (N_792,N_54,N_281);
nor U793 (N_793,N_83,N_290);
and U794 (N_794,N_6,N_274);
nand U795 (N_795,N_325,N_266);
nor U796 (N_796,N_107,N_547);
nor U797 (N_797,N_95,N_612);
nor U798 (N_798,N_398,N_620);
or U799 (N_799,N_645,N_327);
and U800 (N_800,N_23,N_367);
and U801 (N_801,N_488,N_494);
nand U802 (N_802,N_192,N_356);
or U803 (N_803,N_532,N_273);
and U804 (N_804,N_567,N_709);
or U805 (N_805,N_92,N_492);
nor U806 (N_806,N_686,N_476);
or U807 (N_807,N_316,N_411);
xnor U808 (N_808,N_134,N_36);
and U809 (N_809,N_198,N_431);
nor U810 (N_810,N_106,N_453);
or U811 (N_811,N_679,N_401);
nor U812 (N_812,N_529,N_150);
nand U813 (N_813,N_557,N_385);
and U814 (N_814,N_100,N_169);
and U815 (N_815,N_413,N_533);
nand U816 (N_816,N_278,N_70);
or U817 (N_817,N_120,N_148);
nor U818 (N_818,N_339,N_382);
nor U819 (N_819,N_211,N_604);
nand U820 (N_820,N_11,N_587);
nand U821 (N_821,N_420,N_371);
and U822 (N_822,N_88,N_733);
nor U823 (N_823,N_246,N_213);
or U824 (N_824,N_634,N_427);
and U825 (N_825,N_358,N_454);
nand U826 (N_826,N_9,N_183);
and U827 (N_827,N_217,N_540);
nor U828 (N_828,N_419,N_654);
or U829 (N_829,N_682,N_220);
or U830 (N_830,N_234,N_664);
nand U831 (N_831,N_577,N_690);
nor U832 (N_832,N_685,N_293);
and U833 (N_833,N_323,N_99);
and U834 (N_834,N_56,N_282);
and U835 (N_835,N_345,N_4);
or U836 (N_836,N_353,N_542);
and U837 (N_837,N_341,N_517);
and U838 (N_838,N_498,N_91);
nor U839 (N_839,N_463,N_44);
or U840 (N_840,N_222,N_531);
nor U841 (N_841,N_539,N_670);
nand U842 (N_842,N_638,N_128);
or U843 (N_843,N_108,N_394);
and U844 (N_844,N_379,N_186);
nor U845 (N_845,N_10,N_599);
nand U846 (N_846,N_607,N_487);
nor U847 (N_847,N_369,N_734);
nor U848 (N_848,N_110,N_0);
xor U849 (N_849,N_47,N_570);
and U850 (N_850,N_585,N_481);
and U851 (N_851,N_583,N_659);
nor U852 (N_852,N_425,N_97);
and U853 (N_853,N_562,N_746);
nor U854 (N_854,N_5,N_259);
and U855 (N_855,N_386,N_633);
nor U856 (N_856,N_285,N_418);
and U857 (N_857,N_208,N_409);
xnor U858 (N_858,N_523,N_399);
nand U859 (N_859,N_646,N_289);
nand U860 (N_860,N_748,N_28);
or U861 (N_861,N_519,N_569);
nor U862 (N_862,N_609,N_14);
or U863 (N_863,N_336,N_131);
nor U864 (N_864,N_180,N_271);
nand U865 (N_865,N_447,N_38);
nor U866 (N_866,N_42,N_522);
nor U867 (N_867,N_191,N_691);
nor U868 (N_868,N_361,N_441);
nand U869 (N_869,N_82,N_41);
nand U870 (N_870,N_233,N_267);
or U871 (N_871,N_171,N_546);
and U872 (N_872,N_366,N_486);
and U873 (N_873,N_235,N_156);
and U874 (N_874,N_132,N_650);
and U875 (N_875,N_317,N_340);
nor U876 (N_876,N_380,N_319);
and U877 (N_877,N_559,N_669);
and U878 (N_878,N_444,N_588);
or U879 (N_879,N_383,N_296);
or U880 (N_880,N_727,N_695);
or U881 (N_881,N_493,N_743);
xor U882 (N_882,N_741,N_268);
or U883 (N_883,N_680,N_520);
or U884 (N_884,N_270,N_469);
and U885 (N_885,N_138,N_628);
nand U886 (N_886,N_151,N_372);
nand U887 (N_887,N_123,N_33);
nor U888 (N_888,N_142,N_126);
nand U889 (N_889,N_395,N_239);
nand U890 (N_890,N_665,N_558);
nor U891 (N_891,N_455,N_376);
or U892 (N_892,N_30,N_76);
and U893 (N_893,N_105,N_160);
nand U894 (N_894,N_101,N_747);
nand U895 (N_895,N_331,N_631);
nand U896 (N_896,N_359,N_363);
or U897 (N_897,N_593,N_720);
nor U898 (N_898,N_224,N_61);
or U899 (N_899,N_193,N_368);
nand U900 (N_900,N_135,N_145);
and U901 (N_901,N_201,N_745);
nand U902 (N_902,N_674,N_288);
nand U903 (N_903,N_300,N_284);
nor U904 (N_904,N_360,N_161);
nand U905 (N_905,N_637,N_269);
and U906 (N_906,N_111,N_349);
nand U907 (N_907,N_272,N_21);
nand U908 (N_908,N_364,N_79);
nor U909 (N_909,N_303,N_414);
and U910 (N_910,N_449,N_576);
nor U911 (N_911,N_320,N_452);
nand U912 (N_912,N_484,N_417);
nand U913 (N_913,N_742,N_250);
nor U914 (N_914,N_50,N_438);
nor U915 (N_915,N_173,N_229);
or U916 (N_916,N_716,N_537);
and U917 (N_917,N_479,N_381);
and U918 (N_918,N_313,N_700);
and U919 (N_919,N_245,N_545);
nor U920 (N_920,N_254,N_62);
nor U921 (N_921,N_592,N_579);
and U922 (N_922,N_660,N_465);
nand U923 (N_923,N_29,N_37);
or U924 (N_924,N_572,N_321);
nor U925 (N_925,N_672,N_165);
or U926 (N_926,N_698,N_456);
nor U927 (N_927,N_534,N_626);
nor U928 (N_928,N_617,N_109);
or U929 (N_929,N_1,N_603);
nor U930 (N_930,N_194,N_699);
nand U931 (N_931,N_393,N_705);
or U932 (N_932,N_125,N_89);
and U933 (N_933,N_640,N_737);
nand U934 (N_934,N_428,N_505);
nor U935 (N_935,N_715,N_77);
or U936 (N_936,N_666,N_429);
nand U937 (N_937,N_616,N_692);
nor U938 (N_938,N_600,N_578);
or U939 (N_939,N_595,N_90);
nor U940 (N_940,N_636,N_73);
or U941 (N_941,N_661,N_710);
nand U942 (N_942,N_2,N_253);
nor U943 (N_943,N_69,N_580);
nand U944 (N_944,N_139,N_687);
nand U945 (N_945,N_104,N_75);
nand U946 (N_946,N_179,N_644);
nor U947 (N_947,N_346,N_240);
xnor U948 (N_948,N_678,N_223);
nor U949 (N_949,N_348,N_565);
nand U950 (N_950,N_655,N_312);
or U951 (N_951,N_58,N_611);
nor U952 (N_952,N_574,N_721);
and U953 (N_953,N_458,N_474);
nand U954 (N_954,N_730,N_265);
nor U955 (N_955,N_442,N_264);
nor U956 (N_956,N_718,N_495);
or U957 (N_957,N_744,N_68);
nand U958 (N_958,N_287,N_421);
and U959 (N_959,N_738,N_415);
nor U960 (N_960,N_657,N_713);
and U961 (N_961,N_663,N_332);
or U962 (N_962,N_330,N_647);
nand U963 (N_963,N_515,N_103);
nand U964 (N_964,N_236,N_113);
or U965 (N_965,N_377,N_351);
and U966 (N_966,N_681,N_717);
xor U967 (N_967,N_508,N_228);
or U968 (N_968,N_334,N_207);
nor U969 (N_969,N_613,N_129);
or U970 (N_970,N_378,N_181);
and U971 (N_971,N_596,N_85);
and U972 (N_972,N_65,N_497);
nor U973 (N_973,N_189,N_615);
nand U974 (N_974,N_60,N_697);
and U975 (N_975,N_219,N_167);
nand U976 (N_976,N_18,N_114);
and U977 (N_977,N_143,N_555);
xnor U978 (N_978,N_499,N_704);
and U979 (N_979,N_188,N_315);
or U980 (N_980,N_598,N_133);
nor U981 (N_981,N_93,N_237);
nor U982 (N_982,N_244,N_435);
and U983 (N_983,N_170,N_408);
and U984 (N_984,N_324,N_225);
and U985 (N_985,N_308,N_502);
nand U986 (N_986,N_528,N_608);
nor U987 (N_987,N_322,N_594);
nor U988 (N_988,N_196,N_501);
or U989 (N_989,N_525,N_136);
and U990 (N_990,N_157,N_606);
nand U991 (N_991,N_388,N_590);
or U992 (N_992,N_507,N_51);
nor U993 (N_993,N_283,N_202);
nand U994 (N_994,N_602,N_389);
and U995 (N_995,N_218,N_630);
or U996 (N_996,N_500,N_214);
nand U997 (N_997,N_632,N_159);
nand U998 (N_998,N_402,N_601);
and U999 (N_999,N_735,N_280);
xor U1000 (N_1000,N_141,N_541);
or U1001 (N_1001,N_275,N_122);
nand U1002 (N_1002,N_67,N_140);
or U1003 (N_1003,N_168,N_496);
and U1004 (N_1004,N_243,N_683);
nand U1005 (N_1005,N_673,N_467);
and U1006 (N_1006,N_445,N_177);
or U1007 (N_1007,N_554,N_63);
or U1008 (N_1008,N_350,N_450);
nor U1009 (N_1009,N_726,N_354);
and U1010 (N_1010,N_318,N_57);
and U1011 (N_1011,N_335,N_464);
nand U1012 (N_1012,N_530,N_489);
or U1013 (N_1013,N_40,N_649);
and U1014 (N_1014,N_675,N_301);
and U1015 (N_1015,N_209,N_3);
nand U1016 (N_1016,N_306,N_204);
nand U1017 (N_1017,N_357,N_130);
and U1018 (N_1018,N_667,N_564);
nor U1019 (N_1019,N_475,N_392);
or U1020 (N_1020,N_461,N_466);
nor U1021 (N_1021,N_203,N_190);
nor U1022 (N_1022,N_175,N_736);
nor U1023 (N_1023,N_72,N_597);
or U1024 (N_1024,N_121,N_652);
and U1025 (N_1025,N_556,N_560);
nand U1026 (N_1026,N_146,N_355);
nor U1027 (N_1027,N_689,N_295);
or U1028 (N_1028,N_403,N_573);
or U1029 (N_1029,N_205,N_749);
or U1030 (N_1030,N_446,N_310);
nand U1031 (N_1031,N_571,N_568);
or U1032 (N_1032,N_291,N_702);
and U1033 (N_1033,N_149,N_118);
nand U1034 (N_1034,N_676,N_696);
nor U1035 (N_1035,N_365,N_439);
or U1036 (N_1036,N_212,N_261);
or U1037 (N_1037,N_391,N_333);
nor U1038 (N_1038,N_410,N_299);
and U1039 (N_1039,N_277,N_326);
nand U1040 (N_1040,N_8,N_119);
or U1041 (N_1041,N_423,N_586);
or U1042 (N_1042,N_538,N_462);
nand U1043 (N_1043,N_440,N_307);
nor U1044 (N_1044,N_66,N_162);
or U1045 (N_1045,N_485,N_309);
nor U1046 (N_1046,N_512,N_693);
and U1047 (N_1047,N_373,N_405);
nor U1048 (N_1048,N_215,N_712);
and U1049 (N_1049,N_490,N_688);
nor U1050 (N_1050,N_459,N_35);
nand U1051 (N_1051,N_164,N_472);
and U1052 (N_1052,N_591,N_16);
nor U1053 (N_1053,N_197,N_86);
and U1054 (N_1054,N_200,N_115);
nor U1055 (N_1055,N_477,N_729);
nor U1056 (N_1056,N_619,N_623);
or U1057 (N_1057,N_703,N_370);
or U1058 (N_1058,N_84,N_536);
nor U1059 (N_1059,N_94,N_566);
nor U1060 (N_1060,N_45,N_668);
nor U1061 (N_1061,N_286,N_59);
and U1062 (N_1062,N_422,N_524);
and U1063 (N_1063,N_550,N_260);
nand U1064 (N_1064,N_7,N_247);
and U1065 (N_1065,N_677,N_714);
or U1066 (N_1066,N_17,N_48);
nor U1067 (N_1067,N_352,N_230);
nor U1068 (N_1068,N_653,N_621);
or U1069 (N_1069,N_639,N_31);
nor U1070 (N_1070,N_251,N_311);
or U1071 (N_1071,N_43,N_55);
or U1072 (N_1072,N_390,N_13);
or U1073 (N_1073,N_329,N_255);
or U1074 (N_1074,N_46,N_98);
and U1075 (N_1075,N_610,N_504);
nand U1076 (N_1076,N_694,N_328);
and U1077 (N_1077,N_503,N_116);
nand U1078 (N_1078,N_227,N_468);
or U1079 (N_1079,N_701,N_231);
or U1080 (N_1080,N_124,N_648);
and U1081 (N_1081,N_480,N_643);
nor U1082 (N_1082,N_473,N_731);
nor U1083 (N_1083,N_406,N_725);
and U1084 (N_1084,N_279,N_506);
xor U1085 (N_1085,N_412,N_338);
or U1086 (N_1086,N_518,N_144);
and U1087 (N_1087,N_257,N_81);
or U1088 (N_1088,N_155,N_24);
nor U1089 (N_1089,N_581,N_221);
and U1090 (N_1090,N_15,N_448);
nor U1091 (N_1091,N_543,N_102);
nand U1092 (N_1092,N_71,N_384);
nor U1093 (N_1093,N_25,N_430);
nor U1094 (N_1094,N_262,N_629);
nand U1095 (N_1095,N_166,N_216);
nand U1096 (N_1096,N_32,N_26);
and U1097 (N_1097,N_740,N_187);
or U1098 (N_1098,N_551,N_249);
nand U1099 (N_1099,N_374,N_521);
and U1100 (N_1100,N_347,N_342);
nor U1101 (N_1101,N_451,N_294);
nand U1102 (N_1102,N_210,N_470);
and U1103 (N_1103,N_404,N_400);
and U1104 (N_1104,N_64,N_575);
nand U1105 (N_1105,N_407,N_511);
nor U1106 (N_1106,N_206,N_256);
nor U1107 (N_1107,N_527,N_232);
and U1108 (N_1108,N_387,N_163);
or U1109 (N_1109,N_552,N_34);
or U1110 (N_1110,N_706,N_584);
and U1111 (N_1111,N_457,N_658);
or U1112 (N_1112,N_199,N_12);
and U1113 (N_1113,N_723,N_263);
nand U1114 (N_1114,N_622,N_708);
nand U1115 (N_1115,N_516,N_292);
nor U1116 (N_1116,N_117,N_302);
and U1117 (N_1117,N_87,N_252);
nand U1118 (N_1118,N_74,N_526);
or U1119 (N_1119,N_433,N_184);
and U1120 (N_1120,N_625,N_241);
nand U1121 (N_1121,N_614,N_471);
and U1122 (N_1122,N_362,N_297);
or U1123 (N_1123,N_624,N_711);
and U1124 (N_1124,N_258,N_724);
nand U1125 (N_1125,N_272,N_114);
nor U1126 (N_1126,N_533,N_395);
or U1127 (N_1127,N_74,N_124);
nor U1128 (N_1128,N_75,N_151);
or U1129 (N_1129,N_215,N_586);
and U1130 (N_1130,N_287,N_447);
nor U1131 (N_1131,N_555,N_612);
or U1132 (N_1132,N_687,N_434);
nor U1133 (N_1133,N_462,N_413);
or U1134 (N_1134,N_186,N_394);
nor U1135 (N_1135,N_725,N_316);
nand U1136 (N_1136,N_331,N_591);
or U1137 (N_1137,N_22,N_600);
and U1138 (N_1138,N_728,N_546);
or U1139 (N_1139,N_722,N_518);
or U1140 (N_1140,N_135,N_356);
nor U1141 (N_1141,N_69,N_377);
or U1142 (N_1142,N_442,N_63);
xnor U1143 (N_1143,N_181,N_525);
nand U1144 (N_1144,N_401,N_744);
nor U1145 (N_1145,N_366,N_545);
nor U1146 (N_1146,N_175,N_454);
nand U1147 (N_1147,N_136,N_53);
and U1148 (N_1148,N_365,N_140);
nand U1149 (N_1149,N_131,N_37);
and U1150 (N_1150,N_480,N_659);
nor U1151 (N_1151,N_278,N_436);
or U1152 (N_1152,N_187,N_597);
nor U1153 (N_1153,N_423,N_702);
nor U1154 (N_1154,N_247,N_544);
and U1155 (N_1155,N_176,N_462);
and U1156 (N_1156,N_380,N_102);
nor U1157 (N_1157,N_602,N_378);
and U1158 (N_1158,N_317,N_556);
nand U1159 (N_1159,N_427,N_283);
or U1160 (N_1160,N_157,N_635);
nand U1161 (N_1161,N_346,N_587);
nor U1162 (N_1162,N_599,N_612);
and U1163 (N_1163,N_511,N_187);
or U1164 (N_1164,N_744,N_466);
nand U1165 (N_1165,N_374,N_458);
nand U1166 (N_1166,N_290,N_275);
nand U1167 (N_1167,N_600,N_45);
nor U1168 (N_1168,N_749,N_543);
or U1169 (N_1169,N_86,N_408);
nand U1170 (N_1170,N_163,N_27);
xor U1171 (N_1171,N_546,N_621);
xnor U1172 (N_1172,N_76,N_747);
or U1173 (N_1173,N_553,N_71);
or U1174 (N_1174,N_159,N_343);
and U1175 (N_1175,N_361,N_219);
nor U1176 (N_1176,N_82,N_79);
and U1177 (N_1177,N_646,N_598);
and U1178 (N_1178,N_696,N_691);
nand U1179 (N_1179,N_689,N_38);
nand U1180 (N_1180,N_226,N_690);
or U1181 (N_1181,N_394,N_202);
nor U1182 (N_1182,N_693,N_284);
or U1183 (N_1183,N_64,N_282);
and U1184 (N_1184,N_128,N_167);
or U1185 (N_1185,N_190,N_306);
or U1186 (N_1186,N_304,N_348);
nand U1187 (N_1187,N_273,N_594);
and U1188 (N_1188,N_273,N_521);
and U1189 (N_1189,N_124,N_77);
nor U1190 (N_1190,N_556,N_32);
nand U1191 (N_1191,N_449,N_65);
and U1192 (N_1192,N_451,N_14);
and U1193 (N_1193,N_128,N_6);
or U1194 (N_1194,N_494,N_192);
nor U1195 (N_1195,N_370,N_456);
and U1196 (N_1196,N_210,N_277);
and U1197 (N_1197,N_559,N_111);
nand U1198 (N_1198,N_205,N_75);
nand U1199 (N_1199,N_249,N_584);
or U1200 (N_1200,N_213,N_162);
nand U1201 (N_1201,N_343,N_699);
and U1202 (N_1202,N_296,N_495);
or U1203 (N_1203,N_240,N_43);
and U1204 (N_1204,N_636,N_633);
nand U1205 (N_1205,N_3,N_525);
or U1206 (N_1206,N_147,N_330);
nand U1207 (N_1207,N_443,N_679);
and U1208 (N_1208,N_740,N_424);
nor U1209 (N_1209,N_186,N_326);
nand U1210 (N_1210,N_260,N_85);
nor U1211 (N_1211,N_390,N_511);
nor U1212 (N_1212,N_448,N_192);
nor U1213 (N_1213,N_448,N_539);
nand U1214 (N_1214,N_422,N_260);
or U1215 (N_1215,N_212,N_234);
or U1216 (N_1216,N_603,N_635);
nor U1217 (N_1217,N_345,N_405);
and U1218 (N_1218,N_502,N_743);
or U1219 (N_1219,N_746,N_136);
or U1220 (N_1220,N_735,N_676);
nand U1221 (N_1221,N_666,N_163);
nor U1222 (N_1222,N_428,N_627);
and U1223 (N_1223,N_283,N_75);
and U1224 (N_1224,N_271,N_734);
and U1225 (N_1225,N_210,N_160);
or U1226 (N_1226,N_64,N_19);
nor U1227 (N_1227,N_318,N_17);
and U1228 (N_1228,N_692,N_292);
or U1229 (N_1229,N_70,N_156);
xor U1230 (N_1230,N_223,N_457);
and U1231 (N_1231,N_237,N_150);
or U1232 (N_1232,N_468,N_413);
and U1233 (N_1233,N_627,N_743);
or U1234 (N_1234,N_387,N_685);
nor U1235 (N_1235,N_298,N_635);
nor U1236 (N_1236,N_408,N_99);
nor U1237 (N_1237,N_650,N_491);
or U1238 (N_1238,N_277,N_725);
xor U1239 (N_1239,N_448,N_281);
or U1240 (N_1240,N_51,N_457);
nand U1241 (N_1241,N_79,N_438);
or U1242 (N_1242,N_158,N_658);
nand U1243 (N_1243,N_185,N_209);
nand U1244 (N_1244,N_241,N_128);
and U1245 (N_1245,N_676,N_367);
or U1246 (N_1246,N_93,N_599);
nor U1247 (N_1247,N_178,N_469);
or U1248 (N_1248,N_99,N_662);
nor U1249 (N_1249,N_127,N_644);
nor U1250 (N_1250,N_136,N_82);
and U1251 (N_1251,N_60,N_695);
nor U1252 (N_1252,N_20,N_31);
or U1253 (N_1253,N_432,N_211);
nor U1254 (N_1254,N_167,N_338);
and U1255 (N_1255,N_111,N_155);
nor U1256 (N_1256,N_639,N_682);
or U1257 (N_1257,N_389,N_446);
and U1258 (N_1258,N_95,N_343);
nand U1259 (N_1259,N_78,N_292);
nand U1260 (N_1260,N_403,N_267);
or U1261 (N_1261,N_695,N_432);
or U1262 (N_1262,N_132,N_260);
nand U1263 (N_1263,N_167,N_608);
nor U1264 (N_1264,N_673,N_695);
or U1265 (N_1265,N_205,N_644);
or U1266 (N_1266,N_100,N_439);
nand U1267 (N_1267,N_726,N_578);
nand U1268 (N_1268,N_466,N_54);
and U1269 (N_1269,N_46,N_433);
or U1270 (N_1270,N_51,N_714);
or U1271 (N_1271,N_488,N_708);
or U1272 (N_1272,N_359,N_550);
nor U1273 (N_1273,N_298,N_418);
nand U1274 (N_1274,N_683,N_513);
and U1275 (N_1275,N_561,N_565);
or U1276 (N_1276,N_182,N_305);
nand U1277 (N_1277,N_412,N_517);
or U1278 (N_1278,N_280,N_84);
nand U1279 (N_1279,N_483,N_720);
nor U1280 (N_1280,N_570,N_353);
or U1281 (N_1281,N_508,N_136);
nand U1282 (N_1282,N_123,N_703);
or U1283 (N_1283,N_0,N_321);
or U1284 (N_1284,N_409,N_636);
nor U1285 (N_1285,N_438,N_711);
and U1286 (N_1286,N_724,N_497);
nand U1287 (N_1287,N_134,N_544);
nand U1288 (N_1288,N_276,N_690);
nor U1289 (N_1289,N_749,N_610);
or U1290 (N_1290,N_135,N_150);
or U1291 (N_1291,N_380,N_647);
and U1292 (N_1292,N_187,N_690);
or U1293 (N_1293,N_681,N_159);
and U1294 (N_1294,N_563,N_67);
or U1295 (N_1295,N_658,N_662);
nor U1296 (N_1296,N_737,N_721);
or U1297 (N_1297,N_601,N_26);
nor U1298 (N_1298,N_498,N_75);
nor U1299 (N_1299,N_342,N_156);
and U1300 (N_1300,N_630,N_14);
and U1301 (N_1301,N_219,N_289);
or U1302 (N_1302,N_407,N_551);
nand U1303 (N_1303,N_23,N_429);
nor U1304 (N_1304,N_25,N_238);
nand U1305 (N_1305,N_180,N_702);
nor U1306 (N_1306,N_746,N_450);
or U1307 (N_1307,N_662,N_152);
xnor U1308 (N_1308,N_266,N_46);
and U1309 (N_1309,N_356,N_545);
nor U1310 (N_1310,N_624,N_207);
and U1311 (N_1311,N_614,N_546);
or U1312 (N_1312,N_738,N_27);
nor U1313 (N_1313,N_552,N_178);
and U1314 (N_1314,N_19,N_505);
nor U1315 (N_1315,N_273,N_194);
and U1316 (N_1316,N_454,N_661);
nor U1317 (N_1317,N_150,N_615);
nand U1318 (N_1318,N_570,N_304);
xor U1319 (N_1319,N_642,N_650);
or U1320 (N_1320,N_51,N_561);
nand U1321 (N_1321,N_354,N_35);
or U1322 (N_1322,N_263,N_32);
nor U1323 (N_1323,N_344,N_50);
nand U1324 (N_1324,N_738,N_227);
nand U1325 (N_1325,N_638,N_549);
or U1326 (N_1326,N_643,N_728);
nor U1327 (N_1327,N_287,N_729);
or U1328 (N_1328,N_562,N_327);
or U1329 (N_1329,N_323,N_390);
or U1330 (N_1330,N_724,N_259);
nor U1331 (N_1331,N_243,N_742);
nor U1332 (N_1332,N_232,N_403);
nor U1333 (N_1333,N_491,N_593);
xor U1334 (N_1334,N_661,N_146);
nor U1335 (N_1335,N_37,N_616);
nor U1336 (N_1336,N_559,N_100);
nor U1337 (N_1337,N_224,N_618);
or U1338 (N_1338,N_9,N_626);
or U1339 (N_1339,N_286,N_591);
nand U1340 (N_1340,N_222,N_450);
nor U1341 (N_1341,N_327,N_598);
nand U1342 (N_1342,N_357,N_464);
nand U1343 (N_1343,N_387,N_648);
or U1344 (N_1344,N_34,N_52);
nor U1345 (N_1345,N_312,N_375);
and U1346 (N_1346,N_559,N_91);
and U1347 (N_1347,N_742,N_687);
nor U1348 (N_1348,N_123,N_285);
nand U1349 (N_1349,N_643,N_695);
and U1350 (N_1350,N_251,N_443);
or U1351 (N_1351,N_312,N_498);
and U1352 (N_1352,N_54,N_120);
or U1353 (N_1353,N_686,N_582);
and U1354 (N_1354,N_693,N_443);
xor U1355 (N_1355,N_181,N_439);
nand U1356 (N_1356,N_643,N_507);
or U1357 (N_1357,N_323,N_668);
or U1358 (N_1358,N_345,N_404);
or U1359 (N_1359,N_402,N_103);
or U1360 (N_1360,N_663,N_46);
and U1361 (N_1361,N_643,N_404);
xnor U1362 (N_1362,N_627,N_47);
and U1363 (N_1363,N_433,N_140);
nand U1364 (N_1364,N_542,N_432);
nor U1365 (N_1365,N_545,N_514);
nand U1366 (N_1366,N_250,N_286);
nand U1367 (N_1367,N_21,N_197);
nand U1368 (N_1368,N_684,N_71);
and U1369 (N_1369,N_193,N_227);
nand U1370 (N_1370,N_198,N_2);
or U1371 (N_1371,N_479,N_505);
xnor U1372 (N_1372,N_508,N_315);
xnor U1373 (N_1373,N_364,N_396);
and U1374 (N_1374,N_424,N_104);
nor U1375 (N_1375,N_294,N_334);
xor U1376 (N_1376,N_274,N_145);
nand U1377 (N_1377,N_19,N_518);
nor U1378 (N_1378,N_530,N_251);
and U1379 (N_1379,N_325,N_259);
nor U1380 (N_1380,N_391,N_603);
nor U1381 (N_1381,N_545,N_177);
nor U1382 (N_1382,N_472,N_231);
nand U1383 (N_1383,N_631,N_529);
and U1384 (N_1384,N_76,N_413);
nand U1385 (N_1385,N_413,N_313);
nand U1386 (N_1386,N_471,N_17);
or U1387 (N_1387,N_377,N_312);
nor U1388 (N_1388,N_597,N_533);
and U1389 (N_1389,N_101,N_581);
nand U1390 (N_1390,N_710,N_85);
nor U1391 (N_1391,N_488,N_109);
and U1392 (N_1392,N_707,N_373);
or U1393 (N_1393,N_189,N_738);
nand U1394 (N_1394,N_234,N_326);
nor U1395 (N_1395,N_573,N_197);
nor U1396 (N_1396,N_521,N_114);
xnor U1397 (N_1397,N_215,N_11);
or U1398 (N_1398,N_379,N_317);
nor U1399 (N_1399,N_391,N_178);
nor U1400 (N_1400,N_189,N_72);
nor U1401 (N_1401,N_583,N_597);
and U1402 (N_1402,N_181,N_402);
and U1403 (N_1403,N_69,N_375);
nor U1404 (N_1404,N_442,N_712);
nand U1405 (N_1405,N_662,N_668);
nor U1406 (N_1406,N_11,N_742);
nor U1407 (N_1407,N_668,N_631);
nor U1408 (N_1408,N_229,N_612);
nor U1409 (N_1409,N_607,N_525);
nand U1410 (N_1410,N_665,N_492);
nor U1411 (N_1411,N_402,N_153);
or U1412 (N_1412,N_709,N_342);
or U1413 (N_1413,N_119,N_412);
and U1414 (N_1414,N_569,N_51);
nor U1415 (N_1415,N_323,N_536);
or U1416 (N_1416,N_678,N_234);
or U1417 (N_1417,N_372,N_473);
nor U1418 (N_1418,N_333,N_524);
nand U1419 (N_1419,N_694,N_32);
or U1420 (N_1420,N_259,N_109);
or U1421 (N_1421,N_53,N_402);
or U1422 (N_1422,N_56,N_727);
and U1423 (N_1423,N_40,N_91);
or U1424 (N_1424,N_0,N_120);
or U1425 (N_1425,N_594,N_651);
nor U1426 (N_1426,N_649,N_373);
nand U1427 (N_1427,N_536,N_338);
nand U1428 (N_1428,N_272,N_733);
nor U1429 (N_1429,N_393,N_360);
or U1430 (N_1430,N_360,N_83);
and U1431 (N_1431,N_254,N_503);
and U1432 (N_1432,N_165,N_285);
or U1433 (N_1433,N_619,N_466);
nand U1434 (N_1434,N_658,N_629);
nor U1435 (N_1435,N_530,N_574);
or U1436 (N_1436,N_90,N_563);
nor U1437 (N_1437,N_458,N_312);
and U1438 (N_1438,N_68,N_145);
nor U1439 (N_1439,N_303,N_508);
and U1440 (N_1440,N_70,N_259);
or U1441 (N_1441,N_156,N_721);
and U1442 (N_1442,N_637,N_645);
nand U1443 (N_1443,N_495,N_356);
and U1444 (N_1444,N_688,N_371);
and U1445 (N_1445,N_233,N_701);
nand U1446 (N_1446,N_161,N_501);
nor U1447 (N_1447,N_551,N_605);
and U1448 (N_1448,N_134,N_647);
nand U1449 (N_1449,N_101,N_240);
and U1450 (N_1450,N_238,N_292);
nor U1451 (N_1451,N_76,N_633);
xnor U1452 (N_1452,N_584,N_103);
nor U1453 (N_1453,N_574,N_297);
nand U1454 (N_1454,N_131,N_524);
nand U1455 (N_1455,N_507,N_343);
or U1456 (N_1456,N_245,N_175);
and U1457 (N_1457,N_292,N_188);
nand U1458 (N_1458,N_660,N_116);
or U1459 (N_1459,N_704,N_139);
nand U1460 (N_1460,N_268,N_182);
nor U1461 (N_1461,N_445,N_588);
or U1462 (N_1462,N_502,N_241);
nor U1463 (N_1463,N_699,N_57);
nor U1464 (N_1464,N_173,N_523);
and U1465 (N_1465,N_627,N_714);
and U1466 (N_1466,N_172,N_287);
xnor U1467 (N_1467,N_346,N_134);
or U1468 (N_1468,N_197,N_719);
and U1469 (N_1469,N_344,N_653);
nor U1470 (N_1470,N_552,N_714);
nor U1471 (N_1471,N_261,N_456);
nor U1472 (N_1472,N_70,N_379);
nand U1473 (N_1473,N_146,N_204);
nand U1474 (N_1474,N_615,N_423);
nor U1475 (N_1475,N_15,N_714);
or U1476 (N_1476,N_587,N_233);
nor U1477 (N_1477,N_6,N_617);
nand U1478 (N_1478,N_420,N_136);
nor U1479 (N_1479,N_654,N_227);
nor U1480 (N_1480,N_210,N_594);
nor U1481 (N_1481,N_547,N_427);
nand U1482 (N_1482,N_93,N_566);
nor U1483 (N_1483,N_749,N_495);
and U1484 (N_1484,N_536,N_114);
or U1485 (N_1485,N_689,N_263);
nand U1486 (N_1486,N_542,N_517);
and U1487 (N_1487,N_667,N_336);
or U1488 (N_1488,N_29,N_358);
nor U1489 (N_1489,N_458,N_395);
nand U1490 (N_1490,N_370,N_515);
nand U1491 (N_1491,N_360,N_515);
and U1492 (N_1492,N_371,N_640);
and U1493 (N_1493,N_130,N_267);
or U1494 (N_1494,N_175,N_677);
and U1495 (N_1495,N_627,N_626);
nand U1496 (N_1496,N_446,N_480);
nand U1497 (N_1497,N_483,N_593);
and U1498 (N_1498,N_165,N_343);
nand U1499 (N_1499,N_409,N_432);
and U1500 (N_1500,N_1268,N_1002);
nand U1501 (N_1501,N_1165,N_1108);
nand U1502 (N_1502,N_1432,N_785);
and U1503 (N_1503,N_824,N_1475);
nor U1504 (N_1504,N_1219,N_873);
and U1505 (N_1505,N_1383,N_890);
or U1506 (N_1506,N_1469,N_1244);
or U1507 (N_1507,N_1048,N_1222);
or U1508 (N_1508,N_1168,N_1438);
xor U1509 (N_1509,N_1100,N_1425);
or U1510 (N_1510,N_1443,N_1128);
nor U1511 (N_1511,N_972,N_1005);
nor U1512 (N_1512,N_1253,N_1429);
nor U1513 (N_1513,N_885,N_896);
and U1514 (N_1514,N_1391,N_1186);
and U1515 (N_1515,N_1476,N_1171);
and U1516 (N_1516,N_1293,N_1091);
nand U1517 (N_1517,N_1490,N_905);
nor U1518 (N_1518,N_1373,N_1412);
nand U1519 (N_1519,N_1367,N_1081);
nand U1520 (N_1520,N_900,N_1382);
nand U1521 (N_1521,N_986,N_1348);
or U1522 (N_1522,N_848,N_1023);
or U1523 (N_1523,N_1146,N_1021);
nand U1524 (N_1524,N_959,N_1489);
and U1525 (N_1525,N_1182,N_1296);
nand U1526 (N_1526,N_1378,N_862);
or U1527 (N_1527,N_1390,N_792);
nor U1528 (N_1528,N_1319,N_1095);
nor U1529 (N_1529,N_1071,N_876);
and U1530 (N_1530,N_1086,N_1465);
or U1531 (N_1531,N_978,N_1356);
and U1532 (N_1532,N_878,N_807);
nor U1533 (N_1533,N_1089,N_852);
and U1534 (N_1534,N_1326,N_1250);
and U1535 (N_1535,N_1427,N_835);
or U1536 (N_1536,N_1082,N_1450);
nand U1537 (N_1537,N_1050,N_1470);
and U1538 (N_1538,N_818,N_965);
nor U1539 (N_1539,N_899,N_881);
and U1540 (N_1540,N_1175,N_806);
and U1541 (N_1541,N_837,N_1347);
xnor U1542 (N_1542,N_984,N_1158);
and U1543 (N_1543,N_1352,N_1288);
or U1544 (N_1544,N_1085,N_1061);
nor U1545 (N_1545,N_934,N_754);
nor U1546 (N_1546,N_1011,N_1026);
and U1547 (N_1547,N_1112,N_1079);
or U1548 (N_1548,N_1374,N_802);
or U1549 (N_1549,N_1402,N_801);
or U1550 (N_1550,N_774,N_1052);
or U1551 (N_1551,N_751,N_909);
or U1552 (N_1552,N_1466,N_907);
and U1553 (N_1553,N_887,N_1015);
nand U1554 (N_1554,N_863,N_1130);
and U1555 (N_1555,N_990,N_1185);
nor U1556 (N_1556,N_1178,N_1366);
and U1557 (N_1557,N_1148,N_1484);
and U1558 (N_1558,N_1265,N_1109);
and U1559 (N_1559,N_964,N_1313);
nor U1560 (N_1560,N_1216,N_1074);
or U1561 (N_1561,N_969,N_858);
nand U1562 (N_1562,N_1462,N_1436);
and U1563 (N_1563,N_1249,N_836);
and U1564 (N_1564,N_1012,N_825);
or U1565 (N_1565,N_1246,N_1325);
and U1566 (N_1566,N_1426,N_1138);
nor U1567 (N_1567,N_834,N_798);
or U1568 (N_1568,N_989,N_1446);
nor U1569 (N_1569,N_830,N_952);
nor U1570 (N_1570,N_1123,N_1422);
nand U1571 (N_1571,N_1388,N_771);
nand U1572 (N_1572,N_1247,N_1387);
nor U1573 (N_1573,N_924,N_985);
nand U1574 (N_1574,N_1126,N_869);
nand U1575 (N_1575,N_1414,N_1341);
nor U1576 (N_1576,N_1077,N_1202);
and U1577 (N_1577,N_979,N_1097);
nand U1578 (N_1578,N_810,N_1275);
and U1579 (N_1579,N_875,N_1206);
nand U1580 (N_1580,N_1121,N_1283);
and U1581 (N_1581,N_1457,N_1420);
or U1582 (N_1582,N_921,N_947);
and U1583 (N_1583,N_1252,N_1063);
and U1584 (N_1584,N_1447,N_1331);
or U1585 (N_1585,N_1302,N_1029);
nor U1586 (N_1586,N_943,N_1188);
and U1587 (N_1587,N_1020,N_1358);
nor U1588 (N_1588,N_987,N_1167);
nor U1589 (N_1589,N_1025,N_874);
nand U1590 (N_1590,N_1393,N_1073);
nand U1591 (N_1591,N_973,N_1140);
or U1592 (N_1592,N_1280,N_1497);
nand U1593 (N_1593,N_1278,N_1363);
nand U1594 (N_1594,N_1449,N_1212);
nand U1595 (N_1595,N_1267,N_930);
nand U1596 (N_1596,N_1224,N_1306);
and U1597 (N_1597,N_1122,N_1421);
or U1598 (N_1598,N_829,N_1181);
or U1599 (N_1599,N_962,N_1337);
and U1600 (N_1600,N_805,N_1468);
nor U1601 (N_1601,N_941,N_1027);
nand U1602 (N_1602,N_877,N_776);
or U1603 (N_1603,N_1105,N_1481);
nor U1604 (N_1604,N_1389,N_1474);
and U1605 (N_1605,N_1384,N_980);
or U1606 (N_1606,N_1416,N_1149);
and U1607 (N_1607,N_1004,N_1361);
nor U1608 (N_1608,N_1415,N_1180);
nor U1609 (N_1609,N_1159,N_1368);
or U1610 (N_1610,N_820,N_819);
nand U1611 (N_1611,N_1187,N_1134);
or U1612 (N_1612,N_1069,N_1444);
nand U1613 (N_1613,N_1006,N_1228);
or U1614 (N_1614,N_1194,N_1164);
xor U1615 (N_1615,N_1260,N_920);
and U1616 (N_1616,N_767,N_1279);
or U1617 (N_1617,N_1254,N_859);
nor U1618 (N_1618,N_1351,N_1092);
nor U1619 (N_1619,N_1197,N_1036);
nor U1620 (N_1620,N_1031,N_914);
and U1621 (N_1621,N_762,N_1084);
nand U1622 (N_1622,N_1078,N_1324);
or U1623 (N_1623,N_1307,N_853);
nand U1624 (N_1624,N_1016,N_856);
and U1625 (N_1625,N_1120,N_886);
and U1626 (N_1626,N_844,N_1014);
and U1627 (N_1627,N_956,N_1173);
nand U1628 (N_1628,N_1010,N_1292);
or U1629 (N_1629,N_1124,N_864);
and U1630 (N_1630,N_1336,N_789);
and U1631 (N_1631,N_1453,N_1409);
xor U1632 (N_1632,N_1157,N_786);
or U1633 (N_1633,N_1487,N_842);
and U1634 (N_1634,N_1396,N_1170);
or U1635 (N_1635,N_1312,N_1076);
and U1636 (N_1636,N_811,N_895);
or U1637 (N_1637,N_1098,N_1113);
nor U1638 (N_1638,N_888,N_1193);
and U1639 (N_1639,N_940,N_1399);
or U1640 (N_1640,N_1163,N_1131);
nor U1641 (N_1641,N_1299,N_1369);
or U1642 (N_1642,N_1067,N_1225);
nand U1643 (N_1643,N_1377,N_1478);
nor U1644 (N_1644,N_993,N_1329);
nand U1645 (N_1645,N_1150,N_1064);
and U1646 (N_1646,N_1460,N_838);
or U1647 (N_1647,N_832,N_826);
or U1648 (N_1648,N_1259,N_1024);
nor U1649 (N_1649,N_1043,N_1370);
nor U1650 (N_1650,N_1129,N_1322);
or U1651 (N_1651,N_1433,N_1424);
or U1652 (N_1652,N_1235,N_865);
or U1653 (N_1653,N_1471,N_1255);
and U1654 (N_1654,N_1211,N_1332);
or U1655 (N_1655,N_1152,N_1451);
nor U1656 (N_1656,N_946,N_815);
nand U1657 (N_1657,N_775,N_913);
or U1658 (N_1658,N_1458,N_799);
or U1659 (N_1659,N_891,N_1083);
and U1660 (N_1660,N_1217,N_1230);
and U1661 (N_1661,N_1056,N_1135);
or U1662 (N_1662,N_1339,N_931);
nor U1663 (N_1663,N_982,N_937);
nor U1664 (N_1664,N_1117,N_758);
and U1665 (N_1665,N_1153,N_1057);
or U1666 (N_1666,N_768,N_1316);
nor U1667 (N_1667,N_1038,N_1059);
xor U1668 (N_1668,N_816,N_1266);
or U1669 (N_1669,N_823,N_1272);
and U1670 (N_1670,N_1094,N_1488);
or U1671 (N_1671,N_845,N_1435);
and U1672 (N_1672,N_871,N_1115);
and U1673 (N_1673,N_991,N_803);
and U1674 (N_1674,N_1480,N_1297);
nand U1675 (N_1675,N_1214,N_1204);
nand U1676 (N_1676,N_868,N_889);
or U1677 (N_1677,N_897,N_1472);
or U1678 (N_1678,N_1190,N_1037);
or U1679 (N_1679,N_1262,N_939);
or U1680 (N_1680,N_870,N_915);
xnor U1681 (N_1681,N_925,N_1264);
or U1682 (N_1682,N_787,N_957);
nand U1683 (N_1683,N_883,N_998);
or U1684 (N_1684,N_833,N_1287);
and U1685 (N_1685,N_1213,N_794);
or U1686 (N_1686,N_769,N_1009);
nor U1687 (N_1687,N_764,N_1418);
and U1688 (N_1688,N_757,N_1166);
or U1689 (N_1689,N_970,N_1151);
or U1690 (N_1690,N_1053,N_846);
or U1691 (N_1691,N_1406,N_1395);
and U1692 (N_1692,N_1455,N_1479);
or U1693 (N_1693,N_1241,N_1397);
nor U1694 (N_1694,N_1413,N_1137);
nand U1695 (N_1695,N_1353,N_963);
nor U1696 (N_1696,N_1338,N_822);
or U1697 (N_1697,N_1116,N_1405);
and U1698 (N_1698,N_1243,N_928);
nand U1699 (N_1699,N_906,N_1200);
nor U1700 (N_1700,N_988,N_1248);
or U1701 (N_1701,N_1169,N_780);
nor U1702 (N_1702,N_1301,N_821);
nor U1703 (N_1703,N_1147,N_1285);
nor U1704 (N_1704,N_1240,N_849);
xnor U1705 (N_1705,N_994,N_992);
nand U1706 (N_1706,N_1392,N_1162);
nor U1707 (N_1707,N_955,N_1355);
nand U1708 (N_1708,N_983,N_772);
nor U1709 (N_1709,N_1207,N_1298);
and U1710 (N_1710,N_1199,N_1380);
or U1711 (N_1711,N_1417,N_1102);
or U1712 (N_1712,N_1195,N_1018);
or U1713 (N_1713,N_1263,N_1196);
or U1714 (N_1714,N_1454,N_784);
or U1715 (N_1715,N_783,N_1103);
and U1716 (N_1716,N_1104,N_954);
nor U1717 (N_1717,N_945,N_1229);
nand U1718 (N_1718,N_1239,N_1290);
or U1719 (N_1719,N_827,N_1184);
nand U1720 (N_1720,N_1354,N_917);
nor U1721 (N_1721,N_975,N_1289);
nor U1722 (N_1722,N_1286,N_1040);
and U1723 (N_1723,N_1491,N_1440);
nor U1724 (N_1724,N_1046,N_1461);
nor U1725 (N_1725,N_995,N_929);
nor U1726 (N_1726,N_1342,N_966);
and U1727 (N_1727,N_1385,N_1303);
or U1728 (N_1728,N_1172,N_804);
and U1729 (N_1729,N_790,N_857);
or U1730 (N_1730,N_872,N_1428);
and U1731 (N_1731,N_1318,N_1261);
and U1732 (N_1732,N_1256,N_1314);
nor U1733 (N_1733,N_997,N_944);
or U1734 (N_1734,N_766,N_892);
and U1735 (N_1735,N_961,N_1208);
or U1736 (N_1736,N_1408,N_1072);
or U1737 (N_1737,N_1493,N_770);
nand U1738 (N_1738,N_1343,N_1445);
or U1739 (N_1739,N_1189,N_1142);
or U1740 (N_1740,N_1035,N_797);
nand U1741 (N_1741,N_795,N_884);
nand U1742 (N_1742,N_755,N_1281);
nor U1743 (N_1743,N_1411,N_1068);
nand U1744 (N_1744,N_1238,N_1144);
xor U1745 (N_1745,N_1047,N_1357);
and U1746 (N_1746,N_1269,N_840);
or U1747 (N_1747,N_1203,N_1401);
nor U1748 (N_1748,N_1271,N_1226);
or U1749 (N_1749,N_1404,N_855);
nand U1750 (N_1750,N_1101,N_1133);
and U1751 (N_1751,N_1359,N_922);
or U1752 (N_1752,N_1485,N_1274);
nor U1753 (N_1753,N_1335,N_1277);
nand U1754 (N_1754,N_1340,N_1419);
and U1755 (N_1755,N_813,N_981);
nor U1756 (N_1756,N_1410,N_1127);
and U1757 (N_1757,N_1430,N_1209);
nand U1758 (N_1758,N_860,N_760);
nand U1759 (N_1759,N_1156,N_1486);
nand U1760 (N_1760,N_1223,N_791);
nor U1761 (N_1761,N_1107,N_1304);
nor U1762 (N_1762,N_1400,N_1498);
xnor U1763 (N_1763,N_1423,N_1080);
or U1764 (N_1764,N_1441,N_1434);
and U1765 (N_1765,N_1295,N_902);
or U1766 (N_1766,N_763,N_967);
and U1767 (N_1767,N_750,N_1007);
or U1768 (N_1768,N_867,N_1334);
nand U1769 (N_1769,N_1305,N_800);
nor U1770 (N_1770,N_1381,N_1118);
nor U1771 (N_1771,N_839,N_812);
or U1772 (N_1772,N_1119,N_843);
nand U1773 (N_1773,N_1215,N_1448);
nor U1774 (N_1774,N_773,N_1065);
or U1775 (N_1775,N_1231,N_866);
nor U1776 (N_1776,N_765,N_1308);
nand U1777 (N_1777,N_1055,N_1070);
nor U1778 (N_1778,N_1362,N_1315);
or U1779 (N_1779,N_1345,N_1375);
or U1780 (N_1780,N_898,N_1407);
and U1781 (N_1781,N_951,N_1030);
nor U1782 (N_1782,N_911,N_1096);
and U1783 (N_1783,N_1227,N_916);
or U1784 (N_1784,N_1276,N_1350);
or U1785 (N_1785,N_861,N_1183);
nand U1786 (N_1786,N_782,N_926);
or U1787 (N_1787,N_933,N_1364);
nand U1788 (N_1788,N_1191,N_850);
nor U1789 (N_1789,N_919,N_1245);
and U1790 (N_1790,N_949,N_1087);
nor U1791 (N_1791,N_847,N_1003);
nor U1792 (N_1792,N_1032,N_1106);
nor U1793 (N_1793,N_942,N_953);
nor U1794 (N_1794,N_1233,N_1344);
or U1795 (N_1795,N_1022,N_1099);
nor U1796 (N_1796,N_1442,N_976);
nand U1797 (N_1797,N_936,N_971);
nor U1798 (N_1798,N_908,N_793);
nor U1799 (N_1799,N_1258,N_1000);
or U1800 (N_1800,N_1042,N_1282);
or U1801 (N_1801,N_1145,N_1139);
and U1802 (N_1802,N_1062,N_1141);
and U1803 (N_1803,N_808,N_903);
nand U1804 (N_1804,N_1463,N_1088);
nor U1805 (N_1805,N_1349,N_756);
xor U1806 (N_1806,N_1496,N_901);
and U1807 (N_1807,N_1473,N_910);
nand U1808 (N_1808,N_779,N_1394);
nor U1809 (N_1809,N_1372,N_1090);
nor U1810 (N_1810,N_960,N_809);
xnor U1811 (N_1811,N_1093,N_1320);
or U1812 (N_1812,N_1437,N_974);
nor U1813 (N_1813,N_923,N_1317);
nor U1814 (N_1814,N_882,N_1013);
and U1815 (N_1815,N_932,N_1045);
and U1816 (N_1816,N_1431,N_1039);
nand U1817 (N_1817,N_1328,N_999);
nor U1818 (N_1818,N_1232,N_1321);
or U1819 (N_1819,N_904,N_912);
nand U1820 (N_1820,N_1257,N_950);
nand U1821 (N_1821,N_817,N_1398);
nor U1822 (N_1822,N_938,N_1041);
or U1823 (N_1823,N_1310,N_1111);
nand U1824 (N_1824,N_1044,N_1327);
or U1825 (N_1825,N_781,N_1323);
or U1826 (N_1826,N_1205,N_1008);
nor U1827 (N_1827,N_777,N_1154);
or U1828 (N_1828,N_1234,N_1132);
and U1829 (N_1829,N_1494,N_1346);
nor U1830 (N_1830,N_1499,N_918);
or U1831 (N_1831,N_1221,N_1174);
or U1832 (N_1832,N_1218,N_1294);
or U1833 (N_1833,N_1136,N_778);
or U1834 (N_1834,N_1309,N_854);
and U1835 (N_1835,N_1155,N_1459);
and U1836 (N_1836,N_1492,N_1291);
or U1837 (N_1837,N_1192,N_761);
nand U1838 (N_1838,N_1060,N_1177);
or U1839 (N_1839,N_1456,N_1270);
nor U1840 (N_1840,N_977,N_1386);
and U1841 (N_1841,N_1054,N_1464);
and U1842 (N_1842,N_828,N_1452);
nor U1843 (N_1843,N_796,N_1201);
and U1844 (N_1844,N_894,N_1028);
nand U1845 (N_1845,N_927,N_1075);
or U1846 (N_1846,N_1237,N_1198);
nor U1847 (N_1847,N_1236,N_1051);
and U1848 (N_1848,N_1210,N_851);
xnor U1849 (N_1849,N_1033,N_1403);
nand U1850 (N_1850,N_1467,N_1176);
and U1851 (N_1851,N_1273,N_831);
nand U1852 (N_1852,N_1330,N_1220);
or U1853 (N_1853,N_788,N_1058);
or U1854 (N_1854,N_841,N_759);
nor U1855 (N_1855,N_1114,N_752);
nand U1856 (N_1856,N_1477,N_880);
nor U1857 (N_1857,N_1439,N_1311);
or U1858 (N_1858,N_1019,N_1017);
or U1859 (N_1859,N_1284,N_1001);
xnor U1860 (N_1860,N_753,N_1371);
and U1861 (N_1861,N_968,N_958);
and U1862 (N_1862,N_996,N_1482);
nor U1863 (N_1863,N_1066,N_814);
nor U1864 (N_1864,N_1160,N_879);
nor U1865 (N_1865,N_1365,N_1483);
nor U1866 (N_1866,N_1360,N_1143);
nand U1867 (N_1867,N_1034,N_1495);
and U1868 (N_1868,N_1179,N_893);
nand U1869 (N_1869,N_1242,N_1161);
nor U1870 (N_1870,N_1251,N_1110);
and U1871 (N_1871,N_1379,N_1300);
nor U1872 (N_1872,N_948,N_1333);
or U1873 (N_1873,N_1049,N_1376);
nor U1874 (N_1874,N_1125,N_935);
and U1875 (N_1875,N_1318,N_1355);
and U1876 (N_1876,N_1410,N_1291);
or U1877 (N_1877,N_773,N_987);
or U1878 (N_1878,N_1475,N_1243);
and U1879 (N_1879,N_824,N_1091);
nand U1880 (N_1880,N_980,N_929);
nor U1881 (N_1881,N_1357,N_1077);
nor U1882 (N_1882,N_1376,N_1402);
nand U1883 (N_1883,N_1394,N_920);
or U1884 (N_1884,N_1452,N_955);
nand U1885 (N_1885,N_948,N_1245);
nor U1886 (N_1886,N_1491,N_1389);
nand U1887 (N_1887,N_867,N_1487);
or U1888 (N_1888,N_890,N_894);
and U1889 (N_1889,N_984,N_1187);
nand U1890 (N_1890,N_972,N_798);
nor U1891 (N_1891,N_1473,N_1271);
and U1892 (N_1892,N_1345,N_1383);
nor U1893 (N_1893,N_1030,N_1428);
nand U1894 (N_1894,N_1328,N_1164);
nand U1895 (N_1895,N_1126,N_785);
nor U1896 (N_1896,N_1493,N_816);
or U1897 (N_1897,N_958,N_1233);
and U1898 (N_1898,N_759,N_1374);
or U1899 (N_1899,N_1121,N_1056);
nand U1900 (N_1900,N_848,N_1498);
and U1901 (N_1901,N_1425,N_1252);
nand U1902 (N_1902,N_1405,N_999);
nor U1903 (N_1903,N_1232,N_1170);
xnor U1904 (N_1904,N_855,N_785);
or U1905 (N_1905,N_1043,N_1497);
nor U1906 (N_1906,N_1012,N_874);
nor U1907 (N_1907,N_788,N_925);
nand U1908 (N_1908,N_900,N_1289);
and U1909 (N_1909,N_947,N_1071);
and U1910 (N_1910,N_818,N_1270);
nand U1911 (N_1911,N_1217,N_1456);
or U1912 (N_1912,N_896,N_1011);
or U1913 (N_1913,N_1187,N_1158);
nor U1914 (N_1914,N_754,N_881);
nor U1915 (N_1915,N_756,N_990);
or U1916 (N_1916,N_963,N_1236);
nor U1917 (N_1917,N_787,N_932);
or U1918 (N_1918,N_1265,N_1108);
nand U1919 (N_1919,N_1393,N_988);
or U1920 (N_1920,N_1141,N_1159);
and U1921 (N_1921,N_1420,N_850);
nor U1922 (N_1922,N_1407,N_1146);
nand U1923 (N_1923,N_1450,N_890);
and U1924 (N_1924,N_1146,N_1490);
nand U1925 (N_1925,N_760,N_1474);
xor U1926 (N_1926,N_1428,N_965);
nor U1927 (N_1927,N_785,N_1200);
and U1928 (N_1928,N_775,N_1424);
or U1929 (N_1929,N_940,N_1367);
and U1930 (N_1930,N_769,N_991);
nor U1931 (N_1931,N_1288,N_1169);
nand U1932 (N_1932,N_1143,N_1119);
nand U1933 (N_1933,N_1346,N_813);
and U1934 (N_1934,N_1248,N_1032);
nor U1935 (N_1935,N_1136,N_1059);
nor U1936 (N_1936,N_1042,N_935);
and U1937 (N_1937,N_913,N_1257);
nor U1938 (N_1938,N_1326,N_948);
nand U1939 (N_1939,N_1160,N_1088);
nand U1940 (N_1940,N_1374,N_1023);
nand U1941 (N_1941,N_1181,N_919);
nor U1942 (N_1942,N_779,N_999);
nor U1943 (N_1943,N_1378,N_770);
nor U1944 (N_1944,N_760,N_905);
and U1945 (N_1945,N_1079,N_1223);
nor U1946 (N_1946,N_772,N_1141);
nor U1947 (N_1947,N_836,N_1492);
and U1948 (N_1948,N_1314,N_1446);
nor U1949 (N_1949,N_1175,N_1275);
nor U1950 (N_1950,N_930,N_1056);
nand U1951 (N_1951,N_834,N_1059);
nand U1952 (N_1952,N_968,N_1018);
nor U1953 (N_1953,N_854,N_1410);
xor U1954 (N_1954,N_1078,N_1417);
and U1955 (N_1955,N_1411,N_803);
nand U1956 (N_1956,N_996,N_943);
or U1957 (N_1957,N_1047,N_1406);
nand U1958 (N_1958,N_1050,N_766);
nand U1959 (N_1959,N_945,N_884);
nor U1960 (N_1960,N_1325,N_993);
nor U1961 (N_1961,N_889,N_1042);
and U1962 (N_1962,N_1440,N_1220);
nand U1963 (N_1963,N_1099,N_1160);
or U1964 (N_1964,N_1458,N_768);
or U1965 (N_1965,N_1183,N_938);
or U1966 (N_1966,N_1207,N_996);
and U1967 (N_1967,N_934,N_1277);
nand U1968 (N_1968,N_827,N_1403);
or U1969 (N_1969,N_1024,N_940);
nand U1970 (N_1970,N_1354,N_1481);
nand U1971 (N_1971,N_1484,N_765);
nor U1972 (N_1972,N_816,N_1153);
xor U1973 (N_1973,N_1006,N_963);
or U1974 (N_1974,N_1128,N_1036);
nor U1975 (N_1975,N_1173,N_834);
nor U1976 (N_1976,N_1196,N_988);
nor U1977 (N_1977,N_802,N_1097);
and U1978 (N_1978,N_800,N_1135);
nand U1979 (N_1979,N_955,N_1031);
nand U1980 (N_1980,N_1304,N_830);
xor U1981 (N_1981,N_933,N_1063);
and U1982 (N_1982,N_1206,N_978);
nand U1983 (N_1983,N_1021,N_1262);
nand U1984 (N_1984,N_877,N_1488);
nor U1985 (N_1985,N_908,N_769);
or U1986 (N_1986,N_1235,N_870);
and U1987 (N_1987,N_1041,N_1344);
nor U1988 (N_1988,N_882,N_1305);
and U1989 (N_1989,N_1164,N_1203);
nand U1990 (N_1990,N_1026,N_1147);
and U1991 (N_1991,N_1273,N_1480);
or U1992 (N_1992,N_1135,N_1251);
nand U1993 (N_1993,N_1439,N_1070);
and U1994 (N_1994,N_1333,N_1278);
xor U1995 (N_1995,N_1363,N_815);
and U1996 (N_1996,N_911,N_1259);
nor U1997 (N_1997,N_1119,N_1095);
nand U1998 (N_1998,N_946,N_1475);
or U1999 (N_1999,N_1404,N_1066);
nand U2000 (N_2000,N_1242,N_971);
or U2001 (N_2001,N_974,N_789);
and U2002 (N_2002,N_1448,N_1239);
or U2003 (N_2003,N_1424,N_818);
nor U2004 (N_2004,N_1474,N_984);
or U2005 (N_2005,N_1361,N_1294);
nor U2006 (N_2006,N_914,N_964);
nand U2007 (N_2007,N_807,N_1118);
or U2008 (N_2008,N_1481,N_1159);
nand U2009 (N_2009,N_1455,N_856);
and U2010 (N_2010,N_1397,N_1185);
nor U2011 (N_2011,N_864,N_820);
nor U2012 (N_2012,N_912,N_1330);
and U2013 (N_2013,N_1169,N_1462);
and U2014 (N_2014,N_889,N_1360);
and U2015 (N_2015,N_837,N_1142);
and U2016 (N_2016,N_997,N_1454);
and U2017 (N_2017,N_1138,N_1488);
xor U2018 (N_2018,N_1345,N_1065);
nand U2019 (N_2019,N_804,N_1167);
nor U2020 (N_2020,N_1020,N_1094);
and U2021 (N_2021,N_1290,N_1320);
or U2022 (N_2022,N_937,N_1053);
and U2023 (N_2023,N_1139,N_1411);
nand U2024 (N_2024,N_1447,N_1047);
nor U2025 (N_2025,N_1294,N_1304);
nand U2026 (N_2026,N_764,N_1082);
nor U2027 (N_2027,N_795,N_870);
or U2028 (N_2028,N_780,N_998);
nor U2029 (N_2029,N_935,N_1120);
or U2030 (N_2030,N_878,N_1279);
nor U2031 (N_2031,N_1416,N_927);
nor U2032 (N_2032,N_1098,N_1021);
or U2033 (N_2033,N_1378,N_1373);
nand U2034 (N_2034,N_888,N_1377);
nor U2035 (N_2035,N_1342,N_1183);
and U2036 (N_2036,N_829,N_1069);
nand U2037 (N_2037,N_1184,N_1270);
nand U2038 (N_2038,N_1453,N_756);
nor U2039 (N_2039,N_899,N_787);
and U2040 (N_2040,N_1245,N_874);
nor U2041 (N_2041,N_1290,N_1039);
or U2042 (N_2042,N_870,N_1051);
and U2043 (N_2043,N_1146,N_858);
and U2044 (N_2044,N_1160,N_1307);
nand U2045 (N_2045,N_950,N_1370);
and U2046 (N_2046,N_1227,N_997);
and U2047 (N_2047,N_1357,N_1350);
nand U2048 (N_2048,N_1161,N_1111);
or U2049 (N_2049,N_764,N_1254);
or U2050 (N_2050,N_1026,N_1155);
and U2051 (N_2051,N_808,N_1209);
nand U2052 (N_2052,N_1138,N_1235);
nor U2053 (N_2053,N_1344,N_858);
nand U2054 (N_2054,N_1287,N_992);
nor U2055 (N_2055,N_1282,N_1215);
or U2056 (N_2056,N_1096,N_1409);
nor U2057 (N_2057,N_1476,N_1061);
or U2058 (N_2058,N_901,N_1057);
nand U2059 (N_2059,N_775,N_1263);
nor U2060 (N_2060,N_1394,N_1347);
nor U2061 (N_2061,N_864,N_861);
xnor U2062 (N_2062,N_1076,N_993);
nand U2063 (N_2063,N_900,N_1283);
or U2064 (N_2064,N_1333,N_806);
nand U2065 (N_2065,N_1392,N_831);
nand U2066 (N_2066,N_753,N_1379);
nor U2067 (N_2067,N_1170,N_1324);
nand U2068 (N_2068,N_1177,N_1011);
or U2069 (N_2069,N_1422,N_1244);
nand U2070 (N_2070,N_1316,N_1062);
or U2071 (N_2071,N_986,N_1420);
xnor U2072 (N_2072,N_1484,N_1155);
nand U2073 (N_2073,N_1077,N_1133);
nor U2074 (N_2074,N_1010,N_1388);
and U2075 (N_2075,N_899,N_1370);
nand U2076 (N_2076,N_1048,N_1358);
nand U2077 (N_2077,N_1498,N_1010);
or U2078 (N_2078,N_1050,N_1313);
nor U2079 (N_2079,N_822,N_929);
nor U2080 (N_2080,N_1482,N_1211);
and U2081 (N_2081,N_907,N_1333);
nand U2082 (N_2082,N_995,N_894);
or U2083 (N_2083,N_1076,N_1141);
nand U2084 (N_2084,N_960,N_961);
and U2085 (N_2085,N_1414,N_858);
nand U2086 (N_2086,N_1009,N_1211);
nor U2087 (N_2087,N_874,N_1082);
xnor U2088 (N_2088,N_943,N_970);
and U2089 (N_2089,N_1295,N_1419);
or U2090 (N_2090,N_1489,N_1060);
and U2091 (N_2091,N_1498,N_1118);
xnor U2092 (N_2092,N_841,N_939);
nand U2093 (N_2093,N_1010,N_1075);
nor U2094 (N_2094,N_1306,N_1060);
nor U2095 (N_2095,N_1091,N_1449);
nand U2096 (N_2096,N_1109,N_1345);
or U2097 (N_2097,N_1417,N_855);
or U2098 (N_2098,N_1420,N_1013);
or U2099 (N_2099,N_1402,N_855);
nor U2100 (N_2100,N_1178,N_1379);
nor U2101 (N_2101,N_970,N_1200);
and U2102 (N_2102,N_897,N_1039);
nor U2103 (N_2103,N_844,N_1086);
nand U2104 (N_2104,N_874,N_985);
nor U2105 (N_2105,N_1344,N_1353);
nand U2106 (N_2106,N_920,N_837);
and U2107 (N_2107,N_1124,N_1047);
nor U2108 (N_2108,N_1146,N_1132);
or U2109 (N_2109,N_1207,N_1440);
or U2110 (N_2110,N_1101,N_1060);
nand U2111 (N_2111,N_1370,N_836);
and U2112 (N_2112,N_1017,N_1289);
nand U2113 (N_2113,N_1168,N_859);
nand U2114 (N_2114,N_1357,N_988);
nor U2115 (N_2115,N_1396,N_1453);
xor U2116 (N_2116,N_978,N_1133);
or U2117 (N_2117,N_1338,N_1015);
or U2118 (N_2118,N_1078,N_1323);
nand U2119 (N_2119,N_817,N_1033);
nand U2120 (N_2120,N_1028,N_920);
nand U2121 (N_2121,N_1143,N_1004);
and U2122 (N_2122,N_1433,N_893);
nor U2123 (N_2123,N_1169,N_1139);
nor U2124 (N_2124,N_1382,N_1361);
or U2125 (N_2125,N_1327,N_1417);
and U2126 (N_2126,N_1001,N_1349);
or U2127 (N_2127,N_1168,N_1153);
or U2128 (N_2128,N_1269,N_905);
or U2129 (N_2129,N_1155,N_1433);
nand U2130 (N_2130,N_1358,N_857);
nor U2131 (N_2131,N_1033,N_1434);
or U2132 (N_2132,N_1083,N_1461);
and U2133 (N_2133,N_1395,N_1008);
and U2134 (N_2134,N_1225,N_1319);
nand U2135 (N_2135,N_1252,N_844);
or U2136 (N_2136,N_1180,N_1376);
nand U2137 (N_2137,N_990,N_1488);
nand U2138 (N_2138,N_1463,N_1464);
and U2139 (N_2139,N_1108,N_1324);
or U2140 (N_2140,N_1376,N_1092);
nand U2141 (N_2141,N_1219,N_812);
or U2142 (N_2142,N_1386,N_784);
nand U2143 (N_2143,N_770,N_1240);
or U2144 (N_2144,N_760,N_1090);
nand U2145 (N_2145,N_1212,N_863);
or U2146 (N_2146,N_1431,N_1121);
nor U2147 (N_2147,N_1358,N_854);
or U2148 (N_2148,N_852,N_885);
or U2149 (N_2149,N_1165,N_766);
nor U2150 (N_2150,N_1175,N_1022);
nor U2151 (N_2151,N_1328,N_1473);
nor U2152 (N_2152,N_1005,N_1272);
nor U2153 (N_2153,N_824,N_973);
nor U2154 (N_2154,N_1250,N_886);
or U2155 (N_2155,N_994,N_1484);
nor U2156 (N_2156,N_871,N_942);
and U2157 (N_2157,N_1064,N_994);
or U2158 (N_2158,N_1164,N_1449);
and U2159 (N_2159,N_1019,N_1134);
and U2160 (N_2160,N_926,N_1279);
or U2161 (N_2161,N_1035,N_768);
and U2162 (N_2162,N_1324,N_889);
nor U2163 (N_2163,N_1485,N_918);
nor U2164 (N_2164,N_1384,N_1214);
and U2165 (N_2165,N_1428,N_801);
and U2166 (N_2166,N_1292,N_750);
nand U2167 (N_2167,N_821,N_1092);
nor U2168 (N_2168,N_971,N_1203);
or U2169 (N_2169,N_1434,N_1028);
or U2170 (N_2170,N_1303,N_982);
and U2171 (N_2171,N_1001,N_1420);
nand U2172 (N_2172,N_1203,N_809);
nor U2173 (N_2173,N_1440,N_1292);
and U2174 (N_2174,N_1133,N_998);
or U2175 (N_2175,N_776,N_993);
nor U2176 (N_2176,N_763,N_1259);
nor U2177 (N_2177,N_1009,N_1217);
nor U2178 (N_2178,N_902,N_851);
and U2179 (N_2179,N_1283,N_875);
nor U2180 (N_2180,N_944,N_1291);
and U2181 (N_2181,N_1062,N_982);
and U2182 (N_2182,N_752,N_855);
nand U2183 (N_2183,N_1286,N_931);
nor U2184 (N_2184,N_899,N_1008);
nor U2185 (N_2185,N_1056,N_847);
or U2186 (N_2186,N_787,N_845);
and U2187 (N_2187,N_952,N_953);
nand U2188 (N_2188,N_1090,N_779);
nand U2189 (N_2189,N_967,N_866);
nand U2190 (N_2190,N_1475,N_810);
and U2191 (N_2191,N_1353,N_1287);
nor U2192 (N_2192,N_897,N_1232);
nor U2193 (N_2193,N_1273,N_1072);
and U2194 (N_2194,N_1121,N_763);
and U2195 (N_2195,N_1216,N_1351);
and U2196 (N_2196,N_1059,N_1488);
nor U2197 (N_2197,N_1036,N_881);
or U2198 (N_2198,N_1363,N_1405);
nand U2199 (N_2199,N_767,N_780);
nand U2200 (N_2200,N_918,N_1140);
or U2201 (N_2201,N_1403,N_892);
or U2202 (N_2202,N_1076,N_822);
nand U2203 (N_2203,N_1368,N_1091);
nor U2204 (N_2204,N_1426,N_778);
and U2205 (N_2205,N_1031,N_1137);
or U2206 (N_2206,N_1272,N_871);
and U2207 (N_2207,N_1435,N_847);
and U2208 (N_2208,N_1461,N_1155);
or U2209 (N_2209,N_1258,N_852);
nand U2210 (N_2210,N_964,N_1418);
and U2211 (N_2211,N_766,N_1002);
nand U2212 (N_2212,N_1046,N_1182);
nor U2213 (N_2213,N_1461,N_1361);
or U2214 (N_2214,N_1242,N_1258);
and U2215 (N_2215,N_1237,N_1155);
or U2216 (N_2216,N_980,N_1136);
or U2217 (N_2217,N_1027,N_880);
xor U2218 (N_2218,N_1118,N_1260);
or U2219 (N_2219,N_1294,N_1061);
or U2220 (N_2220,N_1209,N_1215);
nand U2221 (N_2221,N_1342,N_858);
nor U2222 (N_2222,N_1110,N_1215);
xnor U2223 (N_2223,N_878,N_1337);
nor U2224 (N_2224,N_979,N_776);
nor U2225 (N_2225,N_1357,N_1163);
nor U2226 (N_2226,N_1077,N_919);
and U2227 (N_2227,N_1406,N_1147);
and U2228 (N_2228,N_1380,N_1016);
or U2229 (N_2229,N_923,N_974);
nor U2230 (N_2230,N_1142,N_1049);
nor U2231 (N_2231,N_1329,N_1249);
or U2232 (N_2232,N_1398,N_940);
and U2233 (N_2233,N_1050,N_1383);
and U2234 (N_2234,N_1132,N_1454);
nor U2235 (N_2235,N_778,N_759);
nand U2236 (N_2236,N_786,N_1498);
or U2237 (N_2237,N_1294,N_908);
nand U2238 (N_2238,N_1152,N_816);
and U2239 (N_2239,N_1335,N_1258);
or U2240 (N_2240,N_1360,N_928);
and U2241 (N_2241,N_1121,N_1087);
nand U2242 (N_2242,N_1266,N_1257);
nor U2243 (N_2243,N_1154,N_1494);
nand U2244 (N_2244,N_1024,N_1364);
or U2245 (N_2245,N_936,N_794);
and U2246 (N_2246,N_1023,N_1420);
nor U2247 (N_2247,N_1011,N_978);
and U2248 (N_2248,N_1339,N_1172);
nand U2249 (N_2249,N_1258,N_845);
nor U2250 (N_2250,N_1716,N_1857);
and U2251 (N_2251,N_2214,N_1930);
nand U2252 (N_2252,N_2128,N_2200);
or U2253 (N_2253,N_2161,N_2087);
nand U2254 (N_2254,N_2219,N_1636);
nand U2255 (N_2255,N_2053,N_1907);
or U2256 (N_2256,N_1964,N_1721);
nand U2257 (N_2257,N_1541,N_2061);
nor U2258 (N_2258,N_1995,N_1823);
nand U2259 (N_2259,N_1934,N_1776);
nor U2260 (N_2260,N_1908,N_2040);
and U2261 (N_2261,N_1531,N_1708);
and U2262 (N_2262,N_1609,N_1566);
nand U2263 (N_2263,N_1789,N_1577);
nor U2264 (N_2264,N_1820,N_1505);
xnor U2265 (N_2265,N_1712,N_2080);
or U2266 (N_2266,N_2198,N_2017);
nor U2267 (N_2267,N_1717,N_1524);
nand U2268 (N_2268,N_1956,N_2036);
or U2269 (N_2269,N_1791,N_1944);
or U2270 (N_2270,N_2137,N_1644);
nand U2271 (N_2271,N_1991,N_1681);
or U2272 (N_2272,N_2136,N_2066);
nor U2273 (N_2273,N_2231,N_1905);
nand U2274 (N_2274,N_2167,N_1549);
and U2275 (N_2275,N_2000,N_2228);
or U2276 (N_2276,N_2181,N_2222);
and U2277 (N_2277,N_1713,N_1616);
and U2278 (N_2278,N_2232,N_1839);
or U2279 (N_2279,N_1884,N_1805);
nand U2280 (N_2280,N_1766,N_2116);
or U2281 (N_2281,N_1928,N_1724);
nor U2282 (N_2282,N_1831,N_1952);
nor U2283 (N_2283,N_1784,N_1570);
nand U2284 (N_2284,N_1645,N_2035);
and U2285 (N_2285,N_1657,N_1601);
or U2286 (N_2286,N_1565,N_1909);
nand U2287 (N_2287,N_1556,N_1591);
nor U2288 (N_2288,N_2224,N_2212);
and U2289 (N_2289,N_1774,N_1604);
or U2290 (N_2290,N_1868,N_1904);
nor U2291 (N_2291,N_2009,N_1573);
nor U2292 (N_2292,N_1850,N_1667);
nand U2293 (N_2293,N_1659,N_2203);
xnor U2294 (N_2294,N_2013,N_2074);
or U2295 (N_2295,N_1661,N_1688);
nor U2296 (N_2296,N_1687,N_1611);
xor U2297 (N_2297,N_1989,N_1792);
or U2298 (N_2298,N_2108,N_2234);
or U2299 (N_2299,N_2183,N_1624);
and U2300 (N_2300,N_2113,N_1899);
xor U2301 (N_2301,N_1590,N_1970);
and U2302 (N_2302,N_1895,N_1523);
nand U2303 (N_2303,N_1802,N_2075);
nand U2304 (N_2304,N_1910,N_2105);
nor U2305 (N_2305,N_1563,N_1870);
nor U2306 (N_2306,N_1918,N_2204);
and U2307 (N_2307,N_2029,N_1711);
or U2308 (N_2308,N_1945,N_1759);
or U2309 (N_2309,N_2059,N_2196);
and U2310 (N_2310,N_1513,N_1927);
nand U2311 (N_2311,N_2072,N_2102);
or U2312 (N_2312,N_1727,N_1822);
or U2313 (N_2313,N_1651,N_2182);
nor U2314 (N_2314,N_2239,N_1740);
or U2315 (N_2315,N_2001,N_2188);
nand U2316 (N_2316,N_1592,N_2099);
and U2317 (N_2317,N_2190,N_1769);
or U2318 (N_2318,N_1979,N_1933);
or U2319 (N_2319,N_1548,N_1569);
and U2320 (N_2320,N_1915,N_1957);
and U2321 (N_2321,N_2071,N_1954);
and U2322 (N_2322,N_1856,N_1693);
or U2323 (N_2323,N_2028,N_1682);
nand U2324 (N_2324,N_1521,N_2127);
and U2325 (N_2325,N_1575,N_2153);
nand U2326 (N_2326,N_2097,N_2078);
and U2327 (N_2327,N_1834,N_1745);
nand U2328 (N_2328,N_1735,N_2191);
nand U2329 (N_2329,N_1939,N_1750);
nand U2330 (N_2330,N_1650,N_1517);
or U2331 (N_2331,N_1818,N_1699);
and U2332 (N_2332,N_1983,N_2245);
nand U2333 (N_2333,N_2151,N_2042);
nand U2334 (N_2334,N_2165,N_1571);
and U2335 (N_2335,N_2133,N_1963);
and U2336 (N_2336,N_1900,N_1793);
nand U2337 (N_2337,N_2207,N_1840);
and U2338 (N_2338,N_1958,N_1935);
nand U2339 (N_2339,N_1720,N_2034);
xnor U2340 (N_2340,N_2062,N_2168);
nand U2341 (N_2341,N_1864,N_2041);
nor U2342 (N_2342,N_1723,N_1754);
nand U2343 (N_2343,N_2077,N_1700);
nor U2344 (N_2344,N_2082,N_1996);
or U2345 (N_2345,N_1536,N_1885);
nand U2346 (N_2346,N_2177,N_1828);
or U2347 (N_2347,N_1937,N_2152);
nor U2348 (N_2348,N_1674,N_1648);
and U2349 (N_2349,N_1883,N_1982);
or U2350 (N_2350,N_1898,N_1528);
or U2351 (N_2351,N_1972,N_1782);
and U2352 (N_2352,N_1732,N_1862);
or U2353 (N_2353,N_1965,N_1518);
and U2354 (N_2354,N_1973,N_1755);
or U2355 (N_2355,N_1603,N_2197);
xor U2356 (N_2356,N_1730,N_2019);
or U2357 (N_2357,N_2115,N_1877);
nor U2358 (N_2358,N_1537,N_1742);
or U2359 (N_2359,N_2103,N_2238);
and U2360 (N_2360,N_1640,N_1562);
or U2361 (N_2361,N_2049,N_2021);
or U2362 (N_2362,N_2123,N_1707);
and U2363 (N_2363,N_2006,N_1701);
nor U2364 (N_2364,N_1837,N_2223);
and U2365 (N_2365,N_2195,N_2032);
nand U2366 (N_2366,N_1623,N_1704);
and U2367 (N_2367,N_1599,N_1653);
and U2368 (N_2368,N_2144,N_1753);
or U2369 (N_2369,N_2106,N_2217);
nand U2370 (N_2370,N_1764,N_1913);
nor U2371 (N_2371,N_1986,N_1586);
and U2372 (N_2372,N_2187,N_2026);
nor U2373 (N_2373,N_1859,N_1627);
and U2374 (N_2374,N_1941,N_1819);
nand U2375 (N_2375,N_1916,N_1737);
nor U2376 (N_2376,N_2159,N_1874);
nand U2377 (N_2377,N_1946,N_2112);
nand U2378 (N_2378,N_2038,N_1760);
or U2379 (N_2379,N_2226,N_1649);
nor U2380 (N_2380,N_1705,N_2056);
and U2381 (N_2381,N_2031,N_1980);
and U2382 (N_2382,N_1550,N_2174);
or U2383 (N_2383,N_1696,N_1635);
nand U2384 (N_2384,N_1912,N_1797);
nor U2385 (N_2385,N_1702,N_2170);
nor U2386 (N_2386,N_2084,N_1654);
nor U2387 (N_2387,N_2037,N_1588);
and U2388 (N_2388,N_2094,N_1998);
nor U2389 (N_2389,N_2155,N_2014);
and U2390 (N_2390,N_2055,N_1781);
nor U2391 (N_2391,N_1765,N_1790);
nor U2392 (N_2392,N_1558,N_2134);
nand U2393 (N_2393,N_1751,N_1576);
and U2394 (N_2394,N_1646,N_1514);
nor U2395 (N_2395,N_1555,N_1960);
or U2396 (N_2396,N_1757,N_2018);
and U2397 (N_2397,N_1775,N_1951);
and U2398 (N_2398,N_1966,N_1943);
or U2399 (N_2399,N_1844,N_1838);
and U2400 (N_2400,N_2098,N_1967);
nor U2401 (N_2401,N_1606,N_2202);
nor U2402 (N_2402,N_1929,N_1610);
nor U2403 (N_2403,N_1660,N_2160);
nor U2404 (N_2404,N_1994,N_1925);
nor U2405 (N_2405,N_1666,N_1572);
or U2406 (N_2406,N_1607,N_1690);
and U2407 (N_2407,N_1799,N_2100);
or U2408 (N_2408,N_1508,N_1999);
or U2409 (N_2409,N_2172,N_1507);
and U2410 (N_2410,N_1851,N_1677);
or U2411 (N_2411,N_2064,N_1785);
or U2412 (N_2412,N_1529,N_1692);
or U2413 (N_2413,N_1917,N_1860);
and U2414 (N_2414,N_1515,N_1605);
nor U2415 (N_2415,N_1655,N_1680);
and U2416 (N_2416,N_1798,N_2109);
and U2417 (N_2417,N_1890,N_1628);
nand U2418 (N_2418,N_1808,N_1892);
nand U2419 (N_2419,N_1530,N_2148);
nand U2420 (N_2420,N_2120,N_1997);
or U2421 (N_2421,N_1580,N_1959);
and U2422 (N_2422,N_1579,N_2068);
nand U2423 (N_2423,N_1694,N_1691);
nand U2424 (N_2424,N_2205,N_2008);
and U2425 (N_2425,N_1891,N_2206);
and U2426 (N_2426,N_1829,N_1990);
nand U2427 (N_2427,N_1843,N_2069);
and U2428 (N_2428,N_2046,N_1647);
or U2429 (N_2429,N_1906,N_1961);
or U2430 (N_2430,N_1686,N_1710);
and U2431 (N_2431,N_2119,N_1719);
nand U2432 (N_2432,N_1893,N_2060);
and U2433 (N_2433,N_2162,N_2145);
nand U2434 (N_2434,N_2089,N_2093);
nand U2435 (N_2435,N_2007,N_1855);
nor U2436 (N_2436,N_1747,N_2176);
nand U2437 (N_2437,N_2010,N_2249);
nand U2438 (N_2438,N_1779,N_1826);
or U2439 (N_2439,N_1709,N_2004);
xor U2440 (N_2440,N_2011,N_1876);
nor U2441 (N_2441,N_1638,N_1615);
and U2442 (N_2442,N_1706,N_1744);
nor U2443 (N_2443,N_1715,N_1672);
or U2444 (N_2444,N_1738,N_2107);
and U2445 (N_2445,N_1526,N_1969);
xnor U2446 (N_2446,N_1950,N_1923);
or U2447 (N_2447,N_1736,N_2233);
nand U2448 (N_2448,N_1949,N_2244);
nor U2449 (N_2449,N_2122,N_2016);
nor U2450 (N_2450,N_1633,N_1585);
nor U2451 (N_2451,N_2070,N_1903);
and U2452 (N_2452,N_1981,N_1617);
or U2453 (N_2453,N_1800,N_1796);
or U2454 (N_2454,N_2057,N_1668);
nand U2455 (N_2455,N_1889,N_1578);
nor U2456 (N_2456,N_1545,N_1564);
nor U2457 (N_2457,N_1938,N_1552);
nor U2458 (N_2458,N_2118,N_2045);
nor U2459 (N_2459,N_2237,N_1602);
or U2460 (N_2460,N_2076,N_2081);
and U2461 (N_2461,N_1920,N_1669);
nor U2462 (N_2462,N_2210,N_2091);
and U2463 (N_2463,N_1777,N_1872);
and U2464 (N_2464,N_1978,N_1863);
nor U2465 (N_2465,N_1542,N_2092);
and U2466 (N_2466,N_2012,N_2243);
or U2467 (N_2467,N_2131,N_1807);
and U2468 (N_2468,N_1675,N_1527);
nor U2469 (N_2469,N_2157,N_2114);
nor U2470 (N_2470,N_1993,N_2175);
nor U2471 (N_2471,N_1932,N_2129);
or U2472 (N_2472,N_2030,N_1984);
nand U2473 (N_2473,N_1504,N_1560);
and U2474 (N_2474,N_1684,N_1783);
nor U2475 (N_2475,N_1652,N_1871);
and U2476 (N_2476,N_1631,N_1503);
and U2477 (N_2477,N_1500,N_1832);
and U2478 (N_2478,N_2088,N_1854);
and U2479 (N_2479,N_1612,N_2229);
nor U2480 (N_2480,N_1940,N_1689);
nor U2481 (N_2481,N_1731,N_1506);
nand U2482 (N_2482,N_1985,N_2158);
and U2483 (N_2483,N_2146,N_1501);
and U2484 (N_2484,N_1845,N_1977);
and U2485 (N_2485,N_1642,N_2216);
and U2486 (N_2486,N_1830,N_1761);
or U2487 (N_2487,N_2051,N_2163);
nor U2488 (N_2488,N_1896,N_1762);
or U2489 (N_2489,N_2022,N_1914);
and U2490 (N_2490,N_1729,N_2135);
nand U2491 (N_2491,N_2058,N_1639);
nor U2492 (N_2492,N_2005,N_1583);
nand U2493 (N_2493,N_2142,N_2140);
or U2494 (N_2494,N_2213,N_1733);
or U2495 (N_2495,N_1811,N_1641);
or U2496 (N_2496,N_2117,N_2130);
or U2497 (N_2497,N_1679,N_1924);
nand U2498 (N_2498,N_2154,N_1544);
or U2499 (N_2499,N_1625,N_1812);
nand U2500 (N_2500,N_1888,N_1894);
nand U2501 (N_2501,N_1598,N_1554);
or U2502 (N_2502,N_1561,N_2166);
nand U2503 (N_2503,N_1559,N_1525);
and U2504 (N_2504,N_1875,N_2192);
or U2505 (N_2505,N_2179,N_2048);
nor U2506 (N_2506,N_1535,N_1768);
or U2507 (N_2507,N_1887,N_1614);
xor U2508 (N_2508,N_1608,N_1847);
and U2509 (N_2509,N_1533,N_2227);
or U2510 (N_2510,N_1835,N_1897);
nand U2511 (N_2511,N_1833,N_1771);
and U2512 (N_2512,N_1848,N_2242);
or U2513 (N_2513,N_2230,N_1502);
and U2514 (N_2514,N_1520,N_1936);
nor U2515 (N_2515,N_2156,N_1620);
or U2516 (N_2516,N_2024,N_1955);
nor U2517 (N_2517,N_2124,N_1516);
nand U2518 (N_2518,N_2208,N_1664);
nand U2519 (N_2519,N_2215,N_1656);
or U2520 (N_2520,N_1534,N_1663);
or U2521 (N_2521,N_1512,N_2209);
and U2522 (N_2522,N_1546,N_1836);
or U2523 (N_2523,N_2090,N_1911);
or U2524 (N_2524,N_1551,N_1522);
or U2525 (N_2525,N_1697,N_1827);
and U2526 (N_2526,N_2033,N_2065);
nand U2527 (N_2527,N_1581,N_1852);
nor U2528 (N_2528,N_1824,N_2044);
nand U2529 (N_2529,N_1795,N_1922);
nor U2530 (N_2530,N_1739,N_1821);
nor U2531 (N_2531,N_1942,N_1749);
nor U2532 (N_2532,N_1746,N_1865);
nand U2533 (N_2533,N_2079,N_2149);
nand U2534 (N_2534,N_2184,N_1589);
nand U2535 (N_2535,N_2020,N_1539);
or U2536 (N_2536,N_2147,N_1511);
or U2537 (N_2537,N_1810,N_1557);
or U2538 (N_2538,N_2139,N_1670);
nor U2539 (N_2539,N_2015,N_1629);
nor U2540 (N_2540,N_1869,N_1553);
and U2541 (N_2541,N_1596,N_1630);
and U2542 (N_2542,N_1976,N_1842);
or U2543 (N_2543,N_1718,N_1921);
nor U2544 (N_2544,N_1597,N_1816);
or U2545 (N_2545,N_2003,N_1814);
nor U2546 (N_2546,N_2111,N_1817);
or U2547 (N_2547,N_1665,N_1695);
nor U2548 (N_2548,N_2150,N_1595);
nand U2549 (N_2549,N_1787,N_1858);
xnor U2550 (N_2550,N_1770,N_2225);
nand U2551 (N_2551,N_2027,N_1987);
nor U2552 (N_2552,N_1866,N_2246);
nor U2553 (N_2553,N_1971,N_1806);
nor U2554 (N_2554,N_1974,N_1621);
and U2555 (N_2555,N_2039,N_1992);
nand U2556 (N_2556,N_1662,N_1778);
nand U2557 (N_2557,N_1634,N_1773);
or U2558 (N_2558,N_1519,N_2201);
and U2559 (N_2559,N_2050,N_2126);
and U2560 (N_2560,N_1613,N_1587);
or U2561 (N_2561,N_1809,N_1879);
or U2562 (N_2562,N_2086,N_2180);
xor U2563 (N_2563,N_1622,N_2185);
and U2564 (N_2564,N_2121,N_1815);
nor U2565 (N_2565,N_2247,N_2141);
nand U2566 (N_2566,N_1867,N_1803);
or U2567 (N_2567,N_1678,N_1538);
nor U2568 (N_2568,N_2025,N_1568);
and U2569 (N_2569,N_2104,N_1846);
and U2570 (N_2570,N_1758,N_1626);
nor U2571 (N_2571,N_1881,N_1671);
xor U2572 (N_2572,N_2002,N_2073);
nor U2573 (N_2573,N_2235,N_1804);
nand U2574 (N_2574,N_1953,N_1926);
nor U2575 (N_2575,N_2218,N_2101);
nand U2576 (N_2576,N_1988,N_2132);
or U2577 (N_2577,N_1726,N_1543);
and U2578 (N_2578,N_1801,N_1532);
nor U2579 (N_2579,N_2169,N_1861);
nand U2580 (N_2580,N_2023,N_1756);
xor U2581 (N_2581,N_2240,N_1873);
nor U2582 (N_2582,N_2052,N_2143);
nand U2583 (N_2583,N_1741,N_1947);
nor U2584 (N_2584,N_1714,N_1919);
or U2585 (N_2585,N_1825,N_1728);
nor U2586 (N_2586,N_2047,N_1673);
and U2587 (N_2587,N_2178,N_1780);
or U2588 (N_2588,N_1594,N_1841);
nand U2589 (N_2589,N_1975,N_1658);
or U2590 (N_2590,N_1725,N_1698);
and U2591 (N_2591,N_1734,N_1547);
nand U2592 (N_2592,N_2125,N_1600);
xnor U2593 (N_2593,N_1968,N_1567);
or U2594 (N_2594,N_1901,N_2063);
or U2595 (N_2595,N_1752,N_1849);
or U2596 (N_2596,N_1880,N_2193);
nand U2597 (N_2597,N_1948,N_2138);
or U2598 (N_2598,N_2110,N_1584);
or U2599 (N_2599,N_2211,N_1767);
and U2600 (N_2600,N_1748,N_1853);
and U2601 (N_2601,N_2054,N_2095);
and U2602 (N_2602,N_2096,N_2189);
nor U2603 (N_2603,N_1786,N_1685);
nor U2604 (N_2604,N_1619,N_2173);
nand U2605 (N_2605,N_1574,N_1676);
nor U2606 (N_2606,N_1637,N_1902);
or U2607 (N_2607,N_2194,N_1510);
nand U2608 (N_2608,N_1878,N_1618);
or U2609 (N_2609,N_2043,N_1632);
xnor U2610 (N_2610,N_1813,N_1743);
nand U2611 (N_2611,N_2171,N_2083);
nand U2612 (N_2612,N_1763,N_1703);
nand U2613 (N_2613,N_1886,N_2241);
and U2614 (N_2614,N_1772,N_2236);
nand U2615 (N_2615,N_1593,N_1582);
or U2616 (N_2616,N_1794,N_2067);
and U2617 (N_2617,N_2199,N_2186);
nand U2618 (N_2618,N_1643,N_2248);
nand U2619 (N_2619,N_1962,N_2221);
or U2620 (N_2620,N_1722,N_1540);
or U2621 (N_2621,N_2220,N_1882);
and U2622 (N_2622,N_1509,N_2085);
nand U2623 (N_2623,N_2164,N_1683);
xor U2624 (N_2624,N_1931,N_1788);
nand U2625 (N_2625,N_1651,N_1704);
nor U2626 (N_2626,N_1872,N_1888);
and U2627 (N_2627,N_2247,N_2239);
nor U2628 (N_2628,N_2083,N_2075);
or U2629 (N_2629,N_1630,N_1584);
and U2630 (N_2630,N_2127,N_2182);
and U2631 (N_2631,N_2095,N_2028);
or U2632 (N_2632,N_2167,N_1809);
nand U2633 (N_2633,N_2172,N_1978);
nand U2634 (N_2634,N_1982,N_2070);
nand U2635 (N_2635,N_1805,N_1647);
or U2636 (N_2636,N_2053,N_1966);
or U2637 (N_2637,N_2101,N_2140);
or U2638 (N_2638,N_1804,N_1975);
and U2639 (N_2639,N_2076,N_1522);
nand U2640 (N_2640,N_1710,N_1633);
nor U2641 (N_2641,N_2032,N_2062);
and U2642 (N_2642,N_1935,N_2038);
and U2643 (N_2643,N_2076,N_1762);
nand U2644 (N_2644,N_2196,N_1646);
and U2645 (N_2645,N_2176,N_2069);
nor U2646 (N_2646,N_2246,N_1517);
or U2647 (N_2647,N_2180,N_2104);
nor U2648 (N_2648,N_2133,N_1790);
nand U2649 (N_2649,N_1889,N_1760);
and U2650 (N_2650,N_2149,N_1540);
or U2651 (N_2651,N_1502,N_2118);
or U2652 (N_2652,N_1692,N_1690);
xor U2653 (N_2653,N_2098,N_1823);
nand U2654 (N_2654,N_1751,N_2139);
nand U2655 (N_2655,N_1757,N_1642);
nor U2656 (N_2656,N_1850,N_1797);
xor U2657 (N_2657,N_2084,N_1743);
nor U2658 (N_2658,N_1668,N_1816);
nand U2659 (N_2659,N_1873,N_1665);
nor U2660 (N_2660,N_1978,N_2126);
and U2661 (N_2661,N_1805,N_2241);
and U2662 (N_2662,N_1640,N_2102);
or U2663 (N_2663,N_1835,N_1535);
nand U2664 (N_2664,N_1900,N_1903);
or U2665 (N_2665,N_2158,N_1737);
nand U2666 (N_2666,N_2000,N_1789);
and U2667 (N_2667,N_1673,N_2010);
nand U2668 (N_2668,N_1537,N_1824);
or U2669 (N_2669,N_1856,N_1508);
or U2670 (N_2670,N_1695,N_1986);
and U2671 (N_2671,N_1533,N_1689);
nor U2672 (N_2672,N_2244,N_1800);
and U2673 (N_2673,N_1632,N_1750);
and U2674 (N_2674,N_1694,N_1612);
nand U2675 (N_2675,N_1640,N_2124);
or U2676 (N_2676,N_2146,N_1896);
and U2677 (N_2677,N_2108,N_2093);
or U2678 (N_2678,N_1843,N_2237);
and U2679 (N_2679,N_1973,N_1902);
and U2680 (N_2680,N_1727,N_2022);
nor U2681 (N_2681,N_1622,N_2196);
nor U2682 (N_2682,N_1517,N_1710);
or U2683 (N_2683,N_1546,N_2122);
or U2684 (N_2684,N_2084,N_1565);
nand U2685 (N_2685,N_1802,N_1794);
nand U2686 (N_2686,N_2161,N_1808);
or U2687 (N_2687,N_1757,N_2095);
and U2688 (N_2688,N_1835,N_1586);
and U2689 (N_2689,N_1816,N_1865);
and U2690 (N_2690,N_1932,N_1877);
and U2691 (N_2691,N_2151,N_1817);
nand U2692 (N_2692,N_1962,N_2143);
nand U2693 (N_2693,N_1732,N_2173);
and U2694 (N_2694,N_1539,N_1655);
nand U2695 (N_2695,N_1861,N_2029);
or U2696 (N_2696,N_2072,N_2079);
and U2697 (N_2697,N_2054,N_1683);
or U2698 (N_2698,N_1864,N_1844);
and U2699 (N_2699,N_2223,N_1761);
and U2700 (N_2700,N_1612,N_1906);
nor U2701 (N_2701,N_1989,N_1888);
nor U2702 (N_2702,N_1815,N_1898);
nand U2703 (N_2703,N_2080,N_1593);
nor U2704 (N_2704,N_1698,N_2046);
and U2705 (N_2705,N_1976,N_1535);
nand U2706 (N_2706,N_2138,N_2000);
or U2707 (N_2707,N_1972,N_1891);
and U2708 (N_2708,N_2226,N_1666);
or U2709 (N_2709,N_1939,N_2072);
or U2710 (N_2710,N_1924,N_1599);
nor U2711 (N_2711,N_1836,N_2066);
xor U2712 (N_2712,N_1524,N_2181);
nor U2713 (N_2713,N_1697,N_1898);
nor U2714 (N_2714,N_2208,N_1551);
or U2715 (N_2715,N_1565,N_1550);
and U2716 (N_2716,N_2102,N_2207);
and U2717 (N_2717,N_1816,N_1995);
nand U2718 (N_2718,N_2094,N_2195);
nand U2719 (N_2719,N_1925,N_2103);
nor U2720 (N_2720,N_2146,N_1964);
or U2721 (N_2721,N_1716,N_1930);
nand U2722 (N_2722,N_1955,N_2068);
and U2723 (N_2723,N_1664,N_1890);
xnor U2724 (N_2724,N_2014,N_1544);
or U2725 (N_2725,N_1782,N_1628);
or U2726 (N_2726,N_1683,N_1721);
and U2727 (N_2727,N_1955,N_1630);
nor U2728 (N_2728,N_1701,N_2190);
nand U2729 (N_2729,N_1823,N_1860);
nor U2730 (N_2730,N_1926,N_1704);
and U2731 (N_2731,N_2073,N_2216);
or U2732 (N_2732,N_1503,N_1504);
and U2733 (N_2733,N_1971,N_1540);
nand U2734 (N_2734,N_1594,N_1937);
or U2735 (N_2735,N_1933,N_1932);
nand U2736 (N_2736,N_1650,N_2120);
nor U2737 (N_2737,N_1954,N_1779);
nand U2738 (N_2738,N_1659,N_1886);
nand U2739 (N_2739,N_2033,N_2217);
nand U2740 (N_2740,N_1536,N_1822);
and U2741 (N_2741,N_1919,N_2069);
and U2742 (N_2742,N_1681,N_1769);
nor U2743 (N_2743,N_1610,N_1579);
or U2744 (N_2744,N_2056,N_1500);
nor U2745 (N_2745,N_2217,N_1518);
or U2746 (N_2746,N_1847,N_2220);
and U2747 (N_2747,N_2089,N_1564);
and U2748 (N_2748,N_2196,N_1518);
nand U2749 (N_2749,N_1934,N_2129);
or U2750 (N_2750,N_1949,N_1786);
nand U2751 (N_2751,N_1557,N_1773);
or U2752 (N_2752,N_2088,N_2073);
or U2753 (N_2753,N_1889,N_1900);
nand U2754 (N_2754,N_1603,N_2021);
and U2755 (N_2755,N_1638,N_2085);
or U2756 (N_2756,N_2213,N_1689);
or U2757 (N_2757,N_1515,N_1529);
and U2758 (N_2758,N_1848,N_2121);
nand U2759 (N_2759,N_2246,N_1530);
and U2760 (N_2760,N_2116,N_1740);
and U2761 (N_2761,N_1891,N_1502);
nor U2762 (N_2762,N_2166,N_2115);
nor U2763 (N_2763,N_1915,N_1598);
and U2764 (N_2764,N_1558,N_1539);
nor U2765 (N_2765,N_1763,N_1722);
nand U2766 (N_2766,N_2216,N_1679);
or U2767 (N_2767,N_1789,N_2174);
nor U2768 (N_2768,N_2010,N_2146);
and U2769 (N_2769,N_1959,N_1736);
or U2770 (N_2770,N_1777,N_1585);
nand U2771 (N_2771,N_1900,N_1651);
nand U2772 (N_2772,N_2040,N_2038);
or U2773 (N_2773,N_1841,N_2217);
or U2774 (N_2774,N_1538,N_1926);
nor U2775 (N_2775,N_1733,N_1798);
or U2776 (N_2776,N_1633,N_1978);
nand U2777 (N_2777,N_2003,N_1815);
nand U2778 (N_2778,N_2157,N_2103);
or U2779 (N_2779,N_2165,N_1766);
or U2780 (N_2780,N_1710,N_1777);
nor U2781 (N_2781,N_1502,N_1917);
nand U2782 (N_2782,N_1618,N_1515);
and U2783 (N_2783,N_2163,N_1792);
nand U2784 (N_2784,N_2047,N_1623);
nor U2785 (N_2785,N_1985,N_2108);
or U2786 (N_2786,N_2226,N_2038);
or U2787 (N_2787,N_2148,N_1645);
xor U2788 (N_2788,N_1506,N_1730);
nor U2789 (N_2789,N_1529,N_2026);
and U2790 (N_2790,N_1665,N_2144);
xnor U2791 (N_2791,N_1784,N_1617);
and U2792 (N_2792,N_1675,N_2167);
and U2793 (N_2793,N_1610,N_1675);
nand U2794 (N_2794,N_1845,N_1844);
or U2795 (N_2795,N_1747,N_1662);
and U2796 (N_2796,N_2145,N_1917);
nand U2797 (N_2797,N_2030,N_1808);
and U2798 (N_2798,N_1726,N_2143);
nor U2799 (N_2799,N_1872,N_1918);
xnor U2800 (N_2800,N_1955,N_2071);
and U2801 (N_2801,N_1602,N_1936);
nor U2802 (N_2802,N_1809,N_2099);
and U2803 (N_2803,N_1783,N_1641);
or U2804 (N_2804,N_1846,N_1997);
nor U2805 (N_2805,N_1748,N_2032);
and U2806 (N_2806,N_2069,N_1701);
nand U2807 (N_2807,N_1743,N_1662);
nand U2808 (N_2808,N_2065,N_2210);
xnor U2809 (N_2809,N_2055,N_1775);
or U2810 (N_2810,N_1517,N_1883);
or U2811 (N_2811,N_1900,N_1577);
or U2812 (N_2812,N_1976,N_2140);
and U2813 (N_2813,N_1909,N_2232);
and U2814 (N_2814,N_1794,N_2087);
and U2815 (N_2815,N_2207,N_1907);
or U2816 (N_2816,N_1631,N_2082);
nor U2817 (N_2817,N_1593,N_2182);
nand U2818 (N_2818,N_1773,N_1971);
nand U2819 (N_2819,N_1526,N_2017);
nor U2820 (N_2820,N_1757,N_1917);
and U2821 (N_2821,N_1535,N_2213);
nand U2822 (N_2822,N_1886,N_2061);
and U2823 (N_2823,N_1728,N_1574);
nand U2824 (N_2824,N_1703,N_1797);
nor U2825 (N_2825,N_2242,N_2181);
nor U2826 (N_2826,N_1920,N_1727);
nand U2827 (N_2827,N_2181,N_1764);
and U2828 (N_2828,N_2117,N_1716);
or U2829 (N_2829,N_1816,N_1777);
nor U2830 (N_2830,N_1758,N_1787);
or U2831 (N_2831,N_1565,N_1543);
nand U2832 (N_2832,N_2078,N_1522);
nor U2833 (N_2833,N_2036,N_1884);
and U2834 (N_2834,N_1670,N_1946);
or U2835 (N_2835,N_1848,N_2061);
nor U2836 (N_2836,N_2151,N_2028);
and U2837 (N_2837,N_2241,N_2215);
and U2838 (N_2838,N_1950,N_2187);
and U2839 (N_2839,N_1900,N_1927);
and U2840 (N_2840,N_1694,N_2039);
nand U2841 (N_2841,N_1926,N_1561);
nor U2842 (N_2842,N_2212,N_1605);
or U2843 (N_2843,N_2124,N_1911);
and U2844 (N_2844,N_1746,N_2163);
and U2845 (N_2845,N_1538,N_1772);
or U2846 (N_2846,N_1705,N_1533);
or U2847 (N_2847,N_1636,N_1780);
nand U2848 (N_2848,N_1886,N_2183);
nor U2849 (N_2849,N_2114,N_2182);
and U2850 (N_2850,N_2191,N_2246);
or U2851 (N_2851,N_1838,N_1940);
and U2852 (N_2852,N_1527,N_1862);
nor U2853 (N_2853,N_1522,N_2028);
nand U2854 (N_2854,N_2208,N_2164);
nor U2855 (N_2855,N_1784,N_1955);
and U2856 (N_2856,N_1822,N_1915);
nor U2857 (N_2857,N_1690,N_1585);
or U2858 (N_2858,N_1887,N_1582);
nand U2859 (N_2859,N_1866,N_1554);
or U2860 (N_2860,N_1956,N_1791);
and U2861 (N_2861,N_1843,N_1770);
nand U2862 (N_2862,N_1788,N_1713);
or U2863 (N_2863,N_1744,N_1950);
or U2864 (N_2864,N_2143,N_1680);
xnor U2865 (N_2865,N_2183,N_1906);
nor U2866 (N_2866,N_1889,N_2165);
and U2867 (N_2867,N_1616,N_1667);
nand U2868 (N_2868,N_2156,N_1945);
or U2869 (N_2869,N_2189,N_2154);
nor U2870 (N_2870,N_1958,N_1691);
or U2871 (N_2871,N_2192,N_1570);
nand U2872 (N_2872,N_1667,N_1822);
nand U2873 (N_2873,N_1937,N_2125);
or U2874 (N_2874,N_1927,N_1781);
nor U2875 (N_2875,N_2247,N_1763);
nor U2876 (N_2876,N_1903,N_1787);
nor U2877 (N_2877,N_1620,N_1693);
nor U2878 (N_2878,N_1705,N_2199);
or U2879 (N_2879,N_1729,N_2166);
nand U2880 (N_2880,N_1768,N_2236);
or U2881 (N_2881,N_2210,N_1666);
xor U2882 (N_2882,N_2238,N_1980);
nand U2883 (N_2883,N_1906,N_2076);
nor U2884 (N_2884,N_2006,N_1815);
or U2885 (N_2885,N_1811,N_2241);
nand U2886 (N_2886,N_2027,N_2029);
xor U2887 (N_2887,N_2224,N_1965);
nand U2888 (N_2888,N_1866,N_1567);
xnor U2889 (N_2889,N_2148,N_1585);
nor U2890 (N_2890,N_2246,N_1956);
nor U2891 (N_2891,N_2091,N_1850);
nand U2892 (N_2892,N_1877,N_1639);
nor U2893 (N_2893,N_2019,N_2094);
and U2894 (N_2894,N_1837,N_1835);
and U2895 (N_2895,N_2221,N_1607);
or U2896 (N_2896,N_1834,N_1537);
nand U2897 (N_2897,N_1505,N_1893);
or U2898 (N_2898,N_1871,N_1512);
xnor U2899 (N_2899,N_1981,N_1833);
nand U2900 (N_2900,N_1999,N_2106);
or U2901 (N_2901,N_1774,N_1570);
and U2902 (N_2902,N_1921,N_1513);
or U2903 (N_2903,N_1719,N_2002);
nor U2904 (N_2904,N_1800,N_2032);
and U2905 (N_2905,N_2130,N_2063);
nand U2906 (N_2906,N_2158,N_2134);
nand U2907 (N_2907,N_1947,N_1744);
xor U2908 (N_2908,N_2127,N_1757);
and U2909 (N_2909,N_2035,N_1586);
and U2910 (N_2910,N_2194,N_1948);
nand U2911 (N_2911,N_1637,N_1692);
nand U2912 (N_2912,N_1632,N_2127);
and U2913 (N_2913,N_2158,N_1880);
nand U2914 (N_2914,N_1556,N_1942);
nand U2915 (N_2915,N_1695,N_1853);
and U2916 (N_2916,N_1904,N_1960);
and U2917 (N_2917,N_2154,N_1830);
nand U2918 (N_2918,N_1705,N_2113);
nor U2919 (N_2919,N_1991,N_1936);
nor U2920 (N_2920,N_1770,N_2101);
and U2921 (N_2921,N_1787,N_1743);
or U2922 (N_2922,N_1507,N_1921);
or U2923 (N_2923,N_2224,N_1876);
nor U2924 (N_2924,N_1524,N_1575);
and U2925 (N_2925,N_1736,N_1980);
nand U2926 (N_2926,N_2147,N_2091);
xor U2927 (N_2927,N_1951,N_1952);
and U2928 (N_2928,N_2024,N_1902);
and U2929 (N_2929,N_2118,N_1727);
or U2930 (N_2930,N_2168,N_1640);
and U2931 (N_2931,N_2106,N_1635);
or U2932 (N_2932,N_2132,N_1848);
or U2933 (N_2933,N_1607,N_1879);
nor U2934 (N_2934,N_1993,N_1639);
nor U2935 (N_2935,N_1660,N_2026);
nor U2936 (N_2936,N_1665,N_1786);
and U2937 (N_2937,N_1963,N_2117);
or U2938 (N_2938,N_2142,N_2064);
or U2939 (N_2939,N_2092,N_1722);
and U2940 (N_2940,N_1912,N_1770);
nand U2941 (N_2941,N_1846,N_2147);
nand U2942 (N_2942,N_2084,N_1846);
nand U2943 (N_2943,N_2159,N_1659);
and U2944 (N_2944,N_1865,N_1567);
and U2945 (N_2945,N_2130,N_1677);
or U2946 (N_2946,N_2104,N_1549);
or U2947 (N_2947,N_1847,N_1875);
nor U2948 (N_2948,N_1906,N_1778);
or U2949 (N_2949,N_1972,N_1606);
nor U2950 (N_2950,N_2103,N_2180);
nor U2951 (N_2951,N_1505,N_1929);
xor U2952 (N_2952,N_1571,N_1838);
nand U2953 (N_2953,N_1928,N_2040);
nand U2954 (N_2954,N_1875,N_2216);
and U2955 (N_2955,N_1995,N_2028);
and U2956 (N_2956,N_1682,N_2025);
and U2957 (N_2957,N_2072,N_1638);
or U2958 (N_2958,N_1593,N_2044);
and U2959 (N_2959,N_1611,N_2155);
and U2960 (N_2960,N_1765,N_1685);
and U2961 (N_2961,N_1633,N_2062);
nand U2962 (N_2962,N_2131,N_1676);
or U2963 (N_2963,N_1635,N_2149);
or U2964 (N_2964,N_1579,N_2195);
and U2965 (N_2965,N_2248,N_1991);
or U2966 (N_2966,N_2104,N_1637);
or U2967 (N_2967,N_1639,N_1587);
nor U2968 (N_2968,N_1982,N_2024);
nand U2969 (N_2969,N_1743,N_2214);
and U2970 (N_2970,N_1959,N_1861);
or U2971 (N_2971,N_1503,N_1519);
nand U2972 (N_2972,N_2086,N_2241);
nor U2973 (N_2973,N_1966,N_2018);
and U2974 (N_2974,N_1701,N_2211);
and U2975 (N_2975,N_2245,N_1834);
nor U2976 (N_2976,N_1694,N_2004);
nand U2977 (N_2977,N_2168,N_1642);
nor U2978 (N_2978,N_1560,N_1757);
nor U2979 (N_2979,N_2156,N_1891);
nand U2980 (N_2980,N_1505,N_1967);
and U2981 (N_2981,N_2185,N_2003);
and U2982 (N_2982,N_1613,N_1944);
nand U2983 (N_2983,N_2248,N_2090);
nor U2984 (N_2984,N_1699,N_1766);
and U2985 (N_2985,N_2107,N_1631);
nand U2986 (N_2986,N_1521,N_2100);
or U2987 (N_2987,N_1940,N_2188);
xor U2988 (N_2988,N_2041,N_1655);
or U2989 (N_2989,N_1597,N_1836);
or U2990 (N_2990,N_1869,N_1905);
and U2991 (N_2991,N_1546,N_2032);
and U2992 (N_2992,N_1925,N_1570);
nor U2993 (N_2993,N_1910,N_1650);
nand U2994 (N_2994,N_1918,N_1621);
and U2995 (N_2995,N_2107,N_2150);
nor U2996 (N_2996,N_2239,N_1764);
nor U2997 (N_2997,N_1599,N_1563);
nor U2998 (N_2998,N_2224,N_1620);
nor U2999 (N_2999,N_2063,N_1840);
or UO_0 (O_0,N_2994,N_2382);
nor UO_1 (O_1,N_2344,N_2761);
and UO_2 (O_2,N_2998,N_2966);
and UO_3 (O_3,N_2885,N_2693);
or UO_4 (O_4,N_2427,N_2339);
nor UO_5 (O_5,N_2640,N_2263);
nor UO_6 (O_6,N_2773,N_2408);
or UO_7 (O_7,N_2791,N_2293);
nand UO_8 (O_8,N_2462,N_2380);
nor UO_9 (O_9,N_2748,N_2886);
or UO_10 (O_10,N_2637,N_2785);
nand UO_11 (O_11,N_2357,N_2682);
nand UO_12 (O_12,N_2337,N_2486);
nand UO_13 (O_13,N_2262,N_2812);
nand UO_14 (O_14,N_2475,N_2655);
or UO_15 (O_15,N_2833,N_2881);
nor UO_16 (O_16,N_2561,N_2618);
nor UO_17 (O_17,N_2976,N_2803);
or UO_18 (O_18,N_2775,N_2711);
and UO_19 (O_19,N_2511,N_2872);
nand UO_20 (O_20,N_2258,N_2741);
nor UO_21 (O_21,N_2632,N_2859);
or UO_22 (O_22,N_2744,N_2534);
nand UO_23 (O_23,N_2954,N_2445);
or UO_24 (O_24,N_2948,N_2464);
or UO_25 (O_25,N_2863,N_2592);
or UO_26 (O_26,N_2436,N_2362);
nor UO_27 (O_27,N_2712,N_2288);
and UO_28 (O_28,N_2788,N_2495);
nor UO_29 (O_29,N_2671,N_2440);
nand UO_30 (O_30,N_2919,N_2694);
or UO_31 (O_31,N_2574,N_2950);
and UO_32 (O_32,N_2937,N_2576);
nand UO_33 (O_33,N_2825,N_2801);
nor UO_34 (O_34,N_2457,N_2975);
or UO_35 (O_35,N_2727,N_2672);
and UO_36 (O_36,N_2333,N_2666);
or UO_37 (O_37,N_2454,N_2680);
or UO_38 (O_38,N_2366,N_2361);
nor UO_39 (O_39,N_2995,N_2928);
and UO_40 (O_40,N_2422,N_2984);
nand UO_41 (O_41,N_2310,N_2912);
nand UO_42 (O_42,N_2709,N_2997);
or UO_43 (O_43,N_2484,N_2721);
and UO_44 (O_44,N_2944,N_2932);
and UO_45 (O_45,N_2483,N_2926);
nor UO_46 (O_46,N_2815,N_2392);
nand UO_47 (O_47,N_2813,N_2479);
or UO_48 (O_48,N_2619,N_2733);
or UO_49 (O_49,N_2804,N_2720);
nor UO_50 (O_50,N_2816,N_2419);
nor UO_51 (O_51,N_2633,N_2875);
or UO_52 (O_52,N_2496,N_2598);
and UO_53 (O_53,N_2424,N_2498);
nor UO_54 (O_54,N_2573,N_2516);
and UO_55 (O_55,N_2299,N_2747);
and UO_56 (O_56,N_2571,N_2442);
or UO_57 (O_57,N_2809,N_2360);
nor UO_58 (O_58,N_2849,N_2965);
and UO_59 (O_59,N_2691,N_2522);
or UO_60 (O_60,N_2379,N_2983);
or UO_61 (O_61,N_2669,N_2609);
nand UO_62 (O_62,N_2867,N_2629);
nand UO_63 (O_63,N_2430,N_2343);
nand UO_64 (O_64,N_2848,N_2331);
nand UO_65 (O_65,N_2557,N_2289);
nor UO_66 (O_66,N_2459,N_2934);
nand UO_67 (O_67,N_2663,N_2644);
nand UO_68 (O_68,N_2473,N_2951);
nand UO_69 (O_69,N_2900,N_2891);
or UO_70 (O_70,N_2477,N_2326);
nand UO_71 (O_71,N_2638,N_2329);
nor UO_72 (O_72,N_2448,N_2665);
nand UO_73 (O_73,N_2469,N_2961);
nor UO_74 (O_74,N_2404,N_2435);
or UO_75 (O_75,N_2981,N_2986);
nor UO_76 (O_76,N_2282,N_2458);
or UO_77 (O_77,N_2355,N_2611);
and UO_78 (O_78,N_2957,N_2896);
nand UO_79 (O_79,N_2898,N_2792);
or UO_80 (O_80,N_2878,N_2635);
or UO_81 (O_81,N_2562,N_2670);
or UO_82 (O_82,N_2295,N_2531);
nand UO_83 (O_83,N_2649,N_2700);
or UO_84 (O_84,N_2342,N_2614);
nand UO_85 (O_85,N_2880,N_2252);
and UO_86 (O_86,N_2385,N_2940);
nand UO_87 (O_87,N_2397,N_2659);
and UO_88 (O_88,N_2735,N_2330);
and UO_89 (O_89,N_2676,N_2309);
nand UO_90 (O_90,N_2656,N_2608);
nand UO_91 (O_91,N_2746,N_2681);
and UO_92 (O_92,N_2322,N_2641);
nor UO_93 (O_93,N_2363,N_2300);
and UO_94 (O_94,N_2958,N_2873);
and UO_95 (O_95,N_2500,N_2536);
nor UO_96 (O_96,N_2959,N_2567);
or UO_97 (O_97,N_2839,N_2643);
nor UO_98 (O_98,N_2956,N_2802);
and UO_99 (O_99,N_2368,N_2850);
nor UO_100 (O_100,N_2999,N_2527);
nor UO_101 (O_101,N_2814,N_2585);
and UO_102 (O_102,N_2841,N_2714);
and UO_103 (O_103,N_2526,N_2367);
or UO_104 (O_104,N_2346,N_2506);
or UO_105 (O_105,N_2616,N_2979);
nor UO_106 (O_106,N_2525,N_2742);
nand UO_107 (O_107,N_2858,N_2467);
and UO_108 (O_108,N_2701,N_2311);
nand UO_109 (O_109,N_2423,N_2854);
nand UO_110 (O_110,N_2468,N_2821);
nor UO_111 (O_111,N_2556,N_2524);
nand UO_112 (O_112,N_2799,N_2726);
nor UO_113 (O_113,N_2780,N_2400);
and UO_114 (O_114,N_2829,N_2630);
nand UO_115 (O_115,N_2260,N_2847);
and UO_116 (O_116,N_2540,N_2504);
and UO_117 (O_117,N_2612,N_2996);
and UO_118 (O_118,N_2989,N_2936);
or UO_119 (O_119,N_2364,N_2767);
and UO_120 (O_120,N_2731,N_2493);
nor UO_121 (O_121,N_2869,N_2931);
or UO_122 (O_122,N_2280,N_2877);
xnor UO_123 (O_123,N_2800,N_2783);
and UO_124 (O_124,N_2543,N_2861);
nand UO_125 (O_125,N_2551,N_2924);
nand UO_126 (O_126,N_2383,N_2320);
and UO_127 (O_127,N_2480,N_2340);
nor UO_128 (O_128,N_2521,N_2563);
xor UO_129 (O_129,N_2617,N_2301);
xor UO_130 (O_130,N_2365,N_2284);
and UO_131 (O_131,N_2316,N_2272);
or UO_132 (O_132,N_2762,N_2276);
or UO_133 (O_133,N_2621,N_2673);
nand UO_134 (O_134,N_2921,N_2358);
or UO_135 (O_135,N_2769,N_2895);
nand UO_136 (O_136,N_2856,N_2377);
and UO_137 (O_137,N_2929,N_2606);
nor UO_138 (O_138,N_2824,N_2810);
or UO_139 (O_139,N_2302,N_2411);
or UO_140 (O_140,N_2933,N_2840);
or UO_141 (O_141,N_2993,N_2667);
nor UO_142 (O_142,N_2760,N_2723);
nand UO_143 (O_143,N_2758,N_2403);
nand UO_144 (O_144,N_2980,N_2507);
nand UO_145 (O_145,N_2582,N_2662);
nor UO_146 (O_146,N_2437,N_2446);
nor UO_147 (O_147,N_2465,N_2555);
nor UO_148 (O_148,N_2345,N_2610);
nand UO_149 (O_149,N_2314,N_2390);
nand UO_150 (O_150,N_2864,N_2580);
and UO_151 (O_151,N_2434,N_2413);
and UO_152 (O_152,N_2432,N_2577);
nand UO_153 (O_153,N_2894,N_2753);
or UO_154 (O_154,N_2418,N_2313);
nor UO_155 (O_155,N_2620,N_2901);
nor UO_156 (O_156,N_2373,N_2692);
and UO_157 (O_157,N_2297,N_2509);
nand UO_158 (O_158,N_2318,N_2636);
and UO_159 (O_159,N_2624,N_2646);
nand UO_160 (O_160,N_2660,N_2684);
and UO_161 (O_161,N_2336,N_2306);
nor UO_162 (O_162,N_2421,N_2907);
and UO_163 (O_163,N_2399,N_2319);
nor UO_164 (O_164,N_2857,N_2830);
and UO_165 (O_165,N_2974,N_2739);
nand UO_166 (O_166,N_2751,N_2826);
or UO_167 (O_167,N_2517,N_2533);
or UO_168 (O_168,N_2528,N_2952);
or UO_169 (O_169,N_2910,N_2560);
and UO_170 (O_170,N_2978,N_2414);
nor UO_171 (O_171,N_2845,N_2906);
nand UO_172 (O_172,N_2552,N_2888);
xor UO_173 (O_173,N_2564,N_2838);
nor UO_174 (O_174,N_2962,N_2372);
nor UO_175 (O_175,N_2729,N_2391);
nand UO_176 (O_176,N_2687,N_2793);
and UO_177 (O_177,N_2764,N_2967);
and UO_178 (O_178,N_2899,N_2325);
and UO_179 (O_179,N_2494,N_2291);
and UO_180 (O_180,N_2811,N_2501);
xnor UO_181 (O_181,N_2294,N_2622);
nor UO_182 (O_182,N_2927,N_2505);
or UO_183 (O_183,N_2451,N_2730);
nor UO_184 (O_184,N_2359,N_2777);
or UO_185 (O_185,N_2642,N_2818);
nand UO_186 (O_186,N_2625,N_2913);
nand UO_187 (O_187,N_2930,N_2759);
and UO_188 (O_188,N_2982,N_2879);
or UO_189 (O_189,N_2710,N_2425);
nand UO_190 (O_190,N_2771,N_2724);
or UO_191 (O_191,N_2737,N_2568);
nand UO_192 (O_192,N_2757,N_2782);
and UO_193 (O_193,N_2449,N_2450);
or UO_194 (O_194,N_2514,N_2503);
or UO_195 (O_195,N_2416,N_2853);
nand UO_196 (O_196,N_2271,N_2969);
nor UO_197 (O_197,N_2914,N_2335);
or UO_198 (O_198,N_2287,N_2513);
or UO_199 (O_199,N_2615,N_2381);
nor UO_200 (O_200,N_2588,N_2452);
nand UO_201 (O_201,N_2596,N_2876);
and UO_202 (O_202,N_2705,N_2808);
nor UO_203 (O_203,N_2402,N_2535);
nor UO_204 (O_204,N_2554,N_2668);
nand UO_205 (O_205,N_2756,N_2796);
nand UO_206 (O_206,N_2321,N_2797);
or UO_207 (O_207,N_2485,N_2652);
and UO_208 (O_208,N_2508,N_2843);
nand UO_209 (O_209,N_2324,N_2407);
or UO_210 (O_210,N_2253,N_2805);
or UO_211 (O_211,N_2920,N_2547);
nand UO_212 (O_212,N_2902,N_2860);
nor UO_213 (O_213,N_2904,N_2332);
nor UO_214 (O_214,N_2781,N_2654);
nor UO_215 (O_215,N_2281,N_2790);
or UO_216 (O_216,N_2278,N_2953);
or UO_217 (O_217,N_2752,N_2916);
or UO_218 (O_218,N_2369,N_2743);
nor UO_219 (O_219,N_2977,N_2678);
and UO_220 (O_220,N_2828,N_2698);
and UO_221 (O_221,N_2417,N_2677);
xor UO_222 (O_222,N_2827,N_2255);
nand UO_223 (O_223,N_2570,N_2817);
and UO_224 (O_224,N_2254,N_2600);
or UO_225 (O_225,N_2602,N_2945);
and UO_226 (O_226,N_2831,N_2572);
nor UO_227 (O_227,N_2715,N_2594);
nand UO_228 (O_228,N_2890,N_2823);
and UO_229 (O_229,N_2482,N_2273);
or UO_230 (O_230,N_2707,N_2444);
nor UO_231 (O_231,N_2703,N_2658);
and UO_232 (O_232,N_2541,N_2639);
nand UO_233 (O_233,N_2664,N_2972);
or UO_234 (O_234,N_2789,N_2530);
nand UO_235 (O_235,N_2779,N_2607);
nor UO_236 (O_236,N_2889,N_2334);
and UO_237 (O_237,N_2702,N_2749);
nand UO_238 (O_238,N_2648,N_2470);
and UO_239 (O_239,N_2460,N_2647);
and UO_240 (O_240,N_2942,N_2341);
nor UO_241 (O_241,N_2695,N_2441);
nand UO_242 (O_242,N_2601,N_2296);
nor UO_243 (O_243,N_2893,N_2431);
and UO_244 (O_244,N_2312,N_2732);
and UO_245 (O_245,N_2415,N_2717);
nand UO_246 (O_246,N_2566,N_2939);
or UO_247 (O_247,N_2964,N_2292);
and UO_248 (O_248,N_2915,N_2683);
or UO_249 (O_249,N_2846,N_2250);
nor UO_250 (O_250,N_2461,N_2489);
nor UO_251 (O_251,N_2519,N_2267);
nor UO_252 (O_252,N_2887,N_2388);
and UO_253 (O_253,N_2699,N_2290);
or UO_254 (O_254,N_2949,N_2581);
nor UO_255 (O_255,N_2386,N_2591);
and UO_256 (O_256,N_2439,N_2532);
nor UO_257 (O_257,N_2370,N_2786);
nand UO_258 (O_258,N_2488,N_2947);
and UO_259 (O_259,N_2943,N_2822);
nor UO_260 (O_260,N_2593,N_2587);
nor UO_261 (O_261,N_2351,N_2453);
nor UO_262 (O_262,N_2918,N_2628);
and UO_263 (O_263,N_2661,N_2938);
nor UO_264 (O_264,N_2935,N_2472);
and UO_265 (O_265,N_2569,N_2352);
and UO_266 (O_266,N_2371,N_2499);
nor UO_267 (O_267,N_2599,N_2807);
nor UO_268 (O_268,N_2868,N_2870);
nand UO_269 (O_269,N_2991,N_2298);
and UO_270 (O_270,N_2548,N_2836);
and UO_271 (O_271,N_2478,N_2565);
and UO_272 (O_272,N_2882,N_2884);
nor UO_273 (O_273,N_2990,N_2597);
xor UO_274 (O_274,N_2406,N_2401);
nor UO_275 (O_275,N_2754,N_2679);
or UO_276 (O_276,N_2674,N_2277);
or UO_277 (O_277,N_2466,N_2835);
nor UO_278 (O_278,N_2350,N_2409);
xor UO_279 (O_279,N_2428,N_2963);
and UO_280 (O_280,N_2871,N_2968);
or UO_281 (O_281,N_2396,N_2257);
and UO_282 (O_282,N_2523,N_2347);
or UO_283 (O_283,N_2897,N_2819);
nor UO_284 (O_284,N_2529,N_2398);
nand UO_285 (O_285,N_2605,N_2837);
or UO_286 (O_286,N_2268,N_2286);
or UO_287 (O_287,N_2559,N_2708);
or UO_288 (O_288,N_2631,N_2410);
and UO_289 (O_289,N_2704,N_2375);
nand UO_290 (O_290,N_2349,N_2553);
nand UO_291 (O_291,N_2586,N_2706);
nor UO_292 (O_292,N_2946,N_2269);
or UO_293 (O_293,N_2653,N_2766);
or UO_294 (O_294,N_2697,N_2327);
nand UO_295 (O_295,N_2909,N_2718);
nand UO_296 (O_296,N_2987,N_2538);
nor UO_297 (O_297,N_2539,N_2520);
or UO_298 (O_298,N_2865,N_2356);
or UO_299 (O_299,N_2719,N_2738);
nor UO_300 (O_300,N_2675,N_2925);
and UO_301 (O_301,N_2443,N_2774);
and UO_302 (O_302,N_2578,N_2626);
and UO_303 (O_303,N_2988,N_2971);
and UO_304 (O_304,N_2651,N_2455);
or UO_305 (O_305,N_2323,N_2716);
nor UO_306 (O_306,N_2405,N_2303);
and UO_307 (O_307,N_2420,N_2512);
nand UO_308 (O_308,N_2795,N_2892);
nor UO_309 (O_309,N_2256,N_2645);
and UO_310 (O_310,N_2595,N_2376);
nand UO_311 (O_311,N_2394,N_2784);
nor UO_312 (O_312,N_2627,N_2515);
or UO_313 (O_313,N_2456,N_2787);
nor UO_314 (O_314,N_2542,N_2842);
nand UO_315 (O_315,N_2603,N_2412);
or UO_316 (O_316,N_2604,N_2471);
and UO_317 (O_317,N_2686,N_2820);
or UO_318 (O_318,N_2261,N_2941);
or UO_319 (O_319,N_2763,N_2279);
nand UO_320 (O_320,N_2696,N_2905);
or UO_321 (O_321,N_2270,N_2510);
nor UO_322 (O_322,N_2579,N_2275);
or UO_323 (O_323,N_2992,N_2722);
or UO_324 (O_324,N_2354,N_2433);
and UO_325 (O_325,N_2688,N_2589);
or UO_326 (O_326,N_2374,N_2264);
xor UO_327 (O_327,N_2985,N_2852);
or UO_328 (O_328,N_2463,N_2348);
nor UO_329 (O_329,N_2844,N_2502);
nor UO_330 (O_330,N_2772,N_2650);
nand UO_331 (O_331,N_2315,N_2970);
or UO_332 (O_332,N_2690,N_2274);
nor UO_333 (O_333,N_2911,N_2917);
or UO_334 (O_334,N_2623,N_2778);
and UO_335 (O_335,N_2491,N_2353);
nand UO_336 (O_336,N_2544,N_2317);
nand UO_337 (O_337,N_2883,N_2728);
nand UO_338 (O_338,N_2308,N_2251);
or UO_339 (O_339,N_2307,N_2393);
nor UO_340 (O_340,N_2776,N_2584);
nor UO_341 (O_341,N_2736,N_2518);
nor UO_342 (O_342,N_2834,N_2832);
and UO_343 (O_343,N_2866,N_2285);
nand UO_344 (O_344,N_2862,N_2794);
nor UO_345 (O_345,N_2851,N_2903);
nand UO_346 (O_346,N_2713,N_2338);
nor UO_347 (O_347,N_2922,N_2583);
nor UO_348 (O_348,N_2389,N_2490);
nand UO_349 (O_349,N_2537,N_2908);
nor UO_350 (O_350,N_2438,N_2745);
nor UO_351 (O_351,N_2265,N_2328);
nand UO_352 (O_352,N_2755,N_2725);
nor UO_353 (O_353,N_2474,N_2497);
or UO_354 (O_354,N_2855,N_2384);
nand UO_355 (O_355,N_2806,N_2550);
nor UO_356 (O_356,N_2770,N_2387);
or UO_357 (O_357,N_2395,N_2447);
nor UO_358 (O_358,N_2750,N_2304);
nand UO_359 (O_359,N_2549,N_2657);
and UO_360 (O_360,N_2487,N_2545);
nand UO_361 (O_361,N_2768,N_2955);
nor UO_362 (O_362,N_2266,N_2575);
and UO_363 (O_363,N_2689,N_2740);
nor UO_364 (O_364,N_2481,N_2476);
nor UO_365 (O_365,N_2546,N_2734);
nand UO_366 (O_366,N_2429,N_2590);
and UO_367 (O_367,N_2685,N_2973);
nor UO_368 (O_368,N_2378,N_2558);
nor UO_369 (O_369,N_2613,N_2305);
nand UO_370 (O_370,N_2259,N_2874);
nor UO_371 (O_371,N_2765,N_2960);
and UO_372 (O_372,N_2426,N_2283);
nor UO_373 (O_373,N_2798,N_2634);
nand UO_374 (O_374,N_2492,N_2923);
xnor UO_375 (O_375,N_2927,N_2404);
nand UO_376 (O_376,N_2592,N_2818);
and UO_377 (O_377,N_2748,N_2296);
and UO_378 (O_378,N_2825,N_2912);
and UO_379 (O_379,N_2854,N_2475);
or UO_380 (O_380,N_2838,N_2935);
and UO_381 (O_381,N_2387,N_2821);
nor UO_382 (O_382,N_2523,N_2937);
and UO_383 (O_383,N_2805,N_2996);
nand UO_384 (O_384,N_2259,N_2534);
and UO_385 (O_385,N_2304,N_2839);
nand UO_386 (O_386,N_2280,N_2544);
nor UO_387 (O_387,N_2438,N_2423);
nor UO_388 (O_388,N_2927,N_2444);
nor UO_389 (O_389,N_2416,N_2426);
nand UO_390 (O_390,N_2312,N_2486);
xnor UO_391 (O_391,N_2338,N_2524);
or UO_392 (O_392,N_2483,N_2681);
nand UO_393 (O_393,N_2571,N_2822);
nor UO_394 (O_394,N_2921,N_2459);
and UO_395 (O_395,N_2871,N_2878);
and UO_396 (O_396,N_2902,N_2371);
nor UO_397 (O_397,N_2822,N_2434);
or UO_398 (O_398,N_2360,N_2754);
nand UO_399 (O_399,N_2774,N_2870);
or UO_400 (O_400,N_2737,N_2467);
nand UO_401 (O_401,N_2931,N_2282);
nand UO_402 (O_402,N_2803,N_2507);
nand UO_403 (O_403,N_2251,N_2538);
or UO_404 (O_404,N_2770,N_2967);
nand UO_405 (O_405,N_2402,N_2567);
nand UO_406 (O_406,N_2929,N_2864);
xor UO_407 (O_407,N_2842,N_2391);
and UO_408 (O_408,N_2259,N_2709);
nand UO_409 (O_409,N_2355,N_2330);
nand UO_410 (O_410,N_2626,N_2763);
nand UO_411 (O_411,N_2254,N_2513);
nor UO_412 (O_412,N_2722,N_2422);
nand UO_413 (O_413,N_2439,N_2351);
nor UO_414 (O_414,N_2815,N_2840);
and UO_415 (O_415,N_2593,N_2397);
nor UO_416 (O_416,N_2583,N_2795);
nand UO_417 (O_417,N_2788,N_2961);
or UO_418 (O_418,N_2943,N_2686);
or UO_419 (O_419,N_2682,N_2341);
or UO_420 (O_420,N_2343,N_2715);
nand UO_421 (O_421,N_2305,N_2317);
and UO_422 (O_422,N_2345,N_2359);
or UO_423 (O_423,N_2412,N_2970);
nand UO_424 (O_424,N_2370,N_2734);
and UO_425 (O_425,N_2737,N_2830);
and UO_426 (O_426,N_2577,N_2357);
nor UO_427 (O_427,N_2343,N_2937);
xor UO_428 (O_428,N_2926,N_2317);
nor UO_429 (O_429,N_2723,N_2852);
xnor UO_430 (O_430,N_2483,N_2285);
and UO_431 (O_431,N_2815,N_2616);
nand UO_432 (O_432,N_2975,N_2437);
or UO_433 (O_433,N_2564,N_2412);
and UO_434 (O_434,N_2909,N_2732);
nand UO_435 (O_435,N_2688,N_2530);
nand UO_436 (O_436,N_2587,N_2848);
or UO_437 (O_437,N_2361,N_2541);
and UO_438 (O_438,N_2960,N_2276);
and UO_439 (O_439,N_2261,N_2713);
or UO_440 (O_440,N_2659,N_2811);
or UO_441 (O_441,N_2434,N_2813);
nand UO_442 (O_442,N_2583,N_2756);
or UO_443 (O_443,N_2424,N_2832);
and UO_444 (O_444,N_2738,N_2896);
and UO_445 (O_445,N_2312,N_2334);
nand UO_446 (O_446,N_2460,N_2943);
nand UO_447 (O_447,N_2510,N_2796);
and UO_448 (O_448,N_2954,N_2477);
nand UO_449 (O_449,N_2698,N_2493);
nand UO_450 (O_450,N_2842,N_2928);
nand UO_451 (O_451,N_2264,N_2516);
or UO_452 (O_452,N_2556,N_2885);
nand UO_453 (O_453,N_2322,N_2430);
and UO_454 (O_454,N_2627,N_2881);
nor UO_455 (O_455,N_2880,N_2585);
nor UO_456 (O_456,N_2696,N_2610);
nand UO_457 (O_457,N_2449,N_2593);
or UO_458 (O_458,N_2971,N_2330);
and UO_459 (O_459,N_2600,N_2973);
nor UO_460 (O_460,N_2384,N_2343);
nor UO_461 (O_461,N_2925,N_2472);
nor UO_462 (O_462,N_2870,N_2997);
nor UO_463 (O_463,N_2498,N_2871);
and UO_464 (O_464,N_2904,N_2397);
and UO_465 (O_465,N_2347,N_2484);
and UO_466 (O_466,N_2613,N_2556);
or UO_467 (O_467,N_2921,N_2490);
and UO_468 (O_468,N_2555,N_2590);
or UO_469 (O_469,N_2283,N_2952);
and UO_470 (O_470,N_2547,N_2543);
and UO_471 (O_471,N_2885,N_2947);
and UO_472 (O_472,N_2358,N_2866);
or UO_473 (O_473,N_2916,N_2803);
and UO_474 (O_474,N_2744,N_2661);
and UO_475 (O_475,N_2496,N_2812);
and UO_476 (O_476,N_2282,N_2964);
or UO_477 (O_477,N_2834,N_2798);
nand UO_478 (O_478,N_2367,N_2980);
nor UO_479 (O_479,N_2564,N_2259);
and UO_480 (O_480,N_2900,N_2943);
nand UO_481 (O_481,N_2684,N_2748);
or UO_482 (O_482,N_2497,N_2692);
and UO_483 (O_483,N_2300,N_2604);
nand UO_484 (O_484,N_2554,N_2713);
nor UO_485 (O_485,N_2311,N_2674);
nor UO_486 (O_486,N_2988,N_2663);
and UO_487 (O_487,N_2501,N_2660);
or UO_488 (O_488,N_2680,N_2355);
nor UO_489 (O_489,N_2418,N_2282);
or UO_490 (O_490,N_2733,N_2517);
or UO_491 (O_491,N_2451,N_2690);
or UO_492 (O_492,N_2308,N_2578);
nor UO_493 (O_493,N_2470,N_2490);
or UO_494 (O_494,N_2921,N_2315);
and UO_495 (O_495,N_2436,N_2420);
nand UO_496 (O_496,N_2546,N_2425);
nand UO_497 (O_497,N_2782,N_2533);
and UO_498 (O_498,N_2896,N_2811);
nor UO_499 (O_499,N_2742,N_2299);
endmodule